module basic_5000_50000_5000_20_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
or U0 (N_0,In_1400,In_4752);
nand U1 (N_1,In_1414,In_4179);
or U2 (N_2,In_869,In_786);
nand U3 (N_3,In_2773,In_3613);
or U4 (N_4,In_1143,In_2358);
and U5 (N_5,In_934,In_4566);
nor U6 (N_6,In_3776,In_3556);
or U7 (N_7,In_2083,In_1033);
or U8 (N_8,In_885,In_1191);
or U9 (N_9,In_3649,In_2486);
nand U10 (N_10,In_1607,In_4280);
nor U11 (N_11,In_873,In_1966);
nand U12 (N_12,In_2745,In_3742);
xor U13 (N_13,In_4596,In_2011);
nand U14 (N_14,In_4562,In_3234);
or U15 (N_15,In_2638,In_1235);
and U16 (N_16,In_402,In_4711);
or U17 (N_17,In_1226,In_2265);
and U18 (N_18,In_3303,In_4198);
or U19 (N_19,In_3521,In_1327);
nor U20 (N_20,In_2619,In_615);
xor U21 (N_21,In_3171,In_4834);
nand U22 (N_22,In_2002,In_4404);
and U23 (N_23,In_2976,In_2445);
xnor U24 (N_24,In_3843,In_4082);
nand U25 (N_25,In_602,In_1670);
nand U26 (N_26,In_166,In_1647);
and U27 (N_27,In_1778,In_1812);
nor U28 (N_28,In_1409,In_3162);
and U29 (N_29,In_824,In_4126);
and U30 (N_30,In_3474,In_2565);
or U31 (N_31,In_1082,In_3980);
xor U32 (N_32,In_266,In_2668);
nand U33 (N_33,In_4309,In_1365);
or U34 (N_34,In_4700,In_2596);
nand U35 (N_35,In_3021,In_1458);
and U36 (N_36,In_3037,In_2851);
nand U37 (N_37,In_3667,In_812);
and U38 (N_38,In_174,In_2622);
nand U39 (N_39,In_2310,In_2537);
and U40 (N_40,In_4153,In_707);
nor U41 (N_41,In_4761,In_3284);
or U42 (N_42,In_1796,In_1698);
nor U43 (N_43,In_2014,In_2664);
or U44 (N_44,In_3460,In_3764);
and U45 (N_45,In_4419,In_1988);
nor U46 (N_46,In_1002,In_2231);
or U47 (N_47,In_4502,In_234);
nand U48 (N_48,In_4889,In_4478);
and U49 (N_49,In_2730,In_3866);
nand U50 (N_50,In_208,In_1364);
or U51 (N_51,In_881,In_3782);
and U52 (N_52,In_4799,In_4918);
or U53 (N_53,In_3401,In_1861);
nor U54 (N_54,In_4655,In_3051);
xnor U55 (N_55,In_4910,In_250);
xnor U56 (N_56,In_3040,In_2292);
nor U57 (N_57,In_2325,In_1029);
or U58 (N_58,In_4358,In_2914);
nand U59 (N_59,In_1528,In_678);
or U60 (N_60,In_541,In_281);
and U61 (N_61,In_159,In_1920);
or U62 (N_62,In_4985,In_1381);
and U63 (N_63,In_341,In_2617);
xnor U64 (N_64,In_3376,In_4218);
or U65 (N_65,In_2508,In_4828);
and U66 (N_66,In_474,In_1268);
nor U67 (N_67,In_2170,In_1883);
nor U68 (N_68,In_72,In_1087);
nand U69 (N_69,In_3741,In_682);
nand U70 (N_70,In_1467,In_4697);
or U71 (N_71,In_4789,In_116);
or U72 (N_72,In_2413,In_3330);
nand U73 (N_73,In_2400,In_4021);
and U74 (N_74,In_1114,In_1272);
nand U75 (N_75,In_2359,In_3525);
nand U76 (N_76,In_2718,In_4670);
nand U77 (N_77,In_332,In_1009);
nand U78 (N_78,In_2320,In_3043);
nand U79 (N_79,In_3213,In_514);
and U80 (N_80,In_1166,In_2236);
and U81 (N_81,In_105,In_4663);
nor U82 (N_82,In_3186,In_4110);
nor U83 (N_83,In_721,In_2516);
and U84 (N_84,In_4346,In_3981);
and U85 (N_85,In_4227,In_4602);
nand U86 (N_86,In_2812,In_3937);
and U87 (N_87,In_2651,In_152);
or U88 (N_88,In_388,In_2807);
xor U89 (N_89,In_4657,In_2691);
nor U90 (N_90,In_333,In_739);
or U91 (N_91,In_2174,In_3624);
xor U92 (N_92,In_1708,In_2841);
and U93 (N_93,In_3299,In_1070);
nand U94 (N_94,In_3635,In_1950);
or U95 (N_95,In_4557,In_2101);
nand U96 (N_96,In_4010,In_4105);
or U97 (N_97,In_2996,In_692);
nand U98 (N_98,In_3932,In_817);
nand U99 (N_99,In_417,In_3489);
or U100 (N_100,In_3601,In_3096);
nor U101 (N_101,In_804,In_2346);
and U102 (N_102,In_4539,In_4268);
nand U103 (N_103,In_3503,In_3222);
xor U104 (N_104,In_4061,In_949);
xnor U105 (N_105,In_1839,In_297);
nor U106 (N_106,In_3602,In_241);
and U107 (N_107,In_3699,In_4031);
nand U108 (N_108,In_4890,In_489);
nor U109 (N_109,In_3951,In_3267);
nor U110 (N_110,In_227,In_238);
nor U111 (N_111,In_3344,In_733);
and U112 (N_112,In_4730,In_289);
nand U113 (N_113,In_4076,In_2015);
and U114 (N_114,In_1225,In_1693);
or U115 (N_115,In_2327,In_114);
and U116 (N_116,In_716,In_1739);
and U117 (N_117,In_4635,In_1896);
nand U118 (N_118,In_3967,In_2073);
nand U119 (N_119,In_932,In_1462);
or U120 (N_120,In_3101,In_981);
nand U121 (N_121,In_565,In_4555);
and U122 (N_122,In_1313,In_4331);
and U123 (N_123,In_625,In_2629);
and U124 (N_124,In_1517,In_2487);
nor U125 (N_125,In_4277,In_1628);
and U126 (N_126,In_39,In_4286);
or U127 (N_127,In_3872,In_2465);
xor U128 (N_128,In_2641,In_2951);
nand U129 (N_129,In_4270,In_419);
nand U130 (N_130,In_4454,In_3170);
or U131 (N_131,In_3459,In_4780);
nand U132 (N_132,In_1952,In_3355);
or U133 (N_133,In_836,In_3530);
and U134 (N_134,In_4293,In_1566);
or U135 (N_135,In_2012,In_3318);
and U136 (N_136,In_3024,In_4666);
and U137 (N_137,In_4370,In_2770);
or U138 (N_138,In_920,In_4222);
nand U139 (N_139,In_2262,In_1475);
nor U140 (N_140,In_179,In_1445);
nand U141 (N_141,In_4690,In_2823);
nor U142 (N_142,In_3528,In_2441);
nand U143 (N_143,In_2125,In_4023);
nand U144 (N_144,In_1489,In_4677);
and U145 (N_145,In_665,In_2559);
nor U146 (N_146,In_2450,In_3871);
nor U147 (N_147,In_2683,In_1250);
nor U148 (N_148,In_638,In_2515);
and U149 (N_149,In_3666,In_1092);
xnor U150 (N_150,In_3368,In_2482);
and U151 (N_151,In_3902,In_4119);
or U152 (N_152,In_2047,In_4745);
nor U153 (N_153,In_3978,In_4742);
or U154 (N_154,In_4764,In_3288);
or U155 (N_155,In_841,In_717);
nand U156 (N_156,In_584,In_2543);
or U157 (N_157,In_3326,In_2068);
and U158 (N_158,In_3795,In_2222);
nor U159 (N_159,In_1416,In_2825);
or U160 (N_160,In_131,In_77);
nand U161 (N_161,In_1339,In_2023);
and U162 (N_162,In_4702,In_1869);
nand U163 (N_163,In_137,In_3590);
xnor U164 (N_164,In_3559,In_3461);
and U165 (N_165,In_979,In_342);
nor U166 (N_166,In_4759,In_4913);
and U167 (N_167,In_3033,In_2127);
and U168 (N_168,In_446,In_3845);
nand U169 (N_169,In_411,In_1929);
and U170 (N_170,In_2200,In_1316);
or U171 (N_171,In_1319,In_2977);
and U172 (N_172,In_4005,In_936);
and U173 (N_173,In_3069,In_761);
nand U174 (N_174,In_1755,In_2250);
xor U175 (N_175,In_1591,In_2892);
and U176 (N_176,In_391,In_783);
nor U177 (N_177,In_394,In_3571);
or U178 (N_178,In_2544,In_4960);
or U179 (N_179,In_3897,In_1516);
or U180 (N_180,In_3523,In_3511);
nor U181 (N_181,In_157,In_1654);
or U182 (N_182,In_3061,In_1027);
and U183 (N_183,In_206,In_3723);
and U184 (N_184,In_4998,In_1435);
and U185 (N_185,In_3923,In_2332);
nor U186 (N_186,In_882,In_4518);
xnor U187 (N_187,In_1592,In_4819);
nand U188 (N_188,In_4736,In_2150);
nand U189 (N_189,In_57,In_654);
and U190 (N_190,In_1903,In_4751);
nor U191 (N_191,In_273,In_1613);
and U192 (N_192,In_4115,In_2653);
or U193 (N_193,In_4907,In_4902);
nor U194 (N_194,In_1137,In_4640);
or U195 (N_195,In_543,In_1997);
nand U196 (N_196,In_3930,In_1404);
and U197 (N_197,In_922,In_2789);
xor U198 (N_198,In_4289,In_1476);
nand U199 (N_199,In_2353,In_987);
xor U200 (N_200,In_2046,In_2104);
and U201 (N_201,In_4629,In_302);
xnor U202 (N_202,In_1408,In_3931);
or U203 (N_203,In_4449,In_4909);
xnor U204 (N_204,In_233,In_2240);
xor U205 (N_205,In_23,In_2258);
or U206 (N_206,In_2178,In_1504);
nand U207 (N_207,In_4090,In_2633);
nand U208 (N_208,In_2331,In_4870);
and U209 (N_209,In_343,In_754);
nor U210 (N_210,In_2452,In_2685);
or U211 (N_211,In_1793,In_4287);
or U212 (N_212,In_3516,In_3022);
and U213 (N_213,In_280,In_4937);
or U214 (N_214,In_1512,In_1285);
nor U215 (N_215,In_4425,In_4647);
nor U216 (N_216,In_532,In_3589);
nand U217 (N_217,In_620,In_3811);
and U218 (N_218,In_3560,In_1434);
and U219 (N_219,In_3997,In_559);
or U220 (N_220,In_570,In_3088);
nand U221 (N_221,In_473,In_1620);
and U222 (N_222,In_1090,In_4573);
and U223 (N_223,In_2409,In_1681);
and U224 (N_224,In_3837,In_3491);
nor U225 (N_225,In_2848,In_915);
or U226 (N_226,In_677,In_1301);
and U227 (N_227,In_4450,In_1579);
or U228 (N_228,In_1483,In_4209);
nand U229 (N_229,In_2733,In_1065);
or U230 (N_230,In_4788,In_2710);
or U231 (N_231,In_3786,In_4698);
and U232 (N_232,In_4935,In_1139);
nand U233 (N_233,In_3893,In_4163);
nor U234 (N_234,In_1849,In_1535);
nand U235 (N_235,In_307,In_3928);
and U236 (N_236,In_606,In_1234);
xnor U237 (N_237,In_2177,In_2172);
nor U238 (N_238,In_1610,In_4324);
nand U239 (N_239,In_4371,In_2202);
nand U240 (N_240,In_4773,In_2899);
xnor U241 (N_241,In_2102,In_1303);
nand U242 (N_242,In_3966,In_2118);
and U243 (N_243,In_3298,In_3456);
nand U244 (N_244,In_1072,In_2189);
or U245 (N_245,In_848,In_3844);
xnor U246 (N_246,In_1187,In_2579);
xor U247 (N_247,In_912,In_4213);
xor U248 (N_248,In_1843,In_2521);
or U249 (N_249,In_2898,In_1656);
or U250 (N_250,In_2694,In_4822);
nor U251 (N_251,In_4554,In_4678);
or U252 (N_252,In_1405,In_1376);
or U253 (N_253,In_1937,In_2490);
and U254 (N_254,In_1100,In_2643);
nand U255 (N_255,In_2607,In_1372);
and U256 (N_256,In_40,In_3550);
nor U257 (N_257,In_4888,In_2035);
nor U258 (N_258,In_210,In_2690);
and U259 (N_259,In_3373,In_4028);
and U260 (N_260,In_994,In_2436);
or U261 (N_261,In_1133,In_2786);
xor U262 (N_262,In_2473,In_47);
nor U263 (N_263,In_3004,In_839);
nor U264 (N_264,In_2693,In_2798);
nand U265 (N_265,In_4569,In_1519);
xnor U266 (N_266,In_4359,In_4380);
or U267 (N_267,In_4336,In_62);
nor U268 (N_268,In_4093,In_2944);
nor U269 (N_269,In_3304,In_765);
and U270 (N_270,In_697,In_1769);
nand U271 (N_271,In_197,In_3791);
or U272 (N_272,In_4187,In_199);
nor U273 (N_273,In_1291,In_3706);
or U274 (N_274,In_4460,In_3231);
nand U275 (N_275,In_2553,In_4703);
nand U276 (N_276,In_464,In_3755);
and U277 (N_277,In_884,In_2484);
nand U278 (N_278,In_4169,In_1794);
or U279 (N_279,In_2961,In_535);
and U280 (N_280,In_907,In_712);
nor U281 (N_281,In_1692,In_1190);
and U282 (N_282,In_3569,In_1240);
or U283 (N_283,In_924,In_4691);
and U284 (N_284,In_3245,In_3858);
and U285 (N_285,In_224,In_1706);
or U286 (N_286,In_4236,In_2679);
nor U287 (N_287,In_4113,In_2984);
nor U288 (N_288,In_4248,In_3718);
or U289 (N_289,In_3011,In_547);
nor U290 (N_290,In_549,In_2119);
nor U291 (N_291,In_1587,In_601);
nand U292 (N_292,In_3434,In_4130);
nand U293 (N_293,In_779,In_3232);
nand U294 (N_294,In_878,In_3929);
nand U295 (N_295,In_310,In_3953);
nor U296 (N_296,In_3309,In_1375);
or U297 (N_297,In_3240,In_4149);
nor U298 (N_298,In_3263,In_594);
nor U299 (N_299,In_4241,In_4284);
and U300 (N_300,In_2031,In_926);
and U301 (N_301,In_1182,In_4796);
or U302 (N_302,In_1781,In_701);
nor U303 (N_303,In_1927,In_3541);
or U304 (N_304,In_168,In_4531);
or U305 (N_305,In_3974,In_3348);
nor U306 (N_306,In_1423,In_1600);
nor U307 (N_307,In_2759,In_1720);
nor U308 (N_308,In_416,In_4977);
nor U309 (N_309,In_4710,In_1465);
nand U310 (N_310,In_3448,In_1917);
nand U311 (N_311,In_4795,In_1678);
nand U312 (N_312,In_3283,In_2243);
xnor U313 (N_313,In_1411,In_1129);
nand U314 (N_314,In_1695,In_916);
xor U315 (N_315,In_4081,In_708);
xor U316 (N_316,In_1771,In_3797);
xnor U317 (N_317,In_1179,In_4911);
and U318 (N_318,In_4856,In_1370);
nand U319 (N_319,In_143,In_4122);
xor U320 (N_320,In_3195,In_2655);
nand U321 (N_321,In_4212,In_1797);
or U322 (N_322,In_1851,In_1683);
and U323 (N_323,In_1184,In_674);
nand U324 (N_324,In_3696,In_1766);
nor U325 (N_325,In_348,In_4194);
nor U326 (N_326,In_3307,In_3411);
xor U327 (N_327,In_65,In_2220);
nand U328 (N_328,In_1563,In_4835);
nand U329 (N_329,In_4316,In_423);
nand U330 (N_330,In_3948,In_2018);
nand U331 (N_331,In_1792,In_3243);
and U332 (N_332,In_3806,In_3648);
nor U333 (N_333,In_1152,In_4747);
nor U334 (N_334,In_367,In_144);
and U335 (N_335,In_3996,In_2697);
nand U336 (N_336,In_1762,In_4995);
nand U337 (N_337,In_316,In_640);
or U338 (N_338,In_583,In_2030);
and U339 (N_339,In_3581,In_4534);
or U340 (N_340,In_436,In_4551);
nand U341 (N_341,In_2025,In_2080);
and U342 (N_342,In_509,In_2362);
or U343 (N_343,In_2645,In_4932);
or U344 (N_344,In_1562,In_4161);
or U345 (N_345,In_123,In_3862);
nor U346 (N_346,In_218,In_1650);
xnor U347 (N_347,In_980,In_1258);
nor U348 (N_348,In_4510,In_3869);
nor U349 (N_349,In_1197,In_1264);
or U350 (N_350,In_578,In_3018);
and U351 (N_351,In_389,In_1325);
and U352 (N_352,In_1457,In_1975);
or U353 (N_353,In_2614,In_1889);
and U354 (N_354,In_2714,In_2322);
nor U355 (N_355,In_753,In_3356);
and U356 (N_356,In_2042,In_792);
and U357 (N_357,In_854,In_3479);
nor U358 (N_358,In_827,In_2161);
nand U359 (N_359,In_4444,In_4857);
or U360 (N_360,In_4642,In_4512);
nand U361 (N_361,In_3744,In_2197);
nand U362 (N_362,In_2503,In_4345);
or U363 (N_363,In_3224,In_3017);
nand U364 (N_364,In_4625,In_2952);
nand U365 (N_365,In_2999,In_4592);
nand U366 (N_366,In_3264,In_3072);
or U367 (N_367,In_2903,In_1761);
or U368 (N_368,In_3239,In_3286);
nor U369 (N_369,In_4471,In_381);
and U370 (N_370,In_3384,In_2425);
or U371 (N_371,In_2299,In_471);
or U372 (N_372,In_2540,In_3086);
and U373 (N_373,In_1902,In_1568);
or U374 (N_374,In_4522,In_3357);
and U375 (N_375,In_1799,In_132);
and U376 (N_376,In_2779,In_1312);
nand U377 (N_377,In_510,In_2483);
nor U378 (N_378,In_3695,In_748);
and U379 (N_379,In_2107,In_3672);
nand U380 (N_380,In_4463,In_229);
nand U381 (N_381,In_1394,In_4328);
xor U382 (N_382,In_1964,In_2708);
and U383 (N_383,In_2148,In_1593);
xnor U384 (N_384,In_3056,In_37);
nand U385 (N_385,In_736,In_3962);
nor U386 (N_386,In_619,In_965);
or U387 (N_387,In_1056,In_862);
nor U388 (N_388,In_866,In_758);
and U389 (N_389,In_2621,In_2140);
xor U390 (N_390,In_3913,In_2138);
nor U391 (N_391,In_2504,In_2344);
or U392 (N_392,In_3241,In_3562);
nand U393 (N_393,In_87,In_1582);
nand U394 (N_394,In_3629,In_3810);
nor U395 (N_395,In_2582,In_3547);
or U396 (N_396,In_2975,In_4542);
or U397 (N_397,In_2211,In_4563);
nand U398 (N_398,In_31,In_2306);
or U399 (N_399,In_1944,In_4473);
nor U400 (N_400,In_2378,In_1709);
and U401 (N_401,In_49,In_2455);
nor U402 (N_402,In_3366,In_4296);
or U403 (N_403,In_1636,In_4408);
and U404 (N_404,In_1001,In_63);
nand U405 (N_405,In_282,In_3181);
nor U406 (N_406,In_3106,In_515);
nor U407 (N_407,In_3099,In_990);
nor U408 (N_408,In_3508,In_1117);
nand U409 (N_409,In_2356,In_4996);
nand U410 (N_410,In_2809,In_4385);
and U411 (N_411,In_34,In_400);
and U412 (N_412,In_2744,In_3394);
nand U413 (N_413,In_1945,In_1806);
or U414 (N_414,In_3614,In_2853);
or U415 (N_415,In_1862,In_1501);
nor U416 (N_416,In_486,In_3148);
nand U417 (N_417,In_3487,In_25);
nor U418 (N_418,In_3204,In_806);
nand U419 (N_419,In_579,In_1808);
and U420 (N_420,In_3596,In_1222);
nand U421 (N_421,In_2769,In_2282);
and U422 (N_422,In_2982,In_1120);
or U423 (N_423,In_2933,In_3007);
nor U424 (N_424,In_4208,In_4981);
and U425 (N_425,In_67,In_1688);
nor U426 (N_426,In_3256,In_3704);
nand U427 (N_427,In_1042,In_3471);
nor U428 (N_428,In_3398,In_913);
and U429 (N_429,In_590,In_481);
xor U430 (N_430,In_1208,In_1942);
nand U431 (N_431,In_2758,In_978);
nand U432 (N_432,In_2647,In_3372);
nand U433 (N_433,In_1194,In_3345);
or U434 (N_434,In_585,In_2603);
nor U435 (N_435,In_6,In_4094);
xnor U436 (N_436,In_4181,In_4574);
nor U437 (N_437,In_15,In_2735);
and U438 (N_438,In_997,In_731);
and U439 (N_439,In_3203,In_562);
or U440 (N_440,In_2350,In_322);
nand U441 (N_441,In_2334,In_3655);
or U442 (N_442,In_4481,In_2144);
and U443 (N_443,In_4606,In_3042);
nand U444 (N_444,In_4442,In_1289);
or U445 (N_445,In_1311,In_4599);
nand U446 (N_446,In_4260,In_58);
nand U447 (N_447,In_2339,In_4047);
or U448 (N_448,In_3029,In_2044);
xor U449 (N_449,In_1022,In_4254);
nand U450 (N_450,In_1478,In_891);
or U451 (N_451,In_1764,In_2987);
xor U452 (N_452,In_2757,In_657);
nor U453 (N_453,In_2936,In_1716);
and U454 (N_454,In_796,In_1488);
xnor U455 (N_455,In_4214,In_3818);
or U456 (N_456,In_3475,In_2437);
or U457 (N_457,In_3733,In_1233);
or U458 (N_458,In_3690,In_2203);
or U459 (N_459,In_4224,In_3386);
nand U460 (N_460,In_3936,In_1112);
nand U461 (N_461,In_749,In_3408);
nor U462 (N_462,In_467,In_4527);
or U463 (N_463,In_893,In_1844);
xnor U464 (N_464,In_204,In_3594);
nor U465 (N_465,In_4836,In_3293);
and U466 (N_466,In_1094,In_3658);
and U467 (N_467,In_2646,In_1733);
or U468 (N_468,In_911,In_3611);
nand U469 (N_469,In_2439,In_633);
nand U470 (N_470,In_1368,In_3631);
nand U471 (N_471,In_3746,In_3289);
or U472 (N_472,In_3127,In_376);
nand U473 (N_473,In_1443,In_2372);
and U474 (N_474,In_1605,In_1686);
xor U475 (N_475,In_954,In_3592);
nor U476 (N_476,In_1257,In_230);
nand U477 (N_477,In_4660,In_1557);
and U478 (N_478,In_4168,In_768);
nand U479 (N_479,In_598,In_2700);
and U480 (N_480,In_1432,In_2003);
nor U481 (N_481,In_3202,In_3053);
nand U482 (N_482,In_203,In_2884);
nor U483 (N_483,In_4680,In_1899);
nor U484 (N_484,In_2205,In_961);
or U485 (N_485,In_781,In_3393);
nor U486 (N_486,In_71,In_1985);
nor U487 (N_487,In_1253,In_718);
or U488 (N_488,In_219,In_1564);
and U489 (N_489,In_4968,In_4276);
or U490 (N_490,In_751,In_3992);
or U491 (N_491,In_1221,In_867);
nand U492 (N_492,In_1900,In_3643);
or U493 (N_493,In_4128,In_3850);
and U494 (N_494,In_4687,In_2591);
or U495 (N_495,In_3796,In_3616);
nor U496 (N_496,In_2624,In_2348);
nor U497 (N_497,In_3917,In_3675);
xnor U498 (N_498,In_2052,In_2935);
and U499 (N_499,In_3295,In_277);
or U500 (N_500,In_3767,In_3312);
and U501 (N_501,In_4084,In_3549);
and U502 (N_502,In_2592,In_3431);
nand U503 (N_503,In_253,In_647);
or U504 (N_504,In_2326,In_1657);
xor U505 (N_505,In_1615,In_399);
nand U506 (N_506,In_4210,In_843);
nand U507 (N_507,In_1943,In_4386);
nor U508 (N_508,In_3066,In_2709);
nor U509 (N_509,In_304,In_1324);
nor U510 (N_510,In_4616,In_1050);
or U511 (N_511,In_1047,In_1992);
nor U512 (N_512,In_1509,In_4390);
and U513 (N_513,In_3082,In_102);
and U514 (N_514,In_2010,In_4022);
and U515 (N_515,In_860,In_3821);
or U516 (N_516,In_641,In_566);
xor U517 (N_517,In_3340,In_3065);
or U518 (N_518,In_1081,In_1697);
and U519 (N_519,In_596,In_4922);
and U520 (N_520,In_4714,In_1876);
and U521 (N_521,In_1634,In_1891);
nor U522 (N_522,In_4252,In_2844);
xor U523 (N_523,In_687,In_4457);
nor U524 (N_524,In_2630,In_2576);
and U525 (N_525,In_3349,In_4676);
nand U526 (N_526,In_4431,In_1779);
and U527 (N_527,In_1121,In_2501);
nor U528 (N_528,In_995,In_4145);
or U529 (N_529,In_3711,In_4921);
or U530 (N_530,In_3462,In_354);
and U531 (N_531,In_4133,In_2678);
nor U532 (N_532,In_1842,In_1663);
and U533 (N_533,In_2587,In_1848);
nand U534 (N_534,In_1960,In_1506);
or U535 (N_535,In_1266,In_4903);
or U536 (N_536,In_4188,In_228);
xor U537 (N_537,In_1346,In_4991);
or U538 (N_538,In_2520,In_93);
and U539 (N_539,In_3023,In_191);
nor U540 (N_540,In_265,In_1469);
or U541 (N_541,In_3944,In_760);
nor U542 (N_542,In_4412,In_3450);
nor U543 (N_543,In_1884,In_729);
or U544 (N_544,In_3276,In_430);
nand U545 (N_545,In_1986,In_4125);
nor U546 (N_546,In_3333,In_2388);
nand U547 (N_547,In_1459,In_499);
and U548 (N_548,In_3313,In_1356);
or U549 (N_549,In_1719,In_4339);
nor U550 (N_550,In_2474,In_1284);
or U551 (N_551,In_3421,In_18);
nor U552 (N_552,In_1712,In_4173);
nor U553 (N_553,In_3009,In_2931);
xor U554 (N_554,In_1213,In_1347);
and U555 (N_555,In_2418,In_931);
nor U556 (N_556,In_1480,In_426);
xor U557 (N_557,In_3465,In_2731);
nor U558 (N_558,In_2857,In_1086);
nor U559 (N_559,In_1643,In_368);
nand U560 (N_560,In_2832,In_209);
or U561 (N_561,In_3734,In_616);
and U562 (N_562,In_4217,In_967);
or U563 (N_563,In_4826,In_4150);
nand U564 (N_564,In_3308,In_3527);
and U565 (N_565,In_4556,In_1109);
or U566 (N_566,In_2865,In_1215);
xor U567 (N_567,In_4776,In_4954);
or U568 (N_568,In_2666,In_3453);
xor U569 (N_569,In_1714,In_2658);
or U570 (N_570,In_2,In_2212);
and U571 (N_571,In_3275,In_3046);
nor U572 (N_572,In_1660,In_4244);
nand U573 (N_573,In_3605,In_1829);
xnor U574 (N_574,In_4801,In_3196);
nand U575 (N_575,In_3422,In_2065);
nor U576 (N_576,In_2640,In_3777);
xnor U577 (N_577,In_3970,In_4480);
and U578 (N_578,In_3972,In_1870);
or U579 (N_579,In_4278,In_895);
nor U580 (N_580,In_2095,In_2434);
or U581 (N_581,In_2882,In_1192);
and U582 (N_582,In_4233,In_3404);
nor U583 (N_583,In_4701,In_3663);
nand U584 (N_584,In_148,In_3364);
and U585 (N_585,In_4343,In_1507);
or U586 (N_586,In_1809,In_3680);
or U587 (N_587,In_3246,In_653);
nor U588 (N_588,In_257,In_4536);
xor U589 (N_589,In_2981,In_2985);
and U590 (N_590,In_4504,In_2235);
xor U591 (N_591,In_1659,In_1773);
nand U592 (N_592,In_2878,In_3747);
or U593 (N_593,In_4853,In_1314);
and U594 (N_594,In_2005,In_2242);
or U595 (N_595,In_3573,In_800);
xnor U596 (N_596,In_3801,In_4506);
nor U597 (N_597,In_2826,In_1957);
xor U598 (N_598,In_4413,In_4477);
nor U599 (N_599,In_2616,In_418);
or U600 (N_600,In_2625,In_2365);
nand U601 (N_601,In_4770,In_3143);
nor U602 (N_602,In_943,In_1401);
nor U603 (N_603,In_1689,In_679);
or U604 (N_604,In_1456,In_1503);
nor U605 (N_605,In_4528,In_2160);
and U606 (N_606,In_244,In_4059);
xnor U607 (N_607,In_2433,In_2573);
and U608 (N_608,In_1188,In_637);
xnor U609 (N_609,In_2020,In_3785);
or U610 (N_610,In_1419,In_1163);
xnor U611 (N_611,In_4892,In_4124);
or U612 (N_612,In_3568,In_276);
nand U613 (N_613,In_3827,In_2995);
nand U614 (N_614,In_2476,In_1195);
nand U615 (N_615,In_2054,In_1293);
nand U616 (N_616,In_4177,In_1262);
nand U617 (N_617,In_4900,In_4581);
nand U618 (N_618,In_90,In_4447);
or U619 (N_619,In_4709,In_3807);
or U620 (N_620,In_531,In_3381);
and U621 (N_621,In_4235,In_4391);
nand U622 (N_622,In_4987,In_3738);
nor U623 (N_623,In_2067,In_1451);
nor U624 (N_624,In_2671,In_1795);
nand U625 (N_625,In_347,In_2239);
and U626 (N_626,In_3494,In_3351);
and U627 (N_627,In_2371,In_516);
nor U628 (N_628,In_1933,In_3038);
nand U629 (N_629,In_2017,In_3273);
nand U630 (N_630,In_198,In_3708);
nand U631 (N_631,In_4044,In_2960);
and U632 (N_632,In_842,In_4230);
or U633 (N_633,In_2147,In_2780);
or U634 (N_634,In_1069,In_4135);
nand U635 (N_635,In_456,In_4334);
nand U636 (N_636,In_3211,In_3419);
nand U637 (N_637,In_852,In_2373);
xnor U638 (N_638,In_2489,In_4199);
nor U639 (N_639,In_763,In_3155);
or U640 (N_640,In_2257,In_84);
or U641 (N_641,In_1136,In_495);
and U642 (N_642,In_4665,In_2957);
nand U643 (N_643,In_974,In_3780);
nor U644 (N_644,In_1583,In_1846);
nor U645 (N_645,In_4971,In_4855);
and U646 (N_646,In_1460,In_1334);
and U647 (N_647,In_4843,In_4410);
xor U648 (N_648,In_4558,In_4363);
nand U649 (N_649,In_1132,In_4852);
and U650 (N_650,In_4429,In_2156);
and U651 (N_651,In_1836,In_3399);
or U652 (N_652,In_540,In_2923);
and U653 (N_653,In_984,In_3320);
and U654 (N_654,In_80,In_2469);
nor U655 (N_655,In_4096,In_735);
nor U656 (N_656,In_1127,In_4317);
and U657 (N_657,In_2777,In_4840);
or U658 (N_658,In_668,In_1546);
nand U659 (N_659,In_2586,In_1544);
or U660 (N_660,In_1156,In_2386);
xor U661 (N_661,In_3792,In_3693);
or U662 (N_662,In_2082,In_948);
and U663 (N_663,In_1329,In_1296);
nand U664 (N_664,In_3646,In_4899);
or U665 (N_665,In_4601,In_4785);
or U666 (N_666,In_4548,In_1831);
or U667 (N_667,In_4139,In_1525);
nor U668 (N_668,In_4018,In_2391);
nand U669 (N_669,In_3910,In_3522);
or U670 (N_670,In_21,In_2990);
nor U671 (N_671,In_4766,In_194);
nand U672 (N_672,In_462,In_2268);
and U673 (N_673,In_1307,In_2091);
and U674 (N_674,In_4654,In_1998);
nor U675 (N_675,In_1020,In_2430);
nor U676 (N_676,In_2803,In_3977);
nand U677 (N_677,In_81,In_1396);
and U678 (N_678,In_1270,In_2699);
and U679 (N_679,In_2126,In_3277);
or U680 (N_680,In_1996,In_905);
nor U681 (N_681,In_1177,In_2379);
or U682 (N_682,In_528,In_556);
and U683 (N_683,In_4962,In_929);
xnor U684 (N_684,In_651,In_3337);
nand U685 (N_685,In_3414,In_909);
nand U686 (N_686,In_2897,In_1826);
nor U687 (N_687,In_1015,In_374);
nor U688 (N_688,In_4472,In_573);
nand U689 (N_689,In_1865,In_46);
nor U690 (N_690,In_1918,In_3689);
nor U691 (N_691,In_3079,In_1577);
xnor U692 (N_692,In_1425,In_1789);
nand U693 (N_693,In_2535,In_3692);
and U694 (N_694,In_3716,In_870);
and U695 (N_695,In_1118,In_3638);
nand U696 (N_696,In_2871,In_3174);
xor U697 (N_697,In_303,In_623);
or U698 (N_698,In_3617,In_4228);
or U699 (N_699,In_3221,In_2263);
nor U700 (N_700,In_3758,In_3583);
nand U701 (N_701,In_207,In_4451);
xor U702 (N_702,In_4393,In_167);
nor U703 (N_703,In_180,In_3242);
nand U704 (N_704,In_656,In_947);
nor U705 (N_705,In_140,In_1248);
xnor U706 (N_706,In_2776,In_4737);
or U707 (N_707,In_4403,In_567);
nand U708 (N_708,In_4781,In_3405);
nand U709 (N_709,In_3950,In_683);
nor U710 (N_710,In_4992,In_3301);
nand U711 (N_711,In_3443,In_3396);
and U712 (N_712,In_54,In_42);
xnor U713 (N_713,In_4823,In_4347);
or U714 (N_714,In_3451,In_4330);
or U715 (N_715,In_4643,In_4099);
nand U716 (N_716,In_164,In_2836);
and U717 (N_717,In_1338,In_1130);
or U718 (N_718,In_1386,In_4906);
nand U719 (N_719,In_3940,In_1422);
or U720 (N_720,In_618,In_2650);
nor U721 (N_721,In_1841,In_2142);
and U722 (N_722,In_2554,In_4738);
xor U723 (N_723,In_3620,In_921);
nand U724 (N_724,In_3724,In_3270);
nand U725 (N_725,In_2447,In_2928);
nand U726 (N_726,In_334,In_3316);
nand U727 (N_727,In_437,In_1742);
or U728 (N_728,In_92,In_3178);
and U729 (N_729,In_4067,In_1915);
nor U730 (N_730,In_849,In_4846);
nand U731 (N_731,In_4934,In_4553);
nand U732 (N_732,In_1271,In_434);
or U733 (N_733,In_314,In_1010);
or U734 (N_734,In_3003,In_4580);
nor U735 (N_735,In_4174,In_1013);
or U736 (N_736,In_2711,In_1625);
and U737 (N_737,In_414,In_1110);
or U738 (N_738,In_553,In_2532);
and U739 (N_739,In_1594,In_2600);
nor U740 (N_740,In_4607,In_4636);
or U741 (N_741,In_447,In_2249);
nor U742 (N_742,In_136,In_3934);
and U743 (N_743,In_4318,In_529);
nand U744 (N_744,In_3714,In_2390);
and U745 (N_745,In_3314,In_1025);
nand U746 (N_746,In_3577,In_4498);
or U747 (N_747,In_497,In_4790);
nand U748 (N_748,In_985,In_4052);
nor U749 (N_749,In_3370,In_3389);
nand U750 (N_750,In_4017,In_1323);
and U751 (N_751,In_4279,In_172);
or U752 (N_752,In_1749,In_4321);
nor U753 (N_753,In_288,In_362);
nor U754 (N_754,In_3452,In_1180);
nor U755 (N_755,In_1154,In_3325);
nor U756 (N_756,In_3062,In_13);
nand U757 (N_757,In_1857,In_433);
nor U758 (N_758,In_4668,In_2915);
or U759 (N_759,In_4196,In_756);
and U760 (N_760,In_287,In_346);
and U761 (N_761,In_3563,In_2198);
or U762 (N_762,In_3493,In_3788);
nand U763 (N_763,In_3676,In_178);
nand U764 (N_764,In_4627,In_511);
nand U765 (N_765,In_3365,In_538);
nor U766 (N_766,In_2120,In_2087);
nand U767 (N_767,In_3469,In_1649);
nor U768 (N_768,In_2224,In_664);
or U769 (N_769,In_3383,In_1715);
nand U770 (N_770,In_2460,In_1178);
nand U771 (N_771,In_4863,In_3026);
or U772 (N_772,In_2111,In_880);
and U773 (N_773,In_2669,In_501);
or U774 (N_774,In_2191,In_291);
nor U775 (N_775,In_2840,In_3436);
nor U776 (N_776,In_358,In_3654);
or U777 (N_777,In_2314,In_4813);
nand U778 (N_778,In_3673,In_188);
or U779 (N_779,In_3778,In_2796);
or U780 (N_780,In_4787,In_1330);
or U781 (N_781,In_2028,In_3904);
or U782 (N_782,In_109,In_1454);
and U783 (N_783,In_1744,In_1612);
nor U784 (N_784,In_1853,In_1561);
xor U785 (N_785,In_3988,In_2096);
nand U786 (N_786,In_1236,In_1084);
nand U787 (N_787,In_4794,In_249);
nor U788 (N_788,In_2199,In_4415);
or U789 (N_789,In_4682,In_4369);
nand U790 (N_790,In_3876,In_2426);
xnor U791 (N_791,In_2463,In_2953);
and U792 (N_792,In_3116,In_2560);
and U793 (N_793,In_4184,In_3554);
xor U794 (N_794,In_4294,In_3535);
nand U795 (N_795,In_2110,In_2333);
or U796 (N_796,In_3371,In_1730);
or U797 (N_797,In_1939,In_1335);
and U798 (N_798,In_3035,In_3670);
nor U799 (N_799,In_1629,In_957);
xor U800 (N_800,In_2956,In_2752);
xnor U801 (N_801,In_4658,In_813);
and U802 (N_802,In_1787,In_4942);
nor U803 (N_803,In_3154,In_2994);
nand U804 (N_804,In_1713,In_1573);
xor U805 (N_805,In_107,In_686);
nor U806 (N_806,In_3544,In_648);
nor U807 (N_807,In_3428,In_4758);
nor U808 (N_808,In_1269,In_3135);
nand U809 (N_809,In_3379,In_2403);
and U810 (N_810,In_4925,In_4232);
or U811 (N_811,In_1652,In_3166);
or U812 (N_812,In_211,In_2458);
or U813 (N_813,In_3763,In_1096);
and U814 (N_814,In_3662,In_4817);
nor U815 (N_815,In_856,In_992);
or U816 (N_816,In_3955,In_2116);
or U817 (N_817,In_3377,In_421);
nand U818 (N_818,In_4990,In_4185);
nand U819 (N_819,In_4713,In_4841);
nor U820 (N_820,In_2880,In_3933);
or U821 (N_821,In_145,In_1273);
or U822 (N_822,In_2924,In_182);
xor U823 (N_823,In_2519,In_2039);
nand U824 (N_824,In_1085,In_384);
and U825 (N_825,In_2084,In_1556);
or U826 (N_826,In_858,In_424);
nor U827 (N_827,In_86,In_4398);
and U828 (N_828,In_3410,In_213);
nor U829 (N_829,In_406,In_1919);
xor U830 (N_830,In_3078,In_1906);
nand U831 (N_831,In_952,In_1723);
and U832 (N_832,In_1924,In_4074);
and U833 (N_833,In_60,In_2571);
or U834 (N_834,In_4605,In_1181);
xor U835 (N_835,In_3715,In_951);
or U836 (N_836,In_1099,In_439);
xor U837 (N_837,In_4917,In_1317);
nor U838 (N_838,In_2584,In_2673);
nand U839 (N_839,In_2190,In_4544);
or U840 (N_840,In_2608,In_121);
or U841 (N_841,In_4368,In_3147);
or U842 (N_842,In_2192,In_95);
and U843 (N_843,In_1554,In_2728);
nor U844 (N_844,In_83,In_3122);
or U845 (N_845,In_2835,In_4065);
or U846 (N_846,In_2815,In_4572);
and U847 (N_847,In_4958,In_2526);
and U848 (N_848,In_2734,In_3539);
nand U849 (N_849,In_3350,In_3892);
nand U850 (N_850,In_1776,In_4783);
nand U851 (N_851,In_1704,In_928);
and U852 (N_852,In_1107,In_4367);
and U853 (N_853,In_493,In_2665);
and U854 (N_854,In_2943,In_855);
nor U855 (N_855,In_807,In_1786);
nor U856 (N_856,In_3362,In_1038);
or U857 (N_857,In_2564,In_32);
or U858 (N_858,In_1491,In_3225);
or U859 (N_859,In_2674,In_1212);
nor U860 (N_860,In_4939,In_4731);
nor U861 (N_861,In_1298,In_2917);
nand U862 (N_862,In_506,In_3885);
and U863 (N_863,In_4373,In_4584);
or U864 (N_864,In_548,In_1369);
or U865 (N_865,In_4062,In_3336);
and U866 (N_866,In_4340,In_2406);
nor U867 (N_867,In_2060,In_1359);
and U868 (N_868,In_2547,In_1062);
nor U869 (N_869,In_4418,In_3499);
nand U870 (N_870,In_3819,In_2829);
nor U871 (N_871,In_4997,In_355);
nor U872 (N_872,In_2716,In_4908);
or U873 (N_873,In_3285,In_4688);
and U874 (N_874,In_3829,In_2123);
nand U875 (N_875,In_4621,In_4978);
or U876 (N_876,In_1604,In_3158);
nor U877 (N_877,In_1838,In_2494);
or U878 (N_878,In_175,In_2947);
and U879 (N_879,In_1753,In_3502);
or U880 (N_880,In_3272,In_2227);
nor U881 (N_881,In_2971,In_2862);
nor U882 (N_882,In_3726,In_3817);
nand U883 (N_883,In_1875,In_4982);
and U884 (N_884,In_1696,In_3039);
xor U885 (N_885,In_2296,In_1286);
or U886 (N_886,In_1682,In_3710);
nor U887 (N_887,In_491,In_2369);
nand U888 (N_888,In_190,In_3612);
nand U889 (N_889,In_2462,In_4038);
and U890 (N_890,In_2756,In_212);
or U891 (N_891,In_3184,In_4507);
nor U892 (N_892,In_2874,In_4274);
or U893 (N_893,In_3175,In_3238);
or U894 (N_894,In_899,In_4458);
and U895 (N_895,In_294,In_2868);
nand U896 (N_896,In_3640,In_675);
xnor U897 (N_897,In_2510,In_3946);
nor U898 (N_898,In_3576,In_4618);
nand U899 (N_899,In_802,In_4333);
nor U900 (N_900,In_1071,In_3339);
nand U901 (N_901,In_2724,In_396);
nor U902 (N_902,In_3449,In_2276);
and U903 (N_903,In_704,In_1169);
nand U904 (N_904,In_1003,In_2066);
nand U905 (N_905,In_4767,In_2077);
nor U906 (N_906,In_2967,In_3006);
or U907 (N_907,In_2929,In_1030);
and U908 (N_908,In_1142,In_784);
nor U909 (N_909,In_1059,In_1981);
and U910 (N_910,In_2207,In_2797);
nor U911 (N_911,In_3713,In_4831);
nor U912 (N_912,In_100,In_2729);
and U913 (N_913,In_1167,In_3808);
and U914 (N_914,In_808,In_4582);
or U915 (N_915,In_1496,In_3943);
or U916 (N_916,In_3750,In_4712);
xnor U917 (N_917,In_120,In_3520);
or U918 (N_918,In_1770,In_4545);
nor U919 (N_919,In_4969,In_3968);
xor U920 (N_920,In_2034,In_235);
and U921 (N_921,In_597,In_2145);
nor U922 (N_922,In_3218,In_305);
or U923 (N_923,In_260,In_1201);
nor U924 (N_924,In_3415,In_35);
xor U925 (N_925,In_220,In_1717);
nor U926 (N_926,In_1868,In_3513);
and U927 (N_927,In_2642,In_457);
nand U928 (N_928,In_150,In_1724);
and U929 (N_929,In_1772,In_183);
nor U930 (N_930,In_4559,In_158);
or U931 (N_931,In_4861,In_2877);
nor U932 (N_932,In_4769,In_1155);
nand U933 (N_933,In_318,In_4880);
nor U934 (N_934,In_4378,In_4191);
and U935 (N_935,In_1134,In_4063);
or U936 (N_936,In_4000,In_2396);
nand U937 (N_937,In_1633,In_4916);
or U938 (N_938,In_1287,In_830);
nor U939 (N_939,In_2580,In_1171);
xnor U940 (N_940,In_3849,In_427);
nor U941 (N_941,In_4308,In_4664);
and U942 (N_942,In_898,In_4176);
nor U943 (N_943,In_3884,In_2846);
nor U944 (N_944,In_2417,In_2478);
nor U945 (N_945,In_1150,In_3545);
nand U946 (N_946,In_3117,In_4205);
or U947 (N_947,In_557,In_1574);
and U948 (N_948,In_2505,In_48);
nand U949 (N_949,In_1148,In_4066);
nand U950 (N_950,In_503,In_1508);
and U951 (N_951,In_3083,In_889);
or U952 (N_952,In_1624,In_4927);
or U953 (N_953,In_4633,In_999);
nor U954 (N_954,In_170,In_4612);
and U955 (N_955,In_3509,In_2790);
and U956 (N_956,In_1701,In_4313);
xnor U957 (N_957,In_3772,In_1147);
and U958 (N_958,In_876,In_925);
nor U959 (N_959,In_3740,In_36);
and U960 (N_960,In_4085,In_1908);
or U961 (N_961,In_2270,In_3651);
xor U962 (N_962,In_403,In_1495);
nand U963 (N_963,In_1202,In_2534);
and U964 (N_964,In_317,In_3311);
and U965 (N_965,In_2251,In_1912);
xnor U966 (N_966,In_1088,In_3369);
nand U967 (N_967,In_4043,In_1231);
nor U968 (N_968,In_2849,In_1391);
nor U969 (N_969,In_4543,In_2561);
nor U970 (N_970,In_3441,In_3472);
and U971 (N_971,In_2467,In_1352);
nor U972 (N_972,In_3429,In_4476);
or U973 (N_973,In_3574,In_2303);
nand U974 (N_974,In_1893,In_1921);
or U975 (N_975,In_563,In_2793);
nor U976 (N_976,In_2180,In_1941);
nor U977 (N_977,In_4546,In_1492);
nand U978 (N_978,In_1961,In_1585);
or U979 (N_979,In_3660,In_3694);
nand U980 (N_980,In_1694,In_3745);
and U981 (N_981,In_3114,In_184);
or U982 (N_982,In_4808,In_1627);
and U983 (N_983,In_4583,In_4941);
and U984 (N_984,In_1863,In_2422);
or U985 (N_985,In_901,In_1642);
nor U986 (N_986,In_1533,In_3762);
and U987 (N_987,In_1955,In_1732);
and U988 (N_988,In_4482,In_3982);
and U989 (N_989,In_2804,In_41);
xnor U990 (N_990,In_3030,In_2550);
nor U991 (N_991,In_2920,In_4275);
and U992 (N_992,In_3199,In_4351);
xnor U993 (N_993,In_1420,In_4862);
nand U994 (N_994,In_4401,In_3842);
xnor U995 (N_995,In_603,In_3519);
or U996 (N_996,In_3064,In_3900);
or U997 (N_997,In_3958,In_900);
and U998 (N_998,In_2290,In_4739);
nor U999 (N_999,In_1800,In_2824);
nor U1000 (N_1000,In_278,In_4674);
xor U1001 (N_1001,In_392,In_4720);
or U1002 (N_1002,In_2335,In_2438);
and U1003 (N_1003,In_3774,In_349);
and U1004 (N_1004,In_2926,In_1076);
or U1005 (N_1005,In_3799,In_769);
and U1006 (N_1006,In_896,In_3119);
and U1007 (N_1007,In_3059,In_3108);
and U1008 (N_1008,In_3800,In_1864);
or U1009 (N_1009,In_2415,In_958);
nor U1010 (N_1010,In_667,In_1350);
xor U1011 (N_1011,In_4575,In_2143);
nand U1012 (N_1012,In_4264,In_1048);
or U1013 (N_1013,In_4928,In_1581);
nor U1014 (N_1014,In_453,In_4092);
nand U1015 (N_1015,In_1935,In_4487);
xnor U1016 (N_1016,In_2680,In_522);
and U1017 (N_1017,In_744,In_3197);
nand U1018 (N_1018,In_195,In_397);
and U1019 (N_1019,In_1466,In_1953);
nand U1020 (N_1020,In_835,In_4366);
and U1021 (N_1021,In_746,In_706);
nor U1022 (N_1022,In_2221,In_3130);
xor U1023 (N_1023,In_2604,In_2583);
and U1024 (N_1024,In_1630,In_722);
nand U1025 (N_1025,In_2761,In_3677);
nand U1026 (N_1026,In_953,In_1599);
or U1027 (N_1027,In_4027,In_4904);
and U1028 (N_1028,In_4820,In_3735);
nand U1029 (N_1029,In_4608,In_4938);
nor U1030 (N_1030,In_2837,In_3625);
or U1031 (N_1031,In_4439,In_2056);
nand U1032 (N_1032,In_1531,In_4384);
xor U1033 (N_1033,In_3478,In_3426);
nand U1034 (N_1034,In_4549,In_3259);
or U1035 (N_1035,In_4651,In_248);
nor U1036 (N_1036,In_3071,In_4866);
or U1037 (N_1037,In_4193,In_2443);
or U1038 (N_1038,In_4497,In_328);
or U1039 (N_1039,In_2246,In_2016);
or U1040 (N_1040,In_1430,In_4189);
and U1041 (N_1041,In_1777,In_2038);
or U1042 (N_1042,In_3597,In_3058);
or U1043 (N_1043,In_859,In_4993);
nand U1044 (N_1044,In_755,In_770);
nand U1045 (N_1045,In_4466,In_4814);
and U1046 (N_1046,In_4100,In_3570);
nand U1047 (N_1047,In_3080,In_2351);
nor U1048 (N_1048,In_4762,In_2392);
or U1049 (N_1049,In_1471,In_4323);
and U1050 (N_1050,In_216,In_2973);
xnor U1051 (N_1051,In_3566,In_551);
nand U1052 (N_1052,In_3717,In_4243);
or U1053 (N_1053,In_2618,In_4129);
and U1054 (N_1054,In_3703,In_271);
or U1055 (N_1055,In_1756,In_1328);
nand U1056 (N_1056,In_2419,In_630);
or U1057 (N_1057,In_2464,In_2963);
nor U1058 (N_1058,In_2252,In_3060);
and U1059 (N_1059,In_459,In_1750);
and U1060 (N_1060,In_4073,In_989);
nor U1061 (N_1061,In_2888,In_1439);
nor U1062 (N_1062,In_2146,In_1763);
nor U1063 (N_1063,In_2538,In_646);
or U1064 (N_1064,In_2416,In_2357);
nor U1065 (N_1065,In_767,In_4040);
xnor U1066 (N_1066,In_3575,In_2449);
and U1067 (N_1067,In_526,In_252);
or U1068 (N_1068,In_299,In_3385);
and U1069 (N_1069,In_3888,In_2374);
or U1070 (N_1070,In_3598,In_4683);
or U1071 (N_1071,In_4155,In_498);
nand U1072 (N_1072,In_2201,In_4973);
and U1073 (N_1073,In_4409,In_4944);
and U1074 (N_1074,In_3665,In_4800);
nand U1075 (N_1075,In_2006,In_3783);
nand U1076 (N_1076,In_3619,In_512);
xnor U1077 (N_1077,In_1976,In_4746);
nor U1078 (N_1078,In_904,In_1645);
nor U1079 (N_1079,In_79,In_484);
and U1080 (N_1080,In_4036,In_3133);
nor U1081 (N_1081,In_3894,In_1224);
and U1082 (N_1082,In_1461,In_3034);
or U1083 (N_1083,In_1871,In_1204);
nand U1084 (N_1084,In_4121,In_829);
nor U1085 (N_1085,In_1982,In_4609);
nor U1086 (N_1086,In_3138,In_1428);
and U1087 (N_1087,In_3769,In_3901);
and U1088 (N_1088,In_4728,In_2749);
or U1089 (N_1089,In_3860,In_2962);
xnor U1090 (N_1090,In_7,In_2907);
and U1091 (N_1091,In_2289,In_4786);
xnor U1092 (N_1092,In_472,In_3300);
and U1093 (N_1093,In_4445,In_639);
nand U1094 (N_1094,In_26,In_3538);
or U1095 (N_1095,In_11,In_3149);
xor U1096 (N_1096,In_74,In_4976);
and U1097 (N_1097,In_3142,In_290);
or U1098 (N_1098,In_1362,In_4116);
nor U1099 (N_1099,In_1444,In_4011);
nor U1100 (N_1100,In_1885,In_4875);
nand U1101 (N_1101,In_2810,In_3650);
nor U1102 (N_1102,In_4579,In_1259);
or U1103 (N_1103,In_508,In_3005);
nor U1104 (N_1104,In_4332,In_255);
nand U1105 (N_1105,In_971,In_142);
or U1106 (N_1106,In_2916,In_3473);
nor U1107 (N_1107,In_14,In_3861);
nor U1108 (N_1108,In_3847,In_2799);
nor U1109 (N_1109,In_2093,In_2682);
nor U1110 (N_1110,In_3500,In_2932);
or U1111 (N_1111,In_2341,In_1515);
nor U1112 (N_1112,In_492,In_2241);
and U1113 (N_1113,In_2309,In_2064);
or U1114 (N_1114,In_4201,In_3388);
nand U1115 (N_1115,In_2196,In_1230);
and U1116 (N_1116,In_3139,In_4740);
nand U1117 (N_1117,In_4042,In_2414);
nand U1118 (N_1118,In_3752,In_2594);
xor U1119 (N_1119,In_1243,In_2867);
and U1120 (N_1120,In_1707,In_2472);
and U1121 (N_1121,In_319,In_3501);
nand U1122 (N_1122,In_865,In_2058);
nand U1123 (N_1123,In_2115,In_1265);
or U1124 (N_1124,In_4433,In_4833);
nand U1125 (N_1125,In_2171,In_996);
nand U1126 (N_1126,In_1014,In_1994);
and U1127 (N_1127,In_192,In_469);
nor U1128 (N_1128,In_3136,In_366);
nand U1129 (N_1129,In_2157,In_2760);
nor U1130 (N_1130,In_4754,In_12);
or U1131 (N_1131,In_4215,In_1691);
xnor U1132 (N_1132,In_2218,In_4652);
nand U1133 (N_1133,In_245,In_4376);
nor U1134 (N_1134,In_2053,In_258);
nand U1135 (N_1135,In_4157,In_286);
or U1136 (N_1136,In_3588,In_3531);
and U1137 (N_1137,In_1498,In_4905);
and U1138 (N_1138,In_1679,In_2791);
nand U1139 (N_1139,In_3041,In_2019);
or U1140 (N_1140,In_3728,In_2283);
or U1141 (N_1141,In_4382,In_4818);
and U1142 (N_1142,In_3212,In_4080);
nand U1143 (N_1143,In_1923,In_3323);
and U1144 (N_1144,In_2105,In_3678);
nand U1145 (N_1145,In_4127,In_3529);
nor U1146 (N_1146,In_4530,In_2461);
or U1147 (N_1147,In_3392,In_4809);
or U1148 (N_1148,In_3835,In_586);
or U1149 (N_1149,In_1847,In_3906);
xnor U1150 (N_1150,In_4850,In_1999);
nand U1151 (N_1151,In_4389,In_3751);
nor U1152 (N_1152,In_89,In_2295);
and U1153 (N_1153,In_1532,In_1718);
or U1154 (N_1154,In_1053,In_9);
or U1155 (N_1155,In_1393,In_1294);
or U1156 (N_1156,In_4251,In_4897);
nand U1157 (N_1157,In_4427,In_115);
nand U1158 (N_1158,In_1910,In_1993);
or U1159 (N_1159,In_962,In_4929);
nand U1160 (N_1160,In_3756,In_4234);
or U1161 (N_1161,In_840,In_4859);
xnor U1162 (N_1162,In_1665,In_3540);
nor U1163 (N_1163,In_28,In_2765);
nor U1164 (N_1164,In_38,In_2628);
nand U1165 (N_1165,In_2662,In_3963);
nand U1166 (N_1166,In_2974,In_4137);
or U1167 (N_1167,In_4729,In_1938);
nor U1168 (N_1168,In_4242,In_1198);
xor U1169 (N_1169,In_435,In_3310);
and U1170 (N_1170,In_3656,In_1687);
nand U1171 (N_1171,In_1565,In_2989);
xor U1172 (N_1172,In_1160,In_4158);
and U1173 (N_1173,In_4257,In_2959);
nand U1174 (N_1174,In_3179,In_1658);
nand U1175 (N_1175,In_1940,In_743);
xor U1176 (N_1176,In_4779,In_117);
or U1177 (N_1177,In_1549,In_3306);
and U1178 (N_1178,In_1536,In_3235);
and U1179 (N_1179,In_3354,In_1482);
nand U1180 (N_1180,In_752,In_1299);
or U1181 (N_1181,In_3367,In_2141);
or U1182 (N_1182,In_4771,In_225);
nor U1183 (N_1183,In_202,In_4741);
nor U1184 (N_1184,In_4068,In_4001);
and U1185 (N_1185,In_2502,In_4322);
or U1186 (N_1186,In_487,In_569);
and U1187 (N_1187,In_803,In_4350);
nand U1188 (N_1188,In_4407,In_3488);
xor U1189 (N_1189,In_2589,In_2024);
xor U1190 (N_1190,In_3214,In_3896);
nand U1191 (N_1191,In_728,In_401);
nand U1192 (N_1192,In_1877,In_451);
xnor U1193 (N_1193,In_4183,In_4681);
and U1194 (N_1194,In_2546,In_930);
nor U1195 (N_1195,In_2387,In_4144);
or U1196 (N_1196,In_3899,In_4337);
or U1197 (N_1197,In_326,In_4812);
and U1198 (N_1198,In_4165,In_4154);
or U1199 (N_1199,In_1251,In_4777);
xnor U1200 (N_1200,In_3548,In_3653);
and U1201 (N_1201,In_3814,In_4893);
xnor U1202 (N_1202,In_4940,In_599);
nand U1203 (N_1203,In_554,In_3200);
or U1204 (N_1204,In_1410,In_2050);
nor U1205 (N_1205,In_4160,In_2945);
and U1206 (N_1206,In_1326,In_2850);
and U1207 (N_1207,In_1128,In_3960);
or U1208 (N_1208,In_3891,In_3012);
and U1209 (N_1209,In_306,In_2336);
nor U1210 (N_1210,In_340,In_4306);
or U1211 (N_1211,In_1377,In_2949);
nor U1212 (N_1212,In_1371,In_2513);
nand U1213 (N_1213,In_2301,In_4053);
and U1214 (N_1214,In_4411,In_3128);
xnor U1215 (N_1215,In_3266,In_1164);
xnor U1216 (N_1216,In_2255,In_4947);
or U1217 (N_1217,In_684,In_2343);
or U1218 (N_1218,In_519,In_2228);
or U1219 (N_1219,In_4540,In_4112);
and U1220 (N_1220,In_950,In_2861);
or U1221 (N_1221,In_4298,In_4077);
nor U1222 (N_1222,In_2950,In_2698);
and U1223 (N_1223,In_2497,In_2112);
and U1224 (N_1224,In_1804,In_4186);
or U1225 (N_1225,In_1361,In_3864);
xnor U1226 (N_1226,In_2681,In_4220);
nand U1227 (N_1227,In_3890,In_4288);
or U1228 (N_1228,In_1631,In_490);
xnor U1229 (N_1229,In_4956,In_713);
nor U1230 (N_1230,In_1049,In_3804);
nor U1231 (N_1231,In_2704,In_3391);
nor U1232 (N_1232,In_222,In_4816);
or U1233 (N_1233,In_2186,In_3526);
nor U1234 (N_1234,In_1474,In_2485);
and U1235 (N_1235,In_2677,In_1887);
nor U1236 (N_1236,In_3870,In_2667);
or U1237 (N_1237,In_344,In_4923);
nor U1238 (N_1238,In_4246,In_2838);
nor U1239 (N_1239,In_4694,In_1173);
nand U1240 (N_1240,In_3076,In_2896);
xor U1241 (N_1241,In_2566,In_1639);
and U1242 (N_1242,In_3533,In_246);
and U1243 (N_1243,In_1990,In_1815);
or U1244 (N_1244,In_582,In_4348);
or U1245 (N_1245,In_3219,In_2260);
or U1246 (N_1246,In_1872,In_4719);
nand U1247 (N_1247,In_2427,In_1802);
and U1248 (N_1248,In_3518,In_4025);
nor U1249 (N_1249,In_574,In_477);
xnor U1250 (N_1250,In_1807,In_2117);
xnor U1251 (N_1251,In_3983,In_2575);
or U1252 (N_1252,In_2795,In_2404);
nor U1253 (N_1253,In_3626,In_4159);
nand U1254 (N_1254,In_1743,In_2649);
xnor U1255 (N_1255,In_4541,In_3089);
and U1256 (N_1256,In_3031,In_2574);
and U1257 (N_1257,In_4171,In_3228);
and U1258 (N_1258,In_3454,In_3578);
or U1259 (N_1259,In_1790,In_2098);
or U1260 (N_1260,In_1486,In_1039);
xor U1261 (N_1261,In_1433,In_1827);
nor U1262 (N_1262,In_4499,In_561);
and U1263 (N_1263,In_3725,In_1227);
nand U1264 (N_1264,In_2500,In_821);
nand U1265 (N_1265,In_737,In_4107);
and U1266 (N_1266,In_1856,In_97);
and U1267 (N_1267,In_4837,In_2539);
or U1268 (N_1268,In_1674,In_4684);
nor U1269 (N_1269,In_2965,In_1685);
and U1270 (N_1270,In_3360,In_4509);
nand U1271 (N_1271,In_2637,In_892);
nor U1272 (N_1272,In_2557,In_825);
or U1273 (N_1273,In_2876,In_1205);
or U1274 (N_1274,In_4400,In_2934);
or U1275 (N_1275,In_311,In_4824);
or U1276 (N_1276,In_44,In_2958);
nor U1277 (N_1277,In_4008,In_631);
nor U1278 (N_1278,In_3052,In_3198);
nor U1279 (N_1279,In_1914,In_4383);
and U1280 (N_1280,In_2533,In_17);
and U1281 (N_1281,In_644,In_3691);
or U1282 (N_1282,In_1621,In_3719);
and U1283 (N_1283,In_4735,In_4064);
nor U1284 (N_1284,In_3016,In_2106);
xor U1285 (N_1285,In_309,In_3084);
xnor U1286 (N_1286,In_4565,In_3131);
nor U1287 (N_1287,In_4949,In_3047);
nand U1288 (N_1288,In_3094,In_955);
and U1289 (N_1289,In_3249,In_3274);
and U1290 (N_1290,In_2768,In_1355);
or U1291 (N_1291,In_2827,In_205);
xor U1292 (N_1292,In_2261,In_1721);
nand U1293 (N_1293,In_4805,In_4943);
nand U1294 (N_1294,In_702,In_3877);
nor U1295 (N_1295,In_383,In_3438);
or U1296 (N_1296,In_3748,In_4631);
nand U1297 (N_1297,In_3517,In_1859);
or U1298 (N_1298,In_2352,In_3201);
nand U1299 (N_1299,In_883,In_1916);
and U1300 (N_1300,In_1635,In_308);
or U1301 (N_1301,In_2639,In_365);
and U1302 (N_1302,In_1229,In_2606);
and U1303 (N_1303,In_410,In_4197);
xnor U1304 (N_1304,In_4521,In_442);
or U1305 (N_1305,In_3664,In_3110);
nor U1306 (N_1306,In_3164,In_3291);
and U1307 (N_1307,In_1586,In_4673);
or U1308 (N_1308,In_3492,In_3440);
nand U1309 (N_1309,In_617,In_1017);
nand U1310 (N_1310,In_2492,In_2873);
nor U1311 (N_1311,In_1470,In_2726);
nand U1312 (N_1312,In_187,In_711);
nand U1313 (N_1313,In_1782,In_129);
nor U1314 (N_1314,In_3,In_3865);
and U1315 (N_1315,In_2927,In_2864);
and U1316 (N_1316,In_3579,In_3446);
nor U1317 (N_1317,In_780,In_1667);
nand U1318 (N_1318,In_2223,In_4537);
nor U1319 (N_1319,In_2173,In_4204);
and U1320 (N_1320,In_3582,In_3585);
and U1321 (N_1321,In_732,In_1214);
nor U1322 (N_1322,In_837,In_4375);
nor U1323 (N_1323,In_3358,In_4919);
nand U1324 (N_1324,In_146,In_4611);
nand U1325 (N_1325,In_4495,In_2894);
or U1326 (N_1326,In_1958,In_2766);
nor U1327 (N_1327,In_1322,In_2360);
and U1328 (N_1328,In_2805,In_3942);
xnor U1329 (N_1329,In_3173,In_1734);
or U1330 (N_1330,In_1576,In_2408);
nand U1331 (N_1331,In_3236,In_3965);
nand U1332 (N_1332,In_894,In_3856);
or U1333 (N_1333,In_485,In_2692);
nor U1334 (N_1334,In_3621,In_1418);
and U1335 (N_1335,In_2204,In_2405);
or U1336 (N_1336,In_542,In_4886);
or U1337 (N_1337,In_2131,In_4304);
nand U1338 (N_1338,In_429,In_3907);
or U1339 (N_1339,In_169,In_2032);
nor U1340 (N_1340,In_4315,In_387);
nor U1341 (N_1341,In_2307,In_1494);
and U1342 (N_1342,In_4034,In_523);
nor U1343 (N_1343,In_1987,In_2743);
xor U1344 (N_1344,In_4692,In_2063);
or U1345 (N_1345,In_1174,In_409);
nor U1346 (N_1346,In_3497,In_104);
nand U1347 (N_1347,In_2089,In_3247);
and U1348 (N_1348,In_4349,In_155);
or U1349 (N_1349,In_370,In_3124);
and U1350 (N_1350,In_4594,In_3599);
or U1351 (N_1351,In_4874,In_670);
xor U1352 (N_1352,In_902,In_460);
and U1353 (N_1353,In_3375,In_2071);
or U1354 (N_1354,In_3883,In_3887);
and U1355 (N_1355,In_412,In_3846);
and U1356 (N_1356,In_4414,In_4434);
or U1357 (N_1357,In_2992,In_2496);
nand U1358 (N_1358,In_4743,In_2858);
or U1359 (N_1359,In_4585,In_3813);
or U1360 (N_1360,In_1551,In_917);
xnor U1361 (N_1361,In_4613,In_2672);
and U1362 (N_1362,In_3485,In_1037);
xnor U1363 (N_1363,In_3361,In_1389);
nor U1364 (N_1364,In_714,In_2787);
and U1365 (N_1365,In_863,In_237);
or U1366 (N_1366,In_2721,In_1453);
nor U1367 (N_1367,In_1520,In_2040);
nor U1368 (N_1368,In_963,In_1089);
and U1369 (N_1369,In_2248,In_1468);
nand U1370 (N_1370,In_2784,In_4392);
or U1371 (N_1371,In_3413,In_3557);
and U1372 (N_1372,In_2661,In_3260);
nor U1373 (N_1373,In_1754,In_1767);
xor U1374 (N_1374,In_438,In_256);
nand U1375 (N_1375,In_964,In_2061);
and U1376 (N_1376,In_2432,In_2828);
nand U1377 (N_1377,In_1651,In_373);
nor U1378 (N_1378,In_4465,In_4123);
or U1379 (N_1379,In_1608,In_1947);
nand U1380 (N_1380,In_3435,In_2152);
nand U1381 (N_1381,In_1584,In_3390);
nor U1382 (N_1382,In_2747,In_4423);
nand U1383 (N_1383,In_2466,In_3506);
xor U1384 (N_1384,In_3922,In_1206);
xor U1385 (N_1385,In_4420,In_3104);
nor U1386 (N_1386,In_593,In_3397);
or U1387 (N_1387,In_4525,In_4591);
nor U1388 (N_1388,In_254,In_3081);
and U1389 (N_1389,In_1731,In_4015);
nor U1390 (N_1390,In_1527,In_1097);
nand U1391 (N_1391,In_330,In_1946);
and U1392 (N_1392,In_3895,In_3606);
nor U1393 (N_1393,In_4039,In_2879);
or U1394 (N_1394,In_1449,In_3882);
nor U1395 (N_1395,In_872,In_2705);
and U1396 (N_1396,In_1380,In_4560);
and U1397 (N_1397,In_2632,In_4356);
nor U1398 (N_1398,In_2706,In_3209);
nor U1399 (N_1399,In_3661,In_448);
or U1400 (N_1400,In_3954,In_3630);
nor U1401 (N_1401,In_3250,In_118);
nor U1402 (N_1402,In_4138,In_1930);
and U1403 (N_1403,In_122,In_3482);
or U1404 (N_1404,In_2213,In_1306);
nor U1405 (N_1405,In_3073,In_3495);
nor U1406 (N_1406,In_4845,In_726);
nand U1407 (N_1407,In_4395,In_2451);
nand U1408 (N_1408,In_2318,In_3177);
nor U1409 (N_1409,In_3766,In_4141);
and U1410 (N_1410,In_3985,In_4648);
nor U1411 (N_1411,In_4054,In_1024);
nand U1412 (N_1412,In_3319,In_3050);
or U1413 (N_1413,In_2377,In_3839);
nor U1414 (N_1414,In_3587,In_4872);
and U1415 (N_1415,In_1680,In_2712);
nand U1416 (N_1416,In_4360,In_4223);
or U1417 (N_1417,In_4513,In_1390);
and U1418 (N_1418,In_4117,In_3113);
nor U1419 (N_1419,In_1580,In_4300);
or U1420 (N_1420,In_444,In_959);
nor U1421 (N_1421,In_262,In_3145);
nor U1422 (N_1422,In_3781,In_20);
nand U1423 (N_1423,In_240,In_3534);
nand U1424 (N_1424,In_4055,In_3609);
nor U1425 (N_1425,In_2244,In_1034);
or U1426 (N_1426,In_1345,In_196);
nor U1427 (N_1427,In_534,In_4405);
or U1428 (N_1428,In_2001,In_2368);
nor U1429 (N_1429,In_4957,In_3730);
or U1430 (N_1430,In_3874,In_1379);
nand U1431 (N_1431,In_3921,In_3863);
nand U1432 (N_1432,In_1254,In_4057);
xnor U1433 (N_1433,In_4792,In_4516);
or U1434 (N_1434,In_4984,In_4967);
nand U1435 (N_1435,In_1759,In_2772);
nand U1436 (N_1436,In_2097,In_1751);
or U1437 (N_1437,In_3153,In_3297);
nor U1438 (N_1438,In_3927,In_2570);
nor U1439 (N_1439,In_2695,In_2572);
and U1440 (N_1440,In_3378,In_3854);
nor U1441 (N_1441,In_3207,In_3163);
or U1442 (N_1442,In_4326,In_2762);
nand U1443 (N_1443,In_445,In_4529);
and U1444 (N_1444,In_1098,In_4329);
nand U1445 (N_1445,In_4325,In_1823);
or U1446 (N_1446,In_345,In_488);
xor U1447 (N_1447,In_3918,In_3105);
nor U1448 (N_1448,In_2885,In_1821);
or U1449 (N_1449,In_3193,In_1246);
nor U1450 (N_1450,In_3558,In_982);
nand U1451 (N_1451,In_2072,In_2872);
nor U1452 (N_1452,In_296,In_1768);
nor U1453 (N_1453,In_1820,In_4492);
or U1454 (N_1454,In_1858,In_1007);
and U1455 (N_1455,In_2814,In_2875);
and U1456 (N_1456,In_500,In_3208);
xnor U1457 (N_1457,In_703,In_475);
nor U1458 (N_1458,In_1558,In_2036);
nor U1459 (N_1459,In_1360,In_4361);
nand U1460 (N_1460,In_2979,In_4030);
and U1461 (N_1461,In_4140,In_1464);
or U1462 (N_1462,In_3220,In_1216);
xnor U1463 (N_1463,In_4705,In_3838);
nand U1464 (N_1464,In_2100,In_2103);
xor U1465 (N_1465,In_3524,In_1737);
and U1466 (N_1466,In_4455,In_3403);
nand U1467 (N_1467,In_4974,In_2128);
nor U1468 (N_1468,In_4075,In_3271);
or U1469 (N_1469,In_3342,In_4106);
xnor U1470 (N_1470,In_3989,In_1542);
or U1471 (N_1471,In_4303,In_2635);
and U1472 (N_1472,In_3591,In_3836);
or U1473 (N_1473,In_4970,In_2788);
or U1474 (N_1474,In_51,In_494);
and U1475 (N_1475,In_937,In_2043);
and U1476 (N_1476,In_1881,In_3070);
nor U1477 (N_1477,In_4979,In_939);
nor U1478 (N_1478,In_2893,In_1019);
nor U1479 (N_1479,In_1783,In_4638);
or U1480 (N_1480,In_4706,In_2175);
nand U1481 (N_1481,In_2495,In_2075);
and U1482 (N_1482,In_103,In_2800);
and U1483 (N_1483,In_1116,In_2964);
nor U1484 (N_1484,In_1882,In_1521);
and U1485 (N_1485,In_3775,In_2910);
and U1486 (N_1486,In_785,In_738);
or U1487 (N_1487,In_2062,In_3999);
and U1488 (N_1488,In_1911,In_2833);
nor U1489 (N_1489,In_3287,In_2774);
and U1490 (N_1490,In_592,In_2259);
nand U1491 (N_1491,In_85,In_3168);
nand U1492 (N_1492,In_1500,In_2986);
nand U1493 (N_1493,In_3121,In_2168);
xor U1494 (N_1494,In_3430,In_3481);
and U1495 (N_1495,In_3722,In_2078);
and U1496 (N_1496,In_1067,In_3761);
nor U1497 (N_1497,In_2905,In_4261);
or U1498 (N_1498,In_4146,In_2158);
or U1499 (N_1499,In_595,In_2159);
or U1500 (N_1500,In_799,In_3085);
xnor U1501 (N_1501,In_4724,In_4748);
nand U1502 (N_1502,In_1138,In_750);
xor U1503 (N_1503,In_1740,In_3784);
nand U1504 (N_1504,In_3749,In_223);
nor U1505 (N_1505,In_1438,In_2165);
nor U1506 (N_1506,In_2215,In_4920);
nand U1507 (N_1507,In_4484,In_3279);
or U1508 (N_1508,In_3618,In_1275);
xnor U1509 (N_1509,In_4959,In_3674);
nand U1510 (N_1510,In_4253,In_1276);
nand U1511 (N_1511,In_3959,In_3268);
nor U1512 (N_1512,In_2457,In_3873);
and U1513 (N_1513,In_976,In_2983);
and U1514 (N_1514,In_775,In_4882);
nand U1515 (N_1515,In_1735,In_3317);
xor U1516 (N_1516,In_3671,In_2737);
nand U1517 (N_1517,In_2133,In_1075);
nand U1518 (N_1518,In_2792,In_564);
nor U1519 (N_1519,In_4838,In_4443);
nand U1520 (N_1520,In_1161,In_2300);
nor U1521 (N_1521,In_2057,In_4267);
and U1522 (N_1522,In_3987,In_4768);
nor U1523 (N_1523,In_2946,In_4131);
nand U1524 (N_1524,In_3412,In_3115);
nor U1525 (N_1525,In_2185,In_2094);
or U1526 (N_1526,In_2742,In_1080);
nor U1527 (N_1527,In_3779,In_3825);
nand U1528 (N_1528,In_527,In_3191);
nor U1529 (N_1529,In_3973,In_4634);
xor U1530 (N_1530,In_2000,In_2599);
and U1531 (N_1531,In_1031,In_4098);
nand U1532 (N_1532,In_2688,In_3150);
nor U1533 (N_1533,In_2930,In_941);
nor U1534 (N_1534,In_4104,In_3183);
nand U1535 (N_1535,In_193,In_580);
nor U1536 (N_1536,In_3294,In_112);
nand U1537 (N_1537,In_3278,In_1726);
nand U1538 (N_1538,In_2286,In_2491);
nor U1539 (N_1539,In_2656,In_2121);
nand U1540 (N_1540,In_3118,In_2429);
and U1541 (N_1541,In_1479,In_2720);
or U1542 (N_1542,In_2839,In_3964);
nand U1543 (N_1543,In_2997,In_3623);
xnor U1544 (N_1544,In_4963,In_3226);
nand U1545 (N_1545,In_3537,In_3636);
and U1546 (N_1546,In_4319,In_3505);
or U1547 (N_1547,In_2108,In_4775);
and U1548 (N_1548,In_2315,In_3439);
and U1549 (N_1549,In_3000,In_4628);
or U1550 (N_1550,In_4983,In_4118);
or U1551 (N_1551,In_3898,In_4301);
nand U1552 (N_1552,In_377,In_4446);
and U1553 (N_1553,In_1653,In_3924);
nand U1554 (N_1554,In_4877,In_2648);
and U1555 (N_1555,In_2518,In_189);
nor U1556 (N_1556,In_805,In_263);
and U1557 (N_1557,In_2822,In_2806);
and U1558 (N_1558,In_3820,In_1032);
and U1559 (N_1559,In_2149,In_2041);
and U1560 (N_1560,In_3878,In_2109);
and U1561 (N_1561,In_1295,In_4653);
xnor U1562 (N_1562,In_4091,In_4086);
or U1563 (N_1563,In_1341,In_2634);
nor U1564 (N_1564,In_2499,In_4952);
nand U1565 (N_1565,In_3464,In_788);
nand U1566 (N_1566,In_2869,In_575);
nand U1567 (N_1567,In_3504,In_2479);
nand U1568 (N_1568,In_1431,In_4014);
nand U1569 (N_1569,In_1427,In_888);
nor U1570 (N_1570,In_2114,In_4708);
xnor U1571 (N_1571,In_1811,In_4136);
xor U1572 (N_1572,In_329,In_2230);
or U1573 (N_1573,In_4871,In_4182);
nor U1574 (N_1574,In_4626,In_1196);
or U1575 (N_1575,In_694,In_1144);
xor U1576 (N_1576,In_4755,In_1382);
xor U1577 (N_1577,In_2689,In_4679);
xor U1578 (N_1578,In_173,In_4134);
nand U1579 (N_1579,In_600,In_2782);
nor U1580 (N_1580,In_3709,In_2055);
nor U1581 (N_1581,In_2381,In_61);
or U1582 (N_1582,In_2702,In_3265);
or U1583 (N_1583,In_663,In_2210);
and U1584 (N_1584,In_1452,In_4240);
nor U1585 (N_1585,In_4505,In_695);
nor U1586 (N_1586,In_2154,In_2611);
nand U1587 (N_1587,In_3831,In_2998);
nor U1588 (N_1588,In_4671,In_1176);
nor U1589 (N_1589,In_315,In_1077);
or U1590 (N_1590,In_468,In_337);
nand U1591 (N_1591,In_2636,In_2552);
nand U1592 (N_1592,In_1572,In_2522);
nor U1593 (N_1593,In_1008,In_4644);
xnor U1594 (N_1594,In_3712,In_4865);
or U1595 (N_1595,In_3561,In_3137);
nor U1596 (N_1596,In_2245,In_181);
nand U1597 (N_1597,In_745,In_3013);
nor U1598 (N_1598,In_1363,In_3971);
nor U1599 (N_1599,In_2442,In_810);
nor U1600 (N_1600,In_4586,In_4723);
and U1601 (N_1601,In_2308,In_2860);
xor U1602 (N_1602,In_3851,In_3920);
nor U1603 (N_1603,In_1833,In_1021);
and U1604 (N_1604,In_1424,In_320);
nor U1605 (N_1605,In_4372,In_2182);
nand U1606 (N_1606,In_2684,In_502);
or U1607 (N_1607,In_3826,In_2187);
and U1608 (N_1608,In_4203,In_2739);
xor U1609 (N_1609,In_890,In_1399);
nand U1610 (N_1610,In_730,In_833);
and U1611 (N_1611,In_555,In_2870);
nor U1612 (N_1612,In_608,In_1669);
nand U1613 (N_1613,In_3352,In_4056);
nand U1614 (N_1614,In_1550,In_3639);
nor U1615 (N_1615,In_4364,In_3852);
nor U1616 (N_1616,In_536,In_3889);
xnor U1617 (N_1617,In_2701,In_3044);
or U1618 (N_1618,In_811,In_1045);
and U1619 (N_1619,In_3417,In_1123);
nor U1620 (N_1620,In_3809,In_4669);
nand U1621 (N_1621,In_2937,In_2395);
nand U1622 (N_1622,In_1623,In_1785);
nor U1623 (N_1623,In_1852,In_2049);
or U1624 (N_1624,In_134,In_3329);
or U1625 (N_1625,In_127,In_2854);
nor U1626 (N_1626,In_4844,In_3647);
or U1627 (N_1627,In_4722,In_2703);
nand U1628 (N_1628,In_3120,In_4355);
nand U1629 (N_1629,In_4806,In_1366);
nand U1630 (N_1630,In_3134,In_3832);
nor U1631 (N_1631,In_1249,In_1814);
xnor U1632 (N_1632,In_823,In_3063);
or U1633 (N_1633,In_3442,In_1290);
and U1634 (N_1634,In_283,In_431);
or U1635 (N_1635,In_1840,In_4438);
nor U1636 (N_1636,In_4440,In_4046);
and U1637 (N_1637,In_1703,In_507);
or U1638 (N_1638,In_331,In_1186);
and U1639 (N_1639,In_846,In_4258);
nand U1640 (N_1640,In_1873,In_4282);
and U1641 (N_1641,In_2022,In_3600);
and U1642 (N_1642,In_3990,In_851);
nor U1643 (N_1643,In_4696,In_972);
or U1644 (N_1644,In_2970,In_2254);
nor U1645 (N_1645,In_3705,In_4604);
and U1646 (N_1646,In_2009,In_747);
or U1647 (N_1647,In_3682,In_1051);
nor U1648 (N_1648,In_1028,In_3683);
or U1649 (N_1649,In_1332,In_3496);
xor U1650 (N_1650,In_622,In_1765);
nand U1651 (N_1651,In_2725,In_4295);
or U1652 (N_1652,In_3261,In_1655);
nor U1653 (N_1653,In_771,In_3727);
or U1654 (N_1654,In_2545,In_2183);
or U1655 (N_1655,In_135,In_2895);
and U1656 (N_1656,In_1398,In_270);
nand U1657 (N_1657,In_1728,In_3281);
nand U1658 (N_1658,In_782,In_4577);
and U1659 (N_1659,In_4019,In_4645);
and U1660 (N_1660,In_2448,In_64);
nor U1661 (N_1661,In_2912,In_4239);
and U1662 (N_1662,In_4102,In_4564);
and U1663 (N_1663,In_844,In_2980);
nand U1664 (N_1664,In_1637,In_3458);
and U1665 (N_1665,In_1043,In_4622);
nor U1666 (N_1666,In_3941,In_27);
or U1667 (N_1667,In_4774,In_4219);
and U1668 (N_1668,In_2514,In_4291);
nor U1669 (N_1669,In_1395,In_4500);
and U1670 (N_1670,In_269,In_589);
nand U1671 (N_1671,In_2181,In_791);
nand U1672 (N_1672,In_4533,In_2615);
nand U1673 (N_1673,In_1725,In_2349);
nand U1674 (N_1674,In_568,In_1095);
xor U1675 (N_1675,In_2267,In_3986);
nand U1676 (N_1676,In_4281,In_2732);
nand U1677 (N_1677,In_2859,In_933);
xor U1678 (N_1678,In_910,In_4269);
xnor U1679 (N_1679,In_1242,In_1309);
and U1680 (N_1680,In_3632,In_160);
nor U1681 (N_1681,In_1936,In_4273);
or U1682 (N_1682,In_3868,In_2536);
nor U1683 (N_1683,In_2783,In_4620);
or U1684 (N_1684,In_2593,In_4195);
xor U1685 (N_1685,In_200,In_2370);
nor U1686 (N_1686,In_2707,In_517);
and U1687 (N_1687,In_2939,In_3036);
or U1688 (N_1688,In_3532,In_1343);
nand U1689 (N_1689,In_3739,In_4470);
xnor U1690 (N_1690,In_3615,In_404);
nand U1691 (N_1691,In_1560,In_815);
nor U1692 (N_1692,In_3230,In_335);
nand U1693 (N_1693,In_3477,In_4342);
or U1694 (N_1694,In_2384,In_4238);
and U1695 (N_1695,In_3551,In_125);
nand U1696 (N_1696,In_632,In_2382);
xor U1697 (N_1697,In_4598,In_3206);
or U1698 (N_1698,In_2338,In_2598);
or U1699 (N_1699,In_4514,In_669);
or U1700 (N_1700,In_3679,In_3979);
and U1701 (N_1701,In_4630,In_740);
or U1702 (N_1702,In_1747,In_2167);
xnor U1703 (N_1703,In_226,In_3759);
nor U1704 (N_1704,In_2891,In_1540);
and U1705 (N_1705,In_4869,In_1984);
or U1706 (N_1706,In_1172,In_1237);
nand U1707 (N_1707,In_2904,In_4646);
or U1708 (N_1708,In_3697,In_242);
nand U1709 (N_1709,In_545,In_3420);
nor U1710 (N_1710,In_3698,In_4072);
or U1711 (N_1711,In_1722,In_2524);
nor U1712 (N_1712,In_3687,In_3141);
or U1713 (N_1713,In_4624,In_4552);
nand U1714 (N_1714,In_1575,In_2748);
or U1715 (N_1715,In_99,In_1481);
or U1716 (N_1716,In_4699,In_4387);
or U1717 (N_1717,In_4033,In_1124);
and U1718 (N_1718,In_3912,In_1093);
nand U1719 (N_1719,In_2139,In_4526);
nor U1720 (N_1720,In_482,In_1497);
xor U1721 (N_1721,In_789,In_3192);
nor U1722 (N_1722,In_4576,In_1774);
nand U1723 (N_1723,In_1145,In_3049);
nor U1724 (N_1724,In_1522,In_2605);
and U1725 (N_1725,In_2955,In_3765);
and U1726 (N_1726,In_4402,In_3480);
or U1727 (N_1727,In_4437,In_4782);
and U1728 (N_1728,In_2275,In_4004);
nor U1729 (N_1729,In_2470,In_797);
nand U1730 (N_1730,In_4111,In_313);
and U1731 (N_1731,In_1041,In_1569);
or U1732 (N_1732,In_1499,In_4980);
nand U1733 (N_1733,In_3555,In_2577);
nor U1734 (N_1734,In_1000,In_4290);
or U1735 (N_1735,In_4206,In_2475);
nor U1736 (N_1736,In_757,In_3855);
nor U1737 (N_1737,In_4285,In_2901);
and U1738 (N_1738,In_386,In_1016);
and U1739 (N_1739,In_2134,In_2906);
or U1740 (N_1740,In_1555,In_3468);
or U1741 (N_1741,In_635,In_2132);
and U1742 (N_1742,In_2361,In_3975);
nand U1743 (N_1743,In_449,In_2340);
or U1744 (N_1744,In_966,In_1664);
nand U1745 (N_1745,In_3048,In_171);
or U1746 (N_1746,In_4070,In_4659);
nand U1747 (N_1747,In_4876,In_339);
nor U1748 (N_1748,In_1641,In_4045);
or U1749 (N_1749,In_4312,In_3363);
nor U1750 (N_1750,In_3736,In_4689);
nor U1751 (N_1751,In_819,In_1101);
nor U1752 (N_1752,In_2029,In_2652);
nand U1753 (N_1753,In_3423,In_2399);
or U1754 (N_1754,In_1426,In_1063);
or U1755 (N_1755,In_4827,In_762);
nor U1756 (N_1756,In_3641,In_1450);
and U1757 (N_1757,In_505,In_2459);
and U1758 (N_1758,In_4811,In_4462);
or U1759 (N_1759,In_4898,In_443);
nand U1760 (N_1760,In_3802,In_3757);
and U1761 (N_1761,In_4002,In_2383);
and U1762 (N_1762,In_1083,In_628);
nor U1763 (N_1763,In_1052,In_2085);
xnor U1764 (N_1764,In_2086,In_4867);
nor U1765 (N_1765,In_4568,In_1058);
and U1766 (N_1766,In_723,In_4120);
xnor U1767 (N_1767,In_4784,In_2453);
nor U1768 (N_1768,In_3753,In_372);
nand U1769 (N_1769,In_4508,In_1968);
nand U1770 (N_1770,In_1278,In_975);
xor U1771 (N_1771,In_4095,In_4501);
or U1772 (N_1772,In_1632,In_476);
nand U1773 (N_1773,In_1983,In_4202);
nand U1774 (N_1774,In_1388,In_2247);
nand U1775 (N_1775,In_215,In_3645);
xor U1776 (N_1776,In_1217,In_4839);
and U1777 (N_1777,In_98,In_110);
and U1778 (N_1778,In_3217,In_919);
nand U1779 (N_1779,In_4567,In_621);
nor U1780 (N_1780,In_357,In_3092);
nor U1781 (N_1781,In_3180,In_1105);
and U1782 (N_1782,In_2304,In_29);
nand U1783 (N_1783,In_3793,In_4600);
and U1784 (N_1784,In_1545,In_4765);
and U1785 (N_1785,In_119,In_395);
nand U1786 (N_1786,In_232,In_4725);
or U1787 (N_1787,In_828,In_2558);
or U1788 (N_1788,In_778,In_425);
and U1789 (N_1789,In_3067,In_3305);
and U1790 (N_1790,In_2556,In_3805);
and U1791 (N_1791,In_1505,In_1552);
nand U1792 (N_1792,In_787,In_3510);
nor U1793 (N_1793,In_3253,In_4428);
nand U1794 (N_1794,In_927,In_2597);
nor U1795 (N_1795,In_3321,In_3125);
nor U1796 (N_1796,In_2402,In_2179);
nor U1797 (N_1797,In_3688,In_2164);
or U1798 (N_1798,In_798,In_2696);
xor U1799 (N_1799,In_3090,In_2909);
and U1800 (N_1800,In_3292,In_2753);
nand U1801 (N_1801,In_2319,In_4753);
or U1802 (N_1802,In_4103,In_1571);
or U1803 (N_1803,In_4734,In_19);
or U1804 (N_1804,In_1310,In_3993);
and U1805 (N_1805,In_4650,In_946);
and U1806 (N_1806,In_3685,In_1972);
xor U1807 (N_1807,In_698,In_642);
nor U1808 (N_1808,In_3822,In_2900);
nor U1809 (N_1809,In_479,In_2922);
nor U1810 (N_1810,In_1926,In_126);
xnor U1811 (N_1811,In_3634,In_1068);
nor U1812 (N_1812,In_1005,In_818);
nor U1813 (N_1813,In_1897,In_897);
nor U1814 (N_1814,In_3172,In_272);
or U1815 (N_1815,In_3498,In_4259);
nor U1816 (N_1816,In_4327,In_4895);
nand U1817 (N_1817,In_1091,In_4152);
nand U1818 (N_1818,In_4951,In_2238);
and U1819 (N_1819,In_4265,In_4013);
and U1820 (N_1820,In_4623,In_3622);
nor U1821 (N_1821,In_2612,In_4041);
nor U1822 (N_1822,In_4221,In_1125);
nor U1823 (N_1823,In_3093,In_3859);
or U1824 (N_1824,In_2863,In_2578);
nand U1825 (N_1825,In_629,In_3644);
or U1826 (N_1826,In_378,In_1974);
nor U1827 (N_1827,In_1989,In_2008);
nor U1828 (N_1828,In_4271,In_1570);
nor U1829 (N_1829,In_2345,In_1609);
and U1830 (N_1830,In_3828,In_1711);
or U1831 (N_1831,In_4550,In_3919);
or U1832 (N_1832,In_3074,In_1493);
xor U1833 (N_1833,In_1567,In_94);
nor U1834 (N_1834,In_1684,In_1402);
nor U1835 (N_1835,In_887,In_53);
nor U1836 (N_1836,In_4488,In_2317);
and U1837 (N_1837,In_1046,In_70);
nand U1838 (N_1838,In_530,In_1559);
nor U1839 (N_1839,In_773,In_1817);
nor U1840 (N_1840,In_942,In_259);
nand U1841 (N_1841,In_2751,In_1165);
or U1842 (N_1842,In_3572,In_4247);
nor U1843 (N_1843,In_4887,In_106);
xor U1844 (N_1844,In_279,In_4132);
nor U1845 (N_1845,In_2166,In_4485);
xor U1846 (N_1846,In_4961,In_1274);
or U1847 (N_1847,In_4936,In_251);
nor U1848 (N_1848,In_970,In_4396);
or U1849 (N_1849,In_2393,In_4381);
nor U1850 (N_1850,In_1490,In_1502);
xor U1851 (N_1851,In_4003,In_1553);
nand U1852 (N_1852,In_2675,In_4804);
nor U1853 (N_1853,In_587,In_2820);
nor U1854 (N_1854,In_2687,In_923);
and U1855 (N_1855,In_2620,In_3343);
nand U1856 (N_1856,In_4707,In_3001);
or U1857 (N_1857,In_3252,In_1320);
nand U1858 (N_1858,In_3949,In_576);
nor U1859 (N_1859,In_82,In_2076);
nor U1860 (N_1860,In_945,In_1485);
nor U1861 (N_1861,In_1970,In_4915);
nand U1862 (N_1862,In_2398,In_4523);
nand U1863 (N_1863,In_4190,In_1668);
xnor U1864 (N_1864,In_201,In_4975);
nand U1865 (N_1865,In_2530,In_1207);
nand U1866 (N_1866,In_504,In_2274);
nor U1867 (N_1867,In_1819,In_300);
nand U1868 (N_1868,In_4435,In_4854);
nand U1869 (N_1869,In_604,In_3684);
and U1870 (N_1870,In_2741,In_1036);
nor U1871 (N_1871,In_3129,In_151);
nand U1872 (N_1872,In_4101,In_2657);
and U1873 (N_1873,In_764,In_1054);
or U1874 (N_1874,In_2312,In_4211);
nand U1875 (N_1875,In_3346,In_940);
or U1876 (N_1876,In_2233,In_1170);
nand U1877 (N_1877,In_4878,In_3302);
nand U1878 (N_1878,In_4394,In_4229);
nand U1879 (N_1879,In_4467,In_4988);
and U1880 (N_1880,In_2555,In_4016);
nor U1881 (N_1881,In_8,In_3514);
nor U1882 (N_1882,In_2659,In_3280);
and U1883 (N_1883,In_2135,In_742);
nor U1884 (N_1884,In_3248,In_1244);
nor U1885 (N_1885,In_1018,In_801);
and U1886 (N_1886,In_2595,In_1995);
or U1887 (N_1887,In_1252,In_2188);
nand U1888 (N_1888,In_613,In_2305);
nand U1889 (N_1889,In_3604,In_671);
nand U1890 (N_1890,In_983,In_2099);
and U1891 (N_1891,In_1736,In_2329);
xor U1892 (N_1892,In_3926,In_2435);
nand U1893 (N_1893,In_809,In_956);
nor U1894 (N_1894,In_1892,In_1526);
and U1895 (N_1895,In_2232,In_2948);
nor U1896 (N_1896,In_3109,In_1595);
and U1897 (N_1897,In_1611,In_1185);
nor U1898 (N_1898,In_3387,In_2746);
and U1899 (N_1899,In_4305,In_1232);
and U1900 (N_1900,In_518,In_5);
xnor U1901 (N_1901,In_149,In_4461);
nand U1902 (N_1902,In_4079,In_4297);
nand U1903 (N_1903,In_1378,In_4424);
nand U1904 (N_1904,In_3490,In_1385);
xnor U1905 (N_1905,In_2517,In_1886);
nand U1906 (N_1906,In_3255,In_3466);
nand U1907 (N_1907,In_1219,In_124);
and U1908 (N_1908,In_375,In_113);
nand U1909 (N_1909,In_30,In_284);
nand U1910 (N_1910,In_3015,In_3353);
nor U1911 (N_1911,In_4192,In_1901);
nor U1912 (N_1912,In_2363,In_1131);
or U1913 (N_1913,In_2411,In_2376);
nand U1914 (N_1914,In_2324,In_1374);
or U1915 (N_1915,In_2890,In_351);
and U1916 (N_1916,In_3720,In_521);
xor U1917 (N_1917,In_4896,In_2454);
and U1918 (N_1918,In_1614,In_1348);
or U1919 (N_1919,In_874,In_2367);
or U1920 (N_1920,In_1832,In_3424);
nand U1921 (N_1921,In_2601,In_3409);
nand U1922 (N_1922,In_4726,In_4885);
and U1923 (N_1923,In_2456,In_2129);
nor U1924 (N_1924,In_1973,In_3915);
nor U1925 (N_1925,In_525,In_1775);
or U1926 (N_1926,In_3875,In_1880);
nand U1927 (N_1927,In_4830,In_3976);
or U1928 (N_1928,In_1928,In_325);
xor U1929 (N_1929,In_4955,In_3798);
or U1930 (N_1930,In_2278,In_4048);
nor U1931 (N_1931,In_676,In_4307);
and U1932 (N_1932,In_2588,In_4756);
and U1933 (N_1933,In_2511,In_3194);
nor U1934 (N_1934,In_2740,In_4858);
and U1935 (N_1935,In_680,In_649);
nor U1936 (N_1936,In_591,In_231);
or U1937 (N_1937,In_360,In_1406);
nor U1938 (N_1938,In_662,In_3637);
and U1939 (N_1939,In_1104,In_776);
or U1940 (N_1940,In_2342,In_537);
nor U1941 (N_1941,In_1798,In_513);
and U1942 (N_1942,In_4109,In_139);
or U1943 (N_1943,In_1925,In_413);
or U1944 (N_1944,In_4448,In_1342);
or U1945 (N_1945,In_1543,In_1666);
nand U1946 (N_1946,In_741,In_4986);
nor U1947 (N_1947,In_1898,In_3057);
or U1948 (N_1948,In_4685,In_688);
nand U1949 (N_1949,In_2644,In_1012);
and U1950 (N_1950,In_3165,In_1931);
xnor U1951 (N_1951,In_1824,In_2092);
and U1952 (N_1952,In_2663,In_614);
nand U1953 (N_1953,In_1102,In_914);
nand U1954 (N_1954,In_1757,In_4167);
nand U1955 (N_1955,In_3227,In_2226);
nor U1956 (N_1956,In_968,In_2563);
nor U1957 (N_1957,In_50,In_1203);
nor U1958 (N_1958,In_1510,In_4432);
xor U1959 (N_1959,In_2921,In_243);
or U1960 (N_1960,In_301,In_2184);
or U1961 (N_1961,In_634,In_4089);
or U1962 (N_1962,In_264,In_111);
and U1963 (N_1963,In_918,In_4881);
or U1964 (N_1964,In_1710,In_4632);
nor U1965 (N_1965,In_2033,In_1228);
xnor U1966 (N_1966,In_2176,In_461);
nor U1967 (N_1967,In_857,In_4578);
and U1968 (N_1968,In_4603,In_3335);
and U1969 (N_1969,In_2256,In_163);
nor U1970 (N_1970,In_4397,In_2512);
nand U1971 (N_1971,In_369,In_1959);
and U1972 (N_1972,In_3834,In_4842);
and U1973 (N_1973,In_285,In_2153);
nor U1974 (N_1974,In_2311,In_4071);
nand U1975 (N_1975,In_2717,In_1626);
nand U1976 (N_1976,In_1040,In_1057);
nor U1977 (N_1977,In_2155,In_4894);
nor U1978 (N_1978,In_3322,In_2347);
or U1979 (N_1979,In_16,In_2808);
nand U1980 (N_1980,In_2843,In_1602);
and U1981 (N_1981,In_1539,In_2991);
nor U1982 (N_1982,In_4717,In_3586);
and U1983 (N_1983,In_2940,In_2394);
or U1984 (N_1984,In_724,In_4156);
nor U1985 (N_1985,In_774,In_2528);
and U1986 (N_1986,In_3867,In_1644);
nand U1987 (N_1987,In_4494,In_1353);
and U1988 (N_1988,In_4474,In_1245);
or U1989 (N_1989,In_1963,In_734);
nand U1990 (N_1990,In_4032,In_1676);
or U1991 (N_1991,In_2287,In_1417);
nand U1992 (N_1992,In_4930,In_2206);
nand U1993 (N_1993,In_4503,In_1340);
xor U1994 (N_1994,In_611,In_1834);
xnor U1995 (N_1995,In_1267,In_2713);
and U1996 (N_1996,In_3425,In_4379);
nor U1997 (N_1997,In_2272,In_3787);
xnor U1998 (N_1998,In_356,In_4829);
or U1999 (N_1999,In_2366,In_1108);
nand U2000 (N_2000,In_4966,In_3020);
nor U2001 (N_2001,In_1748,In_2330);
and U2002 (N_2002,In_4452,In_1727);
or U2003 (N_2003,In_153,In_1126);
nand U2004 (N_2004,In_156,In_1263);
nand U2005 (N_2005,In_969,In_363);
and U2006 (N_2006,In_55,In_4357);
or U2007 (N_2007,In_4570,In_612);
nor U2008 (N_2008,In_1822,In_1854);
or U2009 (N_2009,In_4721,In_1392);
or U2010 (N_2010,In_2424,In_3103);
and U2011 (N_2011,In_2090,In_3237);
nand U2012 (N_2012,In_466,In_1140);
xnor U2013 (N_2013,In_4868,In_3176);
and U2014 (N_2014,In_1302,In_4362);
or U2015 (N_2015,In_1238,In_2819);
nand U2016 (N_2016,In_1113,In_2529);
and U2017 (N_2017,In_935,In_4519);
or U2018 (N_2018,In_76,In_4263);
xor U2019 (N_2019,In_1447,In_2271);
xnor U2020 (N_2020,In_1477,In_441);
nand U2021 (N_2021,In_3916,In_1315);
or U2022 (N_2022,In_2801,In_2911);
or U2023 (N_2023,In_4948,In_3754);
nor U2024 (N_2024,In_1333,In_766);
nand U2025 (N_2025,In_1218,In_689);
xnor U2026 (N_2026,In_908,In_2219);
and U2027 (N_2027,In_650,In_4310);
nand U2028 (N_2028,In_991,In_2277);
nor U2029 (N_2029,In_2993,In_3732);
nor U2030 (N_2030,In_3642,In_455);
nand U2031 (N_2031,In_327,In_3102);
and U2032 (N_2032,In_886,In_2567);
or U2033 (N_2033,In_2480,In_3737);
nand U2034 (N_2034,In_1407,In_1662);
nor U2035 (N_2035,In_3463,In_3564);
nor U2036 (N_2036,In_1297,In_520);
and U2037 (N_2037,In_2007,In_2013);
xnor U2038 (N_2038,In_1239,In_834);
nand U2039 (N_2039,In_3994,In_3402);
xnor U2040 (N_2040,In_2225,In_432);
nand U2041 (N_2041,In_295,In_293);
xor U2042 (N_2042,In_4797,In_661);
and U2043 (N_2043,In_352,In_3512);
and U2044 (N_2044,In_2493,In_3995);
nor U2045 (N_2045,In_2918,In_1888);
nor U2046 (N_2046,In_727,In_440);
xor U2047 (N_2047,In_2654,In_3880);
and U2048 (N_2048,In_1895,In_1962);
nand U2049 (N_2049,In_4619,In_2785);
xor U2050 (N_2050,In_3507,In_1590);
nor U2051 (N_2051,In_3185,In_3476);
and U2052 (N_2052,In_4810,In_1066);
nand U2053 (N_2053,In_1598,In_3282);
nand U2054 (N_2054,In_2719,In_128);
and U2055 (N_2055,In_3984,In_4547);
nand U2056 (N_2056,In_1358,In_2855);
or U2057 (N_2057,In_1199,In_1288);
and U2058 (N_2058,In_3668,In_1894);
or U2059 (N_2059,In_1699,In_2847);
nand U2060 (N_2060,In_2771,In_359);
or U2061 (N_2061,In_1061,In_4757);
nor U2062 (N_2062,In_186,In_463);
or U2063 (N_2063,In_2151,In_4532);
or U2064 (N_2064,In_1106,In_1752);
nor U2065 (N_2065,In_4216,In_1866);
nand U2066 (N_2066,In_1211,In_239);
or U2067 (N_2067,In_478,In_3610);
nand U2068 (N_2068,In_3546,In_1672);
and U2069 (N_2069,In_4535,In_1141);
xor U2070 (N_2070,In_1149,In_1867);
nand U2071 (N_2071,In_696,In_1255);
or U2072 (N_2072,In_2498,In_4926);
nor U2073 (N_2073,In_3911,In_4166);
and U2074 (N_2074,In_4083,In_790);
nor U2075 (N_2075,In_993,In_1321);
nor U2076 (N_2076,In_2723,In_3938);
and U2077 (N_2077,In_2609,In_1956);
xnor U2078 (N_2078,In_4302,In_4416);
nor U2079 (N_2079,In_2727,In_3607);
nor U2080 (N_2080,In_22,In_3881);
and U2081 (N_2081,In_1780,In_3427);
and U2082 (N_2082,In_268,In_577);
nor U2083 (N_2083,In_2813,In_4704);
xor U2084 (N_2084,In_1969,In_3406);
and U2085 (N_2085,In_321,In_324);
nor U2086 (N_2086,In_3552,In_1448);
or U2087 (N_2087,In_1026,In_298);
nor U2088 (N_2088,In_4335,In_4524);
nor U2089 (N_2089,In_78,In_1115);
and U2090 (N_2090,In_2285,In_1463);
nand U2091 (N_2091,In_380,In_1979);
or U2092 (N_2092,In_4791,In_1758);
and U2093 (N_2093,In_4292,In_605);
nor U2094 (N_2094,In_1247,In_1281);
nand U2095 (N_2095,In_4483,In_2428);
or U2096 (N_2096,In_1879,In_1135);
nor U2097 (N_2097,In_2581,In_2842);
nand U2098 (N_2098,In_685,In_1640);
nand U2099 (N_2099,In_4656,In_1103);
nor U2100 (N_2100,In_91,In_2660);
nand U2101 (N_2101,In_1977,In_2364);
or U2102 (N_2102,In_3380,In_3315);
nand U2103 (N_2103,In_4338,In_1373);
nor U2104 (N_2104,In_4051,In_1948);
nand U2105 (N_2105,In_4353,In_960);
nor U2106 (N_2106,In_4341,In_1673);
or U2107 (N_2107,In_4,In_1813);
and U2108 (N_2108,In_3054,In_2302);
nand U2109 (N_2109,In_4793,In_3028);
and U2110 (N_2110,In_4225,In_853);
nor U2111 (N_2111,In_217,In_2845);
nor U2112 (N_2112,In_3484,In_794);
nor U2113 (N_2113,In_3126,In_4148);
nor U2114 (N_2114,In_2631,In_2755);
or U2115 (N_2115,In_4178,In_4597);
nor U2116 (N_2116,In_2323,In_3324);
nor U2117 (N_2117,In_154,In_3729);
xor U2118 (N_2118,In_822,In_2509);
and U2119 (N_2119,In_4453,In_1158);
xor U2120 (N_2120,In_705,In_4693);
and U2121 (N_2121,In_4069,In_2375);
nor U2122 (N_2122,In_2481,In_3395);
nand U2123 (N_2123,In_4972,In_2941);
nand U2124 (N_2124,In_2273,In_2284);
nor U2125 (N_2125,In_1890,In_772);
xor U2126 (N_2126,In_3815,In_1805);
or U2127 (N_2127,In_3447,In_2440);
nand U2128 (N_2128,In_312,In_3189);
nor U2129 (N_2129,In_2590,In_2124);
or U2130 (N_2130,In_4314,In_700);
or U2131 (N_2131,In_3702,In_1534);
nand U2132 (N_2132,In_3157,In_4672);
xor U2133 (N_2133,In_1260,In_2938);
nand U2134 (N_2134,In_1344,In_3633);
nor U2135 (N_2135,In_4595,In_2818);
nand U2136 (N_2136,In_101,In_4479);
nor U2137 (N_2137,In_2280,In_2385);
nand U2138 (N_2138,In_1318,In_3603);
or U2139 (N_2139,In_4931,In_1157);
or U2140 (N_2140,In_1980,In_2298);
or U2141 (N_2141,In_2208,In_1588);
nand U2142 (N_2142,In_2889,In_470);
or U2143 (N_2143,In_3760,In_1200);
or U2144 (N_2144,In_4883,In_3251);
or U2145 (N_2145,In_1079,In_715);
nor U2146 (N_2146,In_1601,In_4164);
nor U2147 (N_2147,In_4426,In_4114);
and U2148 (N_2148,In_719,In_2081);
or U2149 (N_2149,In_4377,In_4914);
nand U2150 (N_2150,In_1619,In_1675);
nand U2151 (N_2151,In_3543,In_4200);
nand U2152 (N_2152,In_1,In_4617);
and U2153 (N_2153,In_96,In_4486);
nor U2154 (N_2154,In_3151,In_2627);
nor U2155 (N_2155,In_973,In_75);
nand U2156 (N_2156,In_1638,In_4207);
and U2157 (N_2157,In_4864,In_1308);
xor U2158 (N_2158,In_1954,In_2902);
nand U2159 (N_2159,In_4924,In_4695);
nor U2160 (N_2160,In_3857,In_1949);
nor U2161 (N_2161,In_673,In_2195);
nand U2162 (N_2162,In_4078,In_1784);
nand U2163 (N_2163,In_1596,In_988);
nor U2164 (N_2164,In_3416,In_2626);
and U2165 (N_2165,In_3132,In_652);
nand U2166 (N_2166,In_1300,In_581);
nor U2167 (N_2167,In_1060,In_4832);
and U2168 (N_2168,In_2423,In_814);
or U2169 (N_2169,In_1618,In_3205);
and U2170 (N_2170,In_1860,In_2389);
and U2171 (N_2171,In_4143,In_2169);
nor U2172 (N_2172,In_1210,In_176);
nand U2173 (N_2173,In_3100,In_3032);
and U2174 (N_2174,In_4615,In_247);
xor U2175 (N_2175,In_759,In_1801);
nor U2176 (N_2176,In_3014,In_1151);
and U2177 (N_2177,In_3840,In_69);
nand U2178 (N_2178,In_1810,In_4245);
nand U2179 (N_2179,In_2079,In_1617);
xor U2180 (N_2180,In_323,In_2446);
nand U2181 (N_2181,In_1878,In_3593);
nand U2182 (N_2182,In_4803,In_59);
nor U2183 (N_2183,In_3823,In_3216);
or U2184 (N_2184,In_4727,In_1648);
nor U2185 (N_2185,In_45,In_3091);
and U2186 (N_2186,In_4237,In_350);
or U2187 (N_2187,In_3223,In_4060);
nor U2188 (N_2188,In_1122,In_1473);
and U2189 (N_2189,In_2130,In_4475);
nor U2190 (N_2190,In_3418,In_3045);
nor U2191 (N_2191,In_2410,In_1589);
xor U2192 (N_2192,In_1487,In_3595);
nand U2193 (N_2193,In_3382,In_3455);
and U2194 (N_2194,In_2778,In_4847);
xor U2195 (N_2195,In_588,In_1223);
nand U2196 (N_2196,In_133,In_3909);
nand U2197 (N_2197,In_2670,In_3400);
xnor U2198 (N_2198,In_275,In_2750);
nor U2199 (N_2199,In_2763,In_353);
xnor U2200 (N_2200,In_1951,In_43);
and U2201 (N_2201,In_1337,In_1616);
nor U2202 (N_2202,In_2775,In_2354);
xor U2203 (N_2203,In_2913,In_3188);
or U2204 (N_2204,In_4732,In_422);
and U2205 (N_2205,In_3159,In_1934);
nor U2206 (N_2206,In_2883,In_4891);
nand U2207 (N_2207,In_4879,In_2137);
or U2208 (N_2208,In_3077,In_2412);
nor U2209 (N_2209,In_1440,In_3008);
nand U2210 (N_2210,In_3098,In_3144);
xor U2211 (N_2211,In_2321,In_4715);
nor U2212 (N_2212,In_3374,In_3407);
xnor U2213 (N_2213,In_371,In_1745);
and U2214 (N_2214,In_3886,In_2781);
nor U2215 (N_2215,In_1421,In_3721);
and U2216 (N_2216,In_3111,In_1193);
nand U2217 (N_2217,In_1965,In_3553);
and U2218 (N_2218,In_1690,In_681);
nor U2219 (N_2219,In_450,In_1904);
or U2220 (N_2220,In_4231,In_4950);
and U2221 (N_2221,In_659,In_3123);
or U2222 (N_2222,In_3608,In_1971);
nand U2223 (N_2223,In_1729,In_2193);
xnor U2224 (N_2224,In_3584,In_2163);
and U2225 (N_2225,In_1700,In_1441);
xor U2226 (N_2226,In_1705,In_1741);
and U2227 (N_2227,In_2328,In_1622);
and U2228 (N_2228,In_4365,In_4999);
or U2229 (N_2229,In_3770,In_699);
nand U2230 (N_2230,In_1541,In_1412);
xor U2231 (N_2231,In_454,In_4511);
and U2232 (N_2232,In_1518,In_826);
nand U2233 (N_2233,In_4953,In_1159);
nor U2234 (N_2234,In_138,In_3580);
or U2235 (N_2235,In_185,In_2966);
nand U2236 (N_2236,In_483,In_1514);
nand U2237 (N_2237,In_793,In_3244);
nor U2238 (N_2238,In_4311,In_1967);
or U2239 (N_2239,In_903,In_1064);
and U2240 (N_2240,In_3467,In_861);
or U2241 (N_2241,In_2229,In_1354);
or U2242 (N_2242,In_1472,In_2253);
xor U2243 (N_2243,In_4778,In_4464);
xor U2244 (N_2244,In_2568,In_4807);
and U2245 (N_2245,In_660,In_3567);
and U2246 (N_2246,In_4050,In_2988);
nor U2247 (N_2247,In_3347,In_1578);
nand U2248 (N_2248,In_10,In_2881);
nor U2249 (N_2249,In_1011,In_3229);
nand U2250 (N_2250,In_2162,In_627);
nand U2251 (N_2251,In_1413,In_1837);
nor U2252 (N_2252,In_66,In_720);
nor U2253 (N_2253,In_407,In_2421);
and U2254 (N_2254,In_4430,In_544);
xnor U2255 (N_2255,In_2355,In_2542);
nand U2256 (N_2256,In_3107,In_4097);
nand U2257 (N_2257,In_3686,In_607);
and U2258 (N_2258,In_3657,In_539);
nand U2259 (N_2259,In_1529,In_452);
nor U2260 (N_2260,In_636,In_1415);
and U2261 (N_2261,In_3969,In_1277);
and U2262 (N_2262,In_4515,In_626);
and U2263 (N_2263,In_2401,In_2821);
nor U2264 (N_2264,In_1403,In_1336);
nor U2265 (N_2265,In_4489,In_2217);
or U2266 (N_2266,In_944,In_1661);
and U2267 (N_2267,In_777,In_4593);
nand U2268 (N_2268,In_398,In_390);
nor U2269 (N_2269,In_4675,In_1845);
nand U2270 (N_2270,In_420,In_4256);
xnor U2271 (N_2271,In_3565,In_1023);
and U2272 (N_2272,In_56,In_1429);
and U2273 (N_2273,In_4421,In_4965);
or U2274 (N_2274,In_1078,In_3652);
nor U2275 (N_2275,In_4026,In_2531);
nand U2276 (N_2276,In_4491,In_214);
and U2277 (N_2277,In_3961,In_1746);
or U2278 (N_2278,In_1978,In_998);
or U2279 (N_2279,In_1791,In_1738);
or U2280 (N_2280,In_3182,In_1220);
and U2281 (N_2281,In_3627,In_643);
xor U2282 (N_2282,In_1153,In_73);
nand U2283 (N_2283,In_2686,In_690);
nor U2284 (N_2284,In_2316,In_645);
nand U2285 (N_2285,In_3140,In_3075);
nand U2286 (N_2286,In_3334,In_33);
xor U2287 (N_2287,In_130,In_2444);
nand U2288 (N_2288,In_4172,In_1850);
nand U2289 (N_2289,In_3841,In_4901);
nand U2290 (N_2290,In_4250,In_4283);
nand U2291 (N_2291,In_3939,In_2817);
xnor U2292 (N_2292,In_1387,In_4088);
nand U2293 (N_2293,In_4175,In_2281);
or U2294 (N_2294,In_2488,In_795);
nand U2295 (N_2295,In_1305,In_68);
or U2296 (N_2296,In_3848,In_1436);
xor U2297 (N_2297,In_3905,In_572);
and U2298 (N_2298,In_458,In_2021);
and U2299 (N_2299,In_4354,In_2623);
nand U2300 (N_2300,In_385,In_546);
nor U2301 (N_2301,In_831,In_4029);
nand U2302 (N_2302,In_274,In_4912);
nand U2303 (N_2303,In_161,In_2738);
and U2304 (N_2304,In_2887,In_4750);
or U2305 (N_2305,In_267,In_4590);
and U2306 (N_2306,In_3833,In_1331);
or U2307 (N_2307,In_1548,In_3486);
nand U2308 (N_2308,In_4946,In_1830);
or U2309 (N_2309,In_3991,In_3187);
nor U2310 (N_2310,In_1907,In_1537);
or U2311 (N_2311,In_986,In_292);
and U2312 (N_2312,In_3945,In_3681);
xnor U2313 (N_2313,In_3327,In_609);
nor U2314 (N_2314,In_4490,In_3341);
and U2315 (N_2315,In_4798,In_3952);
nor U2316 (N_2316,In_2569,In_4686);
or U2317 (N_2317,In_4388,In_2004);
or U2318 (N_2318,In_3824,In_415);
nand U2319 (N_2319,In_4035,In_2069);
nor U2320 (N_2320,In_1006,In_3935);
and U2321 (N_2321,In_2037,In_2816);
nand U2322 (N_2322,In_1055,In_3167);
nand U2323 (N_2323,In_2291,In_3853);
or U2324 (N_2324,In_2610,In_845);
or U2325 (N_2325,In_2978,In_3879);
or U2326 (N_2326,In_3957,In_4825);
nor U2327 (N_2327,In_4170,In_2051);
nor U2328 (N_2328,In_1351,In_2613);
nor U2329 (N_2329,In_655,In_2234);
nor U2330 (N_2330,In_1349,In_1828);
nand U2331 (N_2331,In_4249,In_672);
nand U2332 (N_2332,In_2754,In_4024);
nor U2333 (N_2333,In_4989,In_850);
nor U2334 (N_2334,In_3908,In_2468);
nand U2335 (N_2335,In_2562,In_408);
nand U2336 (N_2336,In_4610,In_4436);
or U2337 (N_2337,In_1991,In_4520);
and U2338 (N_2338,In_4399,In_3338);
or U2339 (N_2339,In_4815,In_1241);
or U2340 (N_2340,In_4058,In_4851);
and U2341 (N_2341,In_2506,In_2288);
nor U2342 (N_2342,In_2925,In_1530);
or U2343 (N_2343,In_610,In_24);
or U2344 (N_2344,In_3914,In_3152);
nor U2345 (N_2345,In_1209,In_3019);
or U2346 (N_2346,In_693,In_2968);
xnor U2347 (N_2347,In_3328,In_1760);
nand U2348 (N_2348,In_1816,In_4802);
xnor U2349 (N_2349,In_2045,In_2074);
and U2350 (N_2350,In_236,In_2856);
nor U2351 (N_2351,In_877,In_4352);
nor U2352 (N_2352,In_4641,In_382);
xor U2353 (N_2353,In_1004,In_2237);
or U2354 (N_2354,In_3947,In_1397);
xnor U2355 (N_2355,In_868,In_2908);
nand U2356 (N_2356,In_1455,In_710);
and U2357 (N_2357,In_2113,In_4151);
xnor U2358 (N_2358,In_1279,In_4299);
and U2359 (N_2359,In_1367,In_1523);
and U2360 (N_2360,In_4716,In_3095);
nand U2361 (N_2361,In_2811,In_3156);
or U2362 (N_2362,In_2209,In_3542);
nand U2363 (N_2363,In_4180,In_2942);
nand U2364 (N_2364,In_3925,In_3296);
xor U2365 (N_2365,In_1788,In_3257);
nand U2366 (N_2366,In_2969,In_1524);
nand U2367 (N_2367,In_3433,In_147);
and U2368 (N_2368,In_3771,In_3332);
nand U2369 (N_2369,In_2027,In_4422);
or U2370 (N_2370,In_4012,In_4933);
or U2371 (N_2371,In_1835,In_3768);
xnor U2372 (N_2372,In_4589,In_3789);
and U2373 (N_2373,In_4272,In_3956);
nor U2374 (N_2374,In_4662,In_428);
and U2375 (N_2375,In_4049,In_1671);
and U2376 (N_2376,In_838,In_3457);
or U2377 (N_2377,In_1074,In_4884);
and U2378 (N_2378,In_3215,In_2293);
nand U2379 (N_2379,In_4468,In_2715);
and U2380 (N_2380,In_847,In_2722);
and U2381 (N_2381,In_1538,In_4417);
or U2382 (N_2382,In_1803,In_165);
nand U2383 (N_2383,In_906,In_2852);
nor U2384 (N_2384,In_4262,In_524);
nand U2385 (N_2385,In_1484,In_4469);
and U2386 (N_2386,In_2026,In_3743);
nand U2387 (N_2387,In_4142,In_2048);
xnor U2388 (N_2388,In_2279,In_4718);
nor U2389 (N_2389,In_2507,In_1603);
and U2390 (N_2390,In_3359,In_3437);
nor U2391 (N_2391,In_550,In_1513);
and U2392 (N_2392,In_2767,In_3331);
or U2393 (N_2393,In_4538,In_0);
or U2394 (N_2394,In_4649,In_4517);
or U2395 (N_2395,In_1905,In_3659);
nor U2396 (N_2396,In_4964,In_2380);
nor U2397 (N_2397,In_2477,In_1044);
or U2398 (N_2398,In_2830,In_336);
nor U2399 (N_2399,In_3112,In_3707);
nand U2400 (N_2400,In_1280,In_4587);
xor U2401 (N_2401,In_3169,In_3160);
and U2402 (N_2402,In_4667,In_2136);
and U2403 (N_2403,In_2676,In_571);
nor U2404 (N_2404,In_3812,In_938);
nor U2405 (N_2405,In_2214,In_4037);
and U2406 (N_2406,In_2525,In_3233);
nor U2407 (N_2407,In_2541,In_3055);
or U2408 (N_2408,In_2122,In_3773);
nand U2409 (N_2409,In_1357,In_4147);
nor U2410 (N_2410,In_3830,In_4009);
nand U2411 (N_2411,In_3002,In_3432);
and U2412 (N_2412,In_1261,In_2523);
nor U2413 (N_2413,In_1146,In_2059);
and U2414 (N_2414,In_1446,In_3794);
nand U2415 (N_2415,In_2794,In_162);
nor U2416 (N_2416,In_864,In_2886);
or U2417 (N_2417,In_4945,In_1646);
and U2418 (N_2418,In_552,In_1855);
nor U2419 (N_2419,In_3669,In_1035);
or U2420 (N_2420,In_3025,In_3254);
nor U2421 (N_2421,In_221,In_4456);
nor U2422 (N_2422,In_4772,In_480);
or U2423 (N_2423,In_2527,In_1874);
nor U2424 (N_2424,In_1304,In_2194);
and U2425 (N_2425,In_4637,In_141);
nor U2426 (N_2426,In_3803,In_2407);
nand U2427 (N_2427,In_3262,In_52);
nand U2428 (N_2428,In_666,In_3816);
nand U2429 (N_2429,In_832,In_3470);
nor U2430 (N_2430,In_2337,In_1282);
nand U2431 (N_2431,In_3536,In_3444);
nand U2432 (N_2432,In_1597,In_2070);
and U2433 (N_2433,In_816,In_4614);
nand U2434 (N_2434,In_3269,In_4763);
or U2435 (N_2435,In_4255,In_2972);
nor U2436 (N_2436,In_2431,In_361);
and U2437 (N_2437,In_4848,In_1702);
xor U2438 (N_2438,In_4006,In_1677);
nand U2439 (N_2439,In_2420,In_4162);
or U2440 (N_2440,In_2266,In_2088);
and U2441 (N_2441,In_1073,In_3445);
or U2442 (N_2442,In_1292,In_3097);
nand U2443 (N_2443,In_1818,In_560);
nor U2444 (N_2444,In_4020,In_1384);
xnor U2445 (N_2445,In_4749,In_558);
or U2446 (N_2446,In_1442,In_3258);
or U2447 (N_2447,In_4226,In_2585);
and U2448 (N_2448,In_177,In_3027);
or U2449 (N_2449,In_4849,In_1119);
nand U2450 (N_2450,In_4374,In_108);
or U2451 (N_2451,In_2294,In_1547);
xnor U2452 (N_2452,In_1183,In_2802);
and U2453 (N_2453,In_3903,In_3483);
or U2454 (N_2454,In_4588,In_3515);
and U2455 (N_2455,In_2866,In_3731);
nor U2456 (N_2456,In_2764,In_4744);
nand U2457 (N_2457,In_2831,In_658);
nand U2458 (N_2458,In_4873,In_977);
nor U2459 (N_2459,In_1606,In_364);
and U2460 (N_2460,In_1825,In_1283);
nor U2461 (N_2461,In_4639,In_1111);
or U2462 (N_2462,In_1256,In_2216);
and U2463 (N_2463,In_4760,In_4571);
nand U2464 (N_2464,In_4406,In_3790);
or U2465 (N_2465,In_4661,In_2602);
nor U2466 (N_2466,In_261,In_3210);
and U2467 (N_2467,In_338,In_393);
and U2468 (N_2468,In_4733,In_2834);
nor U2469 (N_2469,In_4108,In_2297);
or U2470 (N_2470,In_1437,In_2264);
or U2471 (N_2471,In_379,In_820);
nor U2472 (N_2472,In_1189,In_533);
xor U2473 (N_2473,In_875,In_1383);
nand U2474 (N_2474,In_1162,In_3010);
and U2475 (N_2475,In_709,In_4821);
or U2476 (N_2476,In_2954,In_4561);
and U2477 (N_2477,In_1913,In_2736);
nand U2478 (N_2478,In_496,In_3161);
and U2479 (N_2479,In_4087,In_4344);
or U2480 (N_2480,In_2471,In_1168);
nor U2481 (N_2481,In_2919,In_405);
nor U2482 (N_2482,In_4493,In_624);
and U2483 (N_2483,In_1511,In_2549);
nand U2484 (N_2484,In_4459,In_465);
or U2485 (N_2485,In_725,In_2548);
nor U2486 (N_2486,In_3700,In_3190);
or U2487 (N_2487,In_2313,In_1922);
nand U2488 (N_2488,In_4266,In_1932);
nand U2489 (N_2489,In_2397,In_3998);
nor U2490 (N_2490,In_871,In_3068);
nor U2491 (N_2491,In_1909,In_3087);
nor U2492 (N_2492,In_88,In_1175);
nand U2493 (N_2493,In_4994,In_3628);
and U2494 (N_2494,In_2551,In_4860);
xor U2495 (N_2495,In_3290,In_2269);
nor U2496 (N_2496,In_879,In_4320);
and U2497 (N_2497,In_4496,In_3146);
nand U2498 (N_2498,In_3701,In_4007);
or U2499 (N_2499,In_4441,In_691);
nor U2500 (N_2500,N_369,N_868);
nand U2501 (N_2501,N_965,N_653);
nor U2502 (N_2502,N_1127,N_713);
nor U2503 (N_2503,N_399,N_549);
nand U2504 (N_2504,N_154,N_792);
and U2505 (N_2505,N_547,N_1178);
or U2506 (N_2506,N_633,N_1889);
or U2507 (N_2507,N_53,N_2317);
xor U2508 (N_2508,N_1129,N_473);
nor U2509 (N_2509,N_1985,N_1232);
and U2510 (N_2510,N_1528,N_1631);
or U2511 (N_2511,N_854,N_1080);
nor U2512 (N_2512,N_1262,N_1122);
and U2513 (N_2513,N_1871,N_680);
xnor U2514 (N_2514,N_367,N_2297);
nand U2515 (N_2515,N_173,N_102);
or U2516 (N_2516,N_1425,N_1869);
xor U2517 (N_2517,N_614,N_2199);
nor U2518 (N_2518,N_2254,N_1035);
and U2519 (N_2519,N_2218,N_1656);
and U2520 (N_2520,N_1848,N_483);
nand U2521 (N_2521,N_246,N_2001);
or U2522 (N_2522,N_419,N_1926);
nand U2523 (N_2523,N_1841,N_2164);
or U2524 (N_2524,N_708,N_2315);
nand U2525 (N_2525,N_615,N_2337);
nor U2526 (N_2526,N_685,N_801);
and U2527 (N_2527,N_272,N_1521);
xor U2528 (N_2528,N_822,N_668);
nor U2529 (N_2529,N_1752,N_502);
nor U2530 (N_2530,N_412,N_2324);
or U2531 (N_2531,N_1518,N_2059);
nand U2532 (N_2532,N_392,N_2040);
nor U2533 (N_2533,N_247,N_2197);
or U2534 (N_2534,N_1316,N_103);
or U2535 (N_2535,N_266,N_1517);
nand U2536 (N_2536,N_212,N_370);
xor U2537 (N_2537,N_1246,N_1384);
and U2538 (N_2538,N_1060,N_2122);
nand U2539 (N_2539,N_1797,N_1074);
and U2540 (N_2540,N_1005,N_787);
xor U2541 (N_2541,N_990,N_2290);
nor U2542 (N_2542,N_1540,N_703);
or U2543 (N_2543,N_1857,N_887);
nor U2544 (N_2544,N_1557,N_1744);
nand U2545 (N_2545,N_448,N_1583);
nor U2546 (N_2546,N_1390,N_136);
or U2547 (N_2547,N_1681,N_962);
nand U2548 (N_2548,N_955,N_2364);
nand U2549 (N_2549,N_996,N_881);
or U2550 (N_2550,N_979,N_749);
xor U2551 (N_2551,N_357,N_2163);
xor U2552 (N_2552,N_1921,N_984);
and U2553 (N_2553,N_1382,N_640);
nor U2554 (N_2554,N_1929,N_500);
nand U2555 (N_2555,N_1514,N_1441);
xnor U2556 (N_2556,N_960,N_111);
or U2557 (N_2557,N_735,N_494);
and U2558 (N_2558,N_31,N_1864);
and U2559 (N_2559,N_675,N_1312);
and U2560 (N_2560,N_2416,N_2434);
nand U2561 (N_2561,N_1131,N_1628);
and U2562 (N_2562,N_159,N_1618);
nor U2563 (N_2563,N_181,N_991);
or U2564 (N_2564,N_446,N_1894);
nand U2565 (N_2565,N_645,N_1507);
nor U2566 (N_2566,N_1571,N_402);
and U2567 (N_2567,N_175,N_1135);
or U2568 (N_2568,N_2081,N_1655);
nor U2569 (N_2569,N_967,N_332);
nand U2570 (N_2570,N_145,N_1039);
or U2571 (N_2571,N_2128,N_626);
or U2572 (N_2572,N_1919,N_882);
nand U2573 (N_2573,N_1481,N_211);
nand U2574 (N_2574,N_835,N_38);
and U2575 (N_2575,N_24,N_1022);
nand U2576 (N_2576,N_2497,N_742);
xnor U2577 (N_2577,N_436,N_993);
or U2578 (N_2578,N_647,N_1118);
nor U2579 (N_2579,N_1643,N_527);
nand U2580 (N_2580,N_1335,N_216);
and U2581 (N_2581,N_2390,N_805);
nor U2582 (N_2582,N_1215,N_1363);
or U2583 (N_2583,N_2339,N_1527);
and U2584 (N_2584,N_2430,N_2212);
nand U2585 (N_2585,N_852,N_2272);
or U2586 (N_2586,N_699,N_312);
nand U2587 (N_2587,N_1466,N_1368);
or U2588 (N_2588,N_1908,N_586);
xor U2589 (N_2589,N_1463,N_660);
or U2590 (N_2590,N_893,N_1066);
nor U2591 (N_2591,N_2155,N_1480);
or U2592 (N_2592,N_404,N_1069);
and U2593 (N_2593,N_521,N_1222);
or U2594 (N_2594,N_1397,N_936);
or U2595 (N_2595,N_2241,N_2151);
nand U2596 (N_2596,N_1907,N_2093);
nand U2597 (N_2597,N_2246,N_330);
nor U2598 (N_2598,N_2381,N_926);
or U2599 (N_2599,N_550,N_1096);
nor U2600 (N_2600,N_1373,N_2257);
or U2601 (N_2601,N_1298,N_2002);
nand U2602 (N_2602,N_375,N_23);
and U2603 (N_2603,N_1257,N_2355);
or U2604 (N_2604,N_652,N_2062);
nand U2605 (N_2605,N_802,N_1966);
and U2606 (N_2606,N_1709,N_520);
nand U2607 (N_2607,N_2423,N_1145);
or U2608 (N_2608,N_426,N_771);
nand U2609 (N_2609,N_2432,N_978);
and U2610 (N_2610,N_2113,N_463);
nand U2611 (N_2611,N_1151,N_1489);
xnor U2612 (N_2612,N_2465,N_1449);
and U2613 (N_2613,N_1189,N_226);
and U2614 (N_2614,N_661,N_1959);
and U2615 (N_2615,N_982,N_1564);
nor U2616 (N_2616,N_309,N_1333);
nor U2617 (N_2617,N_1522,N_543);
or U2618 (N_2618,N_621,N_331);
nor U2619 (N_2619,N_761,N_2094);
and U2620 (N_2620,N_276,N_78);
nand U2621 (N_2621,N_1467,N_46);
nor U2622 (N_2622,N_2368,N_1679);
nor U2623 (N_2623,N_200,N_1324);
nand U2624 (N_2624,N_1206,N_409);
nor U2625 (N_2625,N_166,N_488);
or U2626 (N_2626,N_1544,N_1295);
or U2627 (N_2627,N_1904,N_149);
or U2628 (N_2628,N_684,N_908);
nand U2629 (N_2629,N_1745,N_2316);
or U2630 (N_2630,N_29,N_1284);
and U2631 (N_2631,N_485,N_1834);
and U2632 (N_2632,N_766,N_1399);
xor U2633 (N_2633,N_1599,N_1837);
and U2634 (N_2634,N_1370,N_2276);
or U2635 (N_2635,N_1386,N_162);
or U2636 (N_2636,N_1121,N_2278);
xnor U2637 (N_2637,N_96,N_2284);
xnor U2638 (N_2638,N_2130,N_658);
or U2639 (N_2639,N_1357,N_806);
nand U2640 (N_2640,N_511,N_1148);
or U2641 (N_2641,N_2038,N_1468);
and U2642 (N_2642,N_254,N_119);
and U2643 (N_2643,N_1100,N_837);
and U2644 (N_2644,N_124,N_731);
or U2645 (N_2645,N_566,N_1790);
and U2646 (N_2646,N_476,N_880);
and U2647 (N_2647,N_465,N_380);
and U2648 (N_2648,N_503,N_1851);
or U2649 (N_2649,N_314,N_2024);
nand U2650 (N_2650,N_2189,N_751);
or U2651 (N_2651,N_1808,N_2017);
nor U2652 (N_2652,N_2314,N_2240);
nand U2653 (N_2653,N_2137,N_1850);
and U2654 (N_2654,N_1041,N_1856);
nor U2655 (N_2655,N_1349,N_1102);
nand U2656 (N_2656,N_1670,N_2484);
xnor U2657 (N_2657,N_1058,N_800);
nand U2658 (N_2658,N_113,N_363);
and U2659 (N_2659,N_1590,N_146);
and U2660 (N_2660,N_2150,N_552);
nand U2661 (N_2661,N_2154,N_2344);
nor U2662 (N_2662,N_1120,N_1139);
nor U2663 (N_2663,N_84,N_2449);
or U2664 (N_2664,N_2329,N_1219);
or U2665 (N_2665,N_1007,N_2299);
or U2666 (N_2666,N_1561,N_657);
nand U2667 (N_2667,N_1493,N_637);
or U2668 (N_2668,N_359,N_1054);
or U2669 (N_2669,N_1989,N_1811);
and U2670 (N_2670,N_321,N_864);
nand U2671 (N_2671,N_1645,N_1037);
nor U2672 (N_2672,N_1799,N_831);
or U2673 (N_2673,N_1830,N_2363);
nor U2674 (N_2674,N_1824,N_395);
or U2675 (N_2675,N_894,N_1296);
and U2676 (N_2676,N_580,N_2296);
xor U2677 (N_2677,N_407,N_1233);
xor U2678 (N_2678,N_946,N_2331);
xnor U2679 (N_2679,N_1347,N_1827);
nor U2680 (N_2680,N_2082,N_885);
xor U2681 (N_2681,N_1785,N_811);
nor U2682 (N_2682,N_1412,N_1482);
or U2683 (N_2683,N_904,N_1710);
nand U2684 (N_2684,N_1696,N_760);
or U2685 (N_2685,N_1458,N_1520);
or U2686 (N_2686,N_1912,N_773);
or U2687 (N_2687,N_1265,N_160);
nand U2688 (N_2688,N_293,N_745);
or U2689 (N_2689,N_1692,N_758);
nand U2690 (N_2690,N_1146,N_459);
xnor U2691 (N_2691,N_1541,N_720);
nand U2692 (N_2692,N_2016,N_1423);
nor U2693 (N_2693,N_423,N_1061);
and U2694 (N_2694,N_1340,N_50);
or U2695 (N_2695,N_2348,N_943);
and U2696 (N_2696,N_1393,N_1539);
and U2697 (N_2697,N_1472,N_2275);
nand U2698 (N_2698,N_539,N_2020);
xnor U2699 (N_2699,N_2459,N_1565);
or U2700 (N_2700,N_1,N_693);
nor U2701 (N_2701,N_232,N_1933);
nand U2702 (N_2702,N_1968,N_1275);
or U2703 (N_2703,N_1250,N_2424);
nand U2704 (N_2704,N_2209,N_2034);
xnor U2705 (N_2705,N_651,N_2433);
and U2706 (N_2706,N_1748,N_2260);
or U2707 (N_2707,N_1923,N_910);
and U2708 (N_2708,N_1334,N_1801);
nand U2709 (N_2709,N_836,N_1276);
or U2710 (N_2710,N_611,N_1639);
nand U2711 (N_2711,N_1981,N_1582);
nor U2712 (N_2712,N_1868,N_2345);
nor U2713 (N_2713,N_1789,N_902);
or U2714 (N_2714,N_2277,N_1788);
xor U2715 (N_2715,N_1636,N_1164);
nand U2716 (N_2716,N_1762,N_2469);
nand U2717 (N_2717,N_1784,N_451);
nand U2718 (N_2718,N_1453,N_1107);
nand U2719 (N_2719,N_1070,N_183);
nand U2720 (N_2720,N_1754,N_1380);
xor U2721 (N_2721,N_1549,N_1516);
nand U2722 (N_2722,N_1918,N_1686);
or U2723 (N_2723,N_1558,N_1783);
or U2724 (N_2724,N_1095,N_403);
or U2725 (N_2725,N_2148,N_1792);
nand U2726 (N_2726,N_378,N_1619);
nand U2727 (N_2727,N_2055,N_1154);
nand U2728 (N_2728,N_1137,N_320);
or U2729 (N_2729,N_487,N_1053);
nand U2730 (N_2730,N_1421,N_2412);
and U2731 (N_2731,N_340,N_772);
or U2732 (N_2732,N_1717,N_525);
or U2733 (N_2733,N_2050,N_1820);
or U2734 (N_2734,N_2443,N_980);
and U2735 (N_2735,N_1774,N_1722);
or U2736 (N_2736,N_2415,N_1727);
or U2737 (N_2737,N_439,N_2077);
nor U2738 (N_2738,N_2420,N_790);
or U2739 (N_2739,N_873,N_1730);
and U2740 (N_2740,N_2255,N_1640);
xnor U2741 (N_2741,N_182,N_1050);
nand U2742 (N_2742,N_2258,N_889);
and U2743 (N_2743,N_1360,N_1875);
nand U2744 (N_2744,N_415,N_1601);
nand U2745 (N_2745,N_351,N_923);
or U2746 (N_2746,N_347,N_1251);
and U2747 (N_2747,N_1647,N_2398);
nor U2748 (N_2748,N_1555,N_1141);
xnor U2749 (N_2749,N_1461,N_2223);
and U2750 (N_2750,N_1270,N_2162);
nor U2751 (N_2751,N_767,N_2244);
nand U2752 (N_2752,N_10,N_2392);
or U2753 (N_2753,N_1642,N_1064);
nor U2754 (N_2754,N_623,N_1993);
and U2755 (N_2755,N_1934,N_1683);
and U2756 (N_2756,N_1142,N_917);
or U2757 (N_2757,N_2338,N_780);
nand U2758 (N_2758,N_757,N_2140);
nand U2759 (N_2759,N_1881,N_275);
and U2760 (N_2760,N_1883,N_1248);
and U2761 (N_2761,N_892,N_1462);
xnor U2762 (N_2762,N_755,N_1650);
and U2763 (N_2763,N_405,N_737);
and U2764 (N_2764,N_1411,N_519);
and U2765 (N_2765,N_695,N_2441);
or U2766 (N_2766,N_2084,N_2108);
nand U2767 (N_2767,N_1828,N_2044);
or U2768 (N_2768,N_215,N_42);
nand U2769 (N_2769,N_1214,N_1318);
and U2770 (N_2770,N_2326,N_1088);
and U2771 (N_2771,N_952,N_76);
xor U2772 (N_2772,N_15,N_2396);
and U2773 (N_2773,N_895,N_1117);
nand U2774 (N_2774,N_915,N_2190);
nand U2775 (N_2775,N_1330,N_2228);
nor U2776 (N_2776,N_2295,N_1773);
and U2777 (N_2777,N_2468,N_849);
and U2778 (N_2778,N_155,N_1627);
nor U2779 (N_2779,N_1017,N_471);
and U2780 (N_2780,N_1303,N_1982);
and U2781 (N_2781,N_1254,N_21);
and U2782 (N_2782,N_1367,N_1537);
nand U2783 (N_2783,N_2135,N_1546);
nor U2784 (N_2784,N_1470,N_663);
nor U2785 (N_2785,N_1417,N_925);
or U2786 (N_2786,N_2173,N_206);
nand U2787 (N_2787,N_1159,N_1319);
nor U2788 (N_2788,N_2032,N_1615);
nand U2789 (N_2789,N_573,N_168);
nor U2790 (N_2790,N_1798,N_1484);
and U2791 (N_2791,N_2175,N_945);
nand U2792 (N_2792,N_1304,N_1720);
nor U2793 (N_2793,N_909,N_214);
and U2794 (N_2794,N_788,N_401);
and U2795 (N_2795,N_1289,N_1294);
or U2796 (N_2796,N_1906,N_798);
xnor U2797 (N_2797,N_605,N_1193);
nor U2798 (N_2798,N_956,N_1306);
nand U2799 (N_2799,N_752,N_1003);
nor U2800 (N_2800,N_365,N_2259);
xor U2801 (N_2801,N_1542,N_2131);
and U2802 (N_2802,N_466,N_1910);
nand U2803 (N_2803,N_1769,N_877);
and U2804 (N_2804,N_1735,N_1002);
nor U2805 (N_2805,N_607,N_1173);
or U2806 (N_2806,N_1958,N_826);
or U2807 (N_2807,N_2047,N_1332);
nor U2808 (N_2808,N_1731,N_1280);
and U2809 (N_2809,N_2022,N_2426);
nor U2810 (N_2810,N_1937,N_932);
and U2811 (N_2811,N_44,N_66);
nand U2812 (N_2812,N_1536,N_2336);
nor U2813 (N_2813,N_432,N_165);
or U2814 (N_2814,N_128,N_32);
nor U2815 (N_2815,N_1447,N_2053);
xor U2816 (N_2816,N_1573,N_2357);
and U2817 (N_2817,N_638,N_1274);
nor U2818 (N_2818,N_2090,N_507);
or U2819 (N_2819,N_1305,N_944);
xnor U2820 (N_2820,N_1728,N_548);
nand U2821 (N_2821,N_1707,N_2429);
xor U2822 (N_2822,N_112,N_736);
or U2823 (N_2823,N_1751,N_1814);
or U2824 (N_2824,N_1526,N_2442);
nand U2825 (N_2825,N_1006,N_1014);
nor U2826 (N_2826,N_475,N_931);
nand U2827 (N_2827,N_793,N_1817);
nor U2828 (N_2828,N_2180,N_271);
nor U2829 (N_2829,N_510,N_2365);
nor U2830 (N_2830,N_1607,N_461);
or U2831 (N_2831,N_1551,N_914);
nor U2832 (N_2832,N_366,N_2097);
nand U2833 (N_2833,N_1048,N_949);
nor U2834 (N_2834,N_568,N_273);
and U2835 (N_2835,N_947,N_495);
nand U2836 (N_2836,N_1580,N_784);
and U2837 (N_2837,N_2498,N_1713);
or U2838 (N_2838,N_1403,N_744);
nand U2839 (N_2839,N_844,N_1083);
xnor U2840 (N_2840,N_334,N_1108);
or U2841 (N_2841,N_1322,N_851);
or U2842 (N_2842,N_863,N_2306);
nand U2843 (N_2843,N_995,N_1201);
nand U2844 (N_2844,N_1140,N_2116);
nor U2845 (N_2845,N_2205,N_2021);
and U2846 (N_2846,N_2438,N_1922);
xor U2847 (N_2847,N_37,N_2192);
nand U2848 (N_2848,N_1073,N_491);
and U2849 (N_2849,N_1896,N_1682);
nor U2850 (N_2850,N_1778,N_1622);
nor U2851 (N_2851,N_185,N_1554);
or U2852 (N_2852,N_498,N_299);
and U2853 (N_2853,N_1396,N_1635);
nand U2854 (N_2854,N_2011,N_408);
nor U2855 (N_2855,N_144,N_1478);
xor U2856 (N_2856,N_928,N_427);
or U2857 (N_2857,N_542,N_1550);
xnor U2858 (N_2858,N_900,N_1202);
or U2859 (N_2859,N_2267,N_1266);
or U2860 (N_2860,N_105,N_939);
nor U2861 (N_2861,N_2301,N_1569);
xnor U2862 (N_2862,N_1822,N_2005);
or U2863 (N_2863,N_2168,N_676);
or U2864 (N_2864,N_65,N_164);
or U2865 (N_2865,N_1990,N_1758);
and U2866 (N_2866,N_1766,N_558);
nor U2867 (N_2867,N_286,N_729);
nand U2868 (N_2868,N_2031,N_1946);
xnor U2869 (N_2869,N_472,N_1132);
nor U2870 (N_2870,N_1701,N_2101);
nand U2871 (N_2871,N_830,N_1459);
xnor U2872 (N_2872,N_2298,N_861);
or U2873 (N_2873,N_1414,N_1043);
or U2874 (N_2874,N_1895,N_1690);
nor U2875 (N_2875,N_17,N_1870);
nor U2876 (N_2876,N_819,N_445);
nand U2877 (N_2877,N_61,N_222);
nand U2878 (N_2878,N_1415,N_1589);
or U2879 (N_2879,N_786,N_1809);
and U2880 (N_2880,N_1000,N_267);
or U2881 (N_2881,N_1501,N_1950);
or U2882 (N_2882,N_1729,N_2479);
xor U2883 (N_2883,N_816,N_2169);
nor U2884 (N_2884,N_493,N_2076);
nor U2885 (N_2885,N_2346,N_1740);
nand U2886 (N_2886,N_1314,N_1917);
or U2887 (N_2887,N_135,N_2211);
and U2888 (N_2888,N_1733,N_346);
and U2889 (N_2889,N_1283,N_610);
nand U2890 (N_2890,N_686,N_2000);
nor U2891 (N_2891,N_1849,N_39);
nor U2892 (N_2892,N_1113,N_783);
xnor U2893 (N_2893,N_177,N_1882);
and U2894 (N_2894,N_462,N_1757);
nor U2895 (N_2895,N_2233,N_1974);
and U2896 (N_2896,N_1831,N_655);
nand U2897 (N_2897,N_217,N_237);
or U2898 (N_2898,N_170,N_2353);
and U2899 (N_2899,N_875,N_479);
xnor U2900 (N_2900,N_297,N_1302);
or U2901 (N_2901,N_2461,N_284);
nor U2902 (N_2902,N_1535,N_1287);
and U2903 (N_2903,N_1358,N_2405);
xor U2904 (N_2904,N_2437,N_1604);
nor U2905 (N_2905,N_509,N_2333);
nand U2906 (N_2906,N_935,N_2492);
and U2907 (N_2907,N_1153,N_782);
or U2908 (N_2908,N_577,N_1225);
and U2909 (N_2909,N_1742,N_1955);
and U2910 (N_2910,N_2487,N_616);
nand U2911 (N_2911,N_1719,N_328);
nand U2912 (N_2912,N_1644,N_2418);
nor U2913 (N_2913,N_253,N_2321);
and U2914 (N_2914,N_1477,N_1229);
or U2915 (N_2915,N_1374,N_517);
nor U2916 (N_2916,N_514,N_1515);
and U2917 (N_2917,N_1559,N_1782);
and U2918 (N_2918,N_1339,N_1512);
nor U2919 (N_2919,N_2366,N_2351);
and U2920 (N_2920,N_1174,N_1285);
and U2921 (N_2921,N_213,N_2170);
xor U2922 (N_2922,N_189,N_624);
and U2923 (N_2923,N_1629,N_799);
nor U2924 (N_2924,N_424,N_474);
nand U2925 (N_2925,N_1965,N_1805);
or U2926 (N_2926,N_2273,N_2120);
nor U2927 (N_2927,N_1443,N_360);
or U2928 (N_2928,N_1715,N_2400);
or U2929 (N_2929,N_690,N_163);
or U2930 (N_2930,N_184,N_564);
or U2931 (N_2931,N_1588,N_977);
nand U2932 (N_2932,N_2358,N_678);
xnor U2933 (N_2933,N_1260,N_1957);
and U2934 (N_2934,N_2499,N_838);
or U2935 (N_2935,N_1490,N_188);
xnor U2936 (N_2936,N_1962,N_1829);
and U2937 (N_2937,N_1776,N_1323);
or U2938 (N_2938,N_1042,N_1085);
and U2939 (N_2939,N_1099,N_2136);
or U2940 (N_2940,N_1420,N_418);
and U2941 (N_2941,N_234,N_1136);
nor U2942 (N_2942,N_282,N_1091);
xnor U2943 (N_2943,N_2323,N_1366);
or U2944 (N_2944,N_1503,N_1847);
or U2945 (N_2945,N_323,N_2349);
xnor U2946 (N_2946,N_1927,N_264);
nor U2947 (N_2947,N_345,N_906);
and U2948 (N_2948,N_594,N_2171);
and U2949 (N_2949,N_508,N_1359);
or U2950 (N_2950,N_2203,N_2312);
xor U2951 (N_2951,N_381,N_879);
nor U2952 (N_2952,N_1637,N_724);
xnor U2953 (N_2953,N_385,N_174);
nand U2954 (N_2954,N_422,N_2256);
nand U2955 (N_2955,N_1658,N_911);
nor U2956 (N_2956,N_1065,N_1577);
nor U2957 (N_2957,N_1903,N_921);
nor U2958 (N_2958,N_1273,N_809);
or U2959 (N_2959,N_719,N_1218);
nor U2960 (N_2960,N_707,N_492);
and U2961 (N_2961,N_571,N_2279);
nor U2962 (N_2962,N_301,N_95);
and U2963 (N_2963,N_827,N_1413);
or U2964 (N_2964,N_171,N_1823);
xor U2965 (N_2965,N_248,N_1175);
and U2966 (N_2966,N_2280,N_1878);
nand U2967 (N_2967,N_1613,N_538);
or U2968 (N_2968,N_1077,N_478);
or U2969 (N_2969,N_523,N_628);
nand U2970 (N_2970,N_2019,N_901);
nor U2971 (N_2971,N_1694,N_1068);
and U2972 (N_2972,N_2393,N_2340);
nor U2973 (N_2973,N_748,N_1353);
or U2974 (N_2974,N_1992,N_64);
nand U2975 (N_2975,N_1021,N_2453);
and U2976 (N_2976,N_537,N_172);
or U2977 (N_2977,N_1932,N_57);
nand U2978 (N_2978,N_1446,N_1891);
and U2979 (N_2979,N_350,N_705);
and U2980 (N_2980,N_1749,N_966);
nand U2981 (N_2981,N_2253,N_1672);
nand U2982 (N_2982,N_2379,N_36);
nand U2983 (N_2983,N_964,N_27);
nand U2984 (N_2984,N_1125,N_1630);
nor U2985 (N_2985,N_1854,N_1369);
or U2986 (N_2986,N_1452,N_2086);
nand U2987 (N_2987,N_438,N_1269);
nor U2988 (N_2988,N_1736,N_2114);
and U2989 (N_2989,N_1646,N_1237);
nand U2990 (N_2990,N_1874,N_2251);
or U2991 (N_2991,N_2036,N_1506);
xor U2992 (N_2992,N_2206,N_2404);
or U2993 (N_2993,N_698,N_1034);
or U2994 (N_2994,N_515,N_20);
nor U2995 (N_2995,N_1952,N_1931);
and U2996 (N_2996,N_1935,N_1597);
xor U2997 (N_2997,N_130,N_1071);
nor U2998 (N_2998,N_296,N_954);
or U2999 (N_2999,N_2224,N_41);
nor U3000 (N_3000,N_1791,N_631);
nor U3001 (N_3001,N_2098,N_871);
and U3002 (N_3002,N_80,N_625);
or U3003 (N_3003,N_289,N_2185);
or U3004 (N_3004,N_143,N_1765);
and U3005 (N_3005,N_2134,N_230);
and U3006 (N_3006,N_2063,N_794);
or U3007 (N_3007,N_1388,N_795);
nor U3008 (N_3008,N_371,N_258);
and U3009 (N_3009,N_1450,N_1807);
nor U3010 (N_3010,N_641,N_1008);
and U3011 (N_3011,N_302,N_2475);
or U3012 (N_3012,N_721,N_2289);
and U3013 (N_3013,N_1133,N_1611);
nor U3014 (N_3014,N_988,N_1570);
and U3015 (N_3015,N_754,N_1530);
or U3016 (N_3016,N_1662,N_1612);
or U3017 (N_3017,N_1244,N_193);
nor U3018 (N_3018,N_516,N_1004);
or U3019 (N_3019,N_732,N_775);
nor U3020 (N_3020,N_1572,N_1325);
or U3021 (N_3021,N_1623,N_2425);
nand U3022 (N_3022,N_2250,N_87);
nor U3023 (N_3023,N_1479,N_2064);
nand U3024 (N_3024,N_1247,N_545);
xor U3025 (N_3025,N_897,N_191);
nand U3026 (N_3026,N_656,N_122);
nor U3027 (N_3027,N_1190,N_2325);
and U3028 (N_3028,N_1015,N_255);
or U3029 (N_3029,N_1885,N_14);
or U3030 (N_3030,N_2310,N_589);
xor U3031 (N_3031,N_2221,N_454);
nand U3032 (N_3032,N_131,N_239);
nor U3033 (N_3033,N_746,N_1652);
nand U3034 (N_3034,N_2422,N_828);
xnor U3035 (N_3035,N_1724,N_1264);
nand U3036 (N_3036,N_1231,N_1001);
xor U3037 (N_3037,N_1203,N_98);
or U3038 (N_3038,N_820,N_349);
xnor U3039 (N_3039,N_219,N_192);
xnor U3040 (N_3040,N_2308,N_1858);
nor U3041 (N_3041,N_2003,N_1212);
or U3042 (N_3042,N_630,N_56);
nand U3043 (N_3043,N_2352,N_1951);
or U3044 (N_3044,N_2490,N_2187);
and U3045 (N_3045,N_28,N_1812);
and U3046 (N_3046,N_575,N_595);
xor U3047 (N_3047,N_602,N_2225);
nor U3048 (N_3048,N_209,N_447);
and U3049 (N_3049,N_627,N_1046);
nand U3050 (N_3050,N_1156,N_2399);
and U3051 (N_3051,N_2145,N_1671);
and U3052 (N_3052,N_743,N_1143);
or U3053 (N_3053,N_1835,N_203);
and U3054 (N_3054,N_1897,N_1429);
and U3055 (N_3055,N_2285,N_1777);
and U3056 (N_3056,N_1106,N_1406);
nand U3057 (N_3057,N_654,N_1914);
nand U3058 (N_3058,N_2458,N_1497);
nand U3059 (N_3059,N_388,N_207);
nor U3060 (N_3060,N_2057,N_1691);
nor U3061 (N_3061,N_560,N_1608);
nand U3062 (N_3062,N_2166,N_74);
or U3063 (N_3063,N_1047,N_2200);
nor U3064 (N_3064,N_2219,N_156);
and U3065 (N_3065,N_1300,N_300);
and U3066 (N_3066,N_1693,N_389);
and U3067 (N_3067,N_1234,N_1451);
nand U3068 (N_3068,N_11,N_1547);
nor U3069 (N_3069,N_1726,N_1925);
or U3070 (N_3070,N_34,N_1031);
and U3071 (N_3071,N_1172,N_1855);
and U3072 (N_3072,N_343,N_2195);
and U3073 (N_3073,N_1045,N_298);
nand U3074 (N_3074,N_2119,N_763);
and U3075 (N_3075,N_778,N_672);
nand U3076 (N_3076,N_565,N_327);
nor U3077 (N_3077,N_1970,N_47);
and U3078 (N_3078,N_109,N_372);
nand U3079 (N_3079,N_992,N_1437);
nor U3080 (N_3080,N_1486,N_1416);
or U3081 (N_3081,N_726,N_903);
or U3082 (N_3082,N_1930,N_229);
and U3083 (N_3083,N_1796,N_1836);
or U3084 (N_3084,N_1702,N_2238);
xnor U3085 (N_3085,N_1948,N_2158);
nor U3086 (N_3086,N_1995,N_581);
nand U3087 (N_3087,N_1427,N_1346);
nor U3088 (N_3088,N_1391,N_1114);
nand U3089 (N_3089,N_2210,N_1400);
nand U3090 (N_3090,N_2350,N_1236);
nor U3091 (N_3091,N_142,N_985);
xnor U3092 (N_3092,N_2009,N_1097);
and U3093 (N_3093,N_1806,N_1695);
or U3094 (N_3094,N_634,N_2463);
and U3095 (N_3095,N_2447,N_1308);
or U3096 (N_3096,N_187,N_629);
nor U3097 (N_3097,N_2235,N_704);
and U3098 (N_3098,N_1119,N_240);
nor U3099 (N_3099,N_1401,N_1843);
xor U3100 (N_3100,N_386,N_1945);
nor U3101 (N_3101,N_1689,N_259);
or U3102 (N_3102,N_1315,N_152);
nand U3103 (N_3103,N_2471,N_1956);
nand U3104 (N_3104,N_919,N_1016);
nand U3105 (N_3105,N_1890,N_1879);
and U3106 (N_3106,N_662,N_2100);
nand U3107 (N_3107,N_2110,N_1152);
nand U3108 (N_3108,N_574,N_1505);
nand U3109 (N_3109,N_1431,N_1755);
nand U3110 (N_3110,N_218,N_148);
and U3111 (N_3111,N_1317,N_1772);
nand U3112 (N_3112,N_92,N_898);
nand U3113 (N_3113,N_1259,N_1055);
or U3114 (N_3114,N_712,N_941);
or U3115 (N_3115,N_6,N_1947);
nor U3116 (N_3116,N_1680,N_1424);
nor U3117 (N_3117,N_1243,N_829);
nor U3118 (N_3118,N_883,N_83);
and U3119 (N_3119,N_431,N_1130);
xnor U3120 (N_3120,N_5,N_591);
and U3121 (N_3121,N_1434,N_2035);
or U3122 (N_3122,N_1078,N_2269);
or U3123 (N_3123,N_1553,N_1086);
or U3124 (N_3124,N_1101,N_1158);
or U3125 (N_3125,N_556,N_700);
nor U3126 (N_3126,N_410,N_1110);
and U3127 (N_3127,N_2229,N_1936);
and U3128 (N_3128,N_823,N_133);
nor U3129 (N_3129,N_1389,N_1291);
or U3130 (N_3130,N_2079,N_768);
nand U3131 (N_3131,N_1861,N_603);
nand U3132 (N_3132,N_1012,N_998);
or U3133 (N_3133,N_82,N_1185);
nor U3134 (N_3134,N_1944,N_270);
nor U3135 (N_3135,N_303,N_2074);
nand U3136 (N_3136,N_669,N_541);
nor U3137 (N_3137,N_2474,N_570);
and U3138 (N_3138,N_2182,N_1737);
nand U3139 (N_3139,N_2141,N_257);
nand U3140 (N_3140,N_455,N_872);
nor U3141 (N_3141,N_1915,N_1093);
and U3142 (N_3142,N_311,N_1838);
xor U3143 (N_3143,N_1706,N_368);
nor U3144 (N_3144,N_118,N_406);
or U3145 (N_3145,N_1587,N_1586);
nor U3146 (N_3146,N_839,N_1029);
or U3147 (N_3147,N_938,N_1375);
nor U3148 (N_3148,N_1621,N_1703);
xor U3149 (N_3149,N_715,N_157);
nand U3150 (N_3150,N_948,N_1455);
or U3151 (N_3151,N_779,N_2291);
nand U3152 (N_3152,N_635,N_151);
and U3153 (N_3153,N_554,N_1938);
and U3154 (N_3154,N_529,N_862);
and U3155 (N_3155,N_1167,N_930);
or U3156 (N_3156,N_1999,N_147);
and U3157 (N_3157,N_63,N_1224);
and U3158 (N_3158,N_1928,N_116);
xnor U3159 (N_3159,N_1980,N_1240);
xnor U3160 (N_3160,N_1651,N_848);
nand U3161 (N_3161,N_2261,N_1892);
and U3162 (N_3162,N_2080,N_522);
nand U3163 (N_3163,N_694,N_45);
nand U3164 (N_3164,N_665,N_1460);
nor U3165 (N_3165,N_905,N_1753);
or U3166 (N_3166,N_2384,N_853);
nor U3167 (N_3167,N_709,N_878);
or U3168 (N_3168,N_382,N_920);
or U3169 (N_3169,N_1418,N_22);
or U3170 (N_3170,N_606,N_1433);
or U3171 (N_3171,N_2476,N_269);
or U3172 (N_3172,N_223,N_1529);
or U3173 (N_3173,N_2431,N_1973);
or U3174 (N_3174,N_813,N_1163);
nor U3175 (N_3175,N_2220,N_587);
nand U3176 (N_3176,N_356,N_1648);
and U3177 (N_3177,N_1770,N_1226);
or U3178 (N_3178,N_1560,N_2380);
nor U3179 (N_3179,N_869,N_1378);
and U3180 (N_3180,N_1103,N_2270);
and U3181 (N_3181,N_339,N_1972);
or U3182 (N_3182,N_961,N_1617);
nand U3183 (N_3183,N_1677,N_2477);
nand U3184 (N_3184,N_430,N_953);
or U3185 (N_3185,N_1723,N_1194);
nor U3186 (N_3186,N_1010,N_759);
or U3187 (N_3187,N_546,N_762);
nor U3188 (N_3188,N_2207,N_86);
and U3189 (N_3189,N_274,N_1469);
and U3190 (N_3190,N_2448,N_134);
and U3191 (N_3191,N_596,N_1448);
nand U3192 (N_3192,N_2049,N_983);
xor U3193 (N_3193,N_2309,N_536);
and U3194 (N_3194,N_1759,N_352);
xnor U3195 (N_3195,N_93,N_572);
nand U3196 (N_3196,N_158,N_482);
and U3197 (N_3197,N_534,N_197);
and U3198 (N_3198,N_1491,N_341);
nor U3199 (N_3199,N_858,N_3);
nor U3200 (N_3200,N_812,N_1354);
xor U3201 (N_3201,N_1839,N_1606);
xnor U3202 (N_3202,N_1768,N_1040);
or U3203 (N_3203,N_1013,N_1543);
nand U3204 (N_3204,N_1803,N_2320);
nor U3205 (N_3205,N_1435,N_71);
or U3206 (N_3206,N_876,N_989);
nor U3207 (N_3207,N_126,N_1059);
and U3208 (N_3208,N_2367,N_1750);
nor U3209 (N_3209,N_460,N_242);
and U3210 (N_3210,N_1997,N_644);
and U3211 (N_3211,N_1678,N_2347);
and U3212 (N_3212,N_2491,N_1057);
nor U3213 (N_3213,N_727,N_2004);
or U3214 (N_3214,N_2167,N_2191);
or U3215 (N_3215,N_1288,N_870);
or U3216 (N_3216,N_1439,N_121);
or U3217 (N_3217,N_2389,N_2071);
and U3218 (N_3218,N_1860,N_1258);
or U3219 (N_3219,N_2354,N_643);
nand U3220 (N_3220,N_781,N_60);
or U3221 (N_3221,N_530,N_1668);
nand U3222 (N_3222,N_927,N_1183);
nand U3223 (N_3223,N_1187,N_319);
and U3224 (N_3224,N_2413,N_2480);
xor U3225 (N_3225,N_1343,N_110);
and U3226 (N_3226,N_2450,N_88);
or U3227 (N_3227,N_2410,N_2010);
nor U3228 (N_3228,N_865,N_316);
or U3229 (N_3229,N_1379,N_723);
and U3230 (N_3230,N_2483,N_486);
and U3231 (N_3231,N_305,N_540);
nand U3232 (N_3232,N_1329,N_13);
and U3233 (N_3233,N_1221,N_1286);
nor U3234 (N_3234,N_1659,N_1741);
xor U3235 (N_3235,N_306,N_2237);
nand U3236 (N_3236,N_1819,N_860);
and U3237 (N_3237,N_1177,N_2362);
nand U3238 (N_3238,N_2159,N_942);
nor U3239 (N_3239,N_4,N_1495);
xor U3240 (N_3240,N_2439,N_1351);
nand U3241 (N_3241,N_2411,N_1780);
nor U3242 (N_3242,N_227,N_1634);
or U3243 (N_3243,N_692,N_2264);
nor U3244 (N_3244,N_1994,N_2294);
and U3245 (N_3245,N_1126,N_697);
or U3246 (N_3246,N_1939,N_533);
and U3247 (N_3247,N_292,N_959);
xnor U3248 (N_3248,N_1134,N_52);
nor U3249 (N_3249,N_2061,N_1591);
nand U3250 (N_3250,N_1653,N_1341);
nand U3251 (N_3251,N_54,N_186);
and U3252 (N_3252,N_2156,N_632);
nor U3253 (N_3253,N_1205,N_376);
nand U3254 (N_3254,N_1211,N_205);
or U3255 (N_3255,N_480,N_1673);
nand U3256 (N_3256,N_2401,N_1863);
nor U3257 (N_3257,N_1230,N_958);
or U3258 (N_3258,N_361,N_1523);
nor U3259 (N_3259,N_2066,N_358);
xor U3260 (N_3260,N_1407,N_2089);
or U3261 (N_3261,N_198,N_1649);
nor U3262 (N_3262,N_1969,N_1877);
nor U3263 (N_3263,N_1104,N_2153);
or U3264 (N_3264,N_470,N_288);
nor U3265 (N_3265,N_618,N_918);
and U3266 (N_3266,N_2012,N_1075);
nand U3267 (N_3267,N_1026,N_1853);
nor U3268 (N_3268,N_2193,N_2454);
nand U3269 (N_3269,N_557,N_2266);
or U3270 (N_3270,N_1872,N_2370);
nor U3271 (N_3271,N_1475,N_642);
nand U3272 (N_3272,N_1361,N_1685);
xnor U3273 (N_3273,N_814,N_457);
nor U3274 (N_3274,N_2455,N_1666);
or U3275 (N_3275,N_2496,N_1483);
and U3276 (N_3276,N_1616,N_1438);
nand U3277 (N_3277,N_2493,N_1504);
and U3278 (N_3278,N_987,N_2123);
nor U3279 (N_3279,N_2414,N_1781);
nor U3280 (N_3280,N_393,N_2092);
or U3281 (N_3281,N_1991,N_687);
and U3282 (N_3282,N_1348,N_807);
nor U3283 (N_3283,N_1337,N_924);
or U3284 (N_3284,N_416,N_2085);
nand U3285 (N_3285,N_562,N_2056);
or U3286 (N_3286,N_261,N_1198);
nor U3287 (N_3287,N_414,N_1816);
nor U3288 (N_3288,N_1840,N_1036);
nor U3289 (N_3289,N_1844,N_1893);
xor U3290 (N_3290,N_1128,N_664);
nand U3291 (N_3291,N_843,N_2106);
nand U3292 (N_3292,N_484,N_2428);
or U3293 (N_3293,N_1025,N_1700);
nand U3294 (N_3294,N_747,N_2014);
and U3295 (N_3295,N_344,N_2408);
nor U3296 (N_3296,N_313,N_2026);
or U3297 (N_3297,N_1665,N_429);
nand U3298 (N_3298,N_2341,N_1654);
xnor U3299 (N_3299,N_2360,N_391);
or U3300 (N_3300,N_290,N_1456);
or U3301 (N_3301,N_2227,N_355);
and U3302 (N_3302,N_2161,N_68);
nor U3303 (N_3303,N_72,N_2083);
xor U3304 (N_3304,N_1245,N_1674);
and U3305 (N_3305,N_2186,N_437);
nand U3306 (N_3306,N_1180,N_139);
nand U3307 (N_3307,N_178,N_691);
or U3308 (N_3308,N_1465,N_834);
nor U3309 (N_3309,N_2133,N_1714);
and U3310 (N_3310,N_2332,N_2111);
and U3311 (N_3311,N_1381,N_25);
nor U3312 (N_3312,N_1667,N_1161);
xnor U3313 (N_3313,N_817,N_601);
or U3314 (N_3314,N_2343,N_1595);
xnor U3315 (N_3315,N_1228,N_674);
or U3316 (N_3316,N_2478,N_913);
nor U3317 (N_3317,N_1365,N_1625);
nand U3318 (N_3318,N_2436,N_153);
nand U3319 (N_3319,N_268,N_2058);
and U3320 (N_3320,N_1310,N_2198);
xor U3321 (N_3321,N_1109,N_201);
and U3322 (N_3322,N_940,N_2283);
nor U3323 (N_3323,N_670,N_1220);
nor U3324 (N_3324,N_916,N_859);
nand U3325 (N_3325,N_2102,N_2263);
or U3326 (N_3326,N_161,N_1009);
nor U3327 (N_3327,N_1256,N_2184);
nor U3328 (N_3328,N_2091,N_1242);
and U3329 (N_3329,N_1402,N_912);
nand U3330 (N_3330,N_2149,N_2070);
nor U3331 (N_3331,N_1199,N_1192);
and U3332 (N_3332,N_326,N_1960);
nor U3333 (N_3333,N_2039,N_1297);
and U3334 (N_3334,N_114,N_636);
and U3335 (N_3335,N_442,N_789);
nand U3336 (N_3336,N_2313,N_1502);
and U3337 (N_3337,N_725,N_450);
xnor U3338 (N_3338,N_287,N_617);
xnor U3339 (N_3339,N_104,N_717);
nor U3340 (N_3340,N_342,N_2495);
and U3341 (N_3341,N_1826,N_2157);
and U3342 (N_3342,N_1176,N_584);
nor U3343 (N_3343,N_318,N_1880);
or U3344 (N_3344,N_285,N_718);
nor U3345 (N_3345,N_1867,N_2231);
and U3346 (N_3346,N_1160,N_9);
nand U3347 (N_3347,N_1633,N_362);
and U3348 (N_3348,N_2369,N_280);
and U3349 (N_3349,N_1763,N_1089);
nand U3350 (N_3350,N_291,N_857);
or U3351 (N_3351,N_1620,N_1208);
nand U3352 (N_3352,N_756,N_141);
nor U3353 (N_3353,N_1290,N_337);
xor U3354 (N_3354,N_2103,N_256);
or U3355 (N_3355,N_769,N_2196);
xnor U3356 (N_3356,N_2023,N_1409);
nor U3357 (N_3357,N_33,N_2395);
nand U3358 (N_3358,N_1454,N_1697);
xor U3359 (N_3359,N_1052,N_1123);
or U3360 (N_3360,N_884,N_70);
nor U3361 (N_3361,N_922,N_1023);
xor U3362 (N_3362,N_578,N_2403);
or U3363 (N_3363,N_612,N_741);
nand U3364 (N_3364,N_384,N_2095);
nand U3365 (N_3365,N_48,N_59);
nor U3366 (N_3366,N_689,N_1171);
and U3367 (N_3367,N_2172,N_117);
nand U3368 (N_3368,N_867,N_1508);
nand U3369 (N_3369,N_2248,N_2048);
nand U3370 (N_3370,N_1200,N_997);
xor U3371 (N_3371,N_929,N_440);
or U3372 (N_3372,N_1609,N_420);
and U3373 (N_3373,N_413,N_649);
or U3374 (N_3374,N_1082,N_2214);
or U3375 (N_3375,N_1513,N_528);
and U3376 (N_3376,N_1311,N_1422);
nor U3377 (N_3377,N_1331,N_2);
nor U3378 (N_3378,N_1532,N_433);
nor U3379 (N_3379,N_1090,N_975);
or U3380 (N_3380,N_1383,N_696);
and U3381 (N_3381,N_770,N_2361);
xnor U3382 (N_3382,N_2125,N_2216);
and U3383 (N_3383,N_1624,N_1660);
and U3384 (N_3384,N_970,N_1942);
nand U3385 (N_3385,N_2078,N_1327);
nor U3386 (N_3386,N_2322,N_411);
nor U3387 (N_3387,N_609,N_933);
nor U3388 (N_3388,N_377,N_2104);
or U3389 (N_3389,N_204,N_277);
nand U3390 (N_3390,N_1887,N_1062);
or U3391 (N_3391,N_2466,N_2188);
nor U3392 (N_3392,N_1350,N_1576);
and U3393 (N_3393,N_1084,N_2319);
nor U3394 (N_3394,N_1352,N_2311);
or U3395 (N_3395,N_2230,N_1899);
nor U3396 (N_3396,N_1272,N_77);
nor U3397 (N_3397,N_994,N_599);
nand U3398 (N_3398,N_1986,N_325);
and U3399 (N_3399,N_753,N_711);
or U3400 (N_3400,N_2456,N_963);
nor U3401 (N_3401,N_241,N_2142);
nand U3402 (N_3402,N_262,N_2132);
and U3403 (N_3403,N_1718,N_89);
nor U3404 (N_3404,N_1473,N_1377);
nor U3405 (N_3405,N_1810,N_2215);
nor U3406 (N_3406,N_79,N_619);
nand U3407 (N_3407,N_896,N_1954);
or U3408 (N_3408,N_1614,N_40);
and U3409 (N_3409,N_1432,N_2176);
and U3410 (N_3410,N_567,N_107);
and U3411 (N_3411,N_210,N_1278);
xnor U3412 (N_3412,N_1961,N_2485);
nor U3413 (N_3413,N_2417,N_856);
nor U3414 (N_3414,N_972,N_1976);
nand U3415 (N_3415,N_2124,N_682);
and U3416 (N_3416,N_468,N_69);
xnor U3417 (N_3417,N_2138,N_2178);
and U3418 (N_3418,N_1499,N_2165);
nor U3419 (N_3419,N_1687,N_1019);
or U3420 (N_3420,N_797,N_2027);
and U3421 (N_3421,N_1675,N_115);
and U3422 (N_3422,N_1866,N_397);
and U3423 (N_3423,N_2068,N_1184);
and U3424 (N_3424,N_477,N_1179);
nand U3425 (N_3425,N_1941,N_840);
or U3426 (N_3426,N_706,N_532);
and U3427 (N_3427,N_1732,N_1028);
nor U3428 (N_3428,N_1699,N_1405);
and U3429 (N_3429,N_1794,N_1168);
nand U3430 (N_3430,N_2305,N_1157);
xor U3431 (N_3431,N_2467,N_585);
and U3432 (N_3432,N_553,N_1725);
or U3433 (N_3433,N_338,N_1592);
nor U3434 (N_3434,N_1585,N_260);
nand U3435 (N_3435,N_2013,N_1063);
nand U3436 (N_3436,N_734,N_1771);
nor U3437 (N_3437,N_2391,N_348);
or U3438 (N_3438,N_456,N_1524);
and U3439 (N_3439,N_1705,N_1216);
or U3440 (N_3440,N_1964,N_501);
or U3441 (N_3441,N_2373,N_1444);
xnor U3442 (N_3442,N_1188,N_1739);
and U3443 (N_3443,N_1602,N_333);
nand U3444 (N_3444,N_390,N_1996);
and U3445 (N_3445,N_1210,N_2226);
xnor U3446 (N_3446,N_1044,N_1967);
xnor U3447 (N_3447,N_2112,N_1704);
nor U3448 (N_3448,N_505,N_738);
and U3449 (N_3449,N_1711,N_176);
or U3450 (N_3450,N_1833,N_1531);
and U3451 (N_3451,N_180,N_968);
nand U3452 (N_3452,N_579,N_2486);
and U3453 (N_3453,N_659,N_1578);
and U3454 (N_3454,N_2271,N_981);
xnor U3455 (N_3455,N_2204,N_441);
and U3456 (N_3456,N_1498,N_1603);
or U3457 (N_3457,N_730,N_1166);
nand U3458 (N_3458,N_1112,N_2472);
nand U3459 (N_3459,N_120,N_1313);
xnor U3460 (N_3460,N_2452,N_1255);
nor U3461 (N_3461,N_1204,N_846);
and U3462 (N_3462,N_2051,N_251);
xnor U3463 (N_3463,N_202,N_8);
nand U3464 (N_3464,N_504,N_597);
and U3465 (N_3465,N_1430,N_1067);
nor U3466 (N_3466,N_1385,N_513);
or U3467 (N_3467,N_604,N_1404);
nand U3468 (N_3468,N_777,N_489);
and U3469 (N_3469,N_710,N_169);
or U3470 (N_3470,N_1584,N_2160);
nand U3471 (N_3471,N_373,N_236);
and U3472 (N_3472,N_2407,N_2060);
nand U3473 (N_3473,N_1328,N_845);
xnor U3474 (N_3474,N_825,N_2371);
nor U3475 (N_3475,N_1496,N_1862);
xor U3476 (N_3476,N_1235,N_106);
xor U3477 (N_3477,N_1815,N_1027);
or U3478 (N_3478,N_1884,N_317);
nor U3479 (N_3479,N_808,N_1494);
and U3480 (N_3480,N_2427,N_1186);
nand U3481 (N_3481,N_512,N_1533);
nand U3482 (N_3482,N_1049,N_1279);
nor U3483 (N_3483,N_1804,N_2375);
nor U3484 (N_3484,N_1445,N_108);
nand U3485 (N_3485,N_1182,N_1876);
and U3486 (N_3486,N_2177,N_1197);
nor U3487 (N_3487,N_97,N_1688);
nor U3488 (N_3488,N_435,N_2304);
nand U3489 (N_3489,N_138,N_750);
and U3490 (N_3490,N_2007,N_551);
and U3491 (N_3491,N_886,N_563);
or U3492 (N_3492,N_1223,N_221);
and U3493 (N_3493,N_1072,N_1111);
nor U3494 (N_3494,N_2018,N_1181);
and U3495 (N_3495,N_75,N_1474);
nor U3496 (N_3496,N_1213,N_140);
and U3497 (N_3497,N_1408,N_1293);
and U3498 (N_3498,N_2300,N_1698);
nand U3499 (N_3499,N_295,N_2451);
nand U3500 (N_3500,N_387,N_2242);
and U3501 (N_3501,N_1227,N_1277);
nand U3502 (N_3502,N_428,N_2482);
or U3503 (N_3503,N_137,N_1832);
nand U3504 (N_3504,N_714,N_2118);
nor U3505 (N_3505,N_1793,N_43);
xor U3506 (N_3506,N_322,N_1813);
and U3507 (N_3507,N_1321,N_2052);
xor U3508 (N_3508,N_2488,N_544);
and U3509 (N_3509,N_1092,N_2265);
and U3510 (N_3510,N_1191,N_646);
nand U3511 (N_3511,N_497,N_2109);
and U3512 (N_3512,N_1641,N_1756);
nand U3513 (N_3513,N_1372,N_481);
and U3514 (N_3514,N_1320,N_1392);
nor U3515 (N_3515,N_499,N_2470);
and U3516 (N_3516,N_1150,N_1567);
or U3517 (N_3517,N_353,N_252);
and U3518 (N_3518,N_1596,N_821);
nand U3519 (N_3519,N_425,N_1859);
nor U3520 (N_3520,N_51,N_1263);
nand U3521 (N_3521,N_1307,N_1116);
xnor U3522 (N_3522,N_531,N_1509);
nor U3523 (N_3523,N_764,N_1292);
nor U3524 (N_3524,N_818,N_1476);
or U3525 (N_3525,N_26,N_1747);
nor U3526 (N_3526,N_971,N_12);
and U3527 (N_3527,N_776,N_1032);
nand U3528 (N_3528,N_2435,N_225);
nand U3529 (N_3529,N_90,N_1105);
nand U3530 (N_3530,N_890,N_336);
nor U3531 (N_3531,N_132,N_1924);
nand U3532 (N_3532,N_167,N_179);
or U3533 (N_3533,N_824,N_716);
nand U3534 (N_3534,N_1165,N_458);
or U3535 (N_3535,N_506,N_1775);
nor U3536 (N_3536,N_2372,N_1795);
nand U3537 (N_3537,N_1760,N_2387);
nand U3538 (N_3538,N_1684,N_2073);
and U3539 (N_3539,N_1395,N_1978);
nand U3540 (N_3540,N_1984,N_1721);
nor U3541 (N_3541,N_2489,N_2328);
nand U3542 (N_3542,N_2174,N_1510);
or U3543 (N_3543,N_2129,N_1708);
and U3544 (N_3544,N_400,N_2075);
nor U3545 (N_3545,N_307,N_374);
or U3546 (N_3546,N_1663,N_1605);
and U3547 (N_3547,N_2232,N_1786);
nand U3548 (N_3548,N_2105,N_129);
nor U3549 (N_3549,N_1364,N_452);
or U3550 (N_3550,N_243,N_310);
nand U3551 (N_3551,N_1568,N_850);
nor U3552 (N_3552,N_1207,N_1574);
and U3553 (N_3553,N_2406,N_1825);
nor U3554 (N_3554,N_2445,N_1436);
nand U3555 (N_3555,N_1238,N_785);
nor U3556 (N_3556,N_2006,N_238);
or U3557 (N_3557,N_101,N_999);
or U3558 (N_3558,N_740,N_576);
or U3559 (N_3559,N_583,N_1345);
or U3560 (N_3560,N_2147,N_1657);
or U3561 (N_3561,N_2222,N_394);
or U3562 (N_3562,N_2117,N_1217);
nand U3563 (N_3563,N_1342,N_2397);
or U3564 (N_3564,N_224,N_2029);
nand U3565 (N_3565,N_0,N_1492);
xor U3566 (N_3566,N_2213,N_2274);
xnor U3567 (N_3567,N_666,N_2146);
nand U3568 (N_3568,N_1901,N_2239);
and U3569 (N_3569,N_2394,N_81);
or U3570 (N_3570,N_281,N_1457);
nor U3571 (N_3571,N_2236,N_1902);
nand U3572 (N_3572,N_907,N_937);
nor U3573 (N_3573,N_1971,N_1563);
nor U3574 (N_3574,N_957,N_569);
nor U3575 (N_3575,N_1398,N_1865);
nand U3576 (N_3576,N_2286,N_976);
nand U3577 (N_3577,N_518,N_592);
and U3578 (N_3578,N_1281,N_524);
nor U3579 (N_3579,N_1488,N_2179);
or U3580 (N_3580,N_1676,N_1282);
or U3581 (N_3581,N_874,N_833);
nand U3582 (N_3582,N_2121,N_245);
or U3583 (N_3583,N_1598,N_1500);
nor U3584 (N_3584,N_888,N_2378);
xnor U3585 (N_3585,N_2382,N_91);
nand U3586 (N_3586,N_2025,N_1087);
nand U3587 (N_3587,N_1664,N_233);
nand U3588 (N_3588,N_2183,N_265);
xor U3589 (N_3589,N_2249,N_2446);
nor U3590 (N_3590,N_2287,N_467);
and U3591 (N_3591,N_1371,N_1746);
nor U3592 (N_3592,N_2444,N_2440);
nand U3593 (N_3593,N_449,N_383);
xnor U3594 (N_3594,N_582,N_1905);
nor U3595 (N_3595,N_608,N_464);
nor U3596 (N_3596,N_55,N_304);
or U3597 (N_3597,N_1842,N_62);
nor U3598 (N_3598,N_688,N_99);
and U3599 (N_3599,N_1953,N_2462);
or U3600 (N_3600,N_94,N_1566);
nor U3601 (N_3601,N_2457,N_1387);
nor U3602 (N_3602,N_1301,N_2402);
xnor U3603 (N_3603,N_434,N_1020);
nand U3604 (N_3604,N_1873,N_19);
nand U3605 (N_3605,N_2262,N_1943);
and U3606 (N_3606,N_2144,N_308);
or U3607 (N_3607,N_1888,N_1241);
and U3608 (N_3608,N_803,N_1846);
nor U3609 (N_3609,N_1338,N_774);
xor U3610 (N_3610,N_1575,N_733);
nor U3611 (N_3611,N_535,N_1716);
xnor U3612 (N_3612,N_194,N_1471);
and U3613 (N_3613,N_1818,N_1051);
nor U3614 (N_3614,N_1761,N_249);
xor U3615 (N_3615,N_1442,N_702);
or U3616 (N_3616,N_1196,N_1767);
and U3617 (N_3617,N_722,N_1511);
and U3618 (N_3618,N_1845,N_417);
or U3619 (N_3619,N_2342,N_85);
and U3620 (N_3620,N_208,N_559);
or U3621 (N_3621,N_1556,N_1098);
nand U3622 (N_3622,N_2096,N_2302);
and U3623 (N_3623,N_620,N_2042);
nor U3624 (N_3624,N_244,N_1162);
nor U3625 (N_3625,N_561,N_2335);
or U3626 (N_3626,N_671,N_1743);
or U3627 (N_3627,N_613,N_2376);
or U3628 (N_3628,N_1712,N_1252);
or U3629 (N_3629,N_1562,N_100);
nor U3630 (N_3630,N_1011,N_1963);
nand U3631 (N_3631,N_679,N_1344);
or U3632 (N_3632,N_2307,N_58);
and U3633 (N_3633,N_2041,N_934);
nor U3634 (N_3634,N_598,N_2088);
and U3635 (N_3635,N_496,N_1170);
and U3636 (N_3636,N_650,N_67);
nor U3637 (N_3637,N_1821,N_622);
or U3638 (N_3638,N_2217,N_2201);
or U3639 (N_3639,N_667,N_974);
nand U3640 (N_3640,N_2409,N_125);
or U3641 (N_3641,N_1979,N_1487);
and U3642 (N_3642,N_2143,N_683);
nor U3643 (N_3643,N_969,N_278);
or U3644 (N_3644,N_2087,N_1410);
or U3645 (N_3645,N_220,N_681);
or U3646 (N_3646,N_329,N_1355);
and U3647 (N_3647,N_231,N_588);
nand U3648 (N_3648,N_354,N_1079);
xor U3649 (N_3649,N_1376,N_1998);
nand U3650 (N_3650,N_1018,N_2069);
xor U3651 (N_3651,N_973,N_73);
nand U3652 (N_3652,N_2152,N_1209);
nand U3653 (N_3653,N_2067,N_526);
nor U3654 (N_3654,N_810,N_855);
or U3655 (N_3655,N_263,N_1115);
or U3656 (N_3656,N_18,N_1920);
nand U3657 (N_3657,N_1940,N_2127);
nand U3658 (N_3658,N_1336,N_1734);
and U3659 (N_3659,N_1977,N_1632);
nand U3660 (N_3660,N_1898,N_1485);
and U3661 (N_3661,N_677,N_1056);
nor U3662 (N_3662,N_2247,N_1038);
and U3663 (N_3663,N_1800,N_2356);
nand U3664 (N_3664,N_639,N_2293);
nor U3665 (N_3665,N_1886,N_1987);
or U3666 (N_3666,N_443,N_1913);
or U3667 (N_3667,N_315,N_2327);
nor U3668 (N_3668,N_1548,N_951);
nand U3669 (N_3669,N_2383,N_590);
and U3670 (N_3670,N_1534,N_728);
or U3671 (N_3671,N_1581,N_1593);
and U3672 (N_3672,N_2374,N_796);
nor U3673 (N_3673,N_2385,N_1909);
nor U3674 (N_3674,N_842,N_2072);
or U3675 (N_3675,N_2046,N_1600);
nand U3676 (N_3676,N_279,N_1094);
nand U3677 (N_3677,N_1545,N_1356);
nor U3678 (N_3678,N_2421,N_2359);
nand U3679 (N_3679,N_1249,N_986);
xor U3680 (N_3680,N_804,N_364);
nor U3681 (N_3681,N_2494,N_2243);
and U3682 (N_3682,N_1916,N_2481);
and U3683 (N_3683,N_2028,N_283);
or U3684 (N_3684,N_199,N_1419);
and U3685 (N_3685,N_1138,N_765);
or U3686 (N_3686,N_2030,N_2115);
and U3687 (N_3687,N_832,N_1440);
xor U3688 (N_3688,N_1900,N_847);
or U3689 (N_3689,N_1949,N_1983);
or U3690 (N_3690,N_1464,N_2292);
and U3691 (N_3691,N_398,N_2330);
xor U3692 (N_3692,N_396,N_1525);
nor U3693 (N_3693,N_2377,N_2008);
or U3694 (N_3694,N_1033,N_235);
nor U3695 (N_3695,N_1426,N_2043);
xor U3696 (N_3696,N_950,N_1195);
nor U3697 (N_3697,N_2194,N_1239);
nor U3698 (N_3698,N_1610,N_2473);
nand U3699 (N_3699,N_2037,N_150);
nor U3700 (N_3700,N_2202,N_2388);
and U3701 (N_3701,N_1988,N_2208);
nand U3702 (N_3702,N_469,N_1024);
or U3703 (N_3703,N_379,N_1268);
or U3704 (N_3704,N_1911,N_1802);
xor U3705 (N_3705,N_335,N_1144);
nor U3706 (N_3706,N_2460,N_2033);
or U3707 (N_3707,N_2252,N_1779);
nor U3708 (N_3708,N_127,N_1519);
nor U3709 (N_3709,N_1594,N_1394);
nor U3710 (N_3710,N_1764,N_600);
nor U3711 (N_3711,N_2045,N_2464);
and U3712 (N_3712,N_2419,N_1147);
nor U3713 (N_3713,N_1579,N_2282);
or U3714 (N_3714,N_2181,N_123);
and U3715 (N_3715,N_324,N_453);
nand U3716 (N_3716,N_1552,N_1267);
xor U3717 (N_3717,N_1326,N_228);
and U3718 (N_3718,N_196,N_1124);
nor U3719 (N_3719,N_490,N_841);
nand U3720 (N_3720,N_899,N_1253);
nor U3721 (N_3721,N_195,N_1638);
or U3722 (N_3722,N_2234,N_1738);
and U3723 (N_3723,N_2139,N_1076);
xnor U3724 (N_3724,N_1309,N_648);
or U3725 (N_3725,N_739,N_593);
nor U3726 (N_3726,N_421,N_2065);
or U3727 (N_3727,N_1626,N_250);
and U3728 (N_3728,N_49,N_673);
and U3729 (N_3729,N_1852,N_2288);
or U3730 (N_3730,N_891,N_190);
nand U3731 (N_3731,N_2318,N_2107);
nor U3732 (N_3732,N_1362,N_1169);
and U3733 (N_3733,N_815,N_1030);
and U3734 (N_3734,N_1661,N_30);
nor U3735 (N_3735,N_1538,N_2126);
nand U3736 (N_3736,N_2281,N_16);
or U3737 (N_3737,N_1787,N_7);
nor U3738 (N_3738,N_444,N_2268);
nor U3739 (N_3739,N_1299,N_701);
and U3740 (N_3740,N_1975,N_2386);
and U3741 (N_3741,N_2054,N_866);
nand U3742 (N_3742,N_1428,N_294);
nor U3743 (N_3743,N_1669,N_2303);
nand U3744 (N_3744,N_1081,N_1149);
and U3745 (N_3745,N_1271,N_2015);
nand U3746 (N_3746,N_791,N_555);
xnor U3747 (N_3747,N_2334,N_35);
nor U3748 (N_3748,N_1261,N_2245);
and U3749 (N_3749,N_2099,N_1155);
and U3750 (N_3750,N_603,N_1294);
and U3751 (N_3751,N_401,N_52);
nor U3752 (N_3752,N_2251,N_1784);
or U3753 (N_3753,N_2362,N_135);
xor U3754 (N_3754,N_1136,N_2393);
and U3755 (N_3755,N_2031,N_1109);
and U3756 (N_3756,N_1958,N_1927);
nor U3757 (N_3757,N_406,N_2232);
nor U3758 (N_3758,N_1510,N_1961);
and U3759 (N_3759,N_695,N_2461);
or U3760 (N_3760,N_739,N_1789);
nand U3761 (N_3761,N_213,N_2198);
and U3762 (N_3762,N_2385,N_978);
nand U3763 (N_3763,N_748,N_389);
and U3764 (N_3764,N_35,N_1821);
and U3765 (N_3765,N_720,N_1727);
nand U3766 (N_3766,N_1171,N_2283);
nand U3767 (N_3767,N_2138,N_407);
nand U3768 (N_3768,N_1145,N_517);
nor U3769 (N_3769,N_924,N_1923);
or U3770 (N_3770,N_584,N_142);
xor U3771 (N_3771,N_889,N_1289);
nor U3772 (N_3772,N_605,N_224);
nand U3773 (N_3773,N_60,N_2178);
or U3774 (N_3774,N_1856,N_1083);
and U3775 (N_3775,N_637,N_1892);
or U3776 (N_3776,N_1369,N_1770);
nand U3777 (N_3777,N_849,N_1593);
nor U3778 (N_3778,N_152,N_2151);
nand U3779 (N_3779,N_1552,N_2204);
nor U3780 (N_3780,N_2438,N_1582);
nor U3781 (N_3781,N_17,N_1800);
or U3782 (N_3782,N_2296,N_910);
or U3783 (N_3783,N_1758,N_554);
or U3784 (N_3784,N_2415,N_1667);
xnor U3785 (N_3785,N_33,N_1174);
nor U3786 (N_3786,N_71,N_334);
nor U3787 (N_3787,N_2303,N_1322);
nor U3788 (N_3788,N_1321,N_675);
and U3789 (N_3789,N_618,N_97);
and U3790 (N_3790,N_114,N_572);
nor U3791 (N_3791,N_1572,N_431);
and U3792 (N_3792,N_648,N_706);
nand U3793 (N_3793,N_1172,N_2339);
nand U3794 (N_3794,N_2129,N_570);
nand U3795 (N_3795,N_229,N_2426);
xnor U3796 (N_3796,N_226,N_172);
xnor U3797 (N_3797,N_694,N_1203);
and U3798 (N_3798,N_81,N_2177);
nor U3799 (N_3799,N_1184,N_1201);
nand U3800 (N_3800,N_2075,N_183);
xnor U3801 (N_3801,N_2154,N_646);
or U3802 (N_3802,N_2156,N_2096);
xnor U3803 (N_3803,N_607,N_1982);
and U3804 (N_3804,N_658,N_599);
or U3805 (N_3805,N_2176,N_2197);
nand U3806 (N_3806,N_707,N_1433);
and U3807 (N_3807,N_802,N_809);
or U3808 (N_3808,N_1679,N_1886);
and U3809 (N_3809,N_1982,N_724);
or U3810 (N_3810,N_2104,N_1109);
and U3811 (N_3811,N_1174,N_1327);
and U3812 (N_3812,N_869,N_360);
or U3813 (N_3813,N_351,N_2462);
nand U3814 (N_3814,N_1591,N_38);
or U3815 (N_3815,N_1763,N_852);
and U3816 (N_3816,N_989,N_1148);
and U3817 (N_3817,N_1954,N_155);
nor U3818 (N_3818,N_1185,N_573);
nor U3819 (N_3819,N_1039,N_2404);
nor U3820 (N_3820,N_141,N_47);
and U3821 (N_3821,N_91,N_23);
nand U3822 (N_3822,N_51,N_1935);
and U3823 (N_3823,N_2226,N_1708);
nand U3824 (N_3824,N_2356,N_1318);
and U3825 (N_3825,N_2250,N_1980);
and U3826 (N_3826,N_1554,N_673);
xnor U3827 (N_3827,N_2253,N_434);
and U3828 (N_3828,N_473,N_1280);
and U3829 (N_3829,N_2074,N_883);
nand U3830 (N_3830,N_1370,N_803);
nor U3831 (N_3831,N_943,N_1918);
or U3832 (N_3832,N_1997,N_671);
nand U3833 (N_3833,N_2204,N_2207);
or U3834 (N_3834,N_478,N_1791);
and U3835 (N_3835,N_2430,N_247);
nand U3836 (N_3836,N_1019,N_574);
or U3837 (N_3837,N_1343,N_1185);
nor U3838 (N_3838,N_931,N_75);
and U3839 (N_3839,N_1859,N_549);
xor U3840 (N_3840,N_670,N_419);
nor U3841 (N_3841,N_1084,N_732);
or U3842 (N_3842,N_191,N_682);
nor U3843 (N_3843,N_342,N_1312);
and U3844 (N_3844,N_2062,N_164);
xor U3845 (N_3845,N_127,N_865);
nor U3846 (N_3846,N_2030,N_1919);
nor U3847 (N_3847,N_139,N_2218);
nand U3848 (N_3848,N_1609,N_977);
nand U3849 (N_3849,N_276,N_1008);
xor U3850 (N_3850,N_147,N_63);
nand U3851 (N_3851,N_33,N_2177);
or U3852 (N_3852,N_1266,N_1681);
or U3853 (N_3853,N_2030,N_1967);
xnor U3854 (N_3854,N_2334,N_848);
xor U3855 (N_3855,N_1177,N_1333);
nand U3856 (N_3856,N_492,N_118);
nand U3857 (N_3857,N_2025,N_1689);
nor U3858 (N_3858,N_2116,N_1095);
nor U3859 (N_3859,N_489,N_1641);
and U3860 (N_3860,N_1464,N_1012);
nor U3861 (N_3861,N_1466,N_1804);
nand U3862 (N_3862,N_1026,N_598);
nor U3863 (N_3863,N_1123,N_1464);
and U3864 (N_3864,N_2084,N_1532);
nand U3865 (N_3865,N_2469,N_1522);
nor U3866 (N_3866,N_1797,N_1914);
nand U3867 (N_3867,N_1060,N_2163);
and U3868 (N_3868,N_932,N_2440);
and U3869 (N_3869,N_1043,N_73);
nor U3870 (N_3870,N_1891,N_757);
nand U3871 (N_3871,N_897,N_2473);
nor U3872 (N_3872,N_1449,N_1761);
nand U3873 (N_3873,N_2151,N_317);
nand U3874 (N_3874,N_1330,N_2497);
or U3875 (N_3875,N_2025,N_2136);
nand U3876 (N_3876,N_2008,N_2068);
nor U3877 (N_3877,N_1586,N_1134);
xor U3878 (N_3878,N_2136,N_858);
nor U3879 (N_3879,N_616,N_1807);
nor U3880 (N_3880,N_1536,N_1823);
and U3881 (N_3881,N_768,N_1721);
nor U3882 (N_3882,N_661,N_1955);
nand U3883 (N_3883,N_1013,N_816);
nand U3884 (N_3884,N_2494,N_1848);
xor U3885 (N_3885,N_1506,N_183);
nor U3886 (N_3886,N_732,N_1235);
xor U3887 (N_3887,N_1182,N_1470);
and U3888 (N_3888,N_1753,N_1844);
or U3889 (N_3889,N_263,N_633);
nand U3890 (N_3890,N_124,N_1786);
nor U3891 (N_3891,N_2438,N_1504);
nand U3892 (N_3892,N_1103,N_2424);
nand U3893 (N_3893,N_2410,N_1199);
nor U3894 (N_3894,N_200,N_1451);
and U3895 (N_3895,N_1983,N_1334);
or U3896 (N_3896,N_58,N_867);
nand U3897 (N_3897,N_1089,N_705);
nand U3898 (N_3898,N_654,N_381);
xor U3899 (N_3899,N_2107,N_1122);
and U3900 (N_3900,N_1938,N_110);
and U3901 (N_3901,N_621,N_742);
nand U3902 (N_3902,N_604,N_440);
nand U3903 (N_3903,N_2314,N_2356);
or U3904 (N_3904,N_747,N_1684);
nand U3905 (N_3905,N_747,N_1790);
nand U3906 (N_3906,N_421,N_1303);
or U3907 (N_3907,N_330,N_2427);
and U3908 (N_3908,N_226,N_1710);
nor U3909 (N_3909,N_405,N_309);
or U3910 (N_3910,N_244,N_1353);
or U3911 (N_3911,N_1221,N_1628);
and U3912 (N_3912,N_1104,N_1006);
or U3913 (N_3913,N_279,N_707);
or U3914 (N_3914,N_1777,N_2115);
nand U3915 (N_3915,N_202,N_1603);
and U3916 (N_3916,N_1626,N_976);
or U3917 (N_3917,N_1634,N_264);
nor U3918 (N_3918,N_1425,N_414);
nand U3919 (N_3919,N_492,N_249);
nor U3920 (N_3920,N_1131,N_1214);
and U3921 (N_3921,N_191,N_2385);
and U3922 (N_3922,N_1318,N_405);
and U3923 (N_3923,N_1471,N_708);
nand U3924 (N_3924,N_1093,N_2466);
nand U3925 (N_3925,N_892,N_1133);
nor U3926 (N_3926,N_2311,N_411);
and U3927 (N_3927,N_1090,N_1571);
nand U3928 (N_3928,N_2486,N_1572);
or U3929 (N_3929,N_2349,N_356);
nor U3930 (N_3930,N_399,N_1479);
nand U3931 (N_3931,N_312,N_559);
xnor U3932 (N_3932,N_1409,N_1941);
nor U3933 (N_3933,N_1861,N_713);
nand U3934 (N_3934,N_1042,N_302);
xnor U3935 (N_3935,N_881,N_1867);
and U3936 (N_3936,N_1184,N_282);
nor U3937 (N_3937,N_1130,N_1961);
xnor U3938 (N_3938,N_1392,N_644);
and U3939 (N_3939,N_637,N_1629);
or U3940 (N_3940,N_328,N_702);
xor U3941 (N_3941,N_1192,N_1507);
nand U3942 (N_3942,N_466,N_1568);
and U3943 (N_3943,N_1302,N_180);
and U3944 (N_3944,N_321,N_946);
or U3945 (N_3945,N_2025,N_1376);
or U3946 (N_3946,N_2310,N_2149);
nand U3947 (N_3947,N_2341,N_2288);
nand U3948 (N_3948,N_628,N_670);
nand U3949 (N_3949,N_234,N_1545);
nor U3950 (N_3950,N_303,N_740);
xor U3951 (N_3951,N_228,N_561);
or U3952 (N_3952,N_527,N_980);
nor U3953 (N_3953,N_2375,N_1767);
or U3954 (N_3954,N_489,N_1820);
nand U3955 (N_3955,N_2340,N_2052);
or U3956 (N_3956,N_345,N_455);
xnor U3957 (N_3957,N_48,N_1254);
or U3958 (N_3958,N_1007,N_89);
and U3959 (N_3959,N_156,N_329);
nand U3960 (N_3960,N_1103,N_583);
nor U3961 (N_3961,N_81,N_1307);
nor U3962 (N_3962,N_1830,N_2199);
and U3963 (N_3963,N_215,N_2435);
or U3964 (N_3964,N_1233,N_434);
or U3965 (N_3965,N_835,N_11);
nor U3966 (N_3966,N_1921,N_897);
nor U3967 (N_3967,N_2236,N_318);
and U3968 (N_3968,N_2231,N_1296);
nor U3969 (N_3969,N_610,N_1544);
xor U3970 (N_3970,N_2191,N_1348);
nor U3971 (N_3971,N_77,N_839);
or U3972 (N_3972,N_1188,N_2112);
and U3973 (N_3973,N_1636,N_934);
xor U3974 (N_3974,N_2198,N_936);
nand U3975 (N_3975,N_1797,N_2493);
nand U3976 (N_3976,N_104,N_2291);
or U3977 (N_3977,N_2039,N_461);
nor U3978 (N_3978,N_1010,N_214);
or U3979 (N_3979,N_2307,N_1156);
or U3980 (N_3980,N_1159,N_1594);
and U3981 (N_3981,N_745,N_2395);
nand U3982 (N_3982,N_268,N_2457);
nand U3983 (N_3983,N_1316,N_1264);
and U3984 (N_3984,N_1468,N_1051);
and U3985 (N_3985,N_2342,N_671);
and U3986 (N_3986,N_1241,N_1642);
and U3987 (N_3987,N_2138,N_1631);
nor U3988 (N_3988,N_2276,N_1413);
and U3989 (N_3989,N_802,N_1754);
nand U3990 (N_3990,N_222,N_1814);
nor U3991 (N_3991,N_1813,N_855);
or U3992 (N_3992,N_693,N_331);
or U3993 (N_3993,N_2222,N_939);
nand U3994 (N_3994,N_2339,N_453);
nand U3995 (N_3995,N_1684,N_166);
or U3996 (N_3996,N_410,N_530);
or U3997 (N_3997,N_26,N_776);
nor U3998 (N_3998,N_2386,N_918);
xnor U3999 (N_3999,N_1864,N_2404);
nand U4000 (N_4000,N_1871,N_449);
and U4001 (N_4001,N_749,N_1615);
nor U4002 (N_4002,N_497,N_568);
or U4003 (N_4003,N_2025,N_970);
or U4004 (N_4004,N_1245,N_193);
nand U4005 (N_4005,N_1540,N_1401);
and U4006 (N_4006,N_1418,N_1730);
nand U4007 (N_4007,N_1443,N_1880);
xor U4008 (N_4008,N_575,N_171);
and U4009 (N_4009,N_722,N_1017);
nand U4010 (N_4010,N_391,N_1833);
nand U4011 (N_4011,N_74,N_753);
xor U4012 (N_4012,N_1917,N_1807);
nand U4013 (N_4013,N_2064,N_957);
or U4014 (N_4014,N_2108,N_1307);
nor U4015 (N_4015,N_2451,N_921);
or U4016 (N_4016,N_1730,N_1575);
or U4017 (N_4017,N_237,N_1408);
nor U4018 (N_4018,N_2267,N_1606);
or U4019 (N_4019,N_1556,N_1198);
nor U4020 (N_4020,N_2421,N_1339);
xor U4021 (N_4021,N_521,N_2330);
and U4022 (N_4022,N_282,N_324);
and U4023 (N_4023,N_2439,N_181);
xor U4024 (N_4024,N_1763,N_2303);
nor U4025 (N_4025,N_173,N_2055);
nor U4026 (N_4026,N_2240,N_1194);
or U4027 (N_4027,N_1834,N_2473);
nor U4028 (N_4028,N_1036,N_1885);
or U4029 (N_4029,N_129,N_1034);
nor U4030 (N_4030,N_19,N_476);
nand U4031 (N_4031,N_627,N_649);
and U4032 (N_4032,N_544,N_955);
nand U4033 (N_4033,N_2485,N_1964);
nor U4034 (N_4034,N_1974,N_1031);
nand U4035 (N_4035,N_1845,N_1639);
nand U4036 (N_4036,N_443,N_1668);
nand U4037 (N_4037,N_8,N_22);
or U4038 (N_4038,N_475,N_2031);
and U4039 (N_4039,N_2330,N_1312);
nand U4040 (N_4040,N_408,N_1301);
nor U4041 (N_4041,N_898,N_291);
nor U4042 (N_4042,N_488,N_2362);
nor U4043 (N_4043,N_930,N_633);
nand U4044 (N_4044,N_2310,N_859);
and U4045 (N_4045,N_805,N_1315);
and U4046 (N_4046,N_706,N_719);
nand U4047 (N_4047,N_728,N_1375);
and U4048 (N_4048,N_613,N_1474);
nand U4049 (N_4049,N_291,N_976);
nor U4050 (N_4050,N_1996,N_1794);
and U4051 (N_4051,N_1939,N_1513);
or U4052 (N_4052,N_807,N_2121);
nand U4053 (N_4053,N_1166,N_436);
nor U4054 (N_4054,N_94,N_1947);
nand U4055 (N_4055,N_2334,N_359);
nand U4056 (N_4056,N_1462,N_2160);
nor U4057 (N_4057,N_961,N_1369);
or U4058 (N_4058,N_2399,N_916);
xor U4059 (N_4059,N_30,N_2361);
xor U4060 (N_4060,N_2256,N_1776);
nor U4061 (N_4061,N_381,N_1716);
xnor U4062 (N_4062,N_504,N_1788);
xor U4063 (N_4063,N_2197,N_1097);
or U4064 (N_4064,N_404,N_932);
nor U4065 (N_4065,N_1547,N_945);
nor U4066 (N_4066,N_2254,N_1545);
or U4067 (N_4067,N_1367,N_309);
or U4068 (N_4068,N_1659,N_345);
nor U4069 (N_4069,N_2384,N_219);
and U4070 (N_4070,N_1865,N_1592);
and U4071 (N_4071,N_645,N_1165);
nor U4072 (N_4072,N_464,N_2383);
nor U4073 (N_4073,N_844,N_649);
xor U4074 (N_4074,N_896,N_958);
or U4075 (N_4075,N_933,N_59);
xor U4076 (N_4076,N_1668,N_207);
or U4077 (N_4077,N_460,N_1343);
or U4078 (N_4078,N_929,N_1020);
nand U4079 (N_4079,N_878,N_904);
nand U4080 (N_4080,N_1974,N_533);
and U4081 (N_4081,N_1412,N_2071);
or U4082 (N_4082,N_1064,N_1464);
and U4083 (N_4083,N_2135,N_300);
nor U4084 (N_4084,N_2283,N_1218);
or U4085 (N_4085,N_716,N_1403);
nor U4086 (N_4086,N_2151,N_1637);
nand U4087 (N_4087,N_2153,N_1);
nor U4088 (N_4088,N_910,N_2384);
and U4089 (N_4089,N_478,N_739);
and U4090 (N_4090,N_1976,N_349);
and U4091 (N_4091,N_682,N_439);
and U4092 (N_4092,N_4,N_1069);
or U4093 (N_4093,N_2368,N_42);
xnor U4094 (N_4094,N_959,N_2205);
nor U4095 (N_4095,N_2073,N_916);
and U4096 (N_4096,N_651,N_1089);
and U4097 (N_4097,N_560,N_1852);
nor U4098 (N_4098,N_1274,N_306);
or U4099 (N_4099,N_2446,N_2437);
nor U4100 (N_4100,N_1613,N_1403);
nand U4101 (N_4101,N_960,N_537);
and U4102 (N_4102,N_903,N_1675);
nand U4103 (N_4103,N_1853,N_2219);
nor U4104 (N_4104,N_2025,N_1301);
nand U4105 (N_4105,N_1834,N_1534);
nand U4106 (N_4106,N_510,N_1954);
nor U4107 (N_4107,N_482,N_530);
nor U4108 (N_4108,N_2033,N_345);
and U4109 (N_4109,N_2440,N_2492);
nand U4110 (N_4110,N_1571,N_1932);
nand U4111 (N_4111,N_243,N_2307);
nor U4112 (N_4112,N_2274,N_1531);
and U4113 (N_4113,N_460,N_486);
nand U4114 (N_4114,N_1789,N_2025);
or U4115 (N_4115,N_1365,N_160);
nand U4116 (N_4116,N_2184,N_1326);
xor U4117 (N_4117,N_1245,N_9);
nor U4118 (N_4118,N_821,N_234);
or U4119 (N_4119,N_1038,N_32);
nor U4120 (N_4120,N_311,N_2318);
or U4121 (N_4121,N_306,N_693);
nor U4122 (N_4122,N_805,N_2359);
nor U4123 (N_4123,N_230,N_1923);
xnor U4124 (N_4124,N_1347,N_436);
and U4125 (N_4125,N_2186,N_1399);
nand U4126 (N_4126,N_338,N_784);
nand U4127 (N_4127,N_735,N_305);
nor U4128 (N_4128,N_1695,N_1277);
nand U4129 (N_4129,N_1474,N_706);
and U4130 (N_4130,N_2346,N_2407);
and U4131 (N_4131,N_1189,N_1958);
nor U4132 (N_4132,N_2341,N_1697);
xnor U4133 (N_4133,N_77,N_2324);
nor U4134 (N_4134,N_245,N_24);
nand U4135 (N_4135,N_794,N_1330);
nand U4136 (N_4136,N_1925,N_1768);
and U4137 (N_4137,N_2388,N_2061);
or U4138 (N_4138,N_656,N_493);
or U4139 (N_4139,N_1731,N_1043);
and U4140 (N_4140,N_464,N_2488);
nand U4141 (N_4141,N_1595,N_1981);
and U4142 (N_4142,N_126,N_1984);
and U4143 (N_4143,N_454,N_1117);
and U4144 (N_4144,N_2450,N_878);
nor U4145 (N_4145,N_1239,N_1548);
nor U4146 (N_4146,N_1545,N_358);
or U4147 (N_4147,N_1940,N_2195);
or U4148 (N_4148,N_1538,N_881);
nor U4149 (N_4149,N_145,N_340);
or U4150 (N_4150,N_1011,N_1364);
or U4151 (N_4151,N_364,N_201);
xor U4152 (N_4152,N_2227,N_1154);
nand U4153 (N_4153,N_2021,N_2388);
nand U4154 (N_4154,N_1352,N_1933);
nor U4155 (N_4155,N_1202,N_1341);
nor U4156 (N_4156,N_2058,N_1528);
and U4157 (N_4157,N_1075,N_223);
or U4158 (N_4158,N_1902,N_1635);
xnor U4159 (N_4159,N_1540,N_1616);
and U4160 (N_4160,N_342,N_1041);
or U4161 (N_4161,N_1507,N_612);
or U4162 (N_4162,N_947,N_2491);
nand U4163 (N_4163,N_204,N_2499);
nor U4164 (N_4164,N_548,N_511);
or U4165 (N_4165,N_2092,N_2323);
or U4166 (N_4166,N_2304,N_401);
xnor U4167 (N_4167,N_2220,N_228);
or U4168 (N_4168,N_1856,N_1635);
and U4169 (N_4169,N_1538,N_2384);
nor U4170 (N_4170,N_849,N_2411);
nand U4171 (N_4171,N_37,N_971);
xnor U4172 (N_4172,N_2325,N_2335);
and U4173 (N_4173,N_891,N_1788);
nand U4174 (N_4174,N_1973,N_946);
nand U4175 (N_4175,N_593,N_1810);
and U4176 (N_4176,N_383,N_1155);
and U4177 (N_4177,N_576,N_738);
or U4178 (N_4178,N_2369,N_2360);
nand U4179 (N_4179,N_2007,N_1860);
and U4180 (N_4180,N_251,N_1907);
xor U4181 (N_4181,N_1125,N_1136);
and U4182 (N_4182,N_310,N_1535);
nand U4183 (N_4183,N_168,N_1893);
and U4184 (N_4184,N_566,N_744);
or U4185 (N_4185,N_1656,N_1892);
and U4186 (N_4186,N_1619,N_1277);
xnor U4187 (N_4187,N_919,N_459);
or U4188 (N_4188,N_1502,N_688);
or U4189 (N_4189,N_655,N_73);
nor U4190 (N_4190,N_2454,N_2499);
xor U4191 (N_4191,N_2160,N_2041);
nor U4192 (N_4192,N_1991,N_1622);
nor U4193 (N_4193,N_289,N_1297);
or U4194 (N_4194,N_1712,N_1186);
or U4195 (N_4195,N_1274,N_2182);
nand U4196 (N_4196,N_1682,N_2215);
or U4197 (N_4197,N_1507,N_925);
nand U4198 (N_4198,N_1266,N_2335);
or U4199 (N_4199,N_2257,N_388);
nand U4200 (N_4200,N_2322,N_218);
or U4201 (N_4201,N_5,N_68);
and U4202 (N_4202,N_564,N_2102);
and U4203 (N_4203,N_1217,N_1406);
nor U4204 (N_4204,N_808,N_2278);
nand U4205 (N_4205,N_665,N_2451);
nor U4206 (N_4206,N_1560,N_2015);
and U4207 (N_4207,N_972,N_1582);
and U4208 (N_4208,N_578,N_2387);
xnor U4209 (N_4209,N_1676,N_2282);
and U4210 (N_4210,N_592,N_753);
or U4211 (N_4211,N_463,N_1091);
nor U4212 (N_4212,N_670,N_652);
xnor U4213 (N_4213,N_1076,N_1227);
nand U4214 (N_4214,N_2340,N_2036);
nor U4215 (N_4215,N_2184,N_1186);
and U4216 (N_4216,N_491,N_913);
and U4217 (N_4217,N_890,N_115);
or U4218 (N_4218,N_2327,N_200);
and U4219 (N_4219,N_2248,N_2465);
or U4220 (N_4220,N_1716,N_1329);
nor U4221 (N_4221,N_1672,N_2256);
nor U4222 (N_4222,N_239,N_184);
and U4223 (N_4223,N_907,N_164);
xnor U4224 (N_4224,N_1868,N_396);
nand U4225 (N_4225,N_923,N_424);
xnor U4226 (N_4226,N_1007,N_13);
xnor U4227 (N_4227,N_135,N_172);
nand U4228 (N_4228,N_2321,N_2318);
nor U4229 (N_4229,N_373,N_1914);
and U4230 (N_4230,N_312,N_824);
nand U4231 (N_4231,N_1383,N_700);
and U4232 (N_4232,N_1830,N_1716);
nor U4233 (N_4233,N_25,N_329);
nand U4234 (N_4234,N_623,N_351);
and U4235 (N_4235,N_625,N_2405);
or U4236 (N_4236,N_976,N_2299);
or U4237 (N_4237,N_1666,N_2111);
or U4238 (N_4238,N_670,N_959);
nor U4239 (N_4239,N_1597,N_656);
or U4240 (N_4240,N_256,N_1325);
and U4241 (N_4241,N_2462,N_2282);
nand U4242 (N_4242,N_653,N_488);
nand U4243 (N_4243,N_954,N_519);
or U4244 (N_4244,N_685,N_1531);
and U4245 (N_4245,N_1416,N_2211);
and U4246 (N_4246,N_1621,N_1903);
nand U4247 (N_4247,N_1248,N_1880);
nand U4248 (N_4248,N_972,N_574);
nor U4249 (N_4249,N_82,N_1139);
nor U4250 (N_4250,N_1626,N_354);
nor U4251 (N_4251,N_310,N_1213);
nand U4252 (N_4252,N_1559,N_1635);
nand U4253 (N_4253,N_110,N_591);
and U4254 (N_4254,N_1192,N_1649);
and U4255 (N_4255,N_893,N_1158);
nor U4256 (N_4256,N_881,N_764);
or U4257 (N_4257,N_613,N_128);
nand U4258 (N_4258,N_1212,N_2295);
or U4259 (N_4259,N_1992,N_1106);
or U4260 (N_4260,N_1050,N_1443);
and U4261 (N_4261,N_973,N_2310);
or U4262 (N_4262,N_1056,N_1229);
or U4263 (N_4263,N_2304,N_1233);
and U4264 (N_4264,N_1630,N_2039);
xnor U4265 (N_4265,N_2229,N_793);
xnor U4266 (N_4266,N_696,N_2237);
nor U4267 (N_4267,N_782,N_652);
xnor U4268 (N_4268,N_1751,N_1169);
and U4269 (N_4269,N_553,N_896);
nor U4270 (N_4270,N_890,N_1880);
nor U4271 (N_4271,N_1232,N_943);
nand U4272 (N_4272,N_1248,N_2160);
nor U4273 (N_4273,N_2430,N_2099);
nor U4274 (N_4274,N_2479,N_575);
or U4275 (N_4275,N_795,N_1705);
xnor U4276 (N_4276,N_540,N_2445);
and U4277 (N_4277,N_859,N_2475);
and U4278 (N_4278,N_2024,N_1476);
nor U4279 (N_4279,N_1959,N_1918);
nor U4280 (N_4280,N_721,N_2064);
and U4281 (N_4281,N_445,N_907);
nand U4282 (N_4282,N_1840,N_2384);
nor U4283 (N_4283,N_1324,N_319);
nand U4284 (N_4284,N_1032,N_1910);
and U4285 (N_4285,N_1892,N_751);
or U4286 (N_4286,N_747,N_659);
nand U4287 (N_4287,N_1022,N_949);
or U4288 (N_4288,N_1219,N_514);
nand U4289 (N_4289,N_3,N_2415);
and U4290 (N_4290,N_989,N_531);
and U4291 (N_4291,N_984,N_2080);
and U4292 (N_4292,N_966,N_143);
nor U4293 (N_4293,N_2094,N_189);
and U4294 (N_4294,N_1329,N_465);
or U4295 (N_4295,N_106,N_1863);
and U4296 (N_4296,N_1377,N_1727);
nor U4297 (N_4297,N_2273,N_1588);
or U4298 (N_4298,N_1252,N_820);
nand U4299 (N_4299,N_2257,N_2366);
and U4300 (N_4300,N_2079,N_1514);
and U4301 (N_4301,N_756,N_1205);
or U4302 (N_4302,N_129,N_1087);
or U4303 (N_4303,N_304,N_4);
nor U4304 (N_4304,N_1384,N_1842);
and U4305 (N_4305,N_230,N_2268);
or U4306 (N_4306,N_650,N_277);
or U4307 (N_4307,N_1124,N_507);
or U4308 (N_4308,N_1183,N_1759);
and U4309 (N_4309,N_1288,N_1176);
and U4310 (N_4310,N_2372,N_933);
nand U4311 (N_4311,N_1949,N_525);
nand U4312 (N_4312,N_891,N_292);
nor U4313 (N_4313,N_407,N_1398);
and U4314 (N_4314,N_1709,N_1646);
xnor U4315 (N_4315,N_243,N_322);
or U4316 (N_4316,N_1449,N_2493);
or U4317 (N_4317,N_378,N_275);
or U4318 (N_4318,N_2240,N_342);
and U4319 (N_4319,N_2459,N_1226);
nand U4320 (N_4320,N_868,N_634);
and U4321 (N_4321,N_1080,N_2380);
or U4322 (N_4322,N_2084,N_1501);
nor U4323 (N_4323,N_1448,N_2179);
nand U4324 (N_4324,N_347,N_31);
or U4325 (N_4325,N_1066,N_1780);
nor U4326 (N_4326,N_1458,N_432);
or U4327 (N_4327,N_733,N_750);
or U4328 (N_4328,N_342,N_1861);
nor U4329 (N_4329,N_2278,N_2133);
nand U4330 (N_4330,N_2087,N_1344);
and U4331 (N_4331,N_739,N_1213);
nor U4332 (N_4332,N_2062,N_2277);
or U4333 (N_4333,N_1149,N_1709);
or U4334 (N_4334,N_1805,N_2449);
nand U4335 (N_4335,N_2044,N_2344);
or U4336 (N_4336,N_350,N_1039);
xnor U4337 (N_4337,N_379,N_1366);
and U4338 (N_4338,N_96,N_1224);
nor U4339 (N_4339,N_869,N_1552);
xor U4340 (N_4340,N_620,N_2029);
or U4341 (N_4341,N_2164,N_1751);
xor U4342 (N_4342,N_2191,N_2334);
nand U4343 (N_4343,N_2112,N_1779);
or U4344 (N_4344,N_2458,N_428);
or U4345 (N_4345,N_650,N_31);
or U4346 (N_4346,N_74,N_1188);
nand U4347 (N_4347,N_458,N_1950);
nand U4348 (N_4348,N_534,N_2226);
nand U4349 (N_4349,N_2407,N_1468);
nand U4350 (N_4350,N_1039,N_715);
nor U4351 (N_4351,N_1500,N_1856);
xnor U4352 (N_4352,N_994,N_1557);
or U4353 (N_4353,N_1194,N_314);
xor U4354 (N_4354,N_982,N_1606);
nor U4355 (N_4355,N_2291,N_2343);
and U4356 (N_4356,N_610,N_956);
nor U4357 (N_4357,N_566,N_857);
or U4358 (N_4358,N_295,N_909);
and U4359 (N_4359,N_1421,N_746);
nor U4360 (N_4360,N_1387,N_2230);
nand U4361 (N_4361,N_803,N_1062);
xor U4362 (N_4362,N_2382,N_1264);
and U4363 (N_4363,N_1152,N_355);
xnor U4364 (N_4364,N_1788,N_2443);
and U4365 (N_4365,N_455,N_539);
or U4366 (N_4366,N_1839,N_650);
xnor U4367 (N_4367,N_1584,N_828);
or U4368 (N_4368,N_1715,N_1501);
or U4369 (N_4369,N_1003,N_1411);
nor U4370 (N_4370,N_323,N_1631);
nand U4371 (N_4371,N_860,N_2207);
and U4372 (N_4372,N_19,N_1610);
and U4373 (N_4373,N_1161,N_2153);
xnor U4374 (N_4374,N_963,N_76);
and U4375 (N_4375,N_1678,N_798);
nand U4376 (N_4376,N_1295,N_253);
nand U4377 (N_4377,N_1151,N_509);
nor U4378 (N_4378,N_834,N_1338);
and U4379 (N_4379,N_1510,N_1007);
and U4380 (N_4380,N_419,N_2309);
nor U4381 (N_4381,N_1788,N_1755);
nand U4382 (N_4382,N_360,N_1324);
nand U4383 (N_4383,N_52,N_67);
xnor U4384 (N_4384,N_1223,N_53);
or U4385 (N_4385,N_1433,N_234);
or U4386 (N_4386,N_364,N_808);
or U4387 (N_4387,N_1032,N_732);
or U4388 (N_4388,N_398,N_1593);
nor U4389 (N_4389,N_279,N_836);
nand U4390 (N_4390,N_995,N_1110);
nand U4391 (N_4391,N_608,N_2268);
and U4392 (N_4392,N_349,N_1798);
or U4393 (N_4393,N_913,N_665);
nand U4394 (N_4394,N_1000,N_127);
and U4395 (N_4395,N_1834,N_2456);
nor U4396 (N_4396,N_1999,N_1263);
or U4397 (N_4397,N_318,N_474);
nor U4398 (N_4398,N_2014,N_1138);
nand U4399 (N_4399,N_1795,N_2090);
nor U4400 (N_4400,N_906,N_2094);
nand U4401 (N_4401,N_1783,N_113);
nor U4402 (N_4402,N_1731,N_1806);
and U4403 (N_4403,N_2032,N_1619);
xnor U4404 (N_4404,N_740,N_134);
and U4405 (N_4405,N_816,N_547);
and U4406 (N_4406,N_91,N_2139);
and U4407 (N_4407,N_279,N_2106);
nand U4408 (N_4408,N_1177,N_383);
or U4409 (N_4409,N_1703,N_2261);
or U4410 (N_4410,N_2055,N_858);
or U4411 (N_4411,N_1426,N_1697);
xor U4412 (N_4412,N_666,N_1926);
nand U4413 (N_4413,N_2240,N_2148);
or U4414 (N_4414,N_2296,N_655);
xor U4415 (N_4415,N_1631,N_484);
or U4416 (N_4416,N_2290,N_777);
or U4417 (N_4417,N_1111,N_150);
nand U4418 (N_4418,N_1966,N_1319);
nand U4419 (N_4419,N_161,N_171);
nand U4420 (N_4420,N_2171,N_2370);
nor U4421 (N_4421,N_1774,N_1823);
and U4422 (N_4422,N_2077,N_305);
nand U4423 (N_4423,N_1476,N_993);
nand U4424 (N_4424,N_361,N_1228);
and U4425 (N_4425,N_887,N_1555);
nor U4426 (N_4426,N_255,N_469);
or U4427 (N_4427,N_2307,N_1877);
nand U4428 (N_4428,N_1927,N_1756);
xnor U4429 (N_4429,N_1053,N_301);
nand U4430 (N_4430,N_1847,N_212);
or U4431 (N_4431,N_483,N_1483);
or U4432 (N_4432,N_1277,N_1640);
or U4433 (N_4433,N_1135,N_451);
nor U4434 (N_4434,N_833,N_133);
nor U4435 (N_4435,N_1556,N_1640);
and U4436 (N_4436,N_1936,N_1130);
or U4437 (N_4437,N_250,N_1879);
or U4438 (N_4438,N_1465,N_450);
nor U4439 (N_4439,N_832,N_729);
nand U4440 (N_4440,N_1771,N_76);
nor U4441 (N_4441,N_1783,N_1164);
nand U4442 (N_4442,N_577,N_1953);
or U4443 (N_4443,N_920,N_2471);
nor U4444 (N_4444,N_387,N_1048);
nand U4445 (N_4445,N_2318,N_26);
nor U4446 (N_4446,N_35,N_212);
nor U4447 (N_4447,N_92,N_757);
nor U4448 (N_4448,N_2111,N_1458);
nand U4449 (N_4449,N_249,N_159);
nor U4450 (N_4450,N_519,N_396);
nand U4451 (N_4451,N_1671,N_446);
and U4452 (N_4452,N_19,N_937);
nand U4453 (N_4453,N_1363,N_959);
xnor U4454 (N_4454,N_467,N_899);
or U4455 (N_4455,N_1582,N_505);
nand U4456 (N_4456,N_1662,N_269);
and U4457 (N_4457,N_1822,N_2192);
or U4458 (N_4458,N_761,N_2044);
and U4459 (N_4459,N_2066,N_1313);
and U4460 (N_4460,N_18,N_661);
nor U4461 (N_4461,N_371,N_2083);
nand U4462 (N_4462,N_1562,N_1721);
nor U4463 (N_4463,N_1362,N_982);
or U4464 (N_4464,N_1372,N_1899);
or U4465 (N_4465,N_1939,N_2497);
nand U4466 (N_4466,N_1456,N_2053);
or U4467 (N_4467,N_1420,N_562);
or U4468 (N_4468,N_125,N_1276);
nor U4469 (N_4469,N_2318,N_1162);
nor U4470 (N_4470,N_2217,N_939);
nand U4471 (N_4471,N_2128,N_531);
nor U4472 (N_4472,N_2364,N_652);
xnor U4473 (N_4473,N_1114,N_2353);
or U4474 (N_4474,N_2376,N_447);
and U4475 (N_4475,N_1021,N_1643);
nand U4476 (N_4476,N_432,N_2258);
or U4477 (N_4477,N_434,N_403);
xnor U4478 (N_4478,N_1117,N_1162);
and U4479 (N_4479,N_1073,N_167);
nor U4480 (N_4480,N_1406,N_1806);
or U4481 (N_4481,N_1535,N_335);
nor U4482 (N_4482,N_712,N_773);
nor U4483 (N_4483,N_1077,N_224);
xnor U4484 (N_4484,N_437,N_2385);
or U4485 (N_4485,N_1712,N_1953);
xnor U4486 (N_4486,N_2307,N_712);
or U4487 (N_4487,N_1246,N_675);
nor U4488 (N_4488,N_1772,N_918);
nand U4489 (N_4489,N_942,N_1675);
or U4490 (N_4490,N_98,N_442);
and U4491 (N_4491,N_1767,N_2348);
xor U4492 (N_4492,N_1845,N_2396);
xnor U4493 (N_4493,N_712,N_2155);
nor U4494 (N_4494,N_1662,N_1902);
nor U4495 (N_4495,N_1208,N_1495);
nor U4496 (N_4496,N_61,N_1163);
nand U4497 (N_4497,N_17,N_1449);
or U4498 (N_4498,N_1806,N_1247);
and U4499 (N_4499,N_2327,N_2097);
nor U4500 (N_4500,N_916,N_2412);
xnor U4501 (N_4501,N_1792,N_2261);
nand U4502 (N_4502,N_1373,N_1473);
xnor U4503 (N_4503,N_8,N_1139);
nor U4504 (N_4504,N_1238,N_2496);
xnor U4505 (N_4505,N_580,N_1554);
or U4506 (N_4506,N_2494,N_1679);
xor U4507 (N_4507,N_342,N_100);
nor U4508 (N_4508,N_1681,N_137);
nand U4509 (N_4509,N_873,N_515);
and U4510 (N_4510,N_1328,N_110);
nor U4511 (N_4511,N_91,N_1423);
and U4512 (N_4512,N_467,N_37);
nand U4513 (N_4513,N_620,N_286);
or U4514 (N_4514,N_523,N_2409);
nand U4515 (N_4515,N_204,N_1245);
nand U4516 (N_4516,N_2135,N_1215);
nand U4517 (N_4517,N_1108,N_53);
or U4518 (N_4518,N_1647,N_1033);
nor U4519 (N_4519,N_320,N_1023);
or U4520 (N_4520,N_2027,N_2319);
nand U4521 (N_4521,N_892,N_1590);
xor U4522 (N_4522,N_2241,N_554);
and U4523 (N_4523,N_2432,N_1366);
nor U4524 (N_4524,N_1237,N_813);
or U4525 (N_4525,N_1946,N_108);
nor U4526 (N_4526,N_1485,N_2463);
nor U4527 (N_4527,N_669,N_1772);
and U4528 (N_4528,N_1805,N_1272);
nor U4529 (N_4529,N_1758,N_1826);
nor U4530 (N_4530,N_1654,N_875);
nor U4531 (N_4531,N_335,N_1628);
or U4532 (N_4532,N_584,N_2130);
nand U4533 (N_4533,N_2330,N_2008);
and U4534 (N_4534,N_2226,N_1386);
nand U4535 (N_4535,N_1736,N_62);
nor U4536 (N_4536,N_2000,N_1687);
xnor U4537 (N_4537,N_2155,N_763);
nor U4538 (N_4538,N_108,N_2362);
or U4539 (N_4539,N_1917,N_15);
nand U4540 (N_4540,N_432,N_565);
nor U4541 (N_4541,N_2295,N_2065);
or U4542 (N_4542,N_1530,N_421);
nor U4543 (N_4543,N_1465,N_585);
xnor U4544 (N_4544,N_1962,N_1168);
and U4545 (N_4545,N_795,N_1179);
nor U4546 (N_4546,N_1195,N_487);
or U4547 (N_4547,N_1570,N_1539);
and U4548 (N_4548,N_832,N_2057);
and U4549 (N_4549,N_1625,N_155);
or U4550 (N_4550,N_801,N_2455);
and U4551 (N_4551,N_1545,N_636);
and U4552 (N_4552,N_1051,N_788);
nand U4553 (N_4553,N_620,N_674);
or U4554 (N_4554,N_790,N_1637);
nand U4555 (N_4555,N_1170,N_580);
nand U4556 (N_4556,N_2092,N_686);
nor U4557 (N_4557,N_1491,N_1074);
nor U4558 (N_4558,N_892,N_1033);
nand U4559 (N_4559,N_1282,N_2173);
nor U4560 (N_4560,N_2389,N_1363);
and U4561 (N_4561,N_64,N_308);
nand U4562 (N_4562,N_290,N_398);
and U4563 (N_4563,N_2269,N_525);
and U4564 (N_4564,N_2082,N_868);
nand U4565 (N_4565,N_2290,N_2020);
nor U4566 (N_4566,N_1607,N_2193);
and U4567 (N_4567,N_2056,N_299);
or U4568 (N_4568,N_670,N_2379);
nor U4569 (N_4569,N_1740,N_2060);
or U4570 (N_4570,N_143,N_1987);
or U4571 (N_4571,N_1726,N_121);
nand U4572 (N_4572,N_1541,N_444);
nor U4573 (N_4573,N_511,N_1775);
and U4574 (N_4574,N_1433,N_569);
xnor U4575 (N_4575,N_683,N_179);
nor U4576 (N_4576,N_1823,N_1355);
or U4577 (N_4577,N_2174,N_310);
xor U4578 (N_4578,N_201,N_509);
or U4579 (N_4579,N_407,N_685);
or U4580 (N_4580,N_1750,N_1473);
nand U4581 (N_4581,N_2012,N_556);
nor U4582 (N_4582,N_1561,N_1772);
and U4583 (N_4583,N_17,N_1316);
nor U4584 (N_4584,N_283,N_753);
or U4585 (N_4585,N_594,N_1055);
and U4586 (N_4586,N_255,N_991);
xnor U4587 (N_4587,N_1169,N_588);
and U4588 (N_4588,N_2169,N_562);
nor U4589 (N_4589,N_2421,N_1081);
nand U4590 (N_4590,N_47,N_1973);
xnor U4591 (N_4591,N_1061,N_2275);
and U4592 (N_4592,N_2114,N_2438);
nor U4593 (N_4593,N_828,N_1972);
or U4594 (N_4594,N_698,N_1394);
nand U4595 (N_4595,N_283,N_361);
or U4596 (N_4596,N_1572,N_1203);
and U4597 (N_4597,N_603,N_1200);
nand U4598 (N_4598,N_725,N_881);
nor U4599 (N_4599,N_1418,N_85);
nor U4600 (N_4600,N_215,N_1491);
or U4601 (N_4601,N_927,N_404);
or U4602 (N_4602,N_2407,N_94);
and U4603 (N_4603,N_2048,N_2112);
nor U4604 (N_4604,N_1315,N_1939);
or U4605 (N_4605,N_4,N_827);
nand U4606 (N_4606,N_639,N_645);
and U4607 (N_4607,N_387,N_1515);
nor U4608 (N_4608,N_1127,N_1480);
or U4609 (N_4609,N_1691,N_178);
nor U4610 (N_4610,N_2421,N_81);
or U4611 (N_4611,N_647,N_2393);
xor U4612 (N_4612,N_1540,N_1479);
nor U4613 (N_4613,N_102,N_2173);
or U4614 (N_4614,N_2299,N_124);
nor U4615 (N_4615,N_2196,N_1456);
nor U4616 (N_4616,N_1205,N_193);
nand U4617 (N_4617,N_2107,N_1943);
or U4618 (N_4618,N_648,N_2354);
and U4619 (N_4619,N_695,N_998);
and U4620 (N_4620,N_602,N_1177);
nand U4621 (N_4621,N_410,N_603);
xor U4622 (N_4622,N_782,N_1890);
or U4623 (N_4623,N_2204,N_272);
nor U4624 (N_4624,N_987,N_1114);
or U4625 (N_4625,N_2472,N_1352);
nor U4626 (N_4626,N_2303,N_1170);
nor U4627 (N_4627,N_626,N_1535);
nor U4628 (N_4628,N_764,N_1770);
and U4629 (N_4629,N_2123,N_692);
and U4630 (N_4630,N_2107,N_1071);
nand U4631 (N_4631,N_160,N_1549);
and U4632 (N_4632,N_1717,N_530);
nor U4633 (N_4633,N_188,N_1480);
nand U4634 (N_4634,N_611,N_2094);
and U4635 (N_4635,N_1225,N_273);
and U4636 (N_4636,N_518,N_1242);
nor U4637 (N_4637,N_1464,N_1275);
nand U4638 (N_4638,N_31,N_285);
nand U4639 (N_4639,N_79,N_1959);
nand U4640 (N_4640,N_545,N_1011);
nand U4641 (N_4641,N_955,N_137);
xnor U4642 (N_4642,N_187,N_2144);
nor U4643 (N_4643,N_1579,N_947);
and U4644 (N_4644,N_372,N_1576);
nand U4645 (N_4645,N_2232,N_1016);
and U4646 (N_4646,N_2330,N_1733);
or U4647 (N_4647,N_331,N_178);
nand U4648 (N_4648,N_2484,N_457);
nor U4649 (N_4649,N_330,N_2173);
nor U4650 (N_4650,N_712,N_143);
nand U4651 (N_4651,N_1276,N_517);
nor U4652 (N_4652,N_1049,N_323);
or U4653 (N_4653,N_501,N_657);
nand U4654 (N_4654,N_759,N_1903);
nor U4655 (N_4655,N_65,N_1163);
and U4656 (N_4656,N_1567,N_1070);
and U4657 (N_4657,N_1541,N_1402);
or U4658 (N_4658,N_1940,N_509);
or U4659 (N_4659,N_945,N_1460);
xnor U4660 (N_4660,N_235,N_1061);
or U4661 (N_4661,N_2382,N_732);
or U4662 (N_4662,N_2216,N_1813);
nand U4663 (N_4663,N_1005,N_1755);
nand U4664 (N_4664,N_1941,N_971);
xor U4665 (N_4665,N_953,N_2039);
nand U4666 (N_4666,N_732,N_531);
or U4667 (N_4667,N_2485,N_805);
xnor U4668 (N_4668,N_1577,N_253);
or U4669 (N_4669,N_1912,N_394);
or U4670 (N_4670,N_1543,N_1973);
and U4671 (N_4671,N_1283,N_140);
or U4672 (N_4672,N_1375,N_331);
and U4673 (N_4673,N_1687,N_619);
xor U4674 (N_4674,N_1575,N_2278);
nand U4675 (N_4675,N_1204,N_1761);
or U4676 (N_4676,N_2345,N_695);
and U4677 (N_4677,N_212,N_463);
and U4678 (N_4678,N_29,N_1454);
nor U4679 (N_4679,N_1778,N_1076);
or U4680 (N_4680,N_1380,N_1675);
nor U4681 (N_4681,N_1017,N_2178);
nand U4682 (N_4682,N_2199,N_2095);
and U4683 (N_4683,N_612,N_757);
nor U4684 (N_4684,N_1386,N_817);
xnor U4685 (N_4685,N_295,N_1731);
nor U4686 (N_4686,N_1192,N_1030);
nor U4687 (N_4687,N_2435,N_1056);
nand U4688 (N_4688,N_2016,N_1953);
nor U4689 (N_4689,N_2009,N_1646);
nor U4690 (N_4690,N_1358,N_1895);
nand U4691 (N_4691,N_1637,N_274);
or U4692 (N_4692,N_1744,N_433);
and U4693 (N_4693,N_536,N_1519);
or U4694 (N_4694,N_1650,N_1647);
nand U4695 (N_4695,N_1226,N_2246);
nor U4696 (N_4696,N_2338,N_2317);
nand U4697 (N_4697,N_2406,N_2141);
or U4698 (N_4698,N_1887,N_1197);
nand U4699 (N_4699,N_77,N_2259);
and U4700 (N_4700,N_1072,N_672);
nand U4701 (N_4701,N_2212,N_2098);
nor U4702 (N_4702,N_2354,N_1341);
nand U4703 (N_4703,N_2174,N_908);
nand U4704 (N_4704,N_1726,N_281);
nand U4705 (N_4705,N_1226,N_1288);
and U4706 (N_4706,N_1562,N_2402);
xor U4707 (N_4707,N_2143,N_2331);
nand U4708 (N_4708,N_338,N_117);
or U4709 (N_4709,N_605,N_2477);
or U4710 (N_4710,N_2245,N_2019);
nand U4711 (N_4711,N_2326,N_806);
or U4712 (N_4712,N_1760,N_129);
and U4713 (N_4713,N_1391,N_394);
and U4714 (N_4714,N_1073,N_976);
xnor U4715 (N_4715,N_58,N_625);
or U4716 (N_4716,N_1687,N_705);
nor U4717 (N_4717,N_717,N_1773);
or U4718 (N_4718,N_193,N_2346);
nor U4719 (N_4719,N_1395,N_1301);
and U4720 (N_4720,N_2186,N_1574);
nor U4721 (N_4721,N_564,N_960);
nand U4722 (N_4722,N_971,N_1723);
or U4723 (N_4723,N_744,N_1777);
nor U4724 (N_4724,N_1692,N_1852);
and U4725 (N_4725,N_2172,N_4);
or U4726 (N_4726,N_1541,N_864);
and U4727 (N_4727,N_1453,N_2077);
or U4728 (N_4728,N_255,N_2384);
nor U4729 (N_4729,N_2305,N_99);
and U4730 (N_4730,N_1233,N_1694);
xnor U4731 (N_4731,N_1441,N_1230);
nor U4732 (N_4732,N_1848,N_160);
and U4733 (N_4733,N_2434,N_1049);
nand U4734 (N_4734,N_594,N_1450);
and U4735 (N_4735,N_1093,N_1807);
xnor U4736 (N_4736,N_468,N_2003);
nor U4737 (N_4737,N_1372,N_1911);
nand U4738 (N_4738,N_1350,N_1885);
nor U4739 (N_4739,N_2475,N_2363);
and U4740 (N_4740,N_2313,N_1486);
nand U4741 (N_4741,N_2064,N_1701);
nor U4742 (N_4742,N_1987,N_2401);
or U4743 (N_4743,N_2367,N_467);
or U4744 (N_4744,N_1542,N_1152);
or U4745 (N_4745,N_2319,N_226);
or U4746 (N_4746,N_1406,N_1342);
nand U4747 (N_4747,N_42,N_2338);
and U4748 (N_4748,N_405,N_1272);
or U4749 (N_4749,N_1230,N_658);
and U4750 (N_4750,N_211,N_1022);
and U4751 (N_4751,N_491,N_401);
xor U4752 (N_4752,N_1633,N_675);
and U4753 (N_4753,N_1990,N_12);
or U4754 (N_4754,N_398,N_762);
nand U4755 (N_4755,N_2444,N_365);
or U4756 (N_4756,N_4,N_1806);
nand U4757 (N_4757,N_1013,N_447);
and U4758 (N_4758,N_1344,N_1508);
nand U4759 (N_4759,N_1837,N_1382);
and U4760 (N_4760,N_1316,N_1059);
nand U4761 (N_4761,N_2151,N_1932);
or U4762 (N_4762,N_737,N_1123);
xor U4763 (N_4763,N_112,N_1427);
nor U4764 (N_4764,N_153,N_609);
nand U4765 (N_4765,N_2248,N_984);
nand U4766 (N_4766,N_2063,N_442);
nand U4767 (N_4767,N_641,N_463);
nand U4768 (N_4768,N_1246,N_228);
or U4769 (N_4769,N_227,N_1443);
nand U4770 (N_4770,N_1450,N_1362);
nand U4771 (N_4771,N_451,N_845);
and U4772 (N_4772,N_2321,N_1274);
nor U4773 (N_4773,N_1238,N_1653);
nor U4774 (N_4774,N_747,N_2287);
or U4775 (N_4775,N_185,N_429);
nor U4776 (N_4776,N_1450,N_237);
nor U4777 (N_4777,N_79,N_2192);
nand U4778 (N_4778,N_1424,N_674);
nor U4779 (N_4779,N_124,N_874);
or U4780 (N_4780,N_1823,N_439);
nand U4781 (N_4781,N_42,N_1885);
nor U4782 (N_4782,N_1367,N_1258);
or U4783 (N_4783,N_1622,N_447);
nand U4784 (N_4784,N_1574,N_2026);
and U4785 (N_4785,N_1664,N_2436);
nand U4786 (N_4786,N_1779,N_2334);
nand U4787 (N_4787,N_1936,N_36);
or U4788 (N_4788,N_1568,N_1100);
and U4789 (N_4789,N_381,N_2416);
nand U4790 (N_4790,N_1309,N_990);
and U4791 (N_4791,N_1309,N_1540);
xor U4792 (N_4792,N_1814,N_1020);
nor U4793 (N_4793,N_2006,N_890);
or U4794 (N_4794,N_560,N_943);
or U4795 (N_4795,N_614,N_762);
nor U4796 (N_4796,N_2372,N_886);
nor U4797 (N_4797,N_73,N_1237);
xor U4798 (N_4798,N_546,N_388);
or U4799 (N_4799,N_848,N_589);
nor U4800 (N_4800,N_968,N_1560);
or U4801 (N_4801,N_101,N_203);
nand U4802 (N_4802,N_723,N_1687);
nor U4803 (N_4803,N_1959,N_966);
nand U4804 (N_4804,N_76,N_842);
or U4805 (N_4805,N_1712,N_2469);
or U4806 (N_4806,N_835,N_1140);
nor U4807 (N_4807,N_1111,N_216);
nor U4808 (N_4808,N_1154,N_2207);
or U4809 (N_4809,N_2401,N_203);
nor U4810 (N_4810,N_621,N_2269);
and U4811 (N_4811,N_1698,N_854);
nor U4812 (N_4812,N_1984,N_1590);
xor U4813 (N_4813,N_2002,N_884);
and U4814 (N_4814,N_2192,N_1641);
nand U4815 (N_4815,N_2193,N_1860);
nor U4816 (N_4816,N_2451,N_1989);
or U4817 (N_4817,N_1610,N_2295);
nand U4818 (N_4818,N_2331,N_401);
nand U4819 (N_4819,N_2421,N_1631);
nor U4820 (N_4820,N_32,N_950);
and U4821 (N_4821,N_1738,N_2493);
and U4822 (N_4822,N_1686,N_1114);
xor U4823 (N_4823,N_135,N_1006);
nor U4824 (N_4824,N_1535,N_656);
xnor U4825 (N_4825,N_1366,N_138);
nand U4826 (N_4826,N_463,N_1486);
or U4827 (N_4827,N_1395,N_1485);
nor U4828 (N_4828,N_32,N_2244);
nand U4829 (N_4829,N_2331,N_1374);
nor U4830 (N_4830,N_1918,N_1977);
nor U4831 (N_4831,N_1716,N_145);
or U4832 (N_4832,N_250,N_1016);
nor U4833 (N_4833,N_2389,N_1813);
nand U4834 (N_4834,N_882,N_2273);
nor U4835 (N_4835,N_1206,N_1475);
and U4836 (N_4836,N_1103,N_828);
or U4837 (N_4837,N_1987,N_831);
nand U4838 (N_4838,N_517,N_166);
or U4839 (N_4839,N_195,N_246);
or U4840 (N_4840,N_2356,N_1391);
and U4841 (N_4841,N_871,N_799);
and U4842 (N_4842,N_2336,N_712);
and U4843 (N_4843,N_1853,N_855);
or U4844 (N_4844,N_1019,N_2406);
or U4845 (N_4845,N_1948,N_1649);
xnor U4846 (N_4846,N_76,N_371);
or U4847 (N_4847,N_2441,N_1285);
and U4848 (N_4848,N_1364,N_543);
or U4849 (N_4849,N_1824,N_459);
nand U4850 (N_4850,N_1602,N_1889);
and U4851 (N_4851,N_1066,N_1165);
xnor U4852 (N_4852,N_788,N_1946);
and U4853 (N_4853,N_1549,N_879);
or U4854 (N_4854,N_1155,N_27);
nor U4855 (N_4855,N_1031,N_1004);
nand U4856 (N_4856,N_1629,N_802);
nor U4857 (N_4857,N_971,N_89);
and U4858 (N_4858,N_2461,N_895);
nand U4859 (N_4859,N_149,N_807);
or U4860 (N_4860,N_1952,N_2066);
nand U4861 (N_4861,N_914,N_1440);
nand U4862 (N_4862,N_1137,N_1486);
nand U4863 (N_4863,N_432,N_2241);
or U4864 (N_4864,N_1592,N_2122);
or U4865 (N_4865,N_1050,N_108);
or U4866 (N_4866,N_1914,N_80);
xnor U4867 (N_4867,N_1888,N_328);
or U4868 (N_4868,N_2446,N_376);
and U4869 (N_4869,N_1225,N_211);
xnor U4870 (N_4870,N_1835,N_749);
nand U4871 (N_4871,N_701,N_1661);
and U4872 (N_4872,N_1499,N_1156);
nor U4873 (N_4873,N_1376,N_145);
nand U4874 (N_4874,N_891,N_1771);
or U4875 (N_4875,N_1224,N_2090);
or U4876 (N_4876,N_1303,N_798);
and U4877 (N_4877,N_2183,N_236);
nand U4878 (N_4878,N_177,N_1357);
nand U4879 (N_4879,N_2316,N_332);
and U4880 (N_4880,N_92,N_774);
nand U4881 (N_4881,N_534,N_1953);
or U4882 (N_4882,N_2107,N_1425);
and U4883 (N_4883,N_1535,N_497);
xor U4884 (N_4884,N_1039,N_193);
and U4885 (N_4885,N_2137,N_475);
nor U4886 (N_4886,N_151,N_1147);
nor U4887 (N_4887,N_765,N_117);
nand U4888 (N_4888,N_2367,N_220);
nor U4889 (N_4889,N_1887,N_1093);
or U4890 (N_4890,N_2436,N_1379);
nor U4891 (N_4891,N_1773,N_2229);
or U4892 (N_4892,N_817,N_2350);
and U4893 (N_4893,N_491,N_798);
and U4894 (N_4894,N_60,N_2243);
or U4895 (N_4895,N_2417,N_610);
xor U4896 (N_4896,N_2439,N_1988);
nand U4897 (N_4897,N_397,N_298);
or U4898 (N_4898,N_209,N_1320);
nand U4899 (N_4899,N_1520,N_869);
nand U4900 (N_4900,N_1879,N_1895);
nand U4901 (N_4901,N_1695,N_1823);
or U4902 (N_4902,N_1981,N_983);
and U4903 (N_4903,N_2359,N_290);
nand U4904 (N_4904,N_2363,N_2319);
or U4905 (N_4905,N_988,N_679);
nor U4906 (N_4906,N_1821,N_679);
or U4907 (N_4907,N_1409,N_2087);
nor U4908 (N_4908,N_322,N_1117);
xnor U4909 (N_4909,N_1855,N_1893);
xor U4910 (N_4910,N_2064,N_867);
nand U4911 (N_4911,N_1961,N_1964);
or U4912 (N_4912,N_1803,N_282);
xor U4913 (N_4913,N_920,N_803);
or U4914 (N_4914,N_1340,N_588);
or U4915 (N_4915,N_1306,N_1992);
nand U4916 (N_4916,N_2317,N_1571);
and U4917 (N_4917,N_362,N_1872);
nor U4918 (N_4918,N_2001,N_748);
and U4919 (N_4919,N_429,N_1772);
or U4920 (N_4920,N_977,N_1257);
or U4921 (N_4921,N_178,N_1967);
or U4922 (N_4922,N_1339,N_1380);
nor U4923 (N_4923,N_1285,N_879);
nor U4924 (N_4924,N_1910,N_2031);
and U4925 (N_4925,N_1979,N_674);
and U4926 (N_4926,N_1240,N_289);
nand U4927 (N_4927,N_841,N_1384);
nor U4928 (N_4928,N_2315,N_1984);
nor U4929 (N_4929,N_2476,N_2424);
and U4930 (N_4930,N_2219,N_1897);
nand U4931 (N_4931,N_1214,N_1856);
and U4932 (N_4932,N_1390,N_1947);
xnor U4933 (N_4933,N_1349,N_989);
nand U4934 (N_4934,N_873,N_1198);
xor U4935 (N_4935,N_1824,N_1779);
nor U4936 (N_4936,N_311,N_132);
nor U4937 (N_4937,N_44,N_1410);
and U4938 (N_4938,N_1028,N_1753);
xor U4939 (N_4939,N_1781,N_1510);
xor U4940 (N_4940,N_2232,N_166);
nor U4941 (N_4941,N_1337,N_39);
nor U4942 (N_4942,N_7,N_1970);
nor U4943 (N_4943,N_1498,N_1888);
nor U4944 (N_4944,N_1732,N_1935);
and U4945 (N_4945,N_1718,N_829);
or U4946 (N_4946,N_496,N_974);
or U4947 (N_4947,N_2141,N_1887);
nor U4948 (N_4948,N_406,N_2412);
xor U4949 (N_4949,N_186,N_1374);
nand U4950 (N_4950,N_529,N_1797);
nor U4951 (N_4951,N_951,N_2244);
nor U4952 (N_4952,N_109,N_907);
nor U4953 (N_4953,N_1030,N_1566);
nor U4954 (N_4954,N_1081,N_474);
xor U4955 (N_4955,N_744,N_1514);
nand U4956 (N_4956,N_2252,N_1018);
or U4957 (N_4957,N_1549,N_535);
and U4958 (N_4958,N_2465,N_1807);
and U4959 (N_4959,N_2179,N_1096);
nor U4960 (N_4960,N_2314,N_417);
nor U4961 (N_4961,N_1669,N_1555);
nand U4962 (N_4962,N_449,N_887);
nand U4963 (N_4963,N_495,N_423);
nor U4964 (N_4964,N_322,N_1588);
xor U4965 (N_4965,N_741,N_1115);
nand U4966 (N_4966,N_765,N_1820);
nand U4967 (N_4967,N_2148,N_406);
nor U4968 (N_4968,N_577,N_1027);
or U4969 (N_4969,N_1004,N_2312);
nor U4970 (N_4970,N_450,N_2427);
nor U4971 (N_4971,N_2258,N_2179);
xor U4972 (N_4972,N_686,N_1485);
and U4973 (N_4973,N_339,N_2034);
and U4974 (N_4974,N_409,N_288);
and U4975 (N_4975,N_1822,N_925);
and U4976 (N_4976,N_183,N_1157);
or U4977 (N_4977,N_2221,N_104);
or U4978 (N_4978,N_1062,N_1185);
or U4979 (N_4979,N_374,N_1767);
nand U4980 (N_4980,N_2357,N_203);
nand U4981 (N_4981,N_1321,N_1951);
nor U4982 (N_4982,N_1877,N_372);
and U4983 (N_4983,N_1722,N_2158);
and U4984 (N_4984,N_2494,N_2210);
or U4985 (N_4985,N_2162,N_1191);
or U4986 (N_4986,N_1290,N_1271);
and U4987 (N_4987,N_2439,N_73);
xor U4988 (N_4988,N_2234,N_646);
or U4989 (N_4989,N_65,N_1205);
nand U4990 (N_4990,N_199,N_1);
nor U4991 (N_4991,N_1917,N_52);
nand U4992 (N_4992,N_2421,N_724);
or U4993 (N_4993,N_508,N_702);
xor U4994 (N_4994,N_2238,N_1135);
and U4995 (N_4995,N_526,N_1187);
or U4996 (N_4996,N_1589,N_1551);
or U4997 (N_4997,N_1521,N_386);
or U4998 (N_4998,N_399,N_736);
and U4999 (N_4999,N_31,N_1544);
or U5000 (N_5000,N_4863,N_3372);
nand U5001 (N_5001,N_4008,N_3390);
nor U5002 (N_5002,N_3504,N_2523);
and U5003 (N_5003,N_4480,N_4819);
nand U5004 (N_5004,N_4133,N_3286);
or U5005 (N_5005,N_4506,N_3215);
or U5006 (N_5006,N_2634,N_2561);
nor U5007 (N_5007,N_4104,N_2677);
nand U5008 (N_5008,N_4013,N_2831);
and U5009 (N_5009,N_3627,N_4259);
and U5010 (N_5010,N_2618,N_4289);
nor U5011 (N_5011,N_4494,N_4434);
nor U5012 (N_5012,N_2579,N_4595);
nor U5013 (N_5013,N_3691,N_4323);
xor U5014 (N_5014,N_4002,N_3053);
or U5015 (N_5015,N_3196,N_3022);
nor U5016 (N_5016,N_3265,N_4797);
nor U5017 (N_5017,N_4182,N_4937);
or U5018 (N_5018,N_4324,N_3400);
nand U5019 (N_5019,N_3929,N_2856);
nand U5020 (N_5020,N_4060,N_2527);
and U5021 (N_5021,N_4774,N_3897);
or U5022 (N_5022,N_4602,N_4792);
nor U5023 (N_5023,N_4743,N_3997);
nor U5024 (N_5024,N_2626,N_3718);
nand U5025 (N_5025,N_3157,N_2845);
nor U5026 (N_5026,N_2762,N_4537);
xnor U5027 (N_5027,N_4096,N_3379);
nand U5028 (N_5028,N_2718,N_2966);
or U5029 (N_5029,N_4229,N_3001);
nor U5030 (N_5030,N_4688,N_4955);
nand U5031 (N_5031,N_3099,N_3154);
and U5032 (N_5032,N_2751,N_3825);
nor U5033 (N_5033,N_4644,N_2591);
nor U5034 (N_5034,N_3738,N_2895);
or U5035 (N_5035,N_4714,N_4226);
nand U5036 (N_5036,N_2608,N_2918);
nor U5037 (N_5037,N_2536,N_2597);
nand U5038 (N_5038,N_4985,N_3343);
and U5039 (N_5039,N_2729,N_3123);
and U5040 (N_5040,N_4521,N_2935);
nor U5041 (N_5041,N_3931,N_4460);
xnor U5042 (N_5042,N_3431,N_2875);
and U5043 (N_5043,N_3850,N_3785);
nor U5044 (N_5044,N_4252,N_3064);
nor U5045 (N_5045,N_2892,N_3707);
or U5046 (N_5046,N_4131,N_3981);
or U5047 (N_5047,N_4691,N_4603);
or U5048 (N_5048,N_4575,N_3571);
nor U5049 (N_5049,N_3685,N_2938);
or U5050 (N_5050,N_3056,N_3983);
and U5051 (N_5051,N_2983,N_4637);
nor U5052 (N_5052,N_4782,N_2768);
nand U5053 (N_5053,N_4286,N_3568);
and U5054 (N_5054,N_3086,N_4940);
nand U5055 (N_5055,N_4152,N_4250);
xnor U5056 (N_5056,N_3529,N_3821);
nor U5057 (N_5057,N_4938,N_2843);
xor U5058 (N_5058,N_3605,N_4146);
nor U5059 (N_5059,N_3739,N_2596);
and U5060 (N_5060,N_4911,N_4206);
nand U5061 (N_5061,N_3153,N_2642);
nor U5062 (N_5062,N_3410,N_4658);
or U5063 (N_5063,N_3904,N_3641);
nand U5064 (N_5064,N_2848,N_4209);
and U5065 (N_5065,N_3509,N_3580);
nand U5066 (N_5066,N_4172,N_4543);
and U5067 (N_5067,N_4760,N_4636);
and U5068 (N_5068,N_2940,N_3798);
xor U5069 (N_5069,N_4785,N_3299);
xnor U5070 (N_5070,N_3743,N_3541);
or U5071 (N_5071,N_4308,N_3827);
nand U5072 (N_5072,N_4655,N_4138);
nand U5073 (N_5073,N_2624,N_2959);
nor U5074 (N_5074,N_3220,N_3492);
or U5075 (N_5075,N_2922,N_4554);
xnor U5076 (N_5076,N_4796,N_3199);
and U5077 (N_5077,N_4459,N_2708);
nand U5078 (N_5078,N_4994,N_4435);
nand U5079 (N_5079,N_3727,N_3511);
nand U5080 (N_5080,N_4372,N_3932);
and U5081 (N_5081,N_3101,N_4099);
and U5082 (N_5082,N_4266,N_2789);
nand U5083 (N_5083,N_3112,N_3019);
nand U5084 (N_5084,N_2697,N_3969);
nor U5085 (N_5085,N_3899,N_3059);
and U5086 (N_5086,N_3693,N_2946);
and U5087 (N_5087,N_3673,N_4256);
and U5088 (N_5088,N_4539,N_2586);
nand U5089 (N_5089,N_4569,N_4367);
nand U5090 (N_5090,N_3214,N_3350);
xor U5091 (N_5091,N_2730,N_3774);
nor U5092 (N_5092,N_2980,N_4184);
and U5093 (N_5093,N_2629,N_4305);
or U5094 (N_5094,N_4223,N_4825);
nand U5095 (N_5095,N_2958,N_2972);
nor U5096 (N_5096,N_3304,N_4734);
and U5097 (N_5097,N_3232,N_3922);
nor U5098 (N_5098,N_2782,N_3733);
nor U5099 (N_5099,N_4814,N_3325);
and U5100 (N_5100,N_2863,N_3439);
nor U5101 (N_5101,N_2851,N_4314);
nor U5102 (N_5102,N_4897,N_4485);
nand U5103 (N_5103,N_4751,N_4878);
or U5104 (N_5104,N_4310,N_2542);
nand U5105 (N_5105,N_4070,N_2585);
xor U5106 (N_5106,N_4034,N_2630);
and U5107 (N_5107,N_3221,N_4377);
nand U5108 (N_5108,N_4306,N_4783);
nor U5109 (N_5109,N_3547,N_3528);
or U5110 (N_5110,N_3510,N_3334);
or U5111 (N_5111,N_3607,N_3702);
or U5112 (N_5112,N_4887,N_2574);
nor U5113 (N_5113,N_4548,N_2802);
or U5114 (N_5114,N_2669,N_3451);
nor U5115 (N_5115,N_2811,N_3044);
nand U5116 (N_5116,N_4667,N_3556);
nor U5117 (N_5117,N_4619,N_2957);
and U5118 (N_5118,N_4492,N_4750);
or U5119 (N_5119,N_3950,N_2567);
nand U5120 (N_5120,N_3858,N_4028);
nand U5121 (N_5121,N_2850,N_3473);
nor U5122 (N_5122,N_4262,N_4513);
nor U5123 (N_5123,N_3616,N_2930);
and U5124 (N_5124,N_4986,N_2776);
nand U5125 (N_5125,N_3082,N_2869);
nor U5126 (N_5126,N_3176,N_4519);
and U5127 (N_5127,N_3364,N_2838);
or U5128 (N_5128,N_3088,N_4536);
and U5129 (N_5129,N_2901,N_4185);
or U5130 (N_5130,N_2520,N_3955);
nor U5131 (N_5131,N_3282,N_3687);
and U5132 (N_5132,N_3952,N_3833);
or U5133 (N_5133,N_4043,N_4907);
nand U5134 (N_5134,N_3946,N_2834);
nor U5135 (N_5135,N_2954,N_4944);
or U5136 (N_5136,N_4534,N_3070);
or U5137 (N_5137,N_4488,N_4959);
nor U5138 (N_5138,N_3107,N_3467);
or U5139 (N_5139,N_2897,N_2594);
and U5140 (N_5140,N_3734,N_4095);
nor U5141 (N_5141,N_3713,N_3182);
nor U5142 (N_5142,N_2943,N_4447);
and U5143 (N_5143,N_3449,N_3939);
nor U5144 (N_5144,N_4711,N_2650);
or U5145 (N_5145,N_4683,N_4061);
or U5146 (N_5146,N_3096,N_3542);
and U5147 (N_5147,N_3330,N_3412);
nor U5148 (N_5148,N_4158,N_4368);
and U5149 (N_5149,N_4469,N_3049);
nand U5150 (N_5150,N_4466,N_4411);
nor U5151 (N_5151,N_3543,N_4420);
xor U5152 (N_5152,N_2704,N_3135);
and U5153 (N_5153,N_2910,N_2949);
nand U5154 (N_5154,N_3396,N_4213);
or U5155 (N_5155,N_2995,N_2735);
and U5156 (N_5156,N_2970,N_3416);
nand U5157 (N_5157,N_4486,N_4437);
and U5158 (N_5158,N_3537,N_2637);
nor U5159 (N_5159,N_3047,N_3573);
and U5160 (N_5160,N_4508,N_4614);
or U5161 (N_5161,N_3434,N_4623);
nor U5162 (N_5162,N_3295,N_3257);
nand U5163 (N_5163,N_3636,N_4850);
or U5164 (N_5164,N_4295,N_4200);
xor U5165 (N_5165,N_2795,N_4894);
and U5166 (N_5166,N_3753,N_2587);
xnor U5167 (N_5167,N_4951,N_3443);
nand U5168 (N_5168,N_3111,N_4765);
or U5169 (N_5169,N_4626,N_3427);
nor U5170 (N_5170,N_4271,N_3912);
nand U5171 (N_5171,N_3776,N_2645);
or U5172 (N_5172,N_4936,N_2500);
and U5173 (N_5173,N_4102,N_2746);
or U5174 (N_5174,N_4518,N_4343);
nor U5175 (N_5175,N_4439,N_4646);
and U5176 (N_5176,N_4870,N_4145);
nand U5177 (N_5177,N_3736,N_4071);
nand U5178 (N_5178,N_4514,N_4909);
or U5179 (N_5179,N_4713,N_4144);
and U5180 (N_5180,N_4076,N_3966);
nor U5181 (N_5181,N_3506,N_2998);
and U5182 (N_5182,N_3784,N_3535);
or U5183 (N_5183,N_2976,N_4352);
and U5184 (N_5184,N_3577,N_4527);
and U5185 (N_5185,N_4772,N_4379);
nor U5186 (N_5186,N_2990,N_3352);
nand U5187 (N_5187,N_4999,N_4895);
and U5188 (N_5188,N_2981,N_4980);
and U5189 (N_5189,N_4078,N_4584);
or U5190 (N_5190,N_3701,N_3889);
nand U5191 (N_5191,N_4596,N_3493);
and U5192 (N_5192,N_3896,N_4925);
nor U5193 (N_5193,N_3575,N_4560);
and U5194 (N_5194,N_4296,N_4784);
xnor U5195 (N_5195,N_3672,N_4981);
or U5196 (N_5196,N_2517,N_2874);
nand U5197 (N_5197,N_4874,N_3495);
xnor U5198 (N_5198,N_2979,N_3208);
or U5199 (N_5199,N_3920,N_2736);
or U5200 (N_5200,N_2670,N_4042);
nand U5201 (N_5201,N_3748,N_3227);
or U5202 (N_5202,N_3591,N_3924);
nand U5203 (N_5203,N_3063,N_3134);
nor U5204 (N_5204,N_4919,N_3081);
nand U5205 (N_5205,N_3140,N_3440);
or U5206 (N_5206,N_2690,N_3598);
or U5207 (N_5207,N_4632,N_3414);
nand U5208 (N_5208,N_3371,N_2506);
and U5209 (N_5209,N_4705,N_3989);
nand U5210 (N_5210,N_3552,N_3383);
or U5211 (N_5211,N_3228,N_4882);
or U5212 (N_5212,N_4605,N_4961);
xor U5213 (N_5213,N_3750,N_4495);
nand U5214 (N_5214,N_3275,N_3035);
nand U5215 (N_5215,N_3793,N_3961);
nand U5216 (N_5216,N_3368,N_2927);
nand U5217 (N_5217,N_4915,N_2806);
and U5218 (N_5218,N_2884,N_2989);
nand U5219 (N_5219,N_4617,N_3645);
nor U5220 (N_5220,N_2625,N_3116);
or U5221 (N_5221,N_3274,N_4048);
nand U5222 (N_5222,N_3630,N_4511);
and U5223 (N_5223,N_2988,N_4701);
nor U5224 (N_5224,N_3557,N_4501);
nand U5225 (N_5225,N_3909,N_4162);
and U5226 (N_5226,N_4253,N_3177);
nor U5227 (N_5227,N_2837,N_4363);
xor U5228 (N_5228,N_4000,N_3464);
or U5229 (N_5229,N_4163,N_2682);
nor U5230 (N_5230,N_3960,N_4197);
nand U5231 (N_5231,N_4572,N_4177);
xnor U5232 (N_5232,N_4094,N_3650);
and U5233 (N_5233,N_3163,N_2524);
nor U5234 (N_5234,N_4516,N_3231);
or U5235 (N_5235,N_4446,N_4015);
nand U5236 (N_5236,N_4824,N_3582);
and U5237 (N_5237,N_3999,N_2633);
nand U5238 (N_5238,N_3518,N_3531);
nor U5239 (N_5239,N_2825,N_3457);
nor U5240 (N_5240,N_3903,N_4888);
and U5241 (N_5241,N_3197,N_3525);
and U5242 (N_5242,N_2687,N_4746);
and U5243 (N_5243,N_4732,N_3040);
nand U5244 (N_5244,N_3115,N_3192);
nor U5245 (N_5245,N_3706,N_3677);
nand U5246 (N_5246,N_3501,N_3052);
nor U5247 (N_5247,N_3174,N_4641);
nor U5248 (N_5248,N_4126,N_4773);
nand U5249 (N_5249,N_4053,N_4578);
and U5250 (N_5250,N_4631,N_3797);
nor U5251 (N_5251,N_2808,N_3033);
or U5252 (N_5252,N_4050,N_4012);
and U5253 (N_5253,N_3988,N_3652);
or U5254 (N_5254,N_4137,N_4427);
nand U5255 (N_5255,N_3809,N_3128);
nor U5256 (N_5256,N_3251,N_3193);
nand U5257 (N_5257,N_4165,N_2747);
or U5258 (N_5258,N_3211,N_3832);
nor U5259 (N_5259,N_3149,N_4913);
nor U5260 (N_5260,N_3122,N_4789);
or U5261 (N_5261,N_4400,N_3009);
and U5262 (N_5262,N_4376,N_3083);
nor U5263 (N_5263,N_2929,N_3884);
or U5264 (N_5264,N_3803,N_4933);
and U5265 (N_5265,N_2842,N_3159);
and U5266 (N_5266,N_4830,N_3164);
and U5267 (N_5267,N_3317,N_3914);
nor U5268 (N_5268,N_3499,N_3497);
nand U5269 (N_5269,N_4726,N_4669);
nand U5270 (N_5270,N_3018,N_3567);
nor U5271 (N_5271,N_3469,N_3016);
and U5272 (N_5272,N_4467,N_4628);
nand U5273 (N_5273,N_4496,N_3055);
nor U5274 (N_5274,N_3735,N_4249);
nor U5275 (N_5275,N_2859,N_4299);
or U5276 (N_5276,N_4033,N_3109);
or U5277 (N_5277,N_3345,N_2676);
and U5278 (N_5278,N_3789,N_4790);
and U5279 (N_5279,N_3977,N_4976);
nand U5280 (N_5280,N_3572,N_3357);
or U5281 (N_5281,N_4020,N_3060);
and U5282 (N_5282,N_4421,N_3054);
and U5283 (N_5283,N_4991,N_3813);
xor U5284 (N_5284,N_3937,N_2857);
nor U5285 (N_5285,N_4026,N_4106);
nor U5286 (N_5286,N_3471,N_3998);
nor U5287 (N_5287,N_2793,N_2840);
or U5288 (N_5288,N_3669,N_3252);
nor U5289 (N_5289,N_3235,N_3381);
or U5290 (N_5290,N_4120,N_4063);
and U5291 (N_5291,N_4901,N_3351);
and U5292 (N_5292,N_3385,N_3610);
nand U5293 (N_5293,N_4448,N_3764);
or U5294 (N_5294,N_2550,N_3113);
and U5295 (N_5295,N_2644,N_3944);
xor U5296 (N_5296,N_2999,N_2692);
nor U5297 (N_5297,N_3302,N_4722);
xor U5298 (N_5298,N_4590,N_3025);
nand U5299 (N_5299,N_4442,N_4872);
nand U5300 (N_5300,N_3462,N_3993);
nand U5301 (N_5301,N_4807,N_3382);
nand U5302 (N_5302,N_4634,N_4649);
and U5303 (N_5303,N_3114,N_3514);
nor U5304 (N_5304,N_4273,N_3039);
nand U5305 (N_5305,N_3415,N_4417);
xor U5306 (N_5306,N_2525,N_3604);
or U5307 (N_5307,N_4652,N_4615);
or U5308 (N_5308,N_3714,N_4221);
nor U5309 (N_5309,N_3625,N_4426);
nor U5310 (N_5310,N_2571,N_3498);
or U5311 (N_5311,N_3237,N_4759);
or U5312 (N_5312,N_3517,N_3285);
and U5313 (N_5313,N_2655,N_4859);
and U5314 (N_5314,N_4087,N_4260);
and U5315 (N_5315,N_4118,N_2750);
nand U5316 (N_5316,N_3705,N_2778);
and U5317 (N_5317,N_4754,N_3386);
nand U5318 (N_5318,N_3484,N_4686);
nand U5319 (N_5319,N_2616,N_3031);
nand U5320 (N_5320,N_2621,N_4633);
nor U5321 (N_5321,N_3034,N_3883);
or U5322 (N_5322,N_3638,N_3500);
and U5323 (N_5323,N_4962,N_4431);
nand U5324 (N_5324,N_4588,N_2662);
and U5325 (N_5325,N_4414,N_3921);
nand U5326 (N_5326,N_3429,N_3586);
nand U5327 (N_5327,N_4207,N_3323);
nor U5328 (N_5328,N_4664,N_3576);
nor U5329 (N_5329,N_2797,N_3256);
xor U5330 (N_5330,N_4809,N_2660);
nand U5331 (N_5331,N_3646,N_3888);
or U5332 (N_5332,N_3779,N_2769);
or U5333 (N_5333,N_4777,N_2559);
and U5334 (N_5334,N_2852,N_2962);
nor U5335 (N_5335,N_2557,N_4027);
and U5336 (N_5336,N_3264,N_3348);
nor U5337 (N_5337,N_4149,N_3654);
or U5338 (N_5338,N_3621,N_4690);
nand U5339 (N_5339,N_2674,N_4418);
or U5340 (N_5340,N_4687,N_3503);
xor U5341 (N_5341,N_3804,N_4160);
or U5342 (N_5342,N_2533,N_4670);
xor U5343 (N_5343,N_4188,N_4550);
and U5344 (N_5344,N_3032,N_2836);
or U5345 (N_5345,N_3548,N_2545);
and U5346 (N_5346,N_2678,N_4503);
nor U5347 (N_5347,N_3085,N_3146);
nor U5348 (N_5348,N_2547,N_4111);
nor U5349 (N_5349,N_3578,N_4350);
or U5350 (N_5350,N_4723,N_4461);
and U5351 (N_5351,N_2753,N_3679);
nor U5352 (N_5352,N_2732,N_3084);
and U5353 (N_5353,N_3767,N_3204);
nor U5354 (N_5354,N_3360,N_4549);
or U5355 (N_5355,N_4598,N_3147);
and U5356 (N_5356,N_3555,N_3108);
nor U5357 (N_5357,N_3068,N_4134);
nand U5358 (N_5358,N_3949,N_2514);
nor U5359 (N_5359,N_4178,N_4761);
or U5360 (N_5360,N_3954,N_4183);
nand U5361 (N_5361,N_3992,N_4164);
nand U5362 (N_5362,N_4468,N_2824);
and U5363 (N_5363,N_4731,N_3963);
nor U5364 (N_5364,N_2512,N_3876);
nand U5365 (N_5365,N_3665,N_3717);
or U5366 (N_5366,N_3117,N_2986);
and U5367 (N_5367,N_4562,N_3709);
and U5368 (N_5368,N_3869,N_2673);
nand U5369 (N_5369,N_2813,N_4862);
nand U5370 (N_5370,N_4240,N_3599);
and U5371 (N_5371,N_2578,N_4405);
xor U5372 (N_5372,N_4861,N_3418);
and U5373 (N_5373,N_4084,N_4808);
and U5374 (N_5374,N_4869,N_3801);
nand U5375 (N_5375,N_2991,N_3234);
nand U5376 (N_5376,N_3491,N_2864);
and U5377 (N_5377,N_3268,N_2641);
nand U5378 (N_5378,N_3162,N_4934);
nand U5379 (N_5379,N_3315,N_3847);
and U5380 (N_5380,N_3751,N_3442);
or U5381 (N_5381,N_3249,N_4279);
or U5382 (N_5382,N_4276,N_3612);
nand U5383 (N_5383,N_2880,N_2893);
nor U5384 (N_5384,N_3682,N_3516);
and U5385 (N_5385,N_3137,N_3593);
nor U5386 (N_5386,N_3786,N_4409);
and U5387 (N_5387,N_4386,N_4583);
and U5388 (N_5388,N_3644,N_4770);
xnor U5389 (N_5389,N_4037,N_4747);
nand U5390 (N_5390,N_3868,N_4136);
xor U5391 (N_5391,N_3704,N_3823);
nor U5392 (N_5392,N_4799,N_2565);
or U5393 (N_5393,N_4170,N_4119);
nand U5394 (N_5394,N_3563,N_3073);
nor U5395 (N_5395,N_2858,N_2713);
and U5396 (N_5396,N_3037,N_3399);
nor U5397 (N_5397,N_4877,N_3581);
and U5398 (N_5398,N_3169,N_2961);
nor U5399 (N_5399,N_3742,N_2612);
nand U5400 (N_5400,N_3316,N_4716);
nand U5401 (N_5401,N_4062,N_2888);
nor U5402 (N_5402,N_3930,N_3843);
and U5403 (N_5403,N_3015,N_3728);
xnor U5404 (N_5404,N_4788,N_3271);
or U5405 (N_5405,N_4660,N_4428);
and U5406 (N_5406,N_3716,N_4471);
nand U5407 (N_5407,N_2590,N_3119);
nor U5408 (N_5408,N_4312,N_4199);
and U5409 (N_5409,N_2919,N_4408);
nand U5410 (N_5410,N_4413,N_4280);
nor U5411 (N_5411,N_4009,N_3446);
and U5412 (N_5412,N_3648,N_3508);
or U5413 (N_5413,N_4357,N_3389);
nand U5414 (N_5414,N_4778,N_4242);
xor U5415 (N_5415,N_4721,N_3405);
nand U5416 (N_5416,N_3747,N_4284);
and U5417 (N_5417,N_2982,N_3800);
nor U5418 (N_5418,N_3408,N_3799);
nand U5419 (N_5419,N_3296,N_3720);
nor U5420 (N_5420,N_2556,N_2656);
nor U5421 (N_5421,N_4843,N_4208);
nand U5422 (N_5422,N_2861,N_4334);
xor U5423 (N_5423,N_4604,N_4960);
or U5424 (N_5424,N_3975,N_2766);
nor U5425 (N_5425,N_3674,N_4231);
and U5426 (N_5426,N_3562,N_3666);
nand U5427 (N_5427,N_3229,N_3318);
nand U5428 (N_5428,N_4975,N_3908);
or U5429 (N_5429,N_3127,N_4107);
nor U5430 (N_5430,N_3928,N_3723);
nor U5431 (N_5431,N_2576,N_3731);
nor U5432 (N_5432,N_4159,N_3816);
and U5433 (N_5433,N_3038,N_3260);
and U5434 (N_5434,N_4873,N_4719);
nand U5435 (N_5435,N_3387,N_4358);
xnor U5436 (N_5436,N_4024,N_2560);
and U5437 (N_5437,N_2604,N_3339);
nor U5438 (N_5438,N_2741,N_4854);
or U5439 (N_5439,N_4553,N_4820);
and U5440 (N_5440,N_4003,N_4456);
and U5441 (N_5441,N_2665,N_3322);
nor U5442 (N_5442,N_3465,N_3363);
nor U5443 (N_5443,N_3239,N_3631);
nor U5444 (N_5444,N_3298,N_4304);
and U5445 (N_5445,N_3306,N_2770);
nor U5446 (N_5446,N_3375,N_3796);
nor U5447 (N_5447,N_2755,N_4031);
and U5448 (N_5448,N_3253,N_2964);
and U5449 (N_5449,N_4504,N_4568);
nand U5450 (N_5450,N_4051,N_3172);
and U5451 (N_5451,N_4717,N_4982);
nand U5452 (N_5452,N_3973,N_4910);
nor U5453 (N_5453,N_4858,N_4211);
nor U5454 (N_5454,N_3588,N_3423);
nand U5455 (N_5455,N_3945,N_4823);
or U5456 (N_5456,N_4900,N_3965);
nor U5457 (N_5457,N_4586,N_3017);
or U5458 (N_5458,N_2743,N_4210);
nand U5459 (N_5459,N_3771,N_4301);
and U5460 (N_5460,N_2829,N_4041);
and U5461 (N_5461,N_3267,N_4059);
and U5462 (N_5462,N_4080,N_4908);
and U5463 (N_5463,N_4114,N_2688);
nand U5464 (N_5464,N_2553,N_4730);
nor U5465 (N_5465,N_4142,N_2715);
nor U5466 (N_5466,N_3324,N_4478);
nand U5467 (N_5467,N_4643,N_3845);
and U5468 (N_5468,N_3028,N_3822);
xor U5469 (N_5469,N_3165,N_4244);
and U5470 (N_5470,N_3029,N_3836);
or U5471 (N_5471,N_4708,N_4073);
xnor U5472 (N_5472,N_3240,N_3042);
and U5473 (N_5473,N_3948,N_4038);
and U5474 (N_5474,N_3692,N_4075);
xor U5475 (N_5475,N_4112,N_2546);
nand U5476 (N_5476,N_3048,N_4684);
nor U5477 (N_5477,N_4443,N_4499);
nand U5478 (N_5478,N_3459,N_4606);
nand U5479 (N_5479,N_4794,N_2728);
nor U5480 (N_5480,N_4689,N_4556);
xor U5481 (N_5481,N_4505,N_4840);
or U5482 (N_5482,N_2686,N_3600);
or U5483 (N_5483,N_4868,N_3168);
and U5484 (N_5484,N_3320,N_3454);
nand U5485 (N_5485,N_3606,N_3321);
nor U5486 (N_5486,N_2771,N_3906);
or U5487 (N_5487,N_2504,N_3815);
or U5488 (N_5488,N_4969,N_4462);
nand U5489 (N_5489,N_3587,N_2904);
and U5490 (N_5490,N_4939,N_3941);
nand U5491 (N_5491,N_3023,N_3241);
xor U5492 (N_5492,N_4179,N_4092);
or U5493 (N_5493,N_2611,N_2785);
and U5494 (N_5494,N_4011,N_2675);
nor U5495 (N_5495,N_4815,N_3513);
nand U5496 (N_5496,N_4693,N_2572);
nand U5497 (N_5497,N_4666,N_4531);
or U5498 (N_5498,N_2994,N_4916);
and U5499 (N_5499,N_4612,N_3148);
and U5500 (N_5500,N_4581,N_2575);
or U5501 (N_5501,N_3925,N_4128);
nand U5502 (N_5502,N_3435,N_4407);
xor U5503 (N_5503,N_3722,N_3183);
nor U5504 (N_5504,N_4831,N_4169);
or U5505 (N_5505,N_4920,N_4851);
xnor U5506 (N_5506,N_3444,N_4673);
and U5507 (N_5507,N_3329,N_4662);
or U5508 (N_5508,N_3838,N_2835);
nand U5509 (N_5509,N_3917,N_3574);
xnor U5510 (N_5510,N_4148,N_2921);
and U5511 (N_5511,N_3002,N_4587);
nor U5512 (N_5512,N_3181,N_3719);
and U5513 (N_5513,N_3634,N_4545);
nand U5514 (N_5514,N_4040,N_4728);
nor U5515 (N_5515,N_4839,N_3765);
or U5516 (N_5516,N_2937,N_4294);
xnor U5517 (N_5517,N_3700,N_3098);
and U5518 (N_5518,N_3075,N_4132);
and U5519 (N_5519,N_3281,N_4838);
nand U5520 (N_5520,N_4391,N_4425);
nor U5521 (N_5521,N_3818,N_3737);
xnor U5522 (N_5522,N_4927,N_4445);
nand U5523 (N_5523,N_3972,N_4573);
nor U5524 (N_5524,N_3795,N_4847);
nand U5525 (N_5525,N_4767,N_4786);
and U5526 (N_5526,N_3526,N_2502);
nor U5527 (N_5527,N_2622,N_3293);
or U5528 (N_5528,N_3987,N_3835);
and U5529 (N_5529,N_4865,N_4006);
and U5530 (N_5530,N_4577,N_4718);
nand U5531 (N_5531,N_4918,N_2589);
nand U5532 (N_5532,N_3470,N_3378);
xnor U5533 (N_5533,N_3900,N_4852);
nand U5534 (N_5534,N_4826,N_4845);
or U5535 (N_5535,N_4194,N_4551);
nor U5536 (N_5536,N_3139,N_3236);
nor U5537 (N_5537,N_4187,N_4766);
and U5538 (N_5538,N_3194,N_3178);
nor U5539 (N_5539,N_4970,N_3065);
xor U5540 (N_5540,N_3030,N_3066);
and U5541 (N_5541,N_4949,N_3894);
or U5542 (N_5542,N_4481,N_4659);
nand U5543 (N_5543,N_4025,N_3061);
nor U5544 (N_5544,N_4237,N_2558);
and U5545 (N_5545,N_4963,N_3212);
or U5546 (N_5546,N_3213,N_4189);
or U5547 (N_5547,N_2950,N_4593);
nand U5548 (N_5548,N_4833,N_4879);
nand U5549 (N_5549,N_4171,N_3620);
xor U5550 (N_5550,N_3676,N_3614);
xor U5551 (N_5551,N_3136,N_2539);
and U5552 (N_5552,N_4054,N_3003);
nand U5553 (N_5553,N_4608,N_3133);
and U5554 (N_5554,N_4699,N_4768);
and U5555 (N_5555,N_4860,N_3310);
nand U5556 (N_5556,N_3554,N_2623);
nor U5557 (N_5557,N_3071,N_4441);
nor U5558 (N_5558,N_2647,N_2780);
nand U5559 (N_5559,N_4457,N_3072);
or U5560 (N_5560,N_4181,N_4509);
or U5561 (N_5561,N_4526,N_4228);
and U5562 (N_5562,N_4086,N_3461);
and U5563 (N_5563,N_3226,N_4594);
nand U5564 (N_5564,N_3284,N_4676);
and U5565 (N_5565,N_2847,N_3486);
or U5566 (N_5566,N_4017,N_3406);
nor U5567 (N_5567,N_4036,N_2631);
xor U5568 (N_5568,N_2740,N_4880);
and U5569 (N_5569,N_2707,N_4668);
nor U5570 (N_5570,N_4234,N_3417);
nor U5571 (N_5571,N_2827,N_3863);
and U5572 (N_5572,N_2951,N_4849);
and U5573 (N_5573,N_4123,N_4898);
xnor U5574 (N_5574,N_3380,N_4798);
and U5575 (N_5575,N_3445,N_3807);
or U5576 (N_5576,N_3354,N_4155);
or U5577 (N_5577,N_2775,N_2552);
and U5578 (N_5578,N_4288,N_4089);
and U5579 (N_5579,N_3840,N_4763);
and U5580 (N_5580,N_3118,N_4044);
nand U5581 (N_5581,N_4281,N_3205);
nor U5582 (N_5582,N_4656,N_2702);
and U5583 (N_5583,N_2549,N_4502);
and U5584 (N_5584,N_3855,N_4948);
nand U5585 (N_5585,N_4758,N_4507);
xor U5586 (N_5586,N_4016,N_4135);
and U5587 (N_5587,N_2978,N_4375);
nor U5588 (N_5588,N_4567,N_2648);
nor U5589 (N_5589,N_3247,N_3632);
xor U5590 (N_5590,N_2737,N_3841);
nor U5591 (N_5591,N_4173,N_3886);
and U5592 (N_5592,N_4337,N_3216);
nand U5593 (N_5593,N_4855,N_3757);
nand U5594 (N_5594,N_2531,N_3647);
nor U5595 (N_5595,N_3655,N_3132);
nand U5596 (N_5596,N_3261,N_2942);
or U5597 (N_5597,N_3481,N_2873);
and U5598 (N_5598,N_3530,N_4315);
xor U5599 (N_5599,N_2807,N_4806);
or U5600 (N_5600,N_2610,N_2725);
nor U5601 (N_5601,N_4388,N_4222);
and U5602 (N_5602,N_3421,N_4320);
and U5603 (N_5603,N_2860,N_3011);
xor U5604 (N_5604,N_2953,N_3689);
xnor U5605 (N_5605,N_4997,N_3681);
or U5606 (N_5606,N_4639,N_3254);
and U5607 (N_5607,N_3512,N_4046);
or U5608 (N_5608,N_3422,N_2534);
and U5609 (N_5609,N_4470,N_3639);
nor U5610 (N_5610,N_2619,N_4045);
nor U5611 (N_5611,N_4167,N_4129);
nor U5612 (N_5612,N_3358,N_3710);
xnor U5613 (N_5613,N_4369,N_3891);
and U5614 (N_5614,N_3198,N_3091);
nor U5615 (N_5615,N_4422,N_3311);
nand U5616 (N_5616,N_3327,N_3775);
nor U5617 (N_5617,N_4647,N_4270);
or U5618 (N_5618,N_4953,N_3426);
or U5619 (N_5619,N_4525,N_4965);
nand U5620 (N_5620,N_2607,N_3595);
or U5621 (N_5621,N_4100,N_4465);
nand U5622 (N_5622,N_4735,N_4109);
or U5623 (N_5623,N_3309,N_4316);
and U5624 (N_5624,N_3255,N_4964);
nor U5625 (N_5625,N_3294,N_3288);
and U5626 (N_5626,N_3430,N_2716);
and U5627 (N_5627,N_3359,N_2635);
xor U5628 (N_5628,N_3394,N_2871);
or U5629 (N_5629,N_2701,N_3043);
and U5630 (N_5630,N_2868,N_4832);
and U5631 (N_5631,N_2761,N_4483);
nand U5632 (N_5632,N_3478,N_3507);
nor U5633 (N_5633,N_3455,N_4559);
nand U5634 (N_5634,N_3892,N_4333);
and U5635 (N_5635,N_3596,N_2664);
nand U5636 (N_5636,N_3926,N_2788);
nor U5637 (N_5637,N_2505,N_2581);
and U5638 (N_5638,N_3523,N_4592);
or U5639 (N_5639,N_4450,N_4335);
or U5640 (N_5640,N_3597,N_4353);
or U5641 (N_5641,N_3515,N_2721);
and U5642 (N_5642,N_2548,N_4336);
nand U5643 (N_5643,N_3207,N_3703);
nor U5644 (N_5644,N_2720,N_2518);
or U5645 (N_5645,N_3258,N_4403);
nor U5646 (N_5646,N_4905,N_4704);
or U5647 (N_5647,N_4698,N_3663);
nand U5648 (N_5648,N_4039,N_4654);
nor U5649 (N_5649,N_4241,N_4813);
nor U5650 (N_5650,N_4444,N_3724);
nor U5651 (N_5651,N_2924,N_4709);
and U5652 (N_5652,N_3697,N_4700);
xnor U5653 (N_5653,N_4300,N_4298);
and U5654 (N_5654,N_3291,N_4725);
or U5655 (N_5655,N_2822,N_4834);
nor U5656 (N_5656,N_2522,N_3970);
xnor U5657 (N_5657,N_2620,N_4057);
and U5658 (N_5658,N_3121,N_2738);
and U5659 (N_5659,N_4220,N_3171);
or U5660 (N_5660,N_3398,N_4844);
and U5661 (N_5661,N_4110,N_3538);
xor U5662 (N_5662,N_2787,N_4979);
or U5663 (N_5663,N_3913,N_3244);
and U5664 (N_5664,N_4010,N_4248);
or U5665 (N_5665,N_2739,N_2544);
nor U5666 (N_5666,N_3678,N_4812);
or U5667 (N_5667,N_3262,N_4219);
xnor U5668 (N_5668,N_3740,N_3328);
nor U5669 (N_5669,N_4835,N_2628);
and U5670 (N_5670,N_4928,N_4769);
and U5671 (N_5671,N_3287,N_2870);
nand U5672 (N_5672,N_3837,N_4941);
nand U5673 (N_5673,N_3027,N_3300);
and U5674 (N_5674,N_3014,N_4487);
and U5675 (N_5675,N_3810,N_4484);
or U5676 (N_5676,N_4520,N_4589);
and U5677 (N_5677,N_2767,N_4214);
nand U5678 (N_5678,N_3413,N_3079);
xor U5679 (N_5679,N_3670,N_4974);
and U5680 (N_5680,N_3520,N_3245);
or U5681 (N_5681,N_2573,N_4795);
and U5682 (N_5682,N_4190,N_4117);
or U5683 (N_5683,N_4049,N_2603);
nand U5684 (N_5684,N_4884,N_4597);
nand U5685 (N_5685,N_2535,N_3867);
nor U5686 (N_5686,N_4365,N_3895);
nor U5687 (N_5687,N_3319,N_2685);
nand U5688 (N_5688,N_4348,N_4098);
nor U5689 (N_5689,N_3209,N_3448);
and U5690 (N_5690,N_2914,N_2841);
nand U5691 (N_5691,N_2805,N_2672);
and U5692 (N_5692,N_2826,N_3715);
xor U5693 (N_5693,N_3062,N_4332);
and U5694 (N_5694,N_2933,N_4474);
or U5695 (N_5695,N_2538,N_2968);
xnor U5696 (N_5696,N_3619,N_4064);
nor U5697 (N_5697,N_4115,N_3860);
and U5698 (N_5698,N_3792,N_2799);
xor U5699 (N_5699,N_4966,N_2510);
nand U5700 (N_5700,N_2781,N_3957);
or U5701 (N_5701,N_4264,N_2666);
nor U5702 (N_5702,N_4945,N_4729);
nand U5703 (N_5703,N_3013,N_4007);
nand U5704 (N_5704,N_4703,N_4139);
nor U5705 (N_5705,N_4775,N_3404);
and U5706 (N_5706,N_4906,N_4331);
nor U5707 (N_5707,N_4585,N_4451);
nor U5708 (N_5708,N_3686,N_4621);
nor U5709 (N_5709,N_3080,N_2671);
xnor U5710 (N_5710,N_3151,N_2653);
nor U5711 (N_5711,N_3374,N_4745);
and U5712 (N_5712,N_2583,N_3012);
nor U5713 (N_5713,N_4946,N_4374);
and U5714 (N_5714,N_3424,N_4821);
nand U5715 (N_5715,N_2947,N_3877);
nand U5716 (N_5716,N_2609,N_3489);
and U5717 (N_5717,N_3721,N_2917);
xor U5718 (N_5718,N_4515,N_3391);
or U5719 (N_5719,N_3708,N_4360);
xor U5720 (N_5720,N_4896,N_3811);
nor U5721 (N_5721,N_4390,N_4463);
and U5722 (N_5722,N_3377,N_2727);
nand U5723 (N_5723,N_2928,N_4021);
nand U5724 (N_5724,N_2744,N_2934);
or U5725 (N_5725,N_3006,N_4954);
nand U5726 (N_5726,N_4303,N_4972);
nand U5727 (N_5727,N_3482,N_3297);
and U5728 (N_5728,N_3688,N_4085);
nand U5729 (N_5729,N_4347,N_2896);
nand U5730 (N_5730,N_4005,N_2882);
or U5731 (N_5731,N_4072,N_4113);
and U5732 (N_5732,N_2639,N_3100);
nand U5733 (N_5733,N_3527,N_4319);
nor U5734 (N_5734,N_2812,N_4362);
nand U5735 (N_5735,N_3104,N_3881);
or U5736 (N_5736,N_2689,N_3898);
nor U5737 (N_5737,N_4014,N_4423);
and U5738 (N_5738,N_2663,N_3982);
nand U5739 (N_5739,N_2820,N_2783);
nor U5740 (N_5740,N_4079,N_3680);
nand U5741 (N_5741,N_3277,N_3093);
nand U5742 (N_5742,N_4528,N_4983);
nand U5743 (N_5743,N_4856,N_4771);
and U5744 (N_5744,N_3918,N_4968);
or U5745 (N_5745,N_3533,N_3524);
nand U5746 (N_5746,N_4875,N_4429);
nor U5747 (N_5747,N_4566,N_3794);
nor U5748 (N_5748,N_4671,N_4533);
and U5749 (N_5749,N_2733,N_4827);
nor U5750 (N_5750,N_4622,N_2915);
or U5751 (N_5751,N_2528,N_2537);
nand U5752 (N_5752,N_4090,N_3560);
nor U5753 (N_5753,N_2582,N_4455);
or U5754 (N_5754,N_3384,N_4245);
xnor U5755 (N_5755,N_4436,N_3760);
nor U5756 (N_5756,N_3290,N_3990);
nor U5757 (N_5757,N_2554,N_4804);
or U5758 (N_5758,N_3656,N_3366);
nor U5759 (N_5759,N_4077,N_3090);
and U5760 (N_5760,N_3626,N_4613);
nand U5761 (N_5761,N_2668,N_3420);
or U5762 (N_5762,N_4154,N_4318);
or U5763 (N_5763,N_4791,N_3788);
nand U5764 (N_5764,N_3566,N_3026);
nand U5765 (N_5765,N_3230,N_4477);
and U5766 (N_5766,N_3808,N_4216);
nand U5767 (N_5767,N_3125,N_3905);
and U5768 (N_5768,N_2891,N_4564);
or U5769 (N_5769,N_3202,N_2798);
and U5770 (N_5770,N_4140,N_3210);
nor U5771 (N_5771,N_3505,N_4512);
nand U5772 (N_5772,N_3830,N_4204);
or U5773 (N_5773,N_3152,N_4889);
and U5774 (N_5774,N_2815,N_3007);
nor U5775 (N_5775,N_2714,N_2532);
and U5776 (N_5776,N_4416,N_4665);
and U5777 (N_5777,N_3087,N_3544);
nand U5778 (N_5778,N_2764,N_4225);
nor U5779 (N_5779,N_4935,N_4212);
nor U5780 (N_5780,N_2925,N_3866);
xnor U5781 (N_5781,N_3155,N_3873);
or U5782 (N_5782,N_3187,N_2636);
and U5783 (N_5783,N_4971,N_3684);
nand U5784 (N_5784,N_4218,N_3092);
nand U5785 (N_5785,N_4618,N_3649);
or U5786 (N_5786,N_3570,N_2569);
nor U5787 (N_5787,N_3141,N_4476);
xor U5788 (N_5788,N_4702,N_2541);
nand U5789 (N_5789,N_3074,N_3008);
or U5790 (N_5790,N_4326,N_4696);
nand U5791 (N_5791,N_4292,N_3479);
and U5792 (N_5792,N_4022,N_3766);
nor U5793 (N_5793,N_4217,N_4793);
nand U5794 (N_5794,N_4779,N_2810);
nor U5795 (N_5795,N_3671,N_3303);
or U5796 (N_5796,N_3401,N_3968);
nand U5797 (N_5797,N_4706,N_3480);
nor U5798 (N_5798,N_4510,N_3200);
and U5799 (N_5799,N_2971,N_3331);
and U5800 (N_5800,N_4694,N_2667);
nand U5801 (N_5801,N_3106,N_4371);
or U5802 (N_5802,N_3996,N_3814);
nand U5803 (N_5803,N_4762,N_3057);
and U5804 (N_5804,N_2566,N_4764);
nor U5805 (N_5805,N_4246,N_4848);
and U5806 (N_5806,N_4893,N_2710);
nand U5807 (N_5807,N_4272,N_3219);
nor U5808 (N_5808,N_3592,N_3675);
nor U5809 (N_5809,N_2907,N_3820);
and U5810 (N_5810,N_4464,N_2599);
nand U5811 (N_5811,N_4392,N_2855);
and U5812 (N_5812,N_4697,N_4269);
nand U5813 (N_5813,N_4921,N_3878);
and U5814 (N_5814,N_3553,N_4493);
nand U5815 (N_5815,N_2772,N_3642);
nand U5816 (N_5816,N_3768,N_4943);
nand U5817 (N_5817,N_3000,N_4876);
and U5818 (N_5818,N_2627,N_3456);
nand U5819 (N_5819,N_4410,N_3558);
nor U5820 (N_5820,N_3643,N_4892);
nand U5821 (N_5821,N_4382,N_4625);
and U5822 (N_5822,N_4235,N_4742);
nor U5823 (N_5823,N_4150,N_2777);
nand U5824 (N_5824,N_3402,N_3875);
or U5825 (N_5825,N_3690,N_3335);
xnor U5826 (N_5826,N_3238,N_4500);
nor U5827 (N_5827,N_3780,N_3901);
and U5828 (N_5828,N_3602,N_2703);
or U5829 (N_5829,N_3138,N_3259);
or U5830 (N_5830,N_4247,N_4952);
nand U5831 (N_5831,N_2696,N_3540);
or U5832 (N_5832,N_3856,N_4389);
and U5833 (N_5833,N_2819,N_4285);
or U5834 (N_5834,N_4942,N_4440);
nor U5835 (N_5835,N_4737,N_2913);
nand U5836 (N_5836,N_4555,N_3851);
and U5837 (N_5837,N_3971,N_3942);
nand U5838 (N_5838,N_3668,N_3487);
xnor U5839 (N_5839,N_3188,N_3828);
nor U5840 (N_5840,N_4330,N_3393);
or U5841 (N_5841,N_3826,N_4682);
and U5842 (N_5842,N_3831,N_4903);
xor U5843 (N_5843,N_2854,N_2680);
or U5844 (N_5844,N_3589,N_2694);
xor U5845 (N_5845,N_4175,N_3985);
nor U5846 (N_5846,N_2757,N_2508);
nor U5847 (N_5847,N_4066,N_3494);
nand U5848 (N_5848,N_2614,N_3667);
nand U5849 (N_5849,N_3885,N_3864);
xor U5850 (N_5850,N_3534,N_3077);
or U5851 (N_5851,N_3224,N_3951);
xnor U5852 (N_5852,N_3893,N_3991);
and U5853 (N_5853,N_2709,N_4215);
nand U5854 (N_5854,N_4890,N_2698);
nand U5855 (N_5855,N_3142,N_4653);
and U5856 (N_5856,N_4720,N_3854);
and U5857 (N_5857,N_3095,N_4359);
nor U5858 (N_5858,N_4756,N_3947);
nand U5859 (N_5859,N_4600,N_2967);
nand U5860 (N_5860,N_2711,N_3611);
and U5861 (N_5861,N_3313,N_2511);
or U5862 (N_5862,N_3824,N_2509);
or U5863 (N_5863,N_3967,N_4105);
or U5864 (N_5864,N_3392,N_3365);
and U5865 (N_5865,N_4541,N_4651);
nand U5866 (N_5866,N_3657,N_4810);
nand U5867 (N_5867,N_2503,N_2593);
and U5868 (N_5868,N_3729,N_4620);
nor U5869 (N_5869,N_3036,N_3150);
nor U5870 (N_5870,N_3103,N_2774);
and U5871 (N_5871,N_4950,N_3995);
xnor U5872 (N_5872,N_3725,N_3879);
and U5873 (N_5873,N_3021,N_3696);
and U5874 (N_5874,N_2866,N_3532);
or U5875 (N_5875,N_4302,N_4680);
nand U5876 (N_5876,N_2568,N_4283);
nand U5877 (N_5877,N_3974,N_2889);
xor U5878 (N_5878,N_3186,N_3301);
xnor U5879 (N_5879,N_2657,N_2993);
or U5880 (N_5880,N_3787,N_4582);
nor U5881 (N_5881,N_4640,N_3919);
nand U5882 (N_5882,N_3622,N_4535);
or U5883 (N_5883,N_4161,N_4561);
nand U5884 (N_5884,N_4097,N_3564);
and U5885 (N_5885,N_4557,N_3936);
or U5886 (N_5886,N_3842,N_4355);
nor U5887 (N_5887,N_2588,N_3160);
nand U5888 (N_5888,N_4282,N_4364);
nor U5889 (N_5889,N_4202,N_4402);
or U5890 (N_5890,N_2790,N_3185);
and U5891 (N_5891,N_2909,N_3355);
nand U5892 (N_5892,N_2844,N_3110);
and U5893 (N_5893,N_4864,N_3628);
nand U5894 (N_5894,N_4322,N_2879);
nor U5895 (N_5895,N_2584,N_3653);
or U5896 (N_5896,N_4001,N_3923);
and U5897 (N_5897,N_3156,N_4967);
nand U5898 (N_5898,N_4195,N_4837);
or U5899 (N_5899,N_3223,N_4317);
or U5900 (N_5900,N_4679,N_3661);
nor U5901 (N_5901,N_4650,N_4993);
and U5902 (N_5902,N_4924,N_3419);
and U5903 (N_5903,N_2955,N_2902);
or U5904 (N_5904,N_4542,N_2800);
or U5905 (N_5905,N_4801,N_4258);
nand U5906 (N_5906,N_2883,N_4692);
nand U5907 (N_5907,N_4291,N_3907);
nand U5908 (N_5908,N_4995,N_3986);
nor U5909 (N_5909,N_3190,N_4309);
and U5910 (N_5910,N_3664,N_2555);
or U5911 (N_5911,N_4883,N_4645);
and U5912 (N_5912,N_2839,N_4661);
nand U5913 (N_5913,N_2699,N_2734);
and U5914 (N_5914,N_2605,N_4156);
nand U5915 (N_5915,N_3067,N_3546);
nor U5916 (N_5916,N_4836,N_3772);
nor U5917 (N_5917,N_3395,N_4290);
nand U5918 (N_5918,N_3640,N_3353);
or U5919 (N_5919,N_4265,N_3872);
nor U5920 (N_5920,N_3770,N_4599);
or U5921 (N_5921,N_3874,N_3076);
and U5922 (N_5922,N_4811,N_2646);
or U5923 (N_5923,N_3617,N_4116);
or U5924 (N_5924,N_3959,N_3938);
and U5925 (N_5925,N_3407,N_2791);
and U5926 (N_5926,N_4393,N_3158);
xor U5927 (N_5927,N_3250,N_4052);
nor U5928 (N_5928,N_3206,N_2801);
or U5929 (N_5929,N_4055,N_4472);
nor U5930 (N_5930,N_2818,N_4278);
nand U5931 (N_5931,N_4239,N_3130);
nor U5932 (N_5932,N_4198,N_4498);
nor U5933 (N_5933,N_2984,N_3749);
xnor U5934 (N_5934,N_3050,N_3058);
or U5935 (N_5935,N_4088,N_2784);
nand U5936 (N_5936,N_2900,N_4987);
nor U5937 (N_5937,N_3475,N_4068);
or U5938 (N_5938,N_4672,N_4947);
nand U5939 (N_5939,N_2706,N_2803);
nand U5940 (N_5940,N_3561,N_4101);
nand U5941 (N_5941,N_3761,N_4192);
xor U5942 (N_5942,N_4396,N_2543);
nor U5943 (N_5943,N_4627,N_4800);
or U5944 (N_5944,N_4430,N_3243);
nor U5945 (N_5945,N_4886,N_4082);
nor U5946 (N_5946,N_3046,N_3857);
xor U5947 (N_5947,N_3460,N_3781);
nor U5948 (N_5948,N_3370,N_2651);
or U5949 (N_5949,N_4740,N_3485);
nand U5950 (N_5950,N_4926,N_4438);
and U5951 (N_5951,N_4108,N_2865);
nand U5952 (N_5952,N_4019,N_4828);
nand U5953 (N_5953,N_4857,N_4984);
xnor U5954 (N_5954,N_3519,N_3089);
nand U5955 (N_5955,N_4176,N_3812);
or U5956 (N_5956,N_2890,N_4203);
nor U5957 (N_5957,N_3342,N_3726);
and U5958 (N_5958,N_3218,N_4151);
xnor U5959 (N_5959,N_2975,N_3201);
nor U5960 (N_5960,N_2872,N_3943);
and U5961 (N_5961,N_2719,N_4546);
nand U5962 (N_5962,N_4677,N_2519);
and U5963 (N_5963,N_3887,N_4547);
nand U5964 (N_5964,N_4366,N_4227);
and U5965 (N_5965,N_3189,N_3312);
and U5966 (N_5966,N_3314,N_3010);
nand U5967 (N_5967,N_3463,N_2748);
and U5968 (N_5968,N_2595,N_3356);
or U5969 (N_5969,N_3496,N_2944);
nand U5970 (N_5970,N_3361,N_4522);
nor U5971 (N_5971,N_4339,N_4325);
xnor U5972 (N_5972,N_4891,N_2941);
nand U5973 (N_5973,N_3978,N_4899);
or U5974 (N_5974,N_2749,N_3292);
nor U5975 (N_5975,N_3539,N_2862);
nor U5976 (N_5976,N_2752,N_3615);
or U5977 (N_5977,N_3276,N_2658);
and U5978 (N_5978,N_3436,N_4180);
nor U5979 (N_5979,N_4083,N_4385);
nor U5980 (N_5980,N_2754,N_4675);
nand U5981 (N_5981,N_2997,N_3934);
or U5982 (N_5982,N_4274,N_4356);
and U5983 (N_5983,N_3004,N_4540);
and U5984 (N_5984,N_4157,N_3332);
or U5985 (N_5985,N_4787,N_2939);
nor U5986 (N_5986,N_3269,N_4601);
nand U5987 (N_5987,N_2515,N_3266);
and U5988 (N_5988,N_4930,N_2773);
nand U5989 (N_5989,N_2804,N_3502);
xnor U5990 (N_5990,N_2885,N_4404);
nor U5991 (N_5991,N_3338,N_3308);
nor U5992 (N_5992,N_2974,N_4313);
or U5993 (N_5993,N_4738,N_4780);
and U5994 (N_5994,N_3437,N_3623);
nor U5995 (N_5995,N_4354,N_3550);
nor U5996 (N_5996,N_3441,N_4529);
nor U5997 (N_5997,N_2577,N_4243);
nor U5998 (N_5998,N_2745,N_4956);
nor U5999 (N_5999,N_4977,N_3453);
nand U6000 (N_6000,N_4230,N_3344);
xor U6001 (N_6001,N_2521,N_4744);
or U6002 (N_6002,N_2712,N_3474);
and U6003 (N_6003,N_4998,N_4275);
nor U6004 (N_6004,N_4958,N_3428);
nor U6005 (N_6005,N_4029,N_2683);
nand U6006 (N_6006,N_3145,N_4842);
or U6007 (N_6007,N_3425,N_2501);
and U6008 (N_6008,N_4370,N_4338);
or U6009 (N_6009,N_3962,N_3005);
nand U6010 (N_6010,N_3635,N_3763);
and U6011 (N_6011,N_4067,N_4524);
or U6012 (N_6012,N_2681,N_4802);
or U6013 (N_6013,N_2936,N_4255);
and U6014 (N_6014,N_4497,N_3769);
and U6015 (N_6015,N_3618,N_4307);
and U6016 (N_6016,N_4871,N_4929);
or U6017 (N_6017,N_3280,N_3175);
nand U6018 (N_6018,N_4074,N_2563);
nand U6019 (N_6019,N_3367,N_4346);
nand U6020 (N_6020,N_3069,N_3712);
nand U6021 (N_6021,N_4866,N_4989);
and U6022 (N_6022,N_2948,N_3683);
or U6023 (N_6023,N_2679,N_4727);
or U6024 (N_6024,N_3433,N_4293);
and U6025 (N_6025,N_3773,N_4611);
nand U6026 (N_6026,N_3438,N_3195);
nor U6027 (N_6027,N_4351,N_3565);
xnor U6028 (N_6028,N_3745,N_4736);
and U6029 (N_6029,N_3848,N_2963);
nand U6030 (N_6030,N_3450,N_4490);
xor U6031 (N_6031,N_4757,N_2920);
nand U6032 (N_6032,N_2760,N_3871);
or U6033 (N_6033,N_4287,N_3173);
nand U6034 (N_6034,N_4629,N_3483);
and U6035 (N_6035,N_3659,N_4990);
nor U6036 (N_6036,N_4193,N_4453);
nand U6037 (N_6037,N_4931,N_3579);
or U6038 (N_6038,N_3373,N_4311);
nor U6039 (N_6039,N_3184,N_2973);
and U6040 (N_6040,N_3468,N_4739);
or U6041 (N_6041,N_4752,N_4384);
or U6042 (N_6042,N_2867,N_3819);
nor U6043 (N_6043,N_3660,N_3933);
nand U6044 (N_6044,N_3203,N_4657);
nor U6045 (N_6045,N_4415,N_3603);
nor U6046 (N_6046,N_2693,N_4268);
nor U6047 (N_6047,N_3658,N_4973);
nand U6048 (N_6048,N_4328,N_2763);
and U6049 (N_6049,N_3409,N_4233);
xor U6050 (N_6050,N_4341,N_4902);
nand U6051 (N_6051,N_2992,N_4380);
and U6052 (N_6052,N_2977,N_4642);
or U6053 (N_6053,N_4816,N_4263);
nand U6054 (N_6054,N_3346,N_4069);
nor U6055 (N_6055,N_2756,N_3984);
and U6056 (N_6056,N_4473,N_2643);
nor U6057 (N_6057,N_4576,N_3129);
nor U6058 (N_6058,N_2853,N_3242);
or U6059 (N_6059,N_2956,N_3466);
nand U6060 (N_6060,N_3273,N_4544);
nand U6061 (N_6061,N_2830,N_4753);
nor U6062 (N_6062,N_4449,N_3935);
xor U6063 (N_6063,N_4458,N_4130);
nand U6064 (N_6064,N_3248,N_3477);
nor U6065 (N_6065,N_4678,N_3161);
xnor U6066 (N_6066,N_3536,N_4395);
nor U6067 (N_6067,N_3452,N_2898);
and U6068 (N_6068,N_4205,N_2923);
and U6069 (N_6069,N_2876,N_2878);
xor U6070 (N_6070,N_2903,N_3217);
nand U6071 (N_6071,N_3336,N_3278);
xnor U6072 (N_6072,N_4398,N_2516);
nand U6073 (N_6073,N_2911,N_3225);
or U6074 (N_6074,N_4818,N_4579);
nand U6075 (N_6075,N_3791,N_3754);
xor U6076 (N_6076,N_3585,N_3994);
xor U6077 (N_6077,N_3759,N_3020);
xnor U6078 (N_6078,N_3882,N_2617);
xnor U6079 (N_6079,N_4591,N_3041);
xor U6080 (N_6080,N_3594,N_4648);
and U6081 (N_6081,N_4143,N_4361);
or U6082 (N_6082,N_4674,N_4387);
nand U6083 (N_6083,N_2823,N_3911);
nand U6084 (N_6084,N_2632,N_2602);
nand U6085 (N_6085,N_4565,N_3601);
and U6086 (N_6086,N_3862,N_2906);
nand U6087 (N_6087,N_3805,N_4238);
nor U6088 (N_6088,N_2786,N_3170);
nand U6089 (N_6089,N_3045,N_3756);
nand U6090 (N_6090,N_4103,N_3844);
nand U6091 (N_6091,N_3559,N_2529);
nand U6092 (N_6092,N_2731,N_2695);
or U6093 (N_6093,N_2659,N_4023);
and U6094 (N_6094,N_4881,N_3307);
or U6095 (N_6095,N_3143,N_2654);
or U6096 (N_6096,N_3337,N_4032);
nand U6097 (N_6097,N_3590,N_3341);
and U6098 (N_6098,N_2987,N_3397);
and U6099 (N_6099,N_4517,N_3105);
nand U6100 (N_6100,N_2899,N_4904);
nor U6101 (N_6101,N_4922,N_3953);
and U6102 (N_6102,N_3326,N_4846);
or U6103 (N_6103,N_2905,N_2507);
and U6104 (N_6104,N_3272,N_4419);
or U6105 (N_6105,N_4748,N_3180);
or U6106 (N_6106,N_4822,N_4741);
and U6107 (N_6107,N_4724,N_4035);
xor U6108 (N_6108,N_2570,N_3762);
nor U6109 (N_6109,N_4412,N_4624);
and U6110 (N_6110,N_3852,N_4153);
and U6111 (N_6111,N_3349,N_3126);
and U6112 (N_6112,N_3637,N_3890);
nor U6113 (N_6113,N_3263,N_4491);
xnor U6114 (N_6114,N_2759,N_3651);
nor U6115 (N_6115,N_3376,N_3744);
nand U6116 (N_6116,N_2684,N_4715);
and U6117 (N_6117,N_4236,N_3024);
xnor U6118 (N_6118,N_3490,N_2833);
or U6119 (N_6119,N_3078,N_3834);
and U6120 (N_6120,N_3166,N_2649);
or U6121 (N_6121,N_3662,N_4630);
or U6122 (N_6122,N_2526,N_4127);
or U6123 (N_6123,N_4755,N_4406);
nor U6124 (N_6124,N_3746,N_2513);
and U6125 (N_6125,N_4399,N_4201);
nand U6126 (N_6126,N_4917,N_2638);
nand U6127 (N_6127,N_2932,N_2691);
nor U6128 (N_6128,N_4749,N_2846);
nand U6129 (N_6129,N_4803,N_2887);
and U6130 (N_6130,N_4532,N_4885);
or U6131 (N_6131,N_3551,N_2540);
nor U6132 (N_6132,N_4710,N_3340);
nand U6133 (N_6133,N_4196,N_4232);
and U6134 (N_6134,N_3940,N_3629);
xor U6135 (N_6135,N_4251,N_3388);
nor U6136 (N_6136,N_4297,N_3458);
and U6137 (N_6137,N_4580,N_4853);
and U6138 (N_6138,N_4373,N_3447);
and U6139 (N_6139,N_3699,N_3916);
nand U6140 (N_6140,N_2562,N_4482);
and U6141 (N_6141,N_4224,N_4329);
nand U6142 (N_6142,N_2700,N_3222);
xor U6143 (N_6143,N_2580,N_4616);
or U6144 (N_6144,N_2724,N_3806);
nand U6145 (N_6145,N_3778,N_2816);
and U6146 (N_6146,N_2598,N_3246);
nand U6147 (N_6147,N_4047,N_3283);
nor U6148 (N_6148,N_3179,N_4733);
and U6149 (N_6149,N_3144,N_4349);
or U6150 (N_6150,N_4489,N_2926);
or U6151 (N_6151,N_3956,N_2530);
or U6152 (N_6152,N_3902,N_2877);
and U6153 (N_6153,N_3233,N_3609);
nor U6154 (N_6154,N_3411,N_2794);
nor U6155 (N_6155,N_3694,N_2705);
and U6156 (N_6156,N_3289,N_2965);
xnor U6157 (N_6157,N_3432,N_2809);
or U6158 (N_6158,N_4432,N_2765);
and U6159 (N_6159,N_4914,N_4186);
or U6160 (N_6160,N_2814,N_3167);
and U6161 (N_6161,N_4321,N_4681);
or U6162 (N_6162,N_4978,N_3124);
nor U6163 (N_6163,N_4817,N_4394);
xor U6164 (N_6164,N_4638,N_3849);
xor U6165 (N_6165,N_2832,N_3711);
and U6166 (N_6166,N_4125,N_4563);
or U6167 (N_6167,N_2931,N_3758);
and U6168 (N_6168,N_3853,N_2952);
nand U6169 (N_6169,N_4433,N_4093);
and U6170 (N_6170,N_3777,N_3120);
nor U6171 (N_6171,N_4475,N_4344);
nor U6172 (N_6172,N_4695,N_4912);
nand U6173 (N_6173,N_4932,N_2726);
nand U6174 (N_6174,N_4174,N_2821);
nand U6175 (N_6175,N_3279,N_2723);
nand U6176 (N_6176,N_4923,N_4574);
nor U6177 (N_6177,N_4191,N_3608);
nand U6178 (N_6178,N_2881,N_3839);
and U6179 (N_6179,N_4277,N_2600);
nor U6180 (N_6180,N_4141,N_4267);
and U6181 (N_6181,N_2894,N_4340);
nand U6182 (N_6182,N_4781,N_3755);
nor U6183 (N_6183,N_3695,N_2564);
nand U6184 (N_6184,N_3829,N_2722);
and U6185 (N_6185,N_4805,N_3488);
and U6186 (N_6186,N_2601,N_3094);
or U6187 (N_6187,N_3817,N_3979);
nor U6188 (N_6188,N_2717,N_2606);
xor U6189 (N_6189,N_4538,N_4635);
or U6190 (N_6190,N_3545,N_4091);
xor U6191 (N_6191,N_3782,N_4996);
nand U6192 (N_6192,N_2742,N_3846);
nor U6193 (N_6193,N_2779,N_3362);
xnor U6194 (N_6194,N_4378,N_2817);
nor U6195 (N_6195,N_2592,N_3347);
nor U6196 (N_6196,N_4776,N_4058);
or U6197 (N_6197,N_4381,N_3880);
or U6198 (N_6198,N_4018,N_4121);
or U6199 (N_6199,N_2551,N_3403);
nor U6200 (N_6200,N_2796,N_3624);
and U6201 (N_6201,N_4004,N_3472);
and U6202 (N_6202,N_2945,N_4081);
nand U6203 (N_6203,N_3915,N_3613);
xor U6204 (N_6204,N_4558,N_4168);
or U6205 (N_6205,N_4454,N_2792);
nor U6206 (N_6206,N_4523,N_2613);
nor U6207 (N_6207,N_3633,N_3051);
and U6208 (N_6208,N_4342,N_3583);
nand U6209 (N_6209,N_4707,N_4609);
xnor U6210 (N_6210,N_4401,N_4166);
xnor U6211 (N_6211,N_3584,N_3333);
and U6212 (N_6212,N_3741,N_2912);
and U6213 (N_6213,N_3976,N_3305);
and U6214 (N_6214,N_3549,N_4056);
or U6215 (N_6215,N_3790,N_3861);
and U6216 (N_6216,N_2661,N_2960);
or U6217 (N_6217,N_3476,N_4479);
nor U6218 (N_6218,N_3732,N_2849);
or U6219 (N_6219,N_4383,N_4607);
xor U6220 (N_6220,N_3980,N_4327);
nor U6221 (N_6221,N_3270,N_4261);
nand U6222 (N_6222,N_4345,N_3730);
or U6223 (N_6223,N_4147,N_3958);
nand U6224 (N_6224,N_4610,N_4988);
and U6225 (N_6225,N_4570,N_2969);
nand U6226 (N_6226,N_4257,N_2886);
nor U6227 (N_6227,N_3865,N_4571);
nand U6228 (N_6228,N_2828,N_4841);
nor U6229 (N_6229,N_4030,N_3097);
xor U6230 (N_6230,N_3191,N_2758);
or U6231 (N_6231,N_3569,N_2652);
or U6232 (N_6232,N_2985,N_2916);
and U6233 (N_6233,N_4254,N_4663);
nand U6234 (N_6234,N_4452,N_4992);
or U6235 (N_6235,N_3131,N_3802);
nor U6236 (N_6236,N_4552,N_4685);
nor U6237 (N_6237,N_3369,N_4530);
nand U6238 (N_6238,N_3521,N_3783);
nand U6239 (N_6239,N_2640,N_4424);
nor U6240 (N_6240,N_4829,N_4867);
and U6241 (N_6241,N_4122,N_3859);
and U6242 (N_6242,N_2996,N_4712);
or U6243 (N_6243,N_3910,N_3752);
nor U6244 (N_6244,N_3870,N_3964);
and U6245 (N_6245,N_3698,N_3927);
xor U6246 (N_6246,N_4957,N_3522);
or U6247 (N_6247,N_4065,N_3102);
xor U6248 (N_6248,N_4397,N_4124);
or U6249 (N_6249,N_2908,N_2615);
xor U6250 (N_6250,N_3084,N_3902);
and U6251 (N_6251,N_3676,N_4623);
nor U6252 (N_6252,N_3002,N_3333);
nand U6253 (N_6253,N_3000,N_4885);
xnor U6254 (N_6254,N_4074,N_3300);
or U6255 (N_6255,N_4299,N_4444);
or U6256 (N_6256,N_2840,N_4225);
or U6257 (N_6257,N_2795,N_4545);
nand U6258 (N_6258,N_3483,N_4321);
or U6259 (N_6259,N_3783,N_3915);
or U6260 (N_6260,N_4771,N_3142);
nor U6261 (N_6261,N_4029,N_3711);
or U6262 (N_6262,N_4009,N_4834);
nor U6263 (N_6263,N_2944,N_3781);
or U6264 (N_6264,N_4543,N_4509);
or U6265 (N_6265,N_4995,N_3552);
nand U6266 (N_6266,N_3959,N_2782);
xor U6267 (N_6267,N_3529,N_2906);
nor U6268 (N_6268,N_2952,N_3901);
nand U6269 (N_6269,N_4986,N_3553);
nor U6270 (N_6270,N_3714,N_2539);
nor U6271 (N_6271,N_4030,N_4222);
xor U6272 (N_6272,N_4453,N_4441);
and U6273 (N_6273,N_3773,N_4104);
or U6274 (N_6274,N_4359,N_4949);
nor U6275 (N_6275,N_3322,N_4335);
nor U6276 (N_6276,N_4044,N_4474);
and U6277 (N_6277,N_3224,N_3569);
nand U6278 (N_6278,N_4722,N_3020);
xnor U6279 (N_6279,N_3411,N_4671);
nor U6280 (N_6280,N_3446,N_3903);
nor U6281 (N_6281,N_4211,N_4964);
nor U6282 (N_6282,N_4119,N_3095);
xor U6283 (N_6283,N_2811,N_3756);
or U6284 (N_6284,N_3231,N_3212);
or U6285 (N_6285,N_3166,N_2569);
nor U6286 (N_6286,N_3062,N_4925);
or U6287 (N_6287,N_3361,N_2893);
nor U6288 (N_6288,N_4065,N_4092);
nor U6289 (N_6289,N_3716,N_2799);
or U6290 (N_6290,N_3614,N_4689);
or U6291 (N_6291,N_2853,N_4545);
and U6292 (N_6292,N_3170,N_2563);
or U6293 (N_6293,N_2866,N_3105);
or U6294 (N_6294,N_3968,N_3914);
nor U6295 (N_6295,N_3350,N_4031);
nand U6296 (N_6296,N_4617,N_3769);
or U6297 (N_6297,N_3746,N_2516);
and U6298 (N_6298,N_3236,N_4544);
nand U6299 (N_6299,N_4302,N_3939);
nor U6300 (N_6300,N_4822,N_3551);
and U6301 (N_6301,N_3539,N_4032);
or U6302 (N_6302,N_2949,N_4953);
nand U6303 (N_6303,N_2704,N_3542);
nor U6304 (N_6304,N_4898,N_2508);
and U6305 (N_6305,N_3839,N_3670);
xnor U6306 (N_6306,N_3137,N_4658);
and U6307 (N_6307,N_2796,N_4110);
nor U6308 (N_6308,N_4550,N_3255);
nor U6309 (N_6309,N_3486,N_2772);
nor U6310 (N_6310,N_4995,N_3832);
nand U6311 (N_6311,N_2673,N_4947);
nor U6312 (N_6312,N_3010,N_2933);
nor U6313 (N_6313,N_2637,N_4214);
nor U6314 (N_6314,N_3830,N_3656);
nand U6315 (N_6315,N_2976,N_3446);
or U6316 (N_6316,N_4741,N_2906);
nand U6317 (N_6317,N_2978,N_3495);
or U6318 (N_6318,N_3619,N_4392);
xor U6319 (N_6319,N_2802,N_4089);
nor U6320 (N_6320,N_4842,N_3457);
xnor U6321 (N_6321,N_3044,N_2697);
nor U6322 (N_6322,N_4317,N_4449);
xor U6323 (N_6323,N_3011,N_4387);
and U6324 (N_6324,N_2651,N_2741);
or U6325 (N_6325,N_3288,N_4253);
or U6326 (N_6326,N_2622,N_4841);
and U6327 (N_6327,N_3928,N_4114);
nand U6328 (N_6328,N_3170,N_3282);
and U6329 (N_6329,N_2849,N_4856);
nand U6330 (N_6330,N_3219,N_4047);
and U6331 (N_6331,N_3637,N_2541);
and U6332 (N_6332,N_2897,N_2818);
nand U6333 (N_6333,N_3491,N_4472);
and U6334 (N_6334,N_4745,N_4230);
and U6335 (N_6335,N_4509,N_3783);
or U6336 (N_6336,N_2621,N_4829);
nand U6337 (N_6337,N_4061,N_2844);
nor U6338 (N_6338,N_4593,N_3088);
nand U6339 (N_6339,N_3090,N_4775);
nand U6340 (N_6340,N_2546,N_3776);
nand U6341 (N_6341,N_4253,N_4219);
nand U6342 (N_6342,N_2702,N_3611);
xnor U6343 (N_6343,N_4850,N_3379);
or U6344 (N_6344,N_3219,N_2500);
or U6345 (N_6345,N_3568,N_2761);
and U6346 (N_6346,N_2689,N_3173);
nor U6347 (N_6347,N_4625,N_3183);
nor U6348 (N_6348,N_2706,N_4725);
and U6349 (N_6349,N_3187,N_3292);
nor U6350 (N_6350,N_4752,N_4506);
nor U6351 (N_6351,N_2711,N_2956);
or U6352 (N_6352,N_4902,N_4550);
and U6353 (N_6353,N_2685,N_4105);
or U6354 (N_6354,N_3902,N_4759);
or U6355 (N_6355,N_2655,N_3508);
and U6356 (N_6356,N_4342,N_3939);
nand U6357 (N_6357,N_2932,N_3286);
or U6358 (N_6358,N_3283,N_3728);
nand U6359 (N_6359,N_3275,N_4770);
and U6360 (N_6360,N_3515,N_3504);
or U6361 (N_6361,N_4095,N_3292);
xor U6362 (N_6362,N_4990,N_4736);
nor U6363 (N_6363,N_2780,N_3687);
nand U6364 (N_6364,N_3988,N_2589);
and U6365 (N_6365,N_3805,N_4115);
and U6366 (N_6366,N_2515,N_2796);
nand U6367 (N_6367,N_3319,N_3808);
nand U6368 (N_6368,N_3126,N_2677);
nand U6369 (N_6369,N_3944,N_2637);
nand U6370 (N_6370,N_2981,N_2830);
or U6371 (N_6371,N_4002,N_4664);
and U6372 (N_6372,N_4988,N_4976);
xnor U6373 (N_6373,N_3484,N_4229);
nand U6374 (N_6374,N_4204,N_3279);
and U6375 (N_6375,N_2714,N_3171);
nand U6376 (N_6376,N_2738,N_4690);
nand U6377 (N_6377,N_4038,N_2927);
nand U6378 (N_6378,N_4303,N_3460);
and U6379 (N_6379,N_3416,N_3508);
or U6380 (N_6380,N_3042,N_3957);
or U6381 (N_6381,N_4301,N_2618);
and U6382 (N_6382,N_3201,N_4983);
nor U6383 (N_6383,N_4943,N_2742);
or U6384 (N_6384,N_3865,N_4756);
and U6385 (N_6385,N_2564,N_3481);
or U6386 (N_6386,N_2674,N_3383);
and U6387 (N_6387,N_2835,N_4343);
xor U6388 (N_6388,N_3276,N_4602);
and U6389 (N_6389,N_4773,N_2967);
and U6390 (N_6390,N_3658,N_4618);
nor U6391 (N_6391,N_4610,N_3762);
and U6392 (N_6392,N_4821,N_4204);
or U6393 (N_6393,N_3702,N_4356);
nand U6394 (N_6394,N_4095,N_4584);
nand U6395 (N_6395,N_3700,N_3511);
nand U6396 (N_6396,N_4994,N_3461);
nor U6397 (N_6397,N_4925,N_4947);
nand U6398 (N_6398,N_3614,N_3776);
and U6399 (N_6399,N_3944,N_4046);
nand U6400 (N_6400,N_3770,N_3582);
nand U6401 (N_6401,N_3656,N_4587);
or U6402 (N_6402,N_4703,N_3476);
and U6403 (N_6403,N_4675,N_3443);
or U6404 (N_6404,N_3704,N_3954);
nand U6405 (N_6405,N_3184,N_4640);
nor U6406 (N_6406,N_3233,N_4912);
nor U6407 (N_6407,N_2964,N_4123);
or U6408 (N_6408,N_2591,N_4902);
nor U6409 (N_6409,N_4868,N_3799);
or U6410 (N_6410,N_4091,N_4468);
or U6411 (N_6411,N_2584,N_4969);
or U6412 (N_6412,N_4686,N_2660);
xor U6413 (N_6413,N_3624,N_4885);
or U6414 (N_6414,N_3963,N_3614);
or U6415 (N_6415,N_2863,N_3450);
and U6416 (N_6416,N_3971,N_4656);
nor U6417 (N_6417,N_4711,N_3796);
nand U6418 (N_6418,N_4856,N_4036);
or U6419 (N_6419,N_3992,N_2923);
nand U6420 (N_6420,N_4287,N_3861);
and U6421 (N_6421,N_3007,N_4015);
or U6422 (N_6422,N_4278,N_4230);
and U6423 (N_6423,N_2984,N_3195);
nor U6424 (N_6424,N_2543,N_4455);
xnor U6425 (N_6425,N_2615,N_4945);
nand U6426 (N_6426,N_2642,N_4333);
nand U6427 (N_6427,N_4137,N_2745);
xnor U6428 (N_6428,N_4030,N_2602);
and U6429 (N_6429,N_4155,N_2647);
or U6430 (N_6430,N_2901,N_3289);
xor U6431 (N_6431,N_4366,N_2545);
nand U6432 (N_6432,N_2542,N_4414);
and U6433 (N_6433,N_3619,N_3776);
and U6434 (N_6434,N_4302,N_4473);
nand U6435 (N_6435,N_2987,N_4608);
xnor U6436 (N_6436,N_3121,N_2793);
or U6437 (N_6437,N_3705,N_4431);
xnor U6438 (N_6438,N_3609,N_3851);
or U6439 (N_6439,N_3756,N_3762);
xor U6440 (N_6440,N_2877,N_4432);
and U6441 (N_6441,N_3140,N_4445);
nand U6442 (N_6442,N_4763,N_4444);
nor U6443 (N_6443,N_3601,N_3706);
and U6444 (N_6444,N_4742,N_3196);
or U6445 (N_6445,N_3131,N_4035);
nor U6446 (N_6446,N_4036,N_2686);
nand U6447 (N_6447,N_3054,N_4223);
nand U6448 (N_6448,N_4930,N_4522);
xor U6449 (N_6449,N_4809,N_2525);
xnor U6450 (N_6450,N_3981,N_4330);
nor U6451 (N_6451,N_4482,N_4650);
nor U6452 (N_6452,N_3225,N_2650);
or U6453 (N_6453,N_4301,N_3729);
nand U6454 (N_6454,N_2503,N_4949);
nor U6455 (N_6455,N_4796,N_3448);
and U6456 (N_6456,N_3073,N_2524);
nor U6457 (N_6457,N_2998,N_2741);
and U6458 (N_6458,N_4319,N_3301);
and U6459 (N_6459,N_3220,N_3173);
or U6460 (N_6460,N_3668,N_3679);
xnor U6461 (N_6461,N_2896,N_2727);
or U6462 (N_6462,N_4679,N_3182);
nand U6463 (N_6463,N_3395,N_4583);
and U6464 (N_6464,N_3410,N_3863);
or U6465 (N_6465,N_3584,N_2694);
nor U6466 (N_6466,N_3700,N_3674);
nor U6467 (N_6467,N_2678,N_2953);
or U6468 (N_6468,N_4745,N_4992);
xor U6469 (N_6469,N_3102,N_3462);
nand U6470 (N_6470,N_3015,N_4628);
xor U6471 (N_6471,N_4735,N_4908);
xnor U6472 (N_6472,N_2743,N_4911);
nor U6473 (N_6473,N_4429,N_4884);
xnor U6474 (N_6474,N_3861,N_4281);
and U6475 (N_6475,N_2561,N_3737);
and U6476 (N_6476,N_2566,N_3529);
or U6477 (N_6477,N_2733,N_4482);
or U6478 (N_6478,N_2963,N_4722);
nor U6479 (N_6479,N_4200,N_3467);
xnor U6480 (N_6480,N_4283,N_4365);
and U6481 (N_6481,N_3847,N_2877);
xor U6482 (N_6482,N_4398,N_2674);
nand U6483 (N_6483,N_2792,N_3033);
nand U6484 (N_6484,N_3058,N_4986);
or U6485 (N_6485,N_4320,N_4414);
nor U6486 (N_6486,N_2573,N_4668);
nand U6487 (N_6487,N_4509,N_2944);
and U6488 (N_6488,N_4755,N_4659);
and U6489 (N_6489,N_3056,N_4566);
nand U6490 (N_6490,N_3960,N_4905);
nand U6491 (N_6491,N_4391,N_3078);
nand U6492 (N_6492,N_3756,N_3686);
nand U6493 (N_6493,N_3066,N_2659);
or U6494 (N_6494,N_3994,N_2856);
nand U6495 (N_6495,N_4062,N_4155);
nor U6496 (N_6496,N_3669,N_2577);
nor U6497 (N_6497,N_3185,N_4792);
nor U6498 (N_6498,N_4504,N_2973);
and U6499 (N_6499,N_3548,N_3989);
or U6500 (N_6500,N_3358,N_4599);
nor U6501 (N_6501,N_3686,N_3996);
nor U6502 (N_6502,N_2501,N_3835);
and U6503 (N_6503,N_4782,N_3281);
and U6504 (N_6504,N_2633,N_3383);
or U6505 (N_6505,N_3011,N_4588);
xor U6506 (N_6506,N_2551,N_3040);
and U6507 (N_6507,N_2520,N_3343);
nand U6508 (N_6508,N_3752,N_3930);
and U6509 (N_6509,N_2646,N_2656);
xor U6510 (N_6510,N_3819,N_4384);
and U6511 (N_6511,N_2987,N_4235);
or U6512 (N_6512,N_4217,N_3794);
nand U6513 (N_6513,N_3467,N_3504);
or U6514 (N_6514,N_3379,N_3279);
and U6515 (N_6515,N_3157,N_4039);
or U6516 (N_6516,N_4709,N_4941);
nand U6517 (N_6517,N_3312,N_3456);
nand U6518 (N_6518,N_4995,N_2723);
xnor U6519 (N_6519,N_4560,N_2894);
nor U6520 (N_6520,N_2888,N_2609);
nand U6521 (N_6521,N_4720,N_3626);
nor U6522 (N_6522,N_3618,N_3316);
nand U6523 (N_6523,N_2566,N_3093);
nor U6524 (N_6524,N_4553,N_3167);
or U6525 (N_6525,N_2510,N_3400);
nand U6526 (N_6526,N_4938,N_3359);
or U6527 (N_6527,N_4621,N_3984);
and U6528 (N_6528,N_4303,N_3275);
and U6529 (N_6529,N_3406,N_2879);
nor U6530 (N_6530,N_4185,N_3436);
nand U6531 (N_6531,N_4587,N_4779);
and U6532 (N_6532,N_4144,N_3392);
and U6533 (N_6533,N_3195,N_3255);
nor U6534 (N_6534,N_3003,N_4804);
nand U6535 (N_6535,N_2622,N_4961);
nand U6536 (N_6536,N_3342,N_2973);
nor U6537 (N_6537,N_3151,N_2902);
and U6538 (N_6538,N_4118,N_2623);
or U6539 (N_6539,N_3239,N_3175);
and U6540 (N_6540,N_3519,N_3189);
nand U6541 (N_6541,N_4428,N_4189);
or U6542 (N_6542,N_4775,N_2797);
or U6543 (N_6543,N_4924,N_4587);
and U6544 (N_6544,N_4420,N_3510);
nor U6545 (N_6545,N_2601,N_3354);
nand U6546 (N_6546,N_4504,N_4216);
xnor U6547 (N_6547,N_2664,N_2799);
xnor U6548 (N_6548,N_3390,N_4118);
and U6549 (N_6549,N_4548,N_2886);
nor U6550 (N_6550,N_3514,N_2905);
nor U6551 (N_6551,N_3040,N_4179);
nor U6552 (N_6552,N_4729,N_4849);
or U6553 (N_6553,N_3018,N_3787);
nor U6554 (N_6554,N_2729,N_3338);
nor U6555 (N_6555,N_2689,N_4927);
and U6556 (N_6556,N_3390,N_3045);
nor U6557 (N_6557,N_3745,N_3928);
or U6558 (N_6558,N_3303,N_4823);
or U6559 (N_6559,N_3049,N_4317);
and U6560 (N_6560,N_4474,N_2668);
nor U6561 (N_6561,N_4054,N_3816);
nor U6562 (N_6562,N_4965,N_2694);
and U6563 (N_6563,N_3855,N_4148);
nor U6564 (N_6564,N_3840,N_4241);
nor U6565 (N_6565,N_4737,N_3861);
or U6566 (N_6566,N_3114,N_3519);
nand U6567 (N_6567,N_3636,N_3792);
or U6568 (N_6568,N_3190,N_3380);
nor U6569 (N_6569,N_4452,N_3581);
or U6570 (N_6570,N_4516,N_3008);
or U6571 (N_6571,N_2873,N_4428);
nor U6572 (N_6572,N_4139,N_4019);
and U6573 (N_6573,N_4434,N_4851);
nor U6574 (N_6574,N_3026,N_2876);
and U6575 (N_6575,N_3372,N_4923);
nand U6576 (N_6576,N_3610,N_3420);
and U6577 (N_6577,N_4415,N_4086);
or U6578 (N_6578,N_3270,N_2922);
or U6579 (N_6579,N_4970,N_4597);
or U6580 (N_6580,N_4137,N_4469);
xor U6581 (N_6581,N_3824,N_3472);
or U6582 (N_6582,N_3352,N_3179);
xnor U6583 (N_6583,N_3288,N_2592);
and U6584 (N_6584,N_3000,N_4559);
nor U6585 (N_6585,N_3268,N_4137);
and U6586 (N_6586,N_3305,N_3179);
nor U6587 (N_6587,N_3237,N_2895);
or U6588 (N_6588,N_4468,N_4070);
or U6589 (N_6589,N_4901,N_2812);
nand U6590 (N_6590,N_3152,N_2946);
or U6591 (N_6591,N_4264,N_4311);
or U6592 (N_6592,N_4943,N_3858);
nand U6593 (N_6593,N_3242,N_4062);
nor U6594 (N_6594,N_3547,N_4195);
nand U6595 (N_6595,N_4413,N_4926);
nor U6596 (N_6596,N_3570,N_3503);
xnor U6597 (N_6597,N_4556,N_3244);
or U6598 (N_6598,N_3385,N_4525);
and U6599 (N_6599,N_3958,N_4169);
or U6600 (N_6600,N_2816,N_3533);
nand U6601 (N_6601,N_2714,N_3176);
xnor U6602 (N_6602,N_3140,N_4222);
nor U6603 (N_6603,N_4441,N_4935);
nor U6604 (N_6604,N_3253,N_4009);
or U6605 (N_6605,N_2909,N_3455);
or U6606 (N_6606,N_4176,N_4726);
and U6607 (N_6607,N_4929,N_3343);
nor U6608 (N_6608,N_4895,N_4593);
xnor U6609 (N_6609,N_4467,N_3615);
nand U6610 (N_6610,N_4810,N_4241);
nor U6611 (N_6611,N_3973,N_4753);
or U6612 (N_6612,N_4046,N_4111);
or U6613 (N_6613,N_4246,N_4483);
nand U6614 (N_6614,N_4758,N_3169);
nor U6615 (N_6615,N_2553,N_3180);
nand U6616 (N_6616,N_4046,N_3031);
nand U6617 (N_6617,N_3285,N_2823);
nor U6618 (N_6618,N_2627,N_3641);
nor U6619 (N_6619,N_4192,N_4700);
nor U6620 (N_6620,N_2530,N_4961);
and U6621 (N_6621,N_4094,N_3160);
xor U6622 (N_6622,N_2707,N_4783);
nand U6623 (N_6623,N_3390,N_3948);
or U6624 (N_6624,N_2598,N_3585);
or U6625 (N_6625,N_3734,N_3421);
nand U6626 (N_6626,N_4143,N_3470);
or U6627 (N_6627,N_3349,N_3388);
nor U6628 (N_6628,N_2817,N_4093);
nand U6629 (N_6629,N_4740,N_3719);
xnor U6630 (N_6630,N_3580,N_3848);
nand U6631 (N_6631,N_4091,N_4726);
and U6632 (N_6632,N_3753,N_4147);
xor U6633 (N_6633,N_3068,N_3098);
and U6634 (N_6634,N_3062,N_2801);
or U6635 (N_6635,N_2939,N_3225);
nor U6636 (N_6636,N_3587,N_4099);
xnor U6637 (N_6637,N_4257,N_3405);
and U6638 (N_6638,N_3959,N_4563);
xor U6639 (N_6639,N_3231,N_4402);
or U6640 (N_6640,N_3628,N_3241);
nor U6641 (N_6641,N_3205,N_3750);
xnor U6642 (N_6642,N_3181,N_3219);
and U6643 (N_6643,N_4818,N_3201);
and U6644 (N_6644,N_2868,N_3209);
or U6645 (N_6645,N_3402,N_2802);
nand U6646 (N_6646,N_3887,N_4050);
or U6647 (N_6647,N_4922,N_4103);
or U6648 (N_6648,N_3027,N_3563);
and U6649 (N_6649,N_4863,N_4699);
nor U6650 (N_6650,N_3751,N_4229);
or U6651 (N_6651,N_4000,N_2898);
and U6652 (N_6652,N_4181,N_2610);
nor U6653 (N_6653,N_3824,N_4238);
nand U6654 (N_6654,N_4059,N_4562);
and U6655 (N_6655,N_4709,N_2779);
or U6656 (N_6656,N_3410,N_3964);
and U6657 (N_6657,N_4869,N_3633);
and U6658 (N_6658,N_3415,N_4173);
nand U6659 (N_6659,N_4797,N_2874);
and U6660 (N_6660,N_2724,N_4673);
xor U6661 (N_6661,N_3393,N_3730);
nand U6662 (N_6662,N_4304,N_4104);
nor U6663 (N_6663,N_3297,N_3668);
or U6664 (N_6664,N_4508,N_3353);
or U6665 (N_6665,N_2536,N_4979);
xnor U6666 (N_6666,N_3773,N_3157);
or U6667 (N_6667,N_4781,N_4719);
xor U6668 (N_6668,N_4669,N_3370);
nor U6669 (N_6669,N_3490,N_4180);
nor U6670 (N_6670,N_3085,N_3091);
or U6671 (N_6671,N_3833,N_3011);
xor U6672 (N_6672,N_3534,N_4064);
or U6673 (N_6673,N_3956,N_2772);
or U6674 (N_6674,N_4483,N_3275);
or U6675 (N_6675,N_3547,N_4176);
nor U6676 (N_6676,N_4914,N_4921);
nand U6677 (N_6677,N_4606,N_4052);
nor U6678 (N_6678,N_4900,N_2501);
xnor U6679 (N_6679,N_3110,N_3283);
or U6680 (N_6680,N_4707,N_3268);
and U6681 (N_6681,N_2938,N_3638);
nand U6682 (N_6682,N_3659,N_3003);
and U6683 (N_6683,N_3238,N_2897);
or U6684 (N_6684,N_3525,N_2944);
nand U6685 (N_6685,N_4166,N_3980);
nand U6686 (N_6686,N_3030,N_2818);
nand U6687 (N_6687,N_3463,N_3864);
and U6688 (N_6688,N_3320,N_3494);
nand U6689 (N_6689,N_4303,N_4626);
nor U6690 (N_6690,N_2663,N_4374);
xnor U6691 (N_6691,N_3298,N_4729);
nor U6692 (N_6692,N_2750,N_4433);
xor U6693 (N_6693,N_3956,N_4880);
xor U6694 (N_6694,N_4580,N_2766);
nor U6695 (N_6695,N_2530,N_3714);
or U6696 (N_6696,N_4461,N_4081);
nand U6697 (N_6697,N_3944,N_4162);
or U6698 (N_6698,N_3971,N_3101);
or U6699 (N_6699,N_4648,N_2683);
nor U6700 (N_6700,N_3844,N_2836);
and U6701 (N_6701,N_3203,N_4211);
and U6702 (N_6702,N_4775,N_3321);
nand U6703 (N_6703,N_4902,N_3027);
nand U6704 (N_6704,N_3732,N_4534);
xnor U6705 (N_6705,N_3330,N_4040);
nand U6706 (N_6706,N_3539,N_3765);
nand U6707 (N_6707,N_4929,N_2613);
xnor U6708 (N_6708,N_3920,N_4292);
xor U6709 (N_6709,N_4085,N_3707);
nor U6710 (N_6710,N_2899,N_4933);
xnor U6711 (N_6711,N_4233,N_2764);
xnor U6712 (N_6712,N_4855,N_4968);
and U6713 (N_6713,N_4417,N_3663);
and U6714 (N_6714,N_2693,N_4364);
nand U6715 (N_6715,N_2971,N_4591);
nor U6716 (N_6716,N_2893,N_3353);
nand U6717 (N_6717,N_2816,N_2927);
xor U6718 (N_6718,N_4457,N_3191);
or U6719 (N_6719,N_3100,N_4122);
and U6720 (N_6720,N_3338,N_3877);
xnor U6721 (N_6721,N_4638,N_4506);
or U6722 (N_6722,N_2792,N_2817);
xor U6723 (N_6723,N_4667,N_4551);
nand U6724 (N_6724,N_3010,N_3539);
and U6725 (N_6725,N_3655,N_3601);
and U6726 (N_6726,N_3747,N_2641);
or U6727 (N_6727,N_3550,N_3484);
nand U6728 (N_6728,N_2631,N_4290);
nand U6729 (N_6729,N_3990,N_4753);
xnor U6730 (N_6730,N_4103,N_2549);
nand U6731 (N_6731,N_3465,N_3575);
nor U6732 (N_6732,N_3749,N_4543);
or U6733 (N_6733,N_3867,N_4178);
xor U6734 (N_6734,N_4834,N_4525);
nand U6735 (N_6735,N_2577,N_3648);
and U6736 (N_6736,N_3918,N_3222);
nor U6737 (N_6737,N_4418,N_3260);
nand U6738 (N_6738,N_4381,N_4470);
or U6739 (N_6739,N_3783,N_4876);
nor U6740 (N_6740,N_4788,N_2962);
or U6741 (N_6741,N_3561,N_4356);
and U6742 (N_6742,N_2662,N_4976);
nor U6743 (N_6743,N_4937,N_2860);
or U6744 (N_6744,N_2535,N_4596);
and U6745 (N_6745,N_2762,N_3818);
nand U6746 (N_6746,N_3757,N_4983);
xor U6747 (N_6747,N_4211,N_3154);
nor U6748 (N_6748,N_2622,N_4219);
or U6749 (N_6749,N_4322,N_3532);
or U6750 (N_6750,N_4543,N_3544);
nand U6751 (N_6751,N_3110,N_3043);
and U6752 (N_6752,N_4221,N_4060);
xnor U6753 (N_6753,N_3196,N_3935);
nand U6754 (N_6754,N_4175,N_2823);
nor U6755 (N_6755,N_3695,N_4541);
xor U6756 (N_6756,N_3187,N_3676);
and U6757 (N_6757,N_3496,N_3383);
nor U6758 (N_6758,N_4244,N_4671);
nor U6759 (N_6759,N_4541,N_4215);
nor U6760 (N_6760,N_3797,N_4761);
xnor U6761 (N_6761,N_2896,N_4874);
nor U6762 (N_6762,N_3230,N_3589);
or U6763 (N_6763,N_4755,N_2952);
and U6764 (N_6764,N_3106,N_3927);
nand U6765 (N_6765,N_3111,N_4164);
nor U6766 (N_6766,N_4339,N_3874);
nand U6767 (N_6767,N_2870,N_4638);
or U6768 (N_6768,N_4593,N_3827);
or U6769 (N_6769,N_3260,N_3422);
or U6770 (N_6770,N_4611,N_4521);
or U6771 (N_6771,N_4125,N_4829);
nor U6772 (N_6772,N_4002,N_3012);
nand U6773 (N_6773,N_4004,N_3419);
nand U6774 (N_6774,N_2958,N_4446);
nand U6775 (N_6775,N_2959,N_3523);
and U6776 (N_6776,N_2766,N_3974);
xnor U6777 (N_6777,N_4790,N_4583);
nand U6778 (N_6778,N_3663,N_4246);
nand U6779 (N_6779,N_4277,N_2904);
and U6780 (N_6780,N_3655,N_3259);
or U6781 (N_6781,N_2519,N_3747);
xor U6782 (N_6782,N_2708,N_3026);
nor U6783 (N_6783,N_3883,N_3940);
and U6784 (N_6784,N_3550,N_3735);
nor U6785 (N_6785,N_2679,N_4238);
nor U6786 (N_6786,N_4438,N_4001);
xnor U6787 (N_6787,N_4483,N_4181);
and U6788 (N_6788,N_2806,N_2627);
xor U6789 (N_6789,N_2523,N_2894);
and U6790 (N_6790,N_4307,N_4990);
nand U6791 (N_6791,N_4828,N_2697);
or U6792 (N_6792,N_2611,N_3310);
and U6793 (N_6793,N_4711,N_3957);
nor U6794 (N_6794,N_2882,N_4346);
or U6795 (N_6795,N_4441,N_3504);
and U6796 (N_6796,N_4034,N_2993);
and U6797 (N_6797,N_2791,N_2617);
nor U6798 (N_6798,N_3218,N_2863);
or U6799 (N_6799,N_3848,N_4624);
and U6800 (N_6800,N_2729,N_4944);
xnor U6801 (N_6801,N_2562,N_3910);
nor U6802 (N_6802,N_3537,N_4813);
nor U6803 (N_6803,N_4592,N_3056);
nand U6804 (N_6804,N_4845,N_3574);
nand U6805 (N_6805,N_3817,N_3045);
nor U6806 (N_6806,N_3583,N_3232);
nor U6807 (N_6807,N_4895,N_2703);
nor U6808 (N_6808,N_3419,N_2697);
xnor U6809 (N_6809,N_3637,N_3845);
xor U6810 (N_6810,N_3543,N_4505);
nor U6811 (N_6811,N_3138,N_4010);
nor U6812 (N_6812,N_3725,N_3396);
nor U6813 (N_6813,N_4890,N_4275);
nor U6814 (N_6814,N_3092,N_2758);
or U6815 (N_6815,N_3137,N_3869);
xor U6816 (N_6816,N_4898,N_4133);
and U6817 (N_6817,N_4363,N_4225);
nand U6818 (N_6818,N_4693,N_4452);
nand U6819 (N_6819,N_4162,N_3284);
nor U6820 (N_6820,N_3242,N_3391);
nor U6821 (N_6821,N_2511,N_4702);
and U6822 (N_6822,N_4772,N_3715);
nor U6823 (N_6823,N_3155,N_3508);
xor U6824 (N_6824,N_3130,N_3056);
and U6825 (N_6825,N_3772,N_4233);
xor U6826 (N_6826,N_2722,N_4212);
nor U6827 (N_6827,N_3726,N_3461);
nor U6828 (N_6828,N_3480,N_4532);
or U6829 (N_6829,N_2846,N_3717);
and U6830 (N_6830,N_4882,N_2636);
and U6831 (N_6831,N_4108,N_4398);
nand U6832 (N_6832,N_3490,N_4946);
xor U6833 (N_6833,N_3605,N_4080);
and U6834 (N_6834,N_4068,N_3474);
and U6835 (N_6835,N_4691,N_3116);
or U6836 (N_6836,N_3673,N_4686);
and U6837 (N_6837,N_3375,N_3953);
and U6838 (N_6838,N_4550,N_3438);
or U6839 (N_6839,N_4705,N_2693);
nor U6840 (N_6840,N_4973,N_4898);
nor U6841 (N_6841,N_3314,N_4905);
nand U6842 (N_6842,N_4458,N_2920);
nand U6843 (N_6843,N_4716,N_3773);
nand U6844 (N_6844,N_4886,N_4970);
xor U6845 (N_6845,N_2566,N_3838);
or U6846 (N_6846,N_3893,N_2522);
nor U6847 (N_6847,N_4082,N_3057);
and U6848 (N_6848,N_4855,N_4957);
or U6849 (N_6849,N_2649,N_4482);
and U6850 (N_6850,N_2695,N_4220);
and U6851 (N_6851,N_3454,N_4600);
or U6852 (N_6852,N_4829,N_4149);
or U6853 (N_6853,N_4484,N_3766);
or U6854 (N_6854,N_2908,N_4382);
or U6855 (N_6855,N_2982,N_3907);
nor U6856 (N_6856,N_3531,N_4324);
or U6857 (N_6857,N_2960,N_4547);
or U6858 (N_6858,N_4349,N_4735);
nor U6859 (N_6859,N_3478,N_4086);
and U6860 (N_6860,N_3165,N_4855);
or U6861 (N_6861,N_4784,N_3710);
nand U6862 (N_6862,N_4859,N_4594);
nor U6863 (N_6863,N_4745,N_4718);
nand U6864 (N_6864,N_3620,N_3616);
or U6865 (N_6865,N_4347,N_3507);
nand U6866 (N_6866,N_3435,N_2786);
nand U6867 (N_6867,N_3820,N_4722);
or U6868 (N_6868,N_4720,N_4474);
and U6869 (N_6869,N_3983,N_3785);
xor U6870 (N_6870,N_3319,N_3474);
xnor U6871 (N_6871,N_4405,N_4928);
nor U6872 (N_6872,N_3971,N_2836);
and U6873 (N_6873,N_4069,N_3127);
nor U6874 (N_6874,N_3362,N_4956);
nor U6875 (N_6875,N_3116,N_3956);
nand U6876 (N_6876,N_4015,N_2983);
and U6877 (N_6877,N_4672,N_3849);
xor U6878 (N_6878,N_4180,N_4286);
or U6879 (N_6879,N_4332,N_3265);
nand U6880 (N_6880,N_4104,N_3741);
or U6881 (N_6881,N_3136,N_4687);
nor U6882 (N_6882,N_3907,N_4033);
and U6883 (N_6883,N_3000,N_4993);
nand U6884 (N_6884,N_4073,N_3684);
or U6885 (N_6885,N_3903,N_4025);
and U6886 (N_6886,N_4600,N_4296);
nor U6887 (N_6887,N_3368,N_4493);
or U6888 (N_6888,N_3797,N_3079);
nand U6889 (N_6889,N_2940,N_3973);
xor U6890 (N_6890,N_2927,N_4493);
nand U6891 (N_6891,N_2744,N_3887);
and U6892 (N_6892,N_3208,N_2723);
nor U6893 (N_6893,N_3426,N_3983);
and U6894 (N_6894,N_3235,N_4037);
and U6895 (N_6895,N_3938,N_2791);
xor U6896 (N_6896,N_3726,N_2694);
xnor U6897 (N_6897,N_4571,N_4583);
and U6898 (N_6898,N_4273,N_3671);
and U6899 (N_6899,N_2679,N_2571);
nand U6900 (N_6900,N_3614,N_4143);
nand U6901 (N_6901,N_4197,N_4157);
or U6902 (N_6902,N_4130,N_4702);
nor U6903 (N_6903,N_2749,N_2815);
and U6904 (N_6904,N_4439,N_3213);
nand U6905 (N_6905,N_3749,N_4900);
xnor U6906 (N_6906,N_4158,N_4231);
nand U6907 (N_6907,N_3592,N_3241);
and U6908 (N_6908,N_3211,N_3258);
or U6909 (N_6909,N_4775,N_4208);
nor U6910 (N_6910,N_4122,N_4937);
and U6911 (N_6911,N_4944,N_3772);
and U6912 (N_6912,N_4481,N_3283);
xor U6913 (N_6913,N_4211,N_3359);
nor U6914 (N_6914,N_3195,N_2536);
nand U6915 (N_6915,N_3584,N_4474);
nor U6916 (N_6916,N_2724,N_2812);
nor U6917 (N_6917,N_3592,N_3058);
nor U6918 (N_6918,N_3151,N_3205);
and U6919 (N_6919,N_4763,N_3498);
nor U6920 (N_6920,N_3006,N_4554);
and U6921 (N_6921,N_2743,N_3946);
and U6922 (N_6922,N_4230,N_2546);
nand U6923 (N_6923,N_3393,N_4155);
nor U6924 (N_6924,N_3376,N_3369);
nor U6925 (N_6925,N_3565,N_2918);
or U6926 (N_6926,N_4496,N_4582);
and U6927 (N_6927,N_4083,N_3451);
nor U6928 (N_6928,N_4817,N_3337);
nand U6929 (N_6929,N_3812,N_4314);
or U6930 (N_6930,N_4745,N_3535);
nor U6931 (N_6931,N_3119,N_4702);
or U6932 (N_6932,N_2628,N_4364);
nand U6933 (N_6933,N_4206,N_3369);
nor U6934 (N_6934,N_4288,N_3301);
or U6935 (N_6935,N_2884,N_4123);
nor U6936 (N_6936,N_3016,N_4393);
nor U6937 (N_6937,N_3776,N_3833);
and U6938 (N_6938,N_3263,N_3791);
or U6939 (N_6939,N_2935,N_4866);
and U6940 (N_6940,N_4076,N_4094);
nor U6941 (N_6941,N_3917,N_3901);
or U6942 (N_6942,N_2863,N_3488);
nor U6943 (N_6943,N_3204,N_4723);
nor U6944 (N_6944,N_3005,N_3395);
nor U6945 (N_6945,N_4857,N_2942);
or U6946 (N_6946,N_4181,N_4809);
or U6947 (N_6947,N_4097,N_3472);
or U6948 (N_6948,N_4321,N_2996);
nand U6949 (N_6949,N_4782,N_2876);
nor U6950 (N_6950,N_4049,N_3239);
and U6951 (N_6951,N_4558,N_2505);
nand U6952 (N_6952,N_3208,N_4246);
and U6953 (N_6953,N_2639,N_4687);
or U6954 (N_6954,N_2713,N_4454);
nor U6955 (N_6955,N_2633,N_2538);
and U6956 (N_6956,N_4639,N_4048);
or U6957 (N_6957,N_4373,N_4454);
nor U6958 (N_6958,N_4486,N_4406);
nor U6959 (N_6959,N_4115,N_4166);
nor U6960 (N_6960,N_2806,N_2825);
nor U6961 (N_6961,N_3111,N_3242);
or U6962 (N_6962,N_3522,N_2799);
or U6963 (N_6963,N_4917,N_2966);
or U6964 (N_6964,N_4759,N_4001);
and U6965 (N_6965,N_4500,N_3225);
nand U6966 (N_6966,N_4389,N_4200);
and U6967 (N_6967,N_4766,N_3170);
and U6968 (N_6968,N_2752,N_4783);
and U6969 (N_6969,N_3081,N_3367);
nand U6970 (N_6970,N_3458,N_2973);
nor U6971 (N_6971,N_4093,N_4625);
and U6972 (N_6972,N_2768,N_4430);
and U6973 (N_6973,N_4972,N_3389);
xor U6974 (N_6974,N_3250,N_2589);
and U6975 (N_6975,N_3604,N_3444);
nand U6976 (N_6976,N_3674,N_4209);
nand U6977 (N_6977,N_3316,N_4114);
nor U6978 (N_6978,N_4555,N_3563);
nor U6979 (N_6979,N_3335,N_4811);
or U6980 (N_6980,N_3522,N_2854);
or U6981 (N_6981,N_3698,N_4770);
and U6982 (N_6982,N_3379,N_3747);
nor U6983 (N_6983,N_4138,N_4443);
xnor U6984 (N_6984,N_2650,N_4076);
or U6985 (N_6985,N_4855,N_4014);
or U6986 (N_6986,N_3875,N_4714);
and U6987 (N_6987,N_4807,N_3289);
and U6988 (N_6988,N_4777,N_4340);
or U6989 (N_6989,N_2634,N_3401);
xor U6990 (N_6990,N_4494,N_3409);
nand U6991 (N_6991,N_4775,N_4273);
or U6992 (N_6992,N_4035,N_3839);
nand U6993 (N_6993,N_2675,N_4006);
or U6994 (N_6994,N_3201,N_2794);
nor U6995 (N_6995,N_3666,N_4276);
nor U6996 (N_6996,N_2516,N_3794);
and U6997 (N_6997,N_4947,N_4636);
or U6998 (N_6998,N_4887,N_4928);
nand U6999 (N_6999,N_3308,N_4298);
xor U7000 (N_7000,N_2754,N_4210);
and U7001 (N_7001,N_3541,N_4202);
nand U7002 (N_7002,N_4502,N_2669);
and U7003 (N_7003,N_4708,N_3383);
or U7004 (N_7004,N_3585,N_3465);
or U7005 (N_7005,N_4925,N_4300);
or U7006 (N_7006,N_3422,N_3107);
nand U7007 (N_7007,N_4249,N_3335);
nor U7008 (N_7008,N_3255,N_4916);
nand U7009 (N_7009,N_4929,N_4885);
or U7010 (N_7010,N_4058,N_3530);
nor U7011 (N_7011,N_4127,N_4870);
xnor U7012 (N_7012,N_4300,N_4975);
or U7013 (N_7013,N_4961,N_4660);
nand U7014 (N_7014,N_4686,N_4951);
or U7015 (N_7015,N_3760,N_4252);
nand U7016 (N_7016,N_3822,N_2838);
nand U7017 (N_7017,N_4389,N_4436);
and U7018 (N_7018,N_4515,N_2893);
and U7019 (N_7019,N_4915,N_4924);
nor U7020 (N_7020,N_4376,N_4980);
and U7021 (N_7021,N_2889,N_2576);
and U7022 (N_7022,N_3363,N_4927);
and U7023 (N_7023,N_3831,N_4314);
nor U7024 (N_7024,N_3961,N_3557);
and U7025 (N_7025,N_3572,N_4218);
and U7026 (N_7026,N_3517,N_2574);
nor U7027 (N_7027,N_2859,N_4379);
and U7028 (N_7028,N_3144,N_3588);
or U7029 (N_7029,N_4105,N_3901);
xnor U7030 (N_7030,N_3237,N_3391);
and U7031 (N_7031,N_3854,N_2878);
nand U7032 (N_7032,N_4619,N_4471);
nand U7033 (N_7033,N_3873,N_4112);
and U7034 (N_7034,N_3677,N_2721);
nor U7035 (N_7035,N_2808,N_4400);
nand U7036 (N_7036,N_3336,N_3799);
or U7037 (N_7037,N_4972,N_3507);
nand U7038 (N_7038,N_4052,N_3229);
xor U7039 (N_7039,N_3269,N_4598);
and U7040 (N_7040,N_3573,N_3239);
and U7041 (N_7041,N_3660,N_3953);
or U7042 (N_7042,N_3915,N_4402);
nor U7043 (N_7043,N_2943,N_4478);
or U7044 (N_7044,N_4900,N_4173);
and U7045 (N_7045,N_3506,N_2568);
nor U7046 (N_7046,N_2574,N_4770);
nor U7047 (N_7047,N_2891,N_2829);
and U7048 (N_7048,N_4181,N_3793);
and U7049 (N_7049,N_3484,N_4387);
or U7050 (N_7050,N_4630,N_2951);
or U7051 (N_7051,N_2800,N_4599);
and U7052 (N_7052,N_2953,N_3840);
or U7053 (N_7053,N_2941,N_2601);
and U7054 (N_7054,N_3596,N_2983);
nand U7055 (N_7055,N_4065,N_2512);
and U7056 (N_7056,N_4151,N_3360);
and U7057 (N_7057,N_3178,N_3272);
xor U7058 (N_7058,N_2983,N_3003);
nor U7059 (N_7059,N_2682,N_2911);
or U7060 (N_7060,N_3385,N_4705);
or U7061 (N_7061,N_3044,N_3916);
or U7062 (N_7062,N_4475,N_3688);
nor U7063 (N_7063,N_4751,N_3106);
and U7064 (N_7064,N_3166,N_2518);
or U7065 (N_7065,N_4652,N_3378);
nor U7066 (N_7066,N_4520,N_2883);
xor U7067 (N_7067,N_2595,N_4517);
or U7068 (N_7068,N_3187,N_3004);
and U7069 (N_7069,N_3468,N_3241);
nand U7070 (N_7070,N_3347,N_3200);
or U7071 (N_7071,N_2611,N_2564);
or U7072 (N_7072,N_3853,N_4135);
nand U7073 (N_7073,N_3932,N_2784);
xor U7074 (N_7074,N_4849,N_4293);
or U7075 (N_7075,N_3739,N_3994);
nor U7076 (N_7076,N_4972,N_4587);
and U7077 (N_7077,N_3002,N_2991);
nor U7078 (N_7078,N_3391,N_4890);
or U7079 (N_7079,N_4088,N_4929);
or U7080 (N_7080,N_3788,N_4562);
nor U7081 (N_7081,N_3174,N_3339);
or U7082 (N_7082,N_3892,N_4325);
xnor U7083 (N_7083,N_2622,N_2572);
or U7084 (N_7084,N_3831,N_4785);
xnor U7085 (N_7085,N_4927,N_4612);
or U7086 (N_7086,N_4407,N_2703);
or U7087 (N_7087,N_2893,N_4791);
or U7088 (N_7088,N_2669,N_4659);
or U7089 (N_7089,N_4229,N_3535);
xor U7090 (N_7090,N_4160,N_3709);
or U7091 (N_7091,N_2924,N_2877);
nor U7092 (N_7092,N_3958,N_2691);
or U7093 (N_7093,N_3653,N_3781);
nand U7094 (N_7094,N_2908,N_3016);
nand U7095 (N_7095,N_2934,N_2812);
and U7096 (N_7096,N_4469,N_3524);
or U7097 (N_7097,N_4903,N_4278);
and U7098 (N_7098,N_3914,N_2768);
and U7099 (N_7099,N_2800,N_4726);
nand U7100 (N_7100,N_4287,N_3768);
nand U7101 (N_7101,N_3276,N_2916);
xor U7102 (N_7102,N_4159,N_3355);
nor U7103 (N_7103,N_4600,N_2726);
nor U7104 (N_7104,N_3261,N_4559);
nor U7105 (N_7105,N_2974,N_2968);
or U7106 (N_7106,N_2772,N_4473);
nand U7107 (N_7107,N_2903,N_4264);
or U7108 (N_7108,N_2516,N_3123);
and U7109 (N_7109,N_3296,N_3829);
xor U7110 (N_7110,N_3802,N_3348);
nor U7111 (N_7111,N_3330,N_3305);
nor U7112 (N_7112,N_2548,N_4177);
nor U7113 (N_7113,N_4706,N_4026);
nand U7114 (N_7114,N_4437,N_2668);
and U7115 (N_7115,N_3096,N_4119);
xnor U7116 (N_7116,N_3321,N_3092);
or U7117 (N_7117,N_3795,N_2906);
xor U7118 (N_7118,N_3799,N_2565);
xor U7119 (N_7119,N_4423,N_3336);
and U7120 (N_7120,N_4318,N_3490);
nor U7121 (N_7121,N_4845,N_3214);
nor U7122 (N_7122,N_4954,N_3620);
or U7123 (N_7123,N_3518,N_4681);
nand U7124 (N_7124,N_3986,N_3944);
or U7125 (N_7125,N_3843,N_3581);
and U7126 (N_7126,N_4062,N_3244);
nor U7127 (N_7127,N_4041,N_3269);
and U7128 (N_7128,N_3045,N_4832);
nor U7129 (N_7129,N_4353,N_4408);
or U7130 (N_7130,N_4864,N_4521);
xnor U7131 (N_7131,N_3059,N_4282);
nand U7132 (N_7132,N_3699,N_4339);
or U7133 (N_7133,N_3656,N_4134);
xor U7134 (N_7134,N_4894,N_2818);
nor U7135 (N_7135,N_4693,N_4065);
xor U7136 (N_7136,N_4176,N_4852);
and U7137 (N_7137,N_3029,N_4100);
nand U7138 (N_7138,N_2524,N_3146);
and U7139 (N_7139,N_2939,N_3255);
or U7140 (N_7140,N_4793,N_3903);
or U7141 (N_7141,N_3781,N_3244);
or U7142 (N_7142,N_3405,N_3638);
nand U7143 (N_7143,N_4223,N_2697);
and U7144 (N_7144,N_4995,N_3108);
nand U7145 (N_7145,N_3624,N_2742);
nand U7146 (N_7146,N_2987,N_3767);
and U7147 (N_7147,N_4038,N_3899);
and U7148 (N_7148,N_2853,N_2734);
xor U7149 (N_7149,N_4239,N_3237);
nand U7150 (N_7150,N_4872,N_4941);
nand U7151 (N_7151,N_2898,N_4939);
and U7152 (N_7152,N_3165,N_4007);
xor U7153 (N_7153,N_4957,N_3880);
nor U7154 (N_7154,N_4448,N_2669);
and U7155 (N_7155,N_4053,N_3938);
and U7156 (N_7156,N_3069,N_3224);
nand U7157 (N_7157,N_3953,N_3449);
nand U7158 (N_7158,N_2756,N_3820);
nor U7159 (N_7159,N_4577,N_3396);
xor U7160 (N_7160,N_4698,N_2863);
xor U7161 (N_7161,N_4739,N_3430);
nand U7162 (N_7162,N_4907,N_3476);
nor U7163 (N_7163,N_4672,N_4085);
nor U7164 (N_7164,N_3189,N_3030);
xor U7165 (N_7165,N_3787,N_3022);
xor U7166 (N_7166,N_3172,N_4184);
or U7167 (N_7167,N_3548,N_4857);
or U7168 (N_7168,N_2559,N_4737);
nor U7169 (N_7169,N_4130,N_4936);
nand U7170 (N_7170,N_4061,N_4713);
or U7171 (N_7171,N_4084,N_2544);
nor U7172 (N_7172,N_4845,N_4549);
or U7173 (N_7173,N_4679,N_2691);
or U7174 (N_7174,N_4581,N_4825);
nor U7175 (N_7175,N_4404,N_4407);
xnor U7176 (N_7176,N_3431,N_3490);
nand U7177 (N_7177,N_4101,N_2599);
and U7178 (N_7178,N_3441,N_2533);
nand U7179 (N_7179,N_3808,N_2826);
or U7180 (N_7180,N_3626,N_3851);
nor U7181 (N_7181,N_3256,N_4391);
nor U7182 (N_7182,N_3627,N_4265);
nand U7183 (N_7183,N_2676,N_2760);
nand U7184 (N_7184,N_3502,N_2641);
or U7185 (N_7185,N_2543,N_2866);
nor U7186 (N_7186,N_4787,N_4367);
or U7187 (N_7187,N_2534,N_3220);
xnor U7188 (N_7188,N_3897,N_3541);
or U7189 (N_7189,N_3081,N_4761);
and U7190 (N_7190,N_4430,N_4401);
xor U7191 (N_7191,N_3325,N_4794);
and U7192 (N_7192,N_4653,N_2914);
nor U7193 (N_7193,N_3419,N_4066);
nor U7194 (N_7194,N_4914,N_3816);
or U7195 (N_7195,N_2771,N_2785);
or U7196 (N_7196,N_3220,N_4246);
and U7197 (N_7197,N_3143,N_3314);
nor U7198 (N_7198,N_3757,N_4987);
xnor U7199 (N_7199,N_2551,N_3675);
nor U7200 (N_7200,N_3638,N_3057);
and U7201 (N_7201,N_4481,N_3667);
nor U7202 (N_7202,N_2516,N_2619);
nor U7203 (N_7203,N_3143,N_4511);
and U7204 (N_7204,N_3281,N_4671);
or U7205 (N_7205,N_2923,N_4778);
or U7206 (N_7206,N_3660,N_3810);
nand U7207 (N_7207,N_3369,N_3924);
nor U7208 (N_7208,N_3643,N_4374);
or U7209 (N_7209,N_4563,N_3582);
and U7210 (N_7210,N_4158,N_4179);
or U7211 (N_7211,N_4694,N_3490);
nand U7212 (N_7212,N_3593,N_4170);
or U7213 (N_7213,N_4152,N_2834);
or U7214 (N_7214,N_4679,N_2749);
nor U7215 (N_7215,N_2584,N_2851);
nor U7216 (N_7216,N_4811,N_4884);
nor U7217 (N_7217,N_2720,N_3513);
or U7218 (N_7218,N_2855,N_4558);
and U7219 (N_7219,N_3488,N_3894);
xnor U7220 (N_7220,N_3946,N_3813);
and U7221 (N_7221,N_4056,N_4078);
nand U7222 (N_7222,N_2998,N_2580);
or U7223 (N_7223,N_2986,N_4917);
nor U7224 (N_7224,N_2736,N_4518);
and U7225 (N_7225,N_4547,N_3554);
and U7226 (N_7226,N_2758,N_2957);
and U7227 (N_7227,N_3257,N_3482);
nand U7228 (N_7228,N_2914,N_3619);
nand U7229 (N_7229,N_2527,N_4287);
and U7230 (N_7230,N_4641,N_2613);
nor U7231 (N_7231,N_3341,N_2552);
nor U7232 (N_7232,N_3667,N_3230);
nor U7233 (N_7233,N_4366,N_2860);
or U7234 (N_7234,N_2910,N_4488);
or U7235 (N_7235,N_2758,N_3982);
or U7236 (N_7236,N_4065,N_3025);
nand U7237 (N_7237,N_4206,N_2874);
xor U7238 (N_7238,N_3747,N_3207);
xnor U7239 (N_7239,N_3589,N_3650);
and U7240 (N_7240,N_2717,N_4349);
nand U7241 (N_7241,N_3071,N_3688);
and U7242 (N_7242,N_4047,N_4705);
nor U7243 (N_7243,N_3563,N_4737);
nor U7244 (N_7244,N_3146,N_3963);
nand U7245 (N_7245,N_3324,N_2519);
or U7246 (N_7246,N_4842,N_4987);
or U7247 (N_7247,N_4593,N_2938);
or U7248 (N_7248,N_2698,N_4900);
and U7249 (N_7249,N_3317,N_4554);
or U7250 (N_7250,N_3088,N_2822);
nor U7251 (N_7251,N_2846,N_2880);
and U7252 (N_7252,N_4909,N_3819);
nand U7253 (N_7253,N_3943,N_4807);
nand U7254 (N_7254,N_4771,N_4886);
xnor U7255 (N_7255,N_3151,N_3641);
nor U7256 (N_7256,N_4824,N_3304);
or U7257 (N_7257,N_3123,N_3516);
or U7258 (N_7258,N_3040,N_3658);
nand U7259 (N_7259,N_4343,N_4372);
and U7260 (N_7260,N_3631,N_3314);
nor U7261 (N_7261,N_4895,N_4625);
nor U7262 (N_7262,N_4229,N_4901);
nor U7263 (N_7263,N_3793,N_4730);
nor U7264 (N_7264,N_2783,N_3275);
or U7265 (N_7265,N_2697,N_4144);
and U7266 (N_7266,N_4325,N_4703);
nor U7267 (N_7267,N_3142,N_4428);
and U7268 (N_7268,N_3767,N_4341);
nor U7269 (N_7269,N_4788,N_3772);
or U7270 (N_7270,N_3172,N_3293);
and U7271 (N_7271,N_3426,N_3991);
and U7272 (N_7272,N_3220,N_3367);
or U7273 (N_7273,N_4897,N_3463);
nand U7274 (N_7274,N_2732,N_4026);
nor U7275 (N_7275,N_3628,N_4599);
nand U7276 (N_7276,N_4654,N_3631);
and U7277 (N_7277,N_4863,N_2690);
nor U7278 (N_7278,N_3731,N_3265);
or U7279 (N_7279,N_4697,N_2500);
and U7280 (N_7280,N_4233,N_2888);
nand U7281 (N_7281,N_4978,N_4566);
nand U7282 (N_7282,N_4899,N_3171);
nand U7283 (N_7283,N_3087,N_3894);
and U7284 (N_7284,N_2540,N_4326);
nand U7285 (N_7285,N_2776,N_4431);
nand U7286 (N_7286,N_3659,N_3515);
and U7287 (N_7287,N_3556,N_2892);
nor U7288 (N_7288,N_3150,N_4871);
nor U7289 (N_7289,N_3954,N_4195);
and U7290 (N_7290,N_2712,N_2792);
nand U7291 (N_7291,N_3865,N_3210);
nand U7292 (N_7292,N_3160,N_4638);
nor U7293 (N_7293,N_4280,N_4479);
nor U7294 (N_7294,N_4735,N_2640);
nor U7295 (N_7295,N_4526,N_4466);
or U7296 (N_7296,N_3926,N_3182);
xnor U7297 (N_7297,N_4119,N_3116);
nor U7298 (N_7298,N_2792,N_2610);
xnor U7299 (N_7299,N_2932,N_3593);
xor U7300 (N_7300,N_2715,N_4124);
or U7301 (N_7301,N_4241,N_2803);
and U7302 (N_7302,N_3519,N_3045);
nand U7303 (N_7303,N_3297,N_4271);
and U7304 (N_7304,N_4692,N_3262);
nand U7305 (N_7305,N_4935,N_2856);
and U7306 (N_7306,N_2551,N_3316);
nand U7307 (N_7307,N_4351,N_2922);
and U7308 (N_7308,N_4096,N_2595);
nand U7309 (N_7309,N_4741,N_4350);
xnor U7310 (N_7310,N_2982,N_3030);
and U7311 (N_7311,N_3451,N_3475);
or U7312 (N_7312,N_2612,N_3199);
nand U7313 (N_7313,N_3121,N_3688);
nand U7314 (N_7314,N_3557,N_4491);
and U7315 (N_7315,N_4677,N_4439);
nand U7316 (N_7316,N_3579,N_3595);
nand U7317 (N_7317,N_3056,N_4343);
or U7318 (N_7318,N_4100,N_3004);
and U7319 (N_7319,N_4793,N_3901);
and U7320 (N_7320,N_3820,N_4730);
nand U7321 (N_7321,N_2607,N_3088);
xnor U7322 (N_7322,N_2679,N_3161);
nor U7323 (N_7323,N_2529,N_3650);
and U7324 (N_7324,N_2887,N_3588);
nand U7325 (N_7325,N_2961,N_3623);
and U7326 (N_7326,N_3659,N_3815);
nor U7327 (N_7327,N_2523,N_4262);
and U7328 (N_7328,N_4997,N_4996);
or U7329 (N_7329,N_4531,N_4746);
or U7330 (N_7330,N_3766,N_4769);
nor U7331 (N_7331,N_3835,N_2725);
nor U7332 (N_7332,N_4808,N_4625);
and U7333 (N_7333,N_2647,N_4597);
or U7334 (N_7334,N_2675,N_4419);
xnor U7335 (N_7335,N_4025,N_3795);
nand U7336 (N_7336,N_2915,N_3638);
nand U7337 (N_7337,N_3437,N_4011);
nor U7338 (N_7338,N_4452,N_4430);
xor U7339 (N_7339,N_3503,N_2996);
nor U7340 (N_7340,N_3647,N_2957);
nor U7341 (N_7341,N_4424,N_3077);
or U7342 (N_7342,N_4001,N_2953);
nand U7343 (N_7343,N_4991,N_4347);
or U7344 (N_7344,N_2939,N_4000);
nor U7345 (N_7345,N_3744,N_3259);
xor U7346 (N_7346,N_4795,N_4307);
and U7347 (N_7347,N_4306,N_3305);
nand U7348 (N_7348,N_4372,N_4168);
xnor U7349 (N_7349,N_4832,N_4200);
nor U7350 (N_7350,N_4711,N_4642);
nor U7351 (N_7351,N_4472,N_4498);
nor U7352 (N_7352,N_3246,N_4777);
or U7353 (N_7353,N_3563,N_3357);
nor U7354 (N_7354,N_4444,N_4991);
or U7355 (N_7355,N_3294,N_3886);
nand U7356 (N_7356,N_3784,N_4469);
nor U7357 (N_7357,N_3796,N_2977);
nand U7358 (N_7358,N_3042,N_4069);
nand U7359 (N_7359,N_4762,N_4188);
and U7360 (N_7360,N_4827,N_4978);
xor U7361 (N_7361,N_3248,N_3208);
and U7362 (N_7362,N_2597,N_4391);
or U7363 (N_7363,N_3327,N_4665);
or U7364 (N_7364,N_3917,N_4885);
or U7365 (N_7365,N_4082,N_4369);
or U7366 (N_7366,N_3963,N_3348);
nand U7367 (N_7367,N_4455,N_3381);
and U7368 (N_7368,N_2504,N_3859);
nor U7369 (N_7369,N_3739,N_2827);
and U7370 (N_7370,N_3083,N_4909);
nand U7371 (N_7371,N_4579,N_3597);
nor U7372 (N_7372,N_3966,N_4070);
nand U7373 (N_7373,N_4184,N_3561);
nand U7374 (N_7374,N_3520,N_3232);
nand U7375 (N_7375,N_4285,N_2728);
or U7376 (N_7376,N_4763,N_4062);
or U7377 (N_7377,N_3405,N_3689);
nor U7378 (N_7378,N_2993,N_4568);
nor U7379 (N_7379,N_3501,N_4230);
nor U7380 (N_7380,N_4060,N_4304);
nor U7381 (N_7381,N_4010,N_2647);
and U7382 (N_7382,N_3467,N_4220);
nand U7383 (N_7383,N_3137,N_4582);
nand U7384 (N_7384,N_4324,N_3466);
nand U7385 (N_7385,N_2808,N_4110);
nand U7386 (N_7386,N_4203,N_2846);
and U7387 (N_7387,N_2522,N_4467);
nand U7388 (N_7388,N_3677,N_4436);
and U7389 (N_7389,N_3949,N_4929);
and U7390 (N_7390,N_4081,N_2976);
or U7391 (N_7391,N_3574,N_4164);
and U7392 (N_7392,N_2799,N_3376);
nand U7393 (N_7393,N_4682,N_4413);
or U7394 (N_7394,N_3859,N_4536);
nor U7395 (N_7395,N_2502,N_3285);
nor U7396 (N_7396,N_3194,N_3637);
and U7397 (N_7397,N_4469,N_3209);
or U7398 (N_7398,N_2952,N_4579);
xnor U7399 (N_7399,N_4193,N_3264);
nand U7400 (N_7400,N_3510,N_3554);
nand U7401 (N_7401,N_2946,N_3318);
nand U7402 (N_7402,N_2586,N_3398);
nand U7403 (N_7403,N_3779,N_3506);
nor U7404 (N_7404,N_3612,N_3545);
and U7405 (N_7405,N_3840,N_4783);
nor U7406 (N_7406,N_4936,N_4908);
nor U7407 (N_7407,N_2792,N_4174);
xnor U7408 (N_7408,N_3790,N_3725);
xor U7409 (N_7409,N_3869,N_3247);
and U7410 (N_7410,N_2537,N_3632);
nand U7411 (N_7411,N_4961,N_2593);
nand U7412 (N_7412,N_4501,N_3035);
xnor U7413 (N_7413,N_2854,N_4433);
nor U7414 (N_7414,N_3745,N_4178);
or U7415 (N_7415,N_3657,N_3471);
nand U7416 (N_7416,N_3577,N_3975);
and U7417 (N_7417,N_4817,N_3600);
or U7418 (N_7418,N_4743,N_4404);
nand U7419 (N_7419,N_2799,N_4509);
xor U7420 (N_7420,N_3871,N_4426);
nor U7421 (N_7421,N_2587,N_2666);
nor U7422 (N_7422,N_2576,N_4656);
xnor U7423 (N_7423,N_4876,N_3968);
xnor U7424 (N_7424,N_4964,N_3161);
or U7425 (N_7425,N_3668,N_4154);
nor U7426 (N_7426,N_3375,N_2975);
and U7427 (N_7427,N_2667,N_2891);
nand U7428 (N_7428,N_3027,N_3020);
xor U7429 (N_7429,N_3649,N_3839);
or U7430 (N_7430,N_2578,N_4973);
xor U7431 (N_7431,N_2623,N_3701);
or U7432 (N_7432,N_4502,N_3648);
nand U7433 (N_7433,N_2752,N_3335);
and U7434 (N_7434,N_4045,N_4588);
nand U7435 (N_7435,N_3227,N_4077);
and U7436 (N_7436,N_3038,N_4232);
or U7437 (N_7437,N_4425,N_3169);
nor U7438 (N_7438,N_3640,N_4533);
and U7439 (N_7439,N_2570,N_3403);
nor U7440 (N_7440,N_4574,N_4438);
nand U7441 (N_7441,N_4134,N_2649);
nand U7442 (N_7442,N_3126,N_3687);
nand U7443 (N_7443,N_2762,N_4671);
nor U7444 (N_7444,N_4274,N_3914);
nor U7445 (N_7445,N_3794,N_4060);
or U7446 (N_7446,N_3026,N_3839);
or U7447 (N_7447,N_2865,N_2872);
nand U7448 (N_7448,N_2730,N_4734);
nor U7449 (N_7449,N_2788,N_4795);
xnor U7450 (N_7450,N_4551,N_4498);
nor U7451 (N_7451,N_4120,N_4274);
nor U7452 (N_7452,N_4177,N_3636);
and U7453 (N_7453,N_3338,N_4144);
nor U7454 (N_7454,N_3600,N_3347);
nor U7455 (N_7455,N_3547,N_4807);
nor U7456 (N_7456,N_3824,N_2632);
nand U7457 (N_7457,N_3612,N_3033);
or U7458 (N_7458,N_4540,N_3809);
or U7459 (N_7459,N_3413,N_4789);
nor U7460 (N_7460,N_4489,N_4896);
nand U7461 (N_7461,N_4022,N_4273);
or U7462 (N_7462,N_4868,N_3652);
xnor U7463 (N_7463,N_4058,N_2703);
or U7464 (N_7464,N_2841,N_2817);
xor U7465 (N_7465,N_4240,N_3280);
xor U7466 (N_7466,N_4077,N_4541);
and U7467 (N_7467,N_3759,N_3207);
or U7468 (N_7468,N_4590,N_3024);
or U7469 (N_7469,N_3056,N_2948);
nor U7470 (N_7470,N_2585,N_4105);
or U7471 (N_7471,N_4755,N_3917);
or U7472 (N_7472,N_4444,N_2922);
or U7473 (N_7473,N_4680,N_2851);
xnor U7474 (N_7474,N_3603,N_2760);
nor U7475 (N_7475,N_4354,N_3258);
and U7476 (N_7476,N_3368,N_4469);
xor U7477 (N_7477,N_3558,N_3070);
or U7478 (N_7478,N_2573,N_4944);
and U7479 (N_7479,N_4213,N_3965);
nand U7480 (N_7480,N_2595,N_4539);
nor U7481 (N_7481,N_4261,N_2787);
nor U7482 (N_7482,N_4858,N_4691);
nand U7483 (N_7483,N_3413,N_3638);
nor U7484 (N_7484,N_4742,N_4042);
xor U7485 (N_7485,N_3478,N_4087);
xnor U7486 (N_7486,N_3451,N_3264);
nand U7487 (N_7487,N_3535,N_4372);
nand U7488 (N_7488,N_4549,N_4046);
nand U7489 (N_7489,N_2598,N_3298);
nand U7490 (N_7490,N_3577,N_4114);
nand U7491 (N_7491,N_4558,N_3908);
nand U7492 (N_7492,N_3268,N_3938);
nand U7493 (N_7493,N_4413,N_4038);
nand U7494 (N_7494,N_4907,N_3211);
nand U7495 (N_7495,N_3997,N_4628);
nand U7496 (N_7496,N_4823,N_2540);
nor U7497 (N_7497,N_2829,N_2894);
nor U7498 (N_7498,N_3576,N_4410);
nor U7499 (N_7499,N_4039,N_4079);
nand U7500 (N_7500,N_7485,N_5150);
and U7501 (N_7501,N_6364,N_6172);
and U7502 (N_7502,N_6730,N_7303);
nor U7503 (N_7503,N_6972,N_5868);
or U7504 (N_7504,N_5862,N_6568);
or U7505 (N_7505,N_6991,N_7041);
and U7506 (N_7506,N_5446,N_6072);
nand U7507 (N_7507,N_7146,N_7169);
nor U7508 (N_7508,N_6235,N_6354);
and U7509 (N_7509,N_5962,N_5182);
nand U7510 (N_7510,N_5222,N_6748);
nand U7511 (N_7511,N_5145,N_6629);
nand U7512 (N_7512,N_6017,N_6092);
nand U7513 (N_7513,N_7015,N_5662);
nand U7514 (N_7514,N_6604,N_7334);
nor U7515 (N_7515,N_7240,N_6382);
nor U7516 (N_7516,N_5611,N_5740);
nor U7517 (N_7517,N_5510,N_6804);
or U7518 (N_7518,N_7217,N_6065);
and U7519 (N_7519,N_6646,N_5299);
and U7520 (N_7520,N_7032,N_5249);
or U7521 (N_7521,N_6101,N_5792);
nor U7522 (N_7522,N_5169,N_6241);
nor U7523 (N_7523,N_7267,N_6381);
or U7524 (N_7524,N_6598,N_5896);
xnor U7525 (N_7525,N_6011,N_6914);
nand U7526 (N_7526,N_5618,N_5649);
nor U7527 (N_7527,N_7079,N_6412);
or U7528 (N_7528,N_5642,N_5289);
nand U7529 (N_7529,N_6705,N_5058);
nor U7530 (N_7530,N_7155,N_5282);
nor U7531 (N_7531,N_6290,N_5790);
or U7532 (N_7532,N_7036,N_5276);
or U7533 (N_7533,N_6607,N_6649);
or U7534 (N_7534,N_5551,N_6619);
xor U7535 (N_7535,N_6859,N_7000);
nand U7536 (N_7536,N_5805,N_7098);
nor U7537 (N_7537,N_5221,N_6137);
nor U7538 (N_7538,N_7450,N_7219);
nor U7539 (N_7539,N_6325,N_6460);
or U7540 (N_7540,N_5542,N_5853);
xnor U7541 (N_7541,N_5309,N_6409);
nand U7542 (N_7542,N_7130,N_7149);
or U7543 (N_7543,N_6784,N_6008);
nand U7544 (N_7544,N_7387,N_6181);
nand U7545 (N_7545,N_5917,N_5823);
and U7546 (N_7546,N_6739,N_5354);
or U7547 (N_7547,N_5831,N_5779);
or U7548 (N_7548,N_5134,N_5116);
and U7549 (N_7549,N_5483,N_5413);
or U7550 (N_7550,N_6342,N_6959);
xnor U7551 (N_7551,N_6756,N_6677);
and U7552 (N_7552,N_5704,N_5439);
or U7553 (N_7553,N_7423,N_5188);
and U7554 (N_7554,N_5357,N_5328);
or U7555 (N_7555,N_6741,N_6673);
nand U7556 (N_7556,N_6868,N_5065);
nand U7557 (N_7557,N_7412,N_5803);
or U7558 (N_7558,N_5969,N_6845);
xnor U7559 (N_7559,N_7115,N_6340);
nor U7560 (N_7560,N_5938,N_5695);
or U7561 (N_7561,N_6519,N_6550);
and U7562 (N_7562,N_6347,N_5488);
nand U7563 (N_7563,N_6171,N_6527);
nand U7564 (N_7564,N_5055,N_7396);
and U7565 (N_7565,N_6539,N_5898);
nand U7566 (N_7566,N_5633,N_5748);
xor U7567 (N_7567,N_7243,N_7173);
and U7568 (N_7568,N_5869,N_6997);
nor U7569 (N_7569,N_7494,N_5669);
nor U7570 (N_7570,N_6714,N_5858);
nor U7571 (N_7571,N_7145,N_6166);
nor U7572 (N_7572,N_5246,N_7301);
or U7573 (N_7573,N_5521,N_5397);
and U7574 (N_7574,N_5172,N_6202);
xnor U7575 (N_7575,N_5423,N_6144);
nor U7576 (N_7576,N_5772,N_6436);
nor U7577 (N_7577,N_5720,N_6272);
xor U7578 (N_7578,N_5924,N_6559);
nor U7579 (N_7579,N_6350,N_7164);
or U7580 (N_7580,N_6599,N_6835);
or U7581 (N_7581,N_6168,N_6492);
nor U7582 (N_7582,N_5122,N_5300);
nor U7583 (N_7583,N_6689,N_6471);
xnor U7584 (N_7584,N_6526,N_6146);
and U7585 (N_7585,N_7213,N_6803);
and U7586 (N_7586,N_6476,N_6555);
nand U7587 (N_7587,N_6333,N_7255);
nor U7588 (N_7588,N_5504,N_5850);
nor U7589 (N_7589,N_6992,N_6737);
nor U7590 (N_7590,N_7109,N_6267);
nand U7591 (N_7591,N_7347,N_6895);
or U7592 (N_7592,N_5900,N_6205);
or U7593 (N_7593,N_5030,N_5495);
nand U7594 (N_7594,N_7226,N_6262);
nor U7595 (N_7595,N_5902,N_6229);
or U7596 (N_7596,N_5247,N_5893);
nand U7597 (N_7597,N_6178,N_6029);
or U7598 (N_7598,N_5255,N_6773);
nand U7599 (N_7599,N_7440,N_6004);
nand U7600 (N_7600,N_6344,N_7043);
or U7601 (N_7601,N_6779,N_5168);
and U7602 (N_7602,N_5745,N_7414);
nor U7603 (N_7603,N_6816,N_5812);
or U7604 (N_7604,N_6678,N_6002);
or U7605 (N_7605,N_7176,N_5700);
nor U7606 (N_7606,N_5787,N_6628);
or U7607 (N_7607,N_7231,N_5294);
and U7608 (N_7608,N_6653,N_6843);
and U7609 (N_7609,N_5179,N_5767);
or U7610 (N_7610,N_6668,N_6270);
and U7611 (N_7611,N_7238,N_7045);
nand U7612 (N_7612,N_6386,N_6510);
or U7613 (N_7613,N_5322,N_6059);
xor U7614 (N_7614,N_5925,N_5444);
and U7615 (N_7615,N_6259,N_5112);
and U7616 (N_7616,N_7214,N_6185);
nand U7617 (N_7617,N_7163,N_6194);
nand U7618 (N_7618,N_6952,N_7478);
or U7619 (N_7619,N_6223,N_5913);
nor U7620 (N_7620,N_5307,N_6359);
nand U7621 (N_7621,N_6749,N_6026);
nand U7622 (N_7622,N_6892,N_5399);
and U7623 (N_7623,N_6341,N_5971);
or U7624 (N_7624,N_5760,N_6005);
and U7625 (N_7625,N_6439,N_6658);
and U7626 (N_7626,N_7187,N_7351);
and U7627 (N_7627,N_6044,N_5911);
or U7628 (N_7628,N_7422,N_6231);
or U7629 (N_7629,N_5127,N_7257);
nand U7630 (N_7630,N_7418,N_5073);
or U7631 (N_7631,N_6230,N_5212);
nor U7632 (N_7632,N_6378,N_6841);
or U7633 (N_7633,N_6879,N_5470);
nor U7634 (N_7634,N_6617,N_6138);
nor U7635 (N_7635,N_6289,N_7196);
xnor U7636 (N_7636,N_7331,N_6576);
xnor U7637 (N_7637,N_7181,N_7336);
nand U7638 (N_7638,N_7017,N_7209);
xnor U7639 (N_7639,N_6732,N_5880);
nor U7640 (N_7640,N_5810,N_5454);
nor U7641 (N_7641,N_6545,N_6942);
nand U7642 (N_7642,N_6414,N_6544);
and U7643 (N_7643,N_6083,N_6516);
nor U7644 (N_7644,N_5199,N_5284);
and U7645 (N_7645,N_6441,N_6571);
nand U7646 (N_7646,N_5340,N_5332);
nor U7647 (N_7647,N_6495,N_5987);
nand U7648 (N_7648,N_7216,N_5820);
and U7649 (N_7649,N_6746,N_6664);
xor U7650 (N_7650,N_6077,N_5614);
and U7651 (N_7651,N_7042,N_5487);
nand U7652 (N_7652,N_5164,N_6045);
nand U7653 (N_7653,N_5106,N_5093);
nor U7654 (N_7654,N_6034,N_6219);
or U7655 (N_7655,N_5100,N_6463);
nor U7656 (N_7656,N_5944,N_5125);
nand U7657 (N_7657,N_7237,N_5796);
nor U7658 (N_7658,N_5665,N_6853);
and U7659 (N_7659,N_6442,N_5102);
and U7660 (N_7660,N_6225,N_6049);
or U7661 (N_7661,N_7111,N_5682);
nand U7662 (N_7662,N_6303,N_6100);
nor U7663 (N_7663,N_6778,N_7378);
nor U7664 (N_7664,N_5866,N_5427);
and U7665 (N_7665,N_5584,N_6175);
nand U7666 (N_7666,N_5142,N_5531);
or U7667 (N_7667,N_7279,N_5697);
and U7668 (N_7668,N_5825,N_6943);
nand U7669 (N_7669,N_5280,N_7479);
or U7670 (N_7670,N_6304,N_5634);
or U7671 (N_7671,N_5723,N_5918);
or U7672 (N_7672,N_6884,N_5729);
nand U7673 (N_7673,N_5652,N_7224);
and U7674 (N_7674,N_7053,N_6679);
xnor U7675 (N_7675,N_7370,N_6661);
or U7676 (N_7676,N_7135,N_5457);
nand U7677 (N_7677,N_6575,N_6372);
nand U7678 (N_7678,N_6944,N_5063);
nand U7679 (N_7679,N_6722,N_6834);
nand U7680 (N_7680,N_6478,N_6917);
or U7681 (N_7681,N_5020,N_6925);
nor U7682 (N_7682,N_6659,N_6594);
nand U7683 (N_7683,N_5845,N_6159);
and U7684 (N_7684,N_5956,N_5851);
or U7685 (N_7685,N_5104,N_5109);
or U7686 (N_7686,N_6240,N_7296);
and U7687 (N_7687,N_5327,N_6709);
or U7688 (N_7688,N_5391,N_6880);
nand U7689 (N_7689,N_5726,N_6491);
and U7690 (N_7690,N_7110,N_5358);
and U7691 (N_7691,N_5534,N_5148);
nand U7692 (N_7692,N_6973,N_6529);
and U7693 (N_7693,N_5854,N_7496);
nand U7694 (N_7694,N_7085,N_5241);
nor U7695 (N_7695,N_6217,N_6208);
xnor U7696 (N_7696,N_5054,N_5032);
or U7697 (N_7697,N_7291,N_5517);
nor U7698 (N_7698,N_7476,N_5429);
nor U7699 (N_7699,N_5067,N_7095);
and U7700 (N_7700,N_5217,N_6788);
nand U7701 (N_7701,N_5691,N_6695);
nand U7702 (N_7702,N_5107,N_6811);
nand U7703 (N_7703,N_7184,N_5573);
nand U7704 (N_7704,N_5047,N_5979);
or U7705 (N_7705,N_7200,N_5556);
or U7706 (N_7706,N_6553,N_5506);
nand U7707 (N_7707,N_7082,N_5929);
nand U7708 (N_7708,N_5747,N_5350);
and U7709 (N_7709,N_7443,N_5958);
and U7710 (N_7710,N_6766,N_6384);
nand U7711 (N_7711,N_5609,N_5046);
or U7712 (N_7712,N_5383,N_5785);
or U7713 (N_7713,N_6875,N_6954);
or U7714 (N_7714,N_5136,N_5033);
or U7715 (N_7715,N_6872,N_6085);
xnor U7716 (N_7716,N_5751,N_6164);
or U7717 (N_7717,N_6213,N_6031);
xnor U7718 (N_7718,N_6762,N_7484);
or U7719 (N_7719,N_7339,N_7268);
nand U7720 (N_7720,N_5507,N_7461);
and U7721 (N_7721,N_6156,N_6951);
nor U7722 (N_7722,N_7261,N_5597);
nand U7723 (N_7723,N_5066,N_6252);
and U7724 (N_7724,N_7349,N_7259);
and U7725 (N_7725,N_5782,N_5064);
and U7726 (N_7726,N_7371,N_7124);
nor U7727 (N_7727,N_6735,N_6353);
xor U7728 (N_7728,N_6455,N_5090);
nor U7729 (N_7729,N_6095,N_6949);
nand U7730 (N_7730,N_7070,N_6306);
nand U7731 (N_7731,N_5764,N_5114);
xor U7732 (N_7732,N_6790,N_6484);
and U7733 (N_7733,N_5436,N_6302);
nor U7734 (N_7734,N_6383,N_6932);
and U7735 (N_7735,N_6890,N_7253);
nor U7736 (N_7736,N_5472,N_5263);
or U7737 (N_7737,N_6919,N_6697);
xor U7738 (N_7738,N_5202,N_5629);
xor U7739 (N_7739,N_5888,N_7235);
and U7740 (N_7740,N_5897,N_6346);
and U7741 (N_7741,N_5267,N_5475);
or U7742 (N_7742,N_6321,N_7493);
nor U7743 (N_7743,N_6182,N_5215);
or U7744 (N_7744,N_7368,N_5563);
or U7745 (N_7745,N_7442,N_5777);
or U7746 (N_7746,N_7193,N_5335);
and U7747 (N_7747,N_7024,N_7080);
nand U7748 (N_7748,N_6468,N_5494);
nor U7749 (N_7749,N_6195,N_6975);
xnor U7750 (N_7750,N_5197,N_6694);
nand U7751 (N_7751,N_6787,N_6525);
or U7752 (N_7752,N_5103,N_6582);
and U7753 (N_7753,N_5019,N_5621);
nor U7754 (N_7754,N_6538,N_5570);
nor U7755 (N_7755,N_5909,N_5497);
and U7756 (N_7756,N_5166,N_6007);
nand U7757 (N_7757,N_6087,N_7067);
xnor U7758 (N_7758,N_7114,N_6196);
nand U7759 (N_7759,N_6109,N_5832);
nand U7760 (N_7760,N_6983,N_5044);
and U7761 (N_7761,N_6127,N_5762);
and U7762 (N_7762,N_6933,N_6977);
nor U7763 (N_7763,N_6871,N_7282);
or U7764 (N_7764,N_5149,N_6842);
and U7765 (N_7765,N_5668,N_5157);
xnor U7766 (N_7766,N_6815,N_6475);
and U7767 (N_7767,N_6636,N_6066);
or U7768 (N_7768,N_6729,N_6897);
and U7769 (N_7769,N_5227,N_6315);
nor U7770 (N_7770,N_5001,N_6685);
nor U7771 (N_7771,N_7435,N_6502);
nor U7772 (N_7772,N_5187,N_5945);
and U7773 (N_7773,N_7160,N_6686);
nand U7774 (N_7774,N_5342,N_6578);
nand U7775 (N_7775,N_5752,N_6363);
and U7776 (N_7776,N_5694,N_6906);
nand U7777 (N_7777,N_7300,N_5130);
or U7778 (N_7778,N_5592,N_5496);
and U7779 (N_7779,N_5941,N_6391);
nand U7780 (N_7780,N_6615,N_5778);
nor U7781 (N_7781,N_5052,N_5463);
nor U7782 (N_7782,N_6512,N_5422);
and U7783 (N_7783,N_5028,N_7254);
or U7784 (N_7784,N_6084,N_6750);
and U7785 (N_7785,N_6404,N_5876);
nand U7786 (N_7786,N_5844,N_5452);
nand U7787 (N_7787,N_6312,N_6624);
xnor U7788 (N_7788,N_7436,N_7452);
xor U7789 (N_7789,N_6752,N_6323);
nand U7790 (N_7790,N_6692,N_6448);
or U7791 (N_7791,N_5657,N_6496);
or U7792 (N_7792,N_5798,N_7195);
nor U7793 (N_7793,N_7104,N_7491);
nand U7794 (N_7794,N_6591,N_6405);
and U7795 (N_7795,N_5206,N_6081);
nand U7796 (N_7796,N_7381,N_6542);
or U7797 (N_7797,N_5549,N_6712);
or U7798 (N_7798,N_5829,N_7121);
or U7799 (N_7799,N_5467,N_5012);
and U7800 (N_7800,N_6129,N_5140);
or U7801 (N_7801,N_5425,N_7180);
nor U7802 (N_7802,N_5639,N_5959);
or U7803 (N_7803,N_6776,N_5339);
nand U7804 (N_7804,N_7358,N_5389);
nand U7805 (N_7805,N_6785,N_6211);
nand U7806 (N_7806,N_5250,N_5324);
xnor U7807 (N_7807,N_5786,N_5297);
or U7808 (N_7808,N_5899,N_7192);
xor U7809 (N_7809,N_6314,N_5827);
nor U7810 (N_7810,N_7321,N_7260);
and U7811 (N_7811,N_7275,N_6560);
or U7812 (N_7812,N_7210,N_6535);
nand U7813 (N_7813,N_6913,N_6939);
nor U7814 (N_7814,N_5161,N_6740);
nor U7815 (N_7815,N_5569,N_6543);
or U7816 (N_7816,N_6062,N_5298);
and U7817 (N_7817,N_6188,N_6955);
nand U7818 (N_7818,N_6206,N_6585);
or U7819 (N_7819,N_6487,N_6430);
xor U7820 (N_7820,N_7475,N_5443);
nand U7821 (N_7821,N_6822,N_5320);
nand U7822 (N_7822,N_6513,N_5572);
or U7823 (N_7823,N_5595,N_5821);
nor U7824 (N_7824,N_6308,N_5582);
nor U7825 (N_7825,N_6108,N_6296);
or U7826 (N_7826,N_7143,N_5338);
nor U7827 (N_7827,N_5501,N_6033);
and U7828 (N_7828,N_7128,N_6387);
and U7829 (N_7829,N_5373,N_6173);
and U7830 (N_7830,N_7140,N_5826);
and U7831 (N_7831,N_5388,N_6866);
xor U7832 (N_7832,N_5756,N_5017);
or U7833 (N_7833,N_5291,N_6286);
or U7834 (N_7834,N_7166,N_6415);
and U7835 (N_7835,N_5603,N_6132);
nor U7836 (N_7836,N_7362,N_6549);
or U7837 (N_7837,N_6258,N_6073);
nand U7838 (N_7838,N_6050,N_6298);
xor U7839 (N_7839,N_6820,N_6375);
nor U7840 (N_7840,N_6078,N_5990);
nor U7841 (N_7841,N_5421,N_6183);
and U7842 (N_7842,N_5456,N_6963);
and U7843 (N_7843,N_6279,N_6288);
nand U7844 (N_7844,N_6757,N_5718);
or U7845 (N_7845,N_6751,N_7252);
and U7846 (N_7846,N_5362,N_6901);
or U7847 (N_7847,N_7465,N_5311);
or U7848 (N_7848,N_6671,N_6855);
and U7849 (N_7849,N_5605,N_6893);
nor U7850 (N_7850,N_6810,N_7059);
xnor U7851 (N_7851,N_5770,N_7338);
nand U7852 (N_7852,N_7401,N_5469);
and U7853 (N_7853,N_5892,N_7474);
xor U7854 (N_7854,N_5374,N_7281);
nand U7855 (N_7855,N_5905,N_6889);
or U7856 (N_7856,N_5708,N_7357);
nor U7857 (N_7857,N_7174,N_5050);
nand U7858 (N_7858,N_6155,N_7467);
nor U7859 (N_7859,N_7118,N_5655);
nand U7860 (N_7860,N_5544,N_5992);
nand U7861 (N_7861,N_5260,N_5735);
and U7862 (N_7862,N_6962,N_5240);
and U7863 (N_7863,N_5673,N_6981);
or U7864 (N_7864,N_6606,N_5970);
nor U7865 (N_7865,N_5783,N_6569);
and U7866 (N_7866,N_6564,N_6858);
or U7867 (N_7867,N_6271,N_5773);
or U7868 (N_7868,N_6479,N_6165);
nand U7869 (N_7869,N_7005,N_7437);
or U7870 (N_7870,N_5021,N_6330);
xnor U7871 (N_7871,N_6522,N_5337);
nand U7872 (N_7872,N_7376,N_6422);
nor U7873 (N_7873,N_6761,N_5165);
or U7874 (N_7874,N_5855,N_5711);
or U7875 (N_7875,N_5286,N_7072);
or U7876 (N_7876,N_5701,N_6110);
or U7877 (N_7877,N_6994,N_6454);
or U7878 (N_7878,N_7352,N_6157);
or U7879 (N_7879,N_7101,N_5623);
and U7880 (N_7880,N_5094,N_5037);
and U7881 (N_7881,N_5524,N_7157);
nor U7882 (N_7882,N_7052,N_5800);
xor U7883 (N_7883,N_5190,N_7318);
and U7884 (N_7884,N_6339,N_7039);
and U7885 (N_7885,N_5589,N_6824);
and U7886 (N_7886,N_5568,N_6399);
and U7887 (N_7887,N_5937,N_5499);
nand U7888 (N_7888,N_6328,N_5465);
nand U7889 (N_7889,N_5119,N_7431);
or U7890 (N_7890,N_6934,N_5061);
and U7891 (N_7891,N_5398,N_6935);
xnor U7892 (N_7892,N_5285,N_5724);
and U7893 (N_7893,N_6300,N_7199);
nor U7894 (N_7894,N_6493,N_5755);
nor U7895 (N_7895,N_5750,N_6310);
and U7896 (N_7896,N_7497,N_6417);
and U7897 (N_7897,N_6584,N_6950);
and U7898 (N_7898,N_7183,N_5194);
or U7899 (N_7899,N_7096,N_6524);
xnor U7900 (N_7900,N_6283,N_7137);
nor U7901 (N_7901,N_5600,N_6852);
xor U7902 (N_7902,N_5163,N_6242);
nand U7903 (N_7903,N_7451,N_6006);
nand U7904 (N_7904,N_7405,N_7141);
nand U7905 (N_7905,N_6427,N_5795);
nand U7906 (N_7906,N_6869,N_7092);
and U7907 (N_7907,N_6228,N_5390);
xnor U7908 (N_7908,N_6851,N_5952);
or U7909 (N_7909,N_6282,N_5181);
nor U7910 (N_7910,N_5930,N_5836);
and U7911 (N_7911,N_5980,N_6540);
and U7912 (N_7912,N_5124,N_7425);
and U7913 (N_7913,N_7159,N_5857);
nand U7914 (N_7914,N_6082,N_6216);
nand U7915 (N_7915,N_6532,N_5833);
xor U7916 (N_7916,N_5434,N_5973);
nor U7917 (N_7917,N_6079,N_5092);
nor U7918 (N_7918,N_5353,N_7463);
nand U7919 (N_7919,N_6700,N_6936);
and U7920 (N_7920,N_5624,N_5110);
or U7921 (N_7921,N_6774,N_5516);
or U7922 (N_7922,N_5403,N_7120);
nand U7923 (N_7923,N_5447,N_6091);
nor U7924 (N_7924,N_5581,N_6248);
nand U7925 (N_7925,N_5325,N_6125);
nand U7926 (N_7926,N_7011,N_6797);
nand U7927 (N_7927,N_6094,N_6051);
nand U7928 (N_7928,N_5640,N_7492);
or U7929 (N_7929,N_6433,N_6876);
or U7930 (N_7930,N_5989,N_5178);
nand U7931 (N_7931,N_7372,N_7189);
or U7932 (N_7932,N_6967,N_5293);
nor U7933 (N_7933,N_5316,N_5226);
and U7934 (N_7934,N_5437,N_5659);
or U7935 (N_7935,N_6385,N_5441);
xnor U7936 (N_7936,N_6621,N_7361);
and U7937 (N_7937,N_7023,N_5170);
and U7938 (N_7938,N_5143,N_5784);
and U7939 (N_7939,N_6902,N_5736);
and U7940 (N_7940,N_7307,N_5801);
and U7941 (N_7941,N_5912,N_7131);
and U7942 (N_7942,N_5401,N_5677);
nor U7943 (N_7943,N_6765,N_5731);
nand U7944 (N_7944,N_5995,N_6369);
nand U7945 (N_7945,N_5641,N_7020);
or U7946 (N_7946,N_6918,N_5643);
and U7947 (N_7947,N_5865,N_6266);
nor U7948 (N_7948,N_6421,N_5920);
and U7949 (N_7949,N_5926,N_6373);
nor U7950 (N_7950,N_7438,N_6048);
nor U7951 (N_7951,N_7360,N_5985);
or U7952 (N_7952,N_6704,N_5988);
nand U7953 (N_7953,N_5746,N_5686);
nor U7954 (N_7954,N_5175,N_6329);
nand U7955 (N_7955,N_7316,N_5481);
nor U7956 (N_7956,N_6970,N_5333);
or U7957 (N_7957,N_7473,N_6257);
or U7958 (N_7958,N_6656,N_5111);
and U7959 (N_7959,N_6253,N_6148);
and U7960 (N_7960,N_5018,N_5367);
nor U7961 (N_7961,N_7037,N_7126);
nand U7962 (N_7962,N_7311,N_6579);
and U7963 (N_7963,N_7292,N_6641);
and U7964 (N_7964,N_6437,N_6307);
or U7965 (N_7965,N_7133,N_7031);
nor U7966 (N_7966,N_5196,N_7054);
nand U7967 (N_7967,N_5585,N_7151);
nand U7968 (N_7968,N_6028,N_5329);
and U7969 (N_7969,N_6141,N_7147);
or U7970 (N_7970,N_5693,N_6899);
or U7971 (N_7971,N_6921,N_6207);
nand U7972 (N_7972,N_6982,N_6911);
and U7973 (N_7973,N_7286,N_6158);
nand U7974 (N_7974,N_5219,N_7211);
nor U7975 (N_7975,N_5098,N_6622);
xnor U7976 (N_7976,N_6601,N_7245);
nor U7977 (N_7977,N_6070,N_6473);
and U7978 (N_7978,N_7276,N_6812);
or U7979 (N_7979,N_5742,N_5982);
and U7980 (N_7980,N_6836,N_5996);
nand U7981 (N_7981,N_6000,N_7197);
nor U7982 (N_7982,N_6500,N_6630);
nand U7983 (N_7983,N_7434,N_5455);
xnor U7984 (N_7984,N_5953,N_5519);
or U7985 (N_7985,N_7134,N_5599);
nor U7986 (N_7986,N_5420,N_7170);
or U7987 (N_7987,N_5843,N_5071);
nor U7988 (N_7988,N_7154,N_6506);
and U7989 (N_7989,N_5056,N_5410);
xnor U7990 (N_7990,N_7326,N_5304);
or U7991 (N_7991,N_5154,N_6764);
nand U7992 (N_7992,N_5211,N_5128);
or U7993 (N_7993,N_6053,N_6801);
nor U7994 (N_7994,N_7250,N_6401);
or U7995 (N_7995,N_6226,N_7317);
and U7996 (N_7996,N_6758,N_6708);
and U7997 (N_7997,N_6126,N_7251);
or U7998 (N_7998,N_6863,N_6464);
xnor U7999 (N_7999,N_6847,N_6638);
nor U8000 (N_8000,N_5198,N_6121);
nand U8001 (N_8001,N_6191,N_5005);
xnor U8002 (N_8002,N_7029,N_6592);
and U8003 (N_8003,N_5292,N_5763);
nand U8004 (N_8004,N_6603,N_6698);
xor U8005 (N_8005,N_5159,N_7350);
nand U8006 (N_8006,N_6010,N_7393);
xor U8007 (N_8007,N_6896,N_5268);
or U8008 (N_8008,N_6016,N_7007);
nor U8009 (N_8009,N_6220,N_6361);
or U8010 (N_8010,N_6703,N_6115);
nand U8011 (N_8011,N_5552,N_5610);
xnor U8012 (N_8012,N_6509,N_5539);
or U8013 (N_8013,N_5312,N_5511);
and U8014 (N_8014,N_6488,N_7421);
nor U8015 (N_8015,N_6458,N_5036);
and U8016 (N_8016,N_5811,N_7274);
or U8017 (N_8017,N_5975,N_5264);
and U8018 (N_8018,N_5068,N_5852);
or U8019 (N_8019,N_6929,N_5998);
nor U8020 (N_8020,N_6514,N_5571);
or U8021 (N_8021,N_5394,N_6197);
nor U8022 (N_8022,N_7456,N_5356);
and U8023 (N_8023,N_6595,N_7466);
nand U8024 (N_8024,N_6222,N_5703);
nand U8025 (N_8025,N_5738,N_5318);
nand U8026 (N_8026,N_7404,N_5553);
xor U8027 (N_8027,N_5015,N_7266);
nor U8028 (N_8028,N_6998,N_5837);
and U8029 (N_8029,N_5654,N_6151);
and U8030 (N_8030,N_5433,N_6411);
nor U8031 (N_8031,N_5416,N_5493);
xor U8032 (N_8032,N_6999,N_7269);
nor U8033 (N_8033,N_5744,N_5809);
nor U8034 (N_8034,N_5698,N_5842);
or U8035 (N_8035,N_6410,N_5626);
nor U8036 (N_8036,N_6301,N_5387);
nand U8037 (N_8037,N_6581,N_6416);
or U8038 (N_8038,N_5039,N_6878);
and U8039 (N_8039,N_5408,N_6444);
and U8040 (N_8040,N_5559,N_6754);
and U8041 (N_8041,N_6986,N_6717);
nor U8042 (N_8042,N_6190,N_6446);
nand U8043 (N_8043,N_5016,N_7384);
nand U8044 (N_8044,N_5991,N_5864);
and U8045 (N_8045,N_5914,N_6681);
nand U8046 (N_8046,N_5118,N_6319);
and U8047 (N_8047,N_6837,N_5797);
or U8048 (N_8048,N_7025,N_6734);
nor U8049 (N_8049,N_6772,N_7429);
or U8050 (N_8050,N_7185,N_6832);
and U8051 (N_8051,N_5229,N_6426);
and U8052 (N_8052,N_6940,N_6965);
or U8053 (N_8053,N_5479,N_6145);
nand U8054 (N_8054,N_5070,N_6915);
nand U8055 (N_8055,N_5051,N_6844);
and U8056 (N_8056,N_5485,N_6783);
nor U8057 (N_8057,N_5806,N_5022);
and U8058 (N_8058,N_5407,N_5514);
nor U8059 (N_8059,N_6727,N_7161);
nand U8060 (N_8060,N_5346,N_6120);
nor U8061 (N_8061,N_6498,N_5722);
nor U8062 (N_8062,N_7319,N_5529);
and U8063 (N_8063,N_5473,N_6715);
nor U8064 (N_8064,N_5345,N_7062);
nand U8065 (N_8065,N_5415,N_6025);
nand U8066 (N_8066,N_5537,N_6554);
and U8067 (N_8067,N_6440,N_5617);
nand U8068 (N_8068,N_6111,N_6809);
nand U8069 (N_8069,N_6152,N_5459);
xnor U8070 (N_8070,N_6922,N_7340);
nor U8071 (N_8071,N_6104,N_5983);
nand U8072 (N_8072,N_6988,N_7264);
or U8073 (N_8073,N_6953,N_7012);
nand U8074 (N_8074,N_5791,N_7201);
nor U8075 (N_8075,N_6637,N_6117);
nor U8076 (N_8076,N_5648,N_6232);
and U8077 (N_8077,N_6987,N_5919);
nor U8078 (N_8078,N_7413,N_6472);
nor U8079 (N_8079,N_5875,N_5838);
xnor U8080 (N_8080,N_7227,N_6075);
xnor U8081 (N_8081,N_5295,N_5628);
and U8082 (N_8082,N_6721,N_5287);
or U8083 (N_8083,N_5236,N_5173);
or U8084 (N_8084,N_6254,N_6140);
nor U8085 (N_8085,N_7411,N_7086);
or U8086 (N_8086,N_5137,N_5776);
nor U8087 (N_8087,N_5461,N_6162);
or U8088 (N_8088,N_7153,N_6702);
and U8089 (N_8089,N_6494,N_5932);
or U8090 (N_8090,N_5513,N_5541);
and U8091 (N_8091,N_5262,N_5828);
xor U8092 (N_8092,N_7178,N_6826);
and U8093 (N_8093,N_5887,N_7288);
nand U8094 (N_8094,N_5231,N_6052);
nor U8095 (N_8095,N_6956,N_6212);
or U8096 (N_8096,N_5370,N_5564);
and U8097 (N_8097,N_6355,N_5619);
nor U8098 (N_8098,N_6295,N_7445);
nand U8099 (N_8099,N_6626,N_6517);
nor U8100 (N_8100,N_6908,N_7388);
or U8101 (N_8101,N_5082,N_7056);
or U8102 (N_8102,N_5527,N_6227);
or U8103 (N_8103,N_5371,N_5025);
nand U8104 (N_8104,N_7284,N_5281);
nand U8105 (N_8105,N_5788,N_6583);
nand U8106 (N_8106,N_5523,N_5808);
nand U8107 (N_8107,N_5158,N_6093);
nor U8108 (N_8108,N_7394,N_5224);
or U8109 (N_8109,N_7408,N_5238);
and U8110 (N_8110,N_5949,N_6612);
nand U8111 (N_8111,N_7094,N_6924);
xor U8112 (N_8112,N_5355,N_7353);
or U8113 (N_8113,N_7258,N_5817);
or U8114 (N_8114,N_5484,N_5663);
nand U8115 (N_8115,N_6640,N_5426);
xor U8116 (N_8116,N_6680,N_6557);
nor U8117 (N_8117,N_5885,N_6076);
or U8118 (N_8118,N_6558,N_6593);
nand U8119 (N_8119,N_7295,N_5027);
nor U8120 (N_8120,N_5895,N_7458);
and U8121 (N_8121,N_7248,N_7483);
xor U8122 (N_8122,N_6759,N_6068);
nor U8123 (N_8123,N_5233,N_7047);
and U8124 (N_8124,N_5879,N_6423);
or U8125 (N_8125,N_6398,N_5505);
xnor U8126 (N_8126,N_5352,N_7191);
nor U8127 (N_8127,N_5840,N_6923);
nand U8128 (N_8128,N_5678,N_5491);
xnor U8129 (N_8129,N_5580,N_6311);
nor U8130 (N_8130,N_6177,N_5176);
nand U8131 (N_8131,N_5315,N_6397);
nand U8132 (N_8132,N_6377,N_5947);
xnor U8133 (N_8133,N_5566,N_5386);
or U8134 (N_8134,N_7165,N_6941);
nand U8135 (N_8135,N_5993,N_5442);
nor U8136 (N_8136,N_5144,N_5059);
nor U8137 (N_8137,N_5977,N_5203);
and U8138 (N_8138,N_7385,N_6018);
nor U8139 (N_8139,N_7335,N_6978);
and U8140 (N_8140,N_7367,N_6828);
nand U8141 (N_8141,N_6037,N_6838);
nand U8142 (N_8142,N_5664,N_5360);
and U8143 (N_8143,N_6930,N_6881);
and U8144 (N_8144,N_5476,N_6660);
or U8145 (N_8145,N_5305,N_6886);
nand U8146 (N_8146,N_6023,N_6780);
and U8147 (N_8147,N_5223,N_7490);
nand U8148 (N_8148,N_6003,N_6523);
or U8149 (N_8149,N_7323,N_7262);
or U8150 (N_8150,N_5135,N_5725);
xor U8151 (N_8151,N_7369,N_5769);
or U8152 (N_8152,N_6352,N_6210);
and U8153 (N_8153,N_7002,N_5536);
or U8154 (N_8154,N_6666,N_7205);
and U8155 (N_8155,N_7232,N_5156);
or U8156 (N_8156,N_6957,N_7172);
nand U8157 (N_8157,N_7499,N_7003);
xnor U8158 (N_8158,N_7299,N_5999);
and U8159 (N_8159,N_6728,N_5847);
nor U8160 (N_8160,N_5627,N_6107);
and U8161 (N_8161,N_6324,N_5954);
nor U8162 (N_8162,N_7363,N_6818);
xnor U8163 (N_8163,N_7327,N_6064);
xnor U8164 (N_8164,N_5319,N_6046);
nor U8165 (N_8165,N_5368,N_7182);
and U8166 (N_8166,N_5209,N_6277);
nor U8167 (N_8167,N_5578,N_6467);
nor U8168 (N_8168,N_5586,N_6418);
nor U8169 (N_8169,N_5321,N_6388);
and U8170 (N_8170,N_5743,N_5269);
nor U8171 (N_8171,N_5123,N_6635);
and U8172 (N_8172,N_7481,N_5780);
nor U8173 (N_8173,N_7239,N_6652);
or U8174 (N_8174,N_6099,N_5372);
or U8175 (N_8175,N_5377,N_6613);
or U8176 (N_8176,N_7298,N_6407);
nor U8177 (N_8177,N_6133,N_5928);
and U8178 (N_8178,N_5859,N_6795);
and U8179 (N_8179,N_5430,N_5688);
nand U8180 (N_8180,N_5602,N_6833);
xnor U8181 (N_8181,N_7087,N_5085);
nand U8182 (N_8182,N_7188,N_5195);
nor U8183 (N_8183,N_5804,N_5038);
and U8184 (N_8184,N_7018,N_5976);
or U8185 (N_8185,N_5771,N_6284);
nor U8186 (N_8186,N_5060,N_6483);
and U8187 (N_8187,N_7342,N_6632);
or U8188 (N_8188,N_5008,N_6305);
or U8189 (N_8189,N_6477,N_5874);
nor U8190 (N_8190,N_5901,N_6588);
nand U8191 (N_8191,N_7150,N_6536);
and U8192 (N_8192,N_7265,N_6521);
nor U8193 (N_8193,N_5789,N_5579);
xor U8194 (N_8194,N_6131,N_5348);
nor U8195 (N_8195,N_5873,N_6293);
xor U8196 (N_8196,N_5482,N_5084);
nor U8197 (N_8197,N_6395,N_6394);
or U8198 (N_8198,N_5449,N_7099);
and U8199 (N_8199,N_5344,N_6547);
and U8200 (N_8200,N_6234,N_6877);
nor U8201 (N_8201,N_7343,N_7069);
nand U8202 (N_8202,N_6103,N_6431);
nor U8203 (N_8203,N_5910,N_6291);
or U8204 (N_8204,N_5967,N_5313);
and U8205 (N_8205,N_7345,N_5613);
xnor U8206 (N_8206,N_6596,N_6747);
or U8207 (N_8207,N_5822,N_5978);
or U8208 (N_8208,N_6041,N_6995);
xor U8209 (N_8209,N_5753,N_5428);
and U8210 (N_8210,N_7022,N_6074);
nand U8211 (N_8211,N_5923,N_5004);
nand U8212 (N_8212,N_7065,N_5675);
nand U8213 (N_8213,N_5512,N_5968);
or U8214 (N_8214,N_6123,N_5132);
nor U8215 (N_8215,N_5207,N_6602);
or U8216 (N_8216,N_5560,N_5278);
nor U8217 (N_8217,N_6657,N_5948);
or U8218 (N_8218,N_6276,N_5296);
or U8219 (N_8219,N_5676,N_6926);
and U8220 (N_8220,N_6675,N_5934);
and U8221 (N_8221,N_6327,N_7105);
nand U8222 (N_8222,N_6263,N_7294);
and U8223 (N_8223,N_6209,N_7380);
and U8224 (N_8224,N_6781,N_5080);
or U8225 (N_8225,N_5121,N_6199);
nand U8226 (N_8226,N_5528,N_6489);
or U8227 (N_8227,N_5251,N_6938);
and U8228 (N_8228,N_5435,N_6256);
nor U8229 (N_8229,N_6552,N_7459);
nor U8230 (N_8230,N_5076,N_7097);
nand U8231 (N_8231,N_7379,N_6112);
or U8232 (N_8232,N_5860,N_5734);
and U8233 (N_8233,N_6281,N_6743);
or U8234 (N_8234,N_6193,N_5147);
nor U8235 (N_8235,N_5414,N_5867);
nor U8236 (N_8236,N_5331,N_7297);
xor U8237 (N_8237,N_6450,N_6910);
or U8238 (N_8238,N_5871,N_5069);
nand U8239 (N_8239,N_6767,N_5088);
and U8240 (N_8240,N_7322,N_7430);
nand U8241 (N_8241,N_7278,N_6245);
or U8242 (N_8242,N_6793,N_6170);
or U8243 (N_8243,N_7194,N_6060);
xnor U8244 (N_8244,N_5235,N_5933);
or U8245 (N_8245,N_6102,N_6586);
or U8246 (N_8246,N_6069,N_7472);
or U8247 (N_8247,N_6763,N_5942);
nor U8248 (N_8248,N_6214,N_6351);
and U8249 (N_8249,N_6204,N_5557);
and U8250 (N_8250,N_6297,N_6665);
or U8251 (N_8251,N_5160,N_7312);
nor U8252 (N_8252,N_5087,N_6299);
or U8253 (N_8253,N_6937,N_5672);
or U8254 (N_8254,N_6813,N_5186);
or U8255 (N_8255,N_7049,N_6246);
nor U8256 (N_8256,N_6334,N_6160);
or U8257 (N_8257,N_7088,N_6831);
nand U8258 (N_8258,N_7495,N_7488);
nand U8259 (N_8259,N_5041,N_5048);
or U8260 (N_8260,N_7091,N_6885);
nor U8261 (N_8261,N_7427,N_6968);
nor U8262 (N_8262,N_6707,N_6888);
or U8263 (N_8263,N_5396,N_5275);
nand U8264 (N_8264,N_5385,N_5670);
nand U8265 (N_8265,N_6742,N_6768);
and U8266 (N_8266,N_7230,N_5042);
or U8267 (N_8267,N_7241,N_5716);
nor U8268 (N_8268,N_6701,N_5220);
and U8269 (N_8269,N_6782,N_6623);
or U8270 (N_8270,N_7089,N_7480);
or U8271 (N_8271,N_6233,N_6777);
nand U8272 (N_8272,N_7075,N_7051);
nor U8273 (N_8273,N_5758,N_6800);
or U8274 (N_8274,N_6775,N_7453);
or U8275 (N_8275,N_5561,N_5303);
xnor U8276 (N_8276,N_6520,N_6186);
nand U8277 (N_8277,N_5903,N_5526);
nor U8278 (N_8278,N_6839,N_6533);
xor U8279 (N_8279,N_5915,N_6503);
nand U8280 (N_8280,N_6786,N_5115);
nand U8281 (N_8281,N_6731,N_5351);
nor U8282 (N_8282,N_5632,N_5814);
nand U8283 (N_8283,N_7035,N_7179);
xnor U8284 (N_8284,N_7407,N_7138);
nand U8285 (N_8285,N_6589,N_7486);
and U8286 (N_8286,N_6755,N_7050);
or U8287 (N_8287,N_6979,N_5105);
nor U8288 (N_8288,N_5245,N_5818);
and U8289 (N_8289,N_6379,N_6447);
or U8290 (N_8290,N_6990,N_6147);
nand U8291 (N_8291,N_7289,N_7365);
or U8292 (N_8292,N_7489,N_6898);
and U8293 (N_8293,N_5471,N_5878);
nor U8294 (N_8294,N_5411,N_6861);
nand U8295 (N_8295,N_5710,N_7014);
and U8296 (N_8296,N_5650,N_7391);
or U8297 (N_8297,N_5432,N_6805);
nand U8298 (N_8298,N_6280,N_6055);
and U8299 (N_8299,N_6650,N_7247);
nor U8300 (N_8300,N_7078,N_5237);
and U8301 (N_8301,N_6699,N_5737);
or U8302 (N_8302,N_6821,N_5393);
and U8303 (N_8303,N_6452,N_6865);
and U8304 (N_8304,N_5886,N_7175);
nor U8305 (N_8305,N_5438,N_5702);
nor U8306 (N_8306,N_7457,N_7468);
nand U8307 (N_8307,N_5192,N_5646);
or U8308 (N_8308,N_6806,N_5205);
nor U8309 (N_8309,N_5644,N_5213);
or U8310 (N_8310,N_5713,N_7113);
nand U8311 (N_8311,N_7030,N_5117);
nor U8312 (N_8312,N_6318,N_6501);
nand U8313 (N_8313,N_5667,N_5014);
or U8314 (N_8314,N_6643,N_6336);
or U8315 (N_8315,N_6163,N_7280);
nand U8316 (N_8316,N_7354,N_6322);
or U8317 (N_8317,N_6706,N_5596);
nor U8318 (N_8318,N_6976,N_6142);
nor U8319 (N_8319,N_6287,N_6180);
and U8320 (N_8320,N_6054,N_5376);
nand U8321 (N_8321,N_5986,N_6425);
nand U8322 (N_8322,N_5392,N_5841);
and U8323 (N_8323,N_7222,N_6798);
xnor U8324 (N_8324,N_5007,N_5216);
and U8325 (N_8325,N_5908,N_5606);
or U8326 (N_8326,N_5877,N_7057);
nor U8327 (N_8327,N_5361,N_6791);
or U8328 (N_8328,N_7203,N_6090);
or U8329 (N_8329,N_5714,N_5464);
or U8330 (N_8330,N_7142,N_5525);
or U8331 (N_8331,N_5906,N_6113);
and U8332 (N_8332,N_5881,N_6469);
or U8333 (N_8333,N_6465,N_5412);
and U8334 (N_8334,N_7382,N_6672);
nor U8335 (N_8335,N_7198,N_6912);
and U8336 (N_8336,N_5965,N_6063);
xor U8337 (N_8337,N_6255,N_7066);
nand U8338 (N_8338,N_7008,N_7333);
nor U8339 (N_8339,N_5593,N_6366);
nand U8340 (N_8340,N_6024,N_5816);
and U8341 (N_8341,N_7324,N_5096);
nand U8342 (N_8342,N_5230,N_5802);
nor U8343 (N_8343,N_5138,N_5616);
xnor U8344 (N_8344,N_7400,N_5266);
or U8345 (N_8345,N_7444,N_5508);
nand U8346 (N_8346,N_7462,N_5002);
nand U8347 (N_8347,N_5598,N_5453);
nand U8348 (N_8348,N_7218,N_6200);
nor U8349 (N_8349,N_5131,N_6931);
nand U8350 (N_8350,N_6662,N_7207);
or U8351 (N_8351,N_6725,N_5257);
nor U8352 (N_8352,N_7033,N_6461);
and U8353 (N_8353,N_6989,N_6663);
or U8354 (N_8354,N_7206,N_6143);
or U8355 (N_8355,N_6089,N_7308);
or U8356 (N_8356,N_5774,N_5343);
nand U8357 (N_8357,N_5045,N_7302);
or U8358 (N_8358,N_6134,N_7415);
nand U8359 (N_8359,N_6459,N_5375);
or U8360 (N_8360,N_6184,N_5935);
nand U8361 (N_8361,N_5940,N_5699);
or U8362 (N_8362,N_6015,N_6116);
or U8363 (N_8363,N_5218,N_6221);
or U8364 (N_8364,N_7283,N_6403);
or U8365 (N_8365,N_6531,N_6470);
or U8366 (N_8366,N_5921,N_7148);
nor U8367 (N_8367,N_7001,N_5283);
nor U8368 (N_8368,N_6676,N_6724);
nand U8369 (N_8369,N_6389,N_7076);
and U8370 (N_8370,N_5502,N_6215);
nand U8371 (N_8371,N_7084,N_5548);
nand U8372 (N_8372,N_7090,N_6357);
nor U8373 (N_8373,N_5607,N_6294);
and U8374 (N_8374,N_7487,N_5258);
and U8375 (N_8375,N_5687,N_6830);
or U8376 (N_8376,N_5741,N_7359);
nand U8377 (N_8377,N_5359,N_7270);
and U8378 (N_8378,N_7228,N_6490);
or U8379 (N_8379,N_6528,N_5306);
and U8380 (N_8380,N_5964,N_7060);
nand U8381 (N_8381,N_6392,N_7144);
nand U8382 (N_8382,N_6887,N_7309);
or U8383 (N_8383,N_5775,N_7310);
or U8384 (N_8384,N_5253,N_6365);
or U8385 (N_8385,N_5049,N_6014);
and U8386 (N_8386,N_7016,N_5963);
nor U8387 (N_8387,N_5075,N_5712);
nor U8388 (N_8388,N_7464,N_5994);
or U8389 (N_8389,N_5477,N_5120);
and U8390 (N_8390,N_7447,N_6827);
nand U8391 (N_8391,N_7455,N_7273);
nand U8392 (N_8392,N_7202,N_5601);
and U8393 (N_8393,N_5174,N_5588);
nand U8394 (N_8394,N_5274,N_7398);
nor U8395 (N_8395,N_6466,N_7171);
or U8396 (N_8396,N_6001,N_5612);
nand U8397 (N_8397,N_7122,N_6408);
and U8398 (N_8398,N_5530,N_6903);
or U8399 (N_8399,N_5872,N_6862);
or U8400 (N_8400,N_6927,N_5366);
and U8401 (N_8401,N_6546,N_7225);
and U8402 (N_8402,N_6249,N_5781);
and U8403 (N_8403,N_6856,N_7220);
nor U8404 (N_8404,N_6860,N_5301);
nand U8405 (N_8405,N_6945,N_7287);
nand U8406 (N_8406,N_5907,N_5533);
nor U8407 (N_8407,N_7346,N_6264);
and U8408 (N_8408,N_5732,N_7064);
or U8409 (N_8409,N_5608,N_6563);
nand U8410 (N_8410,N_6482,N_7063);
nor U8411 (N_8411,N_5567,N_7168);
and U8412 (N_8412,N_6326,N_6443);
and U8413 (N_8413,N_6047,N_5583);
nand U8414 (N_8414,N_5242,N_5418);
nand U8415 (N_8415,N_6850,N_7383);
nor U8416 (N_8416,N_5040,N_6566);
or U8417 (N_8417,N_7329,N_7152);
nand U8418 (N_8418,N_5228,N_6040);
and U8419 (N_8419,N_6434,N_5317);
and U8420 (N_8420,N_6644,N_5927);
xor U8421 (N_8421,N_7136,N_7204);
or U8422 (N_8422,N_5730,N_6275);
nor U8423 (N_8423,N_6038,N_6174);
nand U8424 (N_8424,N_6358,N_6716);
and U8425 (N_8425,N_7125,N_5706);
and U8426 (N_8426,N_5126,N_6572);
and U8427 (N_8427,N_5547,N_7416);
nor U8428 (N_8428,N_7208,N_5010);
or U8429 (N_8429,N_7129,N_6203);
nor U8430 (N_8430,N_6744,N_5894);
nand U8431 (N_8431,N_6236,N_5577);
nor U8432 (N_8432,N_6713,N_5532);
or U8433 (N_8433,N_6198,N_5334);
or U8434 (N_8434,N_5554,N_6067);
nand U8435 (N_8435,N_5023,N_6840);
nand U8436 (N_8436,N_6139,N_6718);
and U8437 (N_8437,N_7386,N_6481);
nor U8438 (N_8438,N_5035,N_7234);
and U8439 (N_8439,N_7498,N_7139);
nand U8440 (N_8440,N_5793,N_5419);
nand U8441 (N_8441,N_7256,N_6690);
nor U8442 (N_8442,N_5330,N_6882);
or U8443 (N_8443,N_6670,N_7271);
nand U8444 (N_8444,N_6406,N_5152);
and U8445 (N_8445,N_7021,N_6574);
nor U8446 (N_8446,N_5405,N_6993);
and U8447 (N_8447,N_5153,N_7215);
nand U8448 (N_8448,N_5727,N_6030);
nor U8449 (N_8449,N_5450,N_6098);
nand U8450 (N_8450,N_5733,N_5256);
or U8451 (N_8451,N_5660,N_6723);
xor U8452 (N_8452,N_5765,N_6187);
xor U8453 (N_8453,N_5239,N_6238);
xor U8454 (N_8454,N_6337,N_5620);
or U8455 (N_8455,N_7009,N_5545);
xnor U8456 (N_8456,N_5326,N_7123);
nand U8457 (N_8457,N_5957,N_5248);
or U8458 (N_8458,N_5636,N_5273);
nor U8459 (N_8459,N_7409,N_5091);
nand U8460 (N_8460,N_6269,N_5685);
nand U8461 (N_8461,N_6349,N_5395);
xor U8462 (N_8462,N_6343,N_6620);
nor U8463 (N_8463,N_7454,N_5141);
and U8464 (N_8464,N_6096,N_6278);
nor U8465 (N_8465,N_6292,N_6614);
xor U8466 (N_8466,N_7100,N_6996);
nand U8467 (N_8467,N_6627,N_6693);
and U8468 (N_8468,N_6900,N_5861);
nor U8469 (N_8469,N_5739,N_7395);
nand U8470 (N_8470,N_5404,N_5232);
nand U8471 (N_8471,N_5108,N_5576);
nor U8472 (N_8472,N_7341,N_6497);
nand U8473 (N_8473,N_6021,N_7446);
or U8474 (N_8474,N_5591,N_6634);
and U8475 (N_8475,N_7328,N_5830);
nor U8476 (N_8476,N_7441,N_7410);
or U8477 (N_8477,N_7040,N_6573);
or U8478 (N_8478,N_7366,N_6792);
xnor U8479 (N_8479,N_7285,N_5252);
nor U8480 (N_8480,N_5575,N_6396);
nor U8481 (N_8481,N_7055,N_5656);
nand U8482 (N_8482,N_5308,N_6474);
nand U8483 (N_8483,N_7058,N_6587);
nor U8484 (N_8484,N_5347,N_6265);
nor U8485 (N_8485,N_5272,N_5696);
and U8486 (N_8486,N_5863,N_6179);
nor U8487 (N_8487,N_6625,N_6883);
nor U8488 (N_8488,N_6948,N_6920);
or U8489 (N_8489,N_6960,N_5766);
nand U8490 (N_8490,N_6043,N_7419);
and U8491 (N_8491,N_7108,N_6631);
nand U8492 (N_8492,N_6570,N_5029);
nand U8493 (N_8493,N_6817,N_6370);
nor U8494 (N_8494,N_6642,N_6771);
xnor U8495 (N_8495,N_5302,N_5631);
or U8496 (N_8496,N_5458,N_6648);
or U8497 (N_8497,N_5171,N_6916);
xnor U8498 (N_8498,N_6453,N_7071);
nand U8499 (N_8499,N_6682,N_6825);
nor U8500 (N_8500,N_7330,N_6909);
nand U8501 (N_8501,N_6167,N_6515);
nor U8502 (N_8502,N_5615,N_5214);
nand U8503 (N_8503,N_5498,N_6338);
or U8504 (N_8504,N_6201,N_7190);
nor U8505 (N_8505,N_5754,N_5807);
and U8506 (N_8506,N_5095,N_5265);
nand U8507 (N_8507,N_7439,N_5480);
xnor U8508 (N_8508,N_6438,N_5208);
and U8509 (N_8509,N_5846,N_6610);
nand U8510 (N_8510,N_6316,N_6770);
or U8511 (N_8511,N_6013,N_5684);
nor U8512 (N_8512,N_5083,N_6332);
xor U8513 (N_8513,N_6429,N_5936);
or U8514 (N_8514,N_6136,N_7290);
nand U8515 (N_8515,N_5400,N_6058);
nand U8516 (N_8516,N_6655,N_5363);
or U8517 (N_8517,N_5590,N_7315);
and U8518 (N_8518,N_6071,N_6251);
nand U8519 (N_8519,N_5683,N_5645);
nor U8520 (N_8520,N_5622,N_7127);
xor U8521 (N_8521,N_6867,N_5072);
nor U8522 (N_8522,N_5870,N_5184);
nand U8523 (N_8523,N_6285,N_6309);
or U8524 (N_8524,N_7356,N_6633);
or U8525 (N_8525,N_5637,N_6130);
nor U8526 (N_8526,N_5204,N_6556);
nor U8527 (N_8527,N_5057,N_6802);
or U8528 (N_8528,N_6618,N_7186);
xnor U8529 (N_8529,N_6022,N_5966);
or U8530 (N_8530,N_6118,N_6360);
or U8531 (N_8531,N_6239,N_6511);
and U8532 (N_8532,N_7355,N_6823);
or U8533 (N_8533,N_6376,N_5077);
and U8534 (N_8534,N_6320,N_6969);
xor U8535 (N_8535,N_5558,N_5653);
or U8536 (N_8536,N_7158,N_7449);
nor U8537 (N_8537,N_5709,N_5515);
xnor U8538 (N_8538,N_7306,N_5794);
nand U8539 (N_8539,N_6808,N_7068);
nand U8540 (N_8540,N_5799,N_5133);
and U8541 (N_8541,N_6189,N_6124);
nor U8542 (N_8542,N_5538,N_6597);
nand U8543 (N_8543,N_6645,N_6449);
nand U8544 (N_8544,N_7221,N_6505);
or U8545 (N_8545,N_5424,N_6485);
xor U8546 (N_8546,N_5189,N_6894);
or U8547 (N_8547,N_6268,N_7223);
or U8548 (N_8548,N_5314,N_5705);
nand U8549 (N_8549,N_6451,N_6042);
nand U8550 (N_8550,N_6243,N_7119);
and U8551 (N_8551,N_5671,N_5177);
nand U8552 (N_8552,N_5379,N_6356);
nand U8553 (N_8553,N_7471,N_6153);
nor U8554 (N_8554,N_6760,N_7006);
and U8555 (N_8555,N_5492,N_5946);
and U8556 (N_8556,N_5409,N_5904);
or U8557 (N_8557,N_5369,N_6374);
nand U8558 (N_8558,N_5647,N_7229);
nand U8559 (N_8559,N_6019,N_6669);
or U8560 (N_8560,N_6435,N_6250);
nor U8561 (N_8561,N_5856,N_5448);
or U8562 (N_8562,N_5382,N_7470);
nor U8563 (N_8563,N_6244,N_6794);
nand U8564 (N_8564,N_7304,N_5234);
or U8565 (N_8565,N_5543,N_5707);
or U8566 (N_8566,N_7399,N_6362);
or U8567 (N_8567,N_6891,N_6738);
nor U8568 (N_8568,N_7034,N_7406);
and U8569 (N_8569,N_5271,N_6846);
and U8570 (N_8570,N_7244,N_6946);
and U8571 (N_8571,N_7432,N_5139);
nand U8572 (N_8572,N_6150,N_6176);
and U8573 (N_8573,N_5666,N_6904);
and U8574 (N_8574,N_6149,N_5151);
or U8575 (N_8575,N_5200,N_5099);
xnor U8576 (N_8576,N_7277,N_5815);
and U8577 (N_8577,N_5984,N_6688);
and U8578 (N_8578,N_5717,N_7013);
nand U8579 (N_8579,N_5244,N_7426);
nand U8580 (N_8580,N_5692,N_6080);
nand U8581 (N_8581,N_7077,N_5972);
nor U8582 (N_8582,N_6061,N_7482);
and U8583 (N_8583,N_6719,N_7337);
or U8584 (N_8584,N_6647,N_5006);
and U8585 (N_8585,N_7477,N_5180);
and U8586 (N_8586,N_5183,N_6984);
and U8587 (N_8587,N_5943,N_5081);
or U8588 (N_8588,N_5451,N_6261);
or U8589 (N_8589,N_7314,N_5550);
nor U8590 (N_8590,N_5960,N_7233);
and U8591 (N_8591,N_5079,N_7433);
nand U8592 (N_8592,N_6348,N_5288);
nor U8593 (N_8593,N_5997,N_6480);
or U8594 (N_8594,N_6726,N_6567);
and U8595 (N_8595,N_6905,N_6551);
xnor U8596 (N_8596,N_6980,N_7375);
or U8597 (N_8597,N_6807,N_5562);
nand U8598 (N_8598,N_6086,N_5721);
xnor U8599 (N_8599,N_7374,N_6710);
nor U8600 (N_8600,N_7397,N_5630);
or U8601 (N_8601,N_6600,N_6486);
nand U8602 (N_8602,N_6562,N_5243);
xnor U8603 (N_8603,N_6119,N_5078);
and U8604 (N_8604,N_5574,N_5546);
and U8605 (N_8605,N_5378,N_6651);
or U8606 (N_8606,N_5011,N_5417);
nand U8607 (N_8607,N_7093,N_6335);
nand U8608 (N_8608,N_5518,N_5813);
and U8609 (N_8609,N_5849,N_5638);
nand U8610 (N_8610,N_7083,N_5466);
and U8611 (N_8611,N_6419,N_6380);
nor U8612 (N_8612,N_7026,N_6687);
or U8613 (N_8613,N_6368,N_6577);
nand U8614 (N_8614,N_6057,N_5185);
and U8615 (N_8615,N_5155,N_6961);
nor U8616 (N_8616,N_6691,N_6097);
and U8617 (N_8617,N_5349,N_7272);
and U8618 (N_8618,N_7162,N_5474);
nor U8619 (N_8619,N_5462,N_7117);
nor U8620 (N_8620,N_5031,N_6616);
and U8621 (N_8621,N_7242,N_7116);
or U8622 (N_8622,N_6864,N_5509);
nand U8623 (N_8623,N_6317,N_6345);
nand U8624 (N_8624,N_5587,N_6745);
nor U8625 (N_8625,N_7044,N_7106);
nor U8626 (N_8626,N_7469,N_5604);
nand U8627 (N_8627,N_5290,N_5761);
nor U8628 (N_8628,N_5489,N_6789);
nand U8629 (N_8629,N_6609,N_5689);
or U8630 (N_8630,N_5961,N_5024);
or U8631 (N_8631,N_5882,N_7389);
nand U8632 (N_8632,N_5034,N_5522);
nor U8633 (N_8633,N_5486,N_7390);
and U8634 (N_8634,N_6639,N_6696);
nand U8635 (N_8635,N_6674,N_7305);
nor U8636 (N_8636,N_7061,N_6928);
nand U8637 (N_8637,N_6402,N_5535);
nor U8638 (N_8638,N_5891,N_6056);
nand U8639 (N_8639,N_7348,N_6966);
nor U8640 (N_8640,N_6605,N_5955);
xnor U8641 (N_8641,N_6907,N_6874);
and U8642 (N_8642,N_6530,N_7177);
and U8643 (N_8643,N_5555,N_6590);
and U8644 (N_8644,N_7460,N_6733);
or U8645 (N_8645,N_5365,N_7048);
or U8646 (N_8646,N_6819,N_7046);
or U8647 (N_8647,N_5009,N_7212);
or U8648 (N_8648,N_5336,N_5279);
xor U8649 (N_8649,N_5402,N_6274);
nor U8650 (N_8650,N_6428,N_5839);
and U8651 (N_8651,N_5824,N_6114);
or U8652 (N_8652,N_7424,N_5884);
nand U8653 (N_8653,N_5883,N_5277);
nor U8654 (N_8654,N_7107,N_6237);
or U8655 (N_8655,N_6854,N_5540);
nand U8656 (N_8656,N_6565,N_5635);
nor U8657 (N_8657,N_6964,N_5406);
xor U8658 (N_8658,N_5146,N_6799);
or U8659 (N_8659,N_6985,N_7246);
nand U8660 (N_8660,N_6683,N_6088);
nand U8661 (N_8661,N_5323,N_5674);
or U8662 (N_8662,N_7417,N_6273);
nor U8663 (N_8663,N_6154,N_5939);
and U8664 (N_8664,N_5951,N_6331);
nand U8665 (N_8665,N_5074,N_7263);
and U8666 (N_8666,N_5848,N_5210);
xnor U8667 (N_8667,N_6849,N_7448);
nor U8668 (N_8668,N_5680,N_5043);
xnor U8669 (N_8669,N_6499,N_6420);
nor U8670 (N_8670,N_5835,N_5759);
xor U8671 (N_8671,N_5000,N_5310);
nor U8672 (N_8672,N_5981,N_5916);
nor U8673 (N_8673,N_6393,N_6445);
nor U8674 (N_8674,N_5225,N_6541);
or U8675 (N_8675,N_7249,N_6260);
nand U8676 (N_8676,N_6548,N_5679);
and U8677 (N_8677,N_5341,N_6814);
and U8678 (N_8678,N_6020,N_7156);
and U8679 (N_8679,N_7112,N_6192);
or U8680 (N_8680,N_7428,N_6947);
nand U8681 (N_8681,N_5254,N_7402);
or U8682 (N_8682,N_6857,N_6684);
and U8683 (N_8683,N_5889,N_6753);
nor U8684 (N_8684,N_6161,N_7325);
or U8685 (N_8685,N_5500,N_6608);
nand U8686 (N_8686,N_6027,N_7027);
or U8687 (N_8687,N_5768,N_5565);
and U8688 (N_8688,N_6462,N_6561);
and U8689 (N_8689,N_5193,N_7073);
nand U8690 (N_8690,N_6507,N_6720);
or U8691 (N_8691,N_7293,N_5478);
or U8692 (N_8692,N_7038,N_5681);
xnor U8693 (N_8693,N_5380,N_6534);
or U8694 (N_8694,N_7364,N_6106);
or U8695 (N_8695,N_6958,N_6218);
and U8696 (N_8696,N_5261,N_5503);
nor U8697 (N_8697,N_5431,N_5890);
or U8698 (N_8698,N_5053,N_5384);
nand U8699 (N_8699,N_5167,N_6537);
nor U8700 (N_8700,N_5460,N_6971);
nor U8701 (N_8701,N_5270,N_6009);
and U8702 (N_8702,N_5931,N_6135);
xor U8703 (N_8703,N_5026,N_6012);
and U8704 (N_8704,N_6654,N_6848);
nor U8705 (N_8705,N_6367,N_5749);
nand U8706 (N_8706,N_5129,N_5950);
nor U8707 (N_8707,N_5658,N_7344);
xor U8708 (N_8708,N_5974,N_5259);
nand U8709 (N_8709,N_6035,N_5097);
and U8710 (N_8710,N_5381,N_7102);
or U8711 (N_8711,N_6413,N_6424);
nor U8712 (N_8712,N_7103,N_7028);
or U8713 (N_8713,N_6974,N_7132);
or U8714 (N_8714,N_7332,N_5728);
and U8715 (N_8715,N_6400,N_5490);
nand U8716 (N_8716,N_6032,N_6224);
or U8717 (N_8717,N_5834,N_5013);
xnor U8718 (N_8718,N_6169,N_5162);
and U8719 (N_8719,N_6667,N_7392);
or U8720 (N_8720,N_6504,N_5201);
or U8721 (N_8721,N_6508,N_5101);
nand U8722 (N_8722,N_6313,N_5003);
nor U8723 (N_8723,N_7019,N_5594);
nor U8724 (N_8724,N_5113,N_6796);
nor U8725 (N_8725,N_5086,N_5468);
nand U8726 (N_8726,N_6105,N_7010);
and U8727 (N_8727,N_7320,N_5715);
and U8728 (N_8728,N_7167,N_6873);
nor U8729 (N_8729,N_6580,N_6870);
and U8730 (N_8730,N_7377,N_5922);
nor U8731 (N_8731,N_5089,N_6247);
xor U8732 (N_8732,N_7373,N_6711);
nor U8733 (N_8733,N_6122,N_6456);
nor U8734 (N_8734,N_6390,N_6611);
and U8735 (N_8735,N_5651,N_5719);
or U8736 (N_8736,N_6432,N_6039);
nor U8737 (N_8737,N_6518,N_7074);
nand U8738 (N_8738,N_7081,N_6128);
nand U8739 (N_8739,N_5690,N_5520);
nor U8740 (N_8740,N_5625,N_7313);
and U8741 (N_8741,N_7420,N_7236);
and U8742 (N_8742,N_7004,N_6371);
and U8743 (N_8743,N_6736,N_6769);
and U8744 (N_8744,N_5062,N_6829);
nand U8745 (N_8745,N_7403,N_6457);
nand U8746 (N_8746,N_5440,N_5191);
xor U8747 (N_8747,N_6036,N_5819);
nand U8748 (N_8748,N_5757,N_5661);
or U8749 (N_8749,N_5445,N_5364);
xor U8750 (N_8750,N_5747,N_6194);
nor U8751 (N_8751,N_6288,N_6432);
xor U8752 (N_8752,N_6138,N_6707);
or U8753 (N_8753,N_6594,N_6603);
nand U8754 (N_8754,N_5857,N_6593);
xnor U8755 (N_8755,N_6522,N_6119);
nand U8756 (N_8756,N_7371,N_5046);
nor U8757 (N_8757,N_5872,N_6800);
nand U8758 (N_8758,N_5284,N_5132);
and U8759 (N_8759,N_5813,N_7031);
and U8760 (N_8760,N_7269,N_7456);
nand U8761 (N_8761,N_7344,N_5751);
nand U8762 (N_8762,N_5363,N_7204);
nand U8763 (N_8763,N_5742,N_7153);
nand U8764 (N_8764,N_5850,N_6863);
and U8765 (N_8765,N_6213,N_6099);
and U8766 (N_8766,N_6786,N_7484);
and U8767 (N_8767,N_5815,N_5426);
nand U8768 (N_8768,N_6580,N_6261);
nor U8769 (N_8769,N_7451,N_7438);
nor U8770 (N_8770,N_5294,N_6621);
or U8771 (N_8771,N_7359,N_6848);
nand U8772 (N_8772,N_5860,N_7145);
xnor U8773 (N_8773,N_6739,N_5975);
and U8774 (N_8774,N_6770,N_7062);
or U8775 (N_8775,N_5564,N_5749);
or U8776 (N_8776,N_6427,N_5054);
or U8777 (N_8777,N_5307,N_5756);
nor U8778 (N_8778,N_6280,N_6422);
or U8779 (N_8779,N_5033,N_7280);
nor U8780 (N_8780,N_6215,N_6466);
nand U8781 (N_8781,N_5274,N_6575);
nand U8782 (N_8782,N_5603,N_7056);
nand U8783 (N_8783,N_5106,N_6492);
or U8784 (N_8784,N_5719,N_7066);
nor U8785 (N_8785,N_5316,N_5360);
nor U8786 (N_8786,N_5998,N_6943);
nand U8787 (N_8787,N_7453,N_5284);
or U8788 (N_8788,N_6306,N_5691);
or U8789 (N_8789,N_6299,N_5138);
or U8790 (N_8790,N_5221,N_5400);
nand U8791 (N_8791,N_6718,N_6380);
nand U8792 (N_8792,N_5694,N_5712);
and U8793 (N_8793,N_6688,N_5713);
and U8794 (N_8794,N_5104,N_5282);
nor U8795 (N_8795,N_5761,N_5856);
nor U8796 (N_8796,N_6033,N_5346);
xnor U8797 (N_8797,N_5283,N_6233);
and U8798 (N_8798,N_7251,N_5430);
or U8799 (N_8799,N_6654,N_7012);
or U8800 (N_8800,N_5149,N_5088);
xor U8801 (N_8801,N_6634,N_6064);
and U8802 (N_8802,N_6657,N_6092);
or U8803 (N_8803,N_7014,N_7325);
nand U8804 (N_8804,N_7198,N_5935);
nor U8805 (N_8805,N_5219,N_6414);
or U8806 (N_8806,N_5857,N_6206);
nand U8807 (N_8807,N_7005,N_6596);
nor U8808 (N_8808,N_6296,N_7014);
nand U8809 (N_8809,N_6379,N_7111);
nor U8810 (N_8810,N_5614,N_6049);
nand U8811 (N_8811,N_6949,N_7490);
nor U8812 (N_8812,N_5283,N_6175);
nor U8813 (N_8813,N_5752,N_6380);
or U8814 (N_8814,N_5165,N_7167);
xnor U8815 (N_8815,N_6907,N_6148);
xor U8816 (N_8816,N_5318,N_6327);
nand U8817 (N_8817,N_7426,N_6809);
nor U8818 (N_8818,N_5055,N_7319);
nand U8819 (N_8819,N_5956,N_5438);
and U8820 (N_8820,N_5533,N_5388);
nand U8821 (N_8821,N_7047,N_6663);
nor U8822 (N_8822,N_7387,N_5635);
and U8823 (N_8823,N_5607,N_6004);
and U8824 (N_8824,N_6511,N_6839);
nor U8825 (N_8825,N_5705,N_6798);
or U8826 (N_8826,N_6228,N_5402);
and U8827 (N_8827,N_5938,N_5849);
nand U8828 (N_8828,N_6913,N_6565);
or U8829 (N_8829,N_6289,N_6252);
nand U8830 (N_8830,N_7009,N_5840);
and U8831 (N_8831,N_5552,N_5205);
or U8832 (N_8832,N_6472,N_6032);
nor U8833 (N_8833,N_5026,N_7347);
or U8834 (N_8834,N_7119,N_6663);
nor U8835 (N_8835,N_6822,N_5951);
nand U8836 (N_8836,N_6019,N_6892);
and U8837 (N_8837,N_5518,N_7202);
xnor U8838 (N_8838,N_7151,N_6891);
nor U8839 (N_8839,N_6946,N_6492);
and U8840 (N_8840,N_7177,N_6821);
and U8841 (N_8841,N_5603,N_6367);
and U8842 (N_8842,N_6446,N_5479);
or U8843 (N_8843,N_7398,N_5361);
and U8844 (N_8844,N_5221,N_7229);
nor U8845 (N_8845,N_5092,N_6116);
nor U8846 (N_8846,N_7452,N_5288);
nand U8847 (N_8847,N_6495,N_6312);
or U8848 (N_8848,N_7113,N_7421);
nor U8849 (N_8849,N_7342,N_6497);
or U8850 (N_8850,N_5543,N_5661);
or U8851 (N_8851,N_6535,N_7248);
and U8852 (N_8852,N_5127,N_5790);
nand U8853 (N_8853,N_7257,N_7254);
nor U8854 (N_8854,N_7073,N_6221);
or U8855 (N_8855,N_6628,N_6442);
nand U8856 (N_8856,N_7315,N_7240);
nand U8857 (N_8857,N_5043,N_7422);
nor U8858 (N_8858,N_5411,N_6701);
or U8859 (N_8859,N_6705,N_5955);
nor U8860 (N_8860,N_7269,N_7022);
or U8861 (N_8861,N_7195,N_6865);
and U8862 (N_8862,N_7340,N_7404);
and U8863 (N_8863,N_6654,N_6674);
nor U8864 (N_8864,N_6127,N_5249);
or U8865 (N_8865,N_5583,N_6222);
or U8866 (N_8866,N_6450,N_5234);
or U8867 (N_8867,N_6211,N_5145);
or U8868 (N_8868,N_5328,N_5788);
xor U8869 (N_8869,N_5583,N_6259);
or U8870 (N_8870,N_7138,N_5043);
and U8871 (N_8871,N_6219,N_5702);
or U8872 (N_8872,N_6612,N_5918);
and U8873 (N_8873,N_5771,N_6661);
or U8874 (N_8874,N_7185,N_5822);
and U8875 (N_8875,N_7218,N_6414);
and U8876 (N_8876,N_5491,N_5922);
nand U8877 (N_8877,N_6909,N_6407);
nand U8878 (N_8878,N_6076,N_6305);
and U8879 (N_8879,N_6253,N_7400);
or U8880 (N_8880,N_5289,N_6374);
and U8881 (N_8881,N_6356,N_6320);
nand U8882 (N_8882,N_5687,N_6675);
nor U8883 (N_8883,N_6448,N_5837);
nand U8884 (N_8884,N_6557,N_6941);
and U8885 (N_8885,N_7304,N_5314);
and U8886 (N_8886,N_6928,N_7093);
nand U8887 (N_8887,N_5628,N_6452);
nor U8888 (N_8888,N_6704,N_6976);
or U8889 (N_8889,N_7247,N_5384);
nand U8890 (N_8890,N_6876,N_6439);
nand U8891 (N_8891,N_6076,N_5040);
nor U8892 (N_8892,N_6064,N_6705);
nor U8893 (N_8893,N_5395,N_6925);
and U8894 (N_8894,N_7010,N_5730);
or U8895 (N_8895,N_7280,N_6896);
nand U8896 (N_8896,N_5228,N_6370);
nor U8897 (N_8897,N_7378,N_6008);
nand U8898 (N_8898,N_5876,N_5367);
or U8899 (N_8899,N_5526,N_6099);
or U8900 (N_8900,N_5353,N_6908);
and U8901 (N_8901,N_6426,N_7471);
and U8902 (N_8902,N_6377,N_6407);
nor U8903 (N_8903,N_7436,N_6686);
and U8904 (N_8904,N_6322,N_5792);
nor U8905 (N_8905,N_6974,N_7327);
xor U8906 (N_8906,N_6169,N_6614);
nand U8907 (N_8907,N_6444,N_6601);
and U8908 (N_8908,N_5989,N_6738);
and U8909 (N_8909,N_5812,N_6750);
or U8910 (N_8910,N_6822,N_6611);
nand U8911 (N_8911,N_6174,N_6388);
and U8912 (N_8912,N_7416,N_6293);
or U8913 (N_8913,N_5087,N_7249);
nor U8914 (N_8914,N_6268,N_6791);
nand U8915 (N_8915,N_7148,N_6072);
xor U8916 (N_8916,N_5561,N_5702);
nor U8917 (N_8917,N_5208,N_6805);
nand U8918 (N_8918,N_6842,N_6934);
and U8919 (N_8919,N_6305,N_5301);
nand U8920 (N_8920,N_7048,N_6119);
nor U8921 (N_8921,N_7128,N_6662);
nor U8922 (N_8922,N_5401,N_5377);
or U8923 (N_8923,N_7319,N_6504);
or U8924 (N_8924,N_7218,N_7475);
and U8925 (N_8925,N_6756,N_6699);
or U8926 (N_8926,N_6624,N_6656);
nand U8927 (N_8927,N_5667,N_7336);
nor U8928 (N_8928,N_6947,N_6113);
nor U8929 (N_8929,N_7094,N_6565);
nor U8930 (N_8930,N_6768,N_7378);
and U8931 (N_8931,N_6168,N_7244);
nor U8932 (N_8932,N_6650,N_7077);
nor U8933 (N_8933,N_6876,N_6210);
nand U8934 (N_8934,N_5083,N_7471);
nor U8935 (N_8935,N_5187,N_6713);
or U8936 (N_8936,N_7271,N_5154);
and U8937 (N_8937,N_7432,N_5573);
xnor U8938 (N_8938,N_7352,N_6658);
xor U8939 (N_8939,N_5141,N_5235);
and U8940 (N_8940,N_7347,N_6968);
nand U8941 (N_8941,N_5690,N_5364);
or U8942 (N_8942,N_5391,N_7268);
nand U8943 (N_8943,N_5768,N_5506);
nand U8944 (N_8944,N_5301,N_5055);
or U8945 (N_8945,N_5455,N_6748);
or U8946 (N_8946,N_5834,N_6147);
nand U8947 (N_8947,N_5117,N_7325);
nand U8948 (N_8948,N_5865,N_7227);
nand U8949 (N_8949,N_5161,N_5916);
or U8950 (N_8950,N_6155,N_5228);
and U8951 (N_8951,N_5608,N_5558);
and U8952 (N_8952,N_5430,N_6421);
xnor U8953 (N_8953,N_5207,N_7479);
or U8954 (N_8954,N_7188,N_6926);
and U8955 (N_8955,N_6837,N_5367);
xor U8956 (N_8956,N_6348,N_7130);
nor U8957 (N_8957,N_6607,N_5147);
or U8958 (N_8958,N_5326,N_5221);
xor U8959 (N_8959,N_7006,N_6105);
and U8960 (N_8960,N_6975,N_6059);
or U8961 (N_8961,N_5305,N_7384);
or U8962 (N_8962,N_6076,N_5753);
and U8963 (N_8963,N_6354,N_6557);
nand U8964 (N_8964,N_6226,N_7004);
and U8965 (N_8965,N_5521,N_5876);
nor U8966 (N_8966,N_6123,N_6684);
and U8967 (N_8967,N_6630,N_6194);
and U8968 (N_8968,N_6395,N_5836);
or U8969 (N_8969,N_6805,N_5905);
nor U8970 (N_8970,N_5949,N_6154);
and U8971 (N_8971,N_6829,N_5395);
nor U8972 (N_8972,N_6418,N_6607);
or U8973 (N_8973,N_6895,N_7212);
nand U8974 (N_8974,N_7250,N_6236);
or U8975 (N_8975,N_5079,N_7198);
or U8976 (N_8976,N_6430,N_7037);
or U8977 (N_8977,N_5144,N_6855);
and U8978 (N_8978,N_5318,N_7405);
nand U8979 (N_8979,N_5919,N_6903);
and U8980 (N_8980,N_7182,N_7177);
or U8981 (N_8981,N_5083,N_5804);
nand U8982 (N_8982,N_6940,N_6148);
nand U8983 (N_8983,N_7134,N_5791);
nand U8984 (N_8984,N_7410,N_6224);
or U8985 (N_8985,N_7059,N_5377);
nor U8986 (N_8986,N_5627,N_6802);
nor U8987 (N_8987,N_6512,N_7489);
and U8988 (N_8988,N_5578,N_5933);
or U8989 (N_8989,N_5418,N_6317);
nor U8990 (N_8990,N_7211,N_5283);
or U8991 (N_8991,N_5113,N_6670);
nor U8992 (N_8992,N_7208,N_5366);
or U8993 (N_8993,N_7278,N_5931);
nand U8994 (N_8994,N_6822,N_6556);
or U8995 (N_8995,N_6062,N_6814);
nand U8996 (N_8996,N_6170,N_6062);
and U8997 (N_8997,N_6754,N_6852);
nor U8998 (N_8998,N_5989,N_6487);
nor U8999 (N_8999,N_5650,N_6954);
xor U9000 (N_9000,N_5055,N_6355);
nand U9001 (N_9001,N_6636,N_5186);
and U9002 (N_9002,N_5869,N_6044);
nand U9003 (N_9003,N_5110,N_6510);
and U9004 (N_9004,N_6988,N_5167);
and U9005 (N_9005,N_5255,N_5603);
nor U9006 (N_9006,N_6751,N_6842);
nand U9007 (N_9007,N_5977,N_6819);
and U9008 (N_9008,N_5126,N_6943);
nor U9009 (N_9009,N_7424,N_7407);
nor U9010 (N_9010,N_6985,N_5672);
and U9011 (N_9011,N_6712,N_6194);
nand U9012 (N_9012,N_5316,N_5772);
and U9013 (N_9013,N_5225,N_6731);
or U9014 (N_9014,N_6698,N_7304);
and U9015 (N_9015,N_7178,N_5531);
nand U9016 (N_9016,N_5136,N_6876);
nor U9017 (N_9017,N_6190,N_6271);
and U9018 (N_9018,N_6882,N_6497);
xor U9019 (N_9019,N_6195,N_7118);
and U9020 (N_9020,N_7117,N_5206);
nand U9021 (N_9021,N_7469,N_7225);
or U9022 (N_9022,N_5547,N_5894);
and U9023 (N_9023,N_5335,N_6405);
nor U9024 (N_9024,N_5415,N_6101);
and U9025 (N_9025,N_5280,N_6889);
nor U9026 (N_9026,N_6570,N_6116);
nor U9027 (N_9027,N_5923,N_5924);
nand U9028 (N_9028,N_5695,N_7317);
nand U9029 (N_9029,N_5602,N_6455);
and U9030 (N_9030,N_5840,N_6153);
nand U9031 (N_9031,N_6708,N_7391);
or U9032 (N_9032,N_7033,N_6035);
or U9033 (N_9033,N_5792,N_5229);
xnor U9034 (N_9034,N_6883,N_6362);
xnor U9035 (N_9035,N_6812,N_7457);
and U9036 (N_9036,N_7165,N_5893);
nand U9037 (N_9037,N_5230,N_5032);
nand U9038 (N_9038,N_7337,N_6155);
or U9039 (N_9039,N_5815,N_7019);
or U9040 (N_9040,N_7439,N_5907);
or U9041 (N_9041,N_7126,N_5961);
nand U9042 (N_9042,N_6017,N_6395);
or U9043 (N_9043,N_6497,N_5728);
nor U9044 (N_9044,N_6235,N_6605);
nor U9045 (N_9045,N_6492,N_6848);
and U9046 (N_9046,N_5047,N_5330);
nand U9047 (N_9047,N_6411,N_6268);
nor U9048 (N_9048,N_5022,N_5093);
and U9049 (N_9049,N_6583,N_6071);
xor U9050 (N_9050,N_6849,N_5459);
xnor U9051 (N_9051,N_7204,N_6381);
or U9052 (N_9052,N_6877,N_5292);
nand U9053 (N_9053,N_5835,N_5755);
nor U9054 (N_9054,N_6942,N_7304);
nor U9055 (N_9055,N_6833,N_6498);
nor U9056 (N_9056,N_6908,N_7423);
nor U9057 (N_9057,N_5853,N_5551);
nor U9058 (N_9058,N_5019,N_5835);
and U9059 (N_9059,N_5467,N_6586);
nand U9060 (N_9060,N_6282,N_5637);
or U9061 (N_9061,N_7321,N_6189);
nand U9062 (N_9062,N_6894,N_6796);
nand U9063 (N_9063,N_5133,N_7064);
xnor U9064 (N_9064,N_7489,N_6619);
and U9065 (N_9065,N_5879,N_5983);
nor U9066 (N_9066,N_6268,N_6647);
and U9067 (N_9067,N_6159,N_6593);
and U9068 (N_9068,N_6162,N_7059);
nor U9069 (N_9069,N_5234,N_5493);
or U9070 (N_9070,N_7059,N_5915);
and U9071 (N_9071,N_7031,N_5769);
or U9072 (N_9072,N_7173,N_6836);
or U9073 (N_9073,N_5777,N_5468);
nand U9074 (N_9074,N_5924,N_5741);
or U9075 (N_9075,N_5997,N_5085);
nor U9076 (N_9076,N_7024,N_6855);
xnor U9077 (N_9077,N_7023,N_5536);
and U9078 (N_9078,N_5730,N_6928);
xor U9079 (N_9079,N_7104,N_6320);
or U9080 (N_9080,N_6790,N_7205);
and U9081 (N_9081,N_5436,N_6371);
and U9082 (N_9082,N_7201,N_6488);
nand U9083 (N_9083,N_5367,N_7134);
nand U9084 (N_9084,N_6625,N_6059);
and U9085 (N_9085,N_5403,N_5291);
nand U9086 (N_9086,N_6451,N_6758);
nor U9087 (N_9087,N_7488,N_5801);
xnor U9088 (N_9088,N_7485,N_5007);
nand U9089 (N_9089,N_5935,N_6703);
or U9090 (N_9090,N_7281,N_6059);
nand U9091 (N_9091,N_5680,N_6280);
nand U9092 (N_9092,N_6135,N_5152);
nor U9093 (N_9093,N_7040,N_5353);
or U9094 (N_9094,N_5756,N_7125);
nor U9095 (N_9095,N_6651,N_6401);
and U9096 (N_9096,N_5072,N_6007);
xnor U9097 (N_9097,N_5705,N_6491);
nand U9098 (N_9098,N_5911,N_6561);
or U9099 (N_9099,N_5497,N_6570);
nand U9100 (N_9100,N_7424,N_6877);
nand U9101 (N_9101,N_5226,N_7155);
nand U9102 (N_9102,N_6407,N_7221);
nand U9103 (N_9103,N_5176,N_6452);
nand U9104 (N_9104,N_5428,N_6012);
and U9105 (N_9105,N_6627,N_5782);
or U9106 (N_9106,N_6130,N_7364);
or U9107 (N_9107,N_5471,N_5986);
nand U9108 (N_9108,N_6998,N_7266);
nand U9109 (N_9109,N_6844,N_7276);
nor U9110 (N_9110,N_7372,N_6589);
or U9111 (N_9111,N_5587,N_6252);
xor U9112 (N_9112,N_5914,N_6093);
nand U9113 (N_9113,N_5367,N_6354);
nor U9114 (N_9114,N_6431,N_7093);
and U9115 (N_9115,N_5403,N_6253);
xnor U9116 (N_9116,N_6981,N_7104);
or U9117 (N_9117,N_6702,N_6455);
xor U9118 (N_9118,N_6981,N_6499);
and U9119 (N_9119,N_5221,N_5619);
nand U9120 (N_9120,N_7400,N_7193);
or U9121 (N_9121,N_5393,N_7340);
or U9122 (N_9122,N_7247,N_6032);
nand U9123 (N_9123,N_6416,N_5355);
or U9124 (N_9124,N_6431,N_6311);
nand U9125 (N_9125,N_6366,N_5377);
nand U9126 (N_9126,N_7493,N_6364);
nor U9127 (N_9127,N_5050,N_7309);
nor U9128 (N_9128,N_6174,N_6606);
and U9129 (N_9129,N_6917,N_5026);
and U9130 (N_9130,N_6813,N_6265);
nand U9131 (N_9131,N_6303,N_5928);
nand U9132 (N_9132,N_5944,N_7152);
nor U9133 (N_9133,N_6666,N_7351);
nand U9134 (N_9134,N_5114,N_7053);
xnor U9135 (N_9135,N_5336,N_5207);
nand U9136 (N_9136,N_6945,N_5847);
and U9137 (N_9137,N_5255,N_5488);
or U9138 (N_9138,N_6269,N_5286);
nor U9139 (N_9139,N_5867,N_6134);
nand U9140 (N_9140,N_5794,N_7209);
or U9141 (N_9141,N_5518,N_7194);
and U9142 (N_9142,N_5223,N_6462);
nand U9143 (N_9143,N_6163,N_5449);
nand U9144 (N_9144,N_5768,N_5690);
nand U9145 (N_9145,N_5483,N_5623);
xnor U9146 (N_9146,N_7111,N_6321);
or U9147 (N_9147,N_6513,N_6656);
and U9148 (N_9148,N_5688,N_5226);
and U9149 (N_9149,N_6305,N_6238);
nand U9150 (N_9150,N_6635,N_6345);
or U9151 (N_9151,N_5705,N_5655);
nor U9152 (N_9152,N_6552,N_7054);
or U9153 (N_9153,N_7470,N_6654);
or U9154 (N_9154,N_6416,N_6439);
xnor U9155 (N_9155,N_5343,N_5565);
nor U9156 (N_9156,N_5950,N_6807);
and U9157 (N_9157,N_6257,N_6042);
nand U9158 (N_9158,N_6717,N_6644);
nor U9159 (N_9159,N_7307,N_5148);
or U9160 (N_9160,N_6164,N_6493);
nand U9161 (N_9161,N_5984,N_7443);
or U9162 (N_9162,N_5651,N_7305);
nor U9163 (N_9163,N_5826,N_7000);
or U9164 (N_9164,N_7164,N_6585);
or U9165 (N_9165,N_6414,N_5615);
and U9166 (N_9166,N_5718,N_6610);
nor U9167 (N_9167,N_7130,N_6382);
or U9168 (N_9168,N_7024,N_7495);
and U9169 (N_9169,N_5474,N_5414);
and U9170 (N_9170,N_5151,N_6110);
or U9171 (N_9171,N_6891,N_6604);
and U9172 (N_9172,N_5333,N_6933);
nor U9173 (N_9173,N_7159,N_6107);
nand U9174 (N_9174,N_6168,N_5174);
xnor U9175 (N_9175,N_6263,N_5216);
nor U9176 (N_9176,N_6875,N_5246);
nor U9177 (N_9177,N_6713,N_6951);
and U9178 (N_9178,N_6769,N_5140);
nand U9179 (N_9179,N_6124,N_5568);
xor U9180 (N_9180,N_6939,N_6964);
or U9181 (N_9181,N_6479,N_5733);
nor U9182 (N_9182,N_6817,N_6432);
and U9183 (N_9183,N_7451,N_6008);
xnor U9184 (N_9184,N_7009,N_7469);
xnor U9185 (N_9185,N_5475,N_5551);
and U9186 (N_9186,N_5331,N_6032);
or U9187 (N_9187,N_5456,N_6253);
xor U9188 (N_9188,N_5718,N_5288);
nand U9189 (N_9189,N_7322,N_5906);
nand U9190 (N_9190,N_7371,N_5288);
or U9191 (N_9191,N_6482,N_6640);
nand U9192 (N_9192,N_7181,N_5635);
and U9193 (N_9193,N_6526,N_5167);
nor U9194 (N_9194,N_6964,N_5577);
nor U9195 (N_9195,N_7098,N_6237);
nor U9196 (N_9196,N_5400,N_6815);
and U9197 (N_9197,N_5535,N_7029);
nor U9198 (N_9198,N_6641,N_7275);
nand U9199 (N_9199,N_6604,N_5015);
or U9200 (N_9200,N_5545,N_6095);
nor U9201 (N_9201,N_5042,N_5106);
nand U9202 (N_9202,N_5463,N_6075);
or U9203 (N_9203,N_5050,N_5529);
nor U9204 (N_9204,N_5327,N_5890);
or U9205 (N_9205,N_7069,N_5765);
or U9206 (N_9206,N_7357,N_7117);
and U9207 (N_9207,N_7103,N_6498);
xnor U9208 (N_9208,N_6761,N_7445);
or U9209 (N_9209,N_7269,N_6408);
and U9210 (N_9210,N_6348,N_6496);
and U9211 (N_9211,N_7286,N_5133);
nor U9212 (N_9212,N_5355,N_6702);
or U9213 (N_9213,N_7063,N_6208);
or U9214 (N_9214,N_6811,N_5895);
xor U9215 (N_9215,N_5231,N_6392);
nand U9216 (N_9216,N_6093,N_5420);
or U9217 (N_9217,N_6747,N_5051);
nand U9218 (N_9218,N_6569,N_5990);
nor U9219 (N_9219,N_6226,N_7443);
nand U9220 (N_9220,N_5130,N_6037);
nor U9221 (N_9221,N_5729,N_7242);
nand U9222 (N_9222,N_6959,N_6282);
nand U9223 (N_9223,N_5885,N_6340);
nor U9224 (N_9224,N_7483,N_5797);
and U9225 (N_9225,N_5181,N_7383);
and U9226 (N_9226,N_7072,N_5535);
nor U9227 (N_9227,N_5229,N_5799);
nor U9228 (N_9228,N_5256,N_7094);
and U9229 (N_9229,N_6337,N_7169);
xnor U9230 (N_9230,N_5184,N_7271);
xnor U9231 (N_9231,N_6269,N_6587);
nor U9232 (N_9232,N_7000,N_5662);
nor U9233 (N_9233,N_5729,N_7013);
nand U9234 (N_9234,N_6021,N_5162);
nor U9235 (N_9235,N_5744,N_5332);
or U9236 (N_9236,N_7038,N_6277);
or U9237 (N_9237,N_6104,N_5175);
and U9238 (N_9238,N_5706,N_5193);
nand U9239 (N_9239,N_5962,N_5552);
nand U9240 (N_9240,N_7157,N_6331);
nor U9241 (N_9241,N_7151,N_7472);
nand U9242 (N_9242,N_5972,N_6285);
nand U9243 (N_9243,N_6543,N_6391);
and U9244 (N_9244,N_5518,N_5109);
and U9245 (N_9245,N_5343,N_6078);
and U9246 (N_9246,N_6430,N_7204);
nand U9247 (N_9247,N_5962,N_5697);
nand U9248 (N_9248,N_5249,N_6436);
and U9249 (N_9249,N_5077,N_6550);
nor U9250 (N_9250,N_5060,N_7185);
nor U9251 (N_9251,N_7357,N_5792);
and U9252 (N_9252,N_5574,N_5381);
and U9253 (N_9253,N_6624,N_7213);
nand U9254 (N_9254,N_7151,N_5233);
and U9255 (N_9255,N_7072,N_5845);
nor U9256 (N_9256,N_5096,N_5296);
or U9257 (N_9257,N_7419,N_6077);
and U9258 (N_9258,N_6516,N_5972);
or U9259 (N_9259,N_6673,N_6012);
nand U9260 (N_9260,N_7180,N_6579);
or U9261 (N_9261,N_6730,N_5330);
and U9262 (N_9262,N_6341,N_5907);
nor U9263 (N_9263,N_5896,N_5836);
xnor U9264 (N_9264,N_6307,N_6710);
or U9265 (N_9265,N_6681,N_5664);
and U9266 (N_9266,N_6552,N_5484);
xnor U9267 (N_9267,N_6438,N_5372);
nand U9268 (N_9268,N_6667,N_6735);
nand U9269 (N_9269,N_6964,N_5461);
and U9270 (N_9270,N_5000,N_6110);
and U9271 (N_9271,N_5874,N_5487);
or U9272 (N_9272,N_5743,N_6790);
nand U9273 (N_9273,N_6221,N_6887);
or U9274 (N_9274,N_5301,N_5011);
nor U9275 (N_9275,N_7356,N_6090);
or U9276 (N_9276,N_5958,N_6258);
nand U9277 (N_9277,N_5213,N_7416);
or U9278 (N_9278,N_6192,N_5592);
xor U9279 (N_9279,N_5626,N_5110);
nor U9280 (N_9280,N_7211,N_6442);
and U9281 (N_9281,N_7467,N_6896);
and U9282 (N_9282,N_5847,N_6178);
and U9283 (N_9283,N_5732,N_6992);
or U9284 (N_9284,N_6354,N_5232);
nand U9285 (N_9285,N_5780,N_6323);
and U9286 (N_9286,N_5535,N_7022);
or U9287 (N_9287,N_5987,N_5118);
nor U9288 (N_9288,N_6501,N_6918);
nand U9289 (N_9289,N_7437,N_5516);
nand U9290 (N_9290,N_6813,N_5179);
nand U9291 (N_9291,N_7329,N_7175);
nand U9292 (N_9292,N_6871,N_5645);
nand U9293 (N_9293,N_5984,N_6513);
and U9294 (N_9294,N_6539,N_5450);
and U9295 (N_9295,N_6525,N_7478);
and U9296 (N_9296,N_6532,N_5091);
and U9297 (N_9297,N_7154,N_7416);
and U9298 (N_9298,N_6643,N_6133);
nand U9299 (N_9299,N_7039,N_7045);
nor U9300 (N_9300,N_6833,N_7051);
or U9301 (N_9301,N_6861,N_5982);
or U9302 (N_9302,N_7393,N_5859);
and U9303 (N_9303,N_5971,N_5357);
or U9304 (N_9304,N_5389,N_7134);
or U9305 (N_9305,N_5359,N_6016);
and U9306 (N_9306,N_6210,N_5635);
nor U9307 (N_9307,N_6955,N_6317);
and U9308 (N_9308,N_6247,N_6239);
or U9309 (N_9309,N_7244,N_7373);
and U9310 (N_9310,N_7069,N_5792);
nand U9311 (N_9311,N_7152,N_6366);
nand U9312 (N_9312,N_6935,N_7037);
nand U9313 (N_9313,N_5054,N_7446);
or U9314 (N_9314,N_5992,N_6703);
or U9315 (N_9315,N_5880,N_7303);
nor U9316 (N_9316,N_5005,N_6606);
or U9317 (N_9317,N_7115,N_5542);
and U9318 (N_9318,N_5902,N_7448);
nor U9319 (N_9319,N_5872,N_6521);
nand U9320 (N_9320,N_5594,N_5816);
and U9321 (N_9321,N_6766,N_5511);
nand U9322 (N_9322,N_5345,N_5457);
or U9323 (N_9323,N_5059,N_5089);
nand U9324 (N_9324,N_7258,N_6628);
or U9325 (N_9325,N_5873,N_6859);
and U9326 (N_9326,N_5741,N_5242);
and U9327 (N_9327,N_6718,N_5438);
nand U9328 (N_9328,N_6238,N_6010);
nor U9329 (N_9329,N_7482,N_6177);
and U9330 (N_9330,N_7024,N_7107);
or U9331 (N_9331,N_5660,N_5515);
nand U9332 (N_9332,N_5590,N_6335);
nand U9333 (N_9333,N_6085,N_6069);
nand U9334 (N_9334,N_5775,N_6452);
nand U9335 (N_9335,N_7488,N_6645);
xnor U9336 (N_9336,N_6716,N_7381);
and U9337 (N_9337,N_7225,N_5585);
nand U9338 (N_9338,N_6052,N_5962);
nor U9339 (N_9339,N_6302,N_5997);
nand U9340 (N_9340,N_7355,N_5465);
and U9341 (N_9341,N_5432,N_7483);
and U9342 (N_9342,N_6000,N_7380);
and U9343 (N_9343,N_6432,N_6490);
or U9344 (N_9344,N_5701,N_6682);
nand U9345 (N_9345,N_7407,N_7357);
nand U9346 (N_9346,N_7292,N_6843);
and U9347 (N_9347,N_5878,N_6533);
and U9348 (N_9348,N_5298,N_5654);
and U9349 (N_9349,N_5621,N_6503);
nand U9350 (N_9350,N_5980,N_7399);
nor U9351 (N_9351,N_5550,N_5517);
and U9352 (N_9352,N_6733,N_5411);
or U9353 (N_9353,N_7204,N_5479);
and U9354 (N_9354,N_5641,N_5897);
or U9355 (N_9355,N_6799,N_6242);
and U9356 (N_9356,N_5843,N_5502);
nand U9357 (N_9357,N_7278,N_5600);
xnor U9358 (N_9358,N_6066,N_5365);
nand U9359 (N_9359,N_5367,N_6003);
nand U9360 (N_9360,N_5765,N_7056);
xnor U9361 (N_9361,N_5180,N_6937);
nand U9362 (N_9362,N_6844,N_6746);
nor U9363 (N_9363,N_6753,N_5360);
nand U9364 (N_9364,N_5244,N_5053);
nand U9365 (N_9365,N_6920,N_6918);
or U9366 (N_9366,N_7237,N_6132);
and U9367 (N_9367,N_7037,N_5767);
or U9368 (N_9368,N_6595,N_5056);
xnor U9369 (N_9369,N_6421,N_6130);
or U9370 (N_9370,N_5471,N_5934);
or U9371 (N_9371,N_5369,N_6102);
and U9372 (N_9372,N_7432,N_5880);
nor U9373 (N_9373,N_6488,N_6195);
and U9374 (N_9374,N_6357,N_5248);
nor U9375 (N_9375,N_5000,N_5370);
or U9376 (N_9376,N_6254,N_6020);
nand U9377 (N_9377,N_5837,N_6774);
nand U9378 (N_9378,N_6622,N_7468);
and U9379 (N_9379,N_6162,N_6480);
or U9380 (N_9380,N_5370,N_5940);
nor U9381 (N_9381,N_6377,N_5591);
xnor U9382 (N_9382,N_7394,N_5256);
nor U9383 (N_9383,N_5760,N_7493);
nand U9384 (N_9384,N_7488,N_5597);
or U9385 (N_9385,N_7062,N_6166);
nor U9386 (N_9386,N_6403,N_6063);
xnor U9387 (N_9387,N_6729,N_7428);
or U9388 (N_9388,N_5247,N_7212);
nand U9389 (N_9389,N_6713,N_6464);
nor U9390 (N_9390,N_5594,N_7322);
xor U9391 (N_9391,N_5676,N_6668);
and U9392 (N_9392,N_5732,N_7438);
xnor U9393 (N_9393,N_7432,N_5794);
nor U9394 (N_9394,N_5561,N_5472);
nor U9395 (N_9395,N_5392,N_7292);
and U9396 (N_9396,N_5264,N_6638);
or U9397 (N_9397,N_6381,N_6089);
xnor U9398 (N_9398,N_5494,N_6670);
or U9399 (N_9399,N_5497,N_6260);
xor U9400 (N_9400,N_5433,N_5354);
and U9401 (N_9401,N_5062,N_7106);
nor U9402 (N_9402,N_5303,N_5163);
and U9403 (N_9403,N_5409,N_6197);
or U9404 (N_9404,N_5414,N_6240);
or U9405 (N_9405,N_6168,N_6852);
nand U9406 (N_9406,N_5833,N_7042);
and U9407 (N_9407,N_6877,N_5497);
nor U9408 (N_9408,N_6784,N_5450);
and U9409 (N_9409,N_6897,N_7330);
nand U9410 (N_9410,N_6167,N_6340);
nand U9411 (N_9411,N_6690,N_6377);
nor U9412 (N_9412,N_7262,N_6408);
or U9413 (N_9413,N_6469,N_6730);
or U9414 (N_9414,N_7390,N_5958);
and U9415 (N_9415,N_7460,N_7385);
and U9416 (N_9416,N_5763,N_5145);
or U9417 (N_9417,N_6232,N_7131);
xor U9418 (N_9418,N_6806,N_5798);
and U9419 (N_9419,N_5967,N_5958);
nand U9420 (N_9420,N_5532,N_5444);
nor U9421 (N_9421,N_6671,N_6885);
nand U9422 (N_9422,N_6237,N_6892);
or U9423 (N_9423,N_6716,N_5585);
nor U9424 (N_9424,N_5519,N_6276);
or U9425 (N_9425,N_5067,N_5981);
nor U9426 (N_9426,N_5739,N_5542);
or U9427 (N_9427,N_6633,N_6368);
nand U9428 (N_9428,N_6370,N_7088);
or U9429 (N_9429,N_5235,N_6767);
nor U9430 (N_9430,N_6585,N_5992);
or U9431 (N_9431,N_6775,N_6773);
xor U9432 (N_9432,N_7495,N_6147);
or U9433 (N_9433,N_5370,N_5463);
nand U9434 (N_9434,N_6785,N_6762);
nor U9435 (N_9435,N_7045,N_5050);
xor U9436 (N_9436,N_6738,N_6951);
or U9437 (N_9437,N_6450,N_5725);
and U9438 (N_9438,N_7084,N_6157);
and U9439 (N_9439,N_5213,N_5358);
nor U9440 (N_9440,N_6361,N_5627);
or U9441 (N_9441,N_6221,N_6019);
nor U9442 (N_9442,N_5141,N_6963);
or U9443 (N_9443,N_6776,N_5007);
nor U9444 (N_9444,N_5863,N_7406);
or U9445 (N_9445,N_7456,N_6212);
nand U9446 (N_9446,N_6423,N_6243);
nor U9447 (N_9447,N_5172,N_6878);
nor U9448 (N_9448,N_5501,N_6637);
nor U9449 (N_9449,N_6577,N_7011);
nor U9450 (N_9450,N_5138,N_6981);
nand U9451 (N_9451,N_6277,N_5361);
xnor U9452 (N_9452,N_6954,N_6404);
nor U9453 (N_9453,N_7257,N_7311);
and U9454 (N_9454,N_6330,N_7356);
and U9455 (N_9455,N_5441,N_6960);
xnor U9456 (N_9456,N_6655,N_7400);
and U9457 (N_9457,N_5345,N_5517);
nand U9458 (N_9458,N_5425,N_5095);
nor U9459 (N_9459,N_5106,N_6597);
nand U9460 (N_9460,N_6007,N_6650);
nor U9461 (N_9461,N_5769,N_5599);
and U9462 (N_9462,N_6797,N_5828);
or U9463 (N_9463,N_6521,N_6368);
and U9464 (N_9464,N_6231,N_7270);
and U9465 (N_9465,N_5940,N_5113);
and U9466 (N_9466,N_6546,N_7036);
or U9467 (N_9467,N_5513,N_5047);
xnor U9468 (N_9468,N_6365,N_5866);
and U9469 (N_9469,N_6287,N_6636);
nor U9470 (N_9470,N_7390,N_6879);
and U9471 (N_9471,N_6779,N_6790);
and U9472 (N_9472,N_5311,N_5152);
nand U9473 (N_9473,N_5013,N_6785);
or U9474 (N_9474,N_5883,N_5175);
nand U9475 (N_9475,N_6732,N_5565);
and U9476 (N_9476,N_5885,N_5817);
or U9477 (N_9477,N_7264,N_6077);
nor U9478 (N_9478,N_5597,N_6382);
xor U9479 (N_9479,N_5455,N_5464);
nand U9480 (N_9480,N_6419,N_5070);
nor U9481 (N_9481,N_6696,N_6143);
xor U9482 (N_9482,N_6485,N_5854);
nor U9483 (N_9483,N_5466,N_6520);
xnor U9484 (N_9484,N_7391,N_7363);
and U9485 (N_9485,N_5793,N_7428);
nand U9486 (N_9486,N_7440,N_5550);
xnor U9487 (N_9487,N_6244,N_6206);
nand U9488 (N_9488,N_6412,N_7243);
xor U9489 (N_9489,N_6637,N_5822);
or U9490 (N_9490,N_6109,N_5594);
xor U9491 (N_9491,N_6662,N_7264);
or U9492 (N_9492,N_5663,N_5018);
nand U9493 (N_9493,N_6593,N_5745);
nand U9494 (N_9494,N_7266,N_5739);
or U9495 (N_9495,N_7281,N_5388);
nor U9496 (N_9496,N_6863,N_5635);
or U9497 (N_9497,N_7439,N_6651);
nor U9498 (N_9498,N_5421,N_5530);
and U9499 (N_9499,N_6366,N_7452);
nand U9500 (N_9500,N_5298,N_5321);
and U9501 (N_9501,N_5894,N_6053);
and U9502 (N_9502,N_5533,N_6755);
or U9503 (N_9503,N_6704,N_6243);
or U9504 (N_9504,N_6460,N_5744);
or U9505 (N_9505,N_6196,N_7257);
nor U9506 (N_9506,N_7094,N_7219);
nor U9507 (N_9507,N_6059,N_5275);
xnor U9508 (N_9508,N_7019,N_7260);
or U9509 (N_9509,N_5842,N_5608);
or U9510 (N_9510,N_6950,N_6319);
and U9511 (N_9511,N_5444,N_5038);
nor U9512 (N_9512,N_5325,N_5633);
nor U9513 (N_9513,N_7417,N_6461);
or U9514 (N_9514,N_7125,N_6350);
and U9515 (N_9515,N_5624,N_6630);
xnor U9516 (N_9516,N_7131,N_6100);
and U9517 (N_9517,N_5596,N_5687);
xnor U9518 (N_9518,N_7043,N_5679);
nand U9519 (N_9519,N_7420,N_5717);
nor U9520 (N_9520,N_5305,N_6393);
or U9521 (N_9521,N_7186,N_5918);
or U9522 (N_9522,N_7430,N_6573);
nand U9523 (N_9523,N_5790,N_6939);
and U9524 (N_9524,N_7346,N_5002);
nor U9525 (N_9525,N_7320,N_6548);
nor U9526 (N_9526,N_5390,N_5109);
or U9527 (N_9527,N_6662,N_6481);
nor U9528 (N_9528,N_6234,N_6015);
and U9529 (N_9529,N_5977,N_5750);
nor U9530 (N_9530,N_6655,N_6846);
and U9531 (N_9531,N_5629,N_6959);
xor U9532 (N_9532,N_5401,N_6931);
and U9533 (N_9533,N_6843,N_7006);
and U9534 (N_9534,N_5238,N_5031);
nand U9535 (N_9535,N_5978,N_5671);
or U9536 (N_9536,N_7267,N_7145);
or U9537 (N_9537,N_5683,N_5739);
or U9538 (N_9538,N_7179,N_5375);
nor U9539 (N_9539,N_5708,N_7091);
nand U9540 (N_9540,N_6114,N_5453);
nand U9541 (N_9541,N_7132,N_7198);
and U9542 (N_9542,N_6399,N_5705);
nor U9543 (N_9543,N_5487,N_6345);
or U9544 (N_9544,N_6230,N_7239);
and U9545 (N_9545,N_6514,N_6811);
nand U9546 (N_9546,N_6833,N_6443);
nor U9547 (N_9547,N_5212,N_7137);
nand U9548 (N_9548,N_6060,N_6889);
or U9549 (N_9549,N_5754,N_5285);
xor U9550 (N_9550,N_7439,N_7486);
nor U9551 (N_9551,N_6456,N_6684);
or U9552 (N_9552,N_6848,N_6601);
and U9553 (N_9553,N_5134,N_6307);
nand U9554 (N_9554,N_5169,N_6593);
xor U9555 (N_9555,N_5015,N_7105);
and U9556 (N_9556,N_7469,N_6189);
nor U9557 (N_9557,N_5990,N_5251);
nand U9558 (N_9558,N_6688,N_5403);
nand U9559 (N_9559,N_7479,N_7350);
and U9560 (N_9560,N_5367,N_5336);
nand U9561 (N_9561,N_7349,N_7041);
or U9562 (N_9562,N_6745,N_6006);
or U9563 (N_9563,N_5032,N_6856);
or U9564 (N_9564,N_5375,N_5412);
nand U9565 (N_9565,N_6777,N_5164);
nor U9566 (N_9566,N_6286,N_6881);
xnor U9567 (N_9567,N_6192,N_5756);
nand U9568 (N_9568,N_5457,N_5224);
xnor U9569 (N_9569,N_6145,N_7465);
or U9570 (N_9570,N_5825,N_5294);
nor U9571 (N_9571,N_6886,N_7097);
or U9572 (N_9572,N_5876,N_6313);
nand U9573 (N_9573,N_6860,N_5589);
and U9574 (N_9574,N_7224,N_6159);
xor U9575 (N_9575,N_5567,N_5026);
xor U9576 (N_9576,N_7131,N_5226);
xnor U9577 (N_9577,N_6620,N_5254);
nor U9578 (N_9578,N_6922,N_5649);
nand U9579 (N_9579,N_6579,N_6805);
or U9580 (N_9580,N_6817,N_5723);
and U9581 (N_9581,N_5684,N_5744);
and U9582 (N_9582,N_5540,N_6077);
and U9583 (N_9583,N_7034,N_6378);
or U9584 (N_9584,N_6277,N_6749);
nand U9585 (N_9585,N_6139,N_5336);
and U9586 (N_9586,N_6332,N_7387);
nor U9587 (N_9587,N_6996,N_5207);
and U9588 (N_9588,N_5303,N_6205);
nor U9589 (N_9589,N_5241,N_5208);
and U9590 (N_9590,N_6828,N_6486);
or U9591 (N_9591,N_6992,N_5595);
and U9592 (N_9592,N_6142,N_6109);
xor U9593 (N_9593,N_6893,N_7248);
or U9594 (N_9594,N_5813,N_5390);
nand U9595 (N_9595,N_6677,N_7379);
and U9596 (N_9596,N_6168,N_5846);
nor U9597 (N_9597,N_5859,N_6646);
nor U9598 (N_9598,N_5992,N_6223);
nand U9599 (N_9599,N_7273,N_6546);
nand U9600 (N_9600,N_7042,N_7401);
or U9601 (N_9601,N_6169,N_6195);
or U9602 (N_9602,N_6024,N_6379);
nor U9603 (N_9603,N_5661,N_6990);
nand U9604 (N_9604,N_6419,N_7277);
nor U9605 (N_9605,N_6965,N_6720);
or U9606 (N_9606,N_7030,N_6325);
and U9607 (N_9607,N_7203,N_7450);
and U9608 (N_9608,N_7124,N_7252);
and U9609 (N_9609,N_6673,N_5857);
and U9610 (N_9610,N_5899,N_6950);
nor U9611 (N_9611,N_6483,N_6957);
and U9612 (N_9612,N_6959,N_7106);
or U9613 (N_9613,N_6425,N_6686);
nor U9614 (N_9614,N_5421,N_7138);
xnor U9615 (N_9615,N_6306,N_5423);
or U9616 (N_9616,N_6941,N_5523);
nand U9617 (N_9617,N_6058,N_7118);
or U9618 (N_9618,N_6137,N_5147);
nor U9619 (N_9619,N_5614,N_7033);
nand U9620 (N_9620,N_5791,N_6729);
or U9621 (N_9621,N_6466,N_6803);
nor U9622 (N_9622,N_7044,N_6414);
nand U9623 (N_9623,N_5582,N_5931);
or U9624 (N_9624,N_5607,N_5256);
nand U9625 (N_9625,N_5064,N_5534);
or U9626 (N_9626,N_6010,N_6999);
or U9627 (N_9627,N_6618,N_7220);
xnor U9628 (N_9628,N_5906,N_5558);
nor U9629 (N_9629,N_5725,N_6950);
nand U9630 (N_9630,N_6118,N_6306);
and U9631 (N_9631,N_5390,N_6471);
nand U9632 (N_9632,N_5266,N_7456);
nand U9633 (N_9633,N_6528,N_5596);
nor U9634 (N_9634,N_6294,N_5291);
nand U9635 (N_9635,N_7416,N_5685);
nor U9636 (N_9636,N_7301,N_5264);
nor U9637 (N_9637,N_6869,N_5796);
and U9638 (N_9638,N_6491,N_6721);
xnor U9639 (N_9639,N_6311,N_7358);
nor U9640 (N_9640,N_6732,N_6792);
nor U9641 (N_9641,N_6324,N_7468);
and U9642 (N_9642,N_6497,N_5188);
nand U9643 (N_9643,N_6394,N_5183);
xnor U9644 (N_9644,N_6057,N_5062);
nand U9645 (N_9645,N_6954,N_5800);
and U9646 (N_9646,N_5070,N_6324);
or U9647 (N_9647,N_7446,N_5089);
nand U9648 (N_9648,N_6236,N_7441);
and U9649 (N_9649,N_6600,N_7348);
and U9650 (N_9650,N_7316,N_5673);
xnor U9651 (N_9651,N_6024,N_6340);
nand U9652 (N_9652,N_5822,N_6913);
or U9653 (N_9653,N_5319,N_6300);
or U9654 (N_9654,N_6824,N_7384);
nand U9655 (N_9655,N_5162,N_6713);
or U9656 (N_9656,N_5373,N_7100);
nor U9657 (N_9657,N_5240,N_5651);
nor U9658 (N_9658,N_6867,N_6205);
nor U9659 (N_9659,N_6721,N_5490);
and U9660 (N_9660,N_6309,N_5828);
and U9661 (N_9661,N_6039,N_5328);
or U9662 (N_9662,N_5183,N_7131);
nand U9663 (N_9663,N_6325,N_5383);
nand U9664 (N_9664,N_6411,N_6846);
nor U9665 (N_9665,N_7048,N_5980);
nor U9666 (N_9666,N_5711,N_7205);
nand U9667 (N_9667,N_5588,N_6392);
or U9668 (N_9668,N_7335,N_6255);
nand U9669 (N_9669,N_6716,N_7217);
and U9670 (N_9670,N_5288,N_7392);
or U9671 (N_9671,N_5501,N_7103);
nor U9672 (N_9672,N_7416,N_5984);
nor U9673 (N_9673,N_7435,N_5955);
xnor U9674 (N_9674,N_6223,N_5294);
nor U9675 (N_9675,N_6961,N_6012);
xnor U9676 (N_9676,N_6122,N_5919);
nor U9677 (N_9677,N_7492,N_6208);
nand U9678 (N_9678,N_5063,N_6547);
nand U9679 (N_9679,N_5739,N_5881);
nor U9680 (N_9680,N_6206,N_6263);
xor U9681 (N_9681,N_5875,N_7445);
nor U9682 (N_9682,N_6584,N_7325);
nor U9683 (N_9683,N_7227,N_5108);
nand U9684 (N_9684,N_5172,N_5225);
nand U9685 (N_9685,N_5033,N_7031);
xor U9686 (N_9686,N_7479,N_6520);
xor U9687 (N_9687,N_6807,N_6985);
nand U9688 (N_9688,N_6913,N_6514);
or U9689 (N_9689,N_5861,N_6755);
nor U9690 (N_9690,N_5843,N_5046);
or U9691 (N_9691,N_6126,N_5528);
or U9692 (N_9692,N_5710,N_5487);
nand U9693 (N_9693,N_5424,N_5371);
nor U9694 (N_9694,N_5454,N_5147);
or U9695 (N_9695,N_5378,N_5531);
and U9696 (N_9696,N_5188,N_7054);
nand U9697 (N_9697,N_6217,N_5275);
or U9698 (N_9698,N_5159,N_6554);
and U9699 (N_9699,N_6229,N_6911);
nor U9700 (N_9700,N_7024,N_5938);
or U9701 (N_9701,N_6508,N_5523);
nand U9702 (N_9702,N_5609,N_5418);
nor U9703 (N_9703,N_5952,N_5642);
nand U9704 (N_9704,N_6097,N_5608);
nor U9705 (N_9705,N_5843,N_6700);
nand U9706 (N_9706,N_6564,N_6823);
and U9707 (N_9707,N_6518,N_5064);
or U9708 (N_9708,N_6385,N_7404);
xor U9709 (N_9709,N_6736,N_7000);
nor U9710 (N_9710,N_5198,N_5532);
or U9711 (N_9711,N_6478,N_6084);
and U9712 (N_9712,N_5666,N_5381);
or U9713 (N_9713,N_5779,N_5381);
nor U9714 (N_9714,N_6558,N_6920);
nand U9715 (N_9715,N_5329,N_6464);
nand U9716 (N_9716,N_5582,N_5585);
nand U9717 (N_9717,N_5499,N_6407);
nand U9718 (N_9718,N_7376,N_5699);
and U9719 (N_9719,N_5345,N_5685);
nor U9720 (N_9720,N_5972,N_5556);
or U9721 (N_9721,N_7232,N_5630);
nor U9722 (N_9722,N_5467,N_6289);
or U9723 (N_9723,N_7262,N_7206);
xnor U9724 (N_9724,N_7111,N_5171);
nor U9725 (N_9725,N_6005,N_5392);
nand U9726 (N_9726,N_6826,N_6645);
nor U9727 (N_9727,N_6553,N_6131);
nor U9728 (N_9728,N_6033,N_6516);
nor U9729 (N_9729,N_5133,N_7086);
nor U9730 (N_9730,N_6207,N_5418);
and U9731 (N_9731,N_6860,N_7416);
nand U9732 (N_9732,N_7299,N_5111);
nand U9733 (N_9733,N_5932,N_6567);
xnor U9734 (N_9734,N_5854,N_7477);
nor U9735 (N_9735,N_7181,N_7051);
or U9736 (N_9736,N_7466,N_7216);
or U9737 (N_9737,N_6279,N_5884);
nor U9738 (N_9738,N_6444,N_6099);
xor U9739 (N_9739,N_5371,N_6574);
nand U9740 (N_9740,N_6730,N_5778);
or U9741 (N_9741,N_5651,N_7397);
nand U9742 (N_9742,N_5827,N_7200);
nor U9743 (N_9743,N_7410,N_5596);
nand U9744 (N_9744,N_6564,N_5470);
or U9745 (N_9745,N_5882,N_5921);
nor U9746 (N_9746,N_5799,N_6645);
or U9747 (N_9747,N_5691,N_6996);
or U9748 (N_9748,N_6262,N_5502);
nor U9749 (N_9749,N_7481,N_7490);
and U9750 (N_9750,N_6125,N_6988);
and U9751 (N_9751,N_6834,N_5240);
nand U9752 (N_9752,N_5463,N_7209);
nand U9753 (N_9753,N_6900,N_6107);
xor U9754 (N_9754,N_6905,N_6813);
or U9755 (N_9755,N_6604,N_5570);
nand U9756 (N_9756,N_5907,N_5502);
nand U9757 (N_9757,N_6463,N_5351);
nand U9758 (N_9758,N_7200,N_6933);
or U9759 (N_9759,N_6403,N_7247);
or U9760 (N_9760,N_6209,N_5205);
nand U9761 (N_9761,N_6072,N_7378);
xor U9762 (N_9762,N_6718,N_6442);
nor U9763 (N_9763,N_6329,N_5529);
nor U9764 (N_9764,N_5636,N_7146);
and U9765 (N_9765,N_6551,N_7051);
nor U9766 (N_9766,N_5778,N_5365);
and U9767 (N_9767,N_6587,N_7218);
and U9768 (N_9768,N_6715,N_7101);
xnor U9769 (N_9769,N_6336,N_7000);
nand U9770 (N_9770,N_6456,N_7420);
or U9771 (N_9771,N_6548,N_6591);
xor U9772 (N_9772,N_6547,N_6078);
nor U9773 (N_9773,N_6075,N_5495);
nor U9774 (N_9774,N_5921,N_5410);
nor U9775 (N_9775,N_6849,N_6152);
nor U9776 (N_9776,N_6521,N_5198);
and U9777 (N_9777,N_5192,N_5379);
nor U9778 (N_9778,N_6962,N_5441);
nor U9779 (N_9779,N_5815,N_7431);
or U9780 (N_9780,N_5468,N_5690);
nand U9781 (N_9781,N_6781,N_6986);
nor U9782 (N_9782,N_7181,N_6049);
and U9783 (N_9783,N_7494,N_6733);
and U9784 (N_9784,N_5748,N_5016);
nand U9785 (N_9785,N_6962,N_5811);
nand U9786 (N_9786,N_6817,N_6969);
or U9787 (N_9787,N_5226,N_5199);
and U9788 (N_9788,N_5549,N_6292);
or U9789 (N_9789,N_6021,N_7231);
and U9790 (N_9790,N_6979,N_6754);
nand U9791 (N_9791,N_7173,N_6794);
and U9792 (N_9792,N_5547,N_7276);
and U9793 (N_9793,N_5983,N_5116);
and U9794 (N_9794,N_5266,N_7008);
and U9795 (N_9795,N_7445,N_6217);
and U9796 (N_9796,N_5686,N_6553);
nand U9797 (N_9797,N_6236,N_6591);
nand U9798 (N_9798,N_6478,N_6167);
nor U9799 (N_9799,N_6972,N_5399);
and U9800 (N_9800,N_5802,N_6912);
and U9801 (N_9801,N_6214,N_7333);
nor U9802 (N_9802,N_5686,N_6295);
or U9803 (N_9803,N_7304,N_5251);
nor U9804 (N_9804,N_5462,N_5880);
nand U9805 (N_9805,N_5418,N_6034);
nand U9806 (N_9806,N_6568,N_5327);
nand U9807 (N_9807,N_5433,N_6698);
nand U9808 (N_9808,N_6848,N_5809);
nand U9809 (N_9809,N_6997,N_5274);
and U9810 (N_9810,N_6482,N_5277);
or U9811 (N_9811,N_5963,N_7289);
nor U9812 (N_9812,N_5051,N_5008);
or U9813 (N_9813,N_5990,N_5253);
nand U9814 (N_9814,N_5915,N_5799);
or U9815 (N_9815,N_6515,N_6173);
and U9816 (N_9816,N_7089,N_7281);
xor U9817 (N_9817,N_6824,N_7304);
or U9818 (N_9818,N_6851,N_7173);
nand U9819 (N_9819,N_6424,N_6962);
nor U9820 (N_9820,N_7473,N_6868);
nand U9821 (N_9821,N_6930,N_5557);
xnor U9822 (N_9822,N_7416,N_6033);
and U9823 (N_9823,N_6968,N_6741);
and U9824 (N_9824,N_6422,N_5981);
and U9825 (N_9825,N_6201,N_6779);
or U9826 (N_9826,N_7086,N_5061);
nand U9827 (N_9827,N_6979,N_7133);
or U9828 (N_9828,N_5213,N_6175);
or U9829 (N_9829,N_6738,N_5711);
or U9830 (N_9830,N_6556,N_5769);
and U9831 (N_9831,N_5108,N_6082);
or U9832 (N_9832,N_6270,N_6092);
and U9833 (N_9833,N_6124,N_7129);
xnor U9834 (N_9834,N_5264,N_6677);
nand U9835 (N_9835,N_6276,N_5711);
and U9836 (N_9836,N_7142,N_6691);
and U9837 (N_9837,N_6027,N_6932);
nor U9838 (N_9838,N_5518,N_7305);
nor U9839 (N_9839,N_6190,N_5236);
nor U9840 (N_9840,N_5696,N_6444);
or U9841 (N_9841,N_6134,N_7271);
and U9842 (N_9842,N_5792,N_6121);
or U9843 (N_9843,N_7446,N_6896);
and U9844 (N_9844,N_6249,N_5336);
nor U9845 (N_9845,N_6932,N_5250);
nor U9846 (N_9846,N_6308,N_5758);
nor U9847 (N_9847,N_6548,N_6036);
nand U9848 (N_9848,N_7197,N_7242);
xor U9849 (N_9849,N_5070,N_5947);
nor U9850 (N_9850,N_5072,N_7151);
or U9851 (N_9851,N_5837,N_5961);
or U9852 (N_9852,N_5699,N_7356);
or U9853 (N_9853,N_5981,N_6028);
and U9854 (N_9854,N_5553,N_6864);
nand U9855 (N_9855,N_5412,N_6846);
nand U9856 (N_9856,N_5613,N_7476);
xnor U9857 (N_9857,N_6461,N_5060);
nand U9858 (N_9858,N_6231,N_6928);
or U9859 (N_9859,N_5953,N_5640);
nor U9860 (N_9860,N_5581,N_5495);
or U9861 (N_9861,N_7289,N_7382);
and U9862 (N_9862,N_5586,N_7091);
nor U9863 (N_9863,N_6615,N_5105);
or U9864 (N_9864,N_5184,N_6351);
nor U9865 (N_9865,N_7193,N_5150);
nor U9866 (N_9866,N_5791,N_5020);
nor U9867 (N_9867,N_6811,N_7338);
or U9868 (N_9868,N_5916,N_6936);
nand U9869 (N_9869,N_5435,N_5011);
nor U9870 (N_9870,N_5593,N_5492);
nor U9871 (N_9871,N_7460,N_7303);
nand U9872 (N_9872,N_5045,N_7283);
and U9873 (N_9873,N_6237,N_7101);
nor U9874 (N_9874,N_5128,N_6729);
or U9875 (N_9875,N_5533,N_7074);
xor U9876 (N_9876,N_7280,N_5658);
or U9877 (N_9877,N_7294,N_5637);
and U9878 (N_9878,N_6972,N_6440);
nor U9879 (N_9879,N_6931,N_6359);
xnor U9880 (N_9880,N_5208,N_5537);
and U9881 (N_9881,N_5861,N_5358);
nand U9882 (N_9882,N_6960,N_6683);
nor U9883 (N_9883,N_6131,N_6394);
and U9884 (N_9884,N_7060,N_5199);
nand U9885 (N_9885,N_5256,N_6311);
nand U9886 (N_9886,N_6456,N_6532);
xor U9887 (N_9887,N_5173,N_6306);
nor U9888 (N_9888,N_6023,N_6381);
or U9889 (N_9889,N_7086,N_7105);
and U9890 (N_9890,N_7413,N_7100);
or U9891 (N_9891,N_6110,N_5547);
or U9892 (N_9892,N_6964,N_6461);
or U9893 (N_9893,N_5559,N_7183);
and U9894 (N_9894,N_6408,N_5214);
nand U9895 (N_9895,N_5353,N_6192);
and U9896 (N_9896,N_7475,N_6805);
and U9897 (N_9897,N_6823,N_7118);
nand U9898 (N_9898,N_7151,N_6477);
or U9899 (N_9899,N_6828,N_5828);
nor U9900 (N_9900,N_6295,N_5652);
nand U9901 (N_9901,N_5839,N_5026);
nor U9902 (N_9902,N_6230,N_6092);
nand U9903 (N_9903,N_6712,N_6700);
xor U9904 (N_9904,N_5361,N_6953);
nand U9905 (N_9905,N_5456,N_5759);
and U9906 (N_9906,N_6418,N_5838);
nor U9907 (N_9907,N_5256,N_6189);
nand U9908 (N_9908,N_6232,N_6024);
xnor U9909 (N_9909,N_5549,N_5651);
nand U9910 (N_9910,N_5576,N_6576);
nand U9911 (N_9911,N_5287,N_6327);
nand U9912 (N_9912,N_6405,N_6302);
or U9913 (N_9913,N_6751,N_6238);
nor U9914 (N_9914,N_6196,N_6337);
nor U9915 (N_9915,N_7374,N_5379);
nor U9916 (N_9916,N_5911,N_7429);
or U9917 (N_9917,N_6207,N_6789);
nor U9918 (N_9918,N_5667,N_5272);
nor U9919 (N_9919,N_5848,N_6176);
nor U9920 (N_9920,N_5973,N_7161);
nor U9921 (N_9921,N_5806,N_6301);
nand U9922 (N_9922,N_5334,N_6256);
nor U9923 (N_9923,N_5544,N_7139);
nor U9924 (N_9924,N_6506,N_7186);
nand U9925 (N_9925,N_7200,N_6544);
and U9926 (N_9926,N_7219,N_6696);
or U9927 (N_9927,N_5482,N_5096);
nand U9928 (N_9928,N_6339,N_5688);
xor U9929 (N_9929,N_5234,N_5996);
nand U9930 (N_9930,N_6628,N_5460);
or U9931 (N_9931,N_7136,N_6320);
or U9932 (N_9932,N_6203,N_6441);
or U9933 (N_9933,N_5353,N_5102);
nor U9934 (N_9934,N_7178,N_6677);
or U9935 (N_9935,N_5857,N_5564);
nand U9936 (N_9936,N_5854,N_5653);
or U9937 (N_9937,N_6701,N_5866);
xor U9938 (N_9938,N_6930,N_7298);
nand U9939 (N_9939,N_5996,N_5188);
nand U9940 (N_9940,N_5774,N_6892);
xor U9941 (N_9941,N_6448,N_7343);
nand U9942 (N_9942,N_6252,N_6495);
nand U9943 (N_9943,N_5956,N_6686);
nand U9944 (N_9944,N_5533,N_6851);
nand U9945 (N_9945,N_6837,N_5419);
and U9946 (N_9946,N_7140,N_5775);
nor U9947 (N_9947,N_6407,N_5843);
and U9948 (N_9948,N_5488,N_7089);
xnor U9949 (N_9949,N_7269,N_6588);
or U9950 (N_9950,N_6138,N_6181);
nand U9951 (N_9951,N_5752,N_5661);
xor U9952 (N_9952,N_5793,N_6868);
nor U9953 (N_9953,N_6727,N_5361);
and U9954 (N_9954,N_6925,N_6888);
xor U9955 (N_9955,N_5697,N_6593);
or U9956 (N_9956,N_5904,N_5493);
and U9957 (N_9957,N_7228,N_5219);
nor U9958 (N_9958,N_5123,N_6113);
nor U9959 (N_9959,N_7420,N_5334);
or U9960 (N_9960,N_5907,N_5170);
and U9961 (N_9961,N_7007,N_5159);
nor U9962 (N_9962,N_6689,N_6096);
nand U9963 (N_9963,N_7340,N_6181);
or U9964 (N_9964,N_6267,N_5529);
nor U9965 (N_9965,N_5057,N_5409);
xor U9966 (N_9966,N_7092,N_5652);
and U9967 (N_9967,N_6792,N_5344);
or U9968 (N_9968,N_6665,N_5889);
nand U9969 (N_9969,N_7254,N_5351);
nand U9970 (N_9970,N_5898,N_7496);
nand U9971 (N_9971,N_7448,N_5264);
and U9972 (N_9972,N_6924,N_6922);
nor U9973 (N_9973,N_7281,N_5455);
nor U9974 (N_9974,N_7346,N_5288);
or U9975 (N_9975,N_6316,N_6626);
or U9976 (N_9976,N_5434,N_5163);
or U9977 (N_9977,N_7243,N_5657);
nor U9978 (N_9978,N_6156,N_5192);
nand U9979 (N_9979,N_7097,N_5067);
nand U9980 (N_9980,N_5612,N_6358);
or U9981 (N_9981,N_6639,N_5888);
and U9982 (N_9982,N_5807,N_6438);
nor U9983 (N_9983,N_7426,N_5679);
nand U9984 (N_9984,N_6068,N_6498);
xnor U9985 (N_9985,N_6063,N_6165);
or U9986 (N_9986,N_5324,N_7475);
nor U9987 (N_9987,N_5603,N_5142);
nand U9988 (N_9988,N_6071,N_5221);
xor U9989 (N_9989,N_5352,N_5772);
or U9990 (N_9990,N_7441,N_5067);
and U9991 (N_9991,N_5593,N_6081);
or U9992 (N_9992,N_6888,N_5422);
and U9993 (N_9993,N_6102,N_5463);
nand U9994 (N_9994,N_6166,N_7212);
and U9995 (N_9995,N_5098,N_7406);
xnor U9996 (N_9996,N_6502,N_5333);
or U9997 (N_9997,N_6702,N_6342);
and U9998 (N_9998,N_6031,N_6957);
nor U9999 (N_9999,N_6957,N_6344);
xnor U10000 (N_10000,N_8557,N_8458);
nand U10001 (N_10001,N_9767,N_9626);
or U10002 (N_10002,N_8115,N_8112);
or U10003 (N_10003,N_7952,N_8298);
xnor U10004 (N_10004,N_9299,N_8377);
nand U10005 (N_10005,N_8305,N_8184);
or U10006 (N_10006,N_7662,N_8495);
nor U10007 (N_10007,N_9474,N_8652);
or U10008 (N_10008,N_7996,N_8380);
nor U10009 (N_10009,N_8438,N_7727);
xor U10010 (N_10010,N_9801,N_8259);
nand U10011 (N_10011,N_7531,N_7638);
nand U10012 (N_10012,N_9557,N_8101);
or U10013 (N_10013,N_8799,N_9857);
or U10014 (N_10014,N_8242,N_9333);
nor U10015 (N_10015,N_8856,N_8983);
nand U10016 (N_10016,N_8333,N_8464);
nor U10017 (N_10017,N_9391,N_7703);
nor U10018 (N_10018,N_8040,N_8805);
nor U10019 (N_10019,N_7873,N_8382);
or U10020 (N_10020,N_7676,N_9561);
or U10021 (N_10021,N_8780,N_7848);
and U10022 (N_10022,N_9027,N_7546);
nor U10023 (N_10023,N_9606,N_7717);
or U10024 (N_10024,N_7992,N_9736);
or U10025 (N_10025,N_9823,N_8054);
or U10026 (N_10026,N_9397,N_9347);
and U10027 (N_10027,N_9791,N_7850);
nor U10028 (N_10028,N_7965,N_9771);
nand U10029 (N_10029,N_7800,N_9264);
or U10030 (N_10030,N_9534,N_9167);
nor U10031 (N_10031,N_8939,N_9655);
xnor U10032 (N_10032,N_8467,N_8235);
and U10033 (N_10033,N_8700,N_8043);
nor U10034 (N_10034,N_8446,N_7766);
xnor U10035 (N_10035,N_7947,N_7978);
and U10036 (N_10036,N_7641,N_9796);
nor U10037 (N_10037,N_9505,N_8255);
or U10038 (N_10038,N_8973,N_9646);
nor U10039 (N_10039,N_8840,N_8689);
nand U10040 (N_10040,N_9401,N_8606);
nand U10041 (N_10041,N_9151,N_8186);
or U10042 (N_10042,N_9670,N_9853);
and U10043 (N_10043,N_7706,N_9128);
nand U10044 (N_10044,N_7645,N_8170);
nor U10045 (N_10045,N_7661,N_7558);
nor U10046 (N_10046,N_9974,N_7984);
nand U10047 (N_10047,N_8809,N_9331);
nand U10048 (N_10048,N_9122,N_8958);
nor U10049 (N_10049,N_9910,N_7514);
nor U10050 (N_10050,N_8474,N_8139);
xor U10051 (N_10051,N_8357,N_7583);
or U10052 (N_10052,N_8231,N_9781);
nand U10053 (N_10053,N_7935,N_7909);
and U10054 (N_10054,N_7521,N_7571);
xor U10055 (N_10055,N_7613,N_8618);
nand U10056 (N_10056,N_9118,N_9713);
or U10057 (N_10057,N_9984,N_9133);
and U10058 (N_10058,N_9916,N_9101);
xnor U10059 (N_10059,N_9111,N_7806);
nand U10060 (N_10060,N_7842,N_7633);
xor U10061 (N_10061,N_9669,N_8472);
nand U10062 (N_10062,N_9918,N_7520);
and U10063 (N_10063,N_9997,N_8179);
or U10064 (N_10064,N_8007,N_7937);
nand U10065 (N_10065,N_9892,N_9532);
xnor U10066 (N_10066,N_7787,N_8926);
nand U10067 (N_10067,N_9510,N_8715);
nor U10068 (N_10068,N_9661,N_8120);
and U10069 (N_10069,N_7733,N_7642);
or U10070 (N_10070,N_9051,N_8864);
and U10071 (N_10071,N_8641,N_7559);
and U10072 (N_10072,N_8642,N_7925);
nor U10073 (N_10073,N_8345,N_9642);
nand U10074 (N_10074,N_7589,N_9224);
or U10075 (N_10075,N_9737,N_9280);
or U10076 (N_10076,N_8267,N_9019);
nand U10077 (N_10077,N_7643,N_7818);
nor U10078 (N_10078,N_7674,N_8005);
nor U10079 (N_10079,N_9537,N_9748);
nor U10080 (N_10080,N_8589,N_9012);
or U10081 (N_10081,N_9536,N_8702);
or U10082 (N_10082,N_9867,N_7636);
or U10083 (N_10083,N_7757,N_8743);
and U10084 (N_10084,N_9378,N_8424);
nand U10085 (N_10085,N_9888,N_9763);
nand U10086 (N_10086,N_8251,N_9805);
nand U10087 (N_10087,N_7913,N_7914);
nor U10088 (N_10088,N_8315,N_8624);
or U10089 (N_10089,N_8062,N_8526);
nor U10090 (N_10090,N_8127,N_9973);
nor U10091 (N_10091,N_7808,N_7711);
nand U10092 (N_10092,N_8519,N_7623);
and U10093 (N_10093,N_8297,N_9475);
nand U10094 (N_10094,N_8797,N_8503);
and U10095 (N_10095,N_9462,N_8277);
or U10096 (N_10096,N_9869,N_9899);
and U10097 (N_10097,N_9950,N_8901);
nor U10098 (N_10098,N_8717,N_8143);
nor U10099 (N_10099,N_7955,N_9086);
nor U10100 (N_10100,N_9559,N_8793);
nor U10101 (N_10101,N_9449,N_8020);
nand U10102 (N_10102,N_9184,N_8528);
and U10103 (N_10103,N_8826,N_9949);
and U10104 (N_10104,N_7905,N_7501);
or U10105 (N_10105,N_8336,N_8321);
and U10106 (N_10106,N_9589,N_8417);
nor U10107 (N_10107,N_8065,N_8951);
or U10108 (N_10108,N_9928,N_7904);
nand U10109 (N_10109,N_9202,N_9564);
nand U10110 (N_10110,N_8655,N_9554);
nand U10111 (N_10111,N_7513,N_9526);
nand U10112 (N_10112,N_9100,N_9487);
nand U10113 (N_10113,N_9313,N_7874);
and U10114 (N_10114,N_9188,N_8995);
xnor U10115 (N_10115,N_8310,N_9567);
or U10116 (N_10116,N_8484,N_9324);
or U10117 (N_10117,N_9983,N_8631);
or U10118 (N_10118,N_8434,N_8969);
xor U10119 (N_10119,N_8736,N_8612);
nor U10120 (N_10120,N_9990,N_7619);
nand U10121 (N_10121,N_8220,N_8695);
and U10122 (N_10122,N_8447,N_8905);
nand U10123 (N_10123,N_9067,N_9206);
xor U10124 (N_10124,N_7979,N_7756);
or U10125 (N_10125,N_9193,N_8899);
or U10126 (N_10126,N_9915,N_7672);
nor U10127 (N_10127,N_8749,N_8018);
or U10128 (N_10128,N_9677,N_8422);
and U10129 (N_10129,N_8930,N_7958);
or U10130 (N_10130,N_7902,N_9760);
or U10131 (N_10131,N_8111,N_7612);
or U10132 (N_10132,N_7760,N_9925);
nor U10133 (N_10133,N_8138,N_7987);
nor U10134 (N_10134,N_9993,N_8405);
and U10135 (N_10135,N_8896,N_8756);
nor U10136 (N_10136,N_7765,N_7886);
nand U10137 (N_10137,N_7741,N_9129);
nand U10138 (N_10138,N_9405,N_8376);
nor U10139 (N_10139,N_7737,N_9229);
nand U10140 (N_10140,N_8466,N_9852);
and U10141 (N_10141,N_8217,N_7782);
nor U10142 (N_10142,N_7567,N_9788);
and U10143 (N_10143,N_9750,N_9587);
nand U10144 (N_10144,N_9716,N_7596);
or U10145 (N_10145,N_7562,N_8802);
nand U10146 (N_10146,N_7815,N_8497);
and U10147 (N_10147,N_9131,N_8538);
xnor U10148 (N_10148,N_7933,N_7863);
and U10149 (N_10149,N_7582,N_9302);
xor U10150 (N_10150,N_7595,N_9814);
nor U10151 (N_10151,N_8868,N_9436);
and U10152 (N_10152,N_8600,N_7893);
nor U10153 (N_10153,N_9211,N_8089);
or U10154 (N_10154,N_8863,N_8762);
nor U10155 (N_10155,N_9595,N_9138);
nand U10156 (N_10156,N_9515,N_7670);
nand U10157 (N_10157,N_7993,N_8692);
and U10158 (N_10158,N_9624,N_7812);
nor U10159 (N_10159,N_7616,N_8653);
and U10160 (N_10160,N_9701,N_7780);
nor U10161 (N_10161,N_7659,N_8694);
nand U10162 (N_10162,N_9715,N_9318);
nor U10163 (N_10163,N_9776,N_8122);
nor U10164 (N_10164,N_9247,N_7897);
and U10165 (N_10165,N_9008,N_7836);
and U10166 (N_10166,N_8857,N_8979);
nand U10167 (N_10167,N_9797,N_9360);
nand U10168 (N_10168,N_9268,N_9733);
and U10169 (N_10169,N_9039,N_9478);
xnor U10170 (N_10170,N_8437,N_9428);
xnor U10171 (N_10171,N_8831,N_9619);
nand U10172 (N_10172,N_7827,N_7868);
and U10173 (N_10173,N_9614,N_9802);
nand U10174 (N_10174,N_8704,N_9375);
nand U10175 (N_10175,N_8536,N_9006);
xnor U10176 (N_10176,N_9519,N_8788);
and U10177 (N_10177,N_7885,N_8019);
nand U10178 (N_10178,N_9352,N_7627);
or U10179 (N_10179,N_8927,N_8426);
xnor U10180 (N_10180,N_9231,N_9696);
and U10181 (N_10181,N_8427,N_9967);
nand U10182 (N_10182,N_7668,N_8287);
or U10183 (N_10183,N_8292,N_9568);
nand U10184 (N_10184,N_8583,N_9469);
or U10185 (N_10185,N_9647,N_8892);
or U10186 (N_10186,N_9609,N_9205);
nand U10187 (N_10187,N_8064,N_8657);
nor U10188 (N_10188,N_7934,N_8032);
and U10189 (N_10189,N_7994,N_8946);
nor U10190 (N_10190,N_7660,N_8888);
nand U10191 (N_10191,N_7912,N_7986);
or U10192 (N_10192,N_8705,N_8090);
and U10193 (N_10193,N_9290,N_8279);
nand U10194 (N_10194,N_7862,N_9803);
or U10195 (N_10195,N_8693,N_9832);
xor U10196 (N_10196,N_9022,N_9693);
nand U10197 (N_10197,N_9521,N_8532);
nand U10198 (N_10198,N_9402,N_9522);
nor U10199 (N_10199,N_8140,N_9187);
nand U10200 (N_10200,N_9107,N_7511);
and U10201 (N_10201,N_8714,N_7607);
nand U10202 (N_10202,N_9682,N_8900);
or U10203 (N_10203,N_9908,N_8052);
nor U10204 (N_10204,N_8258,N_9769);
and U10205 (N_10205,N_8387,N_8911);
and U10206 (N_10206,N_9999,N_9090);
nand U10207 (N_10207,N_9198,N_9203);
xnor U10208 (N_10208,N_7924,N_8419);
and U10209 (N_10209,N_8825,N_8859);
nand U10210 (N_10210,N_9981,N_8713);
or U10211 (N_10211,N_9387,N_8605);
nand U10212 (N_10212,N_7508,N_9498);
xor U10213 (N_10213,N_9450,N_9488);
nor U10214 (N_10214,N_8325,N_8485);
xnor U10215 (N_10215,N_9467,N_9923);
nand U10216 (N_10216,N_8151,N_8607);
nand U10217 (N_10217,N_8662,N_7995);
nand U10218 (N_10218,N_8529,N_7651);
or U10219 (N_10219,N_7680,N_9394);
nand U10220 (N_10220,N_9335,N_9125);
nor U10221 (N_10221,N_8520,N_8081);
nand U10222 (N_10222,N_8209,N_9599);
or U10223 (N_10223,N_7910,N_9062);
nand U10224 (N_10224,N_7870,N_9702);
nor U10225 (N_10225,N_9728,N_8031);
nand U10226 (N_10226,N_9127,N_9607);
or U10227 (N_10227,N_9798,N_7991);
and U10228 (N_10228,N_9884,N_9328);
and U10229 (N_10229,N_7802,N_9858);
xnor U10230 (N_10230,N_8431,N_8898);
nand U10231 (N_10231,N_9476,N_9720);
xor U10232 (N_10232,N_9691,N_9905);
and U10233 (N_10233,N_8820,N_8861);
nor U10234 (N_10234,N_7655,N_7683);
and U10235 (N_10235,N_9850,N_8211);
or U10236 (N_10236,N_9639,N_9348);
nand U10237 (N_10237,N_8636,N_9860);
nor U10238 (N_10238,N_9301,N_9263);
or U10239 (N_10239,N_9085,N_9708);
nand U10240 (N_10240,N_8142,N_8411);
xnor U10241 (N_10241,N_9004,N_8439);
nor U10242 (N_10242,N_9033,N_7517);
xnor U10243 (N_10243,N_8066,N_7795);
nand U10244 (N_10244,N_7872,N_9373);
and U10245 (N_10245,N_8056,N_8649);
nand U10246 (N_10246,N_8171,N_9944);
and U10247 (N_10247,N_9018,N_9800);
nor U10248 (N_10248,N_9779,N_8522);
and U10249 (N_10249,N_9835,N_9902);
nand U10250 (N_10250,N_9755,N_8643);
nand U10251 (N_10251,N_8674,N_7628);
nand U10252 (N_10252,N_8506,N_7677);
and U10253 (N_10253,N_9966,N_8669);
nor U10254 (N_10254,N_8402,N_9920);
and U10255 (N_10255,N_7981,N_8391);
nand U10256 (N_10256,N_8807,N_7743);
nand U10257 (N_10257,N_8549,N_9730);
or U10258 (N_10258,N_8912,N_9023);
or U10259 (N_10259,N_7763,N_8579);
and U10260 (N_10260,N_8189,N_7775);
xnor U10261 (N_10261,N_8765,N_8099);
nor U10262 (N_10262,N_8625,N_7832);
nand U10263 (N_10263,N_7844,N_7723);
nor U10264 (N_10264,N_9729,N_8188);
nand U10265 (N_10265,N_9811,N_8457);
xnor U10266 (N_10266,N_7752,N_8317);
xnor U10267 (N_10267,N_8415,N_9010);
and U10268 (N_10268,N_8542,N_8916);
and U10269 (N_10269,N_9441,N_9180);
nand U10270 (N_10270,N_9117,N_7681);
nand U10271 (N_10271,N_9177,N_8950);
or U10272 (N_10272,N_7635,N_8903);
nor U10273 (N_10273,N_8313,N_9270);
nor U10274 (N_10274,N_7579,N_9414);
xnor U10275 (N_10275,N_8449,N_8275);
and U10276 (N_10276,N_9271,N_7669);
and U10277 (N_10277,N_9723,N_8119);
nor U10278 (N_10278,N_8162,N_9765);
nor U10279 (N_10279,N_7860,N_8760);
nor U10280 (N_10280,N_8319,N_9453);
and U10281 (N_10281,N_8897,N_7930);
nor U10282 (N_10282,N_7799,N_7658);
and U10283 (N_10283,N_9372,N_7997);
nor U10284 (N_10284,N_9120,N_8830);
or U10285 (N_10285,N_9643,N_9032);
nor U10286 (N_10286,N_7900,N_9024);
and U10287 (N_10287,N_9204,N_8568);
and U10288 (N_10288,N_9346,N_7888);
nand U10289 (N_10289,N_9078,N_8726);
xnor U10290 (N_10290,N_9057,N_8751);
xnor U10291 (N_10291,N_8400,N_8410);
and U10292 (N_10292,N_8029,N_7915);
nor U10293 (N_10293,N_9410,N_9936);
and U10294 (N_10294,N_9512,N_8306);
nor U10295 (N_10295,N_8114,N_9278);
or U10296 (N_10296,N_8679,N_7788);
nor U10297 (N_10297,N_9717,N_9049);
nand U10298 (N_10298,N_8499,N_9645);
nor U10299 (N_10299,N_8786,N_9196);
nand U10300 (N_10300,N_9074,N_8635);
and U10301 (N_10301,N_8491,N_7957);
or U10302 (N_10302,N_9272,N_9239);
and U10303 (N_10303,N_8517,N_7881);
or U10304 (N_10304,N_7887,N_7895);
xor U10305 (N_10305,N_7772,N_8902);
nand U10306 (N_10306,N_7774,N_8664);
nand U10307 (N_10307,N_8226,N_8650);
nor U10308 (N_10308,N_8147,N_8166);
and U10309 (N_10309,N_7576,N_9060);
or U10310 (N_10310,N_8048,N_7715);
or U10311 (N_10311,N_8565,N_8659);
or U10312 (N_10312,N_9236,N_8378);
nand U10313 (N_10313,N_8369,N_9444);
or U10314 (N_10314,N_8878,N_8671);
or U10315 (N_10315,N_8634,N_9274);
nand U10316 (N_10316,N_9491,N_7983);
nor U10317 (N_10317,N_9257,N_9005);
nand U10318 (N_10318,N_9254,N_8891);
or U10319 (N_10319,N_8124,N_9460);
or U10320 (N_10320,N_8721,N_9273);
or U10321 (N_10321,N_7804,N_9759);
and U10322 (N_10322,N_9931,N_8706);
nor U10323 (N_10323,N_8362,N_7523);
or U10324 (N_10324,N_9831,N_7516);
or U10325 (N_10325,N_9116,N_8853);
and U10326 (N_10326,N_9359,N_7610);
or U10327 (N_10327,N_7929,N_9115);
and U10328 (N_10328,N_7569,N_9849);
and U10329 (N_10329,N_7691,N_8551);
and U10330 (N_10330,N_8489,N_9937);
xnor U10331 (N_10331,N_8398,N_9790);
nand U10332 (N_10332,N_8510,N_8307);
and U10333 (N_10333,N_9139,N_7649);
nand U10334 (N_10334,N_8294,N_9921);
or U10335 (N_10335,N_9199,N_9584);
nor U10336 (N_10336,N_7949,N_9575);
or U10337 (N_10337,N_9287,N_9745);
or U10338 (N_10338,N_8680,N_7809);
xnor U10339 (N_10339,N_9473,N_9617);
or U10340 (N_10340,N_9421,N_9873);
or U10341 (N_10341,N_7625,N_7586);
nand U10342 (N_10342,N_8418,N_8546);
nand U10343 (N_10343,N_9846,N_7573);
and U10344 (N_10344,N_7506,N_9106);
and U10345 (N_10345,N_7578,N_8597);
xnor U10346 (N_10346,N_8085,N_8573);
xnor U10347 (N_10347,N_8097,N_7530);
and U10348 (N_10348,N_9709,N_9223);
nand U10349 (N_10349,N_7877,N_8036);
or U10350 (N_10350,N_8813,N_8794);
nand U10351 (N_10351,N_8594,N_7859);
nand U10352 (N_10352,N_8789,N_8455);
nand U10353 (N_10353,N_9636,N_9293);
nor U10354 (N_10354,N_9020,N_9784);
or U10355 (N_10355,N_8823,N_9511);
or U10356 (N_10356,N_7847,N_7807);
nor U10357 (N_10357,N_8534,N_8544);
and U10358 (N_10358,N_9212,N_9663);
and U10359 (N_10359,N_8326,N_7906);
and U10360 (N_10360,N_9149,N_9687);
nor U10361 (N_10361,N_9448,N_7563);
nand U10362 (N_10362,N_8723,N_9563);
and U10363 (N_10363,N_7745,N_9897);
or U10364 (N_10364,N_8962,N_9146);
or U10365 (N_10365,N_7833,N_8356);
nand U10366 (N_10366,N_9031,N_8957);
xor U10367 (N_10367,N_9425,N_8476);
nor U10368 (N_10368,N_8207,N_9267);
nand U10369 (N_10369,N_9666,N_9392);
or U10370 (N_10370,N_8498,N_8895);
and U10371 (N_10371,N_9089,N_8027);
or U10372 (N_10372,N_9598,N_9909);
nand U10373 (N_10373,N_7843,N_8541);
xor U10374 (N_10374,N_8550,N_9845);
xnor U10375 (N_10375,N_8963,N_8164);
or U10376 (N_10376,N_9068,N_9256);
and U10377 (N_10377,N_9063,N_9685);
xor U10378 (N_10378,N_8390,N_8562);
xnor U10379 (N_10379,N_8985,N_8365);
nor U10380 (N_10380,N_8450,N_9757);
and U10381 (N_10381,N_9746,N_8639);
nand U10382 (N_10382,N_9383,N_9314);
nor U10383 (N_10383,N_9652,N_8215);
or U10384 (N_10384,N_8684,N_9230);
and U10385 (N_10385,N_8569,N_8701);
or U10386 (N_10386,N_7725,N_7656);
and U10387 (N_10387,N_7713,N_8144);
nand U10388 (N_10388,N_9623,N_7555);
nor U10389 (N_10389,N_9906,N_7601);
nor U10390 (N_10390,N_8848,N_9839);
nor U10391 (N_10391,N_7851,N_7923);
nand U10392 (N_10392,N_8192,N_8137);
and U10393 (N_10393,N_8212,N_8224);
nand U10394 (N_10394,N_7608,N_8953);
nand U10395 (N_10395,N_9471,N_9468);
and U10396 (N_10396,N_7797,N_9385);
or U10397 (N_10397,N_9114,N_9756);
and U10398 (N_10398,N_8197,N_7742);
or U10399 (N_10399,N_8708,N_9732);
or U10400 (N_10400,N_8168,N_9459);
or U10401 (N_10401,N_9964,N_8205);
and U10402 (N_10402,N_9150,N_8332);
and U10403 (N_10403,N_9369,N_8015);
and U10404 (N_10404,N_8854,N_7942);
nand U10405 (N_10405,N_8955,N_9155);
nand U10406 (N_10406,N_9484,N_9251);
nor U10407 (N_10407,N_8533,N_9870);
nor U10408 (N_10408,N_8250,N_8564);
nor U10409 (N_10409,N_8118,N_8158);
and U10410 (N_10410,N_9226,N_8022);
and U10411 (N_10411,N_9327,N_9248);
or U10412 (N_10412,N_8525,N_7554);
nor U10413 (N_10413,N_9282,N_8844);
nor U10414 (N_10414,N_9573,N_9795);
and U10415 (N_10415,N_7789,N_7729);
nand U10416 (N_10416,N_7816,N_7572);
and U10417 (N_10417,N_8910,N_8774);
nor U10418 (N_10418,N_9593,N_9817);
and U10419 (N_10419,N_9946,N_7747);
nand U10420 (N_10420,N_9844,N_8913);
or U10421 (N_10421,N_9935,N_8894);
nor U10422 (N_10422,N_7819,N_8604);
or U10423 (N_10423,N_8682,N_9043);
nand U10424 (N_10424,N_9426,N_7899);
nor U10425 (N_10425,N_8656,N_7716);
nand U10426 (N_10426,N_9000,N_8075);
xor U10427 (N_10427,N_9349,N_9485);
nand U10428 (N_10428,N_9424,N_9955);
xor U10429 (N_10429,N_8136,N_9657);
and U10430 (N_10430,N_7545,N_7931);
nor U10431 (N_10431,N_9588,N_9523);
nor U10432 (N_10432,N_8967,N_9434);
nor U10433 (N_10433,N_9700,N_9040);
nor U10434 (N_10434,N_8026,N_8234);
nor U10435 (N_10435,N_8271,N_9770);
nand U10436 (N_10436,N_8874,N_8595);
nand U10437 (N_10437,N_9939,N_8886);
xnor U10438 (N_10438,N_9752,N_8976);
and U10439 (N_10439,N_7695,N_8560);
and U10440 (N_10440,N_8312,N_9680);
and U10441 (N_10441,N_7823,N_8672);
nand U10442 (N_10442,N_9914,N_9056);
nand U10443 (N_10443,N_9061,N_9244);
or U10444 (N_10444,N_7961,N_8069);
or U10445 (N_10445,N_9225,N_8592);
nor U10446 (N_10446,N_8578,N_9017);
nand U10447 (N_10447,N_7866,N_7820);
and U10448 (N_10448,N_8198,N_8688);
nor U10449 (N_10449,N_8938,N_7693);
and U10450 (N_10450,N_8993,N_7730);
nand U10451 (N_10451,N_8004,N_9079);
nand U10452 (N_10452,N_8727,N_8909);
and U10453 (N_10453,N_8385,N_8448);
nor U10454 (N_10454,N_9152,N_7810);
xnor U10455 (N_10455,N_8556,N_8816);
nand U10456 (N_10456,N_9241,N_9618);
nand U10457 (N_10457,N_8616,N_9605);
or U10458 (N_10458,N_8096,N_8436);
and U10459 (N_10459,N_9296,N_7564);
or U10460 (N_10460,N_7911,N_8998);
and U10461 (N_10461,N_8673,N_8862);
or U10462 (N_10462,N_8965,N_8165);
nor U10463 (N_10463,N_8923,N_7710);
nor U10464 (N_10464,N_7647,N_7654);
and U10465 (N_10465,N_9137,N_8406);
xor U10466 (N_10466,N_8614,N_8442);
xor U10467 (N_10467,N_9092,N_8936);
nand U10468 (N_10468,N_8948,N_7507);
and U10469 (N_10469,N_8473,N_9095);
nor U10470 (N_10470,N_9456,N_7939);
or U10471 (N_10471,N_9253,N_9075);
nand U10472 (N_10472,N_9953,N_8766);
xor U10473 (N_10473,N_7726,N_8470);
xor U10474 (N_10474,N_8545,N_8626);
nor U10475 (N_10475,N_9665,N_8527);
nand U10476 (N_10476,N_7549,N_8591);
or U10477 (N_10477,N_9259,N_9130);
nand U10478 (N_10478,N_7544,N_8091);
nor U10479 (N_10479,N_9896,N_9200);
xor U10480 (N_10480,N_9013,N_8709);
nor U10481 (N_10481,N_8735,N_8157);
and U10482 (N_10482,N_8086,N_8918);
or U10483 (N_10483,N_8960,N_8225);
nor U10484 (N_10484,N_8232,N_8747);
nand U10485 (N_10485,N_8429,N_7560);
nor U10486 (N_10486,N_9439,N_8451);
xor U10487 (N_10487,N_7731,N_8462);
or U10488 (N_10488,N_9361,N_8580);
nor U10489 (N_10489,N_8353,N_9735);
nand U10490 (N_10490,N_7878,N_8346);
nor U10491 (N_10491,N_7689,N_8291);
nand U10492 (N_10492,N_7783,N_9119);
nor U10493 (N_10493,N_7526,N_8057);
or U10494 (N_10494,N_9055,N_9093);
nor U10495 (N_10495,N_8264,N_8053);
nand U10496 (N_10496,N_8453,N_9160);
nor U10497 (N_10497,N_9875,N_7998);
xnor U10498 (N_10498,N_8340,N_7980);
nand U10499 (N_10499,N_7781,N_9166);
nor U10500 (N_10500,N_7951,N_9653);
xor U10501 (N_10501,N_9629,N_8722);
or U10502 (N_10502,N_9651,N_9810);
nor U10503 (N_10503,N_7550,N_9430);
or U10504 (N_10504,N_9613,N_9398);
nor U10505 (N_10505,N_8515,N_8129);
or U10506 (N_10506,N_7945,N_9183);
and U10507 (N_10507,N_7543,N_7896);
xor U10508 (N_10508,N_8237,N_8288);
and U10509 (N_10509,N_8195,N_7841);
nand U10510 (N_10510,N_8024,N_7598);
nor U10511 (N_10511,N_7667,N_9097);
or U10512 (N_10512,N_9047,N_9514);
nor U10513 (N_10513,N_8553,N_8133);
or U10514 (N_10514,N_9232,N_9978);
and U10515 (N_10515,N_8403,N_7972);
nand U10516 (N_10516,N_7966,N_7751);
and U10517 (N_10517,N_7719,N_8163);
nor U10518 (N_10518,N_8640,N_7974);
or U10519 (N_10519,N_9942,N_9841);
or U10520 (N_10520,N_7570,N_9157);
nand U10521 (N_10521,N_9374,N_9604);
or U10522 (N_10522,N_7675,N_9866);
xnor U10523 (N_10523,N_9011,N_8567);
xor U10524 (N_10524,N_8272,N_9099);
or U10525 (N_10525,N_8563,N_9214);
nand U10526 (N_10526,N_8349,N_9726);
and U10527 (N_10527,N_8351,N_8046);
and U10528 (N_10528,N_7814,N_7664);
or U10529 (N_10529,N_7694,N_8102);
and U10530 (N_10530,N_7876,N_8731);
or U10531 (N_10531,N_8461,N_9066);
or U10532 (N_10532,N_8219,N_7614);
nand U10533 (N_10533,N_9321,N_7944);
and U10534 (N_10534,N_9859,N_8008);
nand U10535 (N_10535,N_9812,N_9390);
and U10536 (N_10536,N_8956,N_8608);
nand U10537 (N_10537,N_9281,N_9822);
and U10538 (N_10538,N_9038,N_7518);
and U10539 (N_10539,N_8992,N_9582);
nor U10540 (N_10540,N_7999,N_8044);
xor U10541 (N_10541,N_8284,N_8530);
or U10542 (N_10542,N_8392,N_8238);
nor U10543 (N_10543,N_8698,N_9364);
and U10544 (N_10544,N_9344,N_8987);
nor U10545 (N_10545,N_8877,N_8981);
or U10546 (N_10546,N_8176,N_8227);
and U10547 (N_10547,N_9353,N_9929);
and U10548 (N_10548,N_7976,N_7967);
xor U10549 (N_10549,N_9134,N_8080);
nor U10550 (N_10550,N_7852,N_8621);
and U10551 (N_10551,N_7853,N_9317);
xnor U10552 (N_10552,N_8038,N_8633);
and U10553 (N_10553,N_8931,N_9638);
nor U10554 (N_10554,N_9217,N_9110);
or U10555 (N_10555,N_9890,N_9419);
or U10556 (N_10556,N_9276,N_7988);
nand U10557 (N_10557,N_9601,N_8683);
nor U10558 (N_10558,N_8444,N_9208);
nand U10559 (N_10559,N_7792,N_7500);
and U10560 (N_10560,N_9690,N_8174);
xnor U10561 (N_10561,N_8773,N_8098);
nand U10562 (N_10562,N_9833,N_9179);
nor U10563 (N_10563,N_7556,N_8566);
and U10564 (N_10564,N_9876,N_8827);
or U10565 (N_10565,N_8929,N_9201);
and U10566 (N_10566,N_8504,N_9098);
nand U10567 (N_10567,N_8991,N_7846);
or U10568 (N_10568,N_9783,N_8665);
or U10569 (N_10569,N_9034,N_8984);
xnor U10570 (N_10570,N_8460,N_8710);
nor U10571 (N_10571,N_9773,N_7519);
or U10572 (N_10572,N_9913,N_8216);
nor U10573 (N_10573,N_9124,N_9940);
or U10574 (N_10574,N_8134,N_9332);
and U10575 (N_10575,N_8421,N_8601);
and U10576 (N_10576,N_9297,N_8475);
and U10577 (N_10577,N_9102,N_8067);
or U10578 (N_10578,N_9504,N_7840);
nor U10579 (N_10579,N_7697,N_8304);
nor U10580 (N_10580,N_8374,N_9615);
nor U10581 (N_10581,N_9894,N_8666);
nor U10582 (N_10582,N_9042,N_9751);
and U10583 (N_10583,N_8210,N_9807);
xnor U10584 (N_10584,N_7754,N_7907);
or U10585 (N_10585,N_9874,N_9530);
nor U10586 (N_10586,N_8070,N_8161);
nor U10587 (N_10587,N_8359,N_7960);
or U10588 (N_10588,N_9104,N_8107);
and U10589 (N_10589,N_9911,N_9258);
or U10590 (N_10590,N_9135,N_7696);
nor U10591 (N_10591,N_8443,N_8615);
and U10592 (N_10592,N_8884,N_9540);
xor U10593 (N_10593,N_7620,N_8074);
nor U10594 (N_10594,N_9243,N_8246);
and U10595 (N_10595,N_8087,N_7515);
or U10596 (N_10596,N_9379,N_9722);
nor U10597 (N_10597,N_9501,N_8554);
nor U10598 (N_10598,N_8034,N_8869);
nor U10599 (N_10599,N_9171,N_8971);
nand U10600 (N_10600,N_9877,N_9574);
nor U10601 (N_10601,N_8035,N_8257);
and U10602 (N_10602,N_8806,N_8574);
nand U10603 (N_10603,N_9064,N_9775);
or U10604 (N_10604,N_9627,N_7920);
and U10605 (N_10605,N_8030,N_8845);
nor U10606 (N_10606,N_8331,N_8879);
xor U10607 (N_10607,N_9286,N_8808);
nor U10608 (N_10608,N_9422,N_9793);
nand U10609 (N_10609,N_9819,N_9576);
or U10610 (N_10610,N_9932,N_7786);
and U10611 (N_10611,N_8228,N_9602);
xor U10612 (N_10612,N_9986,N_9987);
nand U10613 (N_10613,N_8803,N_9612);
and U10614 (N_10614,N_7682,N_8887);
nand U10615 (N_10615,N_9592,N_9048);
and U10616 (N_10616,N_9265,N_7884);
nand U10617 (N_10617,N_7824,N_7584);
nand U10618 (N_10618,N_8344,N_8493);
nor U10619 (N_10619,N_9185,N_8882);
or U10620 (N_10620,N_8829,N_8818);
nor U10621 (N_10621,N_9965,N_7634);
and U10622 (N_10622,N_9749,N_8465);
or U10623 (N_10623,N_9956,N_9458);
or U10624 (N_10624,N_9957,N_9934);
or U10625 (N_10625,N_8949,N_8408);
nor U10626 (N_10626,N_8095,N_8758);
or U10627 (N_10627,N_9865,N_8757);
and U10628 (N_10628,N_7502,N_9404);
nand U10629 (N_10629,N_9052,N_7791);
nor U10630 (N_10630,N_9041,N_7509);
nand U10631 (N_10631,N_8796,N_9816);
or U10632 (N_10632,N_7959,N_9380);
and U10633 (N_10633,N_8964,N_9235);
or U10634 (N_10634,N_7605,N_7505);
nand U10635 (N_10635,N_9969,N_9648);
and U10636 (N_10636,N_8972,N_9671);
nand U10637 (N_10637,N_7954,N_7522);
or U10638 (N_10638,N_9632,N_9996);
or U10639 (N_10639,N_8941,N_8646);
or U10640 (N_10640,N_8347,N_8302);
or U10641 (N_10641,N_9650,N_9933);
or U10642 (N_10642,N_9863,N_8016);
or U10643 (N_10643,N_9734,N_9109);
nand U10644 (N_10644,N_8182,N_7773);
or U10645 (N_10645,N_9555,N_9142);
nand U10646 (N_10646,N_8837,N_9579);
or U10647 (N_10647,N_8539,N_8183);
nand U10648 (N_10648,N_9780,N_9323);
nor U10649 (N_10649,N_9371,N_8480);
nand U10650 (N_10650,N_7685,N_8593);
nand U10651 (N_10651,N_9334,N_9195);
or U10652 (N_10652,N_9249,N_9662);
nand U10653 (N_10653,N_7950,N_8083);
nand U10654 (N_10654,N_8017,N_8988);
and U10655 (N_10655,N_9679,N_7835);
nor U10656 (N_10656,N_9881,N_8610);
and U10657 (N_10657,N_9848,N_9727);
xnor U10658 (N_10658,N_8740,N_9084);
or U10659 (N_10659,N_8883,N_8433);
or U10660 (N_10660,N_9053,N_9963);
nand U10661 (N_10661,N_9143,N_8552);
xnor U10662 (N_10662,N_7503,N_7621);
nor U10663 (N_10663,N_7587,N_8501);
nand U10664 (N_10664,N_8678,N_8925);
and U10665 (N_10665,N_9820,N_9316);
or U10666 (N_10666,N_7541,N_9191);
or U10667 (N_10667,N_9399,N_9705);
nand U10668 (N_10668,N_8088,N_8667);
nand U10669 (N_10669,N_8935,N_9156);
nand U10670 (N_10670,N_8716,N_7796);
and U10671 (N_10671,N_8921,N_8543);
nand U10672 (N_10672,N_8523,N_8072);
and U10673 (N_10673,N_9164,N_9220);
nand U10674 (N_10674,N_7561,N_8954);
and U10675 (N_10675,N_8286,N_9562);
nand U10676 (N_10676,N_9368,N_9855);
nor U10677 (N_10677,N_7592,N_8328);
or U10678 (N_10678,N_8777,N_8974);
nand U10679 (N_10679,N_7982,N_7750);
nor U10680 (N_10680,N_7617,N_8880);
or U10681 (N_10681,N_9288,N_8860);
or U10682 (N_10682,N_8875,N_9416);
and U10683 (N_10683,N_9976,N_8637);
or U10684 (N_10684,N_8423,N_8452);
and U10685 (N_10685,N_9329,N_9919);
nor U10686 (N_10686,N_8617,N_7856);
nor U10687 (N_10687,N_8596,N_9420);
nand U10688 (N_10688,N_9945,N_7889);
xnor U10689 (N_10689,N_8093,N_9586);
and U10690 (N_10690,N_7834,N_8441);
nand U10691 (N_10691,N_9695,N_9294);
nor U10692 (N_10692,N_8603,N_7532);
nor U10693 (N_10693,N_8430,N_9707);
xnor U10694 (N_10694,N_7692,N_9002);
and U10695 (N_10695,N_7580,N_8980);
nand U10696 (N_10696,N_8841,N_8511);
or U10697 (N_10697,N_7749,N_8335);
nand U10698 (N_10698,N_9457,N_8940);
nor U10699 (N_10699,N_9437,N_9738);
and U10700 (N_10700,N_9303,N_8194);
and U10701 (N_10701,N_8047,N_9872);
nand U10702 (N_10702,N_9227,N_8628);
or U10703 (N_10703,N_9871,N_8367);
nand U10704 (N_10704,N_9774,N_7857);
nand U10705 (N_10705,N_8668,N_9186);
nand U10706 (N_10706,N_9431,N_9058);
nor U10707 (N_10707,N_9503,N_9351);
nor U10708 (N_10708,N_9172,N_9952);
nand U10709 (N_10709,N_8368,N_7728);
and U10710 (N_10710,N_9544,N_9461);
nand U10711 (N_10711,N_8759,N_7714);
or U10712 (N_10712,N_8748,N_8045);
or U10713 (N_10713,N_8050,N_7890);
and U10714 (N_10714,N_8658,N_8753);
xor U10715 (N_10715,N_9088,N_9815);
and U10716 (N_10716,N_9003,N_9423);
and U10717 (N_10717,N_8274,N_8812);
nand U10718 (N_10718,N_7811,N_9350);
xnor U10719 (N_10719,N_9178,N_8505);
xor U10720 (N_10720,N_7588,N_9408);
nor U10721 (N_10721,N_8320,N_8815);
nor U10722 (N_10722,N_9080,N_9417);
nor U10723 (N_10723,N_9778,N_7637);
nand U10724 (N_10724,N_8076,N_8890);
nor U10725 (N_10725,N_8432,N_7700);
xor U10726 (N_10726,N_7539,N_8490);
nand U10727 (N_10727,N_7948,N_8558);
nor U10728 (N_10728,N_8502,N_9782);
nor U10729 (N_10729,N_9527,N_7552);
and U10730 (N_10730,N_7956,N_9889);
nand U10731 (N_10731,N_7648,N_9985);
nand U10732 (N_10732,N_7603,N_8947);
and U10733 (N_10733,N_7753,N_9363);
nand U10734 (N_10734,N_7712,N_7946);
nor U10735 (N_10735,N_9283,N_9077);
nand U10736 (N_10736,N_8477,N_9250);
and U10737 (N_10737,N_9472,N_8463);
nand U10738 (N_10738,N_9571,N_9818);
xor U10739 (N_10739,N_7985,N_7837);
nor U10740 (N_10740,N_8397,N_7533);
nor U10741 (N_10741,N_8106,N_8889);
and U10742 (N_10742,N_8945,N_8970);
xor U10743 (N_10743,N_8494,N_7528);
and U10744 (N_10744,N_7903,N_8132);
or U10745 (N_10745,N_8907,N_8763);
or U10746 (N_10746,N_7671,N_9830);
nor U10747 (N_10747,N_9388,N_8852);
xor U10748 (N_10748,N_9443,N_9904);
nor U10749 (N_10749,N_7803,N_9943);
nand U10750 (N_10750,N_8630,N_8190);
xor U10751 (N_10751,N_8343,N_9298);
nand U10752 (N_10752,N_7553,N_9838);
nor U10753 (N_10753,N_8598,N_8327);
nor U10754 (N_10754,N_7926,N_8337);
and U10755 (N_10755,N_9234,N_9951);
and U10756 (N_10756,N_7684,N_8039);
nor U10757 (N_10757,N_9979,N_9269);
nand U10758 (N_10758,N_8609,N_8761);
and U10759 (N_10759,N_7854,N_9764);
or U10760 (N_10760,N_9495,N_7646);
xor U10761 (N_10761,N_9558,N_9014);
and U10762 (N_10762,N_8413,N_7928);
or U10763 (N_10763,N_8330,N_9556);
and U10764 (N_10764,N_8180,N_9403);
or U10765 (N_10765,N_8849,N_8835);
nand U10766 (N_10766,N_8703,N_9508);
and U10767 (N_10767,N_8821,N_9429);
or U10768 (N_10768,N_9315,N_9447);
or U10769 (N_10769,N_9432,N_9533);
and U10770 (N_10770,N_9789,N_9381);
xnor U10771 (N_10771,N_9489,N_9072);
nand U10772 (N_10772,N_8061,N_9675);
and U10773 (N_10773,N_7650,N_9393);
or U10774 (N_10774,N_8908,N_8145);
or U10775 (N_10775,N_7770,N_9753);
nand U10776 (N_10776,N_7590,N_7880);
or U10777 (N_10777,N_9882,N_7665);
or U10778 (N_10778,N_7771,N_9496);
or U10779 (N_10779,N_8108,N_9112);
and U10780 (N_10780,N_7798,N_7865);
nand U10781 (N_10781,N_8301,N_8535);
or U10782 (N_10782,N_9113,N_8229);
xor U10783 (N_10783,N_8870,N_8468);
and U10784 (N_10784,N_8663,N_9365);
xnor U10785 (N_10785,N_9787,N_9826);
or U10786 (N_10786,N_8729,N_9541);
nand U10787 (N_10787,N_8719,N_8755);
nand U10788 (N_10788,N_8339,N_9754);
xnor U10789 (N_10789,N_9901,N_7822);
nor U10790 (N_10790,N_8851,N_8110);
nor U10791 (N_10791,N_7720,N_8177);
or U10792 (N_10792,N_8577,N_7892);
and U10793 (N_10793,N_8994,N_8396);
nor U10794 (N_10794,N_8982,N_9828);
and U10795 (N_10795,N_9481,N_8318);
or U10796 (N_10796,N_8629,N_8518);
and U10797 (N_10797,N_9233,N_8316);
nand U10798 (N_10798,N_9600,N_7831);
or U10799 (N_10799,N_9804,N_9898);
xor U10800 (N_10800,N_9147,N_7990);
nor U10801 (N_10801,N_9654,N_9218);
nor U10802 (N_10802,N_9740,N_9837);
nor U10803 (N_10803,N_8154,N_8109);
or U10804 (N_10804,N_7585,N_8058);
nand U10805 (N_10805,N_8943,N_8073);
or U10806 (N_10806,N_9190,N_9121);
and U10807 (N_10807,N_9912,N_7755);
and U10808 (N_10808,N_8150,N_8051);
xor U10809 (N_10809,N_8661,N_8590);
xor U10810 (N_10810,N_8778,N_8627);
nand U10811 (N_10811,N_7864,N_9678);
and U10812 (N_10812,N_9289,N_9548);
nor U10813 (N_10813,N_7829,N_8783);
nand U10814 (N_10814,N_9094,N_8645);
and U10815 (N_10815,N_9037,N_7932);
nand U10816 (N_10816,N_8049,N_8185);
nand U10817 (N_10817,N_8187,N_8128);
or U10818 (N_10818,N_9538,N_7690);
or U10819 (N_10819,N_9930,N_8116);
or U10820 (N_10820,N_9570,N_9785);
xnor U10821 (N_10821,N_7604,N_9689);
and U10822 (N_10822,N_9216,N_7936);
xnor U10823 (N_10823,N_8555,N_8738);
and U10824 (N_10824,N_9887,N_9409);
nor U10825 (N_10825,N_9868,N_9153);
or U10826 (N_10826,N_8126,N_7739);
nor U10827 (N_10827,N_9036,N_8696);
xor U10828 (N_10828,N_9044,N_7718);
nand U10829 (N_10829,N_9182,N_9252);
nand U10830 (N_10830,N_8648,N_9971);
or U10831 (N_10831,N_8370,N_8775);
and U10832 (N_10832,N_9611,N_9572);
xor U10833 (N_10833,N_8690,N_8021);
nand U10834 (N_10834,N_8800,N_9340);
nor U10835 (N_10835,N_9649,N_7524);
nor U10836 (N_10836,N_7529,N_9706);
nand U10837 (N_10837,N_8588,N_9065);
or U10838 (N_10838,N_9998,N_9454);
xnor U10839 (N_10839,N_9747,N_8512);
or U10840 (N_10840,N_9415,N_7746);
nand U10841 (N_10841,N_9007,N_7644);
or U10842 (N_10842,N_8071,N_9207);
xor U10843 (N_10843,N_9493,N_9635);
nor U10844 (N_10844,N_9342,N_7776);
nor U10845 (N_10845,N_8308,N_9338);
and U10846 (N_10846,N_9827,N_9105);
or U10847 (N_10847,N_9354,N_9739);
or U10848 (N_10848,N_9994,N_8804);
nand U10849 (N_10849,N_7548,N_8699);
nor U10850 (N_10850,N_8360,N_8561);
nor U10851 (N_10851,N_7801,N_9021);
or U10852 (N_10852,N_9552,N_8507);
and U10853 (N_10853,N_9210,N_7653);
and U10854 (N_10854,N_9633,N_8213);
nand U10855 (N_10855,N_7883,N_9673);
nor U10856 (N_10856,N_9433,N_8204);
or U10857 (N_10857,N_7779,N_8547);
nand U10858 (N_10858,N_8725,N_7629);
or U10859 (N_10859,N_8836,N_8206);
or U10860 (N_10860,N_7867,N_9616);
or U10861 (N_10861,N_8273,N_7748);
nand U10862 (N_10862,N_8915,N_8524);
nand U10863 (N_10863,N_8334,N_9620);
nand U10864 (N_10864,N_7593,N_8814);
and U10865 (N_10865,N_9644,N_7817);
nor U10866 (N_10866,N_8798,N_9968);
xor U10867 (N_10867,N_8819,N_7794);
nor U10868 (N_10868,N_9608,N_8572);
nand U10869 (N_10869,N_8647,N_9136);
nand U10870 (N_10870,N_8454,N_8300);
nor U10871 (N_10871,N_8324,N_8125);
nor U10872 (N_10872,N_8440,N_9009);
and U10873 (N_10873,N_7538,N_8105);
and U10874 (N_10874,N_7606,N_8214);
and U10875 (N_10875,N_9497,N_8750);
and U10876 (N_10876,N_8379,N_9917);
and U10877 (N_10877,N_9300,N_7591);
nor U10878 (N_10878,N_8077,N_7602);
nor U10879 (N_10879,N_9842,N_8079);
xor U10880 (N_10880,N_9569,N_9358);
or U10881 (N_10881,N_8063,N_7871);
nand U10882 (N_10882,N_9175,N_9144);
nand U10883 (N_10883,N_9566,N_9703);
nand U10884 (N_10884,N_8104,N_8548);
nor U10885 (N_10885,N_9435,N_7964);
nor U10886 (N_10886,N_9291,N_9242);
or U10887 (N_10887,N_7758,N_8230);
xor U10888 (N_10888,N_9886,N_8919);
nand U10889 (N_10889,N_8283,N_8483);
or U10890 (N_10890,N_8303,N_8394);
nor U10891 (N_10891,N_9295,N_8769);
or U10892 (N_10892,N_9880,N_7639);
xnor U10893 (N_10893,N_8745,N_8586);
or U10894 (N_10894,N_7708,N_8782);
and U10895 (N_10895,N_9466,N_7941);
nand U10896 (N_10896,N_7678,N_9477);
or U10897 (N_10897,N_8010,N_8388);
xor U10898 (N_10898,N_9440,N_8383);
and U10899 (N_10899,N_7785,N_9825);
nor U10900 (N_10900,N_8752,N_9900);
nor U10901 (N_10901,N_9103,N_7826);
and U10902 (N_10902,N_8200,N_8584);
nor U10903 (N_10903,N_7975,N_9686);
or U10904 (N_10904,N_9442,N_7759);
or U10905 (N_10905,N_9725,N_7825);
or U10906 (N_10906,N_9320,N_8012);
and U10907 (N_10907,N_9305,N_7736);
nor U10908 (N_10908,N_7919,N_8828);
or U10909 (N_10909,N_8084,N_8770);
or U10910 (N_10910,N_7940,N_7566);
nand U10911 (N_10911,N_8959,N_8350);
nand U10912 (N_10912,N_9046,N_8521);
or U10913 (N_10913,N_8712,N_9343);
nor U10914 (N_10914,N_8479,N_9026);
and U10915 (N_10915,N_7968,N_9255);
xor U10916 (N_10916,N_8638,N_9656);
and U10917 (N_10917,N_9622,N_9834);
and U10918 (N_10918,N_9507,N_9069);
or U10919 (N_10919,N_8707,N_9337);
and U10920 (N_10920,N_9630,N_8268);
nor U10921 (N_10921,N_8435,N_7709);
xor U10922 (N_10922,N_9509,N_9506);
and U10923 (N_10923,N_8871,N_9001);
nand U10924 (N_10924,N_7581,N_9553);
nor U10925 (N_10925,N_8975,N_8933);
and U10926 (N_10926,N_9326,N_8352);
and U10927 (N_10927,N_8175,N_8623);
or U10928 (N_10928,N_8619,N_9479);
or U10929 (N_10929,N_8223,N_8002);
nand U10930 (N_10930,N_8977,N_8420);
and U10931 (N_10931,N_7916,N_7943);
or U10932 (N_10932,N_9813,N_8881);
nand U10933 (N_10933,N_8389,N_8322);
xor U10934 (N_10934,N_8989,N_8570);
nor U10935 (N_10935,N_8754,N_8885);
nor U10936 (N_10936,N_7624,N_9659);
and U10937 (N_10937,N_9411,N_8243);
and U10938 (N_10938,N_8843,N_7568);
nor U10939 (N_10939,N_8266,N_9237);
and U10940 (N_10940,N_8739,N_9948);
and U10941 (N_10941,N_9676,N_9355);
nand U10942 (N_10942,N_8866,N_9025);
nor U10943 (N_10943,N_8261,N_9221);
or U10944 (N_10944,N_9772,N_8772);
and U10945 (N_10945,N_8742,N_9400);
or U10946 (N_10946,N_8003,N_8354);
and U10947 (N_10947,N_8103,N_8509);
and U10948 (N_10948,N_8872,N_7971);
and U10949 (N_10949,N_9091,N_8791);
nor U10950 (N_10950,N_7663,N_8141);
or U10951 (N_10951,N_8787,N_9490);
xnor U10952 (N_10952,N_8937,N_7838);
or U10953 (N_10953,N_8290,N_8269);
nor U10954 (N_10954,N_7632,N_9792);
nor U10955 (N_10955,N_9246,N_8262);
or U10956 (N_10956,N_8309,N_8009);
nand U10957 (N_10957,N_9560,N_8148);
nand U10958 (N_10958,N_9924,N_9045);
and U10959 (N_10959,N_9087,N_7615);
nor U10960 (N_10960,N_9743,N_7882);
or U10961 (N_10961,N_9529,N_8784);
and U10962 (N_10962,N_8893,N_7813);
or U10963 (N_10963,N_9692,N_8146);
nor U10964 (N_10964,N_9535,N_8338);
nand U10965 (N_10965,N_8602,N_8632);
or U10966 (N_10966,N_7901,N_9517);
nand U10967 (N_10967,N_8341,N_7631);
nand U10968 (N_10968,N_9926,N_9389);
and U10969 (N_10969,N_7969,N_8720);
xor U10970 (N_10970,N_9959,N_7599);
nand U10971 (N_10971,N_8513,N_8576);
and U10972 (N_10972,N_9319,N_9843);
nand U10973 (N_10973,N_8482,N_8202);
or U10974 (N_10974,N_9192,N_9029);
nor U10975 (N_10975,N_9427,N_8033);
nand U10976 (N_10976,N_8575,N_8372);
and U10977 (N_10977,N_8932,N_9698);
and U10978 (N_10978,N_9975,N_9163);
nor U10979 (N_10979,N_9854,N_8986);
and U10980 (N_10980,N_8456,N_9464);
nor U10981 (N_10981,N_9549,N_8599);
nand U10982 (N_10982,N_8178,N_9292);
nand U10983 (N_10983,N_8329,N_8289);
nor U10984 (N_10984,N_7821,N_9513);
nor U10985 (N_10985,N_9847,N_8196);
and U10986 (N_10986,N_9628,N_9174);
and U10987 (N_10987,N_9821,N_9480);
or U10988 (N_10988,N_9132,N_7805);
nand U10989 (N_10989,N_7830,N_8810);
or U10990 (N_10990,N_8239,N_9162);
or U10991 (N_10991,N_8741,N_9681);
nand U10992 (N_10992,N_7704,N_9724);
and U10993 (N_10993,N_9777,N_9995);
or U10994 (N_10994,N_8651,N_8373);
nand U10995 (N_10995,N_9719,N_7688);
nand U10996 (N_10996,N_8399,N_9711);
and U10997 (N_10997,N_7898,N_9386);
nand U10998 (N_10998,N_9366,N_9806);
and U10999 (N_10999,N_8691,N_8159);
nand U11000 (N_11000,N_9794,N_9126);
nand U11001 (N_11001,N_8906,N_9194);
xnor U11002 (N_11002,N_8540,N_9308);
and U11003 (N_11003,N_7845,N_8244);
and U11004 (N_11004,N_9158,N_9954);
and U11005 (N_11005,N_9406,N_7721);
nor U11006 (N_11006,N_9660,N_8670);
nor U11007 (N_11007,N_9545,N_8006);
or U11008 (N_11008,N_9640,N_9808);
and U11009 (N_11009,N_9524,N_8832);
or U11010 (N_11010,N_9580,N_9108);
nor U11011 (N_11011,N_7927,N_9499);
and U11012 (N_11012,N_8276,N_8384);
xnor U11013 (N_11013,N_8135,N_9518);
or U11014 (N_11014,N_9637,N_7701);
nand U11015 (N_11015,N_8113,N_8876);
nand U11016 (N_11016,N_8620,N_7699);
or U11017 (N_11017,N_8409,N_8685);
or U11018 (N_11018,N_8922,N_9170);
nand U11019 (N_11019,N_9977,N_9551);
or U11020 (N_11020,N_9015,N_8152);
or U11021 (N_11021,N_9445,N_9325);
or U11022 (N_11022,N_8395,N_8375);
nor U11023 (N_11023,N_8822,N_9285);
and U11024 (N_11024,N_9159,N_8248);
or U11025 (N_11025,N_8414,N_8611);
xnor U11026 (N_11026,N_8393,N_9307);
or U11027 (N_11027,N_9664,N_9674);
nand U11028 (N_11028,N_9988,N_7594);
and U11029 (N_11029,N_7963,N_8404);
and U11030 (N_11030,N_7535,N_8768);
nand U11031 (N_11031,N_8254,N_8361);
xnor U11032 (N_11032,N_9684,N_9721);
nand U11033 (N_11033,N_8000,N_9634);
or U11034 (N_11034,N_8764,N_8697);
nor U11035 (N_11035,N_8252,N_9413);
nand U11036 (N_11036,N_8855,N_7734);
nor U11037 (N_11037,N_9310,N_9096);
nor U11038 (N_11038,N_8644,N_9960);
nand U11039 (N_11039,N_8847,N_8247);
nand U11040 (N_11040,N_9169,N_9197);
or U11041 (N_11041,N_9463,N_9658);
nand U11042 (N_11042,N_7622,N_9581);
or U11043 (N_11043,N_7762,N_9455);
nor U11044 (N_11044,N_9140,N_8767);
xnor U11045 (N_11045,N_9181,N_8445);
nor U11046 (N_11046,N_9059,N_8686);
or U11047 (N_11047,N_7732,N_7778);
or U11048 (N_11048,N_9688,N_9384);
and U11049 (N_11049,N_7565,N_9486);
nor U11050 (N_11050,N_9173,N_8407);
nand U11051 (N_11051,N_8068,N_7769);
nor U11052 (N_11052,N_9494,N_8660);
nor U11053 (N_11053,N_8149,N_9856);
nand U11054 (N_11054,N_9731,N_7547);
xnor U11055 (N_11055,N_9641,N_8728);
nand U11056 (N_11056,N_8730,N_7869);
or U11057 (N_11057,N_9330,N_8282);
xnor U11058 (N_11058,N_8169,N_9376);
or U11059 (N_11059,N_7764,N_8117);
nor U11060 (N_11060,N_9516,N_7744);
nor U11061 (N_11061,N_8342,N_9864);
xor U11062 (N_11062,N_8858,N_8676);
nor U11063 (N_11063,N_9768,N_8280);
nor U11064 (N_11064,N_9992,N_9972);
and U11065 (N_11065,N_8425,N_8236);
nor U11066 (N_11066,N_9938,N_9277);
and U11067 (N_11067,N_9585,N_9883);
nand U11068 (N_11068,N_8531,N_7551);
nor U11069 (N_11069,N_8968,N_8711);
or U11070 (N_11070,N_7575,N_8833);
and U11071 (N_11071,N_9262,N_8245);
nand U11072 (N_11072,N_9465,N_8363);
nor U11073 (N_11073,N_9395,N_9407);
xnor U11074 (N_11074,N_8687,N_9035);
xor U11075 (N_11075,N_9261,N_7652);
nand U11076 (N_11076,N_8193,N_8817);
or U11077 (N_11077,N_8781,N_8260);
nor U11078 (N_11078,N_8401,N_9082);
xor U11079 (N_11079,N_9829,N_7858);
and U11080 (N_11080,N_9418,N_8153);
nor U11081 (N_11081,N_8867,N_8471);
nor U11082 (N_11082,N_7626,N_8156);
nand U11083 (N_11083,N_8160,N_8838);
nand U11084 (N_11084,N_9809,N_7525);
nor U11085 (N_11085,N_8055,N_7977);
or U11086 (N_11086,N_9396,N_9742);
nand U11087 (N_11087,N_8299,N_8779);
nand U11088 (N_11088,N_9367,N_8537);
and U11089 (N_11089,N_9260,N_7768);
and U11090 (N_11090,N_9382,N_9284);
nor U11091 (N_11091,N_8824,N_9962);
nand U11092 (N_11092,N_9861,N_8092);
xnor U11093 (N_11093,N_7707,N_9520);
nand U11094 (N_11094,N_7724,N_8914);
and U11095 (N_11095,N_8917,N_9176);
xor U11096 (N_11096,N_7673,N_8724);
nand U11097 (N_11097,N_9228,N_8924);
xnor U11098 (N_11098,N_7989,N_9712);
nand U11099 (N_11099,N_9697,N_7597);
or U11100 (N_11100,N_7894,N_8366);
nand U11101 (N_11101,N_8014,N_9482);
nand U11102 (N_11102,N_8585,N_9148);
and U11103 (N_11103,N_8037,N_9744);
or U11104 (N_11104,N_8966,N_7630);
and U11105 (N_11105,N_7761,N_8270);
or U11106 (N_11106,N_8082,N_8041);
xor U11107 (N_11107,N_8873,N_9370);
and U11108 (N_11108,N_7917,N_8746);
nand U11109 (N_11109,N_8311,N_8023);
or U11110 (N_11110,N_8459,N_8928);
nand U11111 (N_11111,N_9667,N_8952);
nand U11112 (N_11112,N_9076,N_7640);
and U11113 (N_11113,N_8771,N_8920);
or U11114 (N_11114,N_9050,N_7921);
or U11115 (N_11115,N_7962,N_9222);
nor U11116 (N_11116,N_9893,N_8478);
and U11117 (N_11117,N_7953,N_7784);
nor U11118 (N_11118,N_8790,N_7973);
nor U11119 (N_11119,N_9694,N_8622);
nor U11120 (N_11120,N_9799,N_7574);
nor U11121 (N_11121,N_8123,N_8131);
or U11122 (N_11122,N_9980,N_9470);
nor U11123 (N_11123,N_9539,N_9145);
and U11124 (N_11124,N_8514,N_9028);
nand U11125 (N_11125,N_7609,N_8997);
and U11126 (N_11126,N_8839,N_9941);
nand U11127 (N_11127,N_8371,N_9339);
nor U11128 (N_11128,N_9550,N_9699);
nor U11129 (N_11129,N_8416,N_7828);
nor U11130 (N_11130,N_7657,N_9836);
or U11131 (N_11131,N_8942,N_8488);
nand U11132 (N_11132,N_7875,N_8733);
nor U11133 (N_11133,N_8295,N_9922);
and U11134 (N_11134,N_9543,N_7735);
and U11135 (N_11135,N_7577,N_8904);
and U11136 (N_11136,N_9500,N_7527);
nor U11137 (N_11137,N_9341,N_8428);
nand U11138 (N_11138,N_9311,N_9907);
or U11139 (N_11139,N_9168,N_9879);
nor U11140 (N_11140,N_8961,N_9591);
nand U11141 (N_11141,N_9958,N_9668);
nor U11142 (N_11142,N_8221,N_9578);
nor U11143 (N_11143,N_8481,N_8218);
and U11144 (N_11144,N_7702,N_8785);
and U11145 (N_11145,N_9762,N_9279);
nand U11146 (N_11146,N_8834,N_7861);
xor U11147 (N_11147,N_7611,N_9625);
nor U11148 (N_11148,N_9245,N_9718);
nor U11149 (N_11149,N_7738,N_9631);
xor U11150 (N_11150,N_9165,N_7698);
or U11151 (N_11151,N_8582,N_9903);
nor U11152 (N_11152,N_8201,N_8323);
or U11153 (N_11153,N_9492,N_9213);
or U11154 (N_11154,N_9070,N_8078);
or U11155 (N_11155,N_9947,N_8776);
or U11156 (N_11156,N_8281,N_9683);
or U11157 (N_11157,N_9446,N_8978);
or U11158 (N_11158,N_8042,N_7686);
or U11159 (N_11159,N_8025,N_7879);
nand U11160 (N_11160,N_9991,N_9786);
or U11161 (N_11161,N_8001,N_7536);
or U11162 (N_11162,N_9594,N_7540);
nand U11163 (N_11163,N_9704,N_8100);
nor U11164 (N_11164,N_9603,N_8059);
and U11165 (N_11165,N_8846,N_9141);
or U11166 (N_11166,N_8381,N_8240);
and U11167 (N_11167,N_9123,N_8208);
nand U11168 (N_11168,N_8155,N_9275);
and U11169 (N_11169,N_8492,N_7542);
or U11170 (N_11170,N_7839,N_8469);
and U11171 (N_11171,N_9016,N_9885);
or U11172 (N_11172,N_8181,N_7855);
nand U11173 (N_11173,N_9596,N_8314);
xnor U11174 (N_11174,N_9970,N_8130);
and U11175 (N_11175,N_8996,N_8718);
or U11176 (N_11176,N_8675,N_7534);
and U11177 (N_11177,N_7908,N_8587);
nand U11178 (N_11178,N_8167,N_8278);
and U11179 (N_11179,N_8865,N_8613);
nor U11180 (N_11180,N_7600,N_9961);
or U11181 (N_11181,N_8496,N_9451);
nand U11182 (N_11182,N_9590,N_7687);
or U11183 (N_11183,N_9161,N_9215);
nor U11184 (N_11184,N_8842,N_7790);
and U11185 (N_11185,N_7918,N_8850);
nand U11186 (N_11186,N_8681,N_8734);
or U11187 (N_11187,N_8571,N_9483);
xor U11188 (N_11188,N_7777,N_9546);
nor U11189 (N_11189,N_9531,N_9989);
and U11190 (N_11190,N_8811,N_9542);
nor U11191 (N_11191,N_8348,N_9304);
or U11192 (N_11192,N_8737,N_9357);
nand U11193 (N_11193,N_9306,N_9189);
xnor U11194 (N_11194,N_9547,N_9438);
or U11195 (N_11195,N_8654,N_7666);
and U11196 (N_11196,N_9851,N_9345);
xnor U11197 (N_11197,N_9377,N_8364);
nand U11198 (N_11198,N_9927,N_9452);
and U11199 (N_11199,N_8060,N_9824);
or U11200 (N_11200,N_7740,N_8358);
nand U11201 (N_11201,N_9219,N_8256);
nand U11202 (N_11202,N_8795,N_8581);
nor U11203 (N_11203,N_9525,N_8222);
and U11204 (N_11204,N_9610,N_7891);
xnor U11205 (N_11205,N_8263,N_8508);
or U11206 (N_11206,N_9083,N_8265);
and U11207 (N_11207,N_8355,N_8241);
nor U11208 (N_11208,N_7970,N_9309);
xnor U11209 (N_11209,N_7510,N_8203);
nand U11210 (N_11210,N_7557,N_9336);
and U11211 (N_11211,N_7793,N_8172);
and U11212 (N_11212,N_9741,N_8792);
or U11213 (N_11213,N_8296,N_9073);
or U11214 (N_11214,N_9362,N_8944);
nor U11215 (N_11215,N_9710,N_8801);
nand U11216 (N_11216,N_9240,N_9312);
and U11217 (N_11217,N_9672,N_8013);
xnor U11218 (N_11218,N_7504,N_9758);
nor U11219 (N_11219,N_8173,N_8487);
nand U11220 (N_11220,N_9238,N_9862);
xnor U11221 (N_11221,N_8191,N_9621);
xor U11222 (N_11222,N_8486,N_8285);
nand U11223 (N_11223,N_9840,N_8121);
nor U11224 (N_11224,N_9878,N_9597);
and U11225 (N_11225,N_9895,N_9577);
nand U11226 (N_11226,N_8233,N_8412);
and U11227 (N_11227,N_7705,N_8094);
xnor U11228 (N_11228,N_9266,N_8516);
or U11229 (N_11229,N_8386,N_8011);
or U11230 (N_11230,N_8732,N_8500);
xnor U11231 (N_11231,N_9209,N_9054);
or U11232 (N_11232,N_8744,N_9761);
nor U11233 (N_11233,N_8934,N_7767);
or U11234 (N_11234,N_9528,N_9081);
and U11235 (N_11235,N_7922,N_9766);
or U11236 (N_11236,N_8293,N_9583);
nand U11237 (N_11237,N_9412,N_8249);
or U11238 (N_11238,N_7938,N_9502);
or U11239 (N_11239,N_8028,N_9714);
and U11240 (N_11240,N_7537,N_9982);
and U11241 (N_11241,N_7679,N_9891);
or U11242 (N_11242,N_9565,N_8999);
and U11243 (N_11243,N_9071,N_7849);
and U11244 (N_11244,N_8677,N_9154);
nor U11245 (N_11245,N_7512,N_7722);
nand U11246 (N_11246,N_8199,N_9356);
nor U11247 (N_11247,N_7618,N_9030);
nor U11248 (N_11248,N_8559,N_8990);
and U11249 (N_11249,N_9322,N_8253);
or U11250 (N_11250,N_7783,N_9377);
nor U11251 (N_11251,N_7795,N_9585);
nand U11252 (N_11252,N_8274,N_9081);
nand U11253 (N_11253,N_7581,N_9176);
or U11254 (N_11254,N_7911,N_9775);
and U11255 (N_11255,N_8677,N_8079);
nor U11256 (N_11256,N_8873,N_8956);
or U11257 (N_11257,N_7827,N_9516);
and U11258 (N_11258,N_8991,N_8680);
and U11259 (N_11259,N_9629,N_9440);
or U11260 (N_11260,N_8819,N_7753);
xnor U11261 (N_11261,N_8415,N_8014);
nor U11262 (N_11262,N_7751,N_9410);
nand U11263 (N_11263,N_9661,N_8594);
or U11264 (N_11264,N_7950,N_9345);
or U11265 (N_11265,N_8705,N_9709);
nor U11266 (N_11266,N_8672,N_7715);
nor U11267 (N_11267,N_8979,N_9603);
nand U11268 (N_11268,N_8252,N_8959);
xor U11269 (N_11269,N_9267,N_9572);
nand U11270 (N_11270,N_9785,N_8917);
or U11271 (N_11271,N_8703,N_8201);
xor U11272 (N_11272,N_9850,N_9366);
nor U11273 (N_11273,N_8287,N_9639);
nor U11274 (N_11274,N_9526,N_9882);
or U11275 (N_11275,N_8188,N_9568);
nor U11276 (N_11276,N_8419,N_8778);
or U11277 (N_11277,N_7630,N_8168);
nor U11278 (N_11278,N_9202,N_7713);
and U11279 (N_11279,N_9313,N_8610);
nand U11280 (N_11280,N_9926,N_9662);
and U11281 (N_11281,N_9466,N_7616);
nor U11282 (N_11282,N_8836,N_7952);
or U11283 (N_11283,N_9214,N_9838);
and U11284 (N_11284,N_8191,N_7841);
nand U11285 (N_11285,N_7642,N_8341);
and U11286 (N_11286,N_9926,N_8479);
or U11287 (N_11287,N_8023,N_9186);
nor U11288 (N_11288,N_8361,N_7981);
nor U11289 (N_11289,N_8863,N_9440);
nor U11290 (N_11290,N_8255,N_9971);
nand U11291 (N_11291,N_8882,N_8316);
or U11292 (N_11292,N_7777,N_9430);
nand U11293 (N_11293,N_8247,N_9441);
nor U11294 (N_11294,N_7772,N_9376);
or U11295 (N_11295,N_8456,N_8556);
and U11296 (N_11296,N_9522,N_9818);
and U11297 (N_11297,N_7721,N_9693);
and U11298 (N_11298,N_9787,N_8998);
and U11299 (N_11299,N_8531,N_9418);
and U11300 (N_11300,N_9082,N_7731);
nand U11301 (N_11301,N_9011,N_9029);
xnor U11302 (N_11302,N_8968,N_9605);
nand U11303 (N_11303,N_8348,N_9186);
and U11304 (N_11304,N_8930,N_8778);
or U11305 (N_11305,N_8071,N_9082);
and U11306 (N_11306,N_8655,N_8063);
nand U11307 (N_11307,N_7555,N_9844);
nand U11308 (N_11308,N_9486,N_8286);
nor U11309 (N_11309,N_9392,N_9631);
xor U11310 (N_11310,N_9560,N_8862);
nand U11311 (N_11311,N_8762,N_9210);
xor U11312 (N_11312,N_7968,N_7738);
xnor U11313 (N_11313,N_9574,N_9559);
nand U11314 (N_11314,N_9827,N_8145);
or U11315 (N_11315,N_8350,N_9958);
xnor U11316 (N_11316,N_7685,N_9514);
nand U11317 (N_11317,N_7691,N_8114);
nor U11318 (N_11318,N_7683,N_8930);
and U11319 (N_11319,N_9220,N_8673);
and U11320 (N_11320,N_8319,N_7679);
nor U11321 (N_11321,N_8392,N_8185);
nand U11322 (N_11322,N_7951,N_7777);
nand U11323 (N_11323,N_7911,N_8315);
xnor U11324 (N_11324,N_9471,N_7727);
xnor U11325 (N_11325,N_9249,N_9209);
nor U11326 (N_11326,N_8864,N_7873);
xor U11327 (N_11327,N_8485,N_7632);
or U11328 (N_11328,N_9337,N_8598);
and U11329 (N_11329,N_9150,N_9233);
xnor U11330 (N_11330,N_9090,N_7756);
nand U11331 (N_11331,N_8414,N_8531);
or U11332 (N_11332,N_9102,N_8418);
nand U11333 (N_11333,N_7608,N_8808);
nand U11334 (N_11334,N_7590,N_9975);
nand U11335 (N_11335,N_8320,N_9555);
or U11336 (N_11336,N_8625,N_8899);
and U11337 (N_11337,N_8016,N_8768);
nor U11338 (N_11338,N_9796,N_8288);
nor U11339 (N_11339,N_8454,N_7651);
xnor U11340 (N_11340,N_9131,N_7904);
nor U11341 (N_11341,N_7968,N_9411);
nand U11342 (N_11342,N_9293,N_7914);
nand U11343 (N_11343,N_7570,N_8017);
nand U11344 (N_11344,N_9280,N_8009);
nor U11345 (N_11345,N_8886,N_9094);
or U11346 (N_11346,N_9003,N_7665);
nand U11347 (N_11347,N_7705,N_9898);
nand U11348 (N_11348,N_7841,N_8841);
nand U11349 (N_11349,N_7804,N_8728);
xnor U11350 (N_11350,N_9491,N_8393);
xor U11351 (N_11351,N_8249,N_9268);
or U11352 (N_11352,N_8058,N_7745);
and U11353 (N_11353,N_8665,N_8354);
nor U11354 (N_11354,N_7810,N_9708);
nor U11355 (N_11355,N_9556,N_9442);
or U11356 (N_11356,N_8110,N_8483);
nand U11357 (N_11357,N_9677,N_9628);
or U11358 (N_11358,N_9424,N_9996);
and U11359 (N_11359,N_8540,N_8048);
nor U11360 (N_11360,N_8347,N_9262);
nor U11361 (N_11361,N_8481,N_9188);
or U11362 (N_11362,N_9644,N_9248);
and U11363 (N_11363,N_9741,N_9498);
nand U11364 (N_11364,N_7804,N_8480);
nor U11365 (N_11365,N_9799,N_8876);
nand U11366 (N_11366,N_7834,N_9296);
nor U11367 (N_11367,N_7993,N_7810);
nor U11368 (N_11368,N_8675,N_9231);
or U11369 (N_11369,N_9063,N_7727);
nor U11370 (N_11370,N_7619,N_7628);
and U11371 (N_11371,N_9316,N_9703);
nor U11372 (N_11372,N_7975,N_8354);
or U11373 (N_11373,N_8514,N_8063);
nor U11374 (N_11374,N_8413,N_8561);
and U11375 (N_11375,N_7905,N_7961);
nor U11376 (N_11376,N_9360,N_9975);
or U11377 (N_11377,N_9100,N_7721);
or U11378 (N_11378,N_7877,N_8025);
nand U11379 (N_11379,N_7664,N_9024);
nor U11380 (N_11380,N_9085,N_9597);
nand U11381 (N_11381,N_9334,N_7536);
nand U11382 (N_11382,N_9455,N_9987);
nor U11383 (N_11383,N_7807,N_9044);
nand U11384 (N_11384,N_9253,N_9798);
nand U11385 (N_11385,N_9523,N_9696);
nor U11386 (N_11386,N_8898,N_8704);
or U11387 (N_11387,N_8233,N_7622);
or U11388 (N_11388,N_9980,N_9963);
nor U11389 (N_11389,N_9221,N_7671);
and U11390 (N_11390,N_9705,N_7939);
and U11391 (N_11391,N_9244,N_7859);
nor U11392 (N_11392,N_8235,N_8081);
and U11393 (N_11393,N_8937,N_9860);
and U11394 (N_11394,N_9366,N_8051);
or U11395 (N_11395,N_8937,N_8633);
nand U11396 (N_11396,N_9885,N_9616);
and U11397 (N_11397,N_7557,N_9168);
nor U11398 (N_11398,N_9442,N_8636);
nand U11399 (N_11399,N_9845,N_9983);
nor U11400 (N_11400,N_9584,N_7612);
or U11401 (N_11401,N_7730,N_7586);
nand U11402 (N_11402,N_8107,N_9064);
or U11403 (N_11403,N_9160,N_9181);
nor U11404 (N_11404,N_8202,N_9764);
nand U11405 (N_11405,N_8269,N_9159);
and U11406 (N_11406,N_9682,N_7778);
nand U11407 (N_11407,N_9450,N_8839);
xnor U11408 (N_11408,N_9022,N_8514);
nand U11409 (N_11409,N_7510,N_9381);
or U11410 (N_11410,N_7676,N_8029);
or U11411 (N_11411,N_8319,N_8923);
nand U11412 (N_11412,N_9739,N_8150);
and U11413 (N_11413,N_9170,N_8960);
nor U11414 (N_11414,N_9314,N_7796);
or U11415 (N_11415,N_7510,N_9980);
nand U11416 (N_11416,N_9236,N_9893);
nand U11417 (N_11417,N_7891,N_7830);
nor U11418 (N_11418,N_7891,N_8912);
nor U11419 (N_11419,N_7571,N_9690);
xnor U11420 (N_11420,N_8354,N_9447);
and U11421 (N_11421,N_9723,N_9006);
and U11422 (N_11422,N_9295,N_7624);
nand U11423 (N_11423,N_9255,N_9715);
and U11424 (N_11424,N_9288,N_9353);
and U11425 (N_11425,N_9406,N_9533);
nand U11426 (N_11426,N_8863,N_9464);
and U11427 (N_11427,N_8075,N_9908);
or U11428 (N_11428,N_9022,N_9996);
xor U11429 (N_11429,N_9888,N_8100);
xor U11430 (N_11430,N_9854,N_8760);
nand U11431 (N_11431,N_7581,N_9432);
or U11432 (N_11432,N_7819,N_9623);
nand U11433 (N_11433,N_7946,N_9371);
and U11434 (N_11434,N_9129,N_9267);
nor U11435 (N_11435,N_9607,N_8497);
and U11436 (N_11436,N_8497,N_9442);
nor U11437 (N_11437,N_7545,N_9174);
or U11438 (N_11438,N_9652,N_9098);
xor U11439 (N_11439,N_9072,N_9200);
and U11440 (N_11440,N_7770,N_7749);
and U11441 (N_11441,N_7967,N_9159);
nor U11442 (N_11442,N_8742,N_8681);
nand U11443 (N_11443,N_9718,N_8078);
or U11444 (N_11444,N_9140,N_8893);
and U11445 (N_11445,N_8612,N_8753);
or U11446 (N_11446,N_9044,N_9594);
or U11447 (N_11447,N_7731,N_8456);
and U11448 (N_11448,N_9480,N_8032);
or U11449 (N_11449,N_8673,N_9404);
nand U11450 (N_11450,N_8210,N_9932);
nand U11451 (N_11451,N_8190,N_8227);
nor U11452 (N_11452,N_8007,N_9857);
xnor U11453 (N_11453,N_9558,N_9511);
xnor U11454 (N_11454,N_7762,N_8117);
xor U11455 (N_11455,N_8254,N_8882);
and U11456 (N_11456,N_8607,N_8198);
and U11457 (N_11457,N_8844,N_9142);
nor U11458 (N_11458,N_9088,N_9929);
or U11459 (N_11459,N_8282,N_8929);
nor U11460 (N_11460,N_8266,N_7561);
nor U11461 (N_11461,N_7963,N_9873);
nand U11462 (N_11462,N_9826,N_9597);
nor U11463 (N_11463,N_8266,N_7781);
and U11464 (N_11464,N_8830,N_9519);
nor U11465 (N_11465,N_7623,N_9839);
nand U11466 (N_11466,N_8370,N_9872);
nand U11467 (N_11467,N_9102,N_8189);
nor U11468 (N_11468,N_9840,N_9353);
and U11469 (N_11469,N_8071,N_8152);
nand U11470 (N_11470,N_7540,N_9944);
nand U11471 (N_11471,N_8027,N_8999);
nor U11472 (N_11472,N_8336,N_9593);
nor U11473 (N_11473,N_7986,N_8711);
nand U11474 (N_11474,N_9272,N_9127);
and U11475 (N_11475,N_8462,N_9695);
nor U11476 (N_11476,N_9019,N_9294);
and U11477 (N_11477,N_9163,N_9126);
or U11478 (N_11478,N_8788,N_7519);
nand U11479 (N_11479,N_9589,N_9158);
nand U11480 (N_11480,N_8342,N_9560);
nand U11481 (N_11481,N_9771,N_7523);
and U11482 (N_11482,N_8046,N_9762);
nand U11483 (N_11483,N_9586,N_7657);
nor U11484 (N_11484,N_8493,N_9540);
nor U11485 (N_11485,N_9348,N_8282);
nor U11486 (N_11486,N_8288,N_8733);
and U11487 (N_11487,N_7988,N_8053);
or U11488 (N_11488,N_9982,N_7749);
xor U11489 (N_11489,N_8513,N_8612);
and U11490 (N_11490,N_8982,N_9130);
nand U11491 (N_11491,N_9091,N_9063);
or U11492 (N_11492,N_7512,N_8106);
nor U11493 (N_11493,N_7703,N_8273);
or U11494 (N_11494,N_7518,N_7691);
or U11495 (N_11495,N_7794,N_9002);
or U11496 (N_11496,N_9273,N_9036);
nor U11497 (N_11497,N_9435,N_8757);
or U11498 (N_11498,N_9820,N_8730);
nor U11499 (N_11499,N_8269,N_8691);
nor U11500 (N_11500,N_9220,N_9006);
nor U11501 (N_11501,N_9411,N_7827);
nand U11502 (N_11502,N_9948,N_7923);
xor U11503 (N_11503,N_7558,N_9481);
nor U11504 (N_11504,N_7801,N_8623);
xor U11505 (N_11505,N_9778,N_8206);
nand U11506 (N_11506,N_8737,N_8705);
or U11507 (N_11507,N_8789,N_7576);
nand U11508 (N_11508,N_8760,N_9727);
nand U11509 (N_11509,N_8422,N_9565);
xnor U11510 (N_11510,N_9193,N_9905);
nand U11511 (N_11511,N_8901,N_9752);
xor U11512 (N_11512,N_8406,N_7697);
and U11513 (N_11513,N_8007,N_8603);
nand U11514 (N_11514,N_7745,N_9811);
and U11515 (N_11515,N_9244,N_9057);
and U11516 (N_11516,N_8809,N_9590);
and U11517 (N_11517,N_9143,N_8370);
nor U11518 (N_11518,N_8105,N_9623);
nor U11519 (N_11519,N_7826,N_9457);
and U11520 (N_11520,N_8467,N_9951);
and U11521 (N_11521,N_9402,N_8063);
nand U11522 (N_11522,N_7972,N_8276);
nand U11523 (N_11523,N_9257,N_9017);
nand U11524 (N_11524,N_8537,N_9261);
and U11525 (N_11525,N_9051,N_8795);
nor U11526 (N_11526,N_8988,N_7653);
nor U11527 (N_11527,N_8389,N_9565);
or U11528 (N_11528,N_7929,N_7607);
or U11529 (N_11529,N_8976,N_9718);
xor U11530 (N_11530,N_9371,N_9998);
nand U11531 (N_11531,N_8242,N_9295);
nand U11532 (N_11532,N_9946,N_9259);
nand U11533 (N_11533,N_8453,N_9344);
or U11534 (N_11534,N_8225,N_9327);
and U11535 (N_11535,N_8363,N_8153);
nor U11536 (N_11536,N_8691,N_9166);
nor U11537 (N_11537,N_7843,N_9229);
and U11538 (N_11538,N_9179,N_9620);
nand U11539 (N_11539,N_9394,N_8888);
nor U11540 (N_11540,N_8237,N_7612);
xor U11541 (N_11541,N_9053,N_9702);
nand U11542 (N_11542,N_7546,N_8446);
nand U11543 (N_11543,N_7641,N_9609);
nor U11544 (N_11544,N_9804,N_7915);
or U11545 (N_11545,N_9914,N_8797);
nor U11546 (N_11546,N_7636,N_9027);
nand U11547 (N_11547,N_8091,N_8508);
and U11548 (N_11548,N_8611,N_9429);
nand U11549 (N_11549,N_8173,N_9800);
nor U11550 (N_11550,N_9795,N_9439);
or U11551 (N_11551,N_9795,N_9420);
nand U11552 (N_11552,N_8082,N_7546);
and U11553 (N_11553,N_9132,N_8200);
nor U11554 (N_11554,N_9610,N_9363);
xor U11555 (N_11555,N_9624,N_9303);
nand U11556 (N_11556,N_8396,N_8811);
nand U11557 (N_11557,N_8155,N_8657);
nand U11558 (N_11558,N_8878,N_7637);
xor U11559 (N_11559,N_9867,N_8804);
nor U11560 (N_11560,N_7857,N_8333);
and U11561 (N_11561,N_9318,N_9019);
xor U11562 (N_11562,N_7627,N_7821);
and U11563 (N_11563,N_8950,N_8501);
and U11564 (N_11564,N_9914,N_8497);
nand U11565 (N_11565,N_7622,N_9496);
nor U11566 (N_11566,N_8747,N_8701);
or U11567 (N_11567,N_9197,N_9604);
and U11568 (N_11568,N_9063,N_8981);
nor U11569 (N_11569,N_8582,N_9719);
and U11570 (N_11570,N_9696,N_8308);
nand U11571 (N_11571,N_8214,N_9812);
or U11572 (N_11572,N_9615,N_7940);
nor U11573 (N_11573,N_7773,N_9227);
nor U11574 (N_11574,N_7558,N_8350);
nand U11575 (N_11575,N_8462,N_8248);
nor U11576 (N_11576,N_8625,N_9237);
nor U11577 (N_11577,N_9680,N_8581);
nand U11578 (N_11578,N_9569,N_8440);
or U11579 (N_11579,N_9855,N_7673);
or U11580 (N_11580,N_8599,N_9813);
nand U11581 (N_11581,N_7982,N_7641);
or U11582 (N_11582,N_8121,N_8540);
nand U11583 (N_11583,N_8605,N_7952);
nand U11584 (N_11584,N_9505,N_8339);
xnor U11585 (N_11585,N_8069,N_9783);
nand U11586 (N_11586,N_8197,N_8052);
and U11587 (N_11587,N_7713,N_8699);
nand U11588 (N_11588,N_9731,N_8754);
nand U11589 (N_11589,N_9638,N_7514);
nor U11590 (N_11590,N_9794,N_8773);
nor U11591 (N_11591,N_9474,N_8457);
and U11592 (N_11592,N_9001,N_8835);
or U11593 (N_11593,N_9638,N_7752);
xnor U11594 (N_11594,N_9373,N_9238);
or U11595 (N_11595,N_8287,N_8209);
or U11596 (N_11596,N_9089,N_9649);
or U11597 (N_11597,N_9354,N_8304);
xnor U11598 (N_11598,N_9121,N_9151);
nand U11599 (N_11599,N_7761,N_9279);
and U11600 (N_11600,N_8616,N_8851);
or U11601 (N_11601,N_9118,N_9950);
nand U11602 (N_11602,N_9148,N_8316);
nand U11603 (N_11603,N_9119,N_8042);
nand U11604 (N_11604,N_8468,N_7922);
and U11605 (N_11605,N_7688,N_8306);
nor U11606 (N_11606,N_7756,N_7821);
nor U11607 (N_11607,N_7785,N_9540);
and U11608 (N_11608,N_9703,N_7683);
nor U11609 (N_11609,N_8116,N_8897);
nand U11610 (N_11610,N_7701,N_9883);
and U11611 (N_11611,N_9308,N_9530);
and U11612 (N_11612,N_8546,N_7935);
xnor U11613 (N_11613,N_8141,N_8880);
and U11614 (N_11614,N_8184,N_9059);
or U11615 (N_11615,N_9816,N_7601);
nor U11616 (N_11616,N_8488,N_8897);
or U11617 (N_11617,N_8660,N_9313);
and U11618 (N_11618,N_8508,N_7966);
and U11619 (N_11619,N_9211,N_9901);
nand U11620 (N_11620,N_9705,N_8835);
or U11621 (N_11621,N_8181,N_9056);
xor U11622 (N_11622,N_8822,N_8995);
nand U11623 (N_11623,N_9629,N_8923);
nand U11624 (N_11624,N_9529,N_8234);
xnor U11625 (N_11625,N_9178,N_9328);
and U11626 (N_11626,N_9413,N_8484);
and U11627 (N_11627,N_8430,N_9439);
nor U11628 (N_11628,N_8691,N_8292);
nand U11629 (N_11629,N_9963,N_9155);
and U11630 (N_11630,N_9895,N_9027);
nor U11631 (N_11631,N_8679,N_7552);
xnor U11632 (N_11632,N_8712,N_8437);
nor U11633 (N_11633,N_8721,N_8005);
nor U11634 (N_11634,N_9210,N_7910);
nand U11635 (N_11635,N_8392,N_7703);
nand U11636 (N_11636,N_8766,N_8452);
or U11637 (N_11637,N_9749,N_8677);
nand U11638 (N_11638,N_9026,N_8798);
or U11639 (N_11639,N_7815,N_7935);
or U11640 (N_11640,N_9378,N_9772);
nand U11641 (N_11641,N_7851,N_8891);
or U11642 (N_11642,N_9585,N_9591);
and U11643 (N_11643,N_9698,N_9068);
and U11644 (N_11644,N_9143,N_9317);
or U11645 (N_11645,N_8922,N_7594);
and U11646 (N_11646,N_7987,N_9424);
and U11647 (N_11647,N_7836,N_7614);
and U11648 (N_11648,N_8268,N_7865);
nand U11649 (N_11649,N_8369,N_8360);
or U11650 (N_11650,N_9064,N_8640);
nand U11651 (N_11651,N_9954,N_8021);
and U11652 (N_11652,N_8067,N_9574);
nor U11653 (N_11653,N_9656,N_8089);
nor U11654 (N_11654,N_7725,N_8560);
nand U11655 (N_11655,N_8814,N_8564);
or U11656 (N_11656,N_9744,N_9823);
and U11657 (N_11657,N_8508,N_7979);
nor U11658 (N_11658,N_7531,N_8430);
nand U11659 (N_11659,N_8704,N_9623);
xor U11660 (N_11660,N_9726,N_8470);
nor U11661 (N_11661,N_9781,N_8018);
and U11662 (N_11662,N_7740,N_7521);
and U11663 (N_11663,N_9105,N_9468);
or U11664 (N_11664,N_9435,N_9124);
and U11665 (N_11665,N_9790,N_8343);
or U11666 (N_11666,N_9589,N_8138);
and U11667 (N_11667,N_8076,N_8019);
and U11668 (N_11668,N_8701,N_8912);
and U11669 (N_11669,N_8897,N_9827);
and U11670 (N_11670,N_8274,N_9489);
nand U11671 (N_11671,N_7554,N_7908);
or U11672 (N_11672,N_9437,N_7666);
and U11673 (N_11673,N_9074,N_9478);
xor U11674 (N_11674,N_8883,N_8819);
nor U11675 (N_11675,N_7544,N_7702);
xnor U11676 (N_11676,N_9228,N_8449);
nand U11677 (N_11677,N_9385,N_8378);
xor U11678 (N_11678,N_8718,N_7802);
and U11679 (N_11679,N_7515,N_8144);
nand U11680 (N_11680,N_8004,N_7777);
nand U11681 (N_11681,N_9371,N_8271);
nand U11682 (N_11682,N_9668,N_7646);
nand U11683 (N_11683,N_7979,N_8469);
nor U11684 (N_11684,N_7545,N_8011);
nand U11685 (N_11685,N_9475,N_8889);
or U11686 (N_11686,N_8114,N_9988);
nor U11687 (N_11687,N_7619,N_9888);
nand U11688 (N_11688,N_9043,N_8416);
nor U11689 (N_11689,N_8687,N_8589);
nand U11690 (N_11690,N_9907,N_8872);
or U11691 (N_11691,N_8240,N_8209);
nand U11692 (N_11692,N_8485,N_8608);
or U11693 (N_11693,N_9081,N_7547);
nor U11694 (N_11694,N_8483,N_8722);
and U11695 (N_11695,N_8118,N_8985);
nand U11696 (N_11696,N_8096,N_7582);
nor U11697 (N_11697,N_9131,N_9313);
or U11698 (N_11698,N_8661,N_7872);
nor U11699 (N_11699,N_8412,N_7808);
or U11700 (N_11700,N_9172,N_9103);
nor U11701 (N_11701,N_8053,N_9295);
and U11702 (N_11702,N_8222,N_7795);
and U11703 (N_11703,N_8873,N_8635);
and U11704 (N_11704,N_9627,N_9773);
and U11705 (N_11705,N_8195,N_9811);
nand U11706 (N_11706,N_8988,N_7543);
nor U11707 (N_11707,N_8989,N_7801);
nand U11708 (N_11708,N_8431,N_7851);
nand U11709 (N_11709,N_8083,N_8869);
or U11710 (N_11710,N_9080,N_8496);
and U11711 (N_11711,N_7871,N_9892);
or U11712 (N_11712,N_7596,N_8757);
nor U11713 (N_11713,N_7935,N_9410);
nand U11714 (N_11714,N_9141,N_9176);
and U11715 (N_11715,N_9967,N_8909);
and U11716 (N_11716,N_9354,N_8897);
and U11717 (N_11717,N_8634,N_8334);
nor U11718 (N_11718,N_8831,N_8877);
or U11719 (N_11719,N_8265,N_9997);
nor U11720 (N_11720,N_9550,N_8292);
nor U11721 (N_11721,N_9815,N_7972);
and U11722 (N_11722,N_8575,N_8568);
nand U11723 (N_11723,N_8818,N_8298);
and U11724 (N_11724,N_9266,N_7860);
nor U11725 (N_11725,N_9242,N_9938);
nand U11726 (N_11726,N_8120,N_9149);
or U11727 (N_11727,N_8355,N_9042);
xor U11728 (N_11728,N_7587,N_8452);
xor U11729 (N_11729,N_9930,N_7715);
or U11730 (N_11730,N_8487,N_8236);
nor U11731 (N_11731,N_9916,N_9359);
nand U11732 (N_11732,N_8779,N_9628);
and U11733 (N_11733,N_8821,N_9546);
and U11734 (N_11734,N_8177,N_8816);
and U11735 (N_11735,N_8570,N_7808);
nand U11736 (N_11736,N_7763,N_9036);
nor U11737 (N_11737,N_9751,N_8463);
nand U11738 (N_11738,N_8840,N_8369);
and U11739 (N_11739,N_8617,N_9259);
xor U11740 (N_11740,N_8752,N_8969);
nand U11741 (N_11741,N_9266,N_8567);
or U11742 (N_11742,N_9995,N_9555);
nand U11743 (N_11743,N_9022,N_9319);
or U11744 (N_11744,N_9307,N_8114);
and U11745 (N_11745,N_9803,N_7835);
nand U11746 (N_11746,N_7538,N_9442);
nor U11747 (N_11747,N_8452,N_8863);
nor U11748 (N_11748,N_9992,N_8719);
or U11749 (N_11749,N_9800,N_8436);
and U11750 (N_11750,N_9404,N_8933);
or U11751 (N_11751,N_7838,N_9527);
and U11752 (N_11752,N_9032,N_8386);
nor U11753 (N_11753,N_8274,N_9223);
nor U11754 (N_11754,N_8689,N_8276);
or U11755 (N_11755,N_7686,N_8773);
or U11756 (N_11756,N_9112,N_9479);
nand U11757 (N_11757,N_9290,N_8802);
xor U11758 (N_11758,N_9496,N_9922);
and U11759 (N_11759,N_8552,N_9133);
and U11760 (N_11760,N_8420,N_7963);
and U11761 (N_11761,N_7991,N_8942);
or U11762 (N_11762,N_7626,N_8013);
nand U11763 (N_11763,N_9521,N_8382);
and U11764 (N_11764,N_8176,N_7986);
and U11765 (N_11765,N_7764,N_9954);
and U11766 (N_11766,N_7870,N_9441);
or U11767 (N_11767,N_9620,N_9339);
or U11768 (N_11768,N_9483,N_8154);
nand U11769 (N_11769,N_8586,N_8743);
and U11770 (N_11770,N_7782,N_9972);
xnor U11771 (N_11771,N_9426,N_8268);
xnor U11772 (N_11772,N_7890,N_9082);
and U11773 (N_11773,N_7792,N_9828);
or U11774 (N_11774,N_8070,N_9552);
nor U11775 (N_11775,N_8369,N_7920);
or U11776 (N_11776,N_8869,N_9144);
nor U11777 (N_11777,N_8826,N_8461);
nor U11778 (N_11778,N_8256,N_9126);
or U11779 (N_11779,N_8489,N_8683);
xor U11780 (N_11780,N_9691,N_9537);
and U11781 (N_11781,N_7703,N_7970);
nand U11782 (N_11782,N_8482,N_7897);
nand U11783 (N_11783,N_7572,N_8874);
nand U11784 (N_11784,N_7843,N_9682);
xor U11785 (N_11785,N_7593,N_8097);
nor U11786 (N_11786,N_8706,N_9813);
nor U11787 (N_11787,N_9227,N_9749);
and U11788 (N_11788,N_9241,N_8218);
nor U11789 (N_11789,N_9532,N_8771);
nand U11790 (N_11790,N_9012,N_8156);
nand U11791 (N_11791,N_9595,N_7880);
or U11792 (N_11792,N_8588,N_9956);
and U11793 (N_11793,N_8272,N_9424);
nand U11794 (N_11794,N_8164,N_9439);
xor U11795 (N_11795,N_9359,N_7809);
and U11796 (N_11796,N_9331,N_8490);
or U11797 (N_11797,N_9414,N_8018);
xor U11798 (N_11798,N_8989,N_8089);
and U11799 (N_11799,N_9164,N_9271);
nor U11800 (N_11800,N_8608,N_9197);
nand U11801 (N_11801,N_9684,N_7647);
or U11802 (N_11802,N_9305,N_8095);
or U11803 (N_11803,N_7900,N_9283);
or U11804 (N_11804,N_8628,N_8235);
and U11805 (N_11805,N_7763,N_9503);
nand U11806 (N_11806,N_7903,N_9136);
nor U11807 (N_11807,N_8942,N_8366);
nor U11808 (N_11808,N_9889,N_9270);
and U11809 (N_11809,N_9800,N_7827);
xnor U11810 (N_11810,N_8910,N_9100);
or U11811 (N_11811,N_7557,N_8394);
nand U11812 (N_11812,N_9993,N_9142);
and U11813 (N_11813,N_9723,N_8815);
and U11814 (N_11814,N_8206,N_9957);
xor U11815 (N_11815,N_9969,N_8977);
nand U11816 (N_11816,N_8094,N_9384);
and U11817 (N_11817,N_7827,N_9604);
xor U11818 (N_11818,N_8967,N_8025);
and U11819 (N_11819,N_8294,N_8815);
or U11820 (N_11820,N_8918,N_9946);
or U11821 (N_11821,N_8470,N_9542);
nand U11822 (N_11822,N_7884,N_9283);
and U11823 (N_11823,N_8737,N_9006);
nand U11824 (N_11824,N_9670,N_7806);
or U11825 (N_11825,N_8342,N_9612);
nand U11826 (N_11826,N_8131,N_8686);
and U11827 (N_11827,N_7811,N_9661);
or U11828 (N_11828,N_8487,N_8415);
xor U11829 (N_11829,N_8610,N_8638);
xor U11830 (N_11830,N_9080,N_7934);
or U11831 (N_11831,N_9260,N_7901);
nand U11832 (N_11832,N_8929,N_8163);
xnor U11833 (N_11833,N_9973,N_9898);
and U11834 (N_11834,N_8113,N_9021);
and U11835 (N_11835,N_9044,N_8999);
and U11836 (N_11836,N_8656,N_8505);
or U11837 (N_11837,N_8030,N_8043);
nand U11838 (N_11838,N_7747,N_9861);
nor U11839 (N_11839,N_9715,N_8152);
or U11840 (N_11840,N_9292,N_9667);
nor U11841 (N_11841,N_9482,N_8353);
nand U11842 (N_11842,N_8019,N_8253);
nor U11843 (N_11843,N_9968,N_7721);
nand U11844 (N_11844,N_7909,N_8127);
nor U11845 (N_11845,N_9937,N_8823);
nand U11846 (N_11846,N_9856,N_8064);
nor U11847 (N_11847,N_8833,N_7979);
and U11848 (N_11848,N_7630,N_7825);
or U11849 (N_11849,N_9159,N_7926);
nor U11850 (N_11850,N_8474,N_8734);
or U11851 (N_11851,N_8284,N_8050);
nand U11852 (N_11852,N_8665,N_8168);
and U11853 (N_11853,N_7917,N_9043);
and U11854 (N_11854,N_8586,N_9098);
nand U11855 (N_11855,N_7881,N_8040);
nor U11856 (N_11856,N_9852,N_7762);
and U11857 (N_11857,N_9655,N_9867);
or U11858 (N_11858,N_9888,N_8740);
xor U11859 (N_11859,N_8633,N_7964);
and U11860 (N_11860,N_9584,N_9964);
xnor U11861 (N_11861,N_8385,N_7580);
and U11862 (N_11862,N_7787,N_8095);
and U11863 (N_11863,N_7755,N_8864);
nor U11864 (N_11864,N_8186,N_8781);
nand U11865 (N_11865,N_7523,N_8129);
nand U11866 (N_11866,N_9143,N_8532);
and U11867 (N_11867,N_7711,N_9792);
nor U11868 (N_11868,N_9061,N_9030);
nand U11869 (N_11869,N_7612,N_7800);
nor U11870 (N_11870,N_7832,N_9193);
nand U11871 (N_11871,N_9390,N_8576);
or U11872 (N_11872,N_8655,N_9581);
nand U11873 (N_11873,N_8598,N_8035);
and U11874 (N_11874,N_8464,N_7758);
or U11875 (N_11875,N_9063,N_9758);
and U11876 (N_11876,N_7746,N_9703);
or U11877 (N_11877,N_9990,N_7730);
and U11878 (N_11878,N_7992,N_7777);
nor U11879 (N_11879,N_8916,N_8944);
nor U11880 (N_11880,N_8703,N_8890);
and U11881 (N_11881,N_8577,N_8731);
xor U11882 (N_11882,N_8897,N_8950);
nor U11883 (N_11883,N_8632,N_9656);
xnor U11884 (N_11884,N_7791,N_7634);
nor U11885 (N_11885,N_7920,N_7709);
nor U11886 (N_11886,N_9251,N_7502);
nand U11887 (N_11887,N_8429,N_8378);
nand U11888 (N_11888,N_9507,N_9494);
or U11889 (N_11889,N_8451,N_7734);
and U11890 (N_11890,N_8202,N_8118);
xnor U11891 (N_11891,N_9341,N_7523);
or U11892 (N_11892,N_8997,N_8933);
xnor U11893 (N_11893,N_8940,N_9775);
and U11894 (N_11894,N_8413,N_7976);
or U11895 (N_11895,N_9342,N_9595);
nor U11896 (N_11896,N_9616,N_8215);
nor U11897 (N_11897,N_8519,N_7556);
nand U11898 (N_11898,N_7565,N_8948);
nor U11899 (N_11899,N_7544,N_8872);
and U11900 (N_11900,N_9418,N_9593);
nand U11901 (N_11901,N_9394,N_7555);
nand U11902 (N_11902,N_8172,N_7947);
and U11903 (N_11903,N_9736,N_8361);
or U11904 (N_11904,N_8921,N_7601);
nor U11905 (N_11905,N_8300,N_7875);
or U11906 (N_11906,N_8216,N_9923);
and U11907 (N_11907,N_9915,N_8872);
and U11908 (N_11908,N_8665,N_8427);
nand U11909 (N_11909,N_8863,N_9785);
nand U11910 (N_11910,N_8751,N_8463);
nand U11911 (N_11911,N_9676,N_9803);
nand U11912 (N_11912,N_9047,N_8509);
and U11913 (N_11913,N_9440,N_7634);
or U11914 (N_11914,N_7939,N_9124);
or U11915 (N_11915,N_9454,N_9933);
and U11916 (N_11916,N_9189,N_8376);
nor U11917 (N_11917,N_8524,N_9932);
nor U11918 (N_11918,N_9546,N_8408);
nand U11919 (N_11919,N_9022,N_7815);
nand U11920 (N_11920,N_9401,N_9070);
nand U11921 (N_11921,N_8473,N_9553);
nand U11922 (N_11922,N_8507,N_8614);
and U11923 (N_11923,N_8380,N_7932);
or U11924 (N_11924,N_9754,N_7918);
or U11925 (N_11925,N_9845,N_8693);
and U11926 (N_11926,N_9748,N_9844);
nand U11927 (N_11927,N_8103,N_9295);
or U11928 (N_11928,N_7771,N_8289);
and U11929 (N_11929,N_9363,N_8083);
nor U11930 (N_11930,N_7770,N_8672);
and U11931 (N_11931,N_8904,N_9656);
nor U11932 (N_11932,N_7825,N_7711);
and U11933 (N_11933,N_9318,N_9652);
and U11934 (N_11934,N_9326,N_7912);
nor U11935 (N_11935,N_8445,N_9166);
nand U11936 (N_11936,N_9209,N_7995);
nor U11937 (N_11937,N_9072,N_8491);
nor U11938 (N_11938,N_8434,N_9366);
nand U11939 (N_11939,N_8654,N_8172);
nand U11940 (N_11940,N_9015,N_8665);
nor U11941 (N_11941,N_7539,N_9445);
or U11942 (N_11942,N_7773,N_9221);
or U11943 (N_11943,N_9343,N_9686);
nor U11944 (N_11944,N_9449,N_8737);
or U11945 (N_11945,N_9925,N_9165);
nand U11946 (N_11946,N_9696,N_8604);
or U11947 (N_11947,N_8825,N_9603);
nand U11948 (N_11948,N_9734,N_7927);
and U11949 (N_11949,N_9338,N_8060);
xor U11950 (N_11950,N_8727,N_8172);
and U11951 (N_11951,N_7557,N_8860);
and U11952 (N_11952,N_7610,N_8267);
or U11953 (N_11953,N_8088,N_9439);
nor U11954 (N_11954,N_8863,N_8353);
xor U11955 (N_11955,N_9505,N_8256);
or U11956 (N_11956,N_7559,N_9652);
or U11957 (N_11957,N_9374,N_8008);
or U11958 (N_11958,N_9804,N_9234);
and U11959 (N_11959,N_9143,N_7714);
nand U11960 (N_11960,N_9571,N_9938);
xor U11961 (N_11961,N_8556,N_8798);
nor U11962 (N_11962,N_9873,N_8466);
nand U11963 (N_11963,N_9790,N_7621);
and U11964 (N_11964,N_8528,N_8748);
nand U11965 (N_11965,N_7792,N_8364);
and U11966 (N_11966,N_9428,N_9100);
nand U11967 (N_11967,N_8195,N_7585);
or U11968 (N_11968,N_8986,N_9324);
nand U11969 (N_11969,N_9787,N_8410);
and U11970 (N_11970,N_8448,N_7877);
or U11971 (N_11971,N_7802,N_9957);
nor U11972 (N_11972,N_8644,N_9167);
or U11973 (N_11973,N_9234,N_9414);
and U11974 (N_11974,N_8894,N_8591);
or U11975 (N_11975,N_9551,N_7642);
nand U11976 (N_11976,N_8065,N_8369);
or U11977 (N_11977,N_7906,N_9617);
nand U11978 (N_11978,N_9303,N_7907);
or U11979 (N_11979,N_8536,N_7849);
nand U11980 (N_11980,N_8980,N_9064);
nor U11981 (N_11981,N_9631,N_7901);
xnor U11982 (N_11982,N_7551,N_8199);
nor U11983 (N_11983,N_9897,N_9926);
nor U11984 (N_11984,N_9013,N_8281);
nand U11985 (N_11985,N_9976,N_7576);
and U11986 (N_11986,N_8952,N_9123);
or U11987 (N_11987,N_8356,N_8086);
and U11988 (N_11988,N_9778,N_7705);
nand U11989 (N_11989,N_8863,N_8923);
or U11990 (N_11990,N_9362,N_7570);
or U11991 (N_11991,N_7985,N_9312);
or U11992 (N_11992,N_8547,N_9322);
or U11993 (N_11993,N_8009,N_9041);
nor U11994 (N_11994,N_9681,N_9505);
nor U11995 (N_11995,N_9555,N_8341);
nor U11996 (N_11996,N_9345,N_7541);
nand U11997 (N_11997,N_8349,N_8818);
and U11998 (N_11998,N_9092,N_8201);
or U11999 (N_11999,N_8341,N_9421);
and U12000 (N_12000,N_7792,N_9339);
and U12001 (N_12001,N_8671,N_9286);
nor U12002 (N_12002,N_9987,N_8732);
nor U12003 (N_12003,N_8548,N_7747);
nand U12004 (N_12004,N_9268,N_8667);
nor U12005 (N_12005,N_9353,N_9939);
nand U12006 (N_12006,N_9885,N_9269);
nand U12007 (N_12007,N_8045,N_7831);
nand U12008 (N_12008,N_8844,N_9020);
and U12009 (N_12009,N_9383,N_7578);
and U12010 (N_12010,N_9982,N_8161);
nand U12011 (N_12011,N_9150,N_9776);
nand U12012 (N_12012,N_9236,N_9374);
or U12013 (N_12013,N_8018,N_7725);
nor U12014 (N_12014,N_8614,N_7529);
or U12015 (N_12015,N_9889,N_9549);
nor U12016 (N_12016,N_9729,N_7620);
or U12017 (N_12017,N_9093,N_9502);
and U12018 (N_12018,N_9010,N_8587);
nor U12019 (N_12019,N_7771,N_8015);
or U12020 (N_12020,N_7772,N_9340);
and U12021 (N_12021,N_8436,N_8044);
nand U12022 (N_12022,N_7895,N_9246);
nor U12023 (N_12023,N_8375,N_9450);
xnor U12024 (N_12024,N_9259,N_7860);
nand U12025 (N_12025,N_9863,N_7964);
and U12026 (N_12026,N_9750,N_8690);
and U12027 (N_12027,N_8207,N_8544);
nor U12028 (N_12028,N_9230,N_8028);
and U12029 (N_12029,N_9692,N_7803);
xor U12030 (N_12030,N_7739,N_9560);
and U12031 (N_12031,N_9400,N_8690);
nor U12032 (N_12032,N_8744,N_9509);
or U12033 (N_12033,N_8588,N_8404);
nor U12034 (N_12034,N_8993,N_9784);
nor U12035 (N_12035,N_9950,N_9892);
nor U12036 (N_12036,N_7791,N_9805);
nand U12037 (N_12037,N_8099,N_8289);
nand U12038 (N_12038,N_7761,N_7807);
or U12039 (N_12039,N_8399,N_8968);
xnor U12040 (N_12040,N_8575,N_9364);
and U12041 (N_12041,N_9485,N_8309);
or U12042 (N_12042,N_7664,N_7935);
nand U12043 (N_12043,N_9237,N_7915);
or U12044 (N_12044,N_9822,N_9616);
nor U12045 (N_12045,N_7686,N_9900);
and U12046 (N_12046,N_7691,N_9551);
and U12047 (N_12047,N_7569,N_8332);
nor U12048 (N_12048,N_7992,N_7553);
xor U12049 (N_12049,N_8876,N_7586);
nor U12050 (N_12050,N_8197,N_9169);
and U12051 (N_12051,N_9347,N_8840);
nor U12052 (N_12052,N_7975,N_7647);
nand U12053 (N_12053,N_8394,N_9459);
and U12054 (N_12054,N_7786,N_9513);
and U12055 (N_12055,N_8037,N_7930);
nand U12056 (N_12056,N_9830,N_9045);
xnor U12057 (N_12057,N_7610,N_9313);
or U12058 (N_12058,N_9485,N_9744);
nor U12059 (N_12059,N_8228,N_9900);
nor U12060 (N_12060,N_7706,N_8683);
xnor U12061 (N_12061,N_9873,N_8325);
nor U12062 (N_12062,N_9016,N_8376);
and U12063 (N_12063,N_7886,N_8034);
nor U12064 (N_12064,N_9362,N_8969);
nor U12065 (N_12065,N_8396,N_9794);
and U12066 (N_12066,N_9783,N_7812);
nand U12067 (N_12067,N_9328,N_9446);
nand U12068 (N_12068,N_9474,N_7840);
nor U12069 (N_12069,N_8715,N_8688);
and U12070 (N_12070,N_9629,N_9108);
nor U12071 (N_12071,N_8476,N_9352);
and U12072 (N_12072,N_8964,N_9717);
nand U12073 (N_12073,N_9267,N_7966);
or U12074 (N_12074,N_8189,N_7735);
nor U12075 (N_12075,N_7850,N_7517);
or U12076 (N_12076,N_7980,N_8442);
nand U12077 (N_12077,N_9424,N_8868);
nor U12078 (N_12078,N_9073,N_9369);
or U12079 (N_12079,N_9533,N_9330);
or U12080 (N_12080,N_8739,N_8119);
xor U12081 (N_12081,N_8301,N_7580);
nand U12082 (N_12082,N_9991,N_9125);
and U12083 (N_12083,N_9998,N_9803);
nor U12084 (N_12084,N_9445,N_8603);
nor U12085 (N_12085,N_8533,N_8514);
and U12086 (N_12086,N_9690,N_9545);
and U12087 (N_12087,N_8015,N_9776);
or U12088 (N_12088,N_9816,N_8170);
and U12089 (N_12089,N_9033,N_9999);
and U12090 (N_12090,N_8331,N_9766);
nand U12091 (N_12091,N_7553,N_8255);
and U12092 (N_12092,N_7922,N_9181);
xor U12093 (N_12093,N_9091,N_7758);
nor U12094 (N_12094,N_9446,N_8635);
and U12095 (N_12095,N_8898,N_9997);
or U12096 (N_12096,N_8483,N_7801);
xnor U12097 (N_12097,N_7744,N_9365);
and U12098 (N_12098,N_8553,N_9410);
and U12099 (N_12099,N_8073,N_8014);
nor U12100 (N_12100,N_8533,N_9651);
nor U12101 (N_12101,N_8302,N_8377);
and U12102 (N_12102,N_7551,N_8004);
or U12103 (N_12103,N_8071,N_8096);
xor U12104 (N_12104,N_9207,N_8928);
nand U12105 (N_12105,N_8988,N_9665);
or U12106 (N_12106,N_8675,N_9402);
nand U12107 (N_12107,N_9875,N_9161);
nor U12108 (N_12108,N_8776,N_9627);
nand U12109 (N_12109,N_8550,N_9826);
and U12110 (N_12110,N_8711,N_9019);
nor U12111 (N_12111,N_7739,N_9479);
or U12112 (N_12112,N_9396,N_9667);
xnor U12113 (N_12113,N_9939,N_8020);
or U12114 (N_12114,N_7513,N_8091);
nor U12115 (N_12115,N_9848,N_8318);
nand U12116 (N_12116,N_9949,N_9425);
or U12117 (N_12117,N_8784,N_9517);
xnor U12118 (N_12118,N_9364,N_9453);
nand U12119 (N_12119,N_9236,N_7760);
nor U12120 (N_12120,N_8344,N_8561);
or U12121 (N_12121,N_7508,N_9882);
and U12122 (N_12122,N_8084,N_8417);
nand U12123 (N_12123,N_7605,N_7733);
nor U12124 (N_12124,N_9648,N_7820);
and U12125 (N_12125,N_8692,N_8599);
and U12126 (N_12126,N_9668,N_9555);
nand U12127 (N_12127,N_7573,N_8191);
nand U12128 (N_12128,N_8632,N_8778);
or U12129 (N_12129,N_8339,N_8845);
nand U12130 (N_12130,N_9556,N_7925);
nand U12131 (N_12131,N_9480,N_9877);
nand U12132 (N_12132,N_8326,N_7597);
or U12133 (N_12133,N_9784,N_7833);
nand U12134 (N_12134,N_7550,N_8958);
nor U12135 (N_12135,N_9927,N_8043);
nand U12136 (N_12136,N_9931,N_8847);
nor U12137 (N_12137,N_8354,N_8127);
xnor U12138 (N_12138,N_8905,N_7593);
nor U12139 (N_12139,N_9900,N_8885);
or U12140 (N_12140,N_7975,N_8225);
and U12141 (N_12141,N_8504,N_7948);
xnor U12142 (N_12142,N_8247,N_8487);
nand U12143 (N_12143,N_8052,N_9702);
nand U12144 (N_12144,N_8557,N_9284);
nand U12145 (N_12145,N_8128,N_8457);
and U12146 (N_12146,N_8544,N_8406);
or U12147 (N_12147,N_8283,N_8194);
xor U12148 (N_12148,N_8786,N_7871);
nand U12149 (N_12149,N_9965,N_8289);
or U12150 (N_12150,N_9029,N_9599);
or U12151 (N_12151,N_9952,N_7830);
nand U12152 (N_12152,N_7964,N_8334);
or U12153 (N_12153,N_8928,N_7772);
or U12154 (N_12154,N_8047,N_8341);
and U12155 (N_12155,N_8047,N_8465);
or U12156 (N_12156,N_9509,N_8959);
nor U12157 (N_12157,N_7925,N_9689);
and U12158 (N_12158,N_7565,N_9414);
nand U12159 (N_12159,N_8516,N_9438);
nand U12160 (N_12160,N_7792,N_8960);
and U12161 (N_12161,N_8097,N_8805);
or U12162 (N_12162,N_8034,N_8579);
nand U12163 (N_12163,N_8141,N_9682);
nor U12164 (N_12164,N_7917,N_8935);
and U12165 (N_12165,N_8392,N_9702);
nor U12166 (N_12166,N_8899,N_9492);
or U12167 (N_12167,N_8705,N_9076);
and U12168 (N_12168,N_8861,N_8756);
and U12169 (N_12169,N_9511,N_8993);
nand U12170 (N_12170,N_9983,N_8547);
nand U12171 (N_12171,N_9651,N_7749);
nor U12172 (N_12172,N_9806,N_9592);
nor U12173 (N_12173,N_9463,N_9253);
nor U12174 (N_12174,N_9730,N_8468);
nor U12175 (N_12175,N_8208,N_8087);
and U12176 (N_12176,N_8020,N_8091);
nor U12177 (N_12177,N_8498,N_8226);
or U12178 (N_12178,N_9457,N_7769);
xnor U12179 (N_12179,N_8421,N_8224);
or U12180 (N_12180,N_8128,N_9718);
xnor U12181 (N_12181,N_7785,N_7506);
or U12182 (N_12182,N_9072,N_9947);
or U12183 (N_12183,N_8585,N_9422);
xor U12184 (N_12184,N_9679,N_8666);
and U12185 (N_12185,N_7801,N_8564);
or U12186 (N_12186,N_7976,N_9581);
nor U12187 (N_12187,N_8618,N_8052);
nand U12188 (N_12188,N_8765,N_7642);
and U12189 (N_12189,N_9614,N_8737);
and U12190 (N_12190,N_8316,N_8947);
nor U12191 (N_12191,N_9476,N_9423);
nand U12192 (N_12192,N_8729,N_8199);
nor U12193 (N_12193,N_8658,N_9591);
nor U12194 (N_12194,N_7872,N_8391);
or U12195 (N_12195,N_9984,N_8444);
nor U12196 (N_12196,N_7883,N_9853);
and U12197 (N_12197,N_8292,N_7942);
and U12198 (N_12198,N_7985,N_8056);
and U12199 (N_12199,N_8135,N_8891);
xnor U12200 (N_12200,N_8411,N_9115);
nand U12201 (N_12201,N_8884,N_9701);
xor U12202 (N_12202,N_7940,N_8747);
and U12203 (N_12203,N_8171,N_9606);
or U12204 (N_12204,N_8739,N_9464);
nand U12205 (N_12205,N_9827,N_8687);
or U12206 (N_12206,N_9122,N_8976);
and U12207 (N_12207,N_8737,N_8861);
or U12208 (N_12208,N_9766,N_8731);
nand U12209 (N_12209,N_9794,N_7691);
xor U12210 (N_12210,N_9089,N_9606);
nand U12211 (N_12211,N_9958,N_9965);
nor U12212 (N_12212,N_8243,N_9191);
or U12213 (N_12213,N_8654,N_9905);
and U12214 (N_12214,N_7755,N_9390);
and U12215 (N_12215,N_8774,N_9170);
xor U12216 (N_12216,N_7662,N_9113);
nand U12217 (N_12217,N_9250,N_8605);
nand U12218 (N_12218,N_8135,N_8193);
or U12219 (N_12219,N_9959,N_7893);
nor U12220 (N_12220,N_9143,N_9237);
and U12221 (N_12221,N_8342,N_9089);
nand U12222 (N_12222,N_9085,N_9083);
or U12223 (N_12223,N_7604,N_8328);
xor U12224 (N_12224,N_8673,N_9047);
nand U12225 (N_12225,N_8959,N_9568);
nand U12226 (N_12226,N_7978,N_8243);
and U12227 (N_12227,N_7990,N_7657);
or U12228 (N_12228,N_8729,N_9193);
xnor U12229 (N_12229,N_7898,N_9288);
nand U12230 (N_12230,N_9542,N_7617);
nor U12231 (N_12231,N_8157,N_8045);
nor U12232 (N_12232,N_8763,N_7758);
nor U12233 (N_12233,N_9905,N_7956);
xor U12234 (N_12234,N_8245,N_9826);
nor U12235 (N_12235,N_9059,N_8864);
nand U12236 (N_12236,N_7691,N_8213);
or U12237 (N_12237,N_8738,N_9065);
nand U12238 (N_12238,N_8459,N_8463);
nand U12239 (N_12239,N_7658,N_7839);
and U12240 (N_12240,N_9788,N_9249);
nand U12241 (N_12241,N_7564,N_7506);
nor U12242 (N_12242,N_9090,N_9422);
or U12243 (N_12243,N_9810,N_9946);
nor U12244 (N_12244,N_8159,N_8373);
nand U12245 (N_12245,N_8869,N_9605);
nand U12246 (N_12246,N_7658,N_8094);
nand U12247 (N_12247,N_8406,N_9752);
xnor U12248 (N_12248,N_9362,N_9034);
and U12249 (N_12249,N_8229,N_8589);
nor U12250 (N_12250,N_9489,N_8009);
nor U12251 (N_12251,N_7741,N_9230);
and U12252 (N_12252,N_9646,N_8232);
or U12253 (N_12253,N_7536,N_8991);
nor U12254 (N_12254,N_9745,N_9441);
or U12255 (N_12255,N_9238,N_8539);
and U12256 (N_12256,N_9806,N_8185);
nor U12257 (N_12257,N_9615,N_9271);
nor U12258 (N_12258,N_8796,N_9334);
and U12259 (N_12259,N_9529,N_7805);
or U12260 (N_12260,N_9574,N_8127);
and U12261 (N_12261,N_9145,N_9509);
or U12262 (N_12262,N_9085,N_9548);
or U12263 (N_12263,N_8397,N_8254);
and U12264 (N_12264,N_9207,N_7567);
and U12265 (N_12265,N_7713,N_9712);
and U12266 (N_12266,N_8564,N_8938);
xnor U12267 (N_12267,N_7752,N_9867);
xnor U12268 (N_12268,N_9925,N_8621);
and U12269 (N_12269,N_7605,N_9154);
nand U12270 (N_12270,N_8154,N_8904);
nor U12271 (N_12271,N_7804,N_8489);
or U12272 (N_12272,N_8784,N_8506);
and U12273 (N_12273,N_9851,N_9388);
xnor U12274 (N_12274,N_9660,N_9603);
nand U12275 (N_12275,N_7785,N_8399);
and U12276 (N_12276,N_8988,N_9530);
and U12277 (N_12277,N_7888,N_8884);
or U12278 (N_12278,N_8576,N_8554);
or U12279 (N_12279,N_9786,N_7579);
or U12280 (N_12280,N_8710,N_8031);
nand U12281 (N_12281,N_9253,N_7559);
or U12282 (N_12282,N_8310,N_9931);
nand U12283 (N_12283,N_7505,N_9443);
nor U12284 (N_12284,N_8950,N_8114);
and U12285 (N_12285,N_7938,N_7945);
nand U12286 (N_12286,N_9448,N_7678);
or U12287 (N_12287,N_7652,N_7836);
nor U12288 (N_12288,N_9162,N_9995);
or U12289 (N_12289,N_8293,N_8355);
xnor U12290 (N_12290,N_9241,N_7943);
or U12291 (N_12291,N_7909,N_7952);
nor U12292 (N_12292,N_8661,N_9661);
nor U12293 (N_12293,N_9373,N_9357);
nand U12294 (N_12294,N_9174,N_9962);
nand U12295 (N_12295,N_9834,N_9596);
nand U12296 (N_12296,N_9220,N_9360);
nor U12297 (N_12297,N_7740,N_8735);
and U12298 (N_12298,N_8860,N_7500);
nand U12299 (N_12299,N_9178,N_9782);
nand U12300 (N_12300,N_7712,N_9484);
and U12301 (N_12301,N_8761,N_8685);
or U12302 (N_12302,N_7758,N_7674);
or U12303 (N_12303,N_9532,N_7963);
and U12304 (N_12304,N_9006,N_8907);
or U12305 (N_12305,N_9938,N_8062);
nor U12306 (N_12306,N_7659,N_8063);
xor U12307 (N_12307,N_9248,N_8530);
or U12308 (N_12308,N_9968,N_9902);
nor U12309 (N_12309,N_9679,N_8914);
or U12310 (N_12310,N_9199,N_9118);
nor U12311 (N_12311,N_9736,N_7762);
and U12312 (N_12312,N_9195,N_9729);
or U12313 (N_12313,N_9401,N_8777);
or U12314 (N_12314,N_8758,N_7557);
and U12315 (N_12315,N_9341,N_7528);
or U12316 (N_12316,N_9329,N_7841);
or U12317 (N_12317,N_9789,N_9493);
nand U12318 (N_12318,N_9352,N_8647);
nand U12319 (N_12319,N_9523,N_8177);
nor U12320 (N_12320,N_9470,N_9821);
nand U12321 (N_12321,N_9009,N_9767);
nor U12322 (N_12322,N_9059,N_8546);
and U12323 (N_12323,N_9986,N_9319);
nor U12324 (N_12324,N_9619,N_9323);
or U12325 (N_12325,N_8078,N_8066);
and U12326 (N_12326,N_8339,N_8400);
nor U12327 (N_12327,N_7640,N_8072);
xor U12328 (N_12328,N_7933,N_7743);
nor U12329 (N_12329,N_9714,N_8829);
and U12330 (N_12330,N_9639,N_8105);
nor U12331 (N_12331,N_9878,N_9489);
xor U12332 (N_12332,N_8029,N_8159);
nand U12333 (N_12333,N_9499,N_8881);
nand U12334 (N_12334,N_9446,N_7518);
and U12335 (N_12335,N_8996,N_9112);
or U12336 (N_12336,N_8252,N_8018);
and U12337 (N_12337,N_8488,N_8110);
or U12338 (N_12338,N_8550,N_8109);
nand U12339 (N_12339,N_9302,N_8294);
and U12340 (N_12340,N_8462,N_8120);
nand U12341 (N_12341,N_7939,N_9364);
and U12342 (N_12342,N_8596,N_9212);
and U12343 (N_12343,N_9822,N_7690);
nor U12344 (N_12344,N_7743,N_8267);
and U12345 (N_12345,N_8385,N_9194);
and U12346 (N_12346,N_9790,N_9243);
nor U12347 (N_12347,N_9479,N_8747);
and U12348 (N_12348,N_9814,N_9412);
or U12349 (N_12349,N_8660,N_9886);
nor U12350 (N_12350,N_9024,N_9499);
nor U12351 (N_12351,N_8175,N_9975);
nor U12352 (N_12352,N_9625,N_8042);
and U12353 (N_12353,N_9732,N_7959);
and U12354 (N_12354,N_8798,N_8489);
or U12355 (N_12355,N_7556,N_9535);
or U12356 (N_12356,N_8854,N_9323);
or U12357 (N_12357,N_9353,N_9351);
nor U12358 (N_12358,N_7522,N_7677);
and U12359 (N_12359,N_9766,N_8381);
nand U12360 (N_12360,N_7773,N_9953);
xor U12361 (N_12361,N_9595,N_9212);
or U12362 (N_12362,N_8617,N_8511);
or U12363 (N_12363,N_8450,N_8560);
or U12364 (N_12364,N_8704,N_8354);
and U12365 (N_12365,N_8536,N_9176);
nor U12366 (N_12366,N_9256,N_8957);
and U12367 (N_12367,N_9517,N_8974);
and U12368 (N_12368,N_8603,N_9345);
or U12369 (N_12369,N_8503,N_9679);
nand U12370 (N_12370,N_9538,N_8598);
and U12371 (N_12371,N_9313,N_8022);
or U12372 (N_12372,N_7629,N_9829);
or U12373 (N_12373,N_7754,N_8573);
and U12374 (N_12374,N_9000,N_9637);
nand U12375 (N_12375,N_7530,N_8621);
nor U12376 (N_12376,N_9578,N_8268);
nand U12377 (N_12377,N_8860,N_9203);
or U12378 (N_12378,N_7567,N_7782);
or U12379 (N_12379,N_8064,N_8233);
nand U12380 (N_12380,N_9054,N_8288);
nand U12381 (N_12381,N_9795,N_8756);
and U12382 (N_12382,N_8175,N_9935);
and U12383 (N_12383,N_9204,N_7882);
nand U12384 (N_12384,N_9802,N_9026);
nand U12385 (N_12385,N_9230,N_9729);
and U12386 (N_12386,N_8224,N_8359);
nor U12387 (N_12387,N_8897,N_9568);
nand U12388 (N_12388,N_8486,N_7991);
and U12389 (N_12389,N_8675,N_9517);
and U12390 (N_12390,N_9184,N_9977);
and U12391 (N_12391,N_7677,N_9944);
nand U12392 (N_12392,N_7574,N_9699);
and U12393 (N_12393,N_9788,N_9005);
nand U12394 (N_12394,N_8305,N_9148);
and U12395 (N_12395,N_9298,N_7529);
nor U12396 (N_12396,N_7951,N_9186);
nor U12397 (N_12397,N_8707,N_8641);
and U12398 (N_12398,N_9989,N_9740);
nand U12399 (N_12399,N_8712,N_8847);
or U12400 (N_12400,N_9318,N_9309);
and U12401 (N_12401,N_8744,N_9586);
or U12402 (N_12402,N_8446,N_8335);
or U12403 (N_12403,N_7949,N_9232);
nor U12404 (N_12404,N_8885,N_9572);
or U12405 (N_12405,N_8500,N_8809);
or U12406 (N_12406,N_8843,N_8837);
nor U12407 (N_12407,N_9093,N_7561);
nand U12408 (N_12408,N_9348,N_7952);
and U12409 (N_12409,N_9814,N_9699);
nand U12410 (N_12410,N_8468,N_8561);
nand U12411 (N_12411,N_9877,N_9127);
nor U12412 (N_12412,N_7916,N_9974);
nand U12413 (N_12413,N_7550,N_7955);
nand U12414 (N_12414,N_9475,N_8135);
nand U12415 (N_12415,N_8440,N_8373);
nor U12416 (N_12416,N_8704,N_7824);
xnor U12417 (N_12417,N_9263,N_8213);
nand U12418 (N_12418,N_8039,N_8421);
and U12419 (N_12419,N_8902,N_7972);
and U12420 (N_12420,N_7797,N_7503);
and U12421 (N_12421,N_7727,N_8568);
and U12422 (N_12422,N_8163,N_8928);
or U12423 (N_12423,N_9591,N_9207);
nand U12424 (N_12424,N_9135,N_9922);
nand U12425 (N_12425,N_9145,N_9439);
and U12426 (N_12426,N_9662,N_8593);
nor U12427 (N_12427,N_9517,N_8914);
nand U12428 (N_12428,N_9191,N_8599);
nand U12429 (N_12429,N_9649,N_9148);
xor U12430 (N_12430,N_8739,N_8814);
or U12431 (N_12431,N_8109,N_9374);
nor U12432 (N_12432,N_9269,N_9020);
nand U12433 (N_12433,N_8220,N_7994);
and U12434 (N_12434,N_9012,N_9210);
nor U12435 (N_12435,N_8466,N_9232);
nor U12436 (N_12436,N_9894,N_8269);
and U12437 (N_12437,N_8432,N_7803);
xor U12438 (N_12438,N_9013,N_9493);
nand U12439 (N_12439,N_8634,N_8912);
nand U12440 (N_12440,N_8961,N_9161);
xnor U12441 (N_12441,N_9944,N_7505);
nand U12442 (N_12442,N_9624,N_9543);
or U12443 (N_12443,N_9677,N_9570);
nand U12444 (N_12444,N_9202,N_8446);
and U12445 (N_12445,N_8359,N_7774);
and U12446 (N_12446,N_7800,N_7886);
nor U12447 (N_12447,N_9110,N_8423);
nor U12448 (N_12448,N_9126,N_8769);
or U12449 (N_12449,N_8163,N_9701);
nor U12450 (N_12450,N_7899,N_8521);
or U12451 (N_12451,N_8379,N_9287);
nand U12452 (N_12452,N_9441,N_8094);
xnor U12453 (N_12453,N_9884,N_9814);
and U12454 (N_12454,N_7901,N_8613);
nor U12455 (N_12455,N_9290,N_7950);
nor U12456 (N_12456,N_7542,N_7844);
or U12457 (N_12457,N_8624,N_8696);
xor U12458 (N_12458,N_9091,N_9942);
and U12459 (N_12459,N_8946,N_9272);
and U12460 (N_12460,N_7821,N_8929);
nand U12461 (N_12461,N_9012,N_7961);
nor U12462 (N_12462,N_7520,N_7688);
or U12463 (N_12463,N_9971,N_8349);
nor U12464 (N_12464,N_7717,N_8700);
and U12465 (N_12465,N_8728,N_9233);
nor U12466 (N_12466,N_9934,N_7885);
xor U12467 (N_12467,N_9387,N_9392);
nand U12468 (N_12468,N_9601,N_9218);
nor U12469 (N_12469,N_8151,N_9523);
nor U12470 (N_12470,N_8640,N_8677);
nor U12471 (N_12471,N_9722,N_8929);
or U12472 (N_12472,N_7815,N_9976);
or U12473 (N_12473,N_8408,N_9003);
and U12474 (N_12474,N_9064,N_9608);
nand U12475 (N_12475,N_8436,N_7910);
and U12476 (N_12476,N_7805,N_7571);
nor U12477 (N_12477,N_8707,N_9579);
and U12478 (N_12478,N_8342,N_7641);
xor U12479 (N_12479,N_9959,N_9313);
or U12480 (N_12480,N_9738,N_9210);
and U12481 (N_12481,N_7784,N_7521);
or U12482 (N_12482,N_9754,N_9460);
nand U12483 (N_12483,N_8713,N_9371);
nand U12484 (N_12484,N_9678,N_8318);
nand U12485 (N_12485,N_9971,N_7620);
or U12486 (N_12486,N_9643,N_9577);
and U12487 (N_12487,N_9418,N_8900);
xor U12488 (N_12488,N_8446,N_9931);
nor U12489 (N_12489,N_8695,N_9016);
and U12490 (N_12490,N_8435,N_9190);
or U12491 (N_12491,N_9313,N_8555);
or U12492 (N_12492,N_8930,N_8159);
and U12493 (N_12493,N_9029,N_8103);
nor U12494 (N_12494,N_9047,N_9919);
or U12495 (N_12495,N_8422,N_8604);
and U12496 (N_12496,N_8062,N_9760);
or U12497 (N_12497,N_8086,N_9352);
xor U12498 (N_12498,N_9080,N_8968);
xnor U12499 (N_12499,N_8055,N_9042);
nor U12500 (N_12500,N_11088,N_10355);
nor U12501 (N_12501,N_10178,N_10540);
and U12502 (N_12502,N_12365,N_12383);
and U12503 (N_12503,N_10060,N_10972);
nand U12504 (N_12504,N_10322,N_11074);
and U12505 (N_12505,N_12458,N_10410);
and U12506 (N_12506,N_11060,N_10112);
nor U12507 (N_12507,N_10854,N_10721);
nor U12508 (N_12508,N_10234,N_10361);
nand U12509 (N_12509,N_11653,N_11661);
and U12510 (N_12510,N_11900,N_10369);
nand U12511 (N_12511,N_11085,N_11997);
nor U12512 (N_12512,N_10671,N_10706);
or U12513 (N_12513,N_12133,N_10826);
nor U12514 (N_12514,N_11110,N_10453);
and U12515 (N_12515,N_11474,N_11890);
or U12516 (N_12516,N_12354,N_10227);
nor U12517 (N_12517,N_10358,N_12465);
or U12518 (N_12518,N_11546,N_10067);
nor U12519 (N_12519,N_12497,N_10742);
xor U12520 (N_12520,N_12186,N_10160);
or U12521 (N_12521,N_11993,N_11589);
and U12522 (N_12522,N_10249,N_12243);
and U12523 (N_12523,N_11510,N_11848);
nand U12524 (N_12524,N_12041,N_11933);
xor U12525 (N_12525,N_11023,N_11999);
or U12526 (N_12526,N_10836,N_10535);
nor U12527 (N_12527,N_11923,N_11822);
nor U12528 (N_12528,N_10162,N_12000);
nor U12529 (N_12529,N_10474,N_10376);
and U12530 (N_12530,N_11639,N_11111);
or U12531 (N_12531,N_11073,N_11606);
nor U12532 (N_12532,N_12270,N_11836);
nor U12533 (N_12533,N_11150,N_10277);
nand U12534 (N_12534,N_11191,N_11942);
or U12535 (N_12535,N_11753,N_10991);
nor U12536 (N_12536,N_12391,N_12217);
xor U12537 (N_12537,N_10538,N_11938);
nor U12538 (N_12538,N_10737,N_10301);
nor U12539 (N_12539,N_12165,N_10248);
nand U12540 (N_12540,N_12091,N_12099);
nand U12541 (N_12541,N_12107,N_11185);
or U12542 (N_12542,N_12152,N_11283);
nand U12543 (N_12543,N_12216,N_11193);
or U12544 (N_12544,N_10900,N_10800);
nand U12545 (N_12545,N_10835,N_10061);
or U12546 (N_12546,N_11956,N_11662);
nor U12547 (N_12547,N_11806,N_11791);
and U12548 (N_12548,N_12213,N_11083);
or U12549 (N_12549,N_11790,N_11537);
nand U12550 (N_12550,N_11882,N_11686);
nand U12551 (N_12551,N_12321,N_10755);
nand U12552 (N_12552,N_10000,N_11061);
nand U12553 (N_12553,N_10255,N_11608);
and U12554 (N_12554,N_11226,N_12271);
nand U12555 (N_12555,N_12238,N_10016);
or U12556 (N_12556,N_10774,N_11135);
or U12557 (N_12557,N_11106,N_12159);
or U12558 (N_12558,N_11990,N_10638);
and U12559 (N_12559,N_10910,N_12418);
xnor U12560 (N_12560,N_11177,N_11550);
nor U12561 (N_12561,N_11136,N_12318);
nand U12562 (N_12562,N_10089,N_12363);
nand U12563 (N_12563,N_12495,N_12007);
or U12564 (N_12564,N_11208,N_11300);
xor U12565 (N_12565,N_11406,N_11077);
nand U12566 (N_12566,N_11292,N_11936);
nand U12567 (N_12567,N_10065,N_12226);
xor U12568 (N_12568,N_12036,N_10864);
nor U12569 (N_12569,N_12313,N_11098);
nor U12570 (N_12570,N_12305,N_10004);
and U12571 (N_12571,N_10346,N_11994);
and U12572 (N_12572,N_11582,N_11964);
xnor U12573 (N_12573,N_11097,N_11216);
or U12574 (N_12574,N_11047,N_11579);
xor U12575 (N_12575,N_11909,N_10181);
or U12576 (N_12576,N_12320,N_12436);
and U12577 (N_12577,N_10261,N_11667);
or U12578 (N_12578,N_10224,N_12035);
and U12579 (N_12579,N_11858,N_11516);
and U12580 (N_12580,N_10914,N_10423);
or U12581 (N_12581,N_11812,N_11838);
nor U12582 (N_12582,N_10812,N_11275);
nor U12583 (N_12583,N_12442,N_10516);
and U12584 (N_12584,N_11988,N_12249);
nor U12585 (N_12585,N_12125,N_12002);
or U12586 (N_12586,N_10977,N_11834);
and U12587 (N_12587,N_10806,N_12443);
and U12588 (N_12588,N_10201,N_10300);
nand U12589 (N_12589,N_12204,N_10649);
xor U12590 (N_12590,N_12482,N_11198);
nor U12591 (N_12591,N_11278,N_10905);
nand U12592 (N_12592,N_12116,N_10834);
and U12593 (N_12593,N_12473,N_12046);
or U12594 (N_12594,N_10623,N_11257);
nand U12595 (N_12595,N_10370,N_10487);
and U12596 (N_12596,N_10215,N_11774);
nand U12597 (N_12597,N_11396,N_10558);
nor U12598 (N_12598,N_11468,N_10293);
and U12599 (N_12599,N_11799,N_10982);
and U12600 (N_12600,N_12026,N_10012);
or U12601 (N_12601,N_10377,N_11056);
and U12602 (N_12602,N_11603,N_12456);
or U12603 (N_12603,N_11425,N_11392);
nand U12604 (N_12604,N_10003,N_11120);
nand U12605 (N_12605,N_11766,N_10734);
and U12606 (N_12606,N_11495,N_10843);
nor U12607 (N_12607,N_11915,N_12013);
nor U12608 (N_12608,N_11916,N_10190);
or U12609 (N_12609,N_11013,N_10125);
or U12610 (N_12610,N_12054,N_10478);
and U12611 (N_12611,N_12498,N_11497);
or U12612 (N_12612,N_12156,N_11052);
and U12613 (N_12613,N_12359,N_11144);
nor U12614 (N_12614,N_11003,N_10849);
nor U12615 (N_12615,N_11381,N_12150);
or U12616 (N_12616,N_11683,N_12267);
and U12617 (N_12617,N_10165,N_11911);
nor U12618 (N_12618,N_12220,N_10463);
or U12619 (N_12619,N_10552,N_10015);
and U12620 (N_12620,N_12306,N_10999);
or U12621 (N_12621,N_11006,N_10429);
or U12622 (N_12622,N_12101,N_11256);
and U12623 (N_12623,N_10996,N_11351);
nor U12624 (N_12624,N_11154,N_10640);
nor U12625 (N_12625,N_12048,N_12329);
and U12626 (N_12626,N_10861,N_10823);
nor U12627 (N_12627,N_10564,N_10940);
nand U12628 (N_12628,N_10509,N_10536);
and U12629 (N_12629,N_10484,N_11318);
and U12630 (N_12630,N_11984,N_10339);
and U12631 (N_12631,N_12176,N_10163);
nor U12632 (N_12632,N_11100,N_11702);
and U12633 (N_12633,N_11225,N_11122);
nand U12634 (N_12634,N_11731,N_11515);
xor U12635 (N_12635,N_11271,N_11575);
nand U12636 (N_12636,N_10334,N_12457);
or U12637 (N_12637,N_10508,N_10643);
nand U12638 (N_12638,N_11688,N_11941);
xnor U12639 (N_12639,N_11040,N_11002);
or U12640 (N_12640,N_10777,N_10754);
and U12641 (N_12641,N_11780,N_11247);
nand U12642 (N_12642,N_10064,N_12407);
nand U12643 (N_12643,N_12235,N_10967);
or U12644 (N_12644,N_11856,N_11801);
or U12645 (N_12645,N_10519,N_11531);
and U12646 (N_12646,N_11659,N_10827);
or U12647 (N_12647,N_11195,N_11146);
nor U12648 (N_12648,N_12103,N_12045);
nor U12649 (N_12649,N_11031,N_12352);
and U12650 (N_12650,N_10867,N_11709);
or U12651 (N_12651,N_10135,N_11179);
and U12652 (N_12652,N_11730,N_12266);
nor U12653 (N_12653,N_10081,N_10466);
and U12654 (N_12654,N_10185,N_10929);
xnor U12655 (N_12655,N_10032,N_12346);
nand U12656 (N_12656,N_11249,N_10784);
or U12657 (N_12657,N_11205,N_12301);
nand U12658 (N_12658,N_10889,N_12492);
and U12659 (N_12659,N_12315,N_11412);
and U12660 (N_12660,N_10657,N_12302);
nand U12661 (N_12661,N_12043,N_11171);
or U12662 (N_12662,N_11034,N_12039);
or U12663 (N_12663,N_11761,N_12114);
or U12664 (N_12664,N_10550,N_12225);
and U12665 (N_12665,N_11348,N_10225);
nor U12666 (N_12666,N_10086,N_11927);
or U12667 (N_12667,N_11674,N_12371);
and U12668 (N_12668,N_11959,N_10507);
nand U12669 (N_12669,N_10979,N_10988);
xor U12670 (N_12670,N_10351,N_11728);
nand U12671 (N_12671,N_11295,N_11151);
nor U12672 (N_12672,N_10302,N_11305);
or U12673 (N_12673,N_10359,N_11631);
and U12674 (N_12674,N_11926,N_10780);
and U12675 (N_12675,N_11370,N_10560);
or U12676 (N_12676,N_10476,N_10108);
nor U12677 (N_12677,N_11420,N_11543);
xnor U12678 (N_12678,N_10960,N_11680);
xor U12679 (N_12679,N_11068,N_10821);
nand U12680 (N_12680,N_12239,N_12332);
nor U12681 (N_12681,N_11624,N_12069);
nand U12682 (N_12682,N_10819,N_11798);
or U12683 (N_12683,N_10647,N_11033);
or U12684 (N_12684,N_10354,N_10303);
nor U12685 (N_12685,N_11540,N_11996);
and U12686 (N_12686,N_12262,N_12471);
or U12687 (N_12687,N_12277,N_10214);
and U12688 (N_12688,N_10707,N_11227);
nor U12689 (N_12689,N_10439,N_10789);
or U12690 (N_12690,N_11020,N_11042);
and U12691 (N_12691,N_10438,N_10842);
and U12692 (N_12692,N_12343,N_10412);
nor U12693 (N_12693,N_11689,N_11839);
nand U12694 (N_12694,N_11391,N_10934);
nor U12695 (N_12695,N_11493,N_11706);
or U12696 (N_12696,N_12205,N_10013);
or U12697 (N_12697,N_11867,N_10176);
or U12698 (N_12698,N_10686,N_10228);
or U12699 (N_12699,N_10001,N_10347);
nor U12700 (N_12700,N_10983,N_10936);
and U12701 (N_12701,N_11449,N_11025);
xnor U12702 (N_12702,N_10571,N_12160);
and U12703 (N_12703,N_10697,N_10039);
and U12704 (N_12704,N_10318,N_11700);
or U12705 (N_12705,N_10986,N_12233);
nand U12706 (N_12706,N_11105,N_11324);
and U12707 (N_12707,N_10714,N_10383);
nor U12708 (N_12708,N_11924,N_11577);
nand U12709 (N_12709,N_10437,N_10824);
and U12710 (N_12710,N_10222,N_10129);
nand U12711 (N_12711,N_10947,N_11478);
or U12712 (N_12712,N_11437,N_10079);
nand U12713 (N_12713,N_11560,N_11981);
and U12714 (N_12714,N_10847,N_11765);
and U12715 (N_12715,N_10455,N_11347);
or U12716 (N_12716,N_10544,N_10943);
xnor U12717 (N_12717,N_12276,N_10033);
xor U12718 (N_12718,N_10692,N_10964);
nand U12719 (N_12719,N_11423,N_11861);
and U12720 (N_12720,N_11831,N_10087);
or U12721 (N_12721,N_10773,N_11768);
and U12722 (N_12722,N_10402,N_10586);
or U12723 (N_12723,N_10975,N_10481);
and U12724 (N_12724,N_12435,N_10570);
nor U12725 (N_12725,N_11116,N_11413);
or U12726 (N_12726,N_11431,N_10750);
nand U12727 (N_12727,N_11695,N_11711);
and U12728 (N_12728,N_11961,N_11571);
and U12729 (N_12729,N_10050,N_11417);
xnor U12730 (N_12730,N_10759,N_11217);
nor U12731 (N_12731,N_10950,N_10246);
and U12732 (N_12732,N_10329,N_10708);
and U12733 (N_12733,N_10209,N_10684);
or U12734 (N_12734,N_11279,N_11665);
and U12735 (N_12735,N_12119,N_10080);
nor U12736 (N_12736,N_10328,N_12199);
and U12737 (N_12737,N_10433,N_11937);
nor U12738 (N_12738,N_10593,N_10096);
nand U12739 (N_12739,N_11809,N_11590);
xnor U12740 (N_12740,N_12222,N_12406);
xor U12741 (N_12741,N_12410,N_10186);
nor U12742 (N_12742,N_10631,N_10730);
and U12743 (N_12743,N_11841,N_11134);
nand U12744 (N_12744,N_11573,N_11645);
nor U12745 (N_12745,N_12058,N_10391);
nor U12746 (N_12746,N_12399,N_11276);
or U12747 (N_12747,N_10617,N_10524);
or U12748 (N_12748,N_11340,N_11137);
nand U12749 (N_12749,N_10511,N_10938);
nor U12750 (N_12750,N_10212,N_10633);
or U12751 (N_12751,N_12335,N_11949);
or U12752 (N_12752,N_10898,N_10296);
nor U12753 (N_12753,N_11737,N_11810);
or U12754 (N_12754,N_12430,N_11285);
or U12755 (N_12755,N_10933,N_10373);
or U12756 (N_12756,N_10174,N_12016);
xor U12757 (N_12757,N_10634,N_12398);
nand U12758 (N_12758,N_10574,N_12342);
xor U12759 (N_12759,N_10287,N_11732);
and U12760 (N_12760,N_12072,N_12179);
nand U12761 (N_12761,N_12449,N_11476);
and U12762 (N_12762,N_11442,N_11363);
or U12763 (N_12763,N_12193,N_11299);
or U12764 (N_12764,N_10153,N_10217);
and U12765 (N_12765,N_11749,N_10349);
nand U12766 (N_12766,N_10281,N_11618);
and U12767 (N_12767,N_11201,N_10501);
and U12768 (N_12768,N_10409,N_11830);
nand U12769 (N_12769,N_11113,N_10625);
nand U12770 (N_12770,N_10588,N_12139);
nand U12771 (N_12771,N_11405,N_10314);
nor U12772 (N_12772,N_11188,N_12129);
or U12773 (N_12773,N_12162,N_12453);
nand U12774 (N_12774,N_11508,N_10198);
nor U12775 (N_12775,N_10589,N_12314);
nor U12776 (N_12776,N_11629,N_11311);
nand U12777 (N_12777,N_10719,N_10873);
nor U12778 (N_12778,N_10703,N_12023);
nor U12779 (N_12779,N_10711,N_11585);
or U12780 (N_12780,N_10792,N_11147);
and U12781 (N_12781,N_12260,N_10532);
nand U12782 (N_12782,N_10817,N_11204);
nor U12783 (N_12783,N_10260,N_10272);
or U12784 (N_12784,N_11199,N_10493);
or U12785 (N_12785,N_12396,N_10610);
nor U12786 (N_12786,N_12182,N_10702);
nand U12787 (N_12787,N_10472,N_10119);
or U12788 (N_12788,N_10419,N_11059);
or U12789 (N_12789,N_11072,N_11840);
nor U12790 (N_12790,N_10971,N_12288);
or U12791 (N_12791,N_10688,N_10912);
or U12792 (N_12792,N_12463,N_11473);
and U12793 (N_12793,N_10392,N_10059);
or U12794 (N_12794,N_12382,N_12309);
or U12795 (N_12795,N_11887,N_10642);
or U12796 (N_12796,N_11600,N_12296);
or U12797 (N_12797,N_11635,N_11281);
and U12798 (N_12798,N_12229,N_11443);
and U12799 (N_12799,N_10595,N_10115);
or U12800 (N_12800,N_12474,N_11763);
xnor U12801 (N_12801,N_11559,N_11738);
nand U12802 (N_12802,N_10521,N_11187);
nand U12803 (N_12803,N_11399,N_11541);
or U12804 (N_12804,N_12368,N_12251);
nor U12805 (N_12805,N_11658,N_10627);
and U12806 (N_12806,N_12416,N_10539);
and U12807 (N_12807,N_11597,N_11913);
or U12808 (N_12808,N_12118,N_12149);
nand U12809 (N_12809,N_10626,N_12020);
nand U12810 (N_12810,N_12250,N_10191);
nor U12811 (N_12811,N_11237,N_11162);
or U12812 (N_12812,N_11696,N_11610);
xnor U12813 (N_12813,N_11676,N_10598);
nor U12814 (N_12814,N_10778,N_11844);
nor U12815 (N_12815,N_10751,N_12340);
and U12816 (N_12816,N_10799,N_10208);
nand U12817 (N_12817,N_11084,N_11044);
nand U12818 (N_12818,N_11668,N_12059);
and U12819 (N_12819,N_10257,N_10909);
nor U12820 (N_12820,N_12247,N_11232);
nor U12821 (N_12821,N_10636,N_12010);
nor U12822 (N_12822,N_10757,N_10324);
or U12823 (N_12823,N_12467,N_11192);
or U12824 (N_12824,N_11465,N_10200);
nor U12825 (N_12825,N_10607,N_11734);
xnor U12826 (N_12826,N_12254,N_10426);
or U12827 (N_12827,N_11868,N_10746);
and U12828 (N_12828,N_12263,N_11982);
nand U12829 (N_12829,N_10575,N_10653);
and U12830 (N_12830,N_11236,N_10483);
nand U12831 (N_12831,N_10099,N_12331);
nand U12832 (N_12832,N_12494,N_11733);
and U12833 (N_12833,N_11682,N_11636);
and U12834 (N_12834,N_11595,N_11194);
or U12835 (N_12835,N_11190,N_10116);
nand U12836 (N_12836,N_10105,N_11058);
nand U12837 (N_12837,N_10913,N_11357);
nor U12838 (N_12838,N_11325,N_10791);
or U12839 (N_12839,N_11458,N_12029);
nor U12840 (N_12840,N_12274,N_10815);
and U12841 (N_12841,N_12292,N_11677);
nor U12842 (N_12842,N_11991,N_10689);
and U12843 (N_12843,N_10283,N_12395);
or U12844 (N_12844,N_12174,N_10019);
and U12845 (N_12845,N_11892,N_10504);
and U12846 (N_12846,N_11078,N_12081);
or U12847 (N_12847,N_10926,N_10146);
and U12848 (N_12848,N_11019,N_12245);
nand U12849 (N_12849,N_11588,N_10935);
and U12850 (N_12850,N_12154,N_11436);
nor U12851 (N_12851,N_11920,N_11419);
or U12852 (N_12852,N_11317,N_12481);
nand U12853 (N_12853,N_11342,N_10698);
or U12854 (N_12854,N_10590,N_11714);
nand U12855 (N_12855,N_10366,N_10077);
or U12856 (N_12856,N_10963,N_11211);
nor U12857 (N_12857,N_10704,N_10136);
nand U12858 (N_12858,N_10522,N_11005);
nand U12859 (N_12859,N_10282,N_11845);
nand U12860 (N_12860,N_10054,N_11323);
and U12861 (N_12861,N_10262,N_10883);
xnor U12862 (N_12862,N_10656,N_11592);
or U12863 (N_12863,N_10247,N_10400);
nor U12864 (N_12864,N_11263,N_11966);
nand U12865 (N_12865,N_10903,N_10030);
and U12866 (N_12866,N_11395,N_10078);
or U12867 (N_12867,N_10490,N_10011);
and U12868 (N_12868,N_11759,N_12454);
or U12869 (N_12869,N_12164,N_11879);
xnor U12870 (N_12870,N_10609,N_10491);
nor U12871 (N_12871,N_10743,N_12316);
and U12872 (N_12872,N_10599,N_10342);
xor U12873 (N_12873,N_11037,N_12202);
and U12874 (N_12874,N_10546,N_12240);
and U12875 (N_12875,N_10641,N_11244);
nand U12876 (N_12876,N_11385,N_11306);
nor U12877 (N_12877,N_10145,N_11029);
and U12878 (N_12878,N_12464,N_11980);
or U12879 (N_12879,N_11625,N_12180);
and U12880 (N_12880,N_11905,N_10131);
or U12881 (N_12881,N_10930,N_10434);
or U12882 (N_12882,N_12163,N_11617);
nor U12883 (N_12883,N_10594,N_11017);
and U12884 (N_12884,N_12001,N_11955);
nor U12885 (N_12885,N_11254,N_11987);
nand U12886 (N_12886,N_11943,N_10411);
and U12887 (N_12887,N_10388,N_10492);
or U12888 (N_12888,N_10729,N_11697);
nor U12889 (N_12889,N_10427,N_11796);
nand U12890 (N_12890,N_12362,N_10278);
or U12891 (N_12891,N_12079,N_12447);
nor U12892 (N_12892,N_10728,N_10874);
and U12893 (N_12893,N_10562,N_12369);
nand U12894 (N_12894,N_11335,N_10111);
or U12895 (N_12895,N_10194,N_12378);
and U12896 (N_12896,N_10658,N_12095);
or U12897 (N_12897,N_11649,N_10858);
nor U12898 (N_12898,N_12145,N_11024);
nand U12899 (N_12899,N_10583,N_10235);
or U12900 (N_12900,N_12361,N_11679);
nand U12901 (N_12901,N_11633,N_12425);
and U12902 (N_12902,N_11583,N_11322);
nand U12903 (N_12903,N_10263,N_11609);
nor U12904 (N_12904,N_11654,N_12433);
xor U12905 (N_12905,N_10807,N_12319);
or U12906 (N_12906,N_11398,N_12488);
nand U12907 (N_12907,N_11301,N_11424);
and U12908 (N_12908,N_11175,N_10431);
nor U12909 (N_12909,N_11934,N_11563);
or U12910 (N_12910,N_11797,N_11509);
nor U12911 (N_12911,N_11549,N_11466);
or U12912 (N_12912,N_11358,N_11641);
nand U12913 (N_12913,N_12469,N_11165);
or U12914 (N_12914,N_12144,N_10094);
and U12915 (N_12915,N_11647,N_10315);
nor U12916 (N_12916,N_11373,N_10592);
or U12917 (N_12917,N_12140,N_11026);
or U12918 (N_12918,N_12006,N_11284);
nand U12919 (N_12919,N_10870,N_10816);
nor U12920 (N_12920,N_10371,N_12042);
and U12921 (N_12921,N_11561,N_12431);
or U12922 (N_12922,N_10258,N_12307);
nor U12923 (N_12923,N_10350,N_11555);
nand U12924 (N_12924,N_12078,N_10987);
nor U12925 (N_12925,N_11758,N_11650);
nand U12926 (N_12926,N_10572,N_10223);
and U12927 (N_12927,N_11070,N_12293);
nand U12928 (N_12928,N_10374,N_11393);
nor U12929 (N_12929,N_11849,N_11611);
nor U12930 (N_12930,N_10970,N_12137);
nor U12931 (N_12931,N_10863,N_11788);
nand U12932 (N_12932,N_11881,N_11157);
nand U12933 (N_12933,N_11804,N_11908);
or U12934 (N_12934,N_10764,N_10752);
xnor U12935 (N_12935,N_11713,N_10269);
and U12936 (N_12936,N_10783,N_11729);
nor U12937 (N_12937,N_10868,N_10547);
and U12938 (N_12938,N_11820,N_11904);
nor U12939 (N_12939,N_11968,N_11371);
nand U12940 (N_12940,N_10210,N_11535);
or U12941 (N_12941,N_10932,N_11197);
nand U12942 (N_12942,N_10798,N_11341);
and U12943 (N_12943,N_12478,N_11846);
and U12944 (N_12944,N_11369,N_11664);
xor U12945 (N_12945,N_10820,N_10955);
or U12946 (N_12946,N_10219,N_11894);
nand U12947 (N_12947,N_11490,N_11748);
nor U12948 (N_12948,N_12066,N_12085);
or U12949 (N_12949,N_10968,N_10668);
or U12950 (N_12950,N_10906,N_11117);
xor U12951 (N_12951,N_10330,N_11489);
or U12952 (N_12952,N_10839,N_10533);
or U12953 (N_12953,N_12234,N_10712);
or U12954 (N_12954,N_11539,N_11422);
nor U12955 (N_12955,N_12445,N_11015);
nand U12956 (N_12956,N_12192,N_11945);
nand U12957 (N_12957,N_10083,N_12067);
and U12958 (N_12958,N_11651,N_12232);
nor U12959 (N_12959,N_12284,N_11932);
nand U12960 (N_12960,N_11901,N_10601);
xnor U12961 (N_12961,N_12344,N_10762);
or U12962 (N_12962,N_11605,N_11222);
nor U12963 (N_12963,N_11149,N_10994);
nor U12964 (N_12964,N_10279,N_11621);
or U12965 (N_12965,N_10242,N_11977);
nand U12966 (N_12966,N_10606,N_12452);
nor U12967 (N_12967,N_11627,N_10961);
nor U12968 (N_12968,N_12477,N_10949);
nand U12969 (N_12969,N_10159,N_10573);
nand U12970 (N_12970,N_12051,N_11666);
nor U12971 (N_12971,N_10082,N_10152);
and U12972 (N_12972,N_10788,N_10515);
nand U12973 (N_12973,N_11402,N_11902);
nand U12974 (N_12974,N_12466,N_12328);
and U12975 (N_12975,N_11067,N_10265);
or U12976 (N_12976,N_10090,N_10488);
nand U12977 (N_12977,N_10180,N_10167);
or U12978 (N_12978,N_10962,N_10537);
nor U12979 (N_12979,N_12224,N_10694);
and U12980 (N_12980,N_12387,N_12283);
or U12981 (N_12981,N_12185,N_11958);
or U12982 (N_12982,N_10226,N_12255);
and U12983 (N_12983,N_12201,N_10758);
or U12984 (N_12984,N_10477,N_10899);
nand U12985 (N_12985,N_10204,N_11401);
and U12986 (N_12986,N_10884,N_11764);
nand U12987 (N_12987,N_10304,N_10266);
nor U12988 (N_12988,N_10875,N_10232);
xor U12989 (N_12989,N_10763,N_10475);
or U12990 (N_12990,N_10063,N_12389);
and U12991 (N_12991,N_11862,N_11124);
nand U12992 (N_12992,N_11407,N_11599);
or U12993 (N_12993,N_10765,N_10298);
nor U12994 (N_12994,N_10252,N_11715);
xor U12995 (N_12995,N_12211,N_10271);
nand U12996 (N_12996,N_12261,N_10313);
xnor U12997 (N_12997,N_10319,N_11289);
nor U12998 (N_12998,N_12022,N_10299);
nand U12999 (N_12999,N_11139,N_10288);
and U13000 (N_13000,N_12134,N_11978);
nand U13001 (N_13001,N_10628,N_10352);
or U13002 (N_13002,N_12088,N_11513);
nand U13003 (N_13003,N_10976,N_10744);
and U13004 (N_13004,N_10776,N_10678);
and U13005 (N_13005,N_12440,N_12325);
and U13006 (N_13006,N_12166,N_12275);
nand U13007 (N_13007,N_11346,N_11467);
xor U13008 (N_13008,N_11152,N_10142);
or U13009 (N_13009,N_12244,N_10646);
nor U13010 (N_13010,N_11526,N_10520);
nand U13011 (N_13011,N_12380,N_10654);
and U13012 (N_13012,N_11946,N_11308);
and U13013 (N_13013,N_10958,N_10985);
or U13014 (N_13014,N_12090,N_10379);
or U13015 (N_13015,N_11440,N_10026);
xor U13016 (N_13016,N_12015,N_10221);
nor U13017 (N_13017,N_12050,N_10100);
nand U13018 (N_13018,N_10681,N_11218);
nand U13019 (N_13019,N_11027,N_11228);
and U13020 (N_13020,N_10893,N_11307);
nand U13021 (N_13021,N_12138,N_11757);
nand U13022 (N_13022,N_12167,N_10422);
xor U13023 (N_13023,N_10326,N_11523);
or U13024 (N_13024,N_10771,N_11094);
or U13025 (N_13025,N_10097,N_11062);
and U13026 (N_13026,N_10605,N_10580);
and U13027 (N_13027,N_12074,N_12409);
nand U13028 (N_13028,N_11456,N_12087);
or U13029 (N_13029,N_11525,N_12092);
or U13030 (N_13030,N_10023,N_10937);
xor U13031 (N_13031,N_12366,N_12019);
or U13032 (N_13032,N_11505,N_11562);
nor U13033 (N_13033,N_12056,N_10761);
and U13034 (N_13034,N_10890,N_10723);
nor U13035 (N_13035,N_10556,N_10505);
nand U13036 (N_13036,N_10327,N_11917);
or U13037 (N_13037,N_11903,N_11542);
or U13038 (N_13038,N_10407,N_11008);
and U13039 (N_13039,N_10057,N_11206);
and U13040 (N_13040,N_11328,N_11260);
xor U13041 (N_13041,N_11972,N_10885);
nand U13042 (N_13042,N_10157,N_10622);
nor U13043 (N_13043,N_10333,N_12063);
and U13044 (N_13044,N_10665,N_11004);
and U13045 (N_13045,N_10245,N_10291);
nor U13046 (N_13046,N_11368,N_12060);
or U13047 (N_13047,N_11771,N_12476);
nor U13048 (N_13048,N_10796,N_10741);
nor U13049 (N_13049,N_12127,N_11891);
xnor U13050 (N_13050,N_10687,N_12394);
and U13051 (N_13051,N_12038,N_12040);
and U13052 (N_13052,N_10276,N_10479);
nand U13053 (N_13053,N_10486,N_10393);
or U13054 (N_13054,N_12148,N_11326);
nand U13055 (N_13055,N_10496,N_12128);
or U13056 (N_13056,N_11703,N_11114);
and U13057 (N_13057,N_10196,N_12397);
nor U13058 (N_13058,N_10344,N_12073);
or U13059 (N_13059,N_10017,N_11158);
nand U13060 (N_13060,N_11871,N_11294);
and U13061 (N_13061,N_11472,N_11258);
and U13062 (N_13062,N_11316,N_11051);
nand U13063 (N_13063,N_10154,N_11378);
nor U13064 (N_13064,N_10218,N_11947);
or U13065 (N_13065,N_10335,N_11817);
xnor U13066 (N_13066,N_11320,N_10139);
xor U13067 (N_13067,N_10772,N_11604);
nor U13068 (N_13068,N_11238,N_12280);
or U13069 (N_13069,N_11414,N_11906);
and U13070 (N_13070,N_11534,N_11584);
or U13071 (N_13071,N_12279,N_11118);
nor U13072 (N_13072,N_11251,N_10147);
nand U13073 (N_13073,N_10267,N_11333);
nor U13074 (N_13074,N_10459,N_12076);
and U13075 (N_13075,N_11350,N_11099);
and U13076 (N_13076,N_11598,N_12208);
nor U13077 (N_13077,N_12468,N_12215);
nand U13078 (N_13078,N_12282,N_12401);
nand U13079 (N_13079,N_12143,N_12455);
or U13080 (N_13080,N_12037,N_11364);
nor U13081 (N_13081,N_12379,N_11593);
or U13082 (N_13082,N_10480,N_10084);
or U13083 (N_13083,N_10629,N_11656);
and U13084 (N_13084,N_12299,N_10615);
or U13085 (N_13085,N_10831,N_11016);
nand U13086 (N_13086,N_10639,N_10397);
nor U13087 (N_13087,N_10169,N_11544);
xnor U13088 (N_13088,N_11708,N_10852);
and U13089 (N_13089,N_10871,N_11824);
or U13090 (N_13090,N_11919,N_10454);
nand U13091 (N_13091,N_12422,N_10724);
xnor U13092 (N_13092,N_10207,N_11775);
and U13093 (N_13093,N_10557,N_10417);
or U13094 (N_13094,N_10661,N_10182);
or U13095 (N_13095,N_11475,N_10294);
and U13096 (N_13096,N_10029,N_11821);
and U13097 (N_13097,N_11319,N_10548);
and U13098 (N_13098,N_11224,N_10856);
nand U13099 (N_13099,N_10957,N_11439);
nand U13100 (N_13100,N_11998,N_10673);
or U13101 (N_13101,N_10984,N_12408);
or U13102 (N_13102,N_10473,N_12298);
nand U13103 (N_13103,N_11055,N_11922);
and U13104 (N_13104,N_10797,N_10184);
nor U13105 (N_13105,N_10130,N_10343);
xor U13106 (N_13106,N_10244,N_10506);
and U13107 (N_13107,N_10428,N_11039);
and U13108 (N_13108,N_10632,N_12181);
or U13109 (N_13109,N_11893,N_11172);
nor U13110 (N_13110,N_11471,N_10461);
or U13111 (N_13111,N_10401,N_11685);
nor U13112 (N_13112,N_12106,N_12470);
and U13113 (N_13113,N_10920,N_10448);
xnor U13114 (N_13114,N_11344,N_12175);
or U13115 (N_13115,N_11389,N_10921);
and U13116 (N_13116,N_12417,N_12168);
or U13117 (N_13117,N_12289,N_10043);
xor U13118 (N_13118,N_10882,N_12327);
nand U13119 (N_13119,N_10414,N_10924);
nor U13120 (N_13120,N_10907,N_10756);
and U13121 (N_13121,N_11053,N_10040);
and U13122 (N_13122,N_12281,N_11184);
or U13123 (N_13123,N_10602,N_10896);
xnor U13124 (N_13124,N_12070,N_10725);
nor U13125 (N_13125,N_11046,N_11104);
nand U13126 (N_13126,N_11092,N_10577);
nand U13127 (N_13127,N_10513,N_12253);
or U13128 (N_13128,N_11910,N_11835);
nand U13129 (N_13129,N_11551,N_10172);
and U13130 (N_13130,N_11707,N_11717);
nor U13131 (N_13131,N_12049,N_11638);
nand U13132 (N_13132,N_11855,N_10161);
and U13133 (N_13133,N_10341,N_10464);
nand U13134 (N_13134,N_10362,N_10091);
nand U13135 (N_13135,N_10310,N_12483);
nand U13136 (N_13136,N_10966,N_11545);
nor U13137 (N_13137,N_10555,N_11337);
or U13138 (N_13138,N_11869,N_11057);
and U13139 (N_13139,N_10385,N_10399);
nand U13140 (N_13140,N_10443,N_11536);
and U13141 (N_13141,N_10468,N_10307);
or U13142 (N_13142,N_10166,N_10405);
nor U13143 (N_13143,N_10117,N_12323);
or U13144 (N_13144,N_11479,N_12428);
or U13145 (N_13145,N_12169,N_10444);
nor U13146 (N_13146,N_10220,N_10775);
nand U13147 (N_13147,N_10648,N_11826);
xor U13148 (N_13148,N_11428,N_10360);
xnor U13149 (N_13149,N_11280,N_10738);
nor U13150 (N_13150,N_11829,N_11210);
nand U13151 (N_13151,N_11454,N_10056);
and U13152 (N_13152,N_10804,N_12438);
nand U13153 (N_13153,N_11315,N_12357);
nor U13154 (N_13154,N_12403,N_11642);
nand U13155 (N_13155,N_10902,N_11075);
or U13156 (N_13156,N_11710,N_11298);
or U13157 (N_13157,N_10005,N_10748);
and U13158 (N_13158,N_10931,N_10008);
nand U13159 (N_13159,N_10073,N_11081);
nand U13160 (N_13160,N_11102,N_10954);
or U13161 (N_13161,N_11076,N_12014);
or U13162 (N_13162,N_10916,N_11880);
xnor U13163 (N_13163,N_10470,N_10418);
nor U13164 (N_13164,N_11180,N_10888);
nand U13165 (N_13165,N_10517,N_10578);
and U13166 (N_13166,N_11751,N_12312);
or U13167 (N_13167,N_10897,N_11754);
nor U13168 (N_13168,N_10325,N_11214);
nand U13169 (N_13169,N_11484,N_11760);
nor U13170 (N_13170,N_11547,N_11687);
nor U13171 (N_13171,N_11374,N_12147);
and U13172 (N_13172,N_11447,N_10010);
nand U13173 (N_13173,N_11032,N_10683);
or U13174 (N_13174,N_10482,N_12021);
and U13175 (N_13175,N_10814,N_12124);
nor U13176 (N_13176,N_10320,N_10978);
or U13177 (N_13177,N_12061,N_12402);
or U13178 (N_13178,N_11167,N_11229);
nand U13179 (N_13179,N_11430,N_11512);
nand U13180 (N_13180,N_11345,N_10365);
nor U13181 (N_13181,N_11273,N_12191);
nor U13182 (N_13182,N_11971,N_11189);
nor U13183 (N_13183,N_11663,N_12300);
nor U13184 (N_13184,N_10195,N_10612);
nand U13185 (N_13185,N_11253,N_10074);
or U13186 (N_13186,N_11816,N_11533);
and U13187 (N_13187,N_11223,N_11235);
nand U13188 (N_13188,N_11202,N_10229);
nand U13189 (N_13189,N_11277,N_10382);
and U13190 (N_13190,N_11488,N_11410);
and U13191 (N_13191,N_12218,N_12161);
nor U13192 (N_13192,N_10332,N_12231);
nand U13193 (N_13193,N_10559,N_12426);
nor U13194 (N_13194,N_10810,N_12441);
or U13195 (N_13195,N_10148,N_11853);
nor U13196 (N_13196,N_12415,N_12326);
or U13197 (N_13197,N_11365,N_11678);
xor U13198 (N_13198,N_11309,N_12170);
nor U13199 (N_13199,N_10049,N_11886);
nand U13200 (N_13200,N_10675,N_10596);
nand U13201 (N_13201,N_12171,N_10635);
xor U13202 (N_13202,N_11296,N_12053);
nor U13203 (N_13203,N_11591,N_12113);
or U13204 (N_13204,N_12347,N_10733);
nor U13205 (N_13205,N_12109,N_10803);
nor U13206 (N_13206,N_10098,N_11770);
and U13207 (N_13207,N_10620,N_10833);
or U13208 (N_13208,N_11101,N_11779);
nor U13209 (N_13209,N_11230,N_12324);
or U13210 (N_13210,N_11480,N_11914);
nand U13211 (N_13211,N_10650,N_10268);
or U13212 (N_13212,N_11246,N_10667);
nand U13213 (N_13213,N_11261,N_11178);
and U13214 (N_13214,N_10563,N_11718);
or U13215 (N_13215,N_11452,N_11792);
and U13216 (N_13216,N_11504,N_12439);
nand U13217 (N_13217,N_12256,N_10421);
and U13218 (N_13218,N_11170,N_10811);
and U13219 (N_13219,N_11802,N_12374);
nor U13220 (N_13220,N_11141,N_10323);
or U13221 (N_13221,N_11614,N_12195);
nand U13222 (N_13222,N_11630,N_11036);
or U13223 (N_13223,N_10855,N_12112);
and U13224 (N_13224,N_11164,N_10236);
nor U13225 (N_13225,N_11528,N_10995);
and U13226 (N_13226,N_10384,N_10170);
nor U13227 (N_13227,N_12153,N_11155);
nor U13228 (N_13228,N_11951,N_11724);
xnor U13229 (N_13229,N_11145,N_10998);
and U13230 (N_13230,N_11986,N_11469);
nand U13231 (N_13231,N_11109,N_10127);
or U13232 (N_13232,N_11080,N_11787);
or U13233 (N_13233,N_10150,N_11492);
nand U13234 (N_13234,N_11011,N_10722);
nand U13235 (N_13235,N_10637,N_10525);
xor U13236 (N_13236,N_11288,N_12212);
and U13237 (N_13237,N_11866,N_11827);
and U13238 (N_13238,N_10009,N_12136);
or U13239 (N_13239,N_10510,N_10731);
nand U13240 (N_13240,N_11360,N_10044);
nor U13241 (N_13241,N_11634,N_11503);
nand U13242 (N_13242,N_10837,N_10022);
nor U13243 (N_13243,N_12062,N_10895);
or U13244 (N_13244,N_11451,N_11507);
and U13245 (N_13245,N_11499,N_11698);
nand U13246 (N_13246,N_10530,N_11446);
nand U13247 (N_13247,N_11970,N_12131);
nor U13248 (N_13248,N_10887,N_10183);
nand U13249 (N_13249,N_12386,N_11010);
or U13250 (N_13250,N_10309,N_11481);
nand U13251 (N_13251,N_11940,N_12317);
or U13252 (N_13252,N_10973,N_11564);
xnor U13253 (N_13253,N_10458,N_11252);
nor U13254 (N_13254,N_11607,N_11626);
xnor U13255 (N_13255,N_11948,N_12228);
and U13256 (N_13256,N_11455,N_11756);
nand U13257 (N_13257,N_10345,N_10614);
nor U13258 (N_13258,N_11789,N_10058);
and U13259 (N_13259,N_11762,N_10018);
nand U13260 (N_13260,N_11726,N_10188);
and U13261 (N_13261,N_11735,N_10770);
nor U13262 (N_13262,N_11888,N_10679);
nor U13263 (N_13263,N_10860,N_12499);
nand U13264 (N_13264,N_12117,N_10715);
and U13265 (N_13265,N_10894,N_12273);
and U13266 (N_13266,N_11793,N_11131);
nand U13267 (N_13267,N_12337,N_11161);
xor U13268 (N_13268,N_11159,N_10876);
or U13269 (N_13269,N_10286,N_10338);
nand U13270 (N_13270,N_10616,N_10390);
nand U13271 (N_13271,N_10877,N_10766);
nand U13272 (N_13272,N_10785,N_10192);
and U13273 (N_13273,N_10206,N_12096);
or U13274 (N_13274,N_12258,N_11133);
nor U13275 (N_13275,N_12011,N_11989);
or U13276 (N_13276,N_12265,N_11648);
and U13277 (N_13277,N_11286,N_11030);
nand U13278 (N_13278,N_10237,N_12111);
and U13279 (N_13279,N_10240,N_10760);
and U13280 (N_13280,N_11362,N_12227);
nand U13281 (N_13281,N_10749,N_10233);
or U13282 (N_13282,N_11313,N_11690);
and U13283 (N_13283,N_12203,N_11918);
nand U13284 (N_13284,N_11558,N_11486);
and U13285 (N_13285,N_11091,N_12437);
or U13286 (N_13286,N_12190,N_11640);
and U13287 (N_13287,N_11291,N_12194);
nand U13288 (N_13288,N_11819,N_11628);
nor U13289 (N_13289,N_10254,N_10442);
or U13290 (N_13290,N_11233,N_12025);
xnor U13291 (N_13291,N_11935,N_11864);
nand U13292 (N_13292,N_10311,N_10624);
nor U13293 (N_13293,N_10651,N_11884);
nor U13294 (N_13294,N_10795,N_10969);
xor U13295 (N_13295,N_10663,N_11952);
nand U13296 (N_13296,N_12105,N_11220);
nor U13297 (N_13297,N_10072,N_12479);
nand U13298 (N_13298,N_10848,N_11725);
and U13299 (N_13299,N_12311,N_11657);
nand U13300 (N_13300,N_10713,N_11898);
nor U13301 (N_13301,N_11125,N_10425);
nor U13302 (N_13302,N_10069,N_12491);
nand U13303 (N_13303,N_10526,N_10696);
nand U13304 (N_13304,N_11828,N_10567);
nor U13305 (N_13305,N_11568,N_10020);
and U13306 (N_13306,N_11929,N_12434);
nand U13307 (N_13307,N_10446,N_11883);
nand U13308 (N_13308,N_10440,N_11896);
nor U13309 (N_13309,N_10435,N_12003);
nor U13310 (N_13310,N_12207,N_10830);
nand U13311 (N_13311,N_10685,N_11435);
nor U13312 (N_13312,N_10611,N_11850);
nor U13313 (N_13313,N_12223,N_10878);
nor U13314 (N_13314,N_11409,N_10495);
nor U13315 (N_13315,N_10543,N_11783);
and U13316 (N_13316,N_11973,N_12290);
xnor U13317 (N_13317,N_10199,N_10380);
and U13318 (N_13318,N_11967,N_10337);
nor U13319 (N_13319,N_12475,N_11743);
and U13320 (N_13320,N_10528,N_10565);
nor U13321 (N_13321,N_11587,N_11742);
or U13322 (N_13322,N_11035,N_11699);
and U13323 (N_13323,N_10051,N_11082);
nand U13324 (N_13324,N_11248,N_11115);
nand U13325 (N_13325,N_11366,N_11411);
and U13326 (N_13326,N_10432,N_11837);
nor U13327 (N_13327,N_10832,N_11813);
or U13328 (N_13328,N_11782,N_11786);
nor U13329 (N_13329,N_11416,N_12339);
or U13330 (N_13330,N_11457,N_10168);
nor U13331 (N_13331,N_10216,N_10872);
or U13332 (N_13332,N_11578,N_11153);
nand U13333 (N_13333,N_10993,N_11572);
and U13334 (N_13334,N_12486,N_11721);
nor U13335 (N_13335,N_10113,N_10782);
and U13336 (N_13336,N_11408,N_12236);
nor U13337 (N_13337,N_10948,N_10662);
or U13338 (N_13338,N_12419,N_10494);
or U13339 (N_13339,N_12278,N_12353);
and U13340 (N_13340,N_12370,N_11644);
or U13341 (N_13341,N_11872,N_12373);
nor U13342 (N_13342,N_12077,N_11239);
or U13343 (N_13343,N_10579,N_10841);
nand U13344 (N_13344,N_12345,N_11928);
and U13345 (N_13345,N_12303,N_11863);
xor U13346 (N_13346,N_11143,N_12104);
and U13347 (N_13347,N_10356,N_12057);
and U13348 (N_13348,N_11570,N_12230);
xnor U13349 (N_13349,N_10527,N_10680);
nand U13350 (N_13350,N_10306,N_11310);
nand U13351 (N_13351,N_11312,N_10710);
nand U13352 (N_13352,N_12206,N_12065);
xnor U13353 (N_13353,N_11245,N_11063);
or U13354 (N_13354,N_10107,N_11716);
nand U13355 (N_13355,N_10767,N_11182);
nand U13356 (N_13356,N_10430,N_11390);
or U13357 (N_13357,N_11138,N_12068);
or U13358 (N_13358,N_10846,N_11183);
nor U13359 (N_13359,N_11692,N_12242);
and U13360 (N_13360,N_10851,N_11712);
xnor U13361 (N_13361,N_10420,N_11127);
xnor U13362 (N_13362,N_11684,N_10989);
or U13363 (N_13363,N_11352,N_11885);
nand U13364 (N_13364,N_10672,N_12142);
and U13365 (N_13365,N_10308,N_11574);
xnor U13366 (N_13366,N_12188,N_10853);
or U13367 (N_13367,N_11166,N_10551);
or U13368 (N_13368,N_10289,N_10465);
nor U13369 (N_13369,N_11925,N_12485);
nand U13370 (N_13370,N_10808,N_11221);
nand U13371 (N_13371,N_12030,N_10103);
and U13372 (N_13372,N_11487,N_10965);
xor U13373 (N_13373,N_10693,N_10189);
xor U13374 (N_13374,N_11962,N_11719);
and U13375 (N_13375,N_12071,N_10441);
nand U13376 (N_13376,N_11557,N_11976);
nand U13377 (N_13377,N_10110,N_12120);
and U13378 (N_13378,N_10128,N_10992);
nor U13379 (N_13379,N_11265,N_10253);
or U13380 (N_13380,N_11740,N_11773);
nor U13381 (N_13381,N_12172,N_10512);
xnor U13382 (N_13382,N_10238,N_10052);
or U13383 (N_13383,N_12451,N_10321);
and U13384 (N_13384,N_11377,N_10104);
xor U13385 (N_13385,N_10531,N_12287);
nand U13386 (N_13386,N_11722,N_10561);
nand U13387 (N_13387,N_10880,N_10133);
nor U13388 (N_13388,N_11119,N_12097);
or U13389 (N_13389,N_11794,N_10904);
or U13390 (N_13390,N_11957,N_10034);
nor U13391 (N_13391,N_11931,N_11619);
nor U13392 (N_13392,N_10716,N_11727);
nand U13393 (N_13393,N_12259,N_12272);
xor U13394 (N_13394,N_11336,N_11538);
xnor U13395 (N_13395,N_10035,N_11129);
nor U13396 (N_13396,N_10652,N_11107);
nor U13397 (N_13397,N_10717,N_10122);
and U13398 (N_13398,N_11745,N_11012);
nor U13399 (N_13399,N_10518,N_10372);
nor U13400 (N_13400,N_11815,N_10137);
nand U13401 (N_13401,N_10445,N_11795);
and U13402 (N_13402,N_10357,N_11259);
or U13403 (N_13403,N_12423,N_12178);
and U13404 (N_13404,N_10203,N_11691);
and U13405 (N_13405,N_10953,N_10386);
and U13406 (N_13406,N_12376,N_11897);
and U13407 (N_13407,N_10404,N_11329);
or U13408 (N_13408,N_11418,N_11380);
nor U13409 (N_13409,N_11270,N_10264);
or U13410 (N_13410,N_10118,N_10818);
nor U13411 (N_13411,N_10331,N_11049);
and U13412 (N_13412,N_11123,N_11168);
nand U13413 (N_13413,N_11974,N_10340);
nor U13414 (N_13414,N_12130,N_11269);
nand U13415 (N_13415,N_12421,N_11930);
and U13416 (N_13416,N_11739,N_12151);
and U13417 (N_13417,N_11594,N_10095);
or U13418 (N_13418,N_10939,N_11877);
and U13419 (N_13419,N_10415,N_11130);
nand U13420 (N_13420,N_11394,N_10336);
xnor U13421 (N_13421,N_10469,N_12064);
and U13422 (N_13422,N_10123,N_10828);
nor U13423 (N_13423,N_11847,N_10031);
nor U13424 (N_13424,N_11174,N_11376);
nand U13425 (N_13425,N_11176,N_11009);
and U13426 (N_13426,N_10436,N_11327);
or U13427 (N_13427,N_12089,N_12393);
nor U13428 (N_13428,N_10462,N_12197);
nor U13429 (N_13429,N_11086,N_11207);
and U13430 (N_13430,N_12472,N_12024);
nand U13431 (N_13431,N_10317,N_11601);
nand U13432 (N_13432,N_11669,N_11356);
xor U13433 (N_13433,N_12221,N_10677);
nor U13434 (N_13434,N_11524,N_11382);
and U13435 (N_13435,N_11434,N_11461);
and U13436 (N_13436,N_12033,N_10541);
and U13437 (N_13437,N_10046,N_10701);
xnor U13438 (N_13438,N_11234,N_12484);
and U13439 (N_13439,N_10587,N_10845);
nor U13440 (N_13440,N_11334,N_11979);
nand U13441 (N_13441,N_12126,N_10353);
or U13442 (N_13442,N_10951,N_10941);
nor U13443 (N_13443,N_11498,N_10085);
and U13444 (N_13444,N_10045,N_12356);
and U13445 (N_13445,N_10825,N_12348);
or U13446 (N_13446,N_11874,N_12286);
and U13447 (N_13447,N_10927,N_11483);
or U13448 (N_13448,N_11453,N_12493);
and U13449 (N_13449,N_12080,N_11240);
nor U13450 (N_13450,N_12392,N_10027);
or U13451 (N_13451,N_10581,N_10554);
or U13452 (N_13452,N_11646,N_11383);
nand U13453 (N_13453,N_10241,N_12377);
and U13454 (N_13454,N_10699,N_10690);
nor U13455 (N_13455,N_11670,N_10230);
nand U13456 (N_13456,N_10270,N_10259);
nor U13457 (N_13457,N_11623,N_11255);
nor U13458 (N_13458,N_10790,N_11843);
nor U13459 (N_13459,N_12214,N_10500);
or U13460 (N_13460,N_11889,N_11811);
nand U13461 (N_13461,N_11290,N_11367);
and U13462 (N_13462,N_12082,N_12412);
and U13463 (N_13463,N_11303,N_12367);
xnor U13464 (N_13464,N_12184,N_10387);
nand U13465 (N_13465,N_10802,N_11173);
nand U13466 (N_13466,N_10187,N_11450);
and U13467 (N_13467,N_11266,N_10239);
and U13468 (N_13468,N_10041,N_12173);
and U13469 (N_13469,N_10529,N_11565);
nor U13470 (N_13470,N_10660,N_10735);
nand U13471 (N_13471,N_11693,N_12490);
nor U13472 (N_13472,N_11939,N_10745);
nor U13473 (N_13473,N_10585,N_11470);
nand U13474 (N_13474,N_10919,N_11460);
nand U13475 (N_13475,N_11128,N_10576);
xor U13476 (N_13476,N_10918,N_11463);
nor U13477 (N_13477,N_11282,N_12084);
xnor U13478 (N_13478,N_11349,N_12411);
and U13479 (N_13479,N_10952,N_11953);
nor U13480 (N_13480,N_11386,N_12360);
and U13481 (N_13481,N_11441,N_11506);
and U13482 (N_13482,N_11963,N_10664);
and U13483 (N_13483,N_11242,N_10138);
or U13484 (N_13484,N_10114,N_10007);
nor U13485 (N_13485,N_12157,N_11093);
xor U13486 (N_13486,N_11045,N_10739);
nor U13487 (N_13487,N_11267,N_11293);
nor U13488 (N_13488,N_10088,N_11372);
nand U13489 (N_13489,N_11755,N_10944);
nor U13490 (N_13490,N_11066,N_10348);
or U13491 (N_13491,N_11741,N_11231);
and U13492 (N_13492,N_10149,N_10047);
and U13493 (N_13493,N_11772,N_11339);
nand U13494 (N_13494,N_12123,N_10747);
nand U13495 (N_13495,N_10591,N_10844);
or U13496 (N_13496,N_10140,N_10917);
nor U13497 (N_13497,N_10911,N_10424);
xnor U13498 (N_13498,N_10862,N_10553);
nor U13499 (N_13499,N_10866,N_12446);
nand U13500 (N_13500,N_11652,N_12460);
nor U13501 (N_13501,N_12187,N_12489);
nor U13502 (N_13502,N_11701,N_10584);
or U13503 (N_13503,N_12115,N_11750);
nand U13504 (N_13504,N_11388,N_10805);
xor U13505 (N_13505,N_11415,N_10037);
or U13506 (N_13506,N_11520,N_11502);
and U13507 (N_13507,N_12269,N_12487);
xor U13508 (N_13508,N_10740,N_12237);
xor U13509 (N_13509,N_11992,N_12385);
xor U13510 (N_13510,N_11404,N_11103);
nand U13511 (N_13511,N_12295,N_11069);
and U13512 (N_13512,N_10197,N_10014);
and U13513 (N_13513,N_12432,N_11895);
or U13514 (N_13514,N_11823,N_10859);
and U13515 (N_13515,N_10055,N_10250);
or U13516 (N_13516,N_10143,N_10928);
or U13517 (N_13517,N_12210,N_12496);
xor U13518 (N_13518,N_11694,N_11556);
and U13519 (N_13519,N_11596,N_10193);
nand U13520 (N_13520,N_10408,N_11433);
and U13521 (N_13521,N_10718,N_10002);
or U13522 (N_13522,N_11833,N_11673);
and U13523 (N_13523,N_10171,N_10908);
or U13524 (N_13524,N_10158,N_10545);
nor U13525 (N_13525,N_11445,N_11912);
and U13526 (N_13526,N_12322,N_11637);
nand U13527 (N_13527,N_11803,N_11530);
and U13528 (N_13528,N_11519,N_10036);
or U13529 (N_13529,N_11429,N_10608);
nand U13530 (N_13530,N_12355,N_10822);
and U13531 (N_13531,N_11028,N_10534);
nand U13532 (N_13532,N_10274,N_11643);
nand U13533 (N_13533,N_12338,N_11842);
xnor U13534 (N_13534,N_10881,N_12341);
nor U13535 (N_13535,N_10297,N_10726);
nand U13536 (N_13536,N_10395,N_11805);
nor U13537 (N_13537,N_10644,N_11343);
or U13538 (N_13538,N_12004,N_11160);
nor U13539 (N_13539,N_12055,N_12102);
nor U13540 (N_13540,N_10071,N_12388);
or U13541 (N_13541,N_11995,N_10406);
nor U13542 (N_13542,N_10363,N_10389);
xor U13543 (N_13543,N_11096,N_12209);
and U13544 (N_13544,N_10568,N_11274);
nand U13545 (N_13545,N_12459,N_11736);
nand U13546 (N_13546,N_10457,N_12310);
nand U13547 (N_13547,N_12052,N_10604);
nor U13548 (N_13548,N_11576,N_10720);
nand U13549 (N_13549,N_11907,N_12132);
or U13550 (N_13550,N_11532,N_10523);
and U13551 (N_13551,N_11671,N_11613);
xor U13552 (N_13552,N_10670,N_11196);
or U13553 (N_13553,N_11960,N_11121);
xnor U13554 (N_13554,N_10021,N_12350);
nand U13555 (N_13555,N_10945,N_12108);
or U13556 (N_13556,N_11554,N_11969);
and U13557 (N_13557,N_10682,N_10705);
or U13558 (N_13558,N_11899,N_12400);
or U13559 (N_13559,N_10381,N_11212);
and U13560 (N_13560,N_10946,N_11079);
or U13561 (N_13561,N_11983,N_12390);
or U13562 (N_13562,N_12384,N_10809);
and U13563 (N_13563,N_10793,N_10549);
nand U13564 (N_13564,N_11264,N_11432);
nor U13565 (N_13565,N_10485,N_11330);
nand U13566 (N_13566,N_12334,N_10155);
nand U13567 (N_13567,N_10603,N_12017);
nor U13568 (N_13568,N_11965,N_11529);
and U13569 (N_13569,N_10398,N_10394);
nand U13570 (N_13570,N_12257,N_11485);
nand U13571 (N_13571,N_10121,N_11954);
and U13572 (N_13572,N_10990,N_11209);
nand U13573 (N_13573,N_11511,N_11615);
and U13574 (N_13574,N_12110,N_10786);
nor U13575 (N_13575,N_12246,N_11041);
nor U13576 (N_13576,N_12083,N_11354);
and U13577 (N_13577,N_11262,N_11321);
and U13578 (N_13578,N_10829,N_12005);
and U13579 (N_13579,N_11747,N_11297);
and U13580 (N_13580,N_12183,N_12122);
or U13581 (N_13581,N_10070,N_11353);
or U13582 (N_13582,N_10489,N_10618);
or U13583 (N_13583,N_11169,N_11752);
nor U13584 (N_13584,N_11250,N_11087);
nor U13585 (N_13585,N_12404,N_10038);
and U13586 (N_13586,N_10109,N_10869);
or U13587 (N_13587,N_11126,N_10312);
nand U13588 (N_13588,N_11985,N_11851);
nor U13589 (N_13589,N_12008,N_11064);
and U13590 (N_13590,N_10006,N_10295);
nor U13591 (N_13591,N_10075,N_12075);
or U13592 (N_13592,N_12141,N_10923);
and U13593 (N_13593,N_10621,N_11675);
nor U13594 (N_13594,N_11403,N_10891);
nor U13595 (N_13595,N_10499,N_10231);
or U13596 (N_13596,N_10566,N_12333);
nor U13597 (N_13597,N_10275,N_11464);
and U13598 (N_13598,N_12155,N_11859);
nor U13599 (N_13599,N_10396,N_11426);
nand U13600 (N_13600,N_10915,N_11950);
nor U13601 (N_13601,N_10727,N_10177);
or U13602 (N_13602,N_10497,N_10284);
xor U13603 (N_13603,N_11001,N_11014);
nor U13604 (N_13604,N_11459,N_10141);
xnor U13605 (N_13605,N_10093,N_11375);
or U13606 (N_13606,N_10202,N_11287);
and U13607 (N_13607,N_11272,N_11746);
and U13608 (N_13608,N_11521,N_10700);
nand U13609 (N_13609,N_12448,N_11553);
and U13610 (N_13610,N_12330,N_11215);
or U13611 (N_13611,N_11825,N_10368);
or U13612 (N_13612,N_11586,N_12012);
and U13613 (N_13613,N_10134,N_10942);
and U13614 (N_13614,N_11038,N_10582);
xnor U13615 (N_13615,N_11156,N_10619);
xor U13616 (N_13616,N_12032,N_12450);
and U13617 (N_13617,N_12285,N_11500);
or U13618 (N_13618,N_11108,N_12158);
or U13619 (N_13619,N_10779,N_10467);
and U13620 (N_13620,N_10066,N_10471);
nor U13621 (N_13621,N_10676,N_11860);
nor U13622 (N_13622,N_10503,N_12177);
nor U13623 (N_13623,N_10062,N_12424);
nand U13624 (N_13624,N_11612,N_10413);
xor U13625 (N_13625,N_11807,N_12189);
nor U13626 (N_13626,N_10164,N_11518);
and U13627 (N_13627,N_11785,N_12444);
nor U13628 (N_13628,N_10101,N_11818);
xor U13629 (N_13629,N_11548,N_10416);
and U13630 (N_13630,N_10106,N_11181);
nand U13631 (N_13631,N_11784,N_12034);
nor U13632 (N_13632,N_10630,N_12308);
xnor U13633 (N_13633,N_12413,N_11580);
nand U13634 (N_13634,N_11781,N_11007);
and U13635 (N_13635,N_12294,N_12135);
xor U13636 (N_13636,N_10813,N_10280);
and U13637 (N_13637,N_10502,N_12098);
nand U13638 (N_13638,N_11720,N_11681);
nor U13639 (N_13639,N_10403,N_12414);
or U13640 (N_13640,N_10364,N_10447);
or U13641 (N_13641,N_10243,N_10956);
and U13642 (N_13642,N_10456,N_12349);
and U13643 (N_13643,N_11832,N_10769);
xor U13644 (N_13644,N_12268,N_11065);
or U13645 (N_13645,N_12405,N_10736);
or U13646 (N_13646,N_11219,N_11491);
and U13647 (N_13647,N_10460,N_10645);
and U13648 (N_13648,N_10025,N_10132);
xor U13649 (N_13649,N_10542,N_10850);
nand U13650 (N_13650,N_11514,N_12100);
nor U13651 (N_13651,N_11021,N_11332);
nand U13652 (N_13652,N_11331,N_10211);
xnor U13653 (N_13653,N_11878,N_11089);
or U13654 (N_13654,N_11602,N_10378);
nand U13655 (N_13655,N_10997,N_11444);
xor U13656 (N_13656,N_12044,N_10892);
nand U13657 (N_13657,N_11622,N_11672);
or U13658 (N_13658,N_10092,N_11186);
nor U13659 (N_13659,N_10659,N_12364);
and U13660 (N_13660,N_11705,N_12429);
or U13661 (N_13661,N_11496,N_10076);
or U13662 (N_13662,N_11632,N_11018);
xor U13663 (N_13663,N_11314,N_11379);
or U13664 (N_13664,N_11767,N_10367);
or U13665 (N_13665,N_10256,N_12461);
nand U13666 (N_13666,N_11022,N_12372);
nor U13667 (N_13667,N_10753,N_11769);
nand U13668 (N_13668,N_11142,N_10120);
and U13669 (N_13669,N_10925,N_12358);
and U13670 (N_13670,N_12462,N_10732);
nand U13671 (N_13671,N_11778,N_12047);
or U13672 (N_13672,N_10053,N_11852);
or U13673 (N_13673,N_11243,N_11522);
or U13674 (N_13674,N_12093,N_10151);
nor U13675 (N_13675,N_11921,N_12121);
or U13676 (N_13676,N_11090,N_11744);
nor U13677 (N_13677,N_12196,N_10600);
or U13678 (N_13678,N_10886,N_11361);
xnor U13679 (N_13679,N_10674,N_11873);
nand U13680 (N_13680,N_12248,N_11777);
nand U13681 (N_13681,N_10980,N_10981);
xor U13682 (N_13682,N_10375,N_11050);
and U13683 (N_13683,N_12420,N_12336);
and U13684 (N_13684,N_10213,N_11857);
nand U13685 (N_13685,N_12297,N_10922);
or U13686 (N_13686,N_10102,N_11203);
nand U13687 (N_13687,N_12381,N_11302);
nor U13688 (N_13688,N_12146,N_10801);
or U13689 (N_13689,N_10613,N_10156);
nand U13690 (N_13690,N_11140,N_11048);
and U13691 (N_13691,N_11071,N_12252);
nor U13692 (N_13692,N_10452,N_11427);
or U13693 (N_13693,N_11581,N_11569);
and U13694 (N_13694,N_11338,N_11482);
nand U13695 (N_13695,N_12200,N_11359);
or U13696 (N_13696,N_11213,N_10305);
or U13697 (N_13697,N_11776,N_12427);
nor U13698 (N_13698,N_10569,N_12264);
and U13699 (N_13699,N_12351,N_11975);
and U13700 (N_13700,N_10498,N_11704);
nand U13701 (N_13701,N_10959,N_11566);
or U13702 (N_13702,N_11000,N_10273);
nand U13703 (N_13703,N_10597,N_10042);
nand U13704 (N_13704,N_12018,N_11567);
and U13705 (N_13705,N_11552,N_10691);
nand U13706 (N_13706,N_10175,N_11384);
or U13707 (N_13707,N_10451,N_11477);
and U13708 (N_13708,N_10695,N_10292);
nor U13709 (N_13709,N_12219,N_12304);
or U13710 (N_13710,N_11241,N_10781);
and U13711 (N_13711,N_11854,N_11043);
nor U13712 (N_13712,N_10251,N_10126);
and U13713 (N_13713,N_10290,N_10838);
nor U13714 (N_13714,N_12291,N_10768);
or U13715 (N_13715,N_11800,N_12480);
or U13716 (N_13716,N_10068,N_11268);
nand U13717 (N_13717,N_11723,N_12027);
or U13718 (N_13718,N_11527,N_10655);
or U13719 (N_13719,N_11448,N_10024);
and U13720 (N_13720,N_11517,N_10974);
xor U13721 (N_13721,N_11400,N_11494);
nor U13722 (N_13722,N_10794,N_10124);
nor U13723 (N_13723,N_12028,N_10144);
nor U13724 (N_13724,N_11620,N_11655);
and U13725 (N_13725,N_11200,N_11944);
or U13726 (N_13726,N_10048,N_10901);
or U13727 (N_13727,N_11054,N_11387);
or U13728 (N_13728,N_12031,N_11304);
and U13729 (N_13729,N_10449,N_12241);
nand U13730 (N_13730,N_11501,N_11112);
or U13731 (N_13731,N_10709,N_11132);
and U13732 (N_13732,N_11616,N_11660);
nor U13733 (N_13733,N_10787,N_11095);
nand U13734 (N_13734,N_11163,N_10840);
and U13735 (N_13735,N_10514,N_10173);
nor U13736 (N_13736,N_10316,N_11462);
or U13737 (N_13737,N_10666,N_12094);
and U13738 (N_13738,N_11865,N_10028);
nor U13739 (N_13739,N_10285,N_11148);
nand U13740 (N_13740,N_12375,N_10179);
and U13741 (N_13741,N_11875,N_11397);
nand U13742 (N_13742,N_11876,N_11808);
nand U13743 (N_13743,N_10205,N_12086);
nor U13744 (N_13744,N_10857,N_11814);
nor U13745 (N_13745,N_10450,N_10669);
and U13746 (N_13746,N_12009,N_11438);
nor U13747 (N_13747,N_12198,N_10879);
and U13748 (N_13748,N_11421,N_10865);
xor U13749 (N_13749,N_11870,N_11355);
and U13750 (N_13750,N_11464,N_11083);
and U13751 (N_13751,N_11955,N_10588);
and U13752 (N_13752,N_12408,N_10301);
or U13753 (N_13753,N_12115,N_11338);
nand U13754 (N_13754,N_10137,N_10062);
or U13755 (N_13755,N_11650,N_12095);
nand U13756 (N_13756,N_11199,N_12028);
or U13757 (N_13757,N_12143,N_10505);
nor U13758 (N_13758,N_11317,N_10783);
nand U13759 (N_13759,N_10139,N_11004);
nand U13760 (N_13760,N_10102,N_12148);
and U13761 (N_13761,N_11847,N_11981);
xnor U13762 (N_13762,N_10700,N_10671);
or U13763 (N_13763,N_11052,N_12336);
and U13764 (N_13764,N_10456,N_10923);
and U13765 (N_13765,N_11410,N_10342);
nand U13766 (N_13766,N_12109,N_10424);
and U13767 (N_13767,N_12212,N_10893);
nor U13768 (N_13768,N_12399,N_12077);
nor U13769 (N_13769,N_10805,N_12481);
nor U13770 (N_13770,N_11074,N_10779);
or U13771 (N_13771,N_12202,N_12217);
xor U13772 (N_13772,N_10718,N_12171);
xnor U13773 (N_13773,N_10216,N_10750);
or U13774 (N_13774,N_10977,N_11304);
nor U13775 (N_13775,N_11146,N_12057);
and U13776 (N_13776,N_11499,N_11299);
and U13777 (N_13777,N_10321,N_11702);
or U13778 (N_13778,N_10441,N_12301);
and U13779 (N_13779,N_10032,N_10667);
xnor U13780 (N_13780,N_10388,N_10119);
nand U13781 (N_13781,N_11871,N_10689);
nand U13782 (N_13782,N_11085,N_12094);
nand U13783 (N_13783,N_10658,N_10554);
or U13784 (N_13784,N_10131,N_11802);
or U13785 (N_13785,N_11535,N_10130);
nand U13786 (N_13786,N_11672,N_11089);
nand U13787 (N_13787,N_10825,N_11701);
and U13788 (N_13788,N_10191,N_10173);
nand U13789 (N_13789,N_11241,N_11912);
xor U13790 (N_13790,N_12335,N_11709);
nor U13791 (N_13791,N_11206,N_11612);
nor U13792 (N_13792,N_11137,N_11295);
or U13793 (N_13793,N_12322,N_12002);
or U13794 (N_13794,N_10673,N_12376);
nor U13795 (N_13795,N_11478,N_12265);
xnor U13796 (N_13796,N_11869,N_10155);
nand U13797 (N_13797,N_10437,N_10347);
and U13798 (N_13798,N_11171,N_12258);
and U13799 (N_13799,N_11768,N_11388);
nor U13800 (N_13800,N_12415,N_10338);
nand U13801 (N_13801,N_11509,N_11380);
and U13802 (N_13802,N_10637,N_12183);
nor U13803 (N_13803,N_11984,N_12490);
nor U13804 (N_13804,N_11257,N_12335);
nor U13805 (N_13805,N_10237,N_11888);
nor U13806 (N_13806,N_11861,N_10610);
and U13807 (N_13807,N_12384,N_11208);
nor U13808 (N_13808,N_12165,N_10243);
nor U13809 (N_13809,N_10970,N_11200);
nand U13810 (N_13810,N_10363,N_10400);
or U13811 (N_13811,N_10846,N_10440);
nand U13812 (N_13812,N_12070,N_11011);
and U13813 (N_13813,N_11213,N_10866);
xnor U13814 (N_13814,N_10212,N_11207);
and U13815 (N_13815,N_11864,N_12238);
nand U13816 (N_13816,N_11753,N_11571);
nor U13817 (N_13817,N_11847,N_10856);
nand U13818 (N_13818,N_10564,N_12180);
or U13819 (N_13819,N_11812,N_12038);
nor U13820 (N_13820,N_11853,N_10077);
and U13821 (N_13821,N_10969,N_12295);
xor U13822 (N_13822,N_10713,N_12091);
and U13823 (N_13823,N_12157,N_10391);
and U13824 (N_13824,N_10518,N_10989);
and U13825 (N_13825,N_10931,N_10511);
nor U13826 (N_13826,N_10038,N_11658);
or U13827 (N_13827,N_11063,N_10771);
or U13828 (N_13828,N_12353,N_12132);
nor U13829 (N_13829,N_11725,N_12419);
xnor U13830 (N_13830,N_11778,N_10117);
or U13831 (N_13831,N_10908,N_11679);
and U13832 (N_13832,N_10711,N_12462);
or U13833 (N_13833,N_10223,N_10210);
and U13834 (N_13834,N_10110,N_12113);
nor U13835 (N_13835,N_11009,N_11706);
xor U13836 (N_13836,N_12039,N_11977);
nand U13837 (N_13837,N_11663,N_11079);
or U13838 (N_13838,N_11464,N_11435);
nor U13839 (N_13839,N_10337,N_12092);
and U13840 (N_13840,N_12486,N_10856);
or U13841 (N_13841,N_11836,N_10140);
nor U13842 (N_13842,N_11759,N_11101);
or U13843 (N_13843,N_10782,N_10667);
nand U13844 (N_13844,N_12352,N_12460);
or U13845 (N_13845,N_10060,N_11834);
and U13846 (N_13846,N_10134,N_11950);
nor U13847 (N_13847,N_10691,N_10445);
or U13848 (N_13848,N_10865,N_11021);
or U13849 (N_13849,N_12157,N_11751);
or U13850 (N_13850,N_10367,N_12328);
nand U13851 (N_13851,N_10419,N_10509);
and U13852 (N_13852,N_11826,N_10095);
and U13853 (N_13853,N_10523,N_10883);
nand U13854 (N_13854,N_12093,N_10582);
nor U13855 (N_13855,N_12049,N_11883);
xnor U13856 (N_13856,N_10327,N_10278);
nor U13857 (N_13857,N_10468,N_10506);
xnor U13858 (N_13858,N_10287,N_11131);
and U13859 (N_13859,N_10812,N_11349);
or U13860 (N_13860,N_11088,N_10864);
nor U13861 (N_13861,N_11173,N_10659);
nor U13862 (N_13862,N_10518,N_11920);
nor U13863 (N_13863,N_11131,N_11191);
and U13864 (N_13864,N_10394,N_11419);
and U13865 (N_13865,N_10488,N_12230);
nand U13866 (N_13866,N_11552,N_12417);
and U13867 (N_13867,N_11092,N_11108);
nand U13868 (N_13868,N_12162,N_12351);
nand U13869 (N_13869,N_11717,N_10978);
or U13870 (N_13870,N_10613,N_12410);
nor U13871 (N_13871,N_11190,N_10127);
or U13872 (N_13872,N_10207,N_11742);
xnor U13873 (N_13873,N_10406,N_11869);
and U13874 (N_13874,N_10435,N_11368);
nand U13875 (N_13875,N_11720,N_10739);
nor U13876 (N_13876,N_10380,N_11602);
and U13877 (N_13877,N_10536,N_11413);
nand U13878 (N_13878,N_10727,N_12424);
nor U13879 (N_13879,N_12352,N_10932);
nand U13880 (N_13880,N_12482,N_11167);
and U13881 (N_13881,N_10409,N_10211);
nand U13882 (N_13882,N_11154,N_10255);
xnor U13883 (N_13883,N_11053,N_11008);
or U13884 (N_13884,N_11366,N_12328);
and U13885 (N_13885,N_11423,N_10101);
nor U13886 (N_13886,N_10940,N_11337);
xnor U13887 (N_13887,N_10364,N_10428);
nor U13888 (N_13888,N_12411,N_10338);
nand U13889 (N_13889,N_10668,N_11540);
nand U13890 (N_13890,N_10148,N_12071);
and U13891 (N_13891,N_12039,N_11750);
nor U13892 (N_13892,N_12228,N_11387);
xnor U13893 (N_13893,N_10325,N_10558);
or U13894 (N_13894,N_11169,N_12318);
or U13895 (N_13895,N_11970,N_10717);
and U13896 (N_13896,N_12085,N_12254);
nor U13897 (N_13897,N_11300,N_11792);
and U13898 (N_13898,N_12227,N_11755);
nand U13899 (N_13899,N_11442,N_11610);
and U13900 (N_13900,N_11054,N_12145);
and U13901 (N_13901,N_12456,N_10686);
and U13902 (N_13902,N_12094,N_10930);
nand U13903 (N_13903,N_12115,N_11847);
and U13904 (N_13904,N_12350,N_12235);
nand U13905 (N_13905,N_11529,N_10433);
nand U13906 (N_13906,N_11708,N_11939);
nand U13907 (N_13907,N_10122,N_11973);
nor U13908 (N_13908,N_11831,N_11577);
and U13909 (N_13909,N_12117,N_10598);
nor U13910 (N_13910,N_10675,N_10003);
nor U13911 (N_13911,N_10035,N_12139);
and U13912 (N_13912,N_12025,N_11831);
nand U13913 (N_13913,N_12437,N_10360);
or U13914 (N_13914,N_10271,N_11924);
and U13915 (N_13915,N_12275,N_11181);
xor U13916 (N_13916,N_10508,N_12324);
xor U13917 (N_13917,N_11579,N_10527);
nor U13918 (N_13918,N_12037,N_11935);
or U13919 (N_13919,N_12108,N_10090);
nand U13920 (N_13920,N_10246,N_12344);
and U13921 (N_13921,N_11688,N_11182);
or U13922 (N_13922,N_11897,N_12226);
and U13923 (N_13923,N_11357,N_12460);
nor U13924 (N_13924,N_12365,N_10409);
and U13925 (N_13925,N_11599,N_11542);
and U13926 (N_13926,N_10039,N_11883);
nand U13927 (N_13927,N_11907,N_10067);
or U13928 (N_13928,N_11671,N_10358);
nor U13929 (N_13929,N_11419,N_12342);
nor U13930 (N_13930,N_11918,N_10273);
or U13931 (N_13931,N_10017,N_12113);
nor U13932 (N_13932,N_11982,N_12421);
nand U13933 (N_13933,N_10102,N_11213);
nor U13934 (N_13934,N_12330,N_11772);
or U13935 (N_13935,N_12173,N_10177);
or U13936 (N_13936,N_11161,N_10447);
and U13937 (N_13937,N_11980,N_11020);
nand U13938 (N_13938,N_12082,N_11309);
nand U13939 (N_13939,N_11453,N_11614);
nor U13940 (N_13940,N_11026,N_11793);
and U13941 (N_13941,N_12460,N_12107);
and U13942 (N_13942,N_11928,N_10176);
or U13943 (N_13943,N_10126,N_12128);
and U13944 (N_13944,N_10787,N_10676);
nor U13945 (N_13945,N_12183,N_11066);
and U13946 (N_13946,N_10740,N_11767);
nor U13947 (N_13947,N_12079,N_10453);
nor U13948 (N_13948,N_10784,N_12257);
nor U13949 (N_13949,N_12359,N_11967);
or U13950 (N_13950,N_11565,N_11966);
nor U13951 (N_13951,N_12466,N_10873);
nor U13952 (N_13952,N_11271,N_10264);
and U13953 (N_13953,N_12253,N_10022);
and U13954 (N_13954,N_11807,N_11773);
or U13955 (N_13955,N_11241,N_11737);
or U13956 (N_13956,N_10775,N_12440);
or U13957 (N_13957,N_10918,N_10105);
or U13958 (N_13958,N_12005,N_11707);
nor U13959 (N_13959,N_11341,N_11112);
and U13960 (N_13960,N_10156,N_11726);
and U13961 (N_13961,N_10424,N_10141);
nor U13962 (N_13962,N_11093,N_10855);
nor U13963 (N_13963,N_12280,N_10001);
or U13964 (N_13964,N_10179,N_10487);
and U13965 (N_13965,N_10551,N_10178);
and U13966 (N_13966,N_11305,N_12393);
and U13967 (N_13967,N_10770,N_10669);
xnor U13968 (N_13968,N_10419,N_11390);
nand U13969 (N_13969,N_10219,N_10286);
and U13970 (N_13970,N_11663,N_12127);
or U13971 (N_13971,N_12403,N_11040);
nand U13972 (N_13972,N_11179,N_11810);
or U13973 (N_13973,N_12241,N_12052);
or U13974 (N_13974,N_10325,N_10999);
and U13975 (N_13975,N_11716,N_10355);
or U13976 (N_13976,N_10849,N_10909);
or U13977 (N_13977,N_10433,N_11996);
nand U13978 (N_13978,N_10562,N_11997);
and U13979 (N_13979,N_11841,N_11571);
and U13980 (N_13980,N_10177,N_11238);
nor U13981 (N_13981,N_10145,N_12469);
and U13982 (N_13982,N_10991,N_10813);
or U13983 (N_13983,N_10322,N_10347);
nand U13984 (N_13984,N_11262,N_10236);
xor U13985 (N_13985,N_11357,N_10501);
and U13986 (N_13986,N_12010,N_11070);
and U13987 (N_13987,N_10589,N_10381);
and U13988 (N_13988,N_10443,N_11825);
nand U13989 (N_13989,N_10425,N_10204);
nand U13990 (N_13990,N_11187,N_11992);
and U13991 (N_13991,N_10104,N_10060);
nand U13992 (N_13992,N_10770,N_11209);
nor U13993 (N_13993,N_12494,N_11967);
and U13994 (N_13994,N_11097,N_11972);
nand U13995 (N_13995,N_11114,N_10123);
and U13996 (N_13996,N_12378,N_11507);
or U13997 (N_13997,N_11257,N_10196);
nand U13998 (N_13998,N_11101,N_10983);
nand U13999 (N_13999,N_11343,N_10019);
and U14000 (N_14000,N_12143,N_11006);
nor U14001 (N_14001,N_11301,N_11765);
nor U14002 (N_14002,N_11523,N_10228);
nand U14003 (N_14003,N_11107,N_11593);
or U14004 (N_14004,N_11912,N_10821);
nand U14005 (N_14005,N_11624,N_10895);
nor U14006 (N_14006,N_11550,N_10949);
or U14007 (N_14007,N_11839,N_10907);
and U14008 (N_14008,N_10040,N_10703);
or U14009 (N_14009,N_12204,N_10309);
xor U14010 (N_14010,N_11463,N_11419);
and U14011 (N_14011,N_11662,N_12287);
xnor U14012 (N_14012,N_11752,N_10408);
and U14013 (N_14013,N_11878,N_10330);
nor U14014 (N_14014,N_12133,N_10612);
nand U14015 (N_14015,N_12057,N_10106);
nand U14016 (N_14016,N_11348,N_11530);
nand U14017 (N_14017,N_10922,N_12158);
and U14018 (N_14018,N_11030,N_10610);
or U14019 (N_14019,N_10056,N_10711);
and U14020 (N_14020,N_10089,N_10947);
nor U14021 (N_14021,N_11826,N_10836);
nand U14022 (N_14022,N_12471,N_11376);
nand U14023 (N_14023,N_11824,N_11679);
and U14024 (N_14024,N_12333,N_10851);
and U14025 (N_14025,N_11919,N_12222);
or U14026 (N_14026,N_10073,N_10933);
and U14027 (N_14027,N_11124,N_10922);
nor U14028 (N_14028,N_10604,N_11148);
nand U14029 (N_14029,N_10001,N_10954);
nor U14030 (N_14030,N_10049,N_10956);
nand U14031 (N_14031,N_11734,N_10340);
or U14032 (N_14032,N_11130,N_10999);
nand U14033 (N_14033,N_12209,N_10820);
nand U14034 (N_14034,N_11823,N_10787);
nor U14035 (N_14035,N_10931,N_12409);
and U14036 (N_14036,N_12255,N_10199);
and U14037 (N_14037,N_11865,N_11055);
nor U14038 (N_14038,N_10084,N_10488);
and U14039 (N_14039,N_12001,N_12252);
nand U14040 (N_14040,N_10010,N_11876);
nor U14041 (N_14041,N_11881,N_10746);
nand U14042 (N_14042,N_10616,N_11531);
xor U14043 (N_14043,N_10790,N_11649);
or U14044 (N_14044,N_10299,N_10891);
or U14045 (N_14045,N_10111,N_10035);
nor U14046 (N_14046,N_11868,N_10585);
xor U14047 (N_14047,N_10884,N_12087);
nand U14048 (N_14048,N_10509,N_12361);
and U14049 (N_14049,N_11747,N_10230);
or U14050 (N_14050,N_10685,N_11086);
nor U14051 (N_14051,N_11642,N_10003);
or U14052 (N_14052,N_10044,N_11544);
or U14053 (N_14053,N_11634,N_11084);
nor U14054 (N_14054,N_11636,N_11788);
nand U14055 (N_14055,N_11411,N_10142);
nand U14056 (N_14056,N_11530,N_11242);
and U14057 (N_14057,N_10652,N_11411);
nand U14058 (N_14058,N_11797,N_12204);
nor U14059 (N_14059,N_10167,N_12423);
nand U14060 (N_14060,N_10742,N_11354);
and U14061 (N_14061,N_12349,N_11003);
nor U14062 (N_14062,N_11648,N_10923);
nand U14063 (N_14063,N_10154,N_12395);
nand U14064 (N_14064,N_10774,N_12151);
nand U14065 (N_14065,N_10164,N_10086);
and U14066 (N_14066,N_10952,N_11016);
xnor U14067 (N_14067,N_11019,N_11167);
nand U14068 (N_14068,N_12213,N_10390);
and U14069 (N_14069,N_11545,N_11038);
xnor U14070 (N_14070,N_10691,N_11931);
nand U14071 (N_14071,N_12177,N_10518);
and U14072 (N_14072,N_11662,N_10955);
or U14073 (N_14073,N_11444,N_12027);
nand U14074 (N_14074,N_11039,N_11002);
and U14075 (N_14075,N_11706,N_10686);
nand U14076 (N_14076,N_10180,N_12324);
or U14077 (N_14077,N_10821,N_11326);
nand U14078 (N_14078,N_10014,N_11103);
or U14079 (N_14079,N_11796,N_12445);
nand U14080 (N_14080,N_11465,N_10281);
and U14081 (N_14081,N_11449,N_12156);
and U14082 (N_14082,N_10701,N_12008);
and U14083 (N_14083,N_12181,N_12190);
and U14084 (N_14084,N_11386,N_11621);
nand U14085 (N_14085,N_11239,N_10314);
nor U14086 (N_14086,N_11845,N_12375);
nor U14087 (N_14087,N_12338,N_10694);
or U14088 (N_14088,N_10823,N_11347);
nor U14089 (N_14089,N_10483,N_11655);
and U14090 (N_14090,N_10021,N_10772);
xnor U14091 (N_14091,N_11225,N_10576);
nand U14092 (N_14092,N_11261,N_11968);
nand U14093 (N_14093,N_10153,N_12378);
xor U14094 (N_14094,N_12187,N_11359);
nor U14095 (N_14095,N_10838,N_12304);
nor U14096 (N_14096,N_11925,N_10818);
nand U14097 (N_14097,N_10584,N_10444);
nand U14098 (N_14098,N_10126,N_10894);
nor U14099 (N_14099,N_10557,N_11945);
nor U14100 (N_14100,N_11302,N_10636);
or U14101 (N_14101,N_11122,N_10178);
and U14102 (N_14102,N_11734,N_11350);
xnor U14103 (N_14103,N_10259,N_12051);
xnor U14104 (N_14104,N_10780,N_11770);
nand U14105 (N_14105,N_11628,N_10311);
nand U14106 (N_14106,N_10119,N_11366);
nor U14107 (N_14107,N_10792,N_10777);
nor U14108 (N_14108,N_12332,N_10730);
and U14109 (N_14109,N_10972,N_10653);
nand U14110 (N_14110,N_11065,N_12402);
or U14111 (N_14111,N_10700,N_11546);
nor U14112 (N_14112,N_10242,N_12220);
nand U14113 (N_14113,N_10000,N_11699);
nand U14114 (N_14114,N_10453,N_11878);
xnor U14115 (N_14115,N_10666,N_10905);
nor U14116 (N_14116,N_11164,N_12276);
and U14117 (N_14117,N_10967,N_11996);
or U14118 (N_14118,N_10427,N_10203);
nor U14119 (N_14119,N_12475,N_11546);
nand U14120 (N_14120,N_12362,N_10218);
and U14121 (N_14121,N_12198,N_10089);
nor U14122 (N_14122,N_10309,N_10467);
nand U14123 (N_14123,N_11914,N_10418);
nor U14124 (N_14124,N_11198,N_12330);
xor U14125 (N_14125,N_11308,N_12293);
or U14126 (N_14126,N_11804,N_11334);
or U14127 (N_14127,N_10427,N_12160);
and U14128 (N_14128,N_11111,N_10539);
nand U14129 (N_14129,N_10483,N_12358);
and U14130 (N_14130,N_11517,N_11629);
and U14131 (N_14131,N_11205,N_11291);
nor U14132 (N_14132,N_11137,N_11150);
nor U14133 (N_14133,N_11810,N_12051);
and U14134 (N_14134,N_10612,N_10922);
nand U14135 (N_14135,N_12305,N_12445);
nor U14136 (N_14136,N_11508,N_10203);
nand U14137 (N_14137,N_11139,N_12418);
nor U14138 (N_14138,N_10534,N_10104);
nand U14139 (N_14139,N_11991,N_11385);
xnor U14140 (N_14140,N_10654,N_11898);
nand U14141 (N_14141,N_11064,N_11455);
nor U14142 (N_14142,N_12093,N_12206);
nor U14143 (N_14143,N_11562,N_10716);
nor U14144 (N_14144,N_10622,N_12084);
nand U14145 (N_14145,N_12330,N_11482);
nand U14146 (N_14146,N_10953,N_12250);
nor U14147 (N_14147,N_11715,N_10315);
nor U14148 (N_14148,N_11909,N_10223);
or U14149 (N_14149,N_10343,N_10121);
and U14150 (N_14150,N_12059,N_10552);
and U14151 (N_14151,N_12333,N_11342);
nand U14152 (N_14152,N_10695,N_11646);
nand U14153 (N_14153,N_12279,N_10214);
nor U14154 (N_14154,N_10766,N_12035);
and U14155 (N_14155,N_12179,N_11936);
nor U14156 (N_14156,N_10485,N_12034);
nor U14157 (N_14157,N_10782,N_11485);
nand U14158 (N_14158,N_11116,N_10058);
and U14159 (N_14159,N_11702,N_11359);
nand U14160 (N_14160,N_10703,N_11505);
nor U14161 (N_14161,N_12103,N_11424);
nor U14162 (N_14162,N_10605,N_10288);
and U14163 (N_14163,N_11977,N_10603);
nor U14164 (N_14164,N_11468,N_11215);
or U14165 (N_14165,N_10898,N_10142);
or U14166 (N_14166,N_10662,N_10375);
nand U14167 (N_14167,N_10024,N_11719);
nand U14168 (N_14168,N_11678,N_10927);
and U14169 (N_14169,N_11569,N_11729);
or U14170 (N_14170,N_10920,N_10856);
and U14171 (N_14171,N_12162,N_12150);
nor U14172 (N_14172,N_11626,N_10945);
nor U14173 (N_14173,N_11189,N_11835);
or U14174 (N_14174,N_11645,N_10908);
nand U14175 (N_14175,N_10493,N_10645);
nand U14176 (N_14176,N_12421,N_10796);
and U14177 (N_14177,N_12002,N_11016);
xnor U14178 (N_14178,N_11686,N_10918);
or U14179 (N_14179,N_10915,N_11206);
nor U14180 (N_14180,N_10424,N_11060);
nor U14181 (N_14181,N_10769,N_12208);
nor U14182 (N_14182,N_11325,N_10773);
xor U14183 (N_14183,N_11486,N_10323);
and U14184 (N_14184,N_11760,N_10192);
or U14185 (N_14185,N_11094,N_11800);
or U14186 (N_14186,N_11709,N_11612);
or U14187 (N_14187,N_11724,N_10495);
and U14188 (N_14188,N_11856,N_10950);
or U14189 (N_14189,N_10161,N_11854);
nand U14190 (N_14190,N_11351,N_10283);
and U14191 (N_14191,N_11338,N_11109);
nand U14192 (N_14192,N_10764,N_10221);
xnor U14193 (N_14193,N_10762,N_12052);
xnor U14194 (N_14194,N_10069,N_11919);
or U14195 (N_14195,N_10436,N_11478);
and U14196 (N_14196,N_10731,N_12471);
and U14197 (N_14197,N_11323,N_11992);
nand U14198 (N_14198,N_10701,N_12100);
nor U14199 (N_14199,N_12139,N_10817);
and U14200 (N_14200,N_11866,N_11103);
or U14201 (N_14201,N_12015,N_12268);
nand U14202 (N_14202,N_10649,N_12155);
nor U14203 (N_14203,N_11918,N_11010);
or U14204 (N_14204,N_11263,N_10268);
or U14205 (N_14205,N_12403,N_12360);
nor U14206 (N_14206,N_11603,N_12318);
xor U14207 (N_14207,N_11645,N_12235);
and U14208 (N_14208,N_11313,N_10145);
nor U14209 (N_14209,N_11231,N_11264);
and U14210 (N_14210,N_11681,N_11404);
or U14211 (N_14211,N_10181,N_10547);
or U14212 (N_14212,N_10399,N_10554);
or U14213 (N_14213,N_11959,N_10860);
nand U14214 (N_14214,N_10028,N_12051);
or U14215 (N_14215,N_11893,N_12172);
nand U14216 (N_14216,N_12186,N_11191);
nor U14217 (N_14217,N_10525,N_12108);
or U14218 (N_14218,N_12070,N_10330);
nand U14219 (N_14219,N_12153,N_11576);
or U14220 (N_14220,N_12067,N_11209);
nand U14221 (N_14221,N_10574,N_10864);
nor U14222 (N_14222,N_11734,N_11464);
and U14223 (N_14223,N_10497,N_10858);
and U14224 (N_14224,N_10024,N_10040);
xnor U14225 (N_14225,N_12400,N_12354);
and U14226 (N_14226,N_10388,N_10326);
or U14227 (N_14227,N_10758,N_12236);
or U14228 (N_14228,N_10493,N_12096);
nand U14229 (N_14229,N_11749,N_10098);
and U14230 (N_14230,N_10158,N_10783);
or U14231 (N_14231,N_12149,N_11028);
or U14232 (N_14232,N_12289,N_10433);
nor U14233 (N_14233,N_11218,N_10718);
nor U14234 (N_14234,N_12191,N_10027);
nand U14235 (N_14235,N_12136,N_10196);
nor U14236 (N_14236,N_10355,N_10164);
nor U14237 (N_14237,N_12362,N_11268);
or U14238 (N_14238,N_11059,N_12427);
nor U14239 (N_14239,N_12468,N_11731);
and U14240 (N_14240,N_10549,N_12351);
and U14241 (N_14241,N_11498,N_10525);
nor U14242 (N_14242,N_11150,N_11926);
nor U14243 (N_14243,N_10591,N_11675);
xor U14244 (N_14244,N_11267,N_12044);
and U14245 (N_14245,N_10738,N_10626);
or U14246 (N_14246,N_11701,N_10641);
nand U14247 (N_14247,N_12258,N_10040);
and U14248 (N_14248,N_11367,N_12494);
or U14249 (N_14249,N_11556,N_11330);
xor U14250 (N_14250,N_12390,N_10082);
nand U14251 (N_14251,N_11799,N_10784);
and U14252 (N_14252,N_10225,N_11454);
nand U14253 (N_14253,N_11782,N_12412);
and U14254 (N_14254,N_10681,N_11010);
or U14255 (N_14255,N_10370,N_11494);
nor U14256 (N_14256,N_11563,N_11996);
nor U14257 (N_14257,N_12137,N_11792);
nand U14258 (N_14258,N_12369,N_12145);
nand U14259 (N_14259,N_10922,N_12295);
or U14260 (N_14260,N_10329,N_10815);
or U14261 (N_14261,N_10606,N_11384);
or U14262 (N_14262,N_12338,N_11474);
nor U14263 (N_14263,N_10135,N_10133);
xor U14264 (N_14264,N_10808,N_11284);
xnor U14265 (N_14265,N_10669,N_10213);
or U14266 (N_14266,N_10730,N_10467);
nor U14267 (N_14267,N_10761,N_10694);
and U14268 (N_14268,N_10247,N_12373);
or U14269 (N_14269,N_10033,N_10718);
nor U14270 (N_14270,N_10396,N_11860);
xor U14271 (N_14271,N_11577,N_10866);
or U14272 (N_14272,N_10219,N_10220);
or U14273 (N_14273,N_11564,N_10593);
xor U14274 (N_14274,N_12328,N_10500);
nor U14275 (N_14275,N_12029,N_12106);
nand U14276 (N_14276,N_11345,N_12479);
nor U14277 (N_14277,N_10356,N_10153);
nand U14278 (N_14278,N_11789,N_11681);
xnor U14279 (N_14279,N_11512,N_10855);
nor U14280 (N_14280,N_10453,N_10690);
xnor U14281 (N_14281,N_10546,N_11691);
or U14282 (N_14282,N_11952,N_10570);
nand U14283 (N_14283,N_11638,N_10964);
nor U14284 (N_14284,N_10032,N_12292);
xor U14285 (N_14285,N_12404,N_11200);
nor U14286 (N_14286,N_11039,N_11036);
and U14287 (N_14287,N_11522,N_11817);
and U14288 (N_14288,N_10210,N_10372);
and U14289 (N_14289,N_11600,N_11203);
or U14290 (N_14290,N_10069,N_10591);
or U14291 (N_14291,N_10816,N_11546);
nand U14292 (N_14292,N_12152,N_12255);
and U14293 (N_14293,N_10659,N_10944);
nand U14294 (N_14294,N_11238,N_10196);
xor U14295 (N_14295,N_12440,N_12499);
and U14296 (N_14296,N_10583,N_11146);
nand U14297 (N_14297,N_10281,N_11855);
and U14298 (N_14298,N_12106,N_10508);
nor U14299 (N_14299,N_10860,N_10625);
nand U14300 (N_14300,N_11218,N_11955);
and U14301 (N_14301,N_10705,N_11815);
nor U14302 (N_14302,N_10644,N_10167);
and U14303 (N_14303,N_12055,N_11233);
nor U14304 (N_14304,N_10002,N_10544);
xnor U14305 (N_14305,N_11622,N_12441);
nand U14306 (N_14306,N_11044,N_10084);
or U14307 (N_14307,N_11111,N_10337);
xnor U14308 (N_14308,N_12436,N_12151);
nor U14309 (N_14309,N_10474,N_11313);
or U14310 (N_14310,N_10077,N_10143);
and U14311 (N_14311,N_12388,N_11767);
or U14312 (N_14312,N_11477,N_12492);
or U14313 (N_14313,N_10368,N_11050);
nand U14314 (N_14314,N_11539,N_11164);
and U14315 (N_14315,N_10498,N_11289);
xor U14316 (N_14316,N_10897,N_10205);
or U14317 (N_14317,N_12424,N_10375);
nand U14318 (N_14318,N_12124,N_12290);
nand U14319 (N_14319,N_10669,N_11981);
nand U14320 (N_14320,N_12234,N_11444);
nand U14321 (N_14321,N_10584,N_10690);
or U14322 (N_14322,N_12255,N_11037);
and U14323 (N_14323,N_11789,N_11147);
nand U14324 (N_14324,N_11068,N_11631);
or U14325 (N_14325,N_11026,N_10245);
and U14326 (N_14326,N_11328,N_10599);
and U14327 (N_14327,N_11757,N_11010);
and U14328 (N_14328,N_11030,N_11037);
nand U14329 (N_14329,N_10093,N_10845);
nor U14330 (N_14330,N_10057,N_12355);
nand U14331 (N_14331,N_12102,N_10604);
nand U14332 (N_14332,N_11227,N_10881);
xnor U14333 (N_14333,N_11349,N_10820);
and U14334 (N_14334,N_11429,N_12087);
and U14335 (N_14335,N_10181,N_12260);
and U14336 (N_14336,N_11556,N_12054);
nor U14337 (N_14337,N_12134,N_10247);
and U14338 (N_14338,N_10936,N_10538);
xnor U14339 (N_14339,N_12377,N_11829);
or U14340 (N_14340,N_10949,N_10540);
and U14341 (N_14341,N_10285,N_11482);
or U14342 (N_14342,N_11829,N_10879);
nor U14343 (N_14343,N_11915,N_12257);
or U14344 (N_14344,N_12269,N_10439);
and U14345 (N_14345,N_12239,N_10709);
xor U14346 (N_14346,N_10901,N_12353);
nor U14347 (N_14347,N_11822,N_10557);
and U14348 (N_14348,N_10290,N_12038);
and U14349 (N_14349,N_12371,N_11972);
nor U14350 (N_14350,N_11616,N_11180);
or U14351 (N_14351,N_10251,N_11493);
or U14352 (N_14352,N_11835,N_10003);
or U14353 (N_14353,N_11708,N_11308);
and U14354 (N_14354,N_10653,N_10730);
and U14355 (N_14355,N_10116,N_10724);
xnor U14356 (N_14356,N_11074,N_10237);
nor U14357 (N_14357,N_11856,N_11774);
nand U14358 (N_14358,N_12362,N_12359);
nor U14359 (N_14359,N_11562,N_10331);
nor U14360 (N_14360,N_10706,N_12286);
and U14361 (N_14361,N_11034,N_11947);
nand U14362 (N_14362,N_10635,N_10367);
nor U14363 (N_14363,N_12331,N_12287);
nor U14364 (N_14364,N_10814,N_11311);
or U14365 (N_14365,N_10065,N_12014);
nor U14366 (N_14366,N_12126,N_11702);
nand U14367 (N_14367,N_12368,N_12046);
nor U14368 (N_14368,N_11293,N_11555);
nor U14369 (N_14369,N_10643,N_11476);
nand U14370 (N_14370,N_10829,N_11748);
or U14371 (N_14371,N_10749,N_11102);
nand U14372 (N_14372,N_10611,N_11545);
or U14373 (N_14373,N_12280,N_10092);
and U14374 (N_14374,N_11440,N_10209);
and U14375 (N_14375,N_11402,N_10208);
nor U14376 (N_14376,N_10666,N_11355);
nor U14377 (N_14377,N_10943,N_12060);
nand U14378 (N_14378,N_10301,N_10677);
or U14379 (N_14379,N_11773,N_10577);
or U14380 (N_14380,N_10311,N_10277);
nor U14381 (N_14381,N_11694,N_11587);
or U14382 (N_14382,N_11918,N_11296);
xor U14383 (N_14383,N_11468,N_11122);
or U14384 (N_14384,N_10056,N_11573);
nand U14385 (N_14385,N_11125,N_11368);
nor U14386 (N_14386,N_11291,N_11210);
or U14387 (N_14387,N_11784,N_10137);
and U14388 (N_14388,N_11713,N_11301);
nor U14389 (N_14389,N_11323,N_11079);
and U14390 (N_14390,N_11662,N_11064);
nor U14391 (N_14391,N_12366,N_10622);
nand U14392 (N_14392,N_10021,N_10662);
or U14393 (N_14393,N_10628,N_10594);
nand U14394 (N_14394,N_11019,N_10689);
and U14395 (N_14395,N_10224,N_11859);
or U14396 (N_14396,N_11473,N_10564);
xnor U14397 (N_14397,N_10025,N_11437);
or U14398 (N_14398,N_10794,N_10371);
nor U14399 (N_14399,N_10498,N_10810);
xnor U14400 (N_14400,N_10188,N_12382);
nand U14401 (N_14401,N_10039,N_10947);
nand U14402 (N_14402,N_12370,N_11041);
nor U14403 (N_14403,N_12409,N_12113);
nand U14404 (N_14404,N_12092,N_10621);
nand U14405 (N_14405,N_10567,N_12335);
nand U14406 (N_14406,N_11417,N_11135);
nand U14407 (N_14407,N_10016,N_11520);
or U14408 (N_14408,N_10143,N_11998);
nand U14409 (N_14409,N_11686,N_11523);
nand U14410 (N_14410,N_12271,N_11813);
nand U14411 (N_14411,N_10518,N_11396);
nor U14412 (N_14412,N_11275,N_10054);
or U14413 (N_14413,N_10002,N_10928);
xnor U14414 (N_14414,N_10653,N_10011);
and U14415 (N_14415,N_11436,N_12231);
nand U14416 (N_14416,N_11182,N_11919);
nand U14417 (N_14417,N_11305,N_10390);
or U14418 (N_14418,N_11733,N_11064);
nand U14419 (N_14419,N_11284,N_10956);
nor U14420 (N_14420,N_12200,N_10024);
xnor U14421 (N_14421,N_11801,N_10857);
nor U14422 (N_14422,N_10664,N_11416);
nor U14423 (N_14423,N_10346,N_11019);
nor U14424 (N_14424,N_10790,N_10980);
and U14425 (N_14425,N_12002,N_10000);
nor U14426 (N_14426,N_12362,N_10630);
nand U14427 (N_14427,N_10379,N_12037);
and U14428 (N_14428,N_10529,N_10582);
or U14429 (N_14429,N_10842,N_12158);
nor U14430 (N_14430,N_10636,N_11615);
or U14431 (N_14431,N_11775,N_12177);
nand U14432 (N_14432,N_10760,N_10192);
nand U14433 (N_14433,N_11988,N_10536);
or U14434 (N_14434,N_10417,N_12204);
or U14435 (N_14435,N_12363,N_12148);
or U14436 (N_14436,N_10957,N_11211);
or U14437 (N_14437,N_11854,N_10790);
nor U14438 (N_14438,N_10998,N_11461);
nor U14439 (N_14439,N_11294,N_11177);
nor U14440 (N_14440,N_12300,N_11289);
nor U14441 (N_14441,N_11510,N_10799);
nand U14442 (N_14442,N_12350,N_12388);
nand U14443 (N_14443,N_10735,N_11958);
nand U14444 (N_14444,N_12434,N_11236);
nand U14445 (N_14445,N_11281,N_11948);
xor U14446 (N_14446,N_11493,N_10490);
and U14447 (N_14447,N_11091,N_10990);
nor U14448 (N_14448,N_10965,N_12472);
xnor U14449 (N_14449,N_10925,N_12413);
nand U14450 (N_14450,N_10170,N_11866);
nand U14451 (N_14451,N_10137,N_10999);
nor U14452 (N_14452,N_11080,N_10376);
xnor U14453 (N_14453,N_11256,N_10524);
nand U14454 (N_14454,N_11096,N_10695);
or U14455 (N_14455,N_10181,N_10735);
or U14456 (N_14456,N_11044,N_11016);
and U14457 (N_14457,N_11706,N_12161);
xor U14458 (N_14458,N_10673,N_10262);
and U14459 (N_14459,N_10772,N_10247);
nand U14460 (N_14460,N_11909,N_10299);
and U14461 (N_14461,N_10959,N_10579);
nor U14462 (N_14462,N_11199,N_12085);
xor U14463 (N_14463,N_11362,N_11497);
nor U14464 (N_14464,N_12059,N_12435);
or U14465 (N_14465,N_10873,N_10140);
and U14466 (N_14466,N_12054,N_11009);
nor U14467 (N_14467,N_11423,N_10258);
and U14468 (N_14468,N_11313,N_11346);
or U14469 (N_14469,N_10566,N_11726);
xnor U14470 (N_14470,N_10437,N_10304);
and U14471 (N_14471,N_10641,N_10304);
xnor U14472 (N_14472,N_12422,N_11689);
or U14473 (N_14473,N_11092,N_10942);
xnor U14474 (N_14474,N_10158,N_12367);
xor U14475 (N_14475,N_10203,N_11704);
nand U14476 (N_14476,N_10138,N_10750);
xor U14477 (N_14477,N_10294,N_11187);
nor U14478 (N_14478,N_10534,N_11777);
or U14479 (N_14479,N_10620,N_10613);
and U14480 (N_14480,N_11258,N_10535);
or U14481 (N_14481,N_10310,N_10812);
nand U14482 (N_14482,N_11316,N_11965);
or U14483 (N_14483,N_10332,N_12055);
nand U14484 (N_14484,N_10489,N_11824);
nor U14485 (N_14485,N_12498,N_10632);
nand U14486 (N_14486,N_11133,N_10724);
nor U14487 (N_14487,N_11585,N_11317);
and U14488 (N_14488,N_11041,N_12204);
nand U14489 (N_14489,N_12315,N_10131);
nor U14490 (N_14490,N_12355,N_10792);
nand U14491 (N_14491,N_10484,N_12308);
nor U14492 (N_14492,N_11423,N_10438);
nand U14493 (N_14493,N_12162,N_10832);
or U14494 (N_14494,N_11964,N_10518);
or U14495 (N_14495,N_12074,N_10331);
nor U14496 (N_14496,N_12195,N_12395);
nor U14497 (N_14497,N_12234,N_10059);
xor U14498 (N_14498,N_11299,N_11689);
and U14499 (N_14499,N_10912,N_11306);
or U14500 (N_14500,N_11107,N_11873);
or U14501 (N_14501,N_11596,N_10601);
nor U14502 (N_14502,N_10969,N_10664);
and U14503 (N_14503,N_10604,N_11692);
nand U14504 (N_14504,N_10302,N_11796);
nor U14505 (N_14505,N_12398,N_10588);
nor U14506 (N_14506,N_10229,N_11808);
nor U14507 (N_14507,N_10603,N_11892);
nor U14508 (N_14508,N_10694,N_11958);
nor U14509 (N_14509,N_11244,N_12394);
nor U14510 (N_14510,N_10192,N_10079);
or U14511 (N_14511,N_10275,N_10571);
and U14512 (N_14512,N_11108,N_10669);
nor U14513 (N_14513,N_10215,N_10911);
or U14514 (N_14514,N_10294,N_10516);
nand U14515 (N_14515,N_11677,N_11296);
and U14516 (N_14516,N_11678,N_11658);
or U14517 (N_14517,N_10224,N_11085);
nor U14518 (N_14518,N_11334,N_10673);
or U14519 (N_14519,N_11878,N_12199);
and U14520 (N_14520,N_12470,N_11514);
nor U14521 (N_14521,N_10103,N_10577);
nor U14522 (N_14522,N_11782,N_11093);
and U14523 (N_14523,N_10692,N_12429);
xnor U14524 (N_14524,N_12397,N_10071);
nand U14525 (N_14525,N_10024,N_12162);
or U14526 (N_14526,N_10065,N_12363);
or U14527 (N_14527,N_10697,N_12001);
nor U14528 (N_14528,N_11101,N_11531);
or U14529 (N_14529,N_11825,N_12274);
nand U14530 (N_14530,N_10273,N_10490);
and U14531 (N_14531,N_11054,N_11733);
or U14532 (N_14532,N_10172,N_11786);
nor U14533 (N_14533,N_10646,N_11107);
nand U14534 (N_14534,N_12384,N_10467);
nand U14535 (N_14535,N_12163,N_11710);
nand U14536 (N_14536,N_11089,N_10800);
or U14537 (N_14537,N_11608,N_11379);
and U14538 (N_14538,N_10432,N_10749);
or U14539 (N_14539,N_11133,N_11837);
xnor U14540 (N_14540,N_10162,N_10698);
nor U14541 (N_14541,N_11480,N_12017);
and U14542 (N_14542,N_10669,N_11978);
nand U14543 (N_14543,N_10088,N_11407);
nor U14544 (N_14544,N_10987,N_12323);
nor U14545 (N_14545,N_11587,N_12310);
nor U14546 (N_14546,N_10193,N_11623);
nand U14547 (N_14547,N_12374,N_11974);
nor U14548 (N_14548,N_10499,N_11574);
xnor U14549 (N_14549,N_12448,N_11040);
nor U14550 (N_14550,N_11105,N_11666);
nor U14551 (N_14551,N_10947,N_11977);
nor U14552 (N_14552,N_11872,N_11504);
nand U14553 (N_14553,N_10057,N_11968);
and U14554 (N_14554,N_11180,N_12209);
nand U14555 (N_14555,N_12274,N_10747);
and U14556 (N_14556,N_10803,N_10816);
and U14557 (N_14557,N_12488,N_10096);
nor U14558 (N_14558,N_10196,N_11954);
nor U14559 (N_14559,N_10665,N_11382);
or U14560 (N_14560,N_12328,N_12417);
nand U14561 (N_14561,N_12090,N_12029);
nand U14562 (N_14562,N_11717,N_11496);
nor U14563 (N_14563,N_11193,N_10918);
and U14564 (N_14564,N_10172,N_11243);
nand U14565 (N_14565,N_10615,N_10771);
nor U14566 (N_14566,N_12186,N_10240);
nand U14567 (N_14567,N_10640,N_11098);
nand U14568 (N_14568,N_10526,N_12252);
nor U14569 (N_14569,N_10628,N_12111);
nand U14570 (N_14570,N_10989,N_10010);
or U14571 (N_14571,N_11715,N_11750);
and U14572 (N_14572,N_11853,N_11512);
or U14573 (N_14573,N_12025,N_12315);
or U14574 (N_14574,N_10434,N_11299);
and U14575 (N_14575,N_10372,N_11887);
or U14576 (N_14576,N_10610,N_10108);
nand U14577 (N_14577,N_10047,N_11875);
nand U14578 (N_14578,N_12148,N_12162);
or U14579 (N_14579,N_10322,N_11309);
and U14580 (N_14580,N_11557,N_10594);
nor U14581 (N_14581,N_12152,N_10527);
nor U14582 (N_14582,N_11328,N_11261);
or U14583 (N_14583,N_11561,N_12015);
nor U14584 (N_14584,N_12012,N_12455);
or U14585 (N_14585,N_10519,N_10617);
nand U14586 (N_14586,N_10464,N_11666);
nand U14587 (N_14587,N_12040,N_12224);
nand U14588 (N_14588,N_11207,N_11771);
xnor U14589 (N_14589,N_12066,N_10705);
nand U14590 (N_14590,N_10283,N_12201);
or U14591 (N_14591,N_12254,N_11938);
and U14592 (N_14592,N_10037,N_10931);
or U14593 (N_14593,N_11359,N_10156);
nand U14594 (N_14594,N_10471,N_10147);
nand U14595 (N_14595,N_10356,N_10098);
nand U14596 (N_14596,N_12393,N_10001);
nor U14597 (N_14597,N_10572,N_11321);
or U14598 (N_14598,N_10268,N_10879);
nor U14599 (N_14599,N_10174,N_11506);
or U14600 (N_14600,N_11366,N_10639);
or U14601 (N_14601,N_11309,N_11514);
or U14602 (N_14602,N_12404,N_11397);
or U14603 (N_14603,N_12070,N_11335);
xor U14604 (N_14604,N_10173,N_10361);
or U14605 (N_14605,N_11085,N_12423);
xor U14606 (N_14606,N_11151,N_10129);
or U14607 (N_14607,N_11960,N_10545);
xor U14608 (N_14608,N_10458,N_11367);
or U14609 (N_14609,N_10058,N_10692);
nand U14610 (N_14610,N_10300,N_10059);
or U14611 (N_14611,N_10126,N_10910);
nand U14612 (N_14612,N_11623,N_11663);
xor U14613 (N_14613,N_10992,N_10312);
nand U14614 (N_14614,N_11877,N_10542);
nand U14615 (N_14615,N_10337,N_10479);
nor U14616 (N_14616,N_11629,N_11485);
and U14617 (N_14617,N_10042,N_10950);
nand U14618 (N_14618,N_10555,N_11371);
nor U14619 (N_14619,N_11840,N_10488);
nand U14620 (N_14620,N_10759,N_11512);
or U14621 (N_14621,N_11251,N_11805);
and U14622 (N_14622,N_11051,N_11789);
and U14623 (N_14623,N_12387,N_10097);
xnor U14624 (N_14624,N_11926,N_11853);
nor U14625 (N_14625,N_10516,N_11417);
nand U14626 (N_14626,N_10331,N_12215);
nand U14627 (N_14627,N_10823,N_11285);
nor U14628 (N_14628,N_12457,N_11117);
nor U14629 (N_14629,N_10514,N_11178);
nor U14630 (N_14630,N_12072,N_11036);
xnor U14631 (N_14631,N_10477,N_11796);
nand U14632 (N_14632,N_10088,N_11996);
nand U14633 (N_14633,N_11394,N_11781);
nand U14634 (N_14634,N_10777,N_11160);
and U14635 (N_14635,N_10823,N_12349);
nor U14636 (N_14636,N_10976,N_11344);
nor U14637 (N_14637,N_12399,N_11559);
and U14638 (N_14638,N_11918,N_10167);
or U14639 (N_14639,N_12193,N_10781);
or U14640 (N_14640,N_10476,N_10551);
or U14641 (N_14641,N_10362,N_10626);
nand U14642 (N_14642,N_11917,N_12258);
nor U14643 (N_14643,N_10964,N_10758);
or U14644 (N_14644,N_12065,N_11898);
or U14645 (N_14645,N_12298,N_10659);
or U14646 (N_14646,N_10431,N_10048);
xor U14647 (N_14647,N_11639,N_10510);
and U14648 (N_14648,N_11211,N_10302);
or U14649 (N_14649,N_11208,N_12486);
or U14650 (N_14650,N_11114,N_10739);
nand U14651 (N_14651,N_11053,N_10940);
nor U14652 (N_14652,N_10990,N_10305);
or U14653 (N_14653,N_10493,N_11467);
nor U14654 (N_14654,N_11568,N_10842);
nor U14655 (N_14655,N_11911,N_11353);
or U14656 (N_14656,N_11576,N_12308);
or U14657 (N_14657,N_10707,N_10927);
nor U14658 (N_14658,N_10082,N_10800);
or U14659 (N_14659,N_11519,N_10440);
and U14660 (N_14660,N_11517,N_11512);
nor U14661 (N_14661,N_11750,N_12329);
nand U14662 (N_14662,N_10847,N_12334);
and U14663 (N_14663,N_10546,N_11278);
and U14664 (N_14664,N_10983,N_11228);
or U14665 (N_14665,N_11178,N_11235);
and U14666 (N_14666,N_11957,N_11040);
nor U14667 (N_14667,N_11512,N_10388);
or U14668 (N_14668,N_11150,N_11281);
nand U14669 (N_14669,N_11559,N_12446);
nand U14670 (N_14670,N_12373,N_10079);
nor U14671 (N_14671,N_10233,N_12202);
and U14672 (N_14672,N_11892,N_12499);
and U14673 (N_14673,N_10803,N_11356);
and U14674 (N_14674,N_11237,N_11201);
nand U14675 (N_14675,N_10890,N_11488);
or U14676 (N_14676,N_11562,N_10091);
xnor U14677 (N_14677,N_10165,N_10211);
and U14678 (N_14678,N_11195,N_12258);
nand U14679 (N_14679,N_11591,N_10139);
xor U14680 (N_14680,N_10572,N_12296);
nor U14681 (N_14681,N_10159,N_11774);
nand U14682 (N_14682,N_12323,N_10243);
or U14683 (N_14683,N_10533,N_12083);
xnor U14684 (N_14684,N_10573,N_11283);
nor U14685 (N_14685,N_12111,N_11391);
and U14686 (N_14686,N_10041,N_11990);
nor U14687 (N_14687,N_10914,N_11364);
nor U14688 (N_14688,N_11540,N_12097);
nand U14689 (N_14689,N_11868,N_10851);
nand U14690 (N_14690,N_11984,N_12307);
or U14691 (N_14691,N_12457,N_12410);
nand U14692 (N_14692,N_10022,N_11965);
nor U14693 (N_14693,N_12009,N_11343);
nor U14694 (N_14694,N_12409,N_10242);
or U14695 (N_14695,N_11184,N_12363);
or U14696 (N_14696,N_12232,N_10908);
and U14697 (N_14697,N_11269,N_10025);
xor U14698 (N_14698,N_10137,N_11365);
nor U14699 (N_14699,N_11886,N_11176);
and U14700 (N_14700,N_10175,N_11811);
or U14701 (N_14701,N_11199,N_11373);
or U14702 (N_14702,N_12063,N_11977);
nor U14703 (N_14703,N_11647,N_11222);
nor U14704 (N_14704,N_11605,N_10565);
nand U14705 (N_14705,N_10840,N_11232);
xnor U14706 (N_14706,N_11914,N_10549);
or U14707 (N_14707,N_11242,N_11298);
nand U14708 (N_14708,N_12416,N_10475);
nand U14709 (N_14709,N_10029,N_11830);
or U14710 (N_14710,N_12274,N_11520);
nand U14711 (N_14711,N_11001,N_10637);
nor U14712 (N_14712,N_10789,N_11884);
or U14713 (N_14713,N_11722,N_11946);
nor U14714 (N_14714,N_11868,N_10742);
nor U14715 (N_14715,N_10510,N_10354);
nor U14716 (N_14716,N_10552,N_10256);
nand U14717 (N_14717,N_11443,N_11592);
or U14718 (N_14718,N_11818,N_11203);
nor U14719 (N_14719,N_11106,N_10670);
xnor U14720 (N_14720,N_11941,N_10805);
or U14721 (N_14721,N_11732,N_10243);
nor U14722 (N_14722,N_11860,N_11771);
nand U14723 (N_14723,N_12466,N_10832);
nand U14724 (N_14724,N_11464,N_11233);
nor U14725 (N_14725,N_11891,N_11134);
or U14726 (N_14726,N_11990,N_11214);
or U14727 (N_14727,N_12396,N_11469);
or U14728 (N_14728,N_11019,N_10024);
xor U14729 (N_14729,N_11566,N_10097);
or U14730 (N_14730,N_10518,N_11750);
and U14731 (N_14731,N_12426,N_10216);
nor U14732 (N_14732,N_11766,N_10105);
or U14733 (N_14733,N_11217,N_12342);
xor U14734 (N_14734,N_11799,N_10093);
or U14735 (N_14735,N_11653,N_12420);
nor U14736 (N_14736,N_10692,N_10859);
nor U14737 (N_14737,N_10604,N_11829);
nor U14738 (N_14738,N_11270,N_10775);
nor U14739 (N_14739,N_11710,N_11478);
xor U14740 (N_14740,N_11716,N_11467);
nor U14741 (N_14741,N_12324,N_12100);
or U14742 (N_14742,N_10401,N_10443);
nand U14743 (N_14743,N_11220,N_11803);
and U14744 (N_14744,N_10270,N_10172);
and U14745 (N_14745,N_10326,N_10344);
nor U14746 (N_14746,N_11380,N_12248);
and U14747 (N_14747,N_10527,N_11044);
nand U14748 (N_14748,N_10833,N_11448);
nand U14749 (N_14749,N_10239,N_10843);
or U14750 (N_14750,N_11740,N_10216);
xnor U14751 (N_14751,N_10330,N_11694);
and U14752 (N_14752,N_11767,N_10029);
or U14753 (N_14753,N_11720,N_10953);
nor U14754 (N_14754,N_12365,N_10070);
and U14755 (N_14755,N_12304,N_11284);
nor U14756 (N_14756,N_10875,N_12391);
and U14757 (N_14757,N_11346,N_11400);
or U14758 (N_14758,N_10638,N_10286);
or U14759 (N_14759,N_12132,N_10813);
nand U14760 (N_14760,N_10203,N_10754);
nand U14761 (N_14761,N_12137,N_10411);
nand U14762 (N_14762,N_11388,N_12017);
and U14763 (N_14763,N_11477,N_10782);
nor U14764 (N_14764,N_12406,N_10833);
and U14765 (N_14765,N_11239,N_11491);
and U14766 (N_14766,N_11993,N_12166);
and U14767 (N_14767,N_12455,N_12121);
and U14768 (N_14768,N_10491,N_12363);
and U14769 (N_14769,N_10321,N_10000);
nand U14770 (N_14770,N_11700,N_10281);
xnor U14771 (N_14771,N_11418,N_11960);
or U14772 (N_14772,N_11001,N_11381);
nor U14773 (N_14773,N_10382,N_11500);
or U14774 (N_14774,N_11168,N_11765);
nand U14775 (N_14775,N_10747,N_12287);
nand U14776 (N_14776,N_11956,N_12130);
or U14777 (N_14777,N_11091,N_10400);
or U14778 (N_14778,N_10700,N_11539);
and U14779 (N_14779,N_11886,N_10001);
and U14780 (N_14780,N_10020,N_11109);
nor U14781 (N_14781,N_12338,N_10880);
and U14782 (N_14782,N_11497,N_10079);
nand U14783 (N_14783,N_11994,N_10577);
nor U14784 (N_14784,N_11121,N_11156);
nor U14785 (N_14785,N_10004,N_12128);
and U14786 (N_14786,N_12167,N_11904);
xor U14787 (N_14787,N_10403,N_11161);
nor U14788 (N_14788,N_11122,N_11066);
or U14789 (N_14789,N_10167,N_11385);
xor U14790 (N_14790,N_11185,N_11909);
nand U14791 (N_14791,N_12496,N_12371);
nand U14792 (N_14792,N_10878,N_10373);
nor U14793 (N_14793,N_12308,N_12188);
nand U14794 (N_14794,N_12049,N_12225);
nand U14795 (N_14795,N_10559,N_10733);
nor U14796 (N_14796,N_10869,N_10385);
and U14797 (N_14797,N_11700,N_11526);
nand U14798 (N_14798,N_11945,N_11571);
nand U14799 (N_14799,N_12329,N_10750);
and U14800 (N_14800,N_10228,N_11461);
nor U14801 (N_14801,N_10467,N_11124);
or U14802 (N_14802,N_11067,N_10669);
nor U14803 (N_14803,N_11237,N_10702);
nand U14804 (N_14804,N_11101,N_12139);
nor U14805 (N_14805,N_11819,N_10973);
or U14806 (N_14806,N_11326,N_11778);
and U14807 (N_14807,N_11565,N_10560);
nor U14808 (N_14808,N_11524,N_10959);
nor U14809 (N_14809,N_10153,N_10353);
or U14810 (N_14810,N_10675,N_11479);
and U14811 (N_14811,N_11516,N_10480);
or U14812 (N_14812,N_12086,N_11641);
or U14813 (N_14813,N_11134,N_10414);
or U14814 (N_14814,N_10103,N_12421);
or U14815 (N_14815,N_11311,N_11842);
and U14816 (N_14816,N_11776,N_10215);
and U14817 (N_14817,N_11047,N_10191);
and U14818 (N_14818,N_12188,N_11370);
nand U14819 (N_14819,N_12145,N_10550);
nand U14820 (N_14820,N_10977,N_10998);
nand U14821 (N_14821,N_10058,N_11768);
or U14822 (N_14822,N_12242,N_10420);
xor U14823 (N_14823,N_10958,N_11410);
and U14824 (N_14824,N_11920,N_11581);
nor U14825 (N_14825,N_11739,N_11425);
or U14826 (N_14826,N_12452,N_11873);
nand U14827 (N_14827,N_11788,N_11537);
or U14828 (N_14828,N_10249,N_11713);
nor U14829 (N_14829,N_10861,N_11101);
and U14830 (N_14830,N_10313,N_10675);
nor U14831 (N_14831,N_10826,N_11629);
nor U14832 (N_14832,N_11251,N_11725);
and U14833 (N_14833,N_10044,N_10126);
nor U14834 (N_14834,N_10814,N_11013);
or U14835 (N_14835,N_10447,N_11431);
or U14836 (N_14836,N_11427,N_10857);
or U14837 (N_14837,N_10298,N_11633);
and U14838 (N_14838,N_10561,N_11924);
or U14839 (N_14839,N_12343,N_12361);
and U14840 (N_14840,N_11820,N_11524);
or U14841 (N_14841,N_10205,N_11566);
or U14842 (N_14842,N_10966,N_12045);
and U14843 (N_14843,N_11532,N_11603);
or U14844 (N_14844,N_11135,N_10464);
or U14845 (N_14845,N_11288,N_10118);
xnor U14846 (N_14846,N_11110,N_10576);
and U14847 (N_14847,N_12101,N_12082);
nand U14848 (N_14848,N_11789,N_11102);
or U14849 (N_14849,N_11894,N_10571);
nand U14850 (N_14850,N_12308,N_10200);
or U14851 (N_14851,N_10205,N_11733);
nor U14852 (N_14852,N_11031,N_11223);
and U14853 (N_14853,N_11296,N_11602);
nand U14854 (N_14854,N_12427,N_12283);
xor U14855 (N_14855,N_10369,N_11619);
or U14856 (N_14856,N_11102,N_11888);
or U14857 (N_14857,N_12170,N_12495);
or U14858 (N_14858,N_11485,N_10166);
and U14859 (N_14859,N_11953,N_10150);
xor U14860 (N_14860,N_12205,N_11372);
xnor U14861 (N_14861,N_11824,N_10621);
or U14862 (N_14862,N_11085,N_10673);
nor U14863 (N_14863,N_10195,N_10989);
xor U14864 (N_14864,N_10101,N_11033);
and U14865 (N_14865,N_11625,N_12035);
or U14866 (N_14866,N_10571,N_11435);
nor U14867 (N_14867,N_11941,N_10877);
nor U14868 (N_14868,N_10626,N_11859);
or U14869 (N_14869,N_12004,N_11284);
xnor U14870 (N_14870,N_11927,N_10750);
or U14871 (N_14871,N_11922,N_11042);
or U14872 (N_14872,N_10345,N_10413);
and U14873 (N_14873,N_10024,N_11614);
xnor U14874 (N_14874,N_11651,N_10624);
and U14875 (N_14875,N_10763,N_10786);
nand U14876 (N_14876,N_11583,N_11687);
nor U14877 (N_14877,N_12103,N_11664);
or U14878 (N_14878,N_12257,N_10008);
nor U14879 (N_14879,N_12144,N_10260);
nand U14880 (N_14880,N_11418,N_10075);
nand U14881 (N_14881,N_11152,N_10706);
or U14882 (N_14882,N_10250,N_11375);
nor U14883 (N_14883,N_11304,N_12390);
nand U14884 (N_14884,N_12100,N_11753);
nor U14885 (N_14885,N_10658,N_11356);
nand U14886 (N_14886,N_12217,N_11552);
or U14887 (N_14887,N_10555,N_12437);
and U14888 (N_14888,N_10927,N_11436);
and U14889 (N_14889,N_11177,N_11409);
nor U14890 (N_14890,N_11229,N_10338);
or U14891 (N_14891,N_11687,N_11689);
and U14892 (N_14892,N_11798,N_10774);
nor U14893 (N_14893,N_10394,N_10700);
nand U14894 (N_14894,N_12113,N_12003);
or U14895 (N_14895,N_11413,N_11823);
and U14896 (N_14896,N_11136,N_10498);
or U14897 (N_14897,N_10905,N_11144);
nor U14898 (N_14898,N_10408,N_10605);
or U14899 (N_14899,N_10612,N_11803);
nand U14900 (N_14900,N_11757,N_12452);
and U14901 (N_14901,N_11039,N_11142);
nand U14902 (N_14902,N_11873,N_10279);
and U14903 (N_14903,N_10928,N_10343);
and U14904 (N_14904,N_11935,N_11770);
or U14905 (N_14905,N_10895,N_11873);
or U14906 (N_14906,N_10460,N_12139);
and U14907 (N_14907,N_12220,N_10457);
and U14908 (N_14908,N_11573,N_11767);
nor U14909 (N_14909,N_10439,N_10596);
nand U14910 (N_14910,N_11158,N_10878);
nor U14911 (N_14911,N_10618,N_10980);
nand U14912 (N_14912,N_10624,N_11824);
or U14913 (N_14913,N_10912,N_11447);
or U14914 (N_14914,N_11857,N_12187);
nand U14915 (N_14915,N_12161,N_11574);
nand U14916 (N_14916,N_12216,N_11690);
or U14917 (N_14917,N_10696,N_11526);
xnor U14918 (N_14918,N_11975,N_11907);
nand U14919 (N_14919,N_10693,N_11413);
nor U14920 (N_14920,N_10059,N_10761);
and U14921 (N_14921,N_10568,N_12261);
and U14922 (N_14922,N_10097,N_12198);
nand U14923 (N_14923,N_11092,N_12019);
nand U14924 (N_14924,N_10415,N_10949);
nor U14925 (N_14925,N_10355,N_12364);
nand U14926 (N_14926,N_11387,N_10196);
or U14927 (N_14927,N_11431,N_11879);
or U14928 (N_14928,N_11606,N_11808);
or U14929 (N_14929,N_12097,N_10581);
nor U14930 (N_14930,N_11583,N_12013);
and U14931 (N_14931,N_11939,N_11518);
or U14932 (N_14932,N_11577,N_10995);
or U14933 (N_14933,N_12223,N_10352);
nor U14934 (N_14934,N_11186,N_10858);
and U14935 (N_14935,N_10476,N_10737);
or U14936 (N_14936,N_11232,N_11525);
nand U14937 (N_14937,N_12076,N_10471);
xnor U14938 (N_14938,N_10185,N_10710);
or U14939 (N_14939,N_12014,N_11869);
or U14940 (N_14940,N_12222,N_10738);
nor U14941 (N_14941,N_10911,N_10266);
and U14942 (N_14942,N_10183,N_12168);
or U14943 (N_14943,N_11429,N_10512);
or U14944 (N_14944,N_10152,N_10933);
nand U14945 (N_14945,N_10003,N_11833);
or U14946 (N_14946,N_11937,N_11261);
and U14947 (N_14947,N_10620,N_11762);
or U14948 (N_14948,N_11644,N_10634);
xor U14949 (N_14949,N_12126,N_10550);
and U14950 (N_14950,N_11338,N_10432);
nand U14951 (N_14951,N_11293,N_10753);
or U14952 (N_14952,N_10677,N_11304);
xor U14953 (N_14953,N_11911,N_11913);
nor U14954 (N_14954,N_11847,N_12338);
nor U14955 (N_14955,N_11506,N_10372);
and U14956 (N_14956,N_11600,N_10644);
nor U14957 (N_14957,N_10342,N_12341);
and U14958 (N_14958,N_10877,N_11650);
and U14959 (N_14959,N_12078,N_10942);
nand U14960 (N_14960,N_12325,N_11436);
nand U14961 (N_14961,N_10576,N_10826);
nor U14962 (N_14962,N_10348,N_11824);
xor U14963 (N_14963,N_11896,N_10233);
xnor U14964 (N_14964,N_11985,N_10921);
and U14965 (N_14965,N_10011,N_11695);
or U14966 (N_14966,N_10503,N_11578);
and U14967 (N_14967,N_10764,N_10583);
and U14968 (N_14968,N_12096,N_10397);
and U14969 (N_14969,N_11824,N_10940);
nor U14970 (N_14970,N_11539,N_11526);
nand U14971 (N_14971,N_11524,N_10709);
or U14972 (N_14972,N_11420,N_11710);
nand U14973 (N_14973,N_11891,N_12026);
or U14974 (N_14974,N_10200,N_12043);
and U14975 (N_14975,N_12387,N_10144);
xor U14976 (N_14976,N_11179,N_10703);
nand U14977 (N_14977,N_11844,N_12407);
or U14978 (N_14978,N_10738,N_11064);
or U14979 (N_14979,N_10990,N_10275);
xnor U14980 (N_14980,N_10702,N_12149);
nor U14981 (N_14981,N_10127,N_10096);
xnor U14982 (N_14982,N_10851,N_10496);
nor U14983 (N_14983,N_10983,N_11048);
nor U14984 (N_14984,N_10725,N_10499);
nand U14985 (N_14985,N_12405,N_11209);
nor U14986 (N_14986,N_10475,N_12021);
or U14987 (N_14987,N_11433,N_12463);
nand U14988 (N_14988,N_11213,N_11367);
xor U14989 (N_14989,N_11622,N_11355);
or U14990 (N_14990,N_12257,N_12029);
nor U14991 (N_14991,N_10517,N_10380);
nand U14992 (N_14992,N_11765,N_12100);
nor U14993 (N_14993,N_10272,N_11711);
nor U14994 (N_14994,N_11077,N_10122);
nor U14995 (N_14995,N_12101,N_10842);
nor U14996 (N_14996,N_11235,N_12357);
and U14997 (N_14997,N_12275,N_11069);
nand U14998 (N_14998,N_11638,N_11166);
nor U14999 (N_14999,N_11990,N_10746);
or U15000 (N_15000,N_13691,N_14939);
or U15001 (N_15001,N_14142,N_13377);
nand U15002 (N_15002,N_13216,N_13341);
and U15003 (N_15003,N_12555,N_13943);
nand U15004 (N_15004,N_14234,N_14928);
xor U15005 (N_15005,N_13962,N_14390);
nand U15006 (N_15006,N_14009,N_12815);
and U15007 (N_15007,N_14596,N_14669);
nand U15008 (N_15008,N_13265,N_13048);
nand U15009 (N_15009,N_14582,N_14406);
nand U15010 (N_15010,N_14442,N_14804);
and U15011 (N_15011,N_14682,N_14565);
xnor U15012 (N_15012,N_13653,N_12551);
nand U15013 (N_15013,N_13456,N_13167);
nor U15014 (N_15014,N_12697,N_12674);
nor U15015 (N_15015,N_14289,N_13967);
and U15016 (N_15016,N_14684,N_14308);
nand U15017 (N_15017,N_13482,N_14995);
nand U15018 (N_15018,N_13368,N_13965);
nor U15019 (N_15019,N_13043,N_13840);
or U15020 (N_15020,N_13066,N_14628);
xor U15021 (N_15021,N_14655,N_12964);
nand U15022 (N_15022,N_12514,N_13677);
and U15023 (N_15023,N_12721,N_13000);
nor U15024 (N_15024,N_14452,N_14643);
or U15025 (N_15025,N_14944,N_14242);
and U15026 (N_15026,N_14863,N_13885);
nor U15027 (N_15027,N_14914,N_13547);
and U15028 (N_15028,N_14206,N_14451);
and U15029 (N_15029,N_12925,N_13795);
xor U15030 (N_15030,N_12754,N_14045);
or U15031 (N_15031,N_14803,N_14194);
nand U15032 (N_15032,N_13838,N_12814);
or U15033 (N_15033,N_14150,N_14587);
nand U15034 (N_15034,N_12948,N_13569);
nand U15035 (N_15035,N_14039,N_14575);
nor U15036 (N_15036,N_12919,N_14561);
and U15037 (N_15037,N_14711,N_14794);
nand U15038 (N_15038,N_12795,N_14271);
nor U15039 (N_15039,N_14169,N_12701);
nand U15040 (N_15040,N_13997,N_13219);
or U15041 (N_15041,N_13003,N_12639);
nand U15042 (N_15042,N_13823,N_12520);
nand U15043 (N_15043,N_14338,N_13015);
and U15044 (N_15044,N_12668,N_14522);
or U15045 (N_15045,N_14346,N_12537);
nand U15046 (N_15046,N_14758,N_14245);
or U15047 (N_15047,N_13239,N_13827);
and U15048 (N_15048,N_14300,N_14331);
or U15049 (N_15049,N_13391,N_14704);
and U15050 (N_15050,N_14213,N_14347);
nor U15051 (N_15051,N_14425,N_14648);
nor U15052 (N_15052,N_12531,N_13461);
nor U15053 (N_15053,N_13487,N_13343);
nor U15054 (N_15054,N_12868,N_14267);
and U15055 (N_15055,N_12820,N_13725);
or U15056 (N_15056,N_13690,N_12669);
nor U15057 (N_15057,N_13155,N_13558);
nor U15058 (N_15058,N_14114,N_13350);
xnor U15059 (N_15059,N_13641,N_14641);
or U15060 (N_15060,N_13617,N_13615);
or U15061 (N_15061,N_14906,N_13763);
and U15062 (N_15062,N_14958,N_13836);
nor U15063 (N_15063,N_12633,N_13449);
nand U15064 (N_15064,N_14849,N_13910);
or U15065 (N_15065,N_13776,N_13579);
nor U15066 (N_15066,N_12937,N_13640);
nand U15067 (N_15067,N_12636,N_14841);
and U15068 (N_15068,N_14319,N_14264);
nand U15069 (N_15069,N_13440,N_14443);
nor U15070 (N_15070,N_12768,N_13148);
or U15071 (N_15071,N_14570,N_13489);
or U15072 (N_15072,N_13228,N_14713);
xor U15073 (N_15073,N_12658,N_14580);
or U15074 (N_15074,N_13002,N_14573);
nand U15075 (N_15075,N_12734,N_14756);
or U15076 (N_15076,N_12950,N_13137);
xor U15077 (N_15077,N_12554,N_14612);
or U15078 (N_15078,N_13866,N_14104);
or U15079 (N_15079,N_13915,N_13069);
xnor U15080 (N_15080,N_14401,N_12849);
xor U15081 (N_15081,N_13179,N_14936);
nand U15082 (N_15082,N_14901,N_13597);
and U15083 (N_15083,N_13847,N_14292);
xor U15084 (N_15084,N_14912,N_14523);
and U15085 (N_15085,N_13298,N_13671);
nand U15086 (N_15086,N_13989,N_14809);
nor U15087 (N_15087,N_13050,N_14768);
and U15088 (N_15088,N_12678,N_14248);
nand U15089 (N_15089,N_14501,N_13748);
nor U15090 (N_15090,N_14066,N_14608);
nor U15091 (N_15091,N_14024,N_14383);
nand U15092 (N_15092,N_12751,N_13986);
nand U15093 (N_15093,N_12730,N_13494);
nand U15094 (N_15094,N_13577,N_12650);
nand U15095 (N_15095,N_14447,N_12935);
nand U15096 (N_15096,N_13956,N_13978);
and U15097 (N_15097,N_14847,N_14654);
nand U15098 (N_15098,N_14133,N_12934);
or U15099 (N_15099,N_12878,N_14659);
or U15100 (N_15100,N_14620,N_12931);
or U15101 (N_15101,N_12762,N_13800);
or U15102 (N_15102,N_13764,N_14920);
nand U15103 (N_15103,N_14880,N_12975);
or U15104 (N_15104,N_13474,N_14763);
nand U15105 (N_15105,N_14496,N_13284);
nand U15106 (N_15106,N_13238,N_12728);
nor U15107 (N_15107,N_12804,N_13954);
nor U15108 (N_15108,N_14673,N_14237);
xnor U15109 (N_15109,N_13054,N_14474);
or U15110 (N_15110,N_14773,N_13151);
or U15111 (N_15111,N_13702,N_12602);
xor U15112 (N_15112,N_14785,N_13128);
or U15113 (N_15113,N_13381,N_12606);
nand U15114 (N_15114,N_13512,N_14014);
and U15115 (N_15115,N_12519,N_12969);
nand U15116 (N_15116,N_14858,N_12690);
nand U15117 (N_15117,N_13420,N_12559);
nand U15118 (N_15118,N_13871,N_13273);
and U15119 (N_15119,N_13363,N_12665);
and U15120 (N_15120,N_14305,N_12958);
xnor U15121 (N_15121,N_12769,N_13890);
nand U15122 (N_15122,N_14061,N_13177);
nor U15123 (N_15123,N_14728,N_14293);
or U15124 (N_15124,N_14649,N_12547);
xor U15125 (N_15125,N_13882,N_13629);
xnor U15126 (N_15126,N_12574,N_14355);
xor U15127 (N_15127,N_14008,N_14557);
or U15128 (N_15128,N_14661,N_14887);
nor U15129 (N_15129,N_12998,N_14201);
or U15130 (N_15130,N_14249,N_12563);
and U15131 (N_15131,N_14151,N_14019);
nand U15132 (N_15132,N_12605,N_12899);
and U15133 (N_15133,N_14945,N_13342);
or U15134 (N_15134,N_14075,N_14796);
xor U15135 (N_15135,N_12841,N_13394);
and U15136 (N_15136,N_13110,N_13322);
nor U15137 (N_15137,N_14963,N_12723);
or U15138 (N_15138,N_14179,N_13869);
nor U15139 (N_15139,N_13358,N_14644);
xor U15140 (N_15140,N_14736,N_14697);
or U15141 (N_15141,N_13765,N_14171);
nor U15142 (N_15142,N_12505,N_13451);
or U15143 (N_15143,N_13743,N_12579);
nor U15144 (N_15144,N_12595,N_14994);
or U15145 (N_15145,N_14590,N_13157);
nor U15146 (N_15146,N_13680,N_12764);
xor U15147 (N_15147,N_12576,N_13551);
nand U15148 (N_15148,N_14866,N_13738);
nor U15149 (N_15149,N_14404,N_13016);
or U15150 (N_15150,N_13643,N_14696);
or U15151 (N_15151,N_14772,N_13079);
or U15152 (N_15152,N_14765,N_13162);
or U15153 (N_15153,N_13444,N_13824);
nand U15154 (N_15154,N_14297,N_12616);
or U15155 (N_15155,N_14280,N_12749);
nor U15156 (N_15156,N_13353,N_13888);
nand U15157 (N_15157,N_12586,N_14193);
or U15158 (N_15158,N_14764,N_14145);
nor U15159 (N_15159,N_13211,N_13946);
xnor U15160 (N_15160,N_14411,N_13191);
or U15161 (N_15161,N_13424,N_14329);
nand U15162 (N_15162,N_14957,N_14750);
xnor U15163 (N_15163,N_14134,N_13485);
or U15164 (N_15164,N_14041,N_12530);
nand U15165 (N_15165,N_12737,N_13589);
nand U15166 (N_15166,N_14140,N_14354);
nor U15167 (N_15167,N_14572,N_14089);
or U15168 (N_15168,N_12620,N_13055);
nand U15169 (N_15169,N_14622,N_14291);
or U15170 (N_15170,N_13490,N_13621);
nand U15171 (N_15171,N_14818,N_14702);
and U15172 (N_15172,N_13325,N_13208);
nand U15173 (N_15173,N_13572,N_14219);
and U15174 (N_15174,N_13229,N_14258);
or U15175 (N_15175,N_14170,N_13150);
nor U15176 (N_15176,N_13886,N_13744);
xor U15177 (N_15177,N_13834,N_14893);
and U15178 (N_15178,N_12846,N_14274);
and U15179 (N_15179,N_14015,N_14371);
or U15180 (N_15180,N_14601,N_13672);
or U15181 (N_15181,N_12959,N_13053);
and U15182 (N_15182,N_13430,N_14325);
and U15183 (N_15183,N_14421,N_14011);
nand U15184 (N_15184,N_13185,N_13917);
nand U15185 (N_15185,N_12903,N_13804);
nand U15186 (N_15186,N_14985,N_14480);
nor U15187 (N_15187,N_14605,N_12558);
and U15188 (N_15188,N_12761,N_13721);
and U15189 (N_15189,N_13072,N_14327);
nor U15190 (N_15190,N_14093,N_14202);
or U15191 (N_15191,N_14666,N_13036);
nor U15192 (N_15192,N_14298,N_13518);
nor U15193 (N_15193,N_13614,N_12789);
and U15194 (N_15194,N_14453,N_14059);
nor U15195 (N_15195,N_14969,N_12865);
or U15196 (N_15196,N_13644,N_14328);
or U15197 (N_15197,N_13977,N_14657);
or U15198 (N_15198,N_14252,N_13021);
and U15199 (N_15199,N_12543,N_14177);
or U15200 (N_15200,N_13529,N_12526);
or U15201 (N_15201,N_13876,N_14716);
nor U15202 (N_15202,N_14538,N_14674);
or U15203 (N_15203,N_14568,N_12940);
nor U15204 (N_15204,N_13817,N_14313);
or U15205 (N_15205,N_14902,N_12570);
and U15206 (N_15206,N_12588,N_14854);
nor U15207 (N_15207,N_12511,N_14652);
xor U15208 (N_15208,N_14578,N_13205);
or U15209 (N_15209,N_14576,N_13710);
and U15210 (N_15210,N_14897,N_13779);
xnor U15211 (N_15211,N_14636,N_12827);
nor U15212 (N_15212,N_13771,N_12592);
nor U15213 (N_15213,N_14836,N_12945);
nand U15214 (N_15214,N_13409,N_12743);
nor U15215 (N_15215,N_13094,N_13520);
or U15216 (N_15216,N_13448,N_14820);
or U15217 (N_15217,N_12857,N_13442);
nand U15218 (N_15218,N_14875,N_13913);
and U15219 (N_15219,N_13452,N_12552);
nand U15220 (N_15220,N_14747,N_14934);
xnor U15221 (N_15221,N_12915,N_13887);
nor U15222 (N_15222,N_12837,N_12779);
nand U15223 (N_15223,N_14437,N_14868);
nor U15224 (N_15224,N_13752,N_14873);
nor U15225 (N_15225,N_14118,N_13241);
nand U15226 (N_15226,N_13249,N_12862);
nand U15227 (N_15227,N_13758,N_13545);
nor U15228 (N_15228,N_12741,N_12962);
and U15229 (N_15229,N_14220,N_14633);
nor U15230 (N_15230,N_12744,N_13315);
xnor U15231 (N_15231,N_14679,N_13684);
or U15232 (N_15232,N_13796,N_14161);
xnor U15233 (N_15233,N_13031,N_14976);
nor U15234 (N_15234,N_14068,N_13568);
and U15235 (N_15235,N_14218,N_14921);
nor U15236 (N_15236,N_12680,N_14156);
xnor U15237 (N_15237,N_14732,N_14435);
nand U15238 (N_15238,N_12933,N_12632);
or U15239 (N_15239,N_13147,N_13729);
and U15240 (N_15240,N_13117,N_14852);
nor U15241 (N_15241,N_13659,N_12802);
nand U15242 (N_15242,N_14475,N_14110);
nor U15243 (N_15243,N_13355,N_12770);
and U15244 (N_15244,N_14586,N_13180);
nor U15245 (N_15245,N_12797,N_13080);
or U15246 (N_15246,N_13961,N_12816);
nor U15247 (N_15247,N_14719,N_13385);
and U15248 (N_15248,N_12596,N_14691);
or U15249 (N_15249,N_14498,N_14414);
or U15250 (N_15250,N_14717,N_14671);
and U15251 (N_15251,N_13250,N_14513);
and U15252 (N_15252,N_12939,N_14167);
nand U15253 (N_15253,N_13240,N_13860);
nor U15254 (N_15254,N_14235,N_14367);
nand U15255 (N_15255,N_14368,N_13039);
or U15256 (N_15256,N_13767,N_14438);
or U15257 (N_15257,N_12534,N_14434);
and U15258 (N_15258,N_13559,N_12874);
or U15259 (N_15259,N_12803,N_13332);
nand U15260 (N_15260,N_14216,N_14932);
or U15261 (N_15261,N_14911,N_14079);
nand U15262 (N_15262,N_12805,N_13571);
or U15263 (N_15263,N_13206,N_14828);
or U15264 (N_15264,N_13375,N_12617);
nor U15265 (N_15265,N_13563,N_12818);
nand U15266 (N_15266,N_13495,N_13560);
and U15267 (N_15267,N_13422,N_13272);
or U15268 (N_15268,N_12826,N_13096);
or U15269 (N_15269,N_12686,N_13130);
xor U15270 (N_15270,N_13756,N_13207);
or U15271 (N_15271,N_13406,N_14665);
nor U15272 (N_15272,N_12513,N_14214);
nor U15273 (N_15273,N_14977,N_12810);
nor U15274 (N_15274,N_14953,N_13675);
xnor U15275 (N_15275,N_13881,N_13592);
nand U15276 (N_15276,N_14040,N_14705);
nand U15277 (N_15277,N_12631,N_14970);
nand U15278 (N_15278,N_13670,N_14190);
nand U15279 (N_15279,N_13694,N_13655);
xor U15280 (N_15280,N_14082,N_14834);
and U15281 (N_15281,N_14180,N_13007);
and U15282 (N_15282,N_13580,N_14028);
nor U15283 (N_15283,N_13492,N_14369);
nor U15284 (N_15284,N_12884,N_14613);
nand U15285 (N_15285,N_14023,N_14458);
nand U15286 (N_15286,N_14695,N_12649);
nand U15287 (N_15287,N_13657,N_13283);
or U15288 (N_15288,N_13222,N_13242);
or U15289 (N_15289,N_13753,N_13140);
or U15290 (N_15290,N_14121,N_14625);
or U15291 (N_15291,N_13850,N_13026);
nor U15292 (N_15292,N_12689,N_13372);
nand U15293 (N_15293,N_12822,N_13258);
and U15294 (N_15294,N_14410,N_12788);
and U15295 (N_15295,N_12597,N_14348);
and U15296 (N_15296,N_13479,N_13411);
nor U15297 (N_15297,N_14304,N_13816);
nor U15298 (N_15298,N_13300,N_14004);
nor U15299 (N_15299,N_12654,N_13435);
xor U15300 (N_15300,N_12961,N_13421);
or U15301 (N_15301,N_12640,N_13153);
nor U15302 (N_15302,N_13785,N_13530);
and U15303 (N_15303,N_12577,N_14478);
nand U15304 (N_15304,N_13981,N_14824);
xor U15305 (N_15305,N_14225,N_13646);
nor U15306 (N_15306,N_14923,N_13387);
nand U15307 (N_15307,N_12752,N_14192);
nand U15308 (N_15308,N_13221,N_13471);
nand U15309 (N_15309,N_13062,N_14987);
or U15310 (N_15310,N_13588,N_13286);
nand U15311 (N_15311,N_14098,N_13071);
and U15312 (N_15312,N_14044,N_14783);
and U15313 (N_15313,N_14962,N_14109);
nand U15314 (N_15314,N_14504,N_14314);
xor U15315 (N_15315,N_12807,N_13291);
or U15316 (N_15316,N_13699,N_12828);
and U15317 (N_15317,N_12533,N_13306);
nor U15318 (N_15318,N_13830,N_14900);
or U15319 (N_15319,N_13970,N_14191);
and U15320 (N_15320,N_14814,N_13264);
nor U15321 (N_15321,N_13994,N_12610);
nand U15322 (N_15322,N_13082,N_12974);
nand U15323 (N_15323,N_13552,N_14227);
or U15324 (N_15324,N_13232,N_13851);
or U15325 (N_15325,N_13929,N_13136);
nand U15326 (N_15326,N_13454,N_14833);
nor U15327 (N_15327,N_12589,N_13884);
and U15328 (N_15328,N_12550,N_14154);
xnor U15329 (N_15329,N_12860,N_14483);
nor U15330 (N_15330,N_13303,N_12893);
and U15331 (N_15331,N_14036,N_12707);
xnor U15332 (N_15332,N_13636,N_13109);
and U15333 (N_15333,N_13903,N_13282);
and U15334 (N_15334,N_13786,N_14647);
nand U15335 (N_15335,N_12615,N_14947);
or U15336 (N_15336,N_12825,N_13772);
nand U15337 (N_15337,N_14993,N_13061);
nand U15338 (N_15338,N_14318,N_13792);
and U15339 (N_15339,N_14553,N_13099);
and U15340 (N_15340,N_13747,N_13998);
nand U15341 (N_15341,N_13012,N_14259);
nand U15342 (N_15342,N_14488,N_14047);
or U15343 (N_15343,N_14429,N_14935);
nor U15344 (N_15344,N_14894,N_13092);
xnor U15345 (N_15345,N_14512,N_14835);
and U15346 (N_15346,N_13335,N_13731);
nor U15347 (N_15347,N_13853,N_14006);
nand U15348 (N_15348,N_14153,N_14941);
or U15349 (N_15349,N_12671,N_14574);
or U15350 (N_15350,N_14352,N_12955);
nand U15351 (N_15351,N_13750,N_12502);
nand U15352 (N_15352,N_14738,N_14287);
or U15353 (N_15353,N_13275,N_14164);
and U15354 (N_15354,N_13438,N_13344);
nor U15355 (N_15355,N_13132,N_13849);
nor U15356 (N_15356,N_13013,N_12676);
or U15357 (N_15357,N_13648,N_12838);
or U15358 (N_15358,N_14569,N_14609);
nand U15359 (N_15359,N_14283,N_12685);
or U15360 (N_15360,N_14205,N_13405);
or U15361 (N_15361,N_13959,N_14591);
or U15362 (N_15362,N_14083,N_12796);
xnor U15363 (N_15363,N_12780,N_13619);
and U15364 (N_15364,N_14929,N_13259);
or U15365 (N_15365,N_13714,N_14263);
nand U15366 (N_15366,N_14534,N_14311);
or U15367 (N_15367,N_13526,N_12667);
and U15368 (N_15368,N_14511,N_14116);
or U15369 (N_15369,N_13639,N_13618);
or U15370 (N_15370,N_14869,N_13706);
nor U15371 (N_15371,N_14251,N_13608);
xor U15372 (N_15372,N_14175,N_13466);
nor U15373 (N_15373,N_14725,N_14399);
nor U15374 (N_15374,N_13307,N_14885);
xor U15375 (N_15375,N_13141,N_13364);
and U15376 (N_15376,N_14485,N_13960);
xnor U15377 (N_15377,N_12635,N_14379);
or U15378 (N_15378,N_13832,N_12657);
xnor U15379 (N_15379,N_12835,N_12652);
nor U15380 (N_15380,N_14988,N_14088);
nor U15381 (N_15381,N_14090,N_13941);
or U15382 (N_15382,N_14334,N_13814);
or U15383 (N_15383,N_14418,N_14777);
or U15384 (N_15384,N_12833,N_13201);
or U15385 (N_15385,N_12628,N_12692);
nand U15386 (N_15386,N_14973,N_14690);
xnor U15387 (N_15387,N_14277,N_13052);
nand U15388 (N_15388,N_14279,N_13410);
nor U15389 (N_15389,N_14551,N_13582);
and U15390 (N_15390,N_12850,N_12653);
nand U15391 (N_15391,N_12883,N_14221);
or U15392 (N_15392,N_13908,N_14581);
nor U15393 (N_15393,N_14381,N_13266);
xnor U15394 (N_15394,N_13475,N_13667);
and U15395 (N_15395,N_12549,N_14720);
and U15396 (N_15396,N_13818,N_13121);
and U15397 (N_15397,N_12782,N_12691);
nand U15398 (N_15398,N_12613,N_14158);
nand U15399 (N_15399,N_12517,N_13626);
nand U15400 (N_15400,N_14731,N_12872);
and U15401 (N_15401,N_12986,N_13645);
or U15402 (N_15402,N_13277,N_13843);
xor U15403 (N_15403,N_12786,N_12876);
or U15404 (N_15404,N_14924,N_14247);
nor U15405 (N_15405,N_14617,N_14980);
nor U15406 (N_15406,N_13439,N_14391);
nor U15407 (N_15407,N_13078,N_12619);
and U15408 (N_15408,N_14943,N_14892);
or U15409 (N_15409,N_12800,N_13782);
or U15410 (N_15410,N_13801,N_14256);
or U15411 (N_15411,N_13944,N_13503);
nor U15412 (N_15412,N_13628,N_14843);
and U15413 (N_15413,N_12726,N_13203);
nor U15414 (N_15414,N_13856,N_12963);
nor U15415 (N_15415,N_14398,N_14688);
or U15416 (N_15416,N_14989,N_13927);
or U15417 (N_15417,N_14257,N_14527);
or U15418 (N_15418,N_13757,N_13178);
xor U15419 (N_15419,N_14050,N_13705);
or U15420 (N_15420,N_14281,N_13347);
nor U15421 (N_15421,N_12836,N_13164);
or U15422 (N_15422,N_14779,N_13041);
nand U15423 (N_15423,N_14461,N_14482);
or U15424 (N_15424,N_14365,N_13733);
nor U15425 (N_15425,N_13032,N_13139);
or U15426 (N_15426,N_13415,N_13658);
or U15427 (N_15427,N_12504,N_12834);
and U15428 (N_15428,N_14302,N_14431);
and U15429 (N_15429,N_12968,N_13417);
xnor U15430 (N_15430,N_13085,N_14951);
or U15431 (N_15431,N_13346,N_14959);
xor U15432 (N_15432,N_12947,N_13416);
or U15433 (N_15433,N_13126,N_13168);
nand U15434 (N_15434,N_14322,N_13815);
nand U15435 (N_15435,N_13985,N_13046);
or U15436 (N_15436,N_12867,N_13407);
nor U15437 (N_15437,N_14675,N_12670);
nand U15438 (N_15438,N_14340,N_12627);
nor U15439 (N_15439,N_14749,N_12706);
or U15440 (N_15440,N_13345,N_14559);
nand U15441 (N_15441,N_13635,N_14510);
or U15442 (N_15442,N_14846,N_13649);
or U15443 (N_15443,N_13497,N_14373);
and U15444 (N_15444,N_13980,N_14113);
nand U15445 (N_15445,N_13510,N_12854);
nor U15446 (N_15446,N_12661,N_13361);
nand U15447 (N_15447,N_14931,N_12952);
nor U15448 (N_15448,N_12608,N_13236);
nand U15449 (N_15449,N_13730,N_14394);
xor U15450 (N_15450,N_14490,N_14734);
nand U15451 (N_15451,N_13097,N_14919);
or U15452 (N_15452,N_13642,N_14094);
nor U15453 (N_15453,N_14428,N_14817);
and U15454 (N_15454,N_14739,N_13761);
nor U15455 (N_15455,N_14801,N_14402);
and U15456 (N_15456,N_14471,N_14683);
nand U15457 (N_15457,N_14997,N_13247);
and U15458 (N_15458,N_12532,N_12949);
and U15459 (N_15459,N_14424,N_13175);
nor U15460 (N_15460,N_14775,N_13144);
nor U15461 (N_15461,N_13540,N_14057);
nor U15462 (N_15462,N_14968,N_12708);
or U15463 (N_15463,N_14189,N_14978);
nor U15464 (N_15464,N_14938,N_13057);
nor U15465 (N_15465,N_12573,N_14886);
nor U15466 (N_15466,N_14799,N_14239);
nand U15467 (N_15467,N_13324,N_13114);
or U15468 (N_15468,N_13715,N_14981);
nand U15469 (N_15469,N_12548,N_14624);
and U15470 (N_15470,N_14518,N_13573);
or U15471 (N_15471,N_14427,N_14339);
and U15472 (N_15472,N_12528,N_12888);
nand U15473 (N_15473,N_13855,N_13029);
nand U15474 (N_15474,N_14260,N_13987);
or U15475 (N_15475,N_14455,N_13603);
nand U15476 (N_15476,N_14700,N_13873);
nand U15477 (N_15477,N_13488,N_14528);
nor U15478 (N_15478,N_14844,N_14080);
nand U15479 (N_15479,N_13386,N_12951);
and U15480 (N_15480,N_12845,N_13875);
or U15481 (N_15481,N_14262,N_13297);
nand U15482 (N_15482,N_13477,N_13230);
nor U15483 (N_15483,N_12644,N_14558);
nor U15484 (N_15484,N_14701,N_13251);
or U15485 (N_15485,N_12847,N_14026);
and U15486 (N_15486,N_13637,N_14692);
and U15487 (N_15487,N_14129,N_14433);
nand U15488 (N_15488,N_13576,N_13983);
xnor U15489 (N_15489,N_13686,N_12760);
nor U15490 (N_15490,N_13634,N_12909);
nand U15491 (N_15491,N_14630,N_14069);
nor U15492 (N_15492,N_12582,N_14400);
and U15493 (N_15493,N_14464,N_14627);
nor U15494 (N_15494,N_14806,N_14386);
xnor U15495 (N_15495,N_13351,N_13919);
and U15496 (N_15496,N_13755,N_13696);
nand U15497 (N_15497,N_14484,N_14018);
or U15498 (N_15498,N_14419,N_14529);
and U15499 (N_15499,N_13314,N_12905);
xnor U15500 (N_15500,N_13383,N_13660);
nand U15501 (N_15501,N_12731,N_13171);
or U15502 (N_15502,N_13267,N_14423);
nor U15503 (N_15503,N_12509,N_13458);
nand U15504 (N_15504,N_13189,N_14942);
nand U15505 (N_15505,N_14748,N_14766);
nand U15506 (N_15506,N_14099,N_13703);
nand U15507 (N_15507,N_13524,N_13010);
nor U15508 (N_15508,N_13227,N_14002);
nor U15509 (N_15509,N_13371,N_14672);
and U15510 (N_15510,N_13278,N_13237);
nor U15511 (N_15511,N_13311,N_14030);
nand U15512 (N_15512,N_14831,N_13587);
nand U15513 (N_15513,N_13604,N_14375);
or U15514 (N_15514,N_12594,N_12750);
and U15515 (N_15515,N_14653,N_13596);
nand U15516 (N_15516,N_14729,N_13525);
or U15517 (N_15517,N_13318,N_13709);
and U15518 (N_15518,N_13476,N_12623);
nor U15519 (N_15519,N_14349,N_13065);
or U15520 (N_15520,N_14583,N_13500);
or U15521 (N_15521,N_14462,N_14724);
nor U15522 (N_15522,N_12812,N_14065);
xor U15523 (N_15523,N_14667,N_13357);
nor U15524 (N_15524,N_12946,N_12997);
nand U15525 (N_15525,N_13937,N_14781);
xor U15526 (N_15526,N_12976,N_13483);
xor U15527 (N_15527,N_14905,N_13538);
nor U15528 (N_15528,N_14898,N_12932);
nand U15529 (N_15529,N_14640,N_12659);
or U15530 (N_15530,N_14460,N_14007);
xor U15531 (N_15531,N_13870,N_14309);
and U15532 (N_15532,N_14223,N_12587);
and U15533 (N_15533,N_12882,N_14187);
nand U15534 (N_15534,N_13154,N_14530);
or U15535 (N_15535,N_13839,N_14862);
nor U15536 (N_15536,N_12518,N_14502);
nor U15537 (N_15537,N_14787,N_12508);
nand U15538 (N_15538,N_13067,N_13598);
or U15539 (N_15539,N_14566,N_13907);
and U15540 (N_15540,N_13304,N_13793);
xnor U15541 (N_15541,N_14499,N_13163);
or U15542 (N_15542,N_12618,N_14255);
nor U15543 (N_15543,N_12718,N_14872);
nor U15544 (N_15544,N_13112,N_12638);
xor U15545 (N_15545,N_12675,N_12540);
or U15546 (N_15546,N_13399,N_14182);
nor U15547 (N_15547,N_14477,N_13382);
or U15548 (N_15548,N_12848,N_14965);
or U15549 (N_15549,N_13678,N_13692);
nand U15550 (N_15550,N_12656,N_13398);
nand U15551 (N_15551,N_12572,N_12831);
nand U15552 (N_15552,N_14324,N_14495);
and U15553 (N_15553,N_14983,N_14303);
and U15554 (N_15554,N_13460,N_13292);
and U15555 (N_15555,N_13513,N_14238);
nor U15556 (N_15556,N_13607,N_13950);
nor U15557 (N_15557,N_14544,N_14160);
and U15558 (N_15558,N_13905,N_14058);
nor U15559 (N_15559,N_14366,N_13234);
nor U15560 (N_15560,N_14615,N_13939);
and U15561 (N_15561,N_14735,N_13794);
nand U15562 (N_15562,N_14095,N_13739);
and U15563 (N_15563,N_13688,N_14209);
and U15564 (N_15564,N_13294,N_12539);
or U15565 (N_15565,N_14712,N_14064);
nor U15566 (N_15566,N_12856,N_14122);
nand U15567 (N_15567,N_13214,N_13811);
nand U15568 (N_15568,N_14147,N_13581);
or U15569 (N_15569,N_13700,N_13601);
and U15570 (N_15570,N_12759,N_13627);
nand U15571 (N_15571,N_14326,N_13555);
xor U15572 (N_15572,N_14535,N_13106);
xnor U15573 (N_15573,N_13414,N_14864);
nor U15574 (N_15574,N_12973,N_13682);
xor U15575 (N_15575,N_13182,N_13911);
and U15576 (N_15576,N_12722,N_13975);
and U15577 (N_15577,N_14784,N_14357);
nand U15578 (N_15578,N_14103,N_14541);
and U15579 (N_15579,N_13337,N_13124);
nand U15580 (N_15580,N_13481,N_14853);
or U15581 (N_15581,N_14208,N_12568);
or U15582 (N_15582,N_14607,N_14904);
or U15583 (N_15583,N_14466,N_13537);
nand U15584 (N_15584,N_14403,N_13697);
nor U15585 (N_15585,N_13328,N_14699);
nand U15586 (N_15586,N_13486,N_14276);
and U15587 (N_15587,N_12719,N_13842);
or U15588 (N_15588,N_13561,N_14500);
nand U15589 (N_15589,N_12736,N_13200);
or U15590 (N_15590,N_13436,N_13253);
nor U15591 (N_15591,N_12971,N_14621);
nand U15592 (N_15592,N_12791,N_13244);
nand U15593 (N_15593,N_13491,N_14611);
and U15594 (N_15594,N_12717,N_14708);
and U15595 (N_15595,N_14174,N_12709);
xnor U15596 (N_15596,N_14788,N_14063);
nand U15597 (N_15597,N_14010,N_14888);
nor U15598 (N_15598,N_12724,N_13088);
nor U15599 (N_15599,N_13673,N_14166);
and U15600 (N_15600,N_13075,N_14966);
xnor U15601 (N_15601,N_13101,N_12566);
nand U15602 (N_15602,N_14323,N_12673);
and U15603 (N_15603,N_12702,N_12757);
and U15604 (N_15604,N_14714,N_14417);
nor U15605 (N_15605,N_14233,N_14519);
nand U15606 (N_15606,N_12793,N_12980);
nor U15607 (N_15607,N_14602,N_13852);
nor U15608 (N_15608,N_13622,N_12672);
nand U15609 (N_15609,N_14645,N_13465);
and U15610 (N_15610,N_14086,N_13949);
nor U15611 (N_15611,N_13566,N_12965);
nand U15612 (N_15612,N_12853,N_13519);
nor U15613 (N_15613,N_13698,N_13135);
nand U15614 (N_15614,N_13556,N_14056);
nor U15615 (N_15615,N_12527,N_13567);
nand U15616 (N_15616,N_12604,N_13664);
and U15617 (N_15617,N_14244,N_14884);
or U15618 (N_15618,N_14203,N_13202);
nor U15619 (N_15619,N_14964,N_12535);
or U15620 (N_15620,N_14533,N_14222);
xor U15621 (N_15621,N_14468,N_12981);
nand U15622 (N_15622,N_13844,N_12688);
and U15623 (N_15623,N_12560,N_12683);
xnor U15624 (N_15624,N_13741,N_13701);
nor U15625 (N_15625,N_14102,N_13197);
xnor U15626 (N_15626,N_14635,N_13854);
nand U15627 (N_15627,N_14955,N_13945);
nor U15628 (N_15628,N_13769,N_13810);
nand U15629 (N_15629,N_14038,N_13914);
and U15630 (N_15630,N_14646,N_13656);
and U15631 (N_15631,N_13212,N_13225);
nand U15632 (N_15632,N_14560,N_12712);
or U15633 (N_15633,N_14364,N_13963);
nand U15634 (N_15634,N_12742,N_13433);
nor U15635 (N_15635,N_12637,N_13865);
nor U15636 (N_15636,N_14017,N_14005);
nand U15637 (N_15637,N_12787,N_14584);
nor U15638 (N_15638,N_13742,N_14146);
xor U15639 (N_15639,N_12747,N_12996);
nor U15640 (N_15640,N_13119,N_14703);
xnor U15641 (N_15641,N_13302,N_14465);
nor U15642 (N_15642,N_12809,N_13198);
xnor U15643 (N_15643,N_13923,N_14589);
or U15644 (N_15644,N_14178,N_12625);
and U15645 (N_15645,N_14012,N_13534);
nand U15646 (N_15646,N_13218,N_13496);
or U15647 (N_15647,N_13883,N_13310);
nand U15648 (N_15648,N_12612,N_13784);
nand U15649 (N_15649,N_14930,N_12711);
nand U15650 (N_15650,N_13352,N_13695);
nor U15651 (N_15651,N_14163,N_13204);
and U15652 (N_15652,N_13480,N_12908);
and U15653 (N_15653,N_14415,N_14916);
nand U15654 (N_15654,N_14554,N_13102);
nand U15655 (N_15655,N_14895,N_14998);
nand U15656 (N_15656,N_12641,N_13156);
nor U15657 (N_15657,N_12902,N_13257);
xor U15658 (N_15658,N_13775,N_13143);
nor U15659 (N_15659,N_12599,N_13271);
nor U15660 (N_15660,N_13517,N_12763);
nor U15661 (N_15661,N_14141,N_12503);
or U15662 (N_15662,N_14742,N_14100);
xor U15663 (N_15663,N_14889,N_12808);
nor U15664 (N_15664,N_12694,N_13040);
nor U15665 (N_15665,N_14450,N_14722);
nand U15666 (N_15666,N_14060,N_14971);
nand U15667 (N_15667,N_14780,N_13321);
or U15668 (N_15668,N_12978,N_14927);
xor U15669 (N_15669,N_14405,N_13833);
or U15670 (N_15670,N_14025,N_14922);
xnor U15671 (N_15671,N_14793,N_12651);
nor U15672 (N_15672,N_13789,N_12755);
nand U15673 (N_15673,N_14092,N_14867);
or U15674 (N_15674,N_12611,N_13129);
nand U15675 (N_15675,N_13017,N_13902);
nor U15676 (N_15676,N_14917,N_12607);
nor U15677 (N_15677,N_14155,N_14909);
nand U15678 (N_15678,N_13630,N_12844);
nand U15679 (N_15679,N_14120,N_12544);
and U15680 (N_15680,N_14614,N_12821);
or U15681 (N_15681,N_13327,N_14307);
xor U15682 (N_15682,N_13360,N_14821);
and U15683 (N_15683,N_14562,N_14940);
or U15684 (N_15684,N_12515,N_13380);
and U15685 (N_15685,N_13651,N_13665);
nand U15686 (N_15686,N_14694,N_13781);
xnor U15687 (N_15687,N_14360,N_13428);
nand U15688 (N_15688,N_14320,N_14130);
and U15689 (N_15689,N_13991,N_12601);
nand U15690 (N_15690,N_14588,N_13427);
nor U15691 (N_15691,N_14105,N_14542);
and U15692 (N_15692,N_12994,N_14377);
or U15693 (N_15693,N_14157,N_13425);
or U15694 (N_15694,N_14273,N_13846);
xnor U15695 (N_15695,N_14546,N_13762);
nand U15696 (N_15696,N_13447,N_14476);
nand U15697 (N_15697,N_13390,N_13149);
and U15698 (N_15698,N_12567,N_13624);
and U15699 (N_15699,N_13625,N_14637);
nand U15700 (N_15700,N_12677,N_13766);
and U15701 (N_15701,N_13183,N_13333);
or U15702 (N_15702,N_12662,N_14979);
xnor U15703 (N_15703,N_13095,N_13899);
xnor U15704 (N_15704,N_13858,N_13864);
or U15705 (N_15705,N_14123,N_14376);
and U15706 (N_15706,N_14198,N_14165);
and U15707 (N_15707,N_14333,N_13536);
nor U15708 (N_15708,N_13925,N_13720);
nor U15709 (N_15709,N_13195,N_13933);
or U15710 (N_15710,N_14131,N_13976);
and U15711 (N_15711,N_14778,N_12938);
xnor U15712 (N_15712,N_13274,N_13993);
nand U15713 (N_15713,N_13930,N_13091);
nand U15714 (N_15714,N_13803,N_13431);
nor U15715 (N_15715,N_14001,N_12811);
nor U15716 (N_15716,N_13152,N_12732);
and U15717 (N_15717,N_14350,N_14891);
and U15718 (N_15718,N_13606,N_13770);
and U15719 (N_15719,N_14856,N_13073);
or U15720 (N_15720,N_14552,N_13252);
nand U15721 (N_15721,N_14210,N_14454);
nand U15722 (N_15722,N_12512,N_13366);
and U15723 (N_15723,N_13404,N_13463);
nand U15724 (N_15724,N_13751,N_13279);
or U15725 (N_15725,N_14358,N_14967);
nor U15726 (N_15726,N_12705,N_13254);
or U15727 (N_15727,N_14016,N_12898);
and U15728 (N_15728,N_13125,N_14899);
nor U15729 (N_15729,N_14861,N_14111);
and U15730 (N_15730,N_14752,N_12900);
or U15731 (N_15731,N_14207,N_13533);
nor U15732 (N_15732,N_14996,N_14049);
nor U15733 (N_15733,N_13269,N_12591);
and U15734 (N_15734,N_13432,N_13777);
and U15735 (N_15735,N_13521,N_13170);
or U15736 (N_15736,N_12993,N_12891);
or U15737 (N_15737,N_13403,N_14693);
or U15738 (N_15738,N_13022,N_14631);
nor U15739 (N_15739,N_13246,N_12580);
or U15740 (N_15740,N_13379,N_12507);
xnor U15741 (N_15741,N_13570,N_14361);
nand U15742 (N_15742,N_12614,N_13831);
or U15743 (N_15743,N_14420,N_14789);
nand U15744 (N_15744,N_13260,N_14345);
xor U15745 (N_15745,N_14837,N_14479);
nand U15746 (N_15746,N_13210,N_13504);
nand U15747 (N_15747,N_13472,N_14332);
or U15748 (N_15748,N_13909,N_14850);
or U15749 (N_15749,N_14550,N_13791);
and U15750 (N_15750,N_14879,N_12892);
nand U15751 (N_15751,N_14489,N_13467);
and U15752 (N_15752,N_14830,N_14493);
nor U15753 (N_15753,N_14215,N_14035);
or U15754 (N_15754,N_14228,N_14579);
nand U15755 (N_15755,N_14469,N_14508);
xor U15756 (N_15756,N_14790,N_12866);
xor U15757 (N_15757,N_13243,N_13401);
nand U15758 (N_15758,N_14288,N_12720);
nor U15759 (N_15759,N_14960,N_13138);
nor U15760 (N_15760,N_14555,N_13058);
nand U15761 (N_15761,N_14459,N_13196);
nor U15762 (N_15762,N_14547,N_12629);
or U15763 (N_15763,N_12936,N_14946);
and U15764 (N_15764,N_14343,N_13235);
and U15765 (N_15765,N_12873,N_13122);
nor U15766 (N_15766,N_14991,N_13001);
xnor U15767 (N_15767,N_14925,N_13370);
xor U15768 (N_15768,N_14243,N_14229);
nand U15769 (N_15769,N_13685,N_14548);
and U15770 (N_15770,N_14372,N_13532);
nand U15771 (N_15771,N_13118,N_14974);
or U15772 (N_15772,N_13727,N_13397);
nor U15773 (N_15773,N_14148,N_12989);
and U15774 (N_15774,N_13107,N_14851);
nor U15775 (N_15775,N_14101,N_13502);
xor U15776 (N_15776,N_14396,N_14076);
and U15777 (N_15777,N_14126,N_14585);
nor U15778 (N_15778,N_14676,N_13668);
and U15779 (N_15779,N_13108,N_14592);
or U15780 (N_15780,N_14441,N_13457);
nand U15781 (N_15781,N_12583,N_14825);
nand U15782 (N_15782,N_13453,N_13841);
nor U15783 (N_15783,N_12626,N_13402);
nor U15784 (N_15784,N_12877,N_12875);
nand U15785 (N_15785,N_14409,N_12500);
or U15786 (N_15786,N_14757,N_13590);
and U15787 (N_15787,N_13778,N_12748);
nor U15788 (N_15788,N_14380,N_13938);
nor U15789 (N_15789,N_13464,N_14449);
or U15790 (N_15790,N_13188,N_14278);
and U15791 (N_15791,N_14246,N_13829);
and U15792 (N_15792,N_14819,N_13806);
xnor U15793 (N_15793,N_14549,N_13280);
xor U15794 (N_15794,N_13982,N_14426);
or U15795 (N_15795,N_13224,N_13891);
xor U15796 (N_15796,N_12646,N_14754);
nor U15797 (N_15797,N_14623,N_14275);
and U15798 (N_15798,N_13857,N_14800);
nor U15799 (N_15799,N_14685,N_12879);
and U15800 (N_15800,N_13553,N_12863);
or U15801 (N_15801,N_12861,N_13217);
nor U15802 (N_15802,N_12571,N_14362);
or U15803 (N_15803,N_13223,N_12967);
nor U15804 (N_15804,N_13184,N_14108);
nor U15805 (N_15805,N_13484,N_13340);
or U15806 (N_15806,N_14112,N_14954);
nor U15807 (N_15807,N_14737,N_13133);
nor U15808 (N_15808,N_13924,N_14839);
nand U15809 (N_15809,N_14387,N_12660);
nand U15810 (N_15810,N_13936,N_13105);
and U15811 (N_15811,N_14412,N_13018);
nor U15812 (N_15812,N_12995,N_13774);
nor U15813 (N_15813,N_14597,N_13550);
and U15814 (N_15814,N_12727,N_14933);
nor U15815 (N_15815,N_14707,N_12536);
and U15816 (N_15816,N_14539,N_14168);
nor U15817 (N_15817,N_14062,N_12801);
nor U15818 (N_15818,N_12889,N_13650);
or U15819 (N_15819,N_13728,N_13514);
nor U15820 (N_15820,N_12710,N_13393);
nor U15821 (N_15821,N_12765,N_12663);
xnor U15822 (N_15822,N_13190,N_13359);
nand U15823 (N_15823,N_13493,N_12784);
nor U15824 (N_15824,N_14660,N_12634);
or U15825 (N_15825,N_14043,N_13159);
xnor U15826 (N_15826,N_12885,N_12979);
and U15827 (N_15827,N_13042,N_13892);
nand U15828 (N_15828,N_14265,N_13916);
nor U15829 (N_15829,N_12767,N_13542);
and U15830 (N_15830,N_13600,N_13509);
nand U15831 (N_15831,N_12943,N_14950);
nand U15832 (N_15832,N_13546,N_13922);
nand U15833 (N_15833,N_12881,N_14741);
xor U15834 (N_15834,N_14139,N_14382);
or U15835 (N_15835,N_14577,N_13583);
nor U15836 (N_15836,N_14857,N_12927);
and U15837 (N_15837,N_13362,N_14270);
and U15838 (N_15838,N_13666,N_13068);
nand U15839 (N_15839,N_13093,N_13037);
nand U15840 (N_15840,N_12740,N_12983);
nand U15841 (N_15841,N_13652,N_14286);
xnor U15842 (N_15842,N_13169,N_13783);
and U15843 (N_15843,N_13711,N_14808);
nand U15844 (N_15844,N_13400,N_13330);
nand U15845 (N_15845,N_14771,N_14715);
and U15846 (N_15846,N_13059,N_13988);
nor U15847 (N_15847,N_12817,N_12565);
or U15848 (N_15848,N_13429,N_12895);
or U15849 (N_15849,N_14651,N_13165);
nand U15850 (N_15850,N_12987,N_13878);
and U15851 (N_15851,N_14029,N_13231);
nor U15852 (N_15852,N_13047,N_13564);
nor U15853 (N_15853,N_13541,N_14310);
and U15854 (N_15854,N_13317,N_14473);
nor U15855 (N_15855,N_12556,N_13808);
nand U15856 (N_15856,N_14726,N_14827);
and U15857 (N_15857,N_13798,N_12840);
and U15858 (N_15858,N_13740,N_12645);
and U15859 (N_15859,N_14776,N_13735);
nand U15860 (N_15860,N_14516,N_14294);
or U15861 (N_15861,N_13620,N_14903);
nor U15862 (N_15862,N_14730,N_14759);
nand U15863 (N_15863,N_12842,N_13612);
nand U15864 (N_15864,N_12564,N_13220);
nand U15865 (N_15865,N_14444,N_14106);
xor U15866 (N_15866,N_12970,N_12916);
or U15867 (N_15867,N_13396,N_14224);
or U15868 (N_15868,N_13413,N_14467);
and U15869 (N_15869,N_13104,N_12960);
xor U15870 (N_15870,N_14982,N_12523);
or U15871 (N_15871,N_13984,N_13979);
or U15872 (N_15872,N_14077,N_13194);
or U15873 (N_15873,N_13687,N_14619);
or U15874 (N_15874,N_14027,N_12516);
or U15875 (N_15875,N_13123,N_14037);
or U15876 (N_15876,N_14718,N_12999);
nand U15877 (N_15877,N_12859,N_13193);
or U15878 (N_15878,N_14337,N_14472);
and U15879 (N_15879,N_13874,N_13028);
or U15880 (N_15880,N_14638,N_14436);
or U15881 (N_15881,N_14097,N_12773);
nor U15882 (N_15882,N_14021,N_14604);
and U15883 (N_15883,N_12771,N_13056);
nand U15884 (N_15884,N_12624,N_13378);
nor U15885 (N_15885,N_13384,N_14107);
nor U15886 (N_15886,N_14341,N_13951);
nand U15887 (N_15887,N_12546,N_14197);
and U15888 (N_15888,N_12924,N_13395);
xor U15889 (N_15889,N_12887,N_13861);
or U15890 (N_15890,N_13926,N_14515);
nor U15891 (N_15891,N_13906,N_12914);
or U15892 (N_15892,N_12529,N_13921);
nor U15893 (N_15893,N_13426,N_12642);
nand U15894 (N_15894,N_13008,N_14020);
or U15895 (N_15895,N_13441,N_13586);
or U15896 (N_15896,N_14883,N_14517);
nor U15897 (N_15897,N_12982,N_14204);
nand U15898 (N_15898,N_12829,N_14152);
nand U15899 (N_15899,N_14363,N_13365);
xor U15900 (N_15900,N_14567,N_13797);
and U15901 (N_15901,N_13373,N_13522);
nand U15902 (N_15902,N_14136,N_12666);
and U15903 (N_15903,N_14272,N_13868);
nand U15904 (N_15904,N_14162,N_14791);
nor U15905 (N_15905,N_14316,N_12521);
nand U15906 (N_15906,N_13585,N_14440);
and U15907 (N_15907,N_13034,N_12926);
nand U15908 (N_15908,N_14948,N_13470);
nor U15909 (N_15909,N_13712,N_14003);
and U15910 (N_15910,N_12545,N_14593);
and U15911 (N_15911,N_14301,N_14046);
and U15912 (N_15912,N_13131,N_13948);
xor U15913 (N_15913,N_13952,N_14124);
nand U15914 (N_15914,N_14048,N_14031);
nor U15915 (N_15915,N_14487,N_13263);
or U15916 (N_15916,N_12944,N_13828);
xnor U15917 (N_15917,N_13880,N_13935);
nor U15918 (N_15918,N_14378,N_14642);
nand U15919 (N_15919,N_12806,N_14890);
nor U15920 (N_15920,N_14677,N_13459);
or U15921 (N_15921,N_12990,N_12541);
or U15922 (N_15922,N_12942,N_14990);
xnor U15923 (N_15923,N_12830,N_12753);
nor U15924 (N_15924,N_13276,N_13044);
or U15925 (N_15925,N_12648,N_14710);
nand U15926 (N_15926,N_13931,N_14571);
nand U15927 (N_15927,N_14236,N_14137);
nand U15928 (N_15928,N_13693,N_14826);
nand U15929 (N_15929,N_13215,N_13732);
nor U15930 (N_15930,N_14370,N_13166);
xor U15931 (N_15931,N_14543,N_14448);
xor U15932 (N_15932,N_12775,N_14845);
or U15933 (N_15933,N_13074,N_13565);
nand U15934 (N_15934,N_12603,N_13301);
and U15935 (N_15935,N_14531,N_13134);
and U15936 (N_15936,N_13647,N_13898);
nand U15937 (N_15937,N_13098,N_13100);
and U15938 (N_15938,N_14144,N_13953);
nor U15939 (N_15939,N_13623,N_14000);
or U15940 (N_15940,N_13631,N_14913);
or U15941 (N_15941,N_13848,N_14013);
and U15942 (N_15942,N_14397,N_13103);
or U15943 (N_15943,N_12581,N_14439);
or U15944 (N_15944,N_14336,N_14874);
or U15945 (N_15945,N_14992,N_14698);
nor U15946 (N_15946,N_12561,N_14284);
and U15947 (N_15947,N_13349,N_14486);
nor U15948 (N_15948,N_12890,N_13423);
nand U15949 (N_15949,N_13863,N_13268);
nand U15950 (N_15950,N_12858,N_12735);
nand U15951 (N_15951,N_14594,N_13087);
xnor U15952 (N_15952,N_14525,N_13719);
nand U15953 (N_15953,N_13011,N_14878);
nand U15954 (N_15954,N_13897,N_14782);
nor U15955 (N_15955,N_13064,N_13900);
nand U15956 (N_15956,N_14230,N_14663);
or U15957 (N_15957,N_13030,N_14091);
nand U15958 (N_15958,N_13111,N_13964);
nor U15959 (N_15959,N_12922,N_14721);
xnor U15960 (N_15960,N_12794,N_13116);
nand U15961 (N_15961,N_14389,N_14795);
nor U15962 (N_15962,N_12985,N_14135);
xor U15963 (N_15963,N_14034,N_13528);
xnor U15964 (N_15964,N_13802,N_14149);
and U15965 (N_15965,N_13669,N_13348);
nor U15966 (N_15966,N_14956,N_14070);
and U15967 (N_15967,N_12852,N_13516);
nand U15968 (N_15968,N_12832,N_14430);
nor U15969 (N_15969,N_14395,N_14813);
or U15970 (N_15970,N_13845,N_13319);
nand U15971 (N_15971,N_12930,N_14117);
nand U15972 (N_15972,N_14385,N_13233);
nor U15973 (N_15973,N_14792,N_13127);
nor U15974 (N_15974,N_12739,N_14743);
or U15975 (N_15975,N_14687,N_12600);
or U15976 (N_15976,N_12774,N_13009);
or U15977 (N_15977,N_14681,N_13535);
nor U15978 (N_15978,N_14413,N_12609);
or U15979 (N_15979,N_13070,N_14751);
or U15980 (N_15980,N_14556,N_14632);
nor U15981 (N_15981,N_14618,N_14755);
nand U15982 (N_15982,N_12593,N_12781);
nor U15983 (N_15983,N_13515,N_13611);
nand U15984 (N_15984,N_13973,N_13033);
or U15985 (N_15985,N_12598,N_14172);
or U15986 (N_15986,N_14505,N_13942);
or U15987 (N_15987,N_13872,N_13575);
nor U15988 (N_15988,N_13299,N_14374);
nor U15989 (N_15989,N_14081,N_14503);
and U15990 (N_15990,N_13549,N_13005);
nor U15991 (N_15991,N_13209,N_13038);
xnor U15992 (N_15992,N_13045,N_13947);
or U15993 (N_15993,N_13609,N_14802);
nor U15994 (N_15994,N_13014,N_14598);
and U15995 (N_15995,N_12643,N_14877);
or U15996 (N_15996,N_14926,N_14078);
and U15997 (N_15997,N_13181,N_13826);
nand U15998 (N_15998,N_12896,N_13734);
nor U15999 (N_15999,N_13120,N_12542);
and U16000 (N_16000,N_14838,N_14805);
nand U16001 (N_16001,N_13389,N_14521);
nor U16002 (N_16002,N_13261,N_13726);
nor U16003 (N_16003,N_14232,N_14456);
xnor U16004 (N_16004,N_13248,N_13501);
and U16005 (N_16005,N_14506,N_14356);
or U16006 (N_16006,N_14999,N_13633);
or U16007 (N_16007,N_14786,N_14860);
nor U16008 (N_16008,N_13638,N_14744);
xor U16009 (N_16009,N_14067,N_14159);
nand U16010 (N_16010,N_14285,N_13616);
xor U16011 (N_16011,N_14033,N_14071);
nor U16012 (N_16012,N_12928,N_14603);
and U16013 (N_16013,N_14686,N_14344);
and U16014 (N_16014,N_14908,N_12953);
or U16015 (N_16015,N_13809,N_14882);
xnor U16016 (N_16016,N_14746,N_14727);
nand U16017 (N_16017,N_13192,N_14042);
nand U16018 (N_16018,N_14188,N_13506);
nand U16019 (N_16019,N_13369,N_14815);
xor U16020 (N_16020,N_13499,N_12823);
nand U16021 (N_16021,N_13593,N_13213);
nor U16022 (N_16022,N_12647,N_12772);
nor U16023 (N_16023,N_13505,N_12501);
or U16024 (N_16024,N_12704,N_14446);
xnor U16025 (N_16025,N_14706,N_14599);
or U16026 (N_16026,N_13990,N_13807);
or U16027 (N_16027,N_14072,N_13527);
nor U16028 (N_16028,N_13821,N_13245);
nor U16029 (N_16029,N_13450,N_13006);
nand U16030 (N_16030,N_12729,N_14342);
or U16031 (N_16031,N_14055,N_13704);
nand U16032 (N_16032,N_13090,N_13895);
nand U16033 (N_16033,N_13754,N_13051);
nand U16034 (N_16034,N_14545,N_13724);
nor U16035 (N_16035,N_13287,N_12557);
nor U16036 (N_16036,N_14972,N_13308);
nor U16037 (N_16037,N_13478,N_12851);
xor U16038 (N_16038,N_12525,N_13437);
or U16039 (N_16039,N_13004,N_14975);
or U16040 (N_16040,N_13296,N_13089);
and U16041 (N_16041,N_13173,N_12869);
nand U16042 (N_16042,N_14760,N_12696);
xor U16043 (N_16043,N_13918,N_12695);
nor U16044 (N_16044,N_14384,N_14085);
or U16045 (N_16045,N_13610,N_13312);
xor U16046 (N_16046,N_14176,N_13788);
nor U16047 (N_16047,N_12713,N_14445);
nand U16048 (N_16048,N_13662,N_12630);
or U16049 (N_16049,N_13226,N_14183);
xnor U16050 (N_16050,N_14132,N_14949);
nor U16051 (N_16051,N_14812,N_13115);
nand U16052 (N_16052,N_13446,N_14870);
and U16053 (N_16053,N_13584,N_12506);
and U16054 (N_16054,N_12522,N_12910);
or U16055 (N_16055,N_13035,N_14610);
nand U16056 (N_16056,N_14984,N_13859);
xor U16057 (N_16057,N_14053,N_13024);
xor U16058 (N_16058,N_12921,N_13160);
nand U16059 (N_16059,N_12758,N_14470);
and U16060 (N_16060,N_14626,N_13889);
nor U16061 (N_16061,N_13958,N_13049);
or U16062 (N_16062,N_12917,N_13812);
nand U16063 (N_16063,N_13749,N_12901);
xnor U16064 (N_16064,N_13974,N_14054);
nor U16065 (N_16065,N_14295,N_13408);
nor U16066 (N_16066,N_13605,N_13443);
nand U16067 (N_16067,N_12590,N_13689);
and U16068 (N_16068,N_12954,N_12569);
nand U16069 (N_16069,N_13418,N_13172);
nor U16070 (N_16070,N_14432,N_14634);
and U16071 (N_16071,N_14810,N_13896);
or U16072 (N_16072,N_14865,N_13683);
or U16073 (N_16073,N_14855,N_13928);
nor U16074 (N_16074,N_12991,N_13562);
xnor U16075 (N_16075,N_12871,N_12578);
nand U16076 (N_16076,N_14200,N_14335);
and U16077 (N_16077,N_13813,N_12988);
nor U16078 (N_16078,N_14709,N_14952);
and U16079 (N_16079,N_12585,N_13992);
nor U16080 (N_16080,N_13957,N_14299);
nor U16081 (N_16081,N_13663,N_14761);
or U16082 (N_16082,N_14052,N_14388);
or U16083 (N_16083,N_12776,N_14296);
nand U16084 (N_16084,N_13256,N_13174);
nor U16085 (N_16085,N_13412,N_13877);
and U16086 (N_16086,N_14798,N_13632);
and U16087 (N_16087,N_13820,N_14457);
or U16088 (N_16088,N_13867,N_12715);
nor U16089 (N_16089,N_13674,N_13835);
and U16090 (N_16090,N_13305,N_12700);
and U16091 (N_16091,N_14564,N_14910);
and U16092 (N_16092,N_12956,N_14733);
or U16093 (N_16093,N_13578,N_13338);
nand U16094 (N_16094,N_14915,N_13498);
nand U16095 (N_16095,N_13904,N_14211);
and U16096 (N_16096,N_14315,N_12714);
nand U16097 (N_16097,N_14261,N_13320);
nand U16098 (N_16098,N_14128,N_14173);
nand U16099 (N_16099,N_13462,N_12664);
nand U16100 (N_16100,N_13508,N_14896);
and U16101 (N_16101,N_13158,N_13746);
nor U16102 (N_16102,N_12725,N_14807);
or U16103 (N_16103,N_13329,N_12912);
and U16104 (N_16104,N_13544,N_14492);
nor U16105 (N_16105,N_14217,N_14422);
nor U16106 (N_16106,N_14143,N_14918);
or U16107 (N_16107,N_14125,N_13187);
and U16108 (N_16108,N_12777,N_14250);
or U16109 (N_16109,N_14753,N_13759);
nor U16110 (N_16110,N_13717,N_12880);
or U16111 (N_16111,N_12575,N_14241);
nor U16112 (N_16112,N_12785,N_12824);
nor U16113 (N_16113,N_14881,N_14084);
xor U16114 (N_16114,N_14087,N_13077);
xor U16115 (N_16115,N_14524,N_13595);
nand U16116 (N_16116,N_13837,N_14032);
nand U16117 (N_16117,N_12510,N_14689);
and U16118 (N_16118,N_13523,N_13599);
nand U16119 (N_16119,N_14393,N_14723);
and U16120 (N_16120,N_12682,N_14312);
nand U16121 (N_16121,N_12621,N_13543);
or U16122 (N_16122,N_12918,N_14195);
nor U16123 (N_16123,N_13805,N_14240);
and U16124 (N_16124,N_13270,N_13025);
or U16125 (N_16125,N_12716,N_13023);
or U16126 (N_16126,N_14937,N_13716);
and U16127 (N_16127,N_13199,N_14840);
nor U16128 (N_16128,N_13255,N_12746);
nor U16129 (N_16129,N_12687,N_14762);
and U16130 (N_16130,N_13901,N_13309);
or U16131 (N_16131,N_14226,N_14290);
nor U16132 (N_16132,N_13713,N_12766);
or U16133 (N_16133,N_14509,N_14196);
nand U16134 (N_16134,N_14656,N_14600);
and U16135 (N_16135,N_14138,N_14269);
nor U16136 (N_16136,N_13557,N_14532);
or U16137 (N_16137,N_12984,N_12855);
and U16138 (N_16138,N_14351,N_12792);
nor U16139 (N_16139,N_14407,N_14494);
or U16140 (N_16140,N_13996,N_14330);
and U16141 (N_16141,N_13083,N_14481);
or U16142 (N_16142,N_13356,N_13825);
nor U16143 (N_16143,N_14907,N_14563);
nand U16144 (N_16144,N_14282,N_13708);
nand U16145 (N_16145,N_12886,N_12738);
nor U16146 (N_16146,N_14199,N_13920);
nand U16147 (N_16147,N_13285,N_12655);
nor U16148 (N_16148,N_14266,N_13313);
xor U16149 (N_16149,N_14848,N_13469);
or U16150 (N_16150,N_13176,N_13893);
and U16151 (N_16151,N_13760,N_12584);
nor U16152 (N_16152,N_13574,N_14668);
and U16153 (N_16153,N_12698,N_13722);
nor U16154 (N_16154,N_14507,N_13822);
and U16155 (N_16155,N_13019,N_13745);
nand U16156 (N_16156,N_14823,N_12911);
nor U16157 (N_16157,N_13161,N_14022);
nor U16158 (N_16158,N_12929,N_13879);
nor U16159 (N_16159,N_12870,N_14119);
nand U16160 (N_16160,N_13955,N_14664);
and U16161 (N_16161,N_13334,N_13293);
nand U16162 (N_16162,N_13186,N_14096);
nand U16163 (N_16163,N_13076,N_14650);
nor U16164 (N_16164,N_14832,N_14115);
and U16165 (N_16165,N_13388,N_13799);
nand U16166 (N_16166,N_14986,N_14463);
nor U16167 (N_16167,N_14639,N_13661);
xnor U16168 (N_16168,N_14073,N_12920);
and U16169 (N_16169,N_12894,N_13972);
nor U16170 (N_16170,N_12553,N_13339);
nand U16171 (N_16171,N_14268,N_13934);
nor U16172 (N_16172,N_13084,N_13548);
nand U16173 (N_16173,N_13969,N_12524);
nand U16174 (N_16174,N_14859,N_13736);
nor U16175 (N_16175,N_13787,N_14520);
xor U16176 (N_16176,N_14514,N_13912);
or U16177 (N_16177,N_12972,N_13374);
and U16178 (N_16178,N_13281,N_14670);
nand U16179 (N_16179,N_14074,N_13554);
and U16180 (N_16180,N_13376,N_13894);
nand U16181 (N_16181,N_13966,N_13473);
and U16182 (N_16182,N_13968,N_14491);
nand U16183 (N_16183,N_14678,N_12957);
or U16184 (N_16184,N_14497,N_13354);
nand U16185 (N_16185,N_14254,N_12843);
nand U16186 (N_16186,N_13676,N_13681);
nand U16187 (N_16187,N_12907,N_13027);
nand U16188 (N_16188,N_13289,N_13591);
or U16189 (N_16189,N_14829,N_14629);
nor U16190 (N_16190,N_12693,N_13145);
nor U16191 (N_16191,N_14616,N_12699);
nor U16192 (N_16192,N_12906,N_14416);
nand U16193 (N_16193,N_12679,N_12745);
or U16194 (N_16194,N_13020,N_13419);
xor U16195 (N_16195,N_13780,N_13323);
nor U16196 (N_16196,N_13262,N_12562);
nand U16197 (N_16197,N_14876,N_13434);
nor U16198 (N_16198,N_12790,N_13707);
and U16199 (N_16199,N_13146,N_13290);
or U16200 (N_16200,N_13819,N_12913);
or U16201 (N_16201,N_13367,N_14740);
and U16202 (N_16202,N_13511,N_13507);
or U16203 (N_16203,N_13539,N_12798);
nand U16204 (N_16204,N_13768,N_13679);
nand U16205 (N_16205,N_12783,N_14606);
and U16206 (N_16206,N_12681,N_14745);
or U16207 (N_16207,N_14797,N_14253);
or U16208 (N_16208,N_12839,N_12703);
or U16209 (N_16209,N_14359,N_13971);
nand U16210 (N_16210,N_14184,N_14536);
nor U16211 (N_16211,N_12864,N_14658);
nor U16212 (N_16212,N_14186,N_13602);
xor U16213 (N_16213,N_14181,N_14774);
nand U16214 (N_16214,N_12756,N_13940);
and U16215 (N_16215,N_12799,N_13336);
nand U16216 (N_16216,N_14680,N_13654);
nand U16217 (N_16217,N_13790,N_14540);
nor U16218 (N_16218,N_13392,N_14816);
or U16219 (N_16219,N_13862,N_14408);
xor U16220 (N_16220,N_12778,N_14321);
and U16221 (N_16221,N_12538,N_14353);
nand U16222 (N_16222,N_12819,N_13295);
nand U16223 (N_16223,N_14392,N_14769);
nor U16224 (N_16224,N_14127,N_13718);
nor U16225 (N_16225,N_13594,N_12941);
or U16226 (N_16226,N_14537,N_14770);
or U16227 (N_16227,N_13142,N_13531);
nand U16228 (N_16228,N_12684,N_12897);
or U16229 (N_16229,N_13445,N_14961);
nand U16230 (N_16230,N_14595,N_13455);
and U16231 (N_16231,N_13326,N_12733);
or U16232 (N_16232,N_14212,N_14051);
xor U16233 (N_16233,N_13737,N_14185);
xnor U16234 (N_16234,N_13773,N_12923);
nand U16235 (N_16235,N_14306,N_13723);
nand U16236 (N_16236,N_13995,N_13999);
nor U16237 (N_16237,N_14526,N_13613);
and U16238 (N_16238,N_12992,N_14811);
or U16239 (N_16239,N_13932,N_14317);
and U16240 (N_16240,N_12904,N_13060);
or U16241 (N_16241,N_13113,N_14662);
nand U16242 (N_16242,N_14231,N_13331);
nor U16243 (N_16243,N_14822,N_12966);
nor U16244 (N_16244,N_13288,N_12622);
nor U16245 (N_16245,N_14871,N_12977);
nor U16246 (N_16246,N_14767,N_12813);
and U16247 (N_16247,N_14842,N_13063);
nand U16248 (N_16248,N_13081,N_13086);
nor U16249 (N_16249,N_13316,N_13468);
nor U16250 (N_16250,N_14495,N_13252);
xor U16251 (N_16251,N_13375,N_13421);
nand U16252 (N_16252,N_12613,N_12864);
and U16253 (N_16253,N_12702,N_14857);
or U16254 (N_16254,N_14637,N_14260);
nand U16255 (N_16255,N_12647,N_12724);
and U16256 (N_16256,N_14079,N_13289);
nor U16257 (N_16257,N_13613,N_12731);
and U16258 (N_16258,N_14008,N_12602);
or U16259 (N_16259,N_13336,N_13593);
and U16260 (N_16260,N_13719,N_14888);
or U16261 (N_16261,N_14680,N_13208);
or U16262 (N_16262,N_14892,N_13101);
nor U16263 (N_16263,N_13166,N_14642);
nor U16264 (N_16264,N_14638,N_14610);
or U16265 (N_16265,N_13888,N_13322);
nor U16266 (N_16266,N_14199,N_14370);
nand U16267 (N_16267,N_14938,N_13126);
xnor U16268 (N_16268,N_13434,N_13823);
nor U16269 (N_16269,N_14789,N_14976);
or U16270 (N_16270,N_14222,N_13320);
nand U16271 (N_16271,N_14532,N_13307);
nand U16272 (N_16272,N_14478,N_13644);
nand U16273 (N_16273,N_14391,N_14849);
or U16274 (N_16274,N_13731,N_14716);
xor U16275 (N_16275,N_13817,N_12579);
or U16276 (N_16276,N_13139,N_14082);
or U16277 (N_16277,N_13489,N_14837);
or U16278 (N_16278,N_13994,N_13401);
or U16279 (N_16279,N_14257,N_13214);
or U16280 (N_16280,N_13367,N_14420);
nand U16281 (N_16281,N_13959,N_12911);
or U16282 (N_16282,N_14331,N_12773);
nand U16283 (N_16283,N_14520,N_12974);
nor U16284 (N_16284,N_14988,N_14416);
and U16285 (N_16285,N_14244,N_14261);
and U16286 (N_16286,N_13370,N_13375);
nand U16287 (N_16287,N_13641,N_14031);
and U16288 (N_16288,N_13259,N_12530);
nor U16289 (N_16289,N_14236,N_14064);
nor U16290 (N_16290,N_14981,N_13603);
and U16291 (N_16291,N_12778,N_14742);
nor U16292 (N_16292,N_14270,N_13643);
nor U16293 (N_16293,N_14336,N_13836);
or U16294 (N_16294,N_13443,N_13890);
and U16295 (N_16295,N_13375,N_14000);
or U16296 (N_16296,N_14878,N_14683);
or U16297 (N_16297,N_13498,N_12516);
nor U16298 (N_16298,N_12807,N_13490);
or U16299 (N_16299,N_14116,N_14035);
and U16300 (N_16300,N_13307,N_14977);
and U16301 (N_16301,N_14283,N_14156);
nor U16302 (N_16302,N_13174,N_12576);
and U16303 (N_16303,N_14282,N_14272);
and U16304 (N_16304,N_14831,N_14349);
nand U16305 (N_16305,N_14593,N_13877);
and U16306 (N_16306,N_14704,N_14422);
nor U16307 (N_16307,N_13082,N_14795);
and U16308 (N_16308,N_13700,N_14929);
nand U16309 (N_16309,N_12947,N_12925);
nor U16310 (N_16310,N_12736,N_14715);
nor U16311 (N_16311,N_13432,N_14137);
nor U16312 (N_16312,N_13565,N_13843);
or U16313 (N_16313,N_14963,N_13655);
or U16314 (N_16314,N_13314,N_12649);
or U16315 (N_16315,N_13301,N_14275);
nor U16316 (N_16316,N_14870,N_14204);
and U16317 (N_16317,N_14636,N_14652);
and U16318 (N_16318,N_13622,N_14725);
nor U16319 (N_16319,N_13027,N_14218);
or U16320 (N_16320,N_14292,N_13758);
and U16321 (N_16321,N_13458,N_13495);
nand U16322 (N_16322,N_14385,N_13660);
or U16323 (N_16323,N_14649,N_13001);
xnor U16324 (N_16324,N_14168,N_13108);
xnor U16325 (N_16325,N_12884,N_13514);
or U16326 (N_16326,N_12910,N_14871);
and U16327 (N_16327,N_12812,N_14715);
nor U16328 (N_16328,N_14195,N_13708);
or U16329 (N_16329,N_13778,N_13382);
or U16330 (N_16330,N_14254,N_13301);
and U16331 (N_16331,N_14858,N_12926);
or U16332 (N_16332,N_13854,N_13007);
nor U16333 (N_16333,N_13323,N_14125);
or U16334 (N_16334,N_12827,N_13218);
or U16335 (N_16335,N_13746,N_13573);
nor U16336 (N_16336,N_13448,N_12956);
or U16337 (N_16337,N_13078,N_14981);
nor U16338 (N_16338,N_12957,N_13160);
or U16339 (N_16339,N_12765,N_13013);
nor U16340 (N_16340,N_13912,N_14372);
nor U16341 (N_16341,N_13644,N_14379);
nand U16342 (N_16342,N_12735,N_13077);
and U16343 (N_16343,N_14477,N_13100);
or U16344 (N_16344,N_14302,N_14450);
and U16345 (N_16345,N_13451,N_14540);
and U16346 (N_16346,N_13219,N_14785);
nor U16347 (N_16347,N_12673,N_14259);
and U16348 (N_16348,N_13889,N_14328);
or U16349 (N_16349,N_14365,N_13058);
nor U16350 (N_16350,N_14134,N_14831);
nand U16351 (N_16351,N_14906,N_14606);
xnor U16352 (N_16352,N_13221,N_14292);
xor U16353 (N_16353,N_14427,N_12688);
xor U16354 (N_16354,N_14684,N_14433);
xnor U16355 (N_16355,N_13427,N_13802);
and U16356 (N_16356,N_14444,N_14936);
xnor U16357 (N_16357,N_14080,N_12722);
nor U16358 (N_16358,N_14619,N_14444);
or U16359 (N_16359,N_14004,N_13120);
or U16360 (N_16360,N_12606,N_13840);
xor U16361 (N_16361,N_13148,N_13798);
and U16362 (N_16362,N_14771,N_13181);
and U16363 (N_16363,N_12926,N_13828);
nor U16364 (N_16364,N_14190,N_13268);
and U16365 (N_16365,N_14384,N_13738);
and U16366 (N_16366,N_14644,N_13406);
nor U16367 (N_16367,N_13520,N_14765);
nor U16368 (N_16368,N_13687,N_13985);
nor U16369 (N_16369,N_14793,N_14833);
xor U16370 (N_16370,N_12930,N_14028);
and U16371 (N_16371,N_13076,N_13045);
and U16372 (N_16372,N_14208,N_12547);
nor U16373 (N_16373,N_12859,N_13966);
and U16374 (N_16374,N_13332,N_14642);
or U16375 (N_16375,N_13699,N_13447);
nand U16376 (N_16376,N_13333,N_13610);
or U16377 (N_16377,N_13890,N_13534);
nor U16378 (N_16378,N_14418,N_14526);
or U16379 (N_16379,N_13714,N_14845);
or U16380 (N_16380,N_14187,N_12658);
nor U16381 (N_16381,N_13751,N_14256);
or U16382 (N_16382,N_12984,N_13342);
and U16383 (N_16383,N_14611,N_13110);
nor U16384 (N_16384,N_13791,N_14470);
nand U16385 (N_16385,N_13386,N_13029);
or U16386 (N_16386,N_12845,N_14804);
or U16387 (N_16387,N_13960,N_14039);
nand U16388 (N_16388,N_13531,N_12681);
or U16389 (N_16389,N_13602,N_14447);
nor U16390 (N_16390,N_12534,N_13490);
nand U16391 (N_16391,N_14259,N_13423);
and U16392 (N_16392,N_14902,N_12557);
nand U16393 (N_16393,N_12951,N_13608);
or U16394 (N_16394,N_12983,N_14120);
and U16395 (N_16395,N_13216,N_14746);
or U16396 (N_16396,N_13476,N_12980);
nand U16397 (N_16397,N_14693,N_14781);
nand U16398 (N_16398,N_13973,N_14475);
nor U16399 (N_16399,N_12814,N_14668);
nor U16400 (N_16400,N_12636,N_13093);
xnor U16401 (N_16401,N_13104,N_13612);
nor U16402 (N_16402,N_14706,N_13038);
xor U16403 (N_16403,N_13799,N_14151);
nand U16404 (N_16404,N_14093,N_14383);
or U16405 (N_16405,N_13480,N_14888);
or U16406 (N_16406,N_14754,N_14133);
nor U16407 (N_16407,N_12608,N_14131);
and U16408 (N_16408,N_13923,N_12857);
xor U16409 (N_16409,N_14547,N_13118);
and U16410 (N_16410,N_13287,N_14315);
xor U16411 (N_16411,N_12996,N_14446);
nor U16412 (N_16412,N_13671,N_13069);
nand U16413 (N_16413,N_12975,N_12571);
or U16414 (N_16414,N_14675,N_13156);
nand U16415 (N_16415,N_14286,N_13188);
nand U16416 (N_16416,N_13645,N_13400);
nand U16417 (N_16417,N_14154,N_13286);
and U16418 (N_16418,N_12867,N_12808);
and U16419 (N_16419,N_13385,N_13059);
or U16420 (N_16420,N_12805,N_13381);
nor U16421 (N_16421,N_13661,N_14138);
or U16422 (N_16422,N_13552,N_13000);
nand U16423 (N_16423,N_13213,N_13791);
nor U16424 (N_16424,N_14467,N_14942);
xor U16425 (N_16425,N_12520,N_14978);
or U16426 (N_16426,N_12936,N_14331);
nor U16427 (N_16427,N_13094,N_13963);
xnor U16428 (N_16428,N_12543,N_13411);
or U16429 (N_16429,N_14905,N_14127);
and U16430 (N_16430,N_14652,N_13217);
and U16431 (N_16431,N_14901,N_14917);
or U16432 (N_16432,N_13757,N_14055);
nand U16433 (N_16433,N_14612,N_13249);
and U16434 (N_16434,N_12755,N_13335);
and U16435 (N_16435,N_14113,N_14595);
xor U16436 (N_16436,N_13909,N_14950);
and U16437 (N_16437,N_13000,N_13323);
and U16438 (N_16438,N_14928,N_12949);
nand U16439 (N_16439,N_12799,N_14130);
nand U16440 (N_16440,N_14449,N_14000);
nand U16441 (N_16441,N_13894,N_14804);
nor U16442 (N_16442,N_12534,N_14183);
and U16443 (N_16443,N_14347,N_13276);
nand U16444 (N_16444,N_12949,N_13769);
nand U16445 (N_16445,N_12907,N_13329);
nor U16446 (N_16446,N_14293,N_14988);
nand U16447 (N_16447,N_13075,N_13960);
and U16448 (N_16448,N_14678,N_14722);
xnor U16449 (N_16449,N_13080,N_14814);
and U16450 (N_16450,N_14811,N_12565);
nand U16451 (N_16451,N_14764,N_14756);
xnor U16452 (N_16452,N_13545,N_14166);
and U16453 (N_16453,N_13351,N_14625);
or U16454 (N_16454,N_14128,N_14325);
and U16455 (N_16455,N_14514,N_13255);
or U16456 (N_16456,N_12903,N_12936);
nand U16457 (N_16457,N_13836,N_14527);
nor U16458 (N_16458,N_14480,N_13714);
nor U16459 (N_16459,N_14220,N_14741);
nand U16460 (N_16460,N_14363,N_13115);
and U16461 (N_16461,N_12633,N_14337);
xnor U16462 (N_16462,N_14619,N_13169);
and U16463 (N_16463,N_13691,N_13281);
and U16464 (N_16464,N_14315,N_12949);
nor U16465 (N_16465,N_14566,N_13459);
nor U16466 (N_16466,N_13412,N_12649);
or U16467 (N_16467,N_12962,N_13082);
and U16468 (N_16468,N_14483,N_14215);
nand U16469 (N_16469,N_12634,N_13352);
or U16470 (N_16470,N_13727,N_14711);
and U16471 (N_16471,N_13121,N_14543);
nand U16472 (N_16472,N_14395,N_14074);
or U16473 (N_16473,N_13407,N_13180);
nor U16474 (N_16474,N_12850,N_12787);
and U16475 (N_16475,N_14287,N_13655);
nand U16476 (N_16476,N_12634,N_13520);
nor U16477 (N_16477,N_12816,N_12736);
or U16478 (N_16478,N_13076,N_14626);
or U16479 (N_16479,N_14982,N_13698);
or U16480 (N_16480,N_13078,N_14148);
xnor U16481 (N_16481,N_12937,N_14086);
nand U16482 (N_16482,N_13856,N_13614);
xnor U16483 (N_16483,N_12942,N_14263);
or U16484 (N_16484,N_14988,N_12873);
nor U16485 (N_16485,N_13944,N_13018);
and U16486 (N_16486,N_13178,N_14999);
nor U16487 (N_16487,N_13240,N_14418);
or U16488 (N_16488,N_14035,N_12564);
nor U16489 (N_16489,N_14074,N_14088);
nor U16490 (N_16490,N_13315,N_14889);
nor U16491 (N_16491,N_13122,N_14404);
and U16492 (N_16492,N_12752,N_14829);
and U16493 (N_16493,N_12855,N_13552);
or U16494 (N_16494,N_14880,N_12960);
or U16495 (N_16495,N_13233,N_12804);
nor U16496 (N_16496,N_14016,N_14654);
nand U16497 (N_16497,N_13970,N_14714);
xor U16498 (N_16498,N_14782,N_13769);
or U16499 (N_16499,N_13820,N_13956);
or U16500 (N_16500,N_13211,N_14377);
nand U16501 (N_16501,N_13058,N_13592);
xnor U16502 (N_16502,N_12744,N_13684);
and U16503 (N_16503,N_14703,N_13194);
and U16504 (N_16504,N_12788,N_14013);
nor U16505 (N_16505,N_13213,N_14162);
or U16506 (N_16506,N_14518,N_12751);
or U16507 (N_16507,N_13199,N_12782);
and U16508 (N_16508,N_13222,N_14203);
and U16509 (N_16509,N_14073,N_12835);
nor U16510 (N_16510,N_13870,N_13068);
nor U16511 (N_16511,N_12754,N_14779);
nor U16512 (N_16512,N_12824,N_14904);
nor U16513 (N_16513,N_12971,N_13804);
and U16514 (N_16514,N_13535,N_13410);
and U16515 (N_16515,N_14878,N_13340);
nor U16516 (N_16516,N_14546,N_13043);
or U16517 (N_16517,N_13894,N_13993);
nand U16518 (N_16518,N_12570,N_13785);
nor U16519 (N_16519,N_13658,N_13380);
nor U16520 (N_16520,N_13074,N_14891);
nand U16521 (N_16521,N_12919,N_13038);
or U16522 (N_16522,N_13144,N_13303);
or U16523 (N_16523,N_13536,N_13236);
nand U16524 (N_16524,N_13115,N_14350);
nor U16525 (N_16525,N_13043,N_12590);
nand U16526 (N_16526,N_13003,N_14522);
nand U16527 (N_16527,N_12820,N_13156);
and U16528 (N_16528,N_12782,N_14948);
and U16529 (N_16529,N_13488,N_14627);
xnor U16530 (N_16530,N_14162,N_13200);
nand U16531 (N_16531,N_13010,N_14052);
nor U16532 (N_16532,N_13052,N_13600);
nor U16533 (N_16533,N_13415,N_13584);
nor U16534 (N_16534,N_14212,N_14688);
or U16535 (N_16535,N_13726,N_13978);
or U16536 (N_16536,N_12932,N_13139);
and U16537 (N_16537,N_14929,N_13301);
and U16538 (N_16538,N_14443,N_14913);
nor U16539 (N_16539,N_13688,N_13083);
or U16540 (N_16540,N_13336,N_13539);
xor U16541 (N_16541,N_13368,N_13187);
nor U16542 (N_16542,N_14442,N_13301);
nor U16543 (N_16543,N_12943,N_14217);
nor U16544 (N_16544,N_13147,N_13563);
xnor U16545 (N_16545,N_13246,N_13884);
and U16546 (N_16546,N_14531,N_14669);
and U16547 (N_16547,N_13213,N_14226);
nor U16548 (N_16548,N_14854,N_13573);
nor U16549 (N_16549,N_13454,N_12644);
nand U16550 (N_16550,N_14688,N_14981);
nor U16551 (N_16551,N_14726,N_13127);
nand U16552 (N_16552,N_14696,N_14424);
nor U16553 (N_16553,N_13030,N_14762);
nor U16554 (N_16554,N_13393,N_14229);
and U16555 (N_16555,N_14906,N_12807);
nor U16556 (N_16556,N_13922,N_14454);
nor U16557 (N_16557,N_12746,N_13912);
nand U16558 (N_16558,N_14373,N_14910);
nand U16559 (N_16559,N_12799,N_14451);
and U16560 (N_16560,N_14364,N_12639);
xor U16561 (N_16561,N_13324,N_13446);
nor U16562 (N_16562,N_13059,N_14732);
nor U16563 (N_16563,N_13661,N_14517);
nor U16564 (N_16564,N_12888,N_13289);
and U16565 (N_16565,N_14216,N_13631);
or U16566 (N_16566,N_12605,N_13381);
xor U16567 (N_16567,N_14919,N_12947);
nand U16568 (N_16568,N_13865,N_13768);
nand U16569 (N_16569,N_14826,N_14439);
nand U16570 (N_16570,N_14183,N_14253);
and U16571 (N_16571,N_13364,N_13766);
nand U16572 (N_16572,N_14913,N_14005);
nor U16573 (N_16573,N_13061,N_12811);
nand U16574 (N_16574,N_13790,N_13335);
and U16575 (N_16575,N_13739,N_12864);
and U16576 (N_16576,N_12980,N_14001);
xnor U16577 (N_16577,N_14406,N_13740);
or U16578 (N_16578,N_14481,N_14376);
nor U16579 (N_16579,N_12565,N_14465);
nor U16580 (N_16580,N_12701,N_13410);
nand U16581 (N_16581,N_14993,N_14985);
or U16582 (N_16582,N_14004,N_13628);
nor U16583 (N_16583,N_14599,N_14395);
or U16584 (N_16584,N_12886,N_13501);
nor U16585 (N_16585,N_14819,N_14575);
and U16586 (N_16586,N_14297,N_14784);
nand U16587 (N_16587,N_12540,N_13844);
and U16588 (N_16588,N_13497,N_12805);
or U16589 (N_16589,N_13640,N_13812);
nor U16590 (N_16590,N_14724,N_12562);
or U16591 (N_16591,N_13594,N_13303);
and U16592 (N_16592,N_13946,N_12838);
nand U16593 (N_16593,N_13880,N_13451);
or U16594 (N_16594,N_14241,N_12712);
nor U16595 (N_16595,N_14415,N_13117);
nor U16596 (N_16596,N_13531,N_13123);
and U16597 (N_16597,N_14123,N_13988);
or U16598 (N_16598,N_13652,N_13895);
nor U16599 (N_16599,N_13364,N_13019);
nor U16600 (N_16600,N_14964,N_14824);
and U16601 (N_16601,N_13281,N_14637);
or U16602 (N_16602,N_14356,N_13618);
and U16603 (N_16603,N_12740,N_13505);
or U16604 (N_16604,N_14562,N_14558);
xor U16605 (N_16605,N_13501,N_14124);
and U16606 (N_16606,N_13572,N_13236);
nor U16607 (N_16607,N_14580,N_14862);
nor U16608 (N_16608,N_12892,N_14911);
xor U16609 (N_16609,N_12827,N_14462);
and U16610 (N_16610,N_13535,N_14015);
nor U16611 (N_16611,N_14436,N_14982);
nor U16612 (N_16612,N_12909,N_14354);
nor U16613 (N_16613,N_13991,N_14418);
nor U16614 (N_16614,N_13069,N_12966);
nor U16615 (N_16615,N_13214,N_14147);
nand U16616 (N_16616,N_12661,N_13593);
or U16617 (N_16617,N_14925,N_13082);
nand U16618 (N_16618,N_14355,N_12585);
or U16619 (N_16619,N_14662,N_14241);
xnor U16620 (N_16620,N_13485,N_13041);
or U16621 (N_16621,N_12791,N_12607);
nor U16622 (N_16622,N_13392,N_13198);
nand U16623 (N_16623,N_13329,N_14676);
or U16624 (N_16624,N_14732,N_13573);
and U16625 (N_16625,N_14186,N_12691);
and U16626 (N_16626,N_12838,N_13386);
nand U16627 (N_16627,N_14978,N_13329);
and U16628 (N_16628,N_13955,N_14117);
nor U16629 (N_16629,N_14066,N_13444);
nand U16630 (N_16630,N_13310,N_13223);
or U16631 (N_16631,N_12980,N_14407);
xor U16632 (N_16632,N_13301,N_14093);
and U16633 (N_16633,N_13531,N_13609);
or U16634 (N_16634,N_12755,N_14655);
nor U16635 (N_16635,N_14042,N_13769);
nor U16636 (N_16636,N_13888,N_12554);
and U16637 (N_16637,N_14452,N_14990);
and U16638 (N_16638,N_14776,N_14167);
and U16639 (N_16639,N_14521,N_12556);
or U16640 (N_16640,N_14021,N_14891);
nor U16641 (N_16641,N_13204,N_13893);
nor U16642 (N_16642,N_12770,N_13194);
or U16643 (N_16643,N_13178,N_13640);
or U16644 (N_16644,N_13792,N_13632);
nand U16645 (N_16645,N_13174,N_13459);
or U16646 (N_16646,N_13020,N_13547);
or U16647 (N_16647,N_12889,N_14207);
and U16648 (N_16648,N_13954,N_13505);
and U16649 (N_16649,N_14355,N_14211);
nor U16650 (N_16650,N_13353,N_13072);
or U16651 (N_16651,N_13167,N_14427);
xnor U16652 (N_16652,N_13788,N_13937);
nand U16653 (N_16653,N_14589,N_13319);
and U16654 (N_16654,N_14144,N_12577);
nor U16655 (N_16655,N_13888,N_14115);
xnor U16656 (N_16656,N_14837,N_13313);
and U16657 (N_16657,N_13922,N_13061);
and U16658 (N_16658,N_14022,N_14131);
or U16659 (N_16659,N_14972,N_13553);
xor U16660 (N_16660,N_14912,N_14099);
nor U16661 (N_16661,N_12957,N_14496);
and U16662 (N_16662,N_14065,N_14643);
nand U16663 (N_16663,N_13050,N_12899);
or U16664 (N_16664,N_13194,N_12558);
and U16665 (N_16665,N_12907,N_14644);
or U16666 (N_16666,N_13869,N_12640);
or U16667 (N_16667,N_14963,N_12915);
and U16668 (N_16668,N_13127,N_12586);
nor U16669 (N_16669,N_14563,N_13993);
or U16670 (N_16670,N_13478,N_12628);
xor U16671 (N_16671,N_14774,N_13544);
or U16672 (N_16672,N_12842,N_13389);
and U16673 (N_16673,N_14178,N_14581);
nor U16674 (N_16674,N_14357,N_13292);
xnor U16675 (N_16675,N_14405,N_12856);
and U16676 (N_16676,N_12719,N_13741);
or U16677 (N_16677,N_13981,N_14857);
nand U16678 (N_16678,N_14163,N_14101);
nand U16679 (N_16679,N_14643,N_13874);
nor U16680 (N_16680,N_14527,N_12534);
nand U16681 (N_16681,N_14568,N_13454);
nor U16682 (N_16682,N_13060,N_13320);
xnor U16683 (N_16683,N_13630,N_14450);
or U16684 (N_16684,N_12908,N_14424);
nand U16685 (N_16685,N_13588,N_14935);
or U16686 (N_16686,N_14980,N_12744);
nand U16687 (N_16687,N_14932,N_12728);
and U16688 (N_16688,N_12823,N_12865);
nor U16689 (N_16689,N_12819,N_13871);
nand U16690 (N_16690,N_13721,N_14498);
or U16691 (N_16691,N_14127,N_13551);
nand U16692 (N_16692,N_13399,N_13224);
and U16693 (N_16693,N_14527,N_12576);
xnor U16694 (N_16694,N_14499,N_14809);
or U16695 (N_16695,N_14676,N_14837);
xor U16696 (N_16696,N_14612,N_14961);
or U16697 (N_16697,N_13943,N_13712);
or U16698 (N_16698,N_13333,N_12783);
nor U16699 (N_16699,N_14008,N_13803);
and U16700 (N_16700,N_14115,N_14072);
xnor U16701 (N_16701,N_13026,N_14242);
nor U16702 (N_16702,N_12879,N_12959);
nor U16703 (N_16703,N_12981,N_14229);
or U16704 (N_16704,N_12684,N_13175);
or U16705 (N_16705,N_12851,N_14280);
or U16706 (N_16706,N_14140,N_14742);
or U16707 (N_16707,N_13736,N_13082);
nor U16708 (N_16708,N_12652,N_14900);
xor U16709 (N_16709,N_14103,N_14977);
nand U16710 (N_16710,N_13624,N_13081);
nor U16711 (N_16711,N_13702,N_12548);
and U16712 (N_16712,N_13468,N_14450);
nor U16713 (N_16713,N_13892,N_12900);
and U16714 (N_16714,N_14782,N_12942);
or U16715 (N_16715,N_14476,N_12857);
and U16716 (N_16716,N_13849,N_13801);
nor U16717 (N_16717,N_13365,N_14529);
nand U16718 (N_16718,N_12618,N_12550);
nand U16719 (N_16719,N_13551,N_13419);
or U16720 (N_16720,N_12825,N_14493);
and U16721 (N_16721,N_14697,N_12572);
nor U16722 (N_16722,N_12649,N_14417);
or U16723 (N_16723,N_14381,N_14306);
nor U16724 (N_16724,N_12931,N_13572);
or U16725 (N_16725,N_12838,N_13926);
or U16726 (N_16726,N_14058,N_13031);
or U16727 (N_16727,N_13153,N_13082);
and U16728 (N_16728,N_14721,N_13049);
nor U16729 (N_16729,N_12732,N_12829);
nor U16730 (N_16730,N_14646,N_14056);
nor U16731 (N_16731,N_12698,N_14965);
or U16732 (N_16732,N_14561,N_13164);
nor U16733 (N_16733,N_13471,N_14580);
nand U16734 (N_16734,N_12818,N_12865);
nand U16735 (N_16735,N_14577,N_13630);
and U16736 (N_16736,N_14230,N_14759);
or U16737 (N_16737,N_14165,N_13331);
nor U16738 (N_16738,N_14434,N_13956);
nand U16739 (N_16739,N_12931,N_14475);
nand U16740 (N_16740,N_14107,N_14574);
nand U16741 (N_16741,N_12590,N_13096);
nand U16742 (N_16742,N_14641,N_14225);
nor U16743 (N_16743,N_12657,N_14802);
nor U16744 (N_16744,N_14490,N_12974);
xnor U16745 (N_16745,N_13850,N_13013);
or U16746 (N_16746,N_13972,N_13817);
and U16747 (N_16747,N_13807,N_14922);
nand U16748 (N_16748,N_13261,N_14273);
nor U16749 (N_16749,N_13616,N_13020);
and U16750 (N_16750,N_13479,N_14582);
nand U16751 (N_16751,N_12793,N_14403);
nand U16752 (N_16752,N_13014,N_14713);
nand U16753 (N_16753,N_13146,N_14543);
xor U16754 (N_16754,N_13990,N_14216);
and U16755 (N_16755,N_14491,N_14767);
or U16756 (N_16756,N_12887,N_13060);
nand U16757 (N_16757,N_14729,N_13227);
and U16758 (N_16758,N_13335,N_14037);
nor U16759 (N_16759,N_14108,N_13303);
nor U16760 (N_16760,N_14551,N_13373);
or U16761 (N_16761,N_13746,N_12656);
and U16762 (N_16762,N_13226,N_13002);
nand U16763 (N_16763,N_12937,N_12672);
nand U16764 (N_16764,N_14323,N_14058);
nand U16765 (N_16765,N_13941,N_12729);
or U16766 (N_16766,N_14677,N_13237);
nor U16767 (N_16767,N_14891,N_13859);
or U16768 (N_16768,N_14730,N_14212);
nor U16769 (N_16769,N_13429,N_12717);
and U16770 (N_16770,N_13251,N_14042);
nand U16771 (N_16771,N_12570,N_13956);
or U16772 (N_16772,N_12752,N_13118);
xnor U16773 (N_16773,N_13618,N_13729);
and U16774 (N_16774,N_12834,N_13851);
nor U16775 (N_16775,N_14680,N_13173);
or U16776 (N_16776,N_14334,N_14240);
nand U16777 (N_16777,N_12765,N_14445);
or U16778 (N_16778,N_13111,N_14244);
nand U16779 (N_16779,N_12999,N_14201);
nand U16780 (N_16780,N_14285,N_12539);
nor U16781 (N_16781,N_14546,N_14669);
or U16782 (N_16782,N_14617,N_13096);
and U16783 (N_16783,N_12707,N_13543);
and U16784 (N_16784,N_14404,N_14063);
or U16785 (N_16785,N_14663,N_13217);
and U16786 (N_16786,N_14252,N_14759);
and U16787 (N_16787,N_13694,N_14022);
nand U16788 (N_16788,N_13220,N_12916);
nand U16789 (N_16789,N_13308,N_12800);
nor U16790 (N_16790,N_12841,N_14390);
nor U16791 (N_16791,N_14175,N_13291);
nor U16792 (N_16792,N_14533,N_13375);
nor U16793 (N_16793,N_14344,N_14512);
or U16794 (N_16794,N_13792,N_13887);
nor U16795 (N_16795,N_12701,N_12820);
nand U16796 (N_16796,N_14547,N_13514);
and U16797 (N_16797,N_13930,N_13126);
nor U16798 (N_16798,N_13227,N_12974);
or U16799 (N_16799,N_13692,N_12663);
and U16800 (N_16800,N_13421,N_12687);
xnor U16801 (N_16801,N_14575,N_12833);
xnor U16802 (N_16802,N_12589,N_13792);
nor U16803 (N_16803,N_13648,N_13794);
nor U16804 (N_16804,N_12788,N_12989);
nand U16805 (N_16805,N_13157,N_13933);
or U16806 (N_16806,N_14066,N_14619);
nor U16807 (N_16807,N_13624,N_13940);
nand U16808 (N_16808,N_12968,N_14404);
nand U16809 (N_16809,N_14030,N_12760);
and U16810 (N_16810,N_12942,N_14803);
nand U16811 (N_16811,N_14570,N_14216);
xnor U16812 (N_16812,N_14454,N_14011);
nor U16813 (N_16813,N_14529,N_12916);
nor U16814 (N_16814,N_14965,N_14486);
and U16815 (N_16815,N_13005,N_13562);
or U16816 (N_16816,N_14267,N_13640);
or U16817 (N_16817,N_13600,N_13796);
nor U16818 (N_16818,N_14675,N_14697);
xnor U16819 (N_16819,N_14888,N_13553);
nand U16820 (N_16820,N_13447,N_12690);
and U16821 (N_16821,N_14302,N_12641);
nand U16822 (N_16822,N_14846,N_14667);
nand U16823 (N_16823,N_14533,N_13008);
nand U16824 (N_16824,N_12999,N_13163);
nor U16825 (N_16825,N_13952,N_13845);
xnor U16826 (N_16826,N_14475,N_13433);
nand U16827 (N_16827,N_14634,N_13912);
and U16828 (N_16828,N_14979,N_14811);
and U16829 (N_16829,N_14331,N_12536);
nor U16830 (N_16830,N_14975,N_13436);
and U16831 (N_16831,N_14748,N_13601);
and U16832 (N_16832,N_13645,N_13205);
or U16833 (N_16833,N_14732,N_12755);
nor U16834 (N_16834,N_12839,N_12633);
nand U16835 (N_16835,N_13009,N_14895);
nor U16836 (N_16836,N_14255,N_13537);
and U16837 (N_16837,N_13184,N_13209);
nand U16838 (N_16838,N_13464,N_14367);
nand U16839 (N_16839,N_13633,N_14632);
and U16840 (N_16840,N_13391,N_12602);
and U16841 (N_16841,N_12783,N_14106);
or U16842 (N_16842,N_13898,N_14673);
nand U16843 (N_16843,N_13969,N_14169);
and U16844 (N_16844,N_14810,N_13948);
or U16845 (N_16845,N_12822,N_14755);
xnor U16846 (N_16846,N_12664,N_13788);
or U16847 (N_16847,N_14772,N_13582);
or U16848 (N_16848,N_12941,N_13319);
nand U16849 (N_16849,N_14694,N_14073);
and U16850 (N_16850,N_13032,N_13353);
and U16851 (N_16851,N_12599,N_12801);
nand U16852 (N_16852,N_14452,N_13089);
nand U16853 (N_16853,N_12978,N_13834);
nor U16854 (N_16854,N_12608,N_13555);
or U16855 (N_16855,N_12618,N_13185);
or U16856 (N_16856,N_14842,N_14343);
or U16857 (N_16857,N_14773,N_14046);
nor U16858 (N_16858,N_12566,N_12887);
or U16859 (N_16859,N_14160,N_12670);
nor U16860 (N_16860,N_12992,N_13619);
and U16861 (N_16861,N_14407,N_13405);
nand U16862 (N_16862,N_14894,N_12898);
nor U16863 (N_16863,N_13099,N_14829);
nor U16864 (N_16864,N_13342,N_12598);
xor U16865 (N_16865,N_14038,N_14857);
or U16866 (N_16866,N_14781,N_14643);
nand U16867 (N_16867,N_12919,N_13886);
nor U16868 (N_16868,N_14289,N_14078);
or U16869 (N_16869,N_13547,N_14015);
nand U16870 (N_16870,N_13445,N_14071);
and U16871 (N_16871,N_12526,N_14146);
or U16872 (N_16872,N_13042,N_12947);
nand U16873 (N_16873,N_14713,N_14159);
and U16874 (N_16874,N_13927,N_12952);
or U16875 (N_16875,N_12987,N_14966);
nand U16876 (N_16876,N_13770,N_14612);
or U16877 (N_16877,N_14119,N_13554);
nor U16878 (N_16878,N_14522,N_12836);
nor U16879 (N_16879,N_14325,N_12835);
or U16880 (N_16880,N_13789,N_12807);
nor U16881 (N_16881,N_12579,N_13079);
nand U16882 (N_16882,N_12979,N_12807);
nor U16883 (N_16883,N_13149,N_14829);
and U16884 (N_16884,N_12654,N_14760);
or U16885 (N_16885,N_14312,N_14452);
or U16886 (N_16886,N_14947,N_13034);
or U16887 (N_16887,N_13423,N_13350);
nor U16888 (N_16888,N_14730,N_13161);
and U16889 (N_16889,N_13366,N_13083);
nor U16890 (N_16890,N_14285,N_14664);
nand U16891 (N_16891,N_12834,N_13615);
or U16892 (N_16892,N_12598,N_14386);
nor U16893 (N_16893,N_13198,N_13277);
and U16894 (N_16894,N_12570,N_14491);
or U16895 (N_16895,N_13933,N_14666);
nand U16896 (N_16896,N_14306,N_12963);
and U16897 (N_16897,N_12632,N_13232);
and U16898 (N_16898,N_12970,N_13138);
or U16899 (N_16899,N_12596,N_13788);
xor U16900 (N_16900,N_14459,N_14776);
nor U16901 (N_16901,N_14428,N_14022);
nand U16902 (N_16902,N_14637,N_14158);
nor U16903 (N_16903,N_13889,N_14777);
and U16904 (N_16904,N_13458,N_13630);
and U16905 (N_16905,N_13980,N_13849);
or U16906 (N_16906,N_12698,N_12538);
nor U16907 (N_16907,N_14990,N_12890);
and U16908 (N_16908,N_13397,N_14741);
and U16909 (N_16909,N_13107,N_13849);
nor U16910 (N_16910,N_13844,N_13184);
and U16911 (N_16911,N_14329,N_14961);
nand U16912 (N_16912,N_14503,N_14558);
nor U16913 (N_16913,N_13345,N_13363);
nand U16914 (N_16914,N_14873,N_13866);
xor U16915 (N_16915,N_13010,N_13860);
or U16916 (N_16916,N_13577,N_14747);
xor U16917 (N_16917,N_12533,N_12764);
and U16918 (N_16918,N_14162,N_13456);
nand U16919 (N_16919,N_12841,N_14803);
nor U16920 (N_16920,N_14942,N_14005);
xor U16921 (N_16921,N_14110,N_12806);
and U16922 (N_16922,N_13637,N_12921);
or U16923 (N_16923,N_14164,N_14822);
nand U16924 (N_16924,N_12548,N_14503);
or U16925 (N_16925,N_14801,N_13333);
nand U16926 (N_16926,N_13658,N_13281);
and U16927 (N_16927,N_14101,N_12744);
or U16928 (N_16928,N_12639,N_13569);
or U16929 (N_16929,N_12516,N_14428);
nor U16930 (N_16930,N_14376,N_14854);
nand U16931 (N_16931,N_14924,N_13668);
nor U16932 (N_16932,N_13352,N_14232);
nand U16933 (N_16933,N_14372,N_14542);
xnor U16934 (N_16934,N_14038,N_12928);
nand U16935 (N_16935,N_14404,N_13323);
xor U16936 (N_16936,N_13200,N_14499);
nor U16937 (N_16937,N_14427,N_13858);
and U16938 (N_16938,N_12923,N_14715);
and U16939 (N_16939,N_13706,N_14573);
nand U16940 (N_16940,N_14453,N_12733);
and U16941 (N_16941,N_12858,N_13663);
nor U16942 (N_16942,N_14776,N_13097);
and U16943 (N_16943,N_14939,N_14498);
or U16944 (N_16944,N_14780,N_14256);
or U16945 (N_16945,N_13340,N_12603);
or U16946 (N_16946,N_14176,N_14499);
and U16947 (N_16947,N_14713,N_14340);
or U16948 (N_16948,N_13544,N_13438);
and U16949 (N_16949,N_14572,N_14490);
nor U16950 (N_16950,N_12670,N_12894);
and U16951 (N_16951,N_12917,N_14327);
or U16952 (N_16952,N_14946,N_13434);
nor U16953 (N_16953,N_12940,N_13685);
nor U16954 (N_16954,N_13903,N_13026);
xnor U16955 (N_16955,N_12896,N_13816);
or U16956 (N_16956,N_14262,N_14711);
or U16957 (N_16957,N_14385,N_12606);
and U16958 (N_16958,N_14669,N_14914);
and U16959 (N_16959,N_13183,N_13413);
xor U16960 (N_16960,N_14054,N_13072);
nand U16961 (N_16961,N_12608,N_13605);
or U16962 (N_16962,N_14084,N_14075);
nor U16963 (N_16963,N_14024,N_14722);
or U16964 (N_16964,N_12786,N_14890);
nor U16965 (N_16965,N_14558,N_13769);
or U16966 (N_16966,N_14629,N_13858);
or U16967 (N_16967,N_13676,N_14057);
or U16968 (N_16968,N_12713,N_12951);
nand U16969 (N_16969,N_12890,N_14975);
nor U16970 (N_16970,N_12620,N_14774);
nand U16971 (N_16971,N_13584,N_14694);
or U16972 (N_16972,N_14237,N_14215);
and U16973 (N_16973,N_12601,N_14077);
xnor U16974 (N_16974,N_13477,N_13777);
and U16975 (N_16975,N_12867,N_13159);
nor U16976 (N_16976,N_14122,N_13477);
nand U16977 (N_16977,N_13290,N_13148);
nand U16978 (N_16978,N_13853,N_14883);
or U16979 (N_16979,N_13000,N_12674);
nand U16980 (N_16980,N_14485,N_12813);
or U16981 (N_16981,N_12891,N_13081);
nand U16982 (N_16982,N_13811,N_12826);
nor U16983 (N_16983,N_12909,N_14019);
nand U16984 (N_16984,N_13861,N_14135);
or U16985 (N_16985,N_13785,N_13303);
nand U16986 (N_16986,N_14514,N_12808);
and U16987 (N_16987,N_13200,N_12890);
or U16988 (N_16988,N_14195,N_13674);
nand U16989 (N_16989,N_12829,N_13137);
nand U16990 (N_16990,N_14458,N_14537);
nand U16991 (N_16991,N_13933,N_13421);
xor U16992 (N_16992,N_14041,N_13789);
nand U16993 (N_16993,N_14812,N_14714);
or U16994 (N_16994,N_12903,N_12782);
nand U16995 (N_16995,N_13928,N_14635);
and U16996 (N_16996,N_12829,N_13856);
and U16997 (N_16997,N_14503,N_14190);
nand U16998 (N_16998,N_13910,N_12632);
or U16999 (N_16999,N_13003,N_12649);
nor U17000 (N_17000,N_13664,N_13519);
nand U17001 (N_17001,N_12829,N_14186);
nand U17002 (N_17002,N_13529,N_12530);
nor U17003 (N_17003,N_13415,N_12524);
nor U17004 (N_17004,N_14274,N_12954);
and U17005 (N_17005,N_13500,N_14479);
nor U17006 (N_17006,N_13544,N_14929);
nand U17007 (N_17007,N_14542,N_12943);
nor U17008 (N_17008,N_12750,N_13376);
nand U17009 (N_17009,N_13612,N_14073);
or U17010 (N_17010,N_14351,N_12816);
nor U17011 (N_17011,N_13474,N_14002);
or U17012 (N_17012,N_14657,N_14488);
nor U17013 (N_17013,N_13049,N_14661);
nor U17014 (N_17014,N_14421,N_13017);
nand U17015 (N_17015,N_12793,N_14248);
nor U17016 (N_17016,N_13979,N_13051);
nand U17017 (N_17017,N_12804,N_14251);
nand U17018 (N_17018,N_13891,N_13380);
nand U17019 (N_17019,N_12784,N_13367);
xnor U17020 (N_17020,N_13418,N_13670);
or U17021 (N_17021,N_14574,N_13471);
or U17022 (N_17022,N_13870,N_14836);
nand U17023 (N_17023,N_12669,N_14365);
nand U17024 (N_17024,N_12870,N_14799);
nor U17025 (N_17025,N_14520,N_14013);
or U17026 (N_17026,N_13622,N_12500);
nand U17027 (N_17027,N_14527,N_13704);
nand U17028 (N_17028,N_14081,N_14863);
or U17029 (N_17029,N_13734,N_12704);
nand U17030 (N_17030,N_12539,N_14595);
nor U17031 (N_17031,N_12663,N_13728);
nand U17032 (N_17032,N_14839,N_13904);
nor U17033 (N_17033,N_13529,N_14273);
nand U17034 (N_17034,N_13220,N_14887);
or U17035 (N_17035,N_13363,N_13036);
and U17036 (N_17036,N_13625,N_13373);
and U17037 (N_17037,N_12988,N_13884);
nor U17038 (N_17038,N_13299,N_14644);
xnor U17039 (N_17039,N_12728,N_13212);
nand U17040 (N_17040,N_13604,N_13705);
or U17041 (N_17041,N_12713,N_12828);
nor U17042 (N_17042,N_13600,N_13650);
xnor U17043 (N_17043,N_14197,N_13216);
nor U17044 (N_17044,N_14720,N_12793);
and U17045 (N_17045,N_14979,N_14149);
or U17046 (N_17046,N_12974,N_14238);
or U17047 (N_17047,N_13872,N_14432);
nor U17048 (N_17048,N_14002,N_13643);
nor U17049 (N_17049,N_14287,N_14010);
nor U17050 (N_17050,N_14485,N_14562);
nand U17051 (N_17051,N_14315,N_13167);
xnor U17052 (N_17052,N_12641,N_14416);
or U17053 (N_17053,N_14933,N_14645);
nor U17054 (N_17054,N_14737,N_12577);
and U17055 (N_17055,N_14495,N_12629);
and U17056 (N_17056,N_13268,N_12603);
or U17057 (N_17057,N_14759,N_12737);
and U17058 (N_17058,N_13850,N_13933);
or U17059 (N_17059,N_13453,N_14415);
nand U17060 (N_17060,N_13177,N_12520);
and U17061 (N_17061,N_13053,N_14061);
or U17062 (N_17062,N_13202,N_13908);
or U17063 (N_17063,N_14948,N_14414);
nand U17064 (N_17064,N_13643,N_13225);
nor U17065 (N_17065,N_14161,N_13668);
and U17066 (N_17066,N_14464,N_14773);
and U17067 (N_17067,N_14103,N_12743);
nand U17068 (N_17068,N_13215,N_12592);
and U17069 (N_17069,N_14700,N_14293);
nand U17070 (N_17070,N_14209,N_12652);
nand U17071 (N_17071,N_13135,N_13205);
or U17072 (N_17072,N_12549,N_13912);
and U17073 (N_17073,N_14290,N_14919);
or U17074 (N_17074,N_14732,N_14400);
xnor U17075 (N_17075,N_13055,N_12638);
or U17076 (N_17076,N_14655,N_14851);
or U17077 (N_17077,N_12880,N_14344);
or U17078 (N_17078,N_13717,N_14505);
or U17079 (N_17079,N_13154,N_12579);
nor U17080 (N_17080,N_12892,N_13627);
and U17081 (N_17081,N_12668,N_13723);
nor U17082 (N_17082,N_13946,N_13337);
xnor U17083 (N_17083,N_14085,N_12688);
or U17084 (N_17084,N_12773,N_14227);
or U17085 (N_17085,N_13415,N_14337);
or U17086 (N_17086,N_13726,N_12704);
nand U17087 (N_17087,N_12826,N_12948);
nor U17088 (N_17088,N_14223,N_14802);
or U17089 (N_17089,N_13156,N_13168);
and U17090 (N_17090,N_12711,N_14894);
xor U17091 (N_17091,N_14365,N_13303);
or U17092 (N_17092,N_13162,N_14622);
or U17093 (N_17093,N_14873,N_13281);
nor U17094 (N_17094,N_13923,N_12684);
and U17095 (N_17095,N_12992,N_12601);
nor U17096 (N_17096,N_13261,N_13797);
or U17097 (N_17097,N_14966,N_13913);
and U17098 (N_17098,N_14760,N_13277);
or U17099 (N_17099,N_13054,N_13055);
nor U17100 (N_17100,N_14761,N_14888);
nor U17101 (N_17101,N_13263,N_14903);
nand U17102 (N_17102,N_14799,N_14610);
nand U17103 (N_17103,N_13079,N_13168);
or U17104 (N_17104,N_13381,N_14182);
nand U17105 (N_17105,N_14041,N_13108);
and U17106 (N_17106,N_14347,N_13708);
xor U17107 (N_17107,N_14777,N_13733);
nand U17108 (N_17108,N_14545,N_13011);
nand U17109 (N_17109,N_14865,N_14317);
and U17110 (N_17110,N_14640,N_12711);
nor U17111 (N_17111,N_13566,N_12916);
and U17112 (N_17112,N_14631,N_13167);
nand U17113 (N_17113,N_13100,N_13585);
and U17114 (N_17114,N_14351,N_12560);
nand U17115 (N_17115,N_12754,N_13085);
nor U17116 (N_17116,N_14340,N_13998);
or U17117 (N_17117,N_14133,N_13455);
and U17118 (N_17118,N_13738,N_13756);
or U17119 (N_17119,N_12909,N_12654);
and U17120 (N_17120,N_14483,N_14368);
nand U17121 (N_17121,N_13285,N_13592);
and U17122 (N_17122,N_12591,N_14934);
xor U17123 (N_17123,N_14569,N_13066);
or U17124 (N_17124,N_14636,N_12627);
or U17125 (N_17125,N_13421,N_14984);
nand U17126 (N_17126,N_13878,N_13967);
and U17127 (N_17127,N_13964,N_13473);
nand U17128 (N_17128,N_13536,N_14262);
xor U17129 (N_17129,N_14856,N_13827);
and U17130 (N_17130,N_13695,N_13967);
nand U17131 (N_17131,N_14960,N_14290);
and U17132 (N_17132,N_13258,N_12894);
xor U17133 (N_17133,N_13276,N_13724);
nor U17134 (N_17134,N_14622,N_14583);
or U17135 (N_17135,N_13436,N_14840);
nand U17136 (N_17136,N_13712,N_13715);
and U17137 (N_17137,N_14716,N_13304);
nand U17138 (N_17138,N_14106,N_14268);
nor U17139 (N_17139,N_14986,N_13137);
xor U17140 (N_17140,N_13125,N_14836);
or U17141 (N_17141,N_14458,N_12871);
and U17142 (N_17142,N_12947,N_12599);
nor U17143 (N_17143,N_14638,N_13807);
nor U17144 (N_17144,N_14528,N_14189);
nand U17145 (N_17145,N_13041,N_13189);
or U17146 (N_17146,N_13572,N_13406);
xor U17147 (N_17147,N_14297,N_14138);
nor U17148 (N_17148,N_12914,N_13880);
or U17149 (N_17149,N_13094,N_14025);
and U17150 (N_17150,N_13208,N_12833);
nand U17151 (N_17151,N_13894,N_13178);
or U17152 (N_17152,N_14574,N_14219);
nand U17153 (N_17153,N_12928,N_13167);
and U17154 (N_17154,N_14742,N_12985);
nor U17155 (N_17155,N_14395,N_14679);
nor U17156 (N_17156,N_13448,N_14443);
xnor U17157 (N_17157,N_14616,N_12712);
nor U17158 (N_17158,N_13339,N_14141);
nor U17159 (N_17159,N_13229,N_14371);
xor U17160 (N_17160,N_13711,N_12748);
and U17161 (N_17161,N_13572,N_13083);
or U17162 (N_17162,N_13574,N_12626);
nor U17163 (N_17163,N_14733,N_13015);
nand U17164 (N_17164,N_14025,N_14011);
or U17165 (N_17165,N_13191,N_14709);
and U17166 (N_17166,N_14844,N_13472);
nor U17167 (N_17167,N_13118,N_13599);
and U17168 (N_17168,N_13738,N_12873);
or U17169 (N_17169,N_13026,N_13837);
and U17170 (N_17170,N_13682,N_13325);
and U17171 (N_17171,N_13003,N_12701);
nor U17172 (N_17172,N_12892,N_12656);
nor U17173 (N_17173,N_13033,N_13780);
or U17174 (N_17174,N_14541,N_12557);
nor U17175 (N_17175,N_14014,N_14496);
nor U17176 (N_17176,N_12960,N_13092);
and U17177 (N_17177,N_14000,N_13367);
and U17178 (N_17178,N_13079,N_14485);
or U17179 (N_17179,N_14269,N_13892);
nand U17180 (N_17180,N_14831,N_13916);
and U17181 (N_17181,N_13421,N_13724);
nand U17182 (N_17182,N_12893,N_14335);
xnor U17183 (N_17183,N_13183,N_12509);
nand U17184 (N_17184,N_14879,N_12614);
nand U17185 (N_17185,N_13688,N_14964);
nand U17186 (N_17186,N_14611,N_12581);
nand U17187 (N_17187,N_13638,N_12797);
nand U17188 (N_17188,N_14433,N_13007);
nand U17189 (N_17189,N_14715,N_13659);
and U17190 (N_17190,N_14810,N_12595);
nor U17191 (N_17191,N_14767,N_13211);
or U17192 (N_17192,N_14131,N_13999);
and U17193 (N_17193,N_13388,N_13693);
nor U17194 (N_17194,N_13641,N_13917);
and U17195 (N_17195,N_12862,N_13584);
or U17196 (N_17196,N_14389,N_13463);
or U17197 (N_17197,N_14245,N_14848);
and U17198 (N_17198,N_13181,N_12843);
or U17199 (N_17199,N_12932,N_12702);
nand U17200 (N_17200,N_12587,N_13238);
nor U17201 (N_17201,N_13184,N_14437);
nand U17202 (N_17202,N_12547,N_13769);
xnor U17203 (N_17203,N_13942,N_14632);
and U17204 (N_17204,N_12958,N_12633);
xor U17205 (N_17205,N_14671,N_13882);
or U17206 (N_17206,N_14664,N_13727);
nand U17207 (N_17207,N_13609,N_14488);
and U17208 (N_17208,N_14108,N_14446);
xor U17209 (N_17209,N_14025,N_13063);
nand U17210 (N_17210,N_13080,N_13515);
nor U17211 (N_17211,N_14700,N_14084);
nor U17212 (N_17212,N_14842,N_14868);
or U17213 (N_17213,N_14413,N_12839);
xnor U17214 (N_17214,N_13800,N_14172);
nand U17215 (N_17215,N_14343,N_13473);
and U17216 (N_17216,N_12687,N_13506);
or U17217 (N_17217,N_13020,N_14760);
or U17218 (N_17218,N_13833,N_14495);
nor U17219 (N_17219,N_14563,N_13742);
nand U17220 (N_17220,N_13367,N_13755);
nor U17221 (N_17221,N_14869,N_14781);
nand U17222 (N_17222,N_14850,N_13622);
nor U17223 (N_17223,N_13060,N_12541);
or U17224 (N_17224,N_13419,N_13162);
nor U17225 (N_17225,N_13498,N_12742);
xnor U17226 (N_17226,N_14706,N_14391);
nor U17227 (N_17227,N_14679,N_13593);
and U17228 (N_17228,N_14007,N_12986);
or U17229 (N_17229,N_14415,N_14667);
nor U17230 (N_17230,N_13029,N_14415);
and U17231 (N_17231,N_12584,N_14657);
nand U17232 (N_17232,N_13940,N_12787);
and U17233 (N_17233,N_14922,N_14262);
nand U17234 (N_17234,N_13420,N_14588);
and U17235 (N_17235,N_13361,N_12650);
or U17236 (N_17236,N_13740,N_14935);
and U17237 (N_17237,N_14085,N_13652);
or U17238 (N_17238,N_13095,N_13228);
xnor U17239 (N_17239,N_13173,N_14888);
xor U17240 (N_17240,N_13937,N_14533);
nand U17241 (N_17241,N_14117,N_14920);
and U17242 (N_17242,N_12957,N_13322);
nor U17243 (N_17243,N_14674,N_12681);
nand U17244 (N_17244,N_14349,N_14550);
and U17245 (N_17245,N_14456,N_13297);
xor U17246 (N_17246,N_13504,N_14916);
or U17247 (N_17247,N_13698,N_13978);
nand U17248 (N_17248,N_12647,N_12966);
xnor U17249 (N_17249,N_13421,N_14035);
nor U17250 (N_17250,N_12540,N_12794);
or U17251 (N_17251,N_13723,N_14480);
or U17252 (N_17252,N_12516,N_14349);
or U17253 (N_17253,N_13560,N_13917);
xnor U17254 (N_17254,N_12801,N_12882);
nor U17255 (N_17255,N_12609,N_13884);
and U17256 (N_17256,N_12962,N_14693);
nor U17257 (N_17257,N_12514,N_13530);
nand U17258 (N_17258,N_12719,N_14669);
nand U17259 (N_17259,N_13312,N_13950);
or U17260 (N_17260,N_12508,N_12670);
and U17261 (N_17261,N_12525,N_13950);
nand U17262 (N_17262,N_13862,N_12568);
and U17263 (N_17263,N_13977,N_13648);
or U17264 (N_17264,N_12787,N_12791);
xor U17265 (N_17265,N_13386,N_13300);
and U17266 (N_17266,N_13374,N_12570);
or U17267 (N_17267,N_12668,N_14537);
and U17268 (N_17268,N_14018,N_14148);
or U17269 (N_17269,N_14589,N_13432);
or U17270 (N_17270,N_13085,N_12795);
nor U17271 (N_17271,N_13489,N_12736);
nand U17272 (N_17272,N_13317,N_13795);
or U17273 (N_17273,N_13928,N_14357);
nand U17274 (N_17274,N_13350,N_14122);
nand U17275 (N_17275,N_13191,N_13890);
nor U17276 (N_17276,N_12936,N_14024);
or U17277 (N_17277,N_13848,N_13261);
or U17278 (N_17278,N_13172,N_14253);
nor U17279 (N_17279,N_14808,N_13047);
or U17280 (N_17280,N_12655,N_13159);
and U17281 (N_17281,N_14001,N_13886);
nand U17282 (N_17282,N_14103,N_14084);
and U17283 (N_17283,N_14677,N_12929);
nand U17284 (N_17284,N_14876,N_13197);
and U17285 (N_17285,N_13419,N_13212);
nand U17286 (N_17286,N_13287,N_14993);
nor U17287 (N_17287,N_13946,N_13263);
and U17288 (N_17288,N_13881,N_14887);
or U17289 (N_17289,N_12565,N_12871);
nor U17290 (N_17290,N_14045,N_13098);
nor U17291 (N_17291,N_14004,N_14082);
or U17292 (N_17292,N_13427,N_12965);
or U17293 (N_17293,N_14228,N_13846);
nor U17294 (N_17294,N_14370,N_14227);
nand U17295 (N_17295,N_12728,N_12890);
or U17296 (N_17296,N_14881,N_13580);
nor U17297 (N_17297,N_12542,N_13214);
nor U17298 (N_17298,N_14567,N_13097);
and U17299 (N_17299,N_13728,N_13476);
or U17300 (N_17300,N_14569,N_14371);
nand U17301 (N_17301,N_13435,N_14891);
and U17302 (N_17302,N_13295,N_12684);
and U17303 (N_17303,N_14615,N_14963);
nor U17304 (N_17304,N_13986,N_13698);
and U17305 (N_17305,N_13801,N_13220);
and U17306 (N_17306,N_13074,N_14429);
or U17307 (N_17307,N_13111,N_14533);
and U17308 (N_17308,N_13120,N_13436);
and U17309 (N_17309,N_13468,N_13132);
nand U17310 (N_17310,N_13141,N_13064);
or U17311 (N_17311,N_12615,N_14725);
or U17312 (N_17312,N_13644,N_12725);
xnor U17313 (N_17313,N_12947,N_14597);
or U17314 (N_17314,N_13780,N_13644);
xor U17315 (N_17315,N_14416,N_13439);
nand U17316 (N_17316,N_14851,N_14178);
and U17317 (N_17317,N_13948,N_13554);
nor U17318 (N_17318,N_14986,N_12922);
xnor U17319 (N_17319,N_14677,N_14381);
nor U17320 (N_17320,N_13708,N_13074);
nand U17321 (N_17321,N_14792,N_13551);
nor U17322 (N_17322,N_14325,N_13166);
and U17323 (N_17323,N_14908,N_14218);
nor U17324 (N_17324,N_13218,N_13847);
and U17325 (N_17325,N_14468,N_12689);
nor U17326 (N_17326,N_13908,N_14032);
nor U17327 (N_17327,N_14524,N_14639);
nor U17328 (N_17328,N_13423,N_14834);
or U17329 (N_17329,N_14529,N_13176);
or U17330 (N_17330,N_14878,N_14824);
nor U17331 (N_17331,N_13149,N_13495);
and U17332 (N_17332,N_13769,N_14710);
nor U17333 (N_17333,N_13659,N_13138);
or U17334 (N_17334,N_12990,N_13853);
nand U17335 (N_17335,N_12595,N_13513);
and U17336 (N_17336,N_12781,N_13537);
nor U17337 (N_17337,N_14373,N_13414);
nor U17338 (N_17338,N_14564,N_14379);
or U17339 (N_17339,N_12856,N_14816);
nor U17340 (N_17340,N_14954,N_14143);
nand U17341 (N_17341,N_14689,N_13012);
nor U17342 (N_17342,N_13041,N_14259);
or U17343 (N_17343,N_13533,N_13732);
nand U17344 (N_17344,N_13105,N_12532);
nand U17345 (N_17345,N_14681,N_14545);
nor U17346 (N_17346,N_13180,N_12916);
nor U17347 (N_17347,N_13712,N_13538);
and U17348 (N_17348,N_13476,N_12531);
nor U17349 (N_17349,N_13583,N_13944);
and U17350 (N_17350,N_12670,N_13646);
and U17351 (N_17351,N_12817,N_13651);
or U17352 (N_17352,N_12648,N_13848);
nor U17353 (N_17353,N_14331,N_14149);
or U17354 (N_17354,N_14792,N_12509);
nand U17355 (N_17355,N_14299,N_13730);
nand U17356 (N_17356,N_13732,N_12570);
nand U17357 (N_17357,N_13259,N_13721);
nand U17358 (N_17358,N_14496,N_12519);
or U17359 (N_17359,N_14085,N_14064);
or U17360 (N_17360,N_13425,N_13837);
xor U17361 (N_17361,N_13792,N_13257);
nor U17362 (N_17362,N_12525,N_12887);
or U17363 (N_17363,N_13336,N_12646);
and U17364 (N_17364,N_14939,N_12600);
or U17365 (N_17365,N_13974,N_13226);
xnor U17366 (N_17366,N_12593,N_13676);
nor U17367 (N_17367,N_12653,N_14523);
nor U17368 (N_17368,N_12626,N_12938);
and U17369 (N_17369,N_13646,N_12667);
or U17370 (N_17370,N_13482,N_14898);
and U17371 (N_17371,N_13306,N_13812);
and U17372 (N_17372,N_13625,N_13311);
or U17373 (N_17373,N_13321,N_12793);
and U17374 (N_17374,N_14155,N_13410);
xnor U17375 (N_17375,N_14726,N_12810);
nand U17376 (N_17376,N_14790,N_14691);
and U17377 (N_17377,N_13291,N_13444);
nor U17378 (N_17378,N_13470,N_14881);
or U17379 (N_17379,N_13406,N_14658);
and U17380 (N_17380,N_13357,N_14192);
xor U17381 (N_17381,N_13003,N_13920);
nor U17382 (N_17382,N_14425,N_13792);
or U17383 (N_17383,N_14388,N_14976);
nor U17384 (N_17384,N_13111,N_14521);
or U17385 (N_17385,N_14452,N_14540);
and U17386 (N_17386,N_14976,N_13659);
or U17387 (N_17387,N_14626,N_13046);
nand U17388 (N_17388,N_14034,N_14561);
or U17389 (N_17389,N_13450,N_12798);
nor U17390 (N_17390,N_13473,N_12518);
or U17391 (N_17391,N_13462,N_13492);
nor U17392 (N_17392,N_13138,N_12525);
and U17393 (N_17393,N_12523,N_14061);
and U17394 (N_17394,N_14724,N_13842);
nand U17395 (N_17395,N_14115,N_12514);
and U17396 (N_17396,N_14590,N_13185);
nor U17397 (N_17397,N_14663,N_13672);
nor U17398 (N_17398,N_14286,N_13515);
and U17399 (N_17399,N_12742,N_14648);
nand U17400 (N_17400,N_14198,N_14539);
nor U17401 (N_17401,N_13639,N_14598);
nand U17402 (N_17402,N_14342,N_12844);
nor U17403 (N_17403,N_14961,N_13020);
and U17404 (N_17404,N_12940,N_14957);
nor U17405 (N_17405,N_13721,N_14214);
and U17406 (N_17406,N_14999,N_12767);
and U17407 (N_17407,N_13301,N_14710);
and U17408 (N_17408,N_14959,N_13626);
nor U17409 (N_17409,N_12926,N_14676);
or U17410 (N_17410,N_13274,N_13920);
nand U17411 (N_17411,N_14686,N_12656);
or U17412 (N_17412,N_14161,N_14845);
or U17413 (N_17413,N_13306,N_14246);
nand U17414 (N_17414,N_13935,N_13407);
nand U17415 (N_17415,N_13366,N_14944);
nor U17416 (N_17416,N_14119,N_14206);
and U17417 (N_17417,N_12598,N_14763);
nand U17418 (N_17418,N_14835,N_14438);
xor U17419 (N_17419,N_13708,N_12697);
and U17420 (N_17420,N_12947,N_12884);
xnor U17421 (N_17421,N_14352,N_13891);
and U17422 (N_17422,N_12508,N_12786);
or U17423 (N_17423,N_14157,N_13887);
and U17424 (N_17424,N_14616,N_13115);
and U17425 (N_17425,N_13774,N_14412);
or U17426 (N_17426,N_13761,N_12539);
or U17427 (N_17427,N_12971,N_13067);
and U17428 (N_17428,N_13804,N_12564);
nor U17429 (N_17429,N_13410,N_12691);
or U17430 (N_17430,N_13423,N_12786);
or U17431 (N_17431,N_13359,N_14520);
or U17432 (N_17432,N_14653,N_12774);
xor U17433 (N_17433,N_13974,N_13998);
or U17434 (N_17434,N_14107,N_14322);
nor U17435 (N_17435,N_12972,N_13018);
nand U17436 (N_17436,N_13503,N_13216);
nor U17437 (N_17437,N_12908,N_13589);
nor U17438 (N_17438,N_14017,N_14808);
or U17439 (N_17439,N_14555,N_13534);
and U17440 (N_17440,N_12954,N_14319);
or U17441 (N_17441,N_12913,N_13092);
or U17442 (N_17442,N_13348,N_13918);
nor U17443 (N_17443,N_13934,N_14354);
nor U17444 (N_17444,N_12541,N_13222);
xor U17445 (N_17445,N_12591,N_14286);
or U17446 (N_17446,N_12796,N_14873);
xnor U17447 (N_17447,N_12512,N_14098);
nor U17448 (N_17448,N_12733,N_14540);
or U17449 (N_17449,N_13772,N_13890);
nand U17450 (N_17450,N_14477,N_13395);
and U17451 (N_17451,N_13995,N_12564);
and U17452 (N_17452,N_13070,N_12545);
nand U17453 (N_17453,N_12800,N_14238);
or U17454 (N_17454,N_13893,N_14295);
or U17455 (N_17455,N_13116,N_14092);
nor U17456 (N_17456,N_12758,N_14186);
and U17457 (N_17457,N_13731,N_14829);
xnor U17458 (N_17458,N_13823,N_14270);
and U17459 (N_17459,N_12660,N_13131);
and U17460 (N_17460,N_13484,N_13461);
or U17461 (N_17461,N_14127,N_14630);
nor U17462 (N_17462,N_12906,N_14522);
or U17463 (N_17463,N_14862,N_13597);
nor U17464 (N_17464,N_14269,N_13886);
and U17465 (N_17465,N_13092,N_13474);
nand U17466 (N_17466,N_13418,N_14338);
and U17467 (N_17467,N_13358,N_14855);
and U17468 (N_17468,N_14299,N_12533);
and U17469 (N_17469,N_13804,N_14536);
and U17470 (N_17470,N_14928,N_14924);
and U17471 (N_17471,N_14632,N_14265);
xnor U17472 (N_17472,N_13321,N_13163);
xor U17473 (N_17473,N_14857,N_13186);
nand U17474 (N_17474,N_14321,N_13769);
nor U17475 (N_17475,N_14594,N_13325);
or U17476 (N_17476,N_12985,N_13749);
and U17477 (N_17477,N_12812,N_13361);
and U17478 (N_17478,N_12539,N_14881);
or U17479 (N_17479,N_14160,N_13161);
or U17480 (N_17480,N_13604,N_13124);
xnor U17481 (N_17481,N_12644,N_13039);
xnor U17482 (N_17482,N_14547,N_14036);
and U17483 (N_17483,N_14814,N_14560);
nor U17484 (N_17484,N_12529,N_14482);
nor U17485 (N_17485,N_14791,N_14657);
and U17486 (N_17486,N_13673,N_13572);
and U17487 (N_17487,N_13988,N_14643);
nand U17488 (N_17488,N_13251,N_14335);
xor U17489 (N_17489,N_14967,N_12671);
or U17490 (N_17490,N_12804,N_13175);
nor U17491 (N_17491,N_14054,N_14565);
or U17492 (N_17492,N_13937,N_13338);
nor U17493 (N_17493,N_13084,N_12807);
xnor U17494 (N_17494,N_13408,N_12840);
nor U17495 (N_17495,N_12724,N_13837);
xnor U17496 (N_17496,N_13075,N_13594);
and U17497 (N_17497,N_14437,N_12847);
nor U17498 (N_17498,N_12615,N_14117);
nor U17499 (N_17499,N_12569,N_13863);
nor U17500 (N_17500,N_16049,N_17165);
or U17501 (N_17501,N_17086,N_16787);
and U17502 (N_17502,N_15990,N_16616);
nand U17503 (N_17503,N_17443,N_16457);
nor U17504 (N_17504,N_16680,N_16100);
xnor U17505 (N_17505,N_17450,N_15053);
nand U17506 (N_17506,N_16446,N_16666);
and U17507 (N_17507,N_15564,N_15372);
xnor U17508 (N_17508,N_16917,N_15655);
xor U17509 (N_17509,N_17247,N_16831);
or U17510 (N_17510,N_15957,N_17357);
and U17511 (N_17511,N_15011,N_16816);
and U17512 (N_17512,N_16576,N_16358);
nor U17513 (N_17513,N_15156,N_16878);
nand U17514 (N_17514,N_16552,N_16119);
xor U17515 (N_17515,N_17074,N_16362);
or U17516 (N_17516,N_15084,N_16531);
and U17517 (N_17517,N_16126,N_16571);
nand U17518 (N_17518,N_16428,N_15937);
xor U17519 (N_17519,N_15799,N_16626);
or U17520 (N_17520,N_16866,N_15881);
and U17521 (N_17521,N_17437,N_17238);
nand U17522 (N_17522,N_15229,N_15259);
xor U17523 (N_17523,N_15969,N_17442);
and U17524 (N_17524,N_17024,N_15576);
nand U17525 (N_17525,N_15720,N_17191);
nor U17526 (N_17526,N_15823,N_16954);
nor U17527 (N_17527,N_16633,N_15405);
or U17528 (N_17528,N_16182,N_16276);
and U17529 (N_17529,N_15563,N_16952);
nor U17530 (N_17530,N_15164,N_15092);
nand U17531 (N_17531,N_16823,N_16121);
nor U17532 (N_17532,N_15619,N_15496);
or U17533 (N_17533,N_15559,N_15886);
and U17534 (N_17534,N_17459,N_15843);
or U17535 (N_17535,N_17490,N_16432);
nand U17536 (N_17536,N_16298,N_16903);
nor U17537 (N_17537,N_17255,N_16798);
or U17538 (N_17538,N_17037,N_17361);
nor U17539 (N_17539,N_17108,N_15380);
and U17540 (N_17540,N_16395,N_16240);
or U17541 (N_17541,N_15249,N_16158);
nand U17542 (N_17542,N_16580,N_16111);
nand U17543 (N_17543,N_15914,N_16488);
xnor U17544 (N_17544,N_16169,N_17430);
nand U17545 (N_17545,N_16728,N_16069);
and U17546 (N_17546,N_15299,N_15920);
or U17547 (N_17547,N_17338,N_15636);
nor U17548 (N_17548,N_17197,N_16374);
or U17549 (N_17549,N_16749,N_15208);
or U17550 (N_17550,N_16904,N_16441);
nand U17551 (N_17551,N_16178,N_15946);
and U17552 (N_17552,N_15883,N_16543);
nand U17553 (N_17553,N_15373,N_16538);
or U17554 (N_17554,N_16769,N_15765);
nand U17555 (N_17555,N_16913,N_16645);
xor U17556 (N_17556,N_15007,N_17242);
nor U17557 (N_17557,N_16360,N_16629);
nor U17558 (N_17558,N_17019,N_16064);
or U17559 (N_17559,N_16659,N_16758);
nand U17560 (N_17560,N_16868,N_17184);
xnor U17561 (N_17561,N_17279,N_16415);
nand U17562 (N_17562,N_16375,N_17457);
xor U17563 (N_17563,N_16925,N_15033);
and U17564 (N_17564,N_17201,N_16587);
nand U17565 (N_17565,N_15318,N_16485);
nor U17566 (N_17566,N_17090,N_16458);
nor U17567 (N_17567,N_16167,N_16541);
or U17568 (N_17568,N_17436,N_15044);
nor U17569 (N_17569,N_16955,N_16962);
xnor U17570 (N_17570,N_17033,N_16793);
or U17571 (N_17571,N_15732,N_17458);
and U17572 (N_17572,N_15710,N_16054);
and U17573 (N_17573,N_15970,N_15897);
nor U17574 (N_17574,N_16789,N_15131);
nand U17575 (N_17575,N_15477,N_15449);
nor U17576 (N_17576,N_15360,N_16075);
nand U17577 (N_17577,N_17315,N_16639);
nand U17578 (N_17578,N_15925,N_16459);
or U17579 (N_17579,N_15591,N_15678);
nor U17580 (N_17580,N_17101,N_16802);
nand U17581 (N_17581,N_17252,N_16122);
or U17582 (N_17582,N_17472,N_16526);
nand U17583 (N_17583,N_15932,N_16387);
nor U17584 (N_17584,N_16487,N_15901);
nor U17585 (N_17585,N_15708,N_17312);
nor U17586 (N_17586,N_17114,N_16888);
nor U17587 (N_17587,N_16983,N_16825);
nand U17588 (N_17588,N_15699,N_17131);
and U17589 (N_17589,N_15197,N_15325);
or U17590 (N_17590,N_15460,N_15647);
or U17591 (N_17591,N_17047,N_16186);
or U17592 (N_17592,N_16023,N_17415);
xor U17593 (N_17593,N_15388,N_17395);
nor U17594 (N_17594,N_16514,N_15592);
nor U17595 (N_17595,N_15890,N_17035);
nand U17596 (N_17596,N_16990,N_16112);
or U17597 (N_17597,N_16993,N_17118);
nand U17598 (N_17598,N_15342,N_17155);
xnor U17599 (N_17599,N_16830,N_15841);
xnor U17600 (N_17600,N_16038,N_17115);
and U17601 (N_17601,N_15941,N_15098);
xor U17602 (N_17602,N_15049,N_15158);
or U17603 (N_17603,N_15755,N_17198);
nor U17604 (N_17604,N_15419,N_17025);
or U17605 (N_17605,N_15506,N_16922);
nand U17606 (N_17606,N_16927,N_15238);
xnor U17607 (N_17607,N_17360,N_15550);
nor U17608 (N_17608,N_16607,N_15615);
nor U17609 (N_17609,N_15260,N_15431);
nand U17610 (N_17610,N_17220,N_15387);
or U17611 (N_17611,N_17308,N_16619);
nor U17612 (N_17612,N_17017,N_17029);
and U17613 (N_17613,N_17053,N_16416);
nor U17614 (N_17614,N_16486,N_17205);
nor U17615 (N_17615,N_16846,N_17341);
nor U17616 (N_17616,N_16041,N_16501);
or U17617 (N_17617,N_16942,N_17081);
nand U17618 (N_17618,N_17007,N_15366);
or U17619 (N_17619,N_17211,N_17224);
nor U17620 (N_17620,N_17302,N_15295);
and U17621 (N_17621,N_16776,N_16725);
nand U17622 (N_17622,N_17333,N_15285);
nand U17623 (N_17623,N_16348,N_16767);
or U17624 (N_17624,N_17196,N_16491);
and U17625 (N_17625,N_15484,N_16900);
or U17626 (N_17626,N_16665,N_15005);
or U17627 (N_17627,N_17359,N_16957);
nand U17628 (N_17628,N_15339,N_16693);
or U17629 (N_17629,N_16671,N_16337);
nor U17630 (N_17630,N_15635,N_15779);
nand U17631 (N_17631,N_16430,N_16919);
xnor U17632 (N_17632,N_17468,N_15968);
nand U17633 (N_17633,N_17448,N_16996);
or U17634 (N_17634,N_15492,N_17278);
and U17635 (N_17635,N_16554,N_15784);
and U17636 (N_17636,N_16349,N_16807);
and U17637 (N_17637,N_15715,N_17052);
nand U17638 (N_17638,N_16249,N_16250);
or U17639 (N_17639,N_16701,N_15873);
or U17640 (N_17640,N_15082,N_16120);
xor U17641 (N_17641,N_15054,N_17385);
xor U17642 (N_17642,N_16104,N_16821);
nand U17643 (N_17643,N_15187,N_16448);
and U17644 (N_17644,N_15650,N_17173);
nand U17645 (N_17645,N_16184,N_16586);
and U17646 (N_17646,N_16260,N_17087);
and U17647 (N_17647,N_16176,N_15846);
or U17648 (N_17648,N_15291,N_15314);
and U17649 (N_17649,N_15425,N_16732);
and U17650 (N_17650,N_16709,N_16254);
or U17651 (N_17651,N_15926,N_16735);
or U17652 (N_17652,N_16224,N_16423);
and U17653 (N_17653,N_16067,N_16149);
and U17654 (N_17654,N_17069,N_17065);
nor U17655 (N_17655,N_17319,N_15649);
and U17656 (N_17656,N_17139,N_15143);
and U17657 (N_17657,N_15991,N_16039);
nor U17658 (N_17658,N_16536,N_15250);
and U17659 (N_17659,N_16096,N_16215);
or U17660 (N_17660,N_15488,N_15936);
and U17661 (N_17661,N_17091,N_15258);
or U17662 (N_17662,N_15294,N_15792);
nor U17663 (N_17663,N_16836,N_16608);
or U17664 (N_17664,N_17232,N_15476);
nand U17665 (N_17665,N_15512,N_16946);
xnor U17666 (N_17666,N_15628,N_16390);
nand U17667 (N_17667,N_16193,N_15441);
and U17668 (N_17668,N_16009,N_15704);
and U17669 (N_17669,N_16737,N_17141);
nand U17670 (N_17670,N_17241,N_17147);
or U17671 (N_17671,N_15695,N_17126);
or U17672 (N_17672,N_15927,N_16673);
and U17673 (N_17673,N_17016,N_15434);
nor U17674 (N_17674,N_15370,N_15661);
or U17675 (N_17675,N_15604,N_15903);
xor U17676 (N_17676,N_16440,N_15869);
nor U17677 (N_17677,N_16402,N_17233);
nand U17678 (N_17678,N_17112,N_15834);
xnor U17679 (N_17679,N_16978,N_17051);
and U17680 (N_17680,N_15718,N_15648);
xnor U17681 (N_17681,N_15526,N_17405);
nor U17682 (N_17682,N_16648,N_17445);
nor U17683 (N_17683,N_16961,N_15610);
nand U17684 (N_17684,N_17142,N_15327);
or U17685 (N_17685,N_17296,N_16861);
nor U17686 (N_17686,N_15412,N_17491);
nor U17687 (N_17687,N_17159,N_15919);
nor U17688 (N_17688,N_15787,N_16754);
or U17689 (N_17689,N_15422,N_16013);
or U17690 (N_17690,N_15480,N_16051);
nand U17691 (N_17691,N_16863,N_15984);
nor U17692 (N_17692,N_15411,N_16004);
or U17693 (N_17693,N_16975,N_16509);
nand U17694 (N_17694,N_16472,N_16730);
nor U17695 (N_17695,N_17474,N_16073);
or U17696 (N_17696,N_15482,N_15495);
nor U17697 (N_17697,N_15667,N_16929);
and U17698 (N_17698,N_15875,N_15664);
or U17699 (N_17699,N_15770,N_16980);
or U17700 (N_17700,N_16667,N_16634);
xnor U17701 (N_17701,N_16005,N_15570);
nand U17702 (N_17702,N_16066,N_17272);
nand U17703 (N_17703,N_15467,N_15343);
nand U17704 (N_17704,N_15982,N_16003);
or U17705 (N_17705,N_16194,N_15154);
and U17706 (N_17706,N_16865,N_16532);
xor U17707 (N_17707,N_15983,N_17078);
nand U17708 (N_17708,N_16159,N_15808);
nor U17709 (N_17709,N_16944,N_15048);
nor U17710 (N_17710,N_16095,N_16139);
nand U17711 (N_17711,N_15341,N_15382);
nor U17712 (N_17712,N_17305,N_15288);
and U17713 (N_17713,N_15768,N_15428);
nand U17714 (N_17714,N_16370,N_16653);
nor U17715 (N_17715,N_17077,N_15688);
nand U17716 (N_17716,N_16480,N_16827);
nand U17717 (N_17717,N_17153,N_15107);
nand U17718 (N_17718,N_17493,N_15059);
nor U17719 (N_17719,N_17463,N_16650);
nor U17720 (N_17720,N_17235,N_15446);
nand U17721 (N_17721,N_15735,N_15242);
nand U17722 (N_17722,N_17109,N_15525);
or U17723 (N_17723,N_16553,N_15203);
nand U17724 (N_17724,N_16026,N_15537);
or U17725 (N_17725,N_15629,N_16746);
and U17726 (N_17726,N_17397,N_17396);
nand U17727 (N_17727,N_15786,N_16654);
and U17728 (N_17728,N_15383,N_17079);
or U17729 (N_17729,N_15866,N_15010);
and U17730 (N_17730,N_17410,N_16287);
or U17731 (N_17731,N_15023,N_17329);
and U17732 (N_17732,N_16324,N_16131);
and U17733 (N_17733,N_15255,N_17391);
nand U17734 (N_17734,N_15273,N_15300);
nand U17735 (N_17735,N_16890,N_15944);
or U17736 (N_17736,N_15586,N_16757);
and U17737 (N_17737,N_16133,N_15736);
nand U17738 (N_17738,N_17485,N_17178);
xor U17739 (N_17739,N_17300,N_15188);
xor U17740 (N_17740,N_15035,N_17169);
xnor U17741 (N_17741,N_16811,N_15447);
xor U17742 (N_17742,N_15672,N_16151);
and U17743 (N_17743,N_15297,N_17401);
nor U17744 (N_17744,N_16123,N_15884);
xor U17745 (N_17745,N_16156,N_17054);
nand U17746 (N_17746,N_16199,N_15407);
nor U17747 (N_17747,N_16686,N_15303);
nand U17748 (N_17748,N_16869,N_17163);
nor U17749 (N_17749,N_15381,N_15124);
and U17750 (N_17750,N_15176,N_17085);
nor U17751 (N_17751,N_16308,N_16625);
or U17752 (N_17752,N_15632,N_17031);
and U17753 (N_17753,N_17110,N_16219);
nand U17754 (N_17754,N_16164,N_16562);
xor U17755 (N_17755,N_16338,N_15129);
nor U17756 (N_17756,N_16397,N_16695);
and U17757 (N_17757,N_16867,N_17253);
or U17758 (N_17758,N_16453,N_17044);
nor U17759 (N_17759,N_15752,N_16493);
xor U17760 (N_17760,N_16551,N_16632);
or U17761 (N_17761,N_15270,N_16132);
and U17762 (N_17762,N_16773,N_16325);
and U17763 (N_17763,N_17440,N_15392);
and U17764 (N_17764,N_15729,N_16676);
nor U17765 (N_17765,N_16973,N_16399);
nor U17766 (N_17766,N_15829,N_15783);
and U17767 (N_17767,N_16559,N_17000);
and U17768 (N_17768,N_16766,N_17223);
and U17769 (N_17769,N_16713,N_16268);
and U17770 (N_17770,N_16295,N_15080);
nor U17771 (N_17771,N_15797,N_15277);
or U17772 (N_17772,N_17320,N_17377);
or U17773 (N_17773,N_17323,N_16466);
and U17774 (N_17774,N_16226,N_16826);
xor U17775 (N_17775,N_15885,N_16372);
nand U17776 (N_17776,N_15978,N_15021);
and U17777 (N_17777,N_15414,N_16790);
nor U17778 (N_17778,N_16154,N_16967);
and U17779 (N_17779,N_15772,N_15204);
or U17780 (N_17780,N_16956,N_16649);
and U17781 (N_17781,N_17168,N_16644);
nor U17782 (N_17782,N_15247,N_15620);
nand U17783 (N_17783,N_15409,N_17280);
or U17784 (N_17784,N_15483,N_16855);
or U17785 (N_17785,N_17100,N_15195);
and U17786 (N_17786,N_15962,N_16408);
nor U17787 (N_17787,N_15605,N_16323);
or U17788 (N_17788,N_15089,N_15791);
nand U17789 (N_17789,N_15572,N_15997);
and U17790 (N_17790,N_17406,N_17261);
xor U17791 (N_17791,N_15322,N_17061);
xor U17792 (N_17792,N_15758,N_17137);
nand U17793 (N_17793,N_15583,N_15822);
nor U17794 (N_17794,N_15344,N_15585);
nand U17795 (N_17795,N_15179,N_15026);
and U17796 (N_17796,N_16848,N_15541);
xnor U17797 (N_17797,N_17237,N_17149);
or U17798 (N_17798,N_16839,N_15625);
nand U17799 (N_17799,N_15205,N_15289);
nand U17800 (N_17800,N_16597,N_16436);
nor U17801 (N_17801,N_16443,N_16435);
xor U17802 (N_17802,N_16312,N_17182);
and U17803 (N_17803,N_15111,N_17249);
nand U17804 (N_17804,N_16748,N_15569);
xnor U17805 (N_17805,N_15206,N_16697);
and U17806 (N_17806,N_15478,N_16181);
nand U17807 (N_17807,N_16506,N_17301);
and U17808 (N_17808,N_17370,N_16037);
nor U17809 (N_17809,N_17455,N_15662);
and U17810 (N_17810,N_16280,N_17331);
nor U17811 (N_17811,N_17288,N_15502);
nor U17812 (N_17812,N_16474,N_16342);
nor U17813 (N_17813,N_15364,N_16623);
and U17814 (N_17814,N_16166,N_17476);
nor U17815 (N_17815,N_15220,N_16218);
and U17816 (N_17816,N_16384,N_16462);
nor U17817 (N_17817,N_16282,N_17130);
xor U17818 (N_17818,N_16920,N_15140);
nand U17819 (N_17819,N_16565,N_15511);
nand U17820 (N_17820,N_17045,N_15280);
or U17821 (N_17821,N_16690,N_15102);
and U17822 (N_17822,N_15008,N_17122);
and U17823 (N_17823,N_16489,N_16093);
or U17824 (N_17824,N_16679,N_17478);
nand U17825 (N_17825,N_16707,N_16400);
and U17826 (N_17826,N_16599,N_15095);
nor U17827 (N_17827,N_16788,N_16034);
or U17828 (N_17828,N_16221,N_15232);
or U17829 (N_17829,N_16647,N_15845);
nand U17830 (N_17830,N_16368,N_17022);
and U17831 (N_17831,N_17134,N_16492);
and U17832 (N_17832,N_16561,N_17306);
nor U17833 (N_17833,N_16396,N_16389);
or U17834 (N_17834,N_16365,N_15445);
and U17835 (N_17835,N_17172,N_15106);
and U17836 (N_17836,N_15557,N_15740);
nor U17837 (N_17837,N_16434,N_15423);
nor U17838 (N_17838,N_17386,N_17038);
and U17839 (N_17839,N_15362,N_16476);
nor U17840 (N_17840,N_16621,N_15778);
or U17841 (N_17841,N_17298,N_15726);
or U17842 (N_17842,N_17013,N_15723);
nand U17843 (N_17843,N_16505,N_16481);
nor U17844 (N_17844,N_15621,N_15538);
or U17845 (N_17845,N_16992,N_16135);
nand U17846 (N_17846,N_16378,N_16751);
nand U17847 (N_17847,N_16060,N_16063);
and U17848 (N_17848,N_15612,N_15022);
and U17849 (N_17849,N_17265,N_17117);
or U17850 (N_17850,N_15430,N_15980);
nand U17851 (N_17851,N_17208,N_15336);
and U17852 (N_17852,N_15825,N_16796);
xnor U17853 (N_17853,N_16965,N_17387);
nor U17854 (N_17854,N_16461,N_16943);
and U17855 (N_17855,N_17128,N_15031);
nor U17856 (N_17856,N_15864,N_17473);
nor U17857 (N_17857,N_16893,N_17073);
or U17858 (N_17858,N_17489,N_16622);
and U17859 (N_17859,N_16887,N_15196);
nor U17860 (N_17860,N_15283,N_16048);
or U17861 (N_17861,N_15066,N_15304);
or U17862 (N_17862,N_16563,N_15790);
or U17863 (N_17863,N_17427,N_17152);
nand U17864 (N_17864,N_15858,N_16520);
xnor U17865 (N_17865,N_15630,N_16407);
nor U17866 (N_17866,N_15560,N_15332);
nor U17867 (N_17867,N_16207,N_16529);
or U17868 (N_17868,N_17161,N_16808);
or U17869 (N_17869,N_15210,N_16352);
or U17870 (N_17870,N_16989,N_15674);
nor U17871 (N_17871,N_16074,N_15593);
or U17872 (N_17872,N_16314,N_15065);
or U17873 (N_17873,N_16062,N_15761);
or U17874 (N_17874,N_16874,N_16642);
and U17875 (N_17875,N_15181,N_16015);
nand U17876 (N_17876,N_17006,N_16521);
nand U17877 (N_17877,N_15673,N_15182);
and U17878 (N_17878,N_16142,N_15037);
xor U17879 (N_17879,N_15633,N_15368);
or U17880 (N_17880,N_16190,N_15766);
nand U17881 (N_17881,N_16455,N_16091);
or U17882 (N_17882,N_16870,N_15369);
or U17883 (N_17883,N_16556,N_15105);
or U17884 (N_17884,N_15540,N_15464);
xor U17885 (N_17885,N_16347,N_16760);
nor U17886 (N_17886,N_16367,N_15551);
xor U17887 (N_17887,N_15036,N_16988);
nand U17888 (N_17888,N_15109,N_15677);
or U17889 (N_17889,N_15015,N_15544);
xor U17890 (N_17890,N_17162,N_17321);
nor U17891 (N_17891,N_16165,N_16534);
or U17892 (N_17892,N_16969,N_15151);
nand U17893 (N_17893,N_16351,N_15120);
nor U17894 (N_17894,N_16791,N_15017);
and U17895 (N_17895,N_16637,N_15241);
and U17896 (N_17896,N_15357,N_15075);
nor U17897 (N_17897,N_15532,N_15068);
nand U17898 (N_17898,N_17287,N_16677);
or U17899 (N_17899,N_17451,N_15184);
and U17900 (N_17900,N_16813,N_16089);
nor U17901 (N_17901,N_16163,N_15782);
or U17902 (N_17902,N_17289,N_16698);
or U17903 (N_17903,N_15186,N_15915);
nor U17904 (N_17904,N_15707,N_16590);
and U17905 (N_17905,N_15020,N_15177);
nor U17906 (N_17906,N_15987,N_15073);
xor U17907 (N_17907,N_17375,N_17157);
and U17908 (N_17908,N_15974,N_15833);
nand U17909 (N_17909,N_17462,N_16345);
and U17910 (N_17910,N_17188,N_17324);
and U17911 (N_17911,N_17012,N_15359);
and U17912 (N_17912,N_15333,N_15870);
and U17913 (N_17913,N_15471,N_15389);
nor U17914 (N_17914,N_15032,N_16510);
and U17915 (N_17915,N_15706,N_17380);
nand U17916 (N_17916,N_15236,N_17011);
and U17917 (N_17917,N_15528,N_15663);
or U17918 (N_17918,N_16736,N_15928);
nor U17919 (N_17919,N_15070,N_16941);
nor U17920 (N_17920,N_15958,N_16025);
nor U17921 (N_17921,N_15963,N_16057);
and U17922 (N_17922,N_15933,N_16670);
and U17923 (N_17923,N_17213,N_16406);
and U17924 (N_17924,N_15293,N_15733);
nor U17925 (N_17925,N_15083,N_15623);
xor U17926 (N_17926,N_17292,N_17399);
nor U17927 (N_17927,N_17230,N_15058);
xor U17928 (N_17928,N_17227,N_15317);
nand U17929 (N_17929,N_16635,N_16032);
or U17930 (N_17930,N_17219,N_17040);
nor U17931 (N_17931,N_15321,N_15972);
and U17932 (N_17932,N_16704,N_16923);
xnor U17933 (N_17933,N_16482,N_15950);
and U17934 (N_17934,N_17345,N_16477);
nor U17935 (N_17935,N_15155,N_15762);
or U17936 (N_17936,N_16940,N_16656);
nand U17937 (N_17937,N_16233,N_16101);
and U17938 (N_17938,N_17349,N_16046);
nand U17939 (N_17939,N_16783,N_16265);
and U17940 (N_17940,N_15975,N_16213);
nor U17941 (N_17941,N_15377,N_15505);
nor U17942 (N_17942,N_15754,N_17059);
and U17943 (N_17943,N_16834,N_15596);
nand U17944 (N_17944,N_16382,N_15468);
xor U17945 (N_17945,N_16873,N_17432);
xnor U17946 (N_17946,N_15458,N_16411);
and U17947 (N_17947,N_16953,N_16392);
and U17948 (N_17948,N_16183,N_16099);
nor U17949 (N_17949,N_17175,N_16223);
nor U17950 (N_17950,N_16040,N_15350);
and U17951 (N_17951,N_16257,N_15194);
nand U17952 (N_17952,N_16118,N_15338);
or U17953 (N_17953,N_16202,N_15331);
and U17954 (N_17954,N_17433,N_17060);
and U17955 (N_17955,N_15803,N_16768);
and U17956 (N_17956,N_15088,N_16483);
or U17957 (N_17957,N_15439,N_16533);
or U17958 (N_17958,N_16052,N_16422);
nor U17959 (N_17959,N_15093,N_15349);
and U17960 (N_17960,N_15078,N_16424);
or U17961 (N_17961,N_16499,N_16353);
and U17962 (N_17962,N_15498,N_17167);
xnor U17963 (N_17963,N_16998,N_16090);
or U17964 (N_17964,N_15040,N_16794);
xnor U17965 (N_17965,N_15404,N_15844);
xnor U17966 (N_17966,N_16296,N_15689);
and U17967 (N_17967,N_16404,N_17492);
or U17968 (N_17968,N_17293,N_15878);
or U17969 (N_17969,N_15542,N_15659);
and U17970 (N_17970,N_15329,N_16381);
nor U17971 (N_17971,N_15853,N_17310);
or U17972 (N_17972,N_16883,N_16255);
and U17973 (N_17973,N_16724,N_15069);
nand U17974 (N_17974,N_16750,N_16413);
and U17975 (N_17975,N_16377,N_16935);
nor U17976 (N_17976,N_15218,N_16371);
nand U17977 (N_17977,N_15686,N_15684);
nor U17978 (N_17978,N_17259,N_17113);
nor U17979 (N_17979,N_17276,N_15438);
or U17980 (N_17980,N_16593,N_16752);
nand U17981 (N_17981,N_15753,N_16042);
and U17982 (N_17982,N_16778,N_16712);
nor U17983 (N_17983,N_17304,N_17092);
and U17984 (N_17984,N_15616,N_15192);
and U17985 (N_17985,N_17409,N_15386);
nand U17986 (N_17986,N_15698,N_17277);
nor U17987 (N_17987,N_17199,N_15973);
and U17988 (N_17988,N_17218,N_16875);
nand U17989 (N_17989,N_16539,N_17138);
xnor U17990 (N_17990,N_17394,N_17111);
nand U17991 (N_17991,N_15589,N_17028);
and U17992 (N_17992,N_16449,N_16425);
nand U17993 (N_17993,N_15012,N_16017);
nor U17994 (N_17994,N_16305,N_16837);
or U17995 (N_17995,N_15043,N_16319);
and U17996 (N_17996,N_15437,N_16452);
nand U17997 (N_17997,N_16198,N_16843);
nand U17998 (N_17998,N_17274,N_15268);
nor U17999 (N_17999,N_16244,N_16594);
or U18000 (N_18000,N_17369,N_16911);
nand U18001 (N_18001,N_16427,N_16710);
nand U18002 (N_18002,N_15714,N_16708);
nor U18003 (N_18003,N_16658,N_15062);
nand U18004 (N_18004,N_16854,N_15163);
and U18005 (N_18005,N_16061,N_15309);
and U18006 (N_18006,N_16231,N_15796);
nand U18007 (N_18007,N_15096,N_16496);
and U18008 (N_18008,N_17295,N_15888);
nor U18009 (N_18009,N_16910,N_17140);
nor U18010 (N_18010,N_15815,N_15573);
nand U18011 (N_18011,N_16986,N_15231);
or U18012 (N_18012,N_16687,N_15115);
nand U18013 (N_18013,N_15384,N_16628);
xnor U18014 (N_18014,N_15245,N_15879);
and U18015 (N_18015,N_16784,N_15789);
nand U18016 (N_18016,N_17282,N_16516);
nand U18017 (N_18017,N_15871,N_16274);
or U18018 (N_18018,N_16385,N_15272);
nor U18019 (N_18019,N_16386,N_15262);
or U18020 (N_18020,N_17346,N_16711);
or U18021 (N_18021,N_16558,N_15418);
or U18022 (N_18022,N_15330,N_16088);
and U18023 (N_18023,N_16517,N_17403);
nor U18024 (N_18024,N_16175,N_16617);
or U18025 (N_18025,N_16161,N_15165);
nand U18026 (N_18026,N_15709,N_15479);
nor U18027 (N_18027,N_15114,N_15501);
xor U18028 (N_18028,N_15503,N_15922);
nor U18029 (N_18029,N_15861,N_16264);
and U18030 (N_18030,N_17041,N_17420);
nor U18031 (N_18031,N_15034,N_17482);
nand U18032 (N_18032,N_16733,N_15830);
and U18033 (N_18033,N_15071,N_15466);
nand U18034 (N_18034,N_16478,N_16290);
or U18035 (N_18035,N_17275,N_16380);
nor U18036 (N_18036,N_15904,N_16168);
nor U18037 (N_18037,N_16336,N_15061);
or U18038 (N_18038,N_15051,N_15571);
xor U18039 (N_18039,N_16321,N_15461);
or U18040 (N_18040,N_16723,N_16253);
nand U18041 (N_18041,N_15433,N_17454);
or U18042 (N_18042,N_16661,N_17400);
nor U18043 (N_18043,N_15087,N_16107);
or U18044 (N_18044,N_16852,N_15956);
or U18045 (N_18045,N_15319,N_15452);
nor U18046 (N_18046,N_15444,N_15135);
and U18047 (N_18047,N_15805,N_15896);
nand U18048 (N_18048,N_16320,N_16717);
or U18049 (N_18049,N_15701,N_16252);
or U18050 (N_18050,N_15934,N_17368);
nand U18051 (N_18051,N_16859,N_16300);
nand U18052 (N_18052,N_15948,N_15894);
or U18053 (N_18053,N_16858,N_16817);
nor U18054 (N_18054,N_17251,N_16077);
nor U18055 (N_18055,N_16081,N_15568);
or U18056 (N_18056,N_16614,N_16814);
xnor U18057 (N_18057,N_17055,N_17225);
nor U18058 (N_18058,N_15750,N_16447);
and U18059 (N_18059,N_15774,N_16566);
or U18060 (N_18060,N_16460,N_16885);
or U18061 (N_18061,N_16835,N_16765);
or U18062 (N_18062,N_16546,N_16918);
nor U18063 (N_18063,N_17056,N_15375);
and U18064 (N_18064,N_16484,N_17027);
or U18065 (N_18065,N_16899,N_15465);
and U18066 (N_18066,N_16991,N_16928);
nor U18067 (N_18067,N_16205,N_16086);
or U18068 (N_18068,N_15306,N_15530);
nor U18069 (N_18069,N_15748,N_15801);
or U18070 (N_18070,N_15827,N_16809);
nand U18071 (N_18071,N_15965,N_16256);
or U18072 (N_18072,N_17127,N_16518);
or U18073 (N_18073,N_16589,N_15367);
or U18074 (N_18074,N_16641,N_16419);
or U18075 (N_18075,N_15217,N_16530);
or U18076 (N_18076,N_16437,N_15959);
and U18077 (N_18077,N_15119,N_16682);
and U18078 (N_18078,N_16304,N_16098);
nor U18079 (N_18079,N_15286,N_15246);
xnor U18080 (N_18080,N_16050,N_15345);
and U18081 (N_18081,N_16464,N_16872);
and U18082 (N_18082,N_17136,N_16444);
nor U18083 (N_18083,N_15567,N_17393);
and U18084 (N_18084,N_17486,N_16238);
nor U18085 (N_18085,N_16995,N_16229);
and U18086 (N_18086,N_15737,N_16660);
nand U18087 (N_18087,N_16669,N_16630);
nor U18088 (N_18088,N_16357,N_16124);
and U18089 (N_18089,N_15518,N_16939);
nor U18090 (N_18090,N_15546,N_16445);
nand U18091 (N_18091,N_15942,N_15555);
and U18092 (N_18092,N_15960,N_17133);
nor U18093 (N_18093,N_16010,N_16016);
nor U18094 (N_18094,N_15326,N_16277);
xor U18095 (N_18095,N_16734,N_17195);
and U18096 (N_18096,N_16892,N_15211);
nor U18097 (N_18097,N_16970,N_15390);
nor U18098 (N_18098,N_16542,N_15499);
xor U18099 (N_18099,N_15213,N_17330);
xnor U18100 (N_18100,N_16418,N_16192);
nor U18101 (N_18101,N_17496,N_15906);
nand U18102 (N_18102,N_16979,N_15337);
and U18103 (N_18103,N_15150,N_17093);
nand U18104 (N_18104,N_17334,N_16603);
nor U18105 (N_18105,N_16334,N_16235);
nand U18106 (N_18106,N_15172,N_17384);
nor U18107 (N_18107,N_17094,N_15598);
and U18108 (N_18108,N_15679,N_15191);
or U18109 (N_18109,N_17076,N_17480);
nor U18110 (N_18110,N_15868,N_16335);
xnor U18111 (N_18111,N_15334,N_17236);
or U18112 (N_18112,N_16150,N_15645);
xnor U18113 (N_18113,N_15811,N_17088);
nor U18114 (N_18114,N_16094,N_15697);
nor U18115 (N_18115,N_15256,N_15562);
nand U18116 (N_18116,N_16266,N_15305);
or U18117 (N_18117,N_16810,N_16605);
nand U18118 (N_18118,N_15225,N_17431);
and U18119 (N_18119,N_15907,N_17105);
nor U18120 (N_18120,N_17350,N_17234);
and U18121 (N_18121,N_15307,N_15162);
xor U18122 (N_18122,N_15856,N_16718);
and U18123 (N_18123,N_16102,N_17328);
nor U18124 (N_18124,N_16007,N_16731);
nor U18125 (N_18125,N_16782,N_15584);
or U18126 (N_18126,N_15045,N_16044);
and U18127 (N_18127,N_15081,N_16127);
nor U18128 (N_18128,N_16547,N_15728);
or U18129 (N_18129,N_16844,N_16020);
nor U18130 (N_18130,N_15108,N_15523);
nor U18131 (N_18131,N_15041,N_17291);
and U18132 (N_18132,N_16431,N_15052);
and U18133 (N_18133,N_17388,N_15168);
or U18134 (N_18134,N_17014,N_17156);
nand U18135 (N_18135,N_15455,N_15981);
or U18136 (N_18136,N_16678,N_15346);
nand U18137 (N_18137,N_17257,N_17337);
nor U18138 (N_18138,N_15001,N_16210);
nand U18139 (N_18139,N_16191,N_16618);
or U18140 (N_18140,N_15448,N_16652);
xor U18141 (N_18141,N_15651,N_17362);
xor U18142 (N_18142,N_17202,N_16780);
or U18143 (N_18143,N_15807,N_17464);
or U18144 (N_18144,N_16234,N_17095);
and U18145 (N_18145,N_17461,N_16463);
and U18146 (N_18146,N_15865,N_15515);
xor U18147 (N_18147,N_15376,N_17129);
and U18148 (N_18148,N_15267,N_15624);
nand U18149 (N_18149,N_15857,N_15237);
nand U18150 (N_18150,N_16339,N_15814);
xnor U18151 (N_18151,N_15398,N_16021);
xor U18152 (N_18152,N_16239,N_15029);
nand U18153 (N_18153,N_16771,N_16108);
xnor U18154 (N_18154,N_15378,N_16174);
or U18155 (N_18155,N_17072,N_16997);
and U18156 (N_18156,N_16720,N_17398);
nand U18157 (N_18157,N_16172,N_17186);
nand U18158 (N_18158,N_15281,N_16379);
and U18159 (N_18159,N_15908,N_16646);
nor U18160 (N_18160,N_16894,N_15490);
nor U18161 (N_18161,N_15509,N_15363);
or U18162 (N_18162,N_16291,N_15003);
or U18163 (N_18163,N_16185,N_17273);
nor U18164 (N_18164,N_16588,N_16651);
xnor U18165 (N_18165,N_16045,N_15320);
xnor U18166 (N_18166,N_15086,N_17158);
nor U18167 (N_18167,N_17470,N_15643);
or U18168 (N_18168,N_16053,N_16236);
xor U18169 (N_18169,N_16963,N_16359);
or U18170 (N_18170,N_16110,N_16245);
and U18171 (N_18171,N_15463,N_15396);
nand U18172 (N_18172,N_16170,N_16078);
or U18173 (N_18173,N_15785,N_17120);
nor U18174 (N_18174,N_15275,N_15420);
nor U18175 (N_18175,N_15221,N_15757);
or U18176 (N_18176,N_16468,N_15685);
and U18177 (N_18177,N_15117,N_17467);
or U18178 (N_18178,N_15642,N_16310);
xnor U18179 (N_18179,N_15153,N_16129);
or U18180 (N_18180,N_15575,N_15855);
xor U18181 (N_18181,N_15725,N_16722);
or U18182 (N_18182,N_15828,N_16248);
nor U18183 (N_18183,N_17356,N_16901);
or U18184 (N_18184,N_15921,N_16624);
nand U18185 (N_18185,N_17439,N_17402);
nand U18186 (N_18186,N_17174,N_15738);
and U18187 (N_18187,N_17466,N_16824);
or U18188 (N_18188,N_15485,N_16177);
xor U18189 (N_18189,N_17248,N_16409);
nor U18190 (N_18190,N_15850,N_16162);
nand U18191 (N_18191,N_17030,N_15287);
nor U18192 (N_18192,N_16838,N_15744);
nand U18193 (N_18193,N_16600,N_15693);
nand U18194 (N_18194,N_16879,N_16317);
and U18195 (N_18195,N_15614,N_15756);
nand U18196 (N_18196,N_15999,N_16507);
or U18197 (N_18197,N_15421,N_17452);
or U18198 (N_18198,N_16527,N_17270);
or U18199 (N_18199,N_16433,N_16467);
nand U18200 (N_18200,N_15837,N_15769);
nor U18201 (N_18201,N_16421,N_15279);
or U18202 (N_18202,N_16494,N_17119);
or U18203 (N_18203,N_15100,N_17286);
nor U18204 (N_18204,N_17363,N_16871);
nand U18205 (N_18205,N_16152,N_15116);
or U18206 (N_18206,N_15251,N_15876);
and U18207 (N_18207,N_16832,N_16921);
xnor U18208 (N_18208,N_16092,N_16454);
and U18209 (N_18209,N_15724,N_16511);
and U18210 (N_18210,N_15298,N_16475);
nor U18211 (N_18211,N_16806,N_17425);
nand U18212 (N_18212,N_17154,N_15142);
nor U18213 (N_18213,N_15110,N_17477);
nor U18214 (N_18214,N_17183,N_15751);
nor U18215 (N_18215,N_17046,N_16346);
or U18216 (N_18216,N_16354,N_16114);
xor U18217 (N_18217,N_15125,N_17389);
nand U18218 (N_18218,N_15230,N_16795);
or U18219 (N_18219,N_16891,N_15397);
or U18220 (N_18220,N_16331,N_15099);
nor U18221 (N_18221,N_16528,N_16022);
nand U18222 (N_18222,N_15228,N_16001);
or U18223 (N_18223,N_16815,N_15618);
nor U18224 (N_18224,N_16241,N_17411);
nor U18225 (N_18225,N_16106,N_16141);
and U18226 (N_18226,N_15847,N_17269);
nand U18227 (N_18227,N_15747,N_16915);
and U18228 (N_18228,N_16857,N_16341);
nand U18229 (N_18229,N_16805,N_15057);
and U18230 (N_18230,N_16936,N_15491);
and U18231 (N_18231,N_16525,N_16640);
nor U18232 (N_18232,N_15508,N_15385);
and U18233 (N_18233,N_15527,N_15531);
or U18234 (N_18234,N_16662,N_16716);
nand U18235 (N_18235,N_15159,N_15810);
or U18236 (N_18236,N_15316,N_15459);
xor U18237 (N_18237,N_15955,N_17125);
or U18238 (N_18238,N_15494,N_15076);
and U18239 (N_18239,N_15507,N_15064);
and U18240 (N_18240,N_17005,N_16283);
nand U18241 (N_18241,N_15233,N_15742);
nor U18242 (N_18242,N_15745,N_16270);
and U18243 (N_18243,N_15634,N_17200);
xor U18244 (N_18244,N_15804,N_17210);
and U18245 (N_18245,N_17070,N_16786);
nand U18246 (N_18246,N_17106,N_17283);
and U18247 (N_18247,N_15859,N_17039);
and U18248 (N_18248,N_17271,N_17281);
nor U18249 (N_18249,N_16508,N_15669);
nor U18250 (N_18250,N_15274,N_15977);
nand U18251 (N_18251,N_17160,N_15391);
or U18252 (N_18252,N_16173,N_17231);
nor U18253 (N_18253,N_15644,N_17340);
and U18254 (N_18254,N_16742,N_15891);
nand U18255 (N_18255,N_16113,N_17407);
nor U18256 (N_18256,N_15676,N_16006);
and U18257 (N_18257,N_17245,N_15524);
or U18258 (N_18258,N_16535,N_15637);
nand U18259 (N_18259,N_17063,N_15470);
nand U18260 (N_18260,N_16689,N_15219);
nor U18261 (N_18261,N_15613,N_16138);
or U18262 (N_18262,N_16130,N_15424);
nand U18263 (N_18263,N_15654,N_15882);
or U18264 (N_18264,N_15627,N_15660);
and U18265 (N_18265,N_15821,N_16232);
nand U18266 (N_18266,N_16557,N_16373);
xor U18267 (N_18267,N_17376,N_15379);
and U18268 (N_18268,N_17483,N_15535);
and U18269 (N_18269,N_15079,N_15519);
or U18270 (N_18270,N_16344,N_16540);
and U18271 (N_18271,N_16981,N_15278);
and U18272 (N_18272,N_17209,N_15665);
and U18273 (N_18273,N_16302,N_15652);
nor U18274 (N_18274,N_17204,N_17471);
and U18275 (N_18275,N_16555,N_17193);
or U18276 (N_18276,N_16024,N_15832);
nand U18277 (N_18277,N_17217,N_16497);
nand U18278 (N_18278,N_16318,N_16568);
or U18279 (N_18279,N_15042,N_16908);
nand U18280 (N_18280,N_17189,N_16828);
nor U18281 (N_18281,N_16097,N_16125);
nand U18282 (N_18282,N_15355,N_15493);
and U18283 (N_18283,N_16643,N_15994);
nand U18284 (N_18284,N_15055,N_17034);
or U18285 (N_18285,N_15949,N_15243);
nand U18286 (N_18286,N_16694,N_16949);
nor U18287 (N_18287,N_16675,N_16451);
nor U18288 (N_18288,N_16691,N_16070);
and U18289 (N_18289,N_17096,N_16146);
nor U18290 (N_18290,N_17414,N_16569);
nor U18291 (N_18291,N_15025,N_15517);
nor U18292 (N_18292,N_15028,N_16311);
nand U18293 (N_18293,N_15235,N_15113);
or U18294 (N_18294,N_17228,N_15308);
nor U18295 (N_18295,N_15311,N_15889);
nor U18296 (N_18296,N_16932,N_17344);
xor U18297 (N_18297,N_15590,N_16083);
nor U18298 (N_18298,N_17062,N_17036);
nor U18299 (N_18299,N_16293,N_17067);
or U18300 (N_18300,N_15104,N_17226);
or U18301 (N_18301,N_15854,N_16214);
nor U18302 (N_18302,N_17343,N_16706);
xnor U18303 (N_18303,N_17413,N_17177);
or U18304 (N_18304,N_16195,N_17121);
and U18305 (N_18305,N_15717,N_16316);
or U18306 (N_18306,N_16759,N_15254);
nand U18307 (N_18307,N_17018,N_16059);
and U18308 (N_18308,N_15703,N_16364);
nand U18309 (N_18309,N_17371,N_15986);
xor U18310 (N_18310,N_15356,N_15121);
or U18311 (N_18311,N_16000,N_17348);
xnor U18312 (N_18312,N_16574,N_15966);
xnor U18313 (N_18313,N_17285,N_17434);
and U18314 (N_18314,N_16147,N_16560);
nor U18315 (N_18315,N_15239,N_17404);
and U18316 (N_18316,N_15323,N_16350);
nor U18317 (N_18317,N_16216,N_15160);
nand U18318 (N_18318,N_15126,N_15427);
and U18319 (N_18319,N_15056,N_15565);
xnor U18320 (N_18320,N_16663,N_17042);
nor U18321 (N_18321,N_16672,N_16262);
and U18322 (N_18322,N_15798,N_16664);
and U18323 (N_18323,N_16333,N_16261);
nand U18324 (N_18324,N_17181,N_15134);
xnor U18325 (N_18325,N_16882,N_15899);
and U18326 (N_18326,N_16572,N_16204);
nand U18327 (N_18327,N_16958,N_16140);
nand U18328 (N_18328,N_15207,N_16145);
and U18329 (N_18329,N_16850,N_15989);
or U18330 (N_18330,N_16498,N_16548);
and U18331 (N_18331,N_15269,N_15601);
and U18332 (N_18332,N_15047,N_16747);
and U18333 (N_18333,N_15690,N_15863);
nor U18334 (N_18334,N_15741,N_15147);
and U18335 (N_18335,N_16479,N_17423);
or U18336 (N_18336,N_17099,N_16426);
and U18337 (N_18337,N_15909,N_15013);
or U18338 (N_18338,N_15436,N_16343);
nand U18339 (N_18339,N_16258,N_15209);
xor U18340 (N_18340,N_15402,N_16582);
nand U18341 (N_18341,N_16273,N_15244);
xor U18342 (N_18342,N_17424,N_15887);
or U18343 (N_18343,N_15924,N_16271);
nor U18344 (N_18344,N_16719,N_17032);
or U18345 (N_18345,N_15588,N_16160);
nand U18346 (N_18346,N_16668,N_16018);
or U18347 (N_18347,N_15580,N_16196);
and U18348 (N_18348,N_16502,N_15521);
and U18349 (N_18349,N_15456,N_15967);
xnor U18350 (N_18350,N_15178,N_16087);
xnor U18351 (N_18351,N_15091,N_15848);
or U18352 (N_18352,N_17050,N_17132);
and U18353 (N_18353,N_15417,N_15284);
or U18354 (N_18354,N_16755,N_16657);
nand U18355 (N_18355,N_16959,N_15749);
nor U18356 (N_18356,N_17487,N_15545);
nor U18357 (N_18357,N_16971,N_15534);
and U18358 (N_18358,N_16842,N_17314);
nand U18359 (N_18359,N_17297,N_16601);
nand U18360 (N_18360,N_16627,N_17354);
xnor U18361 (N_18361,N_15510,N_17417);
nand U18362 (N_18362,N_16881,N_16043);
nand U18363 (N_18363,N_15603,N_15161);
or U18364 (N_18364,N_15976,N_15773);
and U18365 (N_18365,N_15719,N_15931);
nand U18366 (N_18366,N_15352,N_15148);
nand U18367 (N_18367,N_15533,N_15199);
nand U18368 (N_18368,N_16412,N_17009);
xor U18369 (N_18369,N_15263,N_16902);
nand U18370 (N_18370,N_16330,N_15167);
and U18371 (N_18371,N_17290,N_17057);
xor U18372 (N_18372,N_16960,N_16537);
and U18373 (N_18373,N_15867,N_16567);
nand U18374 (N_18374,N_15731,N_16136);
or U18375 (N_18375,N_15794,N_15212);
or U18376 (N_18376,N_17107,N_16611);
nor U18377 (N_18377,N_15234,N_15900);
nand U18378 (N_18378,N_17215,N_17083);
nor U18379 (N_18379,N_15935,N_16189);
and U18380 (N_18380,N_16779,N_15240);
nand U18381 (N_18381,N_16309,N_17187);
nand U18382 (N_18382,N_15793,N_15851);
or U18383 (N_18383,N_15009,N_16744);
nand U18384 (N_18384,N_16286,N_16655);
or U18385 (N_18385,N_15954,N_16398);
nor U18386 (N_18386,N_17383,N_17049);
nor U18387 (N_18387,N_16926,N_15429);
nand U18388 (N_18388,N_17416,N_15426);
and U18389 (N_18389,N_16085,N_16267);
or U18390 (N_18390,N_16612,N_16907);
nor U18391 (N_18391,N_15641,N_15497);
and U18392 (N_18392,N_15996,N_15473);
nand U18393 (N_18393,N_17366,N_17135);
xor U18394 (N_18394,N_16948,N_16361);
or U18395 (N_18395,N_17104,N_15347);
nand U18396 (N_18396,N_17381,N_16856);
xnor U18397 (N_18397,N_17313,N_15552);
nand U18398 (N_18398,N_16620,N_15312);
nor U18399 (N_18399,N_16148,N_15964);
or U18400 (N_18400,N_16429,N_16450);
and U18401 (N_18401,N_17082,N_17378);
nor U18402 (N_18402,N_16329,N_16288);
or U18403 (N_18403,N_15536,N_15694);
or U18404 (N_18404,N_15809,N_16761);
or U18405 (N_18405,N_15780,N_15224);
or U18406 (N_18406,N_15892,N_15136);
or U18407 (N_18407,N_17023,N_15722);
xor U18408 (N_18408,N_16227,N_16684);
and U18409 (N_18409,N_15606,N_15712);
or U18410 (N_18410,N_16800,N_15721);
or U18411 (N_18411,N_16934,N_15666);
and U18412 (N_18412,N_16636,N_16171);
nand U18413 (N_18413,N_15227,N_16799);
nor U18414 (N_18414,N_15138,N_17373);
and U18415 (N_18415,N_16490,N_16401);
or U18416 (N_18416,N_16886,N_15365);
nand U18417 (N_18417,N_16703,N_16326);
xnor U18418 (N_18418,N_16847,N_17495);
nor U18419 (N_18419,N_15905,N_17422);
nand U18420 (N_18420,N_16604,N_15351);
and U18421 (N_18421,N_17097,N_17449);
nand U18422 (N_18422,N_17382,N_17465);
and U18423 (N_18423,N_17429,N_16115);
nand U18424 (N_18424,N_16756,N_15400);
nor U18425 (N_18425,N_16072,N_15152);
xnor U18426 (N_18426,N_15824,N_15410);
nand U18427 (N_18427,N_15290,N_16822);
xor U18428 (N_18428,N_15301,N_16984);
nor U18429 (N_18429,N_16729,N_16068);
nand U18430 (N_18430,N_15626,N_16209);
and U18431 (N_18431,N_17367,N_16417);
nand U18432 (N_18432,N_16103,N_17250);
or U18433 (N_18433,N_15826,N_15594);
xnor U18434 (N_18434,N_15006,N_16820);
and U18435 (N_18435,N_16592,N_15328);
nor U18436 (N_18436,N_16246,N_15024);
and U18437 (N_18437,N_16549,N_16383);
xnor U18438 (N_18438,N_16297,N_15800);
and U18439 (N_18439,N_16079,N_16638);
nor U18440 (N_18440,N_15435,N_15739);
nor U18441 (N_18441,N_17116,N_17080);
nand U18442 (N_18442,N_15358,N_16573);
or U18443 (N_18443,N_15504,N_15611);
and U18444 (N_18444,N_17240,N_16977);
and U18445 (N_18445,N_15271,N_15658);
and U18446 (N_18446,N_15600,N_15781);
or U18447 (N_18447,N_15141,N_16157);
and U18448 (N_18448,N_15817,N_15354);
nor U18449 (N_18449,N_15558,N_15556);
xnor U18450 (N_18450,N_15938,N_15137);
nand U18451 (N_18451,N_15816,N_15371);
and U18452 (N_18452,N_16473,N_17258);
or U18453 (N_18453,N_16738,N_16011);
or U18454 (N_18454,N_16860,N_16237);
xor U18455 (N_18455,N_15166,N_16228);
nor U18456 (N_18456,N_15700,N_17004);
xor U18457 (N_18457,N_16897,N_17064);
or U18458 (N_18458,N_15985,N_16327);
or U18459 (N_18459,N_16188,N_16584);
xor U18460 (N_18460,N_15852,N_16564);
nor U18461 (N_18461,N_16739,N_15097);
and U18462 (N_18462,N_17185,N_15574);
or U18463 (N_18463,N_17263,N_15692);
nor U18464 (N_18464,N_17150,N_15453);
nand U18465 (N_18465,N_15818,N_16583);
xor U18466 (N_18466,N_16211,N_17453);
xnor U18467 (N_18467,N_17351,N_16931);
or U18468 (N_18468,N_17326,N_17335);
nand U18469 (N_18469,N_16933,N_15836);
nand U18470 (N_18470,N_16328,N_15705);
nor U18471 (N_18471,N_17020,N_15226);
and U18472 (N_18472,N_16714,N_16456);
or U18473 (N_18473,N_15578,N_15806);
xnor U18474 (N_18474,N_15128,N_16284);
or U18475 (N_18475,N_16974,N_16420);
nand U18476 (N_18476,N_16504,N_16203);
or U18477 (N_18477,N_16201,N_16727);
nor U18478 (N_18478,N_16084,N_17103);
nor U18479 (N_18479,N_15253,N_15157);
nor U18480 (N_18480,N_15746,N_16715);
or U18481 (N_18481,N_15170,N_16674);
or U18482 (N_18482,N_16968,N_16851);
nand U18483 (N_18483,N_16116,N_16578);
nor U18484 (N_18484,N_17355,N_17364);
xor U18485 (N_18485,N_15599,N_17303);
xnor U18486 (N_18486,N_17447,N_17180);
or U18487 (N_18487,N_16206,N_16369);
and U18488 (N_18488,N_15940,N_17221);
and U18489 (N_18489,N_15189,N_15016);
nor U18490 (N_18490,N_15282,N_16606);
nand U18491 (N_18491,N_16909,N_17479);
nand U18492 (N_18492,N_15193,N_16912);
xnor U18493 (N_18493,N_17244,N_16581);
and U18494 (N_18494,N_16610,N_16503);
and U18495 (N_18495,N_16950,N_17021);
nor U18496 (N_18496,N_16056,N_16495);
and U18497 (N_18497,N_16278,N_15038);
xnor U18498 (N_18498,N_17066,N_16994);
nor U18499 (N_18499,N_17026,N_15000);
nand U18500 (N_18500,N_16036,N_16631);
or U18501 (N_18501,N_16058,N_16930);
nand U18502 (N_18502,N_15002,N_16609);
nand U18503 (N_18503,N_16523,N_15395);
nor U18504 (N_18504,N_15597,N_16035);
or U18505 (N_18505,N_15198,N_15067);
and U18506 (N_18506,N_15671,N_17145);
nand U18507 (N_18507,N_17339,N_16366);
xnor U18508 (N_18508,N_16801,N_15656);
nand U18509 (N_18509,N_17267,N_15264);
nor U18510 (N_18510,N_16602,N_15413);
nor U18511 (N_18511,N_15880,N_17222);
nor U18512 (N_18512,N_15514,N_17003);
and U18513 (N_18513,N_15716,N_15513);
nand U18514 (N_18514,N_16699,N_15432);
or U18515 (N_18515,N_16972,N_16155);
nor U18516 (N_18516,N_16208,N_15929);
or U18517 (N_18517,N_15112,N_15123);
and U18518 (N_18518,N_15175,N_16200);
or U18519 (N_18519,N_16804,N_16109);
xnor U18520 (N_18520,N_15839,N_15529);
nor U18521 (N_18521,N_16247,N_15767);
or U18522 (N_18522,N_16470,N_16818);
and U18523 (N_18523,N_17206,N_15248);
nand U18524 (N_18524,N_16987,N_16403);
or U18525 (N_18525,N_16596,N_16772);
or U18526 (N_18526,N_16781,N_17469);
nor U18527 (N_18527,N_17176,N_16812);
or U18528 (N_18528,N_15014,N_16065);
nor U18529 (N_18529,N_15911,N_16777);
nor U18530 (N_18530,N_15898,N_16792);
and U18531 (N_18531,N_16692,N_16579);
or U18532 (N_18532,N_16301,N_17098);
and U18533 (N_18533,N_16785,N_16220);
and U18534 (N_18534,N_15913,N_16585);
xnor U18535 (N_18535,N_16292,N_17426);
or U18536 (N_18536,N_15516,N_17264);
xnor U18537 (N_18537,N_15760,N_15292);
or U18538 (N_18538,N_16938,N_16519);
or U18539 (N_18539,N_17347,N_15617);
nand U18540 (N_18540,N_16315,N_15923);
or U18541 (N_18541,N_16029,N_15127);
xnor U18542 (N_18542,N_16289,N_15174);
xor U18543 (N_18543,N_15118,N_15202);
and U18544 (N_18544,N_16544,N_17456);
nor U18545 (N_18545,N_16797,N_17239);
and U18546 (N_18546,N_17494,N_16819);
or U18547 (N_18547,N_16803,N_17309);
nor U18548 (N_18548,N_15265,N_16222);
xnor U18549 (N_18549,N_16251,N_15486);
nor U18550 (N_18550,N_16982,N_17372);
xor U18551 (N_18551,N_15912,N_16071);
or U18552 (N_18552,N_15691,N_15577);
xnor U18553 (N_18553,N_16014,N_16702);
and U18554 (N_18554,N_17058,N_16153);
nand U18555 (N_18555,N_16833,N_15939);
and U18556 (N_18556,N_15520,N_15171);
nand U18557 (N_18557,N_15681,N_16966);
and U18558 (N_18558,N_17392,N_15103);
and U18559 (N_18559,N_17336,N_16376);
xor U18560 (N_18560,N_16841,N_15696);
or U18561 (N_18561,N_15842,N_15918);
or U18562 (N_18562,N_16117,N_15860);
and U18563 (N_18563,N_17379,N_16524);
and U18564 (N_18564,N_15549,N_15668);
nor U18565 (N_18565,N_15727,N_16143);
or U18566 (N_18566,N_17390,N_16259);
nand U18567 (N_18567,N_15072,N_16008);
nand U18568 (N_18568,N_15296,N_15862);
nor U18569 (N_18569,N_15638,N_15657);
xor U18570 (N_18570,N_16033,N_15711);
nand U18571 (N_18571,N_16027,N_15340);
and U18572 (N_18572,N_15566,N_15335);
and U18573 (N_18573,N_16225,N_15462);
xnor U18574 (N_18574,N_17325,N_16512);
nand U18575 (N_18575,N_15539,N_15840);
nor U18576 (N_18576,N_17260,N_15046);
or U18577 (N_18577,N_15683,N_15063);
nor U18578 (N_18578,N_15085,N_17256);
nand U18579 (N_18579,N_16303,N_17307);
and U18580 (N_18580,N_15132,N_15631);
xnor U18581 (N_18581,N_15457,N_16294);
and U18582 (N_18582,N_15451,N_16212);
xor U18583 (N_18583,N_15893,N_15481);
nor U18584 (N_18584,N_16012,N_17075);
nand U18585 (N_18585,N_17499,N_15543);
nand U18586 (N_18586,N_16410,N_17412);
and U18587 (N_18587,N_16515,N_15872);
and U18588 (N_18588,N_15416,N_15252);
or U18589 (N_18589,N_15930,N_17071);
or U18590 (N_18590,N_17318,N_15200);
xnor U18591 (N_18591,N_16405,N_15101);
or U18592 (N_18592,N_17262,N_16217);
and U18593 (N_18593,N_16829,N_15361);
nor U18594 (N_18594,N_17212,N_15004);
and U18595 (N_18595,N_17164,N_16105);
nand U18596 (N_18596,N_17488,N_15581);
xor U18597 (N_18597,N_16681,N_17327);
nand U18598 (N_18598,N_16263,N_15988);
nor U18599 (N_18599,N_16570,N_15776);
and U18600 (N_18600,N_15522,N_17068);
or U18601 (N_18601,N_15979,N_17317);
nand U18602 (N_18602,N_15640,N_17008);
nand U18603 (N_18603,N_15602,N_16355);
nand U18604 (N_18604,N_15993,N_15185);
nor U18605 (N_18605,N_16179,N_17254);
nor U18606 (N_18606,N_15874,N_15788);
xnor U18607 (N_18607,N_16279,N_15027);
and U18608 (N_18608,N_15474,N_15353);
nand U18609 (N_18609,N_15553,N_17166);
and U18610 (N_18610,N_16999,N_17102);
nand U18611 (N_18611,N_16775,N_16388);
or U18612 (N_18612,N_15548,N_15469);
nand U18613 (N_18613,N_16862,N_16128);
xnor U18614 (N_18614,N_15183,N_16031);
and U18615 (N_18615,N_15579,N_15587);
or U18616 (N_18616,N_15173,N_17089);
and U18617 (N_18617,N_17421,N_16914);
or U18618 (N_18618,N_17179,N_16740);
and U18619 (N_18619,N_17148,N_15992);
nand U18620 (N_18620,N_17203,N_15149);
or U18621 (N_18621,N_15310,N_16895);
nor U18622 (N_18622,N_17484,N_16683);
nor U18623 (N_18623,N_15895,N_15653);
and U18624 (N_18624,N_17144,N_15315);
nor U18625 (N_18625,N_16522,N_15812);
nor U18626 (N_18626,N_16905,N_17194);
nand U18627 (N_18627,N_17002,N_16951);
or U18628 (N_18628,N_17435,N_16976);
and U18629 (N_18629,N_15276,N_15440);
nand U18630 (N_18630,N_15730,N_16180);
and U18631 (N_18631,N_17207,N_17294);
and U18632 (N_18632,N_16082,N_16363);
nand U18633 (N_18633,N_16269,N_16340);
or U18634 (N_18634,N_17151,N_16985);
or U18635 (N_18635,N_16080,N_16272);
and U18636 (N_18636,N_17299,N_16047);
and U18637 (N_18637,N_16439,N_16137);
nor U18638 (N_18638,N_16705,N_15595);
nor U18639 (N_18639,N_16916,N_15313);
or U18640 (N_18640,N_17284,N_16876);
or U18641 (N_18641,N_15910,N_17441);
and U18642 (N_18642,N_16281,N_16356);
and U18643 (N_18643,N_15917,N_16471);
nand U18644 (N_18644,N_16721,N_15902);
nor U18645 (N_18645,N_15838,N_16442);
or U18646 (N_18646,N_15216,N_17084);
and U18647 (N_18647,N_15302,N_15639);
nand U18648 (N_18648,N_15050,N_17481);
or U18649 (N_18649,N_16187,N_15180);
nor U18650 (N_18650,N_17001,N_15399);
nor U18651 (N_18651,N_15018,N_17365);
or U18652 (N_18652,N_16688,N_16577);
nor U18653 (N_18653,N_16030,N_17170);
nor U18654 (N_18654,N_15961,N_16884);
nor U18655 (N_18655,N_15222,N_16394);
or U18656 (N_18656,N_16896,N_17010);
and U18657 (N_18657,N_15947,N_16864);
nand U18658 (N_18658,N_15039,N_15743);
and U18659 (N_18659,N_15214,N_17229);
and U18660 (N_18660,N_15777,N_16889);
and U18661 (N_18661,N_16770,N_15775);
and U18662 (N_18662,N_15916,N_17446);
or U18663 (N_18663,N_15454,N_16575);
and U18664 (N_18664,N_16028,N_15952);
nor U18665 (N_18665,N_16393,N_15802);
and U18666 (N_18666,N_16414,N_17268);
nor U18667 (N_18667,N_15759,N_17418);
nand U18668 (N_18668,N_17048,N_16299);
or U18669 (N_18669,N_15257,N_16391);
xnor U18670 (N_18670,N_15813,N_15442);
nor U18671 (N_18671,N_15130,N_15995);
or U18672 (N_18672,N_17438,N_15500);
nand U18673 (N_18673,N_16741,N_17192);
or U18674 (N_18674,N_16840,N_16700);
nand U18675 (N_18675,N_15609,N_16134);
nand U18676 (N_18676,N_15201,N_15030);
or U18677 (N_18677,N_15415,N_15450);
nand U18678 (N_18678,N_15190,N_15324);
nand U18679 (N_18679,N_17353,N_17043);
and U18680 (N_18680,N_15771,N_16465);
nand U18681 (N_18681,N_17460,N_15472);
nor U18682 (N_18682,N_16615,N_16845);
nor U18683 (N_18683,N_17419,N_15223);
nor U18684 (N_18684,N_15607,N_17358);
nand U18685 (N_18685,N_16307,N_17190);
xor U18686 (N_18686,N_17311,N_16322);
or U18687 (N_18687,N_16853,N_15670);
nor U18688 (N_18688,N_16285,N_17316);
nor U18689 (N_18689,N_17342,N_17143);
or U18690 (N_18690,N_15687,N_15133);
nand U18691 (N_18691,N_17123,N_17146);
and U18692 (N_18692,N_16937,N_16550);
nor U18693 (N_18693,N_15090,N_16332);
nor U18694 (N_18694,N_17171,N_15680);
and U18695 (N_18695,N_15831,N_16898);
xnor U18696 (N_18696,N_17475,N_15374);
and U18697 (N_18697,N_15582,N_15608);
nand U18698 (N_18698,N_15060,N_15139);
nand U18699 (N_18699,N_17015,N_16906);
or U18700 (N_18700,N_16613,N_15734);
nand U18701 (N_18701,N_16313,N_15408);
or U18702 (N_18702,N_15074,N_15849);
nor U18703 (N_18703,N_16945,N_15403);
nor U18704 (N_18704,N_15702,N_16764);
nor U18705 (N_18705,N_15261,N_15713);
or U18706 (N_18706,N_16924,N_15401);
or U18707 (N_18707,N_16595,N_16753);
nand U18708 (N_18708,N_16513,N_16763);
and U18709 (N_18709,N_16197,N_17322);
nor U18710 (N_18710,N_15763,N_16306);
nand U18711 (N_18711,N_16469,N_17266);
xor U18712 (N_18712,N_15819,N_15943);
and U18713 (N_18713,N_16743,N_17374);
xor U18714 (N_18714,N_15835,N_15795);
nand U18715 (N_18715,N_17408,N_15393);
xnor U18716 (N_18716,N_15764,N_16947);
and U18717 (N_18717,N_16696,N_17352);
or U18718 (N_18718,N_15489,N_15820);
nor U18719 (N_18719,N_16877,N_15145);
and U18720 (N_18720,N_15094,N_17428);
nand U18721 (N_18721,N_17243,N_15169);
nor U18722 (N_18722,N_15998,N_17332);
and U18723 (N_18723,N_15971,N_16144);
nor U18724 (N_18724,N_16076,N_16598);
or U18725 (N_18725,N_16745,N_15443);
or U18726 (N_18726,N_16964,N_16242);
nor U18727 (N_18727,N_15675,N_16275);
nor U18728 (N_18728,N_16438,N_17124);
xnor U18729 (N_18729,N_15945,N_16685);
or U18730 (N_18730,N_15266,N_16762);
and U18731 (N_18731,N_15019,N_15622);
or U18732 (N_18732,N_17214,N_17246);
or U18733 (N_18733,N_15394,N_15215);
nand U18734 (N_18734,N_15487,N_16545);
xor U18735 (N_18735,N_15077,N_15682);
nor U18736 (N_18736,N_15406,N_17216);
or U18737 (N_18737,N_16500,N_15951);
xor U18738 (N_18738,N_15646,N_15547);
and U18739 (N_18739,N_16019,N_15122);
and U18740 (N_18740,N_16774,N_15554);
xnor U18741 (N_18741,N_16055,N_15146);
nor U18742 (N_18742,N_16002,N_15144);
nor U18743 (N_18743,N_15561,N_15475);
nor U18744 (N_18744,N_16243,N_17497);
or U18745 (N_18745,N_16230,N_15953);
and U18746 (N_18746,N_16849,N_16726);
nor U18747 (N_18747,N_16591,N_17498);
and U18748 (N_18748,N_17444,N_15877);
nand U18749 (N_18749,N_16880,N_15348);
nand U18750 (N_18750,N_17364,N_16190);
or U18751 (N_18751,N_15152,N_15848);
nand U18752 (N_18752,N_16724,N_16867);
nor U18753 (N_18753,N_16851,N_16581);
nand U18754 (N_18754,N_15325,N_16883);
and U18755 (N_18755,N_17062,N_17221);
or U18756 (N_18756,N_17254,N_16479);
and U18757 (N_18757,N_15691,N_17320);
and U18758 (N_18758,N_15857,N_16372);
and U18759 (N_18759,N_16943,N_16472);
or U18760 (N_18760,N_16958,N_16706);
nand U18761 (N_18761,N_16401,N_15696);
or U18762 (N_18762,N_15248,N_17168);
or U18763 (N_18763,N_15578,N_16171);
and U18764 (N_18764,N_16901,N_15864);
nand U18765 (N_18765,N_16889,N_16149);
nand U18766 (N_18766,N_15889,N_15712);
and U18767 (N_18767,N_17135,N_15920);
and U18768 (N_18768,N_17142,N_16655);
and U18769 (N_18769,N_15400,N_15535);
or U18770 (N_18770,N_16963,N_16986);
xnor U18771 (N_18771,N_17276,N_17009);
nand U18772 (N_18772,N_16137,N_16468);
or U18773 (N_18773,N_16332,N_17355);
nor U18774 (N_18774,N_16919,N_15303);
xor U18775 (N_18775,N_15562,N_17251);
and U18776 (N_18776,N_16671,N_15749);
nand U18777 (N_18777,N_16908,N_15531);
nand U18778 (N_18778,N_15605,N_15429);
nor U18779 (N_18779,N_17308,N_15343);
nor U18780 (N_18780,N_17393,N_15624);
and U18781 (N_18781,N_15741,N_16826);
or U18782 (N_18782,N_15512,N_16552);
nor U18783 (N_18783,N_16762,N_15850);
or U18784 (N_18784,N_15152,N_16877);
nor U18785 (N_18785,N_16070,N_15844);
xnor U18786 (N_18786,N_17200,N_15080);
or U18787 (N_18787,N_16770,N_16886);
nor U18788 (N_18788,N_17058,N_15767);
nor U18789 (N_18789,N_15443,N_17489);
nand U18790 (N_18790,N_16221,N_15362);
and U18791 (N_18791,N_17229,N_17297);
or U18792 (N_18792,N_17267,N_15152);
nor U18793 (N_18793,N_16246,N_17247);
or U18794 (N_18794,N_16692,N_17331);
xnor U18795 (N_18795,N_15464,N_15359);
and U18796 (N_18796,N_15293,N_15061);
and U18797 (N_18797,N_15053,N_17179);
nand U18798 (N_18798,N_17271,N_16440);
xor U18799 (N_18799,N_17494,N_16330);
and U18800 (N_18800,N_17088,N_15899);
xor U18801 (N_18801,N_17391,N_16929);
and U18802 (N_18802,N_15518,N_17086);
and U18803 (N_18803,N_16397,N_17321);
nand U18804 (N_18804,N_16044,N_15347);
and U18805 (N_18805,N_15735,N_15483);
or U18806 (N_18806,N_16832,N_15704);
nand U18807 (N_18807,N_17371,N_17223);
or U18808 (N_18808,N_15950,N_16646);
and U18809 (N_18809,N_16027,N_15806);
and U18810 (N_18810,N_17119,N_15793);
nand U18811 (N_18811,N_17169,N_15366);
xnor U18812 (N_18812,N_16054,N_15230);
nor U18813 (N_18813,N_16464,N_15224);
and U18814 (N_18814,N_15556,N_17121);
nand U18815 (N_18815,N_15381,N_15314);
nor U18816 (N_18816,N_17367,N_16557);
xor U18817 (N_18817,N_15850,N_17078);
nand U18818 (N_18818,N_16577,N_17069);
nor U18819 (N_18819,N_16724,N_16588);
nand U18820 (N_18820,N_15899,N_15129);
nor U18821 (N_18821,N_17455,N_15790);
and U18822 (N_18822,N_15054,N_16580);
nor U18823 (N_18823,N_15138,N_16391);
and U18824 (N_18824,N_17116,N_16246);
nor U18825 (N_18825,N_17404,N_17436);
or U18826 (N_18826,N_15668,N_16434);
nor U18827 (N_18827,N_17122,N_17184);
nand U18828 (N_18828,N_16109,N_15321);
and U18829 (N_18829,N_17451,N_15888);
nand U18830 (N_18830,N_15207,N_15880);
and U18831 (N_18831,N_16055,N_15480);
and U18832 (N_18832,N_15326,N_16881);
nand U18833 (N_18833,N_17384,N_16016);
or U18834 (N_18834,N_16436,N_16803);
nor U18835 (N_18835,N_15935,N_17201);
nor U18836 (N_18836,N_16290,N_17226);
nor U18837 (N_18837,N_17312,N_16672);
xor U18838 (N_18838,N_16064,N_16699);
or U18839 (N_18839,N_16515,N_16846);
and U18840 (N_18840,N_15828,N_16949);
nor U18841 (N_18841,N_17024,N_16437);
or U18842 (N_18842,N_15092,N_16284);
and U18843 (N_18843,N_15645,N_15411);
and U18844 (N_18844,N_16408,N_17226);
xnor U18845 (N_18845,N_16036,N_15551);
or U18846 (N_18846,N_17440,N_17062);
nand U18847 (N_18847,N_15246,N_17326);
nand U18848 (N_18848,N_15350,N_16352);
xor U18849 (N_18849,N_16266,N_16625);
or U18850 (N_18850,N_16471,N_16153);
or U18851 (N_18851,N_15363,N_15726);
and U18852 (N_18852,N_17258,N_16123);
or U18853 (N_18853,N_16788,N_15467);
nor U18854 (N_18854,N_15640,N_16549);
and U18855 (N_18855,N_17090,N_16345);
or U18856 (N_18856,N_16388,N_15266);
and U18857 (N_18857,N_15274,N_17142);
and U18858 (N_18858,N_15240,N_16293);
nor U18859 (N_18859,N_16421,N_16083);
and U18860 (N_18860,N_17198,N_15091);
and U18861 (N_18861,N_15156,N_17256);
and U18862 (N_18862,N_16593,N_16207);
xnor U18863 (N_18863,N_16362,N_15846);
and U18864 (N_18864,N_17149,N_16947);
and U18865 (N_18865,N_17270,N_16726);
xor U18866 (N_18866,N_17141,N_16128);
nor U18867 (N_18867,N_15556,N_16202);
or U18868 (N_18868,N_16113,N_15788);
nand U18869 (N_18869,N_16616,N_16353);
nand U18870 (N_18870,N_16243,N_15696);
nand U18871 (N_18871,N_16178,N_16559);
or U18872 (N_18872,N_16230,N_16312);
or U18873 (N_18873,N_16337,N_16868);
or U18874 (N_18874,N_15988,N_15446);
nor U18875 (N_18875,N_17181,N_16337);
or U18876 (N_18876,N_16682,N_15946);
nor U18877 (N_18877,N_15329,N_16439);
nor U18878 (N_18878,N_15850,N_17340);
or U18879 (N_18879,N_17440,N_15937);
nand U18880 (N_18880,N_15889,N_15042);
and U18881 (N_18881,N_17474,N_16149);
or U18882 (N_18882,N_16483,N_17074);
nor U18883 (N_18883,N_17400,N_16772);
nand U18884 (N_18884,N_15766,N_17168);
xor U18885 (N_18885,N_16337,N_15813);
or U18886 (N_18886,N_15311,N_16657);
or U18887 (N_18887,N_15521,N_16032);
nand U18888 (N_18888,N_15456,N_16478);
nand U18889 (N_18889,N_15225,N_17457);
nor U18890 (N_18890,N_17462,N_16805);
nor U18891 (N_18891,N_15526,N_16585);
and U18892 (N_18892,N_16156,N_16700);
and U18893 (N_18893,N_15552,N_17340);
and U18894 (N_18894,N_17293,N_15600);
nand U18895 (N_18895,N_15695,N_16632);
nand U18896 (N_18896,N_17002,N_15779);
nand U18897 (N_18897,N_15912,N_15479);
nor U18898 (N_18898,N_15941,N_15903);
and U18899 (N_18899,N_15918,N_15003);
or U18900 (N_18900,N_17427,N_15878);
or U18901 (N_18901,N_15966,N_15845);
nor U18902 (N_18902,N_16237,N_15465);
nand U18903 (N_18903,N_15570,N_16181);
or U18904 (N_18904,N_15146,N_15918);
nand U18905 (N_18905,N_16716,N_15306);
nand U18906 (N_18906,N_16235,N_16875);
and U18907 (N_18907,N_15222,N_15120);
or U18908 (N_18908,N_17190,N_16469);
and U18909 (N_18909,N_17415,N_17204);
nand U18910 (N_18910,N_17160,N_16753);
or U18911 (N_18911,N_15111,N_16642);
nand U18912 (N_18912,N_16702,N_16853);
or U18913 (N_18913,N_15750,N_15316);
or U18914 (N_18914,N_17329,N_15551);
nand U18915 (N_18915,N_17075,N_17352);
nor U18916 (N_18916,N_16808,N_17476);
xor U18917 (N_18917,N_15081,N_17237);
nor U18918 (N_18918,N_15475,N_16576);
nand U18919 (N_18919,N_17111,N_16767);
or U18920 (N_18920,N_17264,N_15085);
or U18921 (N_18921,N_16472,N_16939);
nor U18922 (N_18922,N_16387,N_16615);
and U18923 (N_18923,N_16682,N_16412);
nor U18924 (N_18924,N_17335,N_16736);
and U18925 (N_18925,N_15014,N_16124);
nand U18926 (N_18926,N_15331,N_16500);
nor U18927 (N_18927,N_16909,N_15945);
and U18928 (N_18928,N_17317,N_17059);
nand U18929 (N_18929,N_15720,N_15998);
nor U18930 (N_18930,N_15398,N_16080);
nand U18931 (N_18931,N_16312,N_16098);
or U18932 (N_18932,N_15125,N_16145);
nand U18933 (N_18933,N_16786,N_15735);
nand U18934 (N_18934,N_16513,N_17279);
or U18935 (N_18935,N_15727,N_16551);
and U18936 (N_18936,N_16911,N_16892);
xor U18937 (N_18937,N_15995,N_16428);
xor U18938 (N_18938,N_17042,N_17301);
and U18939 (N_18939,N_15567,N_16527);
nor U18940 (N_18940,N_16217,N_15307);
xnor U18941 (N_18941,N_15945,N_16205);
nor U18942 (N_18942,N_16678,N_16544);
xor U18943 (N_18943,N_15969,N_16013);
nor U18944 (N_18944,N_16338,N_16751);
nand U18945 (N_18945,N_16331,N_16000);
nand U18946 (N_18946,N_15926,N_15913);
and U18947 (N_18947,N_15333,N_17344);
and U18948 (N_18948,N_17264,N_17064);
xor U18949 (N_18949,N_15316,N_17098);
and U18950 (N_18950,N_15011,N_15889);
xor U18951 (N_18951,N_15302,N_15948);
and U18952 (N_18952,N_16135,N_17189);
or U18953 (N_18953,N_15576,N_15999);
nand U18954 (N_18954,N_16164,N_15540);
or U18955 (N_18955,N_15335,N_16945);
xnor U18956 (N_18956,N_16839,N_16159);
or U18957 (N_18957,N_15658,N_15002);
xnor U18958 (N_18958,N_15758,N_15511);
nor U18959 (N_18959,N_17370,N_17308);
or U18960 (N_18960,N_17332,N_16130);
and U18961 (N_18961,N_16652,N_17351);
nor U18962 (N_18962,N_17448,N_16907);
nand U18963 (N_18963,N_15964,N_17377);
nor U18964 (N_18964,N_15240,N_17167);
xnor U18965 (N_18965,N_16696,N_15572);
nor U18966 (N_18966,N_16300,N_15858);
nand U18967 (N_18967,N_15994,N_16977);
nor U18968 (N_18968,N_16033,N_17359);
or U18969 (N_18969,N_15176,N_16927);
xnor U18970 (N_18970,N_15622,N_17241);
and U18971 (N_18971,N_17163,N_17374);
and U18972 (N_18972,N_15438,N_17112);
nand U18973 (N_18973,N_17471,N_16493);
and U18974 (N_18974,N_16284,N_15961);
nand U18975 (N_18975,N_15416,N_16876);
nand U18976 (N_18976,N_16929,N_16043);
and U18977 (N_18977,N_16904,N_16834);
and U18978 (N_18978,N_17496,N_16242);
xor U18979 (N_18979,N_16025,N_17119);
nor U18980 (N_18980,N_16679,N_15685);
or U18981 (N_18981,N_15558,N_17439);
or U18982 (N_18982,N_17173,N_17486);
nand U18983 (N_18983,N_16238,N_16599);
or U18984 (N_18984,N_15728,N_16619);
xnor U18985 (N_18985,N_16626,N_16406);
or U18986 (N_18986,N_17140,N_16363);
and U18987 (N_18987,N_15206,N_16121);
nor U18988 (N_18988,N_16799,N_16865);
nor U18989 (N_18989,N_16339,N_15746);
nor U18990 (N_18990,N_15992,N_16961);
nor U18991 (N_18991,N_16633,N_15594);
nor U18992 (N_18992,N_15906,N_15009);
nand U18993 (N_18993,N_15908,N_16014);
or U18994 (N_18994,N_16952,N_15420);
nand U18995 (N_18995,N_16744,N_16752);
and U18996 (N_18996,N_16602,N_15252);
xnor U18997 (N_18997,N_16335,N_16929);
nand U18998 (N_18998,N_16235,N_15729);
or U18999 (N_18999,N_16452,N_15060);
or U19000 (N_19000,N_17320,N_17177);
xor U19001 (N_19001,N_15417,N_16662);
nor U19002 (N_19002,N_16486,N_15290);
or U19003 (N_19003,N_16702,N_17003);
xor U19004 (N_19004,N_16213,N_17040);
nor U19005 (N_19005,N_16722,N_15301);
or U19006 (N_19006,N_17103,N_15057);
xor U19007 (N_19007,N_16352,N_15815);
xnor U19008 (N_19008,N_15533,N_16875);
nand U19009 (N_19009,N_16625,N_17397);
nor U19010 (N_19010,N_15073,N_15698);
and U19011 (N_19011,N_15281,N_15001);
nand U19012 (N_19012,N_16602,N_15392);
or U19013 (N_19013,N_16034,N_17332);
nand U19014 (N_19014,N_17025,N_16226);
nand U19015 (N_19015,N_15031,N_16145);
nor U19016 (N_19016,N_16994,N_16879);
nor U19017 (N_19017,N_15332,N_17225);
nand U19018 (N_19018,N_15090,N_15285);
nor U19019 (N_19019,N_15290,N_15928);
nand U19020 (N_19020,N_16558,N_16304);
xnor U19021 (N_19021,N_17386,N_15918);
or U19022 (N_19022,N_15619,N_16172);
nor U19023 (N_19023,N_15078,N_15144);
or U19024 (N_19024,N_17405,N_15153);
nand U19025 (N_19025,N_16959,N_15560);
or U19026 (N_19026,N_15581,N_17254);
nand U19027 (N_19027,N_15747,N_16902);
and U19028 (N_19028,N_16000,N_15111);
xor U19029 (N_19029,N_15900,N_15734);
nand U19030 (N_19030,N_16765,N_17189);
nor U19031 (N_19031,N_16512,N_15543);
or U19032 (N_19032,N_16210,N_15363);
nand U19033 (N_19033,N_16536,N_15647);
nand U19034 (N_19034,N_15209,N_16717);
nand U19035 (N_19035,N_15376,N_15067);
and U19036 (N_19036,N_15842,N_17026);
and U19037 (N_19037,N_17273,N_15501);
or U19038 (N_19038,N_17020,N_15034);
nor U19039 (N_19039,N_16904,N_16330);
and U19040 (N_19040,N_17335,N_15416);
nand U19041 (N_19041,N_16066,N_17419);
xnor U19042 (N_19042,N_15497,N_16784);
or U19043 (N_19043,N_16251,N_16772);
nor U19044 (N_19044,N_17395,N_17139);
nand U19045 (N_19045,N_15057,N_16976);
and U19046 (N_19046,N_16017,N_15048);
nand U19047 (N_19047,N_15738,N_15036);
nand U19048 (N_19048,N_16421,N_15705);
nand U19049 (N_19049,N_16553,N_16430);
and U19050 (N_19050,N_15952,N_15911);
or U19051 (N_19051,N_17190,N_17301);
nand U19052 (N_19052,N_17494,N_15640);
xor U19053 (N_19053,N_15718,N_15325);
nor U19054 (N_19054,N_15814,N_15022);
nor U19055 (N_19055,N_15839,N_15599);
or U19056 (N_19056,N_16841,N_15536);
or U19057 (N_19057,N_16751,N_15801);
nand U19058 (N_19058,N_17230,N_16784);
nor U19059 (N_19059,N_15741,N_16911);
xnor U19060 (N_19060,N_16098,N_16911);
nand U19061 (N_19061,N_16444,N_17177);
and U19062 (N_19062,N_15558,N_15144);
or U19063 (N_19063,N_17231,N_15888);
or U19064 (N_19064,N_16362,N_15820);
and U19065 (N_19065,N_15791,N_15734);
nand U19066 (N_19066,N_17302,N_15760);
and U19067 (N_19067,N_16849,N_15644);
and U19068 (N_19068,N_15385,N_16095);
nand U19069 (N_19069,N_16319,N_16956);
nor U19070 (N_19070,N_16096,N_16450);
and U19071 (N_19071,N_16568,N_15764);
nand U19072 (N_19072,N_16645,N_15975);
nor U19073 (N_19073,N_17434,N_17243);
nor U19074 (N_19074,N_15269,N_15432);
or U19075 (N_19075,N_15919,N_17055);
or U19076 (N_19076,N_15548,N_15785);
or U19077 (N_19077,N_15583,N_15883);
and U19078 (N_19078,N_16838,N_16994);
or U19079 (N_19079,N_16927,N_15133);
or U19080 (N_19080,N_15853,N_16981);
and U19081 (N_19081,N_15496,N_16945);
nand U19082 (N_19082,N_16878,N_16680);
nand U19083 (N_19083,N_15240,N_16873);
or U19084 (N_19084,N_17012,N_17371);
nor U19085 (N_19085,N_16160,N_15061);
and U19086 (N_19086,N_16933,N_15856);
nor U19087 (N_19087,N_16886,N_17025);
or U19088 (N_19088,N_17032,N_15145);
nor U19089 (N_19089,N_16610,N_15851);
nor U19090 (N_19090,N_15871,N_16562);
and U19091 (N_19091,N_16950,N_16667);
and U19092 (N_19092,N_15792,N_15533);
nand U19093 (N_19093,N_15872,N_17074);
nor U19094 (N_19094,N_16550,N_15003);
nor U19095 (N_19095,N_15740,N_16942);
and U19096 (N_19096,N_15424,N_15610);
or U19097 (N_19097,N_17154,N_17494);
or U19098 (N_19098,N_15526,N_17054);
and U19099 (N_19099,N_15173,N_16276);
nor U19100 (N_19100,N_15199,N_17116);
nor U19101 (N_19101,N_16780,N_15313);
xor U19102 (N_19102,N_17498,N_15812);
or U19103 (N_19103,N_16735,N_15180);
or U19104 (N_19104,N_15135,N_15550);
nand U19105 (N_19105,N_15163,N_16901);
or U19106 (N_19106,N_15827,N_16570);
and U19107 (N_19107,N_15722,N_17105);
or U19108 (N_19108,N_16389,N_16531);
or U19109 (N_19109,N_16503,N_15416);
nor U19110 (N_19110,N_15504,N_17309);
xnor U19111 (N_19111,N_16455,N_16055);
nor U19112 (N_19112,N_16527,N_15854);
or U19113 (N_19113,N_16063,N_16038);
nor U19114 (N_19114,N_17200,N_17034);
xor U19115 (N_19115,N_17263,N_15633);
nand U19116 (N_19116,N_17227,N_16391);
nor U19117 (N_19117,N_16279,N_15468);
nand U19118 (N_19118,N_17458,N_16104);
nand U19119 (N_19119,N_16121,N_17392);
nor U19120 (N_19120,N_15871,N_17316);
nand U19121 (N_19121,N_17378,N_16334);
or U19122 (N_19122,N_15098,N_15339);
nor U19123 (N_19123,N_17015,N_17445);
nor U19124 (N_19124,N_15844,N_15525);
nor U19125 (N_19125,N_16488,N_16279);
and U19126 (N_19126,N_16387,N_16482);
nand U19127 (N_19127,N_16888,N_15854);
nand U19128 (N_19128,N_15274,N_16802);
nand U19129 (N_19129,N_17275,N_15631);
and U19130 (N_19130,N_15969,N_16390);
nor U19131 (N_19131,N_15034,N_15487);
or U19132 (N_19132,N_15476,N_16869);
xor U19133 (N_19133,N_15495,N_17101);
or U19134 (N_19134,N_15237,N_15696);
xnor U19135 (N_19135,N_17430,N_15665);
nor U19136 (N_19136,N_17410,N_15087);
and U19137 (N_19137,N_16893,N_15867);
xnor U19138 (N_19138,N_16514,N_17077);
and U19139 (N_19139,N_16580,N_16397);
nor U19140 (N_19140,N_17160,N_15795);
nor U19141 (N_19141,N_16088,N_15134);
or U19142 (N_19142,N_15471,N_16126);
nor U19143 (N_19143,N_15815,N_17271);
or U19144 (N_19144,N_16352,N_15273);
and U19145 (N_19145,N_16533,N_15758);
or U19146 (N_19146,N_16565,N_17032);
nor U19147 (N_19147,N_16306,N_15146);
nand U19148 (N_19148,N_16929,N_17160);
nand U19149 (N_19149,N_17105,N_17284);
nor U19150 (N_19150,N_16388,N_15913);
nand U19151 (N_19151,N_15430,N_16533);
nor U19152 (N_19152,N_16383,N_16038);
and U19153 (N_19153,N_16735,N_16145);
nor U19154 (N_19154,N_15128,N_15382);
or U19155 (N_19155,N_16916,N_15357);
or U19156 (N_19156,N_15702,N_15099);
nor U19157 (N_19157,N_17412,N_16698);
and U19158 (N_19158,N_15954,N_16057);
or U19159 (N_19159,N_17018,N_15966);
nor U19160 (N_19160,N_15392,N_17429);
xnor U19161 (N_19161,N_16093,N_17011);
nor U19162 (N_19162,N_15443,N_15222);
nor U19163 (N_19163,N_15793,N_15117);
and U19164 (N_19164,N_16565,N_16300);
nor U19165 (N_19165,N_16259,N_16790);
nor U19166 (N_19166,N_16444,N_15590);
nor U19167 (N_19167,N_17209,N_16547);
nand U19168 (N_19168,N_16148,N_16998);
and U19169 (N_19169,N_16156,N_16408);
and U19170 (N_19170,N_15125,N_16960);
or U19171 (N_19171,N_16124,N_15299);
and U19172 (N_19172,N_16617,N_16960);
nor U19173 (N_19173,N_15385,N_15098);
nand U19174 (N_19174,N_15476,N_16442);
nor U19175 (N_19175,N_16129,N_16185);
and U19176 (N_19176,N_16232,N_17187);
nor U19177 (N_19177,N_15550,N_17329);
or U19178 (N_19178,N_16141,N_17320);
or U19179 (N_19179,N_17174,N_17321);
and U19180 (N_19180,N_15764,N_15654);
nand U19181 (N_19181,N_15538,N_15832);
nor U19182 (N_19182,N_16202,N_17050);
xor U19183 (N_19183,N_16501,N_15134);
or U19184 (N_19184,N_16922,N_15787);
nor U19185 (N_19185,N_16422,N_16000);
or U19186 (N_19186,N_16714,N_16038);
and U19187 (N_19187,N_15440,N_15541);
or U19188 (N_19188,N_16350,N_17223);
xnor U19189 (N_19189,N_16057,N_15158);
nand U19190 (N_19190,N_16048,N_15427);
nand U19191 (N_19191,N_16202,N_17155);
and U19192 (N_19192,N_17369,N_15123);
nand U19193 (N_19193,N_15061,N_16885);
or U19194 (N_19194,N_15493,N_16328);
nor U19195 (N_19195,N_16920,N_15711);
nor U19196 (N_19196,N_16857,N_16422);
nor U19197 (N_19197,N_15604,N_16624);
and U19198 (N_19198,N_17384,N_16873);
and U19199 (N_19199,N_16486,N_16296);
nand U19200 (N_19200,N_15021,N_15006);
nand U19201 (N_19201,N_15154,N_17031);
or U19202 (N_19202,N_16295,N_16368);
or U19203 (N_19203,N_15579,N_16340);
nand U19204 (N_19204,N_15794,N_15942);
nand U19205 (N_19205,N_17022,N_16682);
nor U19206 (N_19206,N_15843,N_15608);
and U19207 (N_19207,N_16442,N_15489);
or U19208 (N_19208,N_16476,N_16219);
nand U19209 (N_19209,N_15615,N_17095);
or U19210 (N_19210,N_17081,N_15413);
nor U19211 (N_19211,N_17042,N_15134);
xor U19212 (N_19212,N_15541,N_16865);
nand U19213 (N_19213,N_16019,N_17469);
and U19214 (N_19214,N_16095,N_16610);
nor U19215 (N_19215,N_17416,N_16625);
nand U19216 (N_19216,N_15471,N_15465);
nor U19217 (N_19217,N_15247,N_15196);
nand U19218 (N_19218,N_16322,N_16984);
or U19219 (N_19219,N_15064,N_16088);
and U19220 (N_19220,N_16054,N_16472);
and U19221 (N_19221,N_15708,N_16568);
nor U19222 (N_19222,N_17226,N_16477);
or U19223 (N_19223,N_16321,N_15416);
nand U19224 (N_19224,N_15654,N_17229);
or U19225 (N_19225,N_15852,N_17089);
or U19226 (N_19226,N_15393,N_17395);
nand U19227 (N_19227,N_16296,N_16251);
and U19228 (N_19228,N_16432,N_16179);
nand U19229 (N_19229,N_17402,N_16382);
nor U19230 (N_19230,N_15194,N_16259);
nand U19231 (N_19231,N_15103,N_16261);
or U19232 (N_19232,N_17451,N_15248);
or U19233 (N_19233,N_17323,N_17260);
or U19234 (N_19234,N_15699,N_17349);
or U19235 (N_19235,N_15676,N_15766);
nor U19236 (N_19236,N_15124,N_15094);
and U19237 (N_19237,N_16651,N_16780);
or U19238 (N_19238,N_16918,N_16640);
xnor U19239 (N_19239,N_16222,N_16622);
and U19240 (N_19240,N_16717,N_15083);
or U19241 (N_19241,N_16977,N_15497);
or U19242 (N_19242,N_16652,N_16753);
or U19243 (N_19243,N_16513,N_16009);
nor U19244 (N_19244,N_15987,N_16603);
and U19245 (N_19245,N_17238,N_16879);
nand U19246 (N_19246,N_15886,N_17042);
and U19247 (N_19247,N_15153,N_16514);
or U19248 (N_19248,N_17274,N_15736);
nor U19249 (N_19249,N_16738,N_15531);
nand U19250 (N_19250,N_16863,N_15421);
nand U19251 (N_19251,N_15971,N_17160);
nor U19252 (N_19252,N_16496,N_16478);
nor U19253 (N_19253,N_17084,N_17408);
or U19254 (N_19254,N_15605,N_16882);
nor U19255 (N_19255,N_16073,N_17011);
or U19256 (N_19256,N_15559,N_17324);
nor U19257 (N_19257,N_15233,N_16182);
nor U19258 (N_19258,N_16319,N_15147);
or U19259 (N_19259,N_15654,N_17129);
and U19260 (N_19260,N_15822,N_17469);
nor U19261 (N_19261,N_16107,N_16671);
or U19262 (N_19262,N_17005,N_16191);
nand U19263 (N_19263,N_16065,N_16888);
nor U19264 (N_19264,N_15610,N_15191);
nand U19265 (N_19265,N_16151,N_15420);
nand U19266 (N_19266,N_17061,N_15777);
or U19267 (N_19267,N_15402,N_17428);
or U19268 (N_19268,N_17254,N_17209);
xnor U19269 (N_19269,N_15784,N_17153);
xor U19270 (N_19270,N_17475,N_16904);
and U19271 (N_19271,N_16853,N_16179);
xor U19272 (N_19272,N_17210,N_15874);
nor U19273 (N_19273,N_16117,N_16751);
and U19274 (N_19274,N_17342,N_17228);
nor U19275 (N_19275,N_16615,N_16669);
nor U19276 (N_19276,N_16935,N_15529);
nand U19277 (N_19277,N_15749,N_17280);
or U19278 (N_19278,N_16472,N_15670);
and U19279 (N_19279,N_15409,N_16987);
nor U19280 (N_19280,N_17170,N_17167);
nor U19281 (N_19281,N_17292,N_15575);
or U19282 (N_19282,N_15028,N_16693);
and U19283 (N_19283,N_16443,N_15808);
or U19284 (N_19284,N_15016,N_16075);
nand U19285 (N_19285,N_16555,N_16537);
or U19286 (N_19286,N_16297,N_15501);
and U19287 (N_19287,N_15469,N_15370);
nand U19288 (N_19288,N_17242,N_16134);
xor U19289 (N_19289,N_15819,N_16903);
or U19290 (N_19290,N_15150,N_15442);
nand U19291 (N_19291,N_15290,N_15785);
nand U19292 (N_19292,N_16253,N_16006);
and U19293 (N_19293,N_16610,N_16436);
nand U19294 (N_19294,N_15297,N_16913);
and U19295 (N_19295,N_16937,N_15419);
and U19296 (N_19296,N_15557,N_15625);
or U19297 (N_19297,N_16482,N_15479);
nand U19298 (N_19298,N_15757,N_16578);
and U19299 (N_19299,N_16027,N_16924);
nor U19300 (N_19300,N_16743,N_16632);
nand U19301 (N_19301,N_16847,N_15778);
and U19302 (N_19302,N_15205,N_16994);
xor U19303 (N_19303,N_17378,N_16211);
and U19304 (N_19304,N_16836,N_16299);
nand U19305 (N_19305,N_15913,N_17222);
nand U19306 (N_19306,N_15561,N_16415);
or U19307 (N_19307,N_17210,N_15371);
xnor U19308 (N_19308,N_17428,N_17254);
or U19309 (N_19309,N_15286,N_15890);
nand U19310 (N_19310,N_15603,N_17429);
nor U19311 (N_19311,N_15242,N_15983);
nor U19312 (N_19312,N_17059,N_15326);
or U19313 (N_19313,N_16600,N_16910);
nand U19314 (N_19314,N_15664,N_15839);
or U19315 (N_19315,N_15897,N_15353);
nor U19316 (N_19316,N_17196,N_17375);
or U19317 (N_19317,N_16598,N_15370);
or U19318 (N_19318,N_17314,N_16921);
or U19319 (N_19319,N_15602,N_16907);
xor U19320 (N_19320,N_16332,N_15703);
and U19321 (N_19321,N_15593,N_15165);
nand U19322 (N_19322,N_16476,N_17284);
nand U19323 (N_19323,N_15811,N_16491);
and U19324 (N_19324,N_15980,N_16555);
nor U19325 (N_19325,N_17012,N_17412);
nor U19326 (N_19326,N_16826,N_15799);
and U19327 (N_19327,N_17367,N_15394);
nor U19328 (N_19328,N_16849,N_15693);
or U19329 (N_19329,N_15952,N_15514);
nor U19330 (N_19330,N_15567,N_15195);
nor U19331 (N_19331,N_15297,N_17342);
nor U19332 (N_19332,N_16632,N_15137);
nand U19333 (N_19333,N_15986,N_16943);
xnor U19334 (N_19334,N_15069,N_15271);
nand U19335 (N_19335,N_16926,N_17319);
nor U19336 (N_19336,N_16084,N_17320);
nor U19337 (N_19337,N_15257,N_16515);
or U19338 (N_19338,N_15956,N_16407);
nor U19339 (N_19339,N_17300,N_17330);
nand U19340 (N_19340,N_17213,N_15438);
or U19341 (N_19341,N_16764,N_16596);
nand U19342 (N_19342,N_16177,N_16735);
or U19343 (N_19343,N_15524,N_15649);
nor U19344 (N_19344,N_15176,N_16388);
nor U19345 (N_19345,N_16761,N_15247);
and U19346 (N_19346,N_17213,N_15940);
nand U19347 (N_19347,N_17420,N_16501);
nor U19348 (N_19348,N_16717,N_16571);
or U19349 (N_19349,N_17467,N_17160);
and U19350 (N_19350,N_16667,N_17412);
nor U19351 (N_19351,N_15267,N_16340);
nand U19352 (N_19352,N_16964,N_16613);
and U19353 (N_19353,N_15158,N_15185);
or U19354 (N_19354,N_16855,N_17129);
and U19355 (N_19355,N_15787,N_16835);
nor U19356 (N_19356,N_16508,N_16932);
nand U19357 (N_19357,N_15417,N_15005);
xnor U19358 (N_19358,N_16619,N_17176);
or U19359 (N_19359,N_15993,N_16133);
nand U19360 (N_19360,N_16614,N_15198);
nand U19361 (N_19361,N_16664,N_16396);
nor U19362 (N_19362,N_15167,N_16995);
or U19363 (N_19363,N_17002,N_16563);
nor U19364 (N_19364,N_15688,N_15387);
nor U19365 (N_19365,N_15802,N_16985);
and U19366 (N_19366,N_15776,N_15878);
nor U19367 (N_19367,N_16731,N_17100);
or U19368 (N_19368,N_17145,N_17335);
or U19369 (N_19369,N_15391,N_15711);
nand U19370 (N_19370,N_15384,N_16216);
nand U19371 (N_19371,N_15980,N_17487);
xor U19372 (N_19372,N_17367,N_15461);
nor U19373 (N_19373,N_17384,N_16321);
or U19374 (N_19374,N_17101,N_15739);
and U19375 (N_19375,N_17140,N_16812);
and U19376 (N_19376,N_16379,N_16780);
or U19377 (N_19377,N_15759,N_15336);
and U19378 (N_19378,N_17465,N_16297);
xor U19379 (N_19379,N_16866,N_17285);
nor U19380 (N_19380,N_15515,N_15556);
and U19381 (N_19381,N_15558,N_16276);
nand U19382 (N_19382,N_16044,N_16030);
and U19383 (N_19383,N_16846,N_16828);
nor U19384 (N_19384,N_16928,N_16228);
nor U19385 (N_19385,N_16255,N_16658);
or U19386 (N_19386,N_16113,N_15573);
nor U19387 (N_19387,N_16966,N_16163);
nand U19388 (N_19388,N_15942,N_15252);
nor U19389 (N_19389,N_17169,N_16591);
or U19390 (N_19390,N_16986,N_15299);
and U19391 (N_19391,N_15685,N_16220);
or U19392 (N_19392,N_15438,N_15371);
xnor U19393 (N_19393,N_15812,N_15607);
nor U19394 (N_19394,N_17381,N_16818);
or U19395 (N_19395,N_15909,N_16685);
nand U19396 (N_19396,N_15034,N_16455);
nor U19397 (N_19397,N_15460,N_17395);
and U19398 (N_19398,N_16470,N_16112);
or U19399 (N_19399,N_16074,N_15130);
nand U19400 (N_19400,N_15361,N_16309);
or U19401 (N_19401,N_17196,N_16285);
nor U19402 (N_19402,N_15925,N_17266);
nor U19403 (N_19403,N_17270,N_17409);
and U19404 (N_19404,N_15752,N_16695);
or U19405 (N_19405,N_16642,N_16895);
or U19406 (N_19406,N_16323,N_16899);
or U19407 (N_19407,N_17257,N_15410);
or U19408 (N_19408,N_16718,N_16449);
or U19409 (N_19409,N_15776,N_16781);
nand U19410 (N_19410,N_17316,N_16311);
nand U19411 (N_19411,N_17311,N_16512);
nand U19412 (N_19412,N_15623,N_17077);
or U19413 (N_19413,N_16196,N_16493);
nand U19414 (N_19414,N_16702,N_15637);
or U19415 (N_19415,N_16331,N_17288);
nand U19416 (N_19416,N_17207,N_17304);
and U19417 (N_19417,N_16279,N_15629);
and U19418 (N_19418,N_16387,N_17458);
nand U19419 (N_19419,N_15221,N_16265);
nand U19420 (N_19420,N_17243,N_16096);
nand U19421 (N_19421,N_17466,N_15840);
or U19422 (N_19422,N_17225,N_15351);
xnor U19423 (N_19423,N_16522,N_16083);
and U19424 (N_19424,N_16653,N_17157);
nand U19425 (N_19425,N_16147,N_16721);
nor U19426 (N_19426,N_15715,N_15621);
or U19427 (N_19427,N_15872,N_16007);
and U19428 (N_19428,N_16541,N_15661);
or U19429 (N_19429,N_15613,N_16629);
or U19430 (N_19430,N_16564,N_15469);
or U19431 (N_19431,N_16569,N_16102);
or U19432 (N_19432,N_16458,N_17306);
and U19433 (N_19433,N_15784,N_16796);
or U19434 (N_19434,N_16076,N_15891);
or U19435 (N_19435,N_15638,N_16666);
nor U19436 (N_19436,N_17292,N_16102);
nand U19437 (N_19437,N_15322,N_16297);
or U19438 (N_19438,N_15996,N_16786);
nor U19439 (N_19439,N_15637,N_17326);
or U19440 (N_19440,N_15533,N_16596);
and U19441 (N_19441,N_16469,N_16283);
nor U19442 (N_19442,N_16849,N_15852);
or U19443 (N_19443,N_16725,N_16295);
xnor U19444 (N_19444,N_15826,N_15145);
nand U19445 (N_19445,N_15095,N_16614);
nor U19446 (N_19446,N_16295,N_16573);
nor U19447 (N_19447,N_16141,N_16098);
and U19448 (N_19448,N_17040,N_15516);
nor U19449 (N_19449,N_15721,N_16049);
or U19450 (N_19450,N_16056,N_15766);
and U19451 (N_19451,N_17484,N_15279);
or U19452 (N_19452,N_17017,N_17263);
nand U19453 (N_19453,N_15828,N_16191);
nor U19454 (N_19454,N_15724,N_17203);
nor U19455 (N_19455,N_16689,N_16458);
nor U19456 (N_19456,N_16402,N_15051);
and U19457 (N_19457,N_15008,N_17431);
and U19458 (N_19458,N_16909,N_16872);
and U19459 (N_19459,N_15091,N_15059);
or U19460 (N_19460,N_15283,N_15140);
or U19461 (N_19461,N_15751,N_15099);
or U19462 (N_19462,N_17369,N_16568);
nor U19463 (N_19463,N_15216,N_16154);
and U19464 (N_19464,N_15425,N_15534);
and U19465 (N_19465,N_17248,N_15169);
nor U19466 (N_19466,N_15987,N_15325);
nor U19467 (N_19467,N_15247,N_15781);
or U19468 (N_19468,N_16956,N_16217);
or U19469 (N_19469,N_15326,N_15946);
nand U19470 (N_19470,N_15982,N_15571);
nand U19471 (N_19471,N_17075,N_15494);
xor U19472 (N_19472,N_15136,N_17340);
nor U19473 (N_19473,N_17477,N_16165);
or U19474 (N_19474,N_17090,N_15945);
nor U19475 (N_19475,N_16917,N_16349);
nor U19476 (N_19476,N_15554,N_17460);
or U19477 (N_19477,N_15407,N_17087);
and U19478 (N_19478,N_16197,N_16149);
nand U19479 (N_19479,N_16964,N_16021);
nor U19480 (N_19480,N_15160,N_16667);
and U19481 (N_19481,N_15015,N_16996);
and U19482 (N_19482,N_15123,N_16647);
nor U19483 (N_19483,N_16168,N_15175);
nand U19484 (N_19484,N_17176,N_16841);
and U19485 (N_19485,N_16419,N_15327);
xnor U19486 (N_19486,N_15290,N_17200);
and U19487 (N_19487,N_17288,N_16794);
and U19488 (N_19488,N_15189,N_17216);
nor U19489 (N_19489,N_16921,N_17101);
nor U19490 (N_19490,N_15631,N_16962);
and U19491 (N_19491,N_16568,N_16647);
nor U19492 (N_19492,N_15622,N_15442);
or U19493 (N_19493,N_16355,N_16966);
nor U19494 (N_19494,N_17413,N_15033);
or U19495 (N_19495,N_15227,N_15699);
or U19496 (N_19496,N_16091,N_16458);
and U19497 (N_19497,N_16130,N_16795);
nor U19498 (N_19498,N_17482,N_15383);
and U19499 (N_19499,N_17018,N_15954);
nor U19500 (N_19500,N_16398,N_16816);
nor U19501 (N_19501,N_16143,N_16405);
or U19502 (N_19502,N_17417,N_16812);
nor U19503 (N_19503,N_15681,N_17142);
nand U19504 (N_19504,N_16253,N_16592);
nand U19505 (N_19505,N_15726,N_15880);
and U19506 (N_19506,N_17201,N_15965);
or U19507 (N_19507,N_16074,N_17027);
nor U19508 (N_19508,N_17485,N_16572);
and U19509 (N_19509,N_16413,N_16837);
and U19510 (N_19510,N_17316,N_15519);
or U19511 (N_19511,N_15718,N_16746);
xor U19512 (N_19512,N_15158,N_16324);
and U19513 (N_19513,N_17071,N_15758);
nand U19514 (N_19514,N_15029,N_15760);
or U19515 (N_19515,N_17110,N_17467);
or U19516 (N_19516,N_16112,N_15274);
nand U19517 (N_19517,N_17368,N_17322);
and U19518 (N_19518,N_16138,N_15323);
or U19519 (N_19519,N_17451,N_15867);
and U19520 (N_19520,N_15607,N_16475);
and U19521 (N_19521,N_17483,N_15315);
nand U19522 (N_19522,N_15070,N_17123);
nand U19523 (N_19523,N_16128,N_16585);
nand U19524 (N_19524,N_15885,N_16501);
nor U19525 (N_19525,N_16751,N_15669);
nor U19526 (N_19526,N_16468,N_15800);
nand U19527 (N_19527,N_16653,N_15773);
nor U19528 (N_19528,N_16365,N_17223);
and U19529 (N_19529,N_15387,N_17257);
xnor U19530 (N_19530,N_15380,N_16188);
nand U19531 (N_19531,N_15256,N_17498);
and U19532 (N_19532,N_17040,N_16772);
and U19533 (N_19533,N_16658,N_16836);
and U19534 (N_19534,N_15500,N_15381);
nor U19535 (N_19535,N_15012,N_15403);
or U19536 (N_19536,N_15885,N_16134);
nand U19537 (N_19537,N_15307,N_16564);
nor U19538 (N_19538,N_15439,N_16931);
nor U19539 (N_19539,N_17396,N_17372);
xnor U19540 (N_19540,N_17075,N_17323);
xnor U19541 (N_19541,N_16337,N_16106);
nor U19542 (N_19542,N_16127,N_15175);
and U19543 (N_19543,N_17324,N_16079);
xnor U19544 (N_19544,N_16916,N_17071);
nor U19545 (N_19545,N_17441,N_15762);
or U19546 (N_19546,N_16314,N_15296);
xor U19547 (N_19547,N_15635,N_15803);
or U19548 (N_19548,N_15079,N_16846);
xnor U19549 (N_19549,N_15816,N_16843);
and U19550 (N_19550,N_15221,N_16694);
or U19551 (N_19551,N_16467,N_15971);
or U19552 (N_19552,N_17423,N_15902);
xor U19553 (N_19553,N_17143,N_15700);
and U19554 (N_19554,N_16787,N_17164);
and U19555 (N_19555,N_16166,N_17300);
nand U19556 (N_19556,N_16458,N_15457);
or U19557 (N_19557,N_15233,N_17071);
xnor U19558 (N_19558,N_15659,N_17245);
and U19559 (N_19559,N_16010,N_15322);
nor U19560 (N_19560,N_15363,N_16884);
nand U19561 (N_19561,N_17042,N_15936);
or U19562 (N_19562,N_17455,N_15271);
or U19563 (N_19563,N_15391,N_15911);
nor U19564 (N_19564,N_15894,N_15962);
nor U19565 (N_19565,N_15945,N_16817);
nor U19566 (N_19566,N_15883,N_15990);
nor U19567 (N_19567,N_15619,N_17040);
nor U19568 (N_19568,N_15446,N_16793);
and U19569 (N_19569,N_16086,N_16087);
xor U19570 (N_19570,N_15971,N_17389);
or U19571 (N_19571,N_15163,N_16021);
and U19572 (N_19572,N_17480,N_15222);
nor U19573 (N_19573,N_16808,N_16194);
nand U19574 (N_19574,N_16385,N_16533);
nand U19575 (N_19575,N_16820,N_15396);
nand U19576 (N_19576,N_15132,N_16950);
and U19577 (N_19577,N_17026,N_15894);
or U19578 (N_19578,N_17463,N_15044);
or U19579 (N_19579,N_16199,N_15752);
nor U19580 (N_19580,N_17331,N_15864);
or U19581 (N_19581,N_15526,N_16035);
nand U19582 (N_19582,N_16790,N_15542);
nand U19583 (N_19583,N_16257,N_15146);
nor U19584 (N_19584,N_15187,N_17285);
and U19585 (N_19585,N_15610,N_15133);
or U19586 (N_19586,N_16242,N_15590);
nor U19587 (N_19587,N_16384,N_15664);
nand U19588 (N_19588,N_17456,N_16793);
nand U19589 (N_19589,N_15829,N_15288);
or U19590 (N_19590,N_15559,N_15582);
and U19591 (N_19591,N_15399,N_16243);
nand U19592 (N_19592,N_15126,N_15496);
or U19593 (N_19593,N_15520,N_15202);
and U19594 (N_19594,N_16325,N_16571);
nand U19595 (N_19595,N_16741,N_17409);
and U19596 (N_19596,N_15965,N_16095);
or U19597 (N_19597,N_16379,N_16032);
nand U19598 (N_19598,N_17442,N_15268);
or U19599 (N_19599,N_15685,N_16881);
and U19600 (N_19600,N_16349,N_17340);
nor U19601 (N_19601,N_16528,N_15636);
and U19602 (N_19602,N_16917,N_15769);
nand U19603 (N_19603,N_16619,N_16859);
and U19604 (N_19604,N_16543,N_16289);
and U19605 (N_19605,N_15527,N_17222);
and U19606 (N_19606,N_15229,N_16108);
nor U19607 (N_19607,N_16577,N_16538);
or U19608 (N_19608,N_16139,N_17450);
nor U19609 (N_19609,N_15846,N_15301);
xnor U19610 (N_19610,N_15331,N_15323);
xor U19611 (N_19611,N_15673,N_16130);
and U19612 (N_19612,N_16396,N_16372);
nor U19613 (N_19613,N_17104,N_16596);
or U19614 (N_19614,N_17034,N_15556);
or U19615 (N_19615,N_15817,N_17436);
or U19616 (N_19616,N_17328,N_15096);
or U19617 (N_19617,N_16258,N_16239);
nand U19618 (N_19618,N_15411,N_17350);
xor U19619 (N_19619,N_15917,N_16494);
nor U19620 (N_19620,N_16173,N_15643);
or U19621 (N_19621,N_15771,N_15502);
or U19622 (N_19622,N_16331,N_16618);
nand U19623 (N_19623,N_17474,N_15026);
nor U19624 (N_19624,N_15367,N_16806);
and U19625 (N_19625,N_16158,N_16577);
or U19626 (N_19626,N_17292,N_16034);
nor U19627 (N_19627,N_15036,N_16622);
and U19628 (N_19628,N_15369,N_17266);
nand U19629 (N_19629,N_16652,N_16945);
or U19630 (N_19630,N_16736,N_15714);
and U19631 (N_19631,N_17277,N_15403);
xnor U19632 (N_19632,N_15096,N_15746);
nor U19633 (N_19633,N_16572,N_15926);
nand U19634 (N_19634,N_16466,N_15635);
or U19635 (N_19635,N_16307,N_15631);
and U19636 (N_19636,N_16522,N_16143);
or U19637 (N_19637,N_15880,N_16143);
nor U19638 (N_19638,N_16494,N_17489);
nand U19639 (N_19639,N_16076,N_16910);
nor U19640 (N_19640,N_16896,N_17137);
or U19641 (N_19641,N_17164,N_15130);
xnor U19642 (N_19642,N_16455,N_15830);
or U19643 (N_19643,N_16679,N_16127);
nor U19644 (N_19644,N_15624,N_16487);
xnor U19645 (N_19645,N_16446,N_16416);
nand U19646 (N_19646,N_16212,N_16812);
nand U19647 (N_19647,N_15453,N_15002);
nand U19648 (N_19648,N_17026,N_15299);
xor U19649 (N_19649,N_17391,N_15334);
nor U19650 (N_19650,N_16056,N_15103);
nand U19651 (N_19651,N_17256,N_17177);
xor U19652 (N_19652,N_15523,N_16985);
or U19653 (N_19653,N_16399,N_16565);
and U19654 (N_19654,N_15503,N_16002);
or U19655 (N_19655,N_17340,N_15984);
nor U19656 (N_19656,N_17384,N_16215);
xnor U19657 (N_19657,N_15022,N_15849);
or U19658 (N_19658,N_15747,N_15525);
nand U19659 (N_19659,N_15867,N_15349);
or U19660 (N_19660,N_15122,N_15341);
or U19661 (N_19661,N_15592,N_16932);
nand U19662 (N_19662,N_15661,N_15371);
xnor U19663 (N_19663,N_17441,N_15347);
or U19664 (N_19664,N_15710,N_15780);
nor U19665 (N_19665,N_16054,N_16033);
and U19666 (N_19666,N_17244,N_16715);
nand U19667 (N_19667,N_15895,N_16735);
nor U19668 (N_19668,N_15907,N_16284);
and U19669 (N_19669,N_17189,N_15618);
and U19670 (N_19670,N_16493,N_17020);
xnor U19671 (N_19671,N_15278,N_17374);
and U19672 (N_19672,N_17437,N_16708);
or U19673 (N_19673,N_15890,N_16158);
nand U19674 (N_19674,N_16745,N_16697);
nor U19675 (N_19675,N_16236,N_17153);
nor U19676 (N_19676,N_16605,N_16148);
or U19677 (N_19677,N_15459,N_15637);
nor U19678 (N_19678,N_16170,N_17451);
xnor U19679 (N_19679,N_17262,N_15081);
nand U19680 (N_19680,N_16154,N_15918);
xor U19681 (N_19681,N_15792,N_15375);
nand U19682 (N_19682,N_16932,N_15660);
xor U19683 (N_19683,N_17037,N_16838);
xnor U19684 (N_19684,N_16244,N_15774);
and U19685 (N_19685,N_16110,N_16575);
nor U19686 (N_19686,N_16399,N_15643);
nand U19687 (N_19687,N_15054,N_15640);
or U19688 (N_19688,N_16207,N_15604);
nand U19689 (N_19689,N_15225,N_16254);
or U19690 (N_19690,N_15364,N_16224);
nor U19691 (N_19691,N_15879,N_16572);
nor U19692 (N_19692,N_17417,N_15234);
nand U19693 (N_19693,N_16240,N_16948);
nand U19694 (N_19694,N_16732,N_17497);
nor U19695 (N_19695,N_15943,N_17378);
and U19696 (N_19696,N_16347,N_15135);
nand U19697 (N_19697,N_16941,N_17054);
and U19698 (N_19698,N_16339,N_16617);
or U19699 (N_19699,N_17041,N_16628);
and U19700 (N_19700,N_16966,N_17378);
nand U19701 (N_19701,N_15370,N_15382);
or U19702 (N_19702,N_17256,N_16072);
or U19703 (N_19703,N_15030,N_16555);
nand U19704 (N_19704,N_15401,N_17028);
and U19705 (N_19705,N_16261,N_16927);
xor U19706 (N_19706,N_17249,N_16167);
xor U19707 (N_19707,N_15854,N_17399);
xor U19708 (N_19708,N_17470,N_15923);
nand U19709 (N_19709,N_15623,N_15855);
and U19710 (N_19710,N_17130,N_15148);
and U19711 (N_19711,N_15862,N_16951);
nand U19712 (N_19712,N_15316,N_16843);
or U19713 (N_19713,N_15371,N_15685);
nand U19714 (N_19714,N_17395,N_16366);
nor U19715 (N_19715,N_15416,N_16664);
nor U19716 (N_19716,N_17335,N_15848);
and U19717 (N_19717,N_16046,N_15325);
xor U19718 (N_19718,N_16645,N_16607);
nor U19719 (N_19719,N_15504,N_15115);
nor U19720 (N_19720,N_15972,N_15391);
or U19721 (N_19721,N_15236,N_16579);
or U19722 (N_19722,N_16420,N_16440);
xor U19723 (N_19723,N_16281,N_17474);
and U19724 (N_19724,N_16865,N_17191);
nor U19725 (N_19725,N_17365,N_15869);
xnor U19726 (N_19726,N_15742,N_15839);
nand U19727 (N_19727,N_15741,N_15602);
nor U19728 (N_19728,N_15080,N_16811);
and U19729 (N_19729,N_16325,N_15518);
and U19730 (N_19730,N_15564,N_17087);
nor U19731 (N_19731,N_16484,N_15621);
nor U19732 (N_19732,N_16626,N_15748);
nor U19733 (N_19733,N_17124,N_16492);
nor U19734 (N_19734,N_17140,N_17150);
nand U19735 (N_19735,N_15316,N_15383);
nand U19736 (N_19736,N_16943,N_17173);
nand U19737 (N_19737,N_16924,N_16822);
nor U19738 (N_19738,N_17306,N_15567);
and U19739 (N_19739,N_15987,N_16947);
nand U19740 (N_19740,N_15675,N_17199);
and U19741 (N_19741,N_15546,N_15500);
nor U19742 (N_19742,N_16183,N_16411);
and U19743 (N_19743,N_16664,N_15410);
or U19744 (N_19744,N_15018,N_16845);
or U19745 (N_19745,N_17394,N_16538);
or U19746 (N_19746,N_17025,N_16334);
or U19747 (N_19747,N_17409,N_17135);
nand U19748 (N_19748,N_17115,N_16171);
nor U19749 (N_19749,N_15620,N_16860);
nand U19750 (N_19750,N_16179,N_16815);
or U19751 (N_19751,N_17492,N_15568);
nand U19752 (N_19752,N_15043,N_15073);
or U19753 (N_19753,N_17263,N_16377);
nand U19754 (N_19754,N_15737,N_16860);
nor U19755 (N_19755,N_15396,N_16167);
or U19756 (N_19756,N_15273,N_17022);
or U19757 (N_19757,N_16738,N_16498);
nor U19758 (N_19758,N_17093,N_16141);
nor U19759 (N_19759,N_16849,N_16888);
nand U19760 (N_19760,N_16183,N_16968);
nor U19761 (N_19761,N_15929,N_15801);
nand U19762 (N_19762,N_15634,N_16895);
or U19763 (N_19763,N_15921,N_17465);
nor U19764 (N_19764,N_16531,N_16924);
or U19765 (N_19765,N_16533,N_15795);
nand U19766 (N_19766,N_16447,N_16745);
nor U19767 (N_19767,N_17215,N_16252);
nand U19768 (N_19768,N_17292,N_16028);
or U19769 (N_19769,N_15983,N_17123);
xnor U19770 (N_19770,N_15335,N_16970);
nor U19771 (N_19771,N_16979,N_16790);
nor U19772 (N_19772,N_16232,N_15500);
nand U19773 (N_19773,N_15558,N_16611);
nor U19774 (N_19774,N_15747,N_15038);
or U19775 (N_19775,N_15192,N_16113);
nor U19776 (N_19776,N_17142,N_16868);
nor U19777 (N_19777,N_16168,N_15300);
or U19778 (N_19778,N_16631,N_15860);
nor U19779 (N_19779,N_16262,N_17216);
nor U19780 (N_19780,N_16135,N_17040);
or U19781 (N_19781,N_16460,N_16807);
and U19782 (N_19782,N_15800,N_16891);
nor U19783 (N_19783,N_17463,N_15133);
nor U19784 (N_19784,N_16047,N_15923);
and U19785 (N_19785,N_16787,N_15137);
or U19786 (N_19786,N_16616,N_15699);
or U19787 (N_19787,N_16593,N_15729);
or U19788 (N_19788,N_16922,N_16488);
or U19789 (N_19789,N_16629,N_16260);
or U19790 (N_19790,N_17061,N_16206);
nand U19791 (N_19791,N_15544,N_15488);
nand U19792 (N_19792,N_17028,N_16145);
nor U19793 (N_19793,N_15054,N_17416);
nor U19794 (N_19794,N_16102,N_16290);
or U19795 (N_19795,N_15782,N_17251);
and U19796 (N_19796,N_15954,N_15730);
or U19797 (N_19797,N_15352,N_16474);
nor U19798 (N_19798,N_17047,N_15127);
or U19799 (N_19799,N_15365,N_15357);
nand U19800 (N_19800,N_16412,N_16391);
and U19801 (N_19801,N_17193,N_16717);
and U19802 (N_19802,N_16250,N_16410);
and U19803 (N_19803,N_15885,N_15376);
or U19804 (N_19804,N_16558,N_16985);
nand U19805 (N_19805,N_16526,N_16789);
and U19806 (N_19806,N_16116,N_16348);
nor U19807 (N_19807,N_15667,N_15027);
and U19808 (N_19808,N_16876,N_16520);
or U19809 (N_19809,N_15534,N_17162);
or U19810 (N_19810,N_16911,N_15608);
and U19811 (N_19811,N_16719,N_17370);
or U19812 (N_19812,N_17344,N_15618);
nor U19813 (N_19813,N_17220,N_16795);
nand U19814 (N_19814,N_15018,N_17191);
xnor U19815 (N_19815,N_15691,N_16907);
xnor U19816 (N_19816,N_15679,N_15590);
or U19817 (N_19817,N_16744,N_15513);
or U19818 (N_19818,N_16818,N_16141);
xnor U19819 (N_19819,N_16859,N_16308);
xor U19820 (N_19820,N_16159,N_16248);
and U19821 (N_19821,N_17353,N_16078);
or U19822 (N_19822,N_16145,N_16219);
or U19823 (N_19823,N_15423,N_15298);
nor U19824 (N_19824,N_16981,N_15140);
xnor U19825 (N_19825,N_16343,N_15706);
nand U19826 (N_19826,N_16518,N_17498);
and U19827 (N_19827,N_15314,N_16601);
xor U19828 (N_19828,N_15928,N_15732);
nand U19829 (N_19829,N_16270,N_17364);
and U19830 (N_19830,N_15753,N_15819);
and U19831 (N_19831,N_16159,N_15024);
nor U19832 (N_19832,N_16654,N_15855);
nand U19833 (N_19833,N_16743,N_17247);
nand U19834 (N_19834,N_15796,N_15909);
or U19835 (N_19835,N_16633,N_16520);
nor U19836 (N_19836,N_16463,N_16700);
or U19837 (N_19837,N_17180,N_15105);
nor U19838 (N_19838,N_15482,N_15224);
or U19839 (N_19839,N_15694,N_16985);
nand U19840 (N_19840,N_15433,N_15581);
nand U19841 (N_19841,N_16509,N_16073);
nor U19842 (N_19842,N_15707,N_15933);
xor U19843 (N_19843,N_16060,N_16632);
nand U19844 (N_19844,N_15907,N_17246);
and U19845 (N_19845,N_15985,N_15016);
nand U19846 (N_19846,N_15914,N_15993);
and U19847 (N_19847,N_15905,N_16661);
nor U19848 (N_19848,N_16328,N_15061);
nand U19849 (N_19849,N_15698,N_16867);
nand U19850 (N_19850,N_15585,N_17215);
nand U19851 (N_19851,N_15717,N_16150);
nand U19852 (N_19852,N_17368,N_15408);
or U19853 (N_19853,N_15860,N_15501);
or U19854 (N_19854,N_15698,N_16357);
and U19855 (N_19855,N_16396,N_16340);
and U19856 (N_19856,N_16293,N_15029);
or U19857 (N_19857,N_15945,N_16286);
xnor U19858 (N_19858,N_17187,N_17462);
nor U19859 (N_19859,N_16933,N_17198);
xor U19860 (N_19860,N_17020,N_17093);
nor U19861 (N_19861,N_15343,N_16627);
and U19862 (N_19862,N_15499,N_15634);
nand U19863 (N_19863,N_15999,N_16812);
nand U19864 (N_19864,N_16627,N_15931);
nand U19865 (N_19865,N_16758,N_16222);
and U19866 (N_19866,N_16048,N_15849);
and U19867 (N_19867,N_16491,N_16317);
and U19868 (N_19868,N_16897,N_15336);
nand U19869 (N_19869,N_16294,N_16359);
nand U19870 (N_19870,N_17448,N_16802);
and U19871 (N_19871,N_17289,N_15725);
and U19872 (N_19872,N_17007,N_16464);
or U19873 (N_19873,N_16117,N_16668);
nor U19874 (N_19874,N_17374,N_17199);
and U19875 (N_19875,N_17297,N_17448);
or U19876 (N_19876,N_15389,N_16309);
nand U19877 (N_19877,N_16705,N_15625);
nor U19878 (N_19878,N_17178,N_16839);
and U19879 (N_19879,N_16524,N_16937);
xnor U19880 (N_19880,N_15855,N_16056);
nor U19881 (N_19881,N_15914,N_17093);
or U19882 (N_19882,N_17376,N_16315);
and U19883 (N_19883,N_15773,N_17492);
and U19884 (N_19884,N_16815,N_16346);
nand U19885 (N_19885,N_16387,N_15324);
or U19886 (N_19886,N_15169,N_17019);
nor U19887 (N_19887,N_15510,N_15794);
nand U19888 (N_19888,N_17142,N_16482);
or U19889 (N_19889,N_16084,N_15058);
nand U19890 (N_19890,N_16264,N_15649);
xnor U19891 (N_19891,N_17064,N_15396);
and U19892 (N_19892,N_16429,N_16879);
nor U19893 (N_19893,N_17060,N_15025);
xnor U19894 (N_19894,N_17287,N_16092);
and U19895 (N_19895,N_15131,N_16203);
and U19896 (N_19896,N_17058,N_15550);
or U19897 (N_19897,N_15333,N_16813);
nand U19898 (N_19898,N_15497,N_16165);
or U19899 (N_19899,N_15652,N_15817);
nand U19900 (N_19900,N_17064,N_16932);
nor U19901 (N_19901,N_15606,N_15121);
nand U19902 (N_19902,N_15272,N_16426);
xnor U19903 (N_19903,N_16690,N_15543);
and U19904 (N_19904,N_15355,N_15698);
and U19905 (N_19905,N_17161,N_15050);
and U19906 (N_19906,N_16994,N_16439);
and U19907 (N_19907,N_17357,N_16858);
or U19908 (N_19908,N_16104,N_17070);
nand U19909 (N_19909,N_15403,N_15247);
nor U19910 (N_19910,N_17311,N_16100);
and U19911 (N_19911,N_15747,N_15690);
nand U19912 (N_19912,N_17483,N_16081);
and U19913 (N_19913,N_15395,N_16408);
nand U19914 (N_19914,N_15769,N_15521);
and U19915 (N_19915,N_16379,N_15037);
and U19916 (N_19916,N_16783,N_16935);
nand U19917 (N_19917,N_16436,N_15764);
nand U19918 (N_19918,N_15556,N_16381);
and U19919 (N_19919,N_17124,N_16202);
or U19920 (N_19920,N_16831,N_16494);
and U19921 (N_19921,N_15425,N_16006);
and U19922 (N_19922,N_16613,N_15603);
and U19923 (N_19923,N_16607,N_16115);
nand U19924 (N_19924,N_15222,N_15099);
nor U19925 (N_19925,N_15012,N_16881);
nor U19926 (N_19926,N_17217,N_16827);
nand U19927 (N_19927,N_17327,N_16249);
or U19928 (N_19928,N_16358,N_15403);
and U19929 (N_19929,N_15542,N_15109);
and U19930 (N_19930,N_16517,N_17471);
nand U19931 (N_19931,N_17185,N_15323);
and U19932 (N_19932,N_15638,N_16396);
and U19933 (N_19933,N_16224,N_16789);
and U19934 (N_19934,N_16613,N_16115);
nand U19935 (N_19935,N_17455,N_16158);
or U19936 (N_19936,N_15619,N_16819);
xor U19937 (N_19937,N_16486,N_15634);
nand U19938 (N_19938,N_15033,N_16916);
or U19939 (N_19939,N_16725,N_15321);
nand U19940 (N_19940,N_17401,N_16014);
nor U19941 (N_19941,N_15640,N_17128);
or U19942 (N_19942,N_17272,N_16980);
or U19943 (N_19943,N_16317,N_16807);
xnor U19944 (N_19944,N_16414,N_15371);
nand U19945 (N_19945,N_16702,N_15885);
or U19946 (N_19946,N_15648,N_16706);
nor U19947 (N_19947,N_16173,N_15541);
nor U19948 (N_19948,N_16482,N_16138);
nand U19949 (N_19949,N_17028,N_16397);
nor U19950 (N_19950,N_16392,N_16417);
nor U19951 (N_19951,N_16454,N_17235);
nor U19952 (N_19952,N_15763,N_16787);
nor U19953 (N_19953,N_17372,N_15775);
xor U19954 (N_19954,N_15835,N_17026);
nand U19955 (N_19955,N_16570,N_17294);
nor U19956 (N_19956,N_15314,N_15442);
nor U19957 (N_19957,N_15716,N_15528);
and U19958 (N_19958,N_15305,N_16944);
xnor U19959 (N_19959,N_17430,N_17433);
and U19960 (N_19960,N_16470,N_16157);
and U19961 (N_19961,N_15845,N_16122);
nor U19962 (N_19962,N_15326,N_16640);
nor U19963 (N_19963,N_15728,N_15088);
and U19964 (N_19964,N_16235,N_16189);
and U19965 (N_19965,N_15079,N_15792);
nand U19966 (N_19966,N_16268,N_15137);
nor U19967 (N_19967,N_16867,N_17238);
nand U19968 (N_19968,N_15095,N_17342);
and U19969 (N_19969,N_17347,N_15564);
nor U19970 (N_19970,N_16818,N_16203);
and U19971 (N_19971,N_16745,N_16460);
nand U19972 (N_19972,N_15529,N_15177);
and U19973 (N_19973,N_16182,N_15717);
nand U19974 (N_19974,N_17300,N_16835);
and U19975 (N_19975,N_16703,N_15219);
or U19976 (N_19976,N_15632,N_15151);
and U19977 (N_19977,N_16585,N_15290);
and U19978 (N_19978,N_16890,N_16578);
nand U19979 (N_19979,N_17007,N_16002);
nand U19980 (N_19980,N_16386,N_17131);
nand U19981 (N_19981,N_17444,N_15530);
and U19982 (N_19982,N_15673,N_15349);
nand U19983 (N_19983,N_15264,N_16459);
or U19984 (N_19984,N_16662,N_16129);
nor U19985 (N_19985,N_17044,N_15575);
or U19986 (N_19986,N_15961,N_16690);
or U19987 (N_19987,N_15787,N_17298);
nor U19988 (N_19988,N_17380,N_15875);
nor U19989 (N_19989,N_15221,N_15463);
or U19990 (N_19990,N_15507,N_16294);
and U19991 (N_19991,N_15679,N_15055);
xor U19992 (N_19992,N_15573,N_15410);
nor U19993 (N_19993,N_15061,N_16737);
xor U19994 (N_19994,N_16779,N_16162);
xnor U19995 (N_19995,N_15762,N_16233);
or U19996 (N_19996,N_17367,N_16618);
nand U19997 (N_19997,N_16076,N_17044);
xnor U19998 (N_19998,N_15056,N_16787);
or U19999 (N_19999,N_15675,N_17198);
or U20000 (N_20000,N_18848,N_17566);
nand U20001 (N_20001,N_19204,N_18511);
nor U20002 (N_20002,N_18075,N_17836);
nor U20003 (N_20003,N_17998,N_19459);
nand U20004 (N_20004,N_18351,N_17701);
nand U20005 (N_20005,N_17588,N_19071);
and U20006 (N_20006,N_19480,N_18258);
or U20007 (N_20007,N_18913,N_19721);
xor U20008 (N_20008,N_17586,N_19093);
nand U20009 (N_20009,N_19696,N_18325);
or U20010 (N_20010,N_17983,N_17709);
and U20011 (N_20011,N_18694,N_17605);
nor U20012 (N_20012,N_19416,N_18000);
nor U20013 (N_20013,N_19560,N_19143);
nor U20014 (N_20014,N_18407,N_18699);
or U20015 (N_20015,N_18425,N_18763);
nor U20016 (N_20016,N_18376,N_17662);
nor U20017 (N_20017,N_19491,N_18235);
or U20018 (N_20018,N_19965,N_19487);
nand U20019 (N_20019,N_19021,N_18459);
and U20020 (N_20020,N_18035,N_19177);
or U20021 (N_20021,N_19938,N_18536);
nand U20022 (N_20022,N_19354,N_18462);
and U20023 (N_20023,N_17890,N_19345);
nand U20024 (N_20024,N_18573,N_19181);
or U20025 (N_20025,N_18179,N_18401);
and U20026 (N_20026,N_18271,N_18309);
nor U20027 (N_20027,N_18305,N_18321);
xor U20028 (N_20028,N_19090,N_19189);
nor U20029 (N_20029,N_18787,N_19078);
xor U20030 (N_20030,N_18803,N_18116);
or U20031 (N_20031,N_19474,N_17914);
or U20032 (N_20032,N_19584,N_17885);
or U20033 (N_20033,N_19170,N_18361);
and U20034 (N_20034,N_18941,N_17531);
or U20035 (N_20035,N_18284,N_19147);
nand U20036 (N_20036,N_18302,N_18864);
and U20037 (N_20037,N_18624,N_17827);
and U20038 (N_20038,N_19278,N_19771);
xor U20039 (N_20039,N_17667,N_19044);
nor U20040 (N_20040,N_18051,N_18426);
nand U20041 (N_20041,N_19984,N_18731);
or U20042 (N_20042,N_18532,N_19522);
xnor U20043 (N_20043,N_17535,N_18147);
nor U20044 (N_20044,N_17670,N_18703);
or U20045 (N_20045,N_18835,N_18533);
xor U20046 (N_20046,N_19464,N_17769);
and U20047 (N_20047,N_18831,N_17750);
nand U20048 (N_20048,N_17600,N_17934);
nand U20049 (N_20049,N_18087,N_19113);
xor U20050 (N_20050,N_17894,N_19850);
or U20051 (N_20051,N_19698,N_18571);
or U20052 (N_20052,N_17778,N_19551);
nor U20053 (N_20053,N_17919,N_19971);
and U20054 (N_20054,N_19864,N_19081);
or U20055 (N_20055,N_18754,N_18828);
and U20056 (N_20056,N_19267,N_19695);
nor U20057 (N_20057,N_19663,N_18987);
or U20058 (N_20058,N_18945,N_19558);
nor U20059 (N_20059,N_18278,N_18254);
or U20060 (N_20060,N_18454,N_17755);
or U20061 (N_20061,N_17892,N_19532);
nor U20062 (N_20062,N_17936,N_18950);
or U20063 (N_20063,N_18995,N_18193);
nand U20064 (N_20064,N_19132,N_19748);
and U20065 (N_20065,N_17607,N_19219);
nor U20066 (N_20066,N_18553,N_19228);
and U20067 (N_20067,N_19401,N_18349);
xor U20068 (N_20068,N_19791,N_19571);
nor U20069 (N_20069,N_19383,N_19531);
or U20070 (N_20070,N_19272,N_18921);
nand U20071 (N_20071,N_19035,N_18496);
and U20072 (N_20072,N_18198,N_19307);
or U20073 (N_20073,N_18209,N_19066);
nand U20074 (N_20074,N_19207,N_17813);
and U20075 (N_20075,N_19392,N_19171);
or U20076 (N_20076,N_19706,N_19178);
or U20077 (N_20077,N_18617,N_18839);
or U20078 (N_20078,N_17632,N_19646);
or U20079 (N_20079,N_18634,N_18974);
nor U20080 (N_20080,N_18800,N_19167);
nand U20081 (N_20081,N_18140,N_17807);
and U20082 (N_20082,N_18970,N_17805);
nor U20083 (N_20083,N_18919,N_18282);
nand U20084 (N_20084,N_19585,N_19039);
nor U20085 (N_20085,N_18001,N_18976);
xnor U20086 (N_20086,N_18447,N_18393);
nor U20087 (N_20087,N_17939,N_19277);
and U20088 (N_20088,N_19175,N_19588);
xnor U20089 (N_20089,N_18679,N_18312);
or U20090 (N_20090,N_18888,N_19719);
xnor U20091 (N_20091,N_18324,N_17528);
nand U20092 (N_20092,N_19820,N_18547);
nand U20093 (N_20093,N_19319,N_17958);
nand U20094 (N_20094,N_19273,N_19340);
or U20095 (N_20095,N_19376,N_19570);
or U20096 (N_20096,N_19947,N_19854);
nand U20097 (N_20097,N_18266,N_19155);
nand U20098 (N_20098,N_19783,N_19727);
nand U20099 (N_20099,N_19431,N_17513);
or U20100 (N_20100,N_18063,N_18755);
nand U20101 (N_20101,N_18236,N_17689);
nand U20102 (N_20102,N_17694,N_18172);
nor U20103 (N_20103,N_18287,N_17738);
nor U20104 (N_20104,N_19420,N_18643);
xnor U20105 (N_20105,N_18636,N_17754);
nor U20106 (N_20106,N_18390,N_19036);
nor U20107 (N_20107,N_19242,N_18957);
nand U20108 (N_20108,N_18182,N_18940);
nand U20109 (N_20109,N_19765,N_18036);
nor U20110 (N_20110,N_19799,N_18315);
or U20111 (N_20111,N_18463,N_18473);
xnor U20112 (N_20112,N_17516,N_19598);
and U20113 (N_20113,N_18242,N_17906);
and U20114 (N_20114,N_19789,N_19003);
nand U20115 (N_20115,N_18181,N_18263);
nand U20116 (N_20116,N_18444,N_19438);
and U20117 (N_20117,N_18389,N_19852);
nand U20118 (N_20118,N_19573,N_18827);
xor U20119 (N_20119,N_18613,N_17596);
or U20120 (N_20120,N_18489,N_18227);
or U20121 (N_20121,N_18412,N_18470);
nor U20122 (N_20122,N_19263,N_19357);
nor U20123 (N_20123,N_18234,N_19845);
nand U20124 (N_20124,N_18949,N_18188);
xnor U20125 (N_20125,N_18863,N_19952);
and U20126 (N_20126,N_17636,N_17940);
and U20127 (N_20127,N_18770,N_19083);
xor U20128 (N_20128,N_18790,N_18501);
and U20129 (N_20129,N_19266,N_19973);
nor U20130 (N_20130,N_18373,N_19746);
and U20131 (N_20131,N_19575,N_19441);
nand U20132 (N_20132,N_19708,N_19085);
or U20133 (N_20133,N_19792,N_19369);
or U20134 (N_20134,N_18285,N_18169);
or U20135 (N_20135,N_17883,N_17590);
nor U20136 (N_20136,N_19561,N_19704);
and U20137 (N_20137,N_19740,N_19492);
and U20138 (N_20138,N_18434,N_19607);
and U20139 (N_20139,N_17597,N_19130);
or U20140 (N_20140,N_19014,N_18020);
or U20141 (N_20141,N_19700,N_19484);
xnor U20142 (N_20142,N_17567,N_17749);
and U20143 (N_20143,N_19139,N_17860);
nand U20144 (N_20144,N_17942,N_19202);
and U20145 (N_20145,N_17688,N_18436);
nor U20146 (N_20146,N_17602,N_18934);
and U20147 (N_20147,N_19890,N_17806);
or U20148 (N_20148,N_18798,N_19903);
nand U20149 (N_20149,N_19099,N_19931);
or U20150 (N_20150,N_19255,N_19754);
nor U20151 (N_20151,N_19126,N_18824);
xnor U20152 (N_20152,N_18241,N_17945);
nand U20153 (N_20153,N_17665,N_18616);
nand U20154 (N_20154,N_19174,N_17580);
or U20155 (N_20155,N_19751,N_18021);
nand U20156 (N_20156,N_17820,N_17796);
or U20157 (N_20157,N_19312,N_19161);
and U20158 (N_20158,N_19853,N_18158);
and U20159 (N_20159,N_18549,N_17925);
nand U20160 (N_20160,N_17843,N_18838);
xor U20161 (N_20161,N_19285,N_19736);
or U20162 (N_20162,N_18186,N_18967);
nor U20163 (N_20163,N_19144,N_19054);
nor U20164 (N_20164,N_19098,N_19301);
nor U20165 (N_20165,N_19887,N_18993);
nand U20166 (N_20166,N_19807,N_19196);
nand U20167 (N_20167,N_19001,N_19333);
or U20168 (N_20168,N_18204,N_17589);
nor U20169 (N_20169,N_19197,N_18490);
nor U20170 (N_20170,N_19550,N_17723);
nor U20171 (N_20171,N_19388,N_18966);
or U20172 (N_20172,N_19992,N_17727);
xor U20173 (N_20173,N_19670,N_18658);
nand U20174 (N_20174,N_19612,N_17871);
or U20175 (N_20175,N_19300,N_19406);
or U20176 (N_20176,N_18767,N_19371);
or U20177 (N_20177,N_18165,N_19712);
nor U20178 (N_20178,N_18003,N_19688);
and U20179 (N_20179,N_18255,N_19215);
nor U20180 (N_20180,N_18938,N_18103);
or U20181 (N_20181,N_18073,N_18216);
nor U20182 (N_20182,N_17963,N_17610);
nor U20183 (N_20183,N_18692,N_18556);
and U20184 (N_20184,N_18019,N_19628);
nor U20185 (N_20185,N_19953,N_18356);
xor U20186 (N_20186,N_19988,N_18881);
and U20187 (N_20187,N_19008,N_19534);
nor U20188 (N_20188,N_19785,N_18269);
and U20189 (N_20189,N_19270,N_18429);
or U20190 (N_20190,N_17646,N_18207);
nor U20191 (N_20191,N_17592,N_19805);
or U20192 (N_20192,N_19722,N_19390);
and U20193 (N_20193,N_19918,N_18933);
nand U20194 (N_20194,N_17664,N_17540);
nand U20195 (N_20195,N_19037,N_19798);
nand U20196 (N_20196,N_19284,N_19456);
or U20197 (N_20197,N_18205,N_18479);
xor U20198 (N_20198,N_18590,N_19959);
or U20199 (N_20199,N_18068,N_18522);
nand U20200 (N_20200,N_18598,N_19855);
or U20201 (N_20201,N_19146,N_19298);
or U20202 (N_20202,N_18722,N_18728);
xor U20203 (N_20203,N_19836,N_19259);
nand U20204 (N_20204,N_19368,N_19104);
and U20205 (N_20205,N_17537,N_19955);
or U20206 (N_20206,N_18101,N_19960);
or U20207 (N_20207,N_17917,N_19764);
nor U20208 (N_20208,N_18145,N_18879);
nand U20209 (N_20209,N_19562,N_19823);
or U20210 (N_20210,N_17708,N_19367);
or U20211 (N_20211,N_18719,N_18920);
nor U20212 (N_20212,N_19999,N_19544);
and U20213 (N_20213,N_17888,N_17552);
and U20214 (N_20214,N_17676,N_17645);
and U20215 (N_20215,N_19508,N_18203);
or U20216 (N_20216,N_19811,N_18622);
or U20217 (N_20217,N_18820,N_17553);
and U20218 (N_20218,N_19034,N_19385);
or U20219 (N_20219,N_19088,N_17526);
xnor U20220 (N_20220,N_18502,N_18753);
or U20221 (N_20221,N_18564,N_19778);
xnor U20222 (N_20222,N_19210,N_17832);
xor U20223 (N_20223,N_19028,N_18519);
nor U20224 (N_20224,N_17993,N_18895);
or U20225 (N_20225,N_19338,N_19762);
nor U20226 (N_20226,N_18917,N_19389);
nand U20227 (N_20227,N_18815,N_19757);
nor U20228 (N_20228,N_18570,N_17818);
or U20229 (N_20229,N_18276,N_17969);
nor U20230 (N_20230,N_19061,N_18651);
nand U20231 (N_20231,N_19941,N_18701);
nand U20232 (N_20232,N_18922,N_18525);
or U20233 (N_20233,N_17899,N_19423);
nand U20234 (N_20234,N_17821,N_19684);
nor U20235 (N_20235,N_19797,N_18008);
and U20236 (N_20236,N_19543,N_17995);
nand U20237 (N_20237,N_18210,N_19308);
xor U20238 (N_20238,N_18334,N_17720);
or U20239 (N_20239,N_18856,N_19914);
nand U20240 (N_20240,N_17788,N_19068);
or U20241 (N_20241,N_17621,N_19651);
xnor U20242 (N_20242,N_19833,N_19363);
and U20243 (N_20243,N_19411,N_19726);
and U20244 (N_20244,N_19690,N_18142);
and U20245 (N_20245,N_18743,N_19501);
nand U20246 (N_20246,N_17595,N_19950);
nor U20247 (N_20247,N_18138,N_18033);
nor U20248 (N_20248,N_19701,N_19927);
and U20249 (N_20249,N_17800,N_19634);
nand U20250 (N_20250,N_19224,N_18369);
or U20251 (N_20251,N_18503,N_19148);
nor U20252 (N_20252,N_18723,N_18277);
nand U20253 (N_20253,N_17608,N_19258);
or U20254 (N_20254,N_17681,N_18673);
or U20255 (N_20255,N_17956,N_19176);
and U20256 (N_20256,N_19232,N_17524);
nor U20257 (N_20257,N_18343,N_19107);
nor U20258 (N_20258,N_18682,N_18690);
or U20259 (N_20259,N_19583,N_19460);
nor U20260 (N_20260,N_17633,N_19309);
nor U20261 (N_20261,N_17938,N_18792);
xnor U20262 (N_20262,N_17911,N_19691);
nand U20263 (N_20263,N_17866,N_19288);
xor U20264 (N_20264,N_19872,N_18977);
and U20265 (N_20265,N_19164,N_19576);
nor U20266 (N_20266,N_17859,N_18543);
nor U20267 (N_20267,N_19605,N_19303);
nand U20268 (N_20268,N_18223,N_19849);
or U20269 (N_20269,N_18776,N_19946);
nand U20270 (N_20270,N_19949,N_17954);
nand U20271 (N_20271,N_19533,N_17710);
and U20272 (N_20272,N_19814,N_17519);
or U20273 (N_20273,N_18702,N_18202);
or U20274 (N_20274,N_17725,N_18265);
or U20275 (N_20275,N_18894,N_19112);
and U20276 (N_20276,N_18497,N_18903);
nand U20277 (N_20277,N_18100,N_18166);
nor U20278 (N_20278,N_18481,N_19466);
or U20279 (N_20279,N_19647,N_17649);
nand U20280 (N_20280,N_19316,N_18833);
and U20281 (N_20281,N_19010,N_19602);
and U20282 (N_20282,N_19212,N_18378);
nor U20283 (N_20283,N_18898,N_19655);
and U20284 (N_20284,N_18161,N_19640);
xnor U20285 (N_20285,N_19517,N_18715);
nand U20286 (N_20286,N_18906,N_19816);
nor U20287 (N_20287,N_19923,N_17564);
and U20288 (N_20288,N_17760,N_18836);
or U20289 (N_20289,N_18576,N_18187);
nand U20290 (N_20290,N_19252,N_17627);
or U20291 (N_20291,N_17762,N_19100);
and U20292 (N_20292,N_19116,N_19402);
nor U20293 (N_20293,N_18678,N_18717);
nand U20294 (N_20294,N_18959,N_19409);
or U20295 (N_20295,N_17948,N_18294);
nand U20296 (N_20296,N_18244,N_17669);
and U20297 (N_20297,N_19289,N_18086);
xor U20298 (N_20298,N_18875,N_18546);
nor U20299 (N_20299,N_17643,N_18289);
nor U20300 (N_20300,N_18245,N_17699);
and U20301 (N_20301,N_18850,N_17541);
or U20302 (N_20302,N_18327,N_18756);
and U20303 (N_20303,N_19117,N_19617);
nand U20304 (N_20304,N_18148,N_19115);
xor U20305 (N_20305,N_18925,N_19079);
nor U20306 (N_20306,N_18119,N_17781);
nor U20307 (N_20307,N_18718,N_19683);
and U20308 (N_20308,N_18652,N_17895);
or U20309 (N_20309,N_17802,N_19019);
nor U20310 (N_20310,N_17848,N_18301);
nor U20311 (N_20311,N_19557,N_17828);
nor U20312 (N_20312,N_18588,N_18027);
nor U20313 (N_20313,N_19672,N_19221);
nor U20314 (N_20314,N_19172,N_18541);
and U20315 (N_20315,N_19828,N_18883);
xor U20316 (N_20316,N_18232,N_19463);
nor U20317 (N_20317,N_19377,N_18128);
xor U20318 (N_20318,N_19720,N_18286);
or U20319 (N_20319,N_19049,N_19384);
xnor U20320 (N_20320,N_17555,N_18025);
or U20321 (N_20321,N_19025,N_18706);
or U20322 (N_20322,N_17622,N_17522);
nor U20323 (N_20323,N_18929,N_17858);
or U20324 (N_20324,N_18102,N_18983);
nor U20325 (N_20325,N_19292,N_19535);
and U20326 (N_20326,N_18346,N_18319);
or U20327 (N_20327,N_18239,N_18880);
nor U20328 (N_20328,N_19554,N_18821);
or U20329 (N_20329,N_18859,N_19843);
nand U20330 (N_20330,N_18493,N_18350);
nand U20331 (N_20331,N_19447,N_19936);
nand U20332 (N_20332,N_18120,N_18830);
nand U20333 (N_20333,N_19494,N_19566);
nor U20334 (N_20334,N_19419,N_19993);
nor U20335 (N_20335,N_18799,N_17950);
and U20336 (N_20336,N_18782,N_17539);
nor U20337 (N_20337,N_17514,N_17657);
and U20338 (N_20338,N_19041,N_19227);
nand U20339 (N_20339,N_19847,N_18752);
nor U20340 (N_20340,N_19179,N_18411);
or U20341 (N_20341,N_17976,N_19458);
or U20342 (N_20342,N_19865,N_19793);
nand U20343 (N_20343,N_18619,N_17873);
nor U20344 (N_20344,N_19022,N_19069);
nand U20345 (N_20345,N_19205,N_18381);
nor U20346 (N_20346,N_19268,N_18861);
nand U20347 (N_20347,N_18288,N_18762);
nand U20348 (N_20348,N_18353,N_18458);
and U20349 (N_20349,N_19404,N_18639);
and U20350 (N_20350,N_17502,N_18078);
nor U20351 (N_20351,N_19582,N_17982);
nor U20352 (N_20352,N_17511,N_19618);
or U20353 (N_20353,N_19702,N_19842);
and U20354 (N_20354,N_17574,N_18342);
and U20355 (N_20355,N_17856,N_19649);
or U20356 (N_20356,N_19777,N_19011);
or U20357 (N_20357,N_17599,N_18733);
nor U20358 (N_20358,N_19831,N_19603);
nand U20359 (N_20359,N_19526,N_18744);
nor U20360 (N_20360,N_18046,N_18013);
nor U20361 (N_20361,N_17671,N_17570);
or U20362 (N_20362,N_18646,N_19826);
or U20363 (N_20363,N_19211,N_17913);
nand U20364 (N_20364,N_19525,N_19859);
nor U20365 (N_20365,N_18954,N_19193);
nand U20366 (N_20366,N_18539,N_17826);
or U20367 (N_20367,N_17816,N_19291);
and U20368 (N_20368,N_19318,N_18889);
and U20369 (N_20369,N_18779,N_18592);
nor U20370 (N_20370,N_19063,N_19087);
xor U20371 (N_20371,N_17978,N_18251);
nor U20372 (N_20372,N_18430,N_17810);
or U20373 (N_20373,N_19505,N_19567);
nor U20374 (N_20374,N_17683,N_19863);
nor U20375 (N_20375,N_18738,N_19326);
nor U20376 (N_20376,N_18247,N_17970);
and U20377 (N_20377,N_17901,N_18695);
or U20378 (N_20378,N_19006,N_18672);
or U20379 (N_20379,N_19124,N_18781);
nor U20380 (N_20380,N_19446,N_18228);
or U20381 (N_20381,N_19926,N_19062);
xnor U20382 (N_20382,N_18386,N_18670);
nand U20383 (N_20383,N_19137,N_19020);
or U20384 (N_20384,N_18229,N_18272);
and U20385 (N_20385,N_17967,N_19269);
and U20386 (N_20386,N_17761,N_17558);
nand U20387 (N_20387,N_19709,N_18777);
xor U20388 (N_20388,N_19874,N_17837);
nand U20389 (N_20389,N_18985,N_18797);
nand U20390 (N_20390,N_18133,N_18494);
xor U20391 (N_20391,N_19775,N_17730);
nand U20392 (N_20392,N_17663,N_18191);
nand U20393 (N_20393,N_17903,N_17690);
nand U20394 (N_20394,N_17579,N_18213);
xnor U20395 (N_20395,N_17943,N_18914);
or U20396 (N_20396,N_18813,N_19445);
nor U20397 (N_20397,N_19023,N_19685);
and U20398 (N_20398,N_18184,N_19436);
and U20399 (N_20399,N_18478,N_19784);
xor U20400 (N_20400,N_18852,N_19238);
nand U20401 (N_20401,N_18874,N_19944);
and U20402 (N_20402,N_19832,N_18642);
nor U20403 (N_20403,N_19165,N_18091);
nor U20404 (N_20404,N_18153,N_19387);
xor U20405 (N_20405,N_18629,N_18841);
and U20406 (N_20406,N_17655,N_18780);
nor U20407 (N_20407,N_17784,N_17759);
or U20408 (N_20408,N_19970,N_18558);
nand U20409 (N_20409,N_19779,N_19669);
nand U20410 (N_20410,N_18721,N_18300);
nand U20411 (N_20411,N_17752,N_17547);
and U20412 (N_20412,N_19325,N_18860);
and U20413 (N_20413,N_18468,N_19689);
and U20414 (N_20414,N_18061,N_18404);
nor U20415 (N_20415,N_17507,N_19660);
nor U20416 (N_20416,N_18846,N_19609);
or U20417 (N_20417,N_19900,N_19499);
nand U20418 (N_20418,N_18697,N_19449);
and U20419 (N_20419,N_17659,N_17915);
nor U20420 (N_20420,N_17520,N_17581);
nor U20421 (N_20421,N_17787,N_19190);
or U20422 (N_20422,N_18457,N_19313);
and U20423 (N_20423,N_18275,N_19752);
xnor U20424 (N_20424,N_17672,N_18329);
nor U20425 (N_20425,N_19795,N_17594);
nand U20426 (N_20426,N_18132,N_17732);
nor U20427 (N_20427,N_19974,N_18391);
and U20428 (N_20428,N_18891,N_19052);
nor U20429 (N_20429,N_18845,N_17576);
and U20430 (N_20430,N_18238,N_17613);
xnor U20431 (N_20431,N_18341,N_19507);
nand U20432 (N_20432,N_18840,N_18545);
xor U20433 (N_20433,N_19933,N_17606);
xnor U20434 (N_20434,N_19744,N_19675);
nor U20435 (N_20435,N_18322,N_19009);
nor U20436 (N_20436,N_17960,N_19145);
nand U20437 (N_20437,N_17550,N_19929);
or U20438 (N_20438,N_18870,N_19747);
or U20439 (N_20439,N_19482,N_19662);
or U20440 (N_20440,N_18606,N_17735);
nor U20441 (N_20441,N_17704,N_19483);
nand U20442 (N_20442,N_18750,N_18387);
and U20443 (N_20443,N_19468,N_17897);
and U20444 (N_20444,N_17734,N_18778);
nor U20445 (N_20445,N_18865,N_18605);
nand U20446 (N_20446,N_17677,N_18893);
and U20447 (N_20447,N_17624,N_18514);
or U20448 (N_20448,N_17905,N_19064);
or U20449 (N_20449,N_17501,N_19195);
or U20450 (N_20450,N_18971,N_19815);
nand U20451 (N_20451,N_17509,N_18997);
or U20452 (N_20452,N_19342,N_19750);
xnor U20453 (N_20453,N_17833,N_18992);
nand U20454 (N_20454,N_17881,N_18467);
or U20455 (N_20455,N_19496,N_19587);
nor U20456 (N_20456,N_18657,N_18460);
nor U20457 (N_20457,N_18215,N_18164);
or U20458 (N_20458,N_19599,N_17935);
nor U20459 (N_20459,N_19344,N_18012);
xor U20460 (N_20460,N_19086,N_18359);
nand U20461 (N_20461,N_18095,N_19703);
and U20462 (N_20462,N_19366,N_18045);
nand U20463 (N_20463,N_19808,N_18347);
nand U20464 (N_20464,N_18620,N_17584);
nand U20465 (N_20465,N_18612,N_17907);
nor U20466 (N_20466,N_19804,N_19254);
and U20467 (N_20467,N_18082,N_19932);
and U20468 (N_20468,N_18952,N_19964);
and U20469 (N_20469,N_19065,N_19412);
nand U20470 (N_20470,N_17630,N_19559);
nand U20471 (N_20471,N_19774,N_19626);
nand U20472 (N_20472,N_18632,N_17678);
and U20473 (N_20473,N_19790,N_17684);
nand U20474 (N_20474,N_18786,N_19614);
nand U20475 (N_20475,N_19593,N_19030);
nand U20476 (N_20476,N_19051,N_18360);
nand U20477 (N_20477,N_18871,N_17992);
or U20478 (N_20478,N_17951,N_18844);
nor U20479 (N_20479,N_19237,N_18469);
nand U20480 (N_20480,N_17941,N_19514);
or U20481 (N_20481,N_18607,N_17985);
nor U20482 (N_20482,N_18002,N_18908);
nor U20483 (N_20483,N_18167,N_18810);
nor U20484 (N_20484,N_19897,N_18355);
nor U20485 (N_20485,N_17965,N_17611);
nor U20486 (N_20486,N_19260,N_19395);
or U20487 (N_20487,N_18726,N_19231);
nand U20488 (N_20488,N_18890,N_17577);
nor U20489 (N_20489,N_18584,N_18623);
nand U20490 (N_20490,N_18071,N_19265);
nand U20491 (N_20491,N_17568,N_17598);
xor U20492 (N_20492,N_18270,N_19091);
or U20493 (N_20493,N_18633,N_19432);
nand U20494 (N_20494,N_18981,N_18455);
nand U20495 (N_20495,N_19156,N_18591);
and U20496 (N_20496,N_18047,N_19930);
nand U20497 (N_20497,N_18575,N_17685);
or U20498 (N_20498,N_17889,N_18281);
or U20499 (N_20499,N_19844,N_19142);
nor U20500 (N_20500,N_17647,N_17578);
and U20501 (N_20501,N_18878,N_17542);
and U20502 (N_20502,N_17674,N_19128);
and U20503 (N_20503,N_18687,N_18998);
xnor U20504 (N_20504,N_19686,N_18260);
nor U20505 (N_20505,N_18956,N_19994);
nand U20506 (N_20506,N_18943,N_18383);
nand U20507 (N_20507,N_19657,N_18370);
nor U20508 (N_20508,N_18405,N_18816);
and U20509 (N_20509,N_19433,N_17949);
nor U20510 (N_20510,N_19214,N_19578);
xnor U20511 (N_20511,N_19641,N_18099);
nor U20512 (N_20512,N_19129,N_18011);
or U20513 (N_20513,N_19408,N_19539);
nand U20514 (N_20514,N_19841,N_17711);
and U20515 (N_20515,N_19336,N_19677);
xor U20516 (N_20516,N_19261,N_17625);
nand U20517 (N_20517,N_19188,N_18038);
nor U20518 (N_20518,N_18385,N_19473);
nor U20519 (N_20519,N_19943,N_18683);
nor U20520 (N_20520,N_19996,N_17532);
nor U20521 (N_20521,N_17920,N_17614);
nand U20522 (N_20522,N_18667,N_17554);
nand U20523 (N_20523,N_17637,N_19209);
and U20524 (N_20524,N_17991,N_19796);
and U20525 (N_20525,N_19782,N_17615);
or U20526 (N_20526,N_18015,N_18771);
and U20527 (N_20527,N_17990,N_18572);
and U20528 (N_20528,N_19475,N_19426);
and U20529 (N_20529,N_17544,N_18433);
and U20530 (N_20530,N_18604,N_19725);
nor U20531 (N_20531,N_18747,N_19297);
xnor U20532 (N_20532,N_19302,N_19118);
and U20533 (N_20533,N_17795,N_17634);
nand U20534 (N_20534,N_19761,N_18026);
and U20535 (N_20535,N_18825,N_18094);
or U20536 (N_20536,N_17523,N_18445);
or U20537 (N_20537,N_18451,N_18923);
nor U20538 (N_20538,N_19329,N_17679);
nand U20539 (N_20539,N_19733,N_18654);
or U20540 (N_20540,N_19427,N_17994);
nand U20541 (N_20541,N_18332,N_18508);
nand U20542 (N_20542,N_18554,N_18413);
and U20543 (N_20543,N_19939,N_19668);
or U20544 (N_20544,N_18137,N_18076);
xnor U20545 (N_20545,N_18936,N_18946);
nand U20546 (N_20546,N_17571,N_18579);
and U20547 (N_20547,N_18964,N_17693);
and U20548 (N_20548,N_19935,N_18626);
or U20549 (N_20549,N_19581,N_18710);
nor U20550 (N_20550,N_18680,N_17656);
nand U20551 (N_20551,N_18443,N_19809);
or U20552 (N_20552,N_18018,N_19380);
nand U20553 (N_20553,N_19040,N_17814);
nor U20554 (N_20554,N_18307,N_18980);
nor U20555 (N_20555,N_18224,N_19274);
nand U20556 (N_20556,N_19552,N_19478);
nor U20557 (N_20557,N_19157,N_18905);
and U20558 (N_20558,N_18696,N_18190);
nand U20559 (N_20559,N_18973,N_18568);
and U20560 (N_20560,N_19359,N_19961);
nor U20561 (N_20561,N_19027,N_17904);
nor U20562 (N_20562,N_17870,N_18448);
or U20563 (N_20563,N_18037,N_18318);
and U20564 (N_20564,N_19563,N_19403);
nor U20565 (N_20565,N_18023,N_18089);
or U20566 (N_20566,N_19169,N_18380);
or U20567 (N_20567,N_18937,N_17686);
xor U20568 (N_20568,N_19495,N_17853);
or U20569 (N_20569,N_17812,N_18292);
xor U20570 (N_20570,N_17786,N_17801);
nor U20571 (N_20571,N_18339,N_17715);
or U20572 (N_20572,N_18326,N_18614);
nor U20573 (N_20573,N_18331,N_18608);
nand U20574 (N_20574,N_19892,N_18053);
and U20575 (N_20575,N_19589,N_19017);
and U20576 (N_20576,N_18513,N_19358);
and U20577 (N_20577,N_19737,N_18127);
nand U20578 (N_20578,N_19162,N_19679);
nand U20579 (N_20579,N_18283,N_18032);
nand U20580 (N_20580,N_19835,N_19742);
nor U20581 (N_20581,N_19007,N_19912);
and U20582 (N_20582,N_17747,N_19067);
and U20583 (N_20583,N_19718,N_19812);
and U20584 (N_20584,N_19472,N_17887);
and U20585 (N_20585,N_19904,N_17700);
or U20586 (N_20586,N_19882,N_18492);
nor U20587 (N_20587,N_18534,N_19180);
xor U20588 (N_20588,N_18093,N_19998);
nand U20589 (N_20589,N_18736,N_17642);
nor U20590 (N_20590,N_18066,N_18656);
or U20591 (N_20591,N_19606,N_18274);
nor U20592 (N_20592,N_18211,N_18371);
and U20593 (N_20593,N_18958,N_19317);
or U20594 (N_20594,N_19600,N_19574);
xnor U20595 (N_20595,N_17543,N_18662);
nand U20596 (N_20596,N_18328,N_18842);
nand U20597 (N_20597,N_19666,N_18237);
nand U20598 (N_20598,N_19378,N_19131);
or U20599 (N_20599,N_19518,N_19281);
and U20600 (N_20600,N_19208,N_18907);
nor U20601 (N_20601,N_18440,N_17530);
or U20602 (N_20602,N_18942,N_17631);
nor U20603 (N_20603,N_18569,N_17744);
nor U20604 (N_20604,N_19072,N_19895);
and U20605 (N_20605,N_19519,N_19370);
xnor U20606 (N_20606,N_19975,N_17640);
nor U20607 (N_20607,N_18807,N_19327);
and U20608 (N_20608,N_18765,N_19310);
nand U20609 (N_20609,N_19694,N_17799);
and U20610 (N_20610,N_18773,N_19356);
or U20611 (N_20611,N_18377,N_18996);
nand U20612 (N_20612,N_17979,N_17609);
or U20613 (N_20613,N_19095,N_18560);
or U20614 (N_20614,N_19697,N_19906);
xnor U20615 (N_20615,N_18313,N_18124);
nor U20616 (N_20616,N_19594,N_18439);
or U20617 (N_20617,N_19758,N_19611);
nor U20618 (N_20618,N_17648,N_19199);
xor U20619 (N_20619,N_18107,N_18524);
xnor U20620 (N_20620,N_18437,N_19879);
nor U20621 (N_20621,N_19159,N_18498);
or U20622 (N_20622,N_18125,N_19958);
or U20623 (N_20623,N_19510,N_19565);
and U20624 (N_20624,N_19141,N_19591);
nor U20625 (N_20625,N_18637,N_18295);
and U20626 (N_20626,N_18984,N_19362);
xor U20627 (N_20627,N_18183,N_18542);
nand U20628 (N_20628,N_17668,N_19435);
nor U20629 (N_20629,N_17721,N_18293);
nor U20630 (N_20630,N_19246,N_18685);
or U20631 (N_20631,N_18826,N_18899);
and U20632 (N_20632,N_19194,N_17884);
xor U20633 (N_20633,N_19294,N_17714);
or U20634 (N_20634,N_19123,N_17823);
nor U20635 (N_20635,N_18877,N_17852);
nand U20636 (N_20636,N_18136,N_19084);
nand U20637 (N_20637,N_19149,N_19033);
nor U20638 (N_20638,N_19692,N_18005);
nand U20639 (N_20639,N_18280,N_17536);
nor U20640 (N_20640,N_19957,N_19968);
nor U20641 (N_20641,N_19353,N_17773);
xor U20642 (N_20642,N_18601,N_19105);
nor U20643 (N_20643,N_18600,N_19983);
or U20644 (N_20644,N_18175,N_19153);
nand U20645 (N_20645,N_18796,N_17933);
or U20646 (N_20646,N_18482,N_19470);
or U20647 (N_20647,N_18394,N_18126);
and U20648 (N_20648,N_19631,N_19621);
and U20649 (N_20649,N_19322,N_18171);
or U20650 (N_20650,N_17712,N_18837);
xor U20651 (N_20651,N_18586,N_19074);
nand U20652 (N_20652,N_19060,N_18240);
nand U20653 (N_20653,N_19568,N_19056);
nand U20654 (N_20654,N_19756,N_18348);
nor U20655 (N_20655,N_17811,N_17525);
xor U20656 (N_20656,N_19538,N_18225);
or U20657 (N_20657,N_19114,N_19693);
or U20658 (N_20658,N_19106,N_19714);
nand U20659 (N_20659,N_19150,N_18994);
xnor U20660 (N_20660,N_19158,N_17822);
nand U20661 (N_20661,N_18812,N_17557);
nor U20662 (N_20662,N_19004,N_19883);
and U20663 (N_20663,N_19528,N_17964);
nand U20664 (N_20664,N_19241,N_18267);
and U20665 (N_20665,N_19880,N_18675);
or U20666 (N_20666,N_17893,N_18259);
nand U20667 (N_20667,N_19448,N_19885);
nand U20668 (N_20668,N_19908,N_18587);
xnor U20669 (N_20669,N_18931,N_19645);
nand U20670 (N_20670,N_18146,N_19763);
xnor U20671 (N_20671,N_19861,N_18686);
or U20672 (N_20672,N_19682,N_17777);
nor U20673 (N_20673,N_17538,N_17687);
xor U20674 (N_20674,N_18111,N_18466);
nand U20675 (N_20675,N_17804,N_18074);
nand U20676 (N_20676,N_19945,N_18222);
nand U20677 (N_20677,N_19223,N_18523);
nor U20678 (N_20678,N_19638,N_19553);
nor U20679 (N_20679,N_18372,N_17505);
nor U20680 (N_20680,N_19825,N_17875);
nand U20681 (N_20681,N_19375,N_18517);
or U20682 (N_20682,N_17959,N_19332);
or U20683 (N_20683,N_19515,N_19160);
and U20684 (N_20684,N_19321,N_19942);
or U20685 (N_20685,N_17751,N_18808);
xor U20686 (N_20686,N_19818,N_18150);
and U20687 (N_20687,N_18358,N_19991);
nor U20688 (N_20688,N_18791,N_19956);
nand U20689 (N_20689,N_18230,N_17876);
nand U20690 (N_20690,N_17575,N_18544);
nand U20691 (N_20691,N_17729,N_19341);
and U20692 (N_20692,N_18088,N_19819);
nor U20693 (N_20693,N_17741,N_19296);
xor U20694 (N_20694,N_18054,N_18062);
nand U20695 (N_20695,N_19891,N_18299);
nand U20696 (N_20696,N_18246,N_18582);
or U20697 (N_20697,N_18660,N_17587);
nor U20698 (N_20698,N_18611,N_19355);
and U20699 (N_20699,N_18784,N_19636);
or U20700 (N_20700,N_19545,N_17909);
or U20701 (N_20701,N_19622,N_17660);
nor U20702 (N_20702,N_19940,N_18399);
nand U20703 (N_20703,N_19857,N_18832);
and U20704 (N_20704,N_18530,N_19830);
nand U20705 (N_20705,N_18262,N_19422);
nor U20706 (N_20706,N_18252,N_17854);
nand U20707 (N_20707,N_18602,N_18991);
nor U20708 (N_20708,N_17529,N_19119);
or U20709 (N_20709,N_18450,N_18410);
nand U20710 (N_20710,N_18603,N_18700);
and U20711 (N_20711,N_19125,N_18418);
nor U20712 (N_20712,N_19462,N_19601);
and U20713 (N_20713,N_18655,N_18308);
nand U20714 (N_20714,N_18990,N_18402);
or U20715 (N_20715,N_19979,N_17930);
and U20716 (N_20716,N_19225,N_18935);
or U20717 (N_20717,N_18843,N_19262);
and U20718 (N_20718,N_17999,N_18851);
nand U20719 (N_20719,N_18868,N_18904);
nand U20720 (N_20720,N_18397,N_19894);
or U20721 (N_20721,N_19026,N_17977);
nand U20722 (N_20722,N_19871,N_19810);
or U20723 (N_20723,N_17987,N_19920);
or U20724 (N_20724,N_19787,N_19092);
nor U20725 (N_20725,N_18173,N_18220);
nor U20726 (N_20726,N_18398,N_17798);
or U20727 (N_20727,N_18438,N_19613);
xnor U20728 (N_20728,N_19485,N_19829);
nor U20729 (N_20729,N_19910,N_19497);
nand U20730 (N_20730,N_19184,N_18357);
or U20731 (N_20731,N_18367,N_18423);
nand U20732 (N_20732,N_19875,N_19015);
xnor U20733 (N_20733,N_18317,N_19415);
nor U20734 (N_20734,N_19905,N_19122);
xnor U20735 (N_20735,N_19152,N_18461);
nor U20736 (N_20736,N_17616,N_19282);
nand U20737 (N_20737,N_18583,N_18337);
nor U20738 (N_20738,N_18531,N_17706);
nand U20739 (N_20739,N_18866,N_19236);
nand U20740 (N_20740,N_18764,N_19523);
or U20741 (N_20741,N_18574,N_18345);
and U20742 (N_20742,N_19245,N_18911);
or U20743 (N_20743,N_18809,N_18298);
nor U20744 (N_20744,N_18528,N_17716);
nor U20745 (N_20745,N_17953,N_18735);
nand U20746 (N_20746,N_19760,N_17722);
nand U20747 (N_20747,N_18406,N_18648);
nand U20748 (N_20748,N_19806,N_18344);
nor U20749 (N_20749,N_18192,N_19101);
and U20750 (N_20750,N_18420,N_18296);
or U20751 (N_20751,N_19848,N_18677);
or U20752 (N_20752,N_19753,N_18691);
and U20753 (N_20753,N_18811,N_19133);
or U20754 (N_20754,N_17707,N_18176);
xor U20755 (N_20755,N_17651,N_17790);
nor U20756 (N_20756,N_19909,N_17737);
nor U20757 (N_20757,N_17698,N_17868);
and U20758 (N_20758,N_17989,N_19869);
nand U20759 (N_20759,N_19102,N_18157);
nand U20760 (N_20760,N_19759,N_18927);
xor U20761 (N_20761,N_18761,N_18080);
nand U20762 (N_20762,N_18561,N_19328);
nand U20763 (N_20763,N_17830,N_18195);
xnor U20764 (N_20764,N_18214,N_18212);
and U20765 (N_20765,N_19000,N_19524);
xnor U20766 (N_20766,N_17867,N_19339);
nor U20767 (N_20767,N_18689,N_17782);
and U20768 (N_20768,N_19656,N_19365);
or U20769 (N_20769,N_19741,N_18595);
and U20770 (N_20770,N_19453,N_19976);
nor U20771 (N_20771,N_18751,N_18669);
and U20772 (N_20772,N_18330,N_19024);
and U20773 (N_20773,N_17872,N_17556);
and U20774 (N_20774,N_19250,N_19455);
or U20775 (N_20775,N_17736,N_18151);
xnor U20776 (N_20776,N_19769,N_19440);
nor U20777 (N_20777,N_19951,N_18031);
and U20778 (N_20778,N_18665,N_18039);
nand U20779 (N_20779,N_18847,N_18714);
and U20780 (N_20780,N_17984,N_18724);
and U20781 (N_20781,N_19481,N_19513);
nand U20782 (N_20782,N_19521,N_19699);
nand U20783 (N_20783,N_17783,N_18794);
nand U20784 (N_20784,N_18823,N_17705);
nand U20785 (N_20785,N_18593,N_17745);
nand U20786 (N_20786,N_18961,N_17944);
nand U20787 (N_20787,N_18814,N_19109);
nand U20788 (N_20788,N_18291,N_19579);
or U20789 (N_20789,N_17809,N_18520);
nor U20790 (N_20790,N_19776,N_17815);
and U20791 (N_20791,N_19780,N_18708);
xor U20792 (N_20792,N_19421,N_19234);
nand U20793 (N_20793,N_18769,N_17864);
and U20794 (N_20794,N_18540,N_18709);
and U20795 (N_20795,N_19635,N_18666);
or U20796 (N_20796,N_19077,N_17918);
and U20797 (N_20797,N_18323,N_19346);
and U20798 (N_20798,N_19821,N_18030);
nand U20799 (N_20799,N_18647,N_18618);
or U20800 (N_20800,N_19541,N_18416);
nor U20801 (N_20801,N_17923,N_17695);
or U20802 (N_20802,N_19766,N_19884);
xor U20803 (N_20803,N_17740,N_19788);
and U20804 (N_20804,N_19548,N_18999);
xor U20805 (N_20805,N_18452,N_19846);
or U20806 (N_20806,N_19331,N_17764);
xor U20807 (N_20807,N_17628,N_19428);
nand U20808 (N_20808,N_18510,N_17988);
and U20809 (N_20809,N_18793,N_19629);
and U20810 (N_20810,N_19642,N_19488);
and U20811 (N_20811,N_19186,N_18926);
nor U20812 (N_20812,N_18876,N_19711);
or U20813 (N_20813,N_19443,N_17503);
nor U20814 (N_20814,N_19969,N_18599);
nor U20815 (N_20815,N_18340,N_17929);
and U20816 (N_20816,N_18048,N_19610);
or U20817 (N_20817,N_17808,N_19503);
xnor U20818 (N_20818,N_19643,N_19967);
or U20819 (N_20819,N_17910,N_18365);
nor U20820 (N_20820,N_18644,N_17673);
or U20821 (N_20821,N_17927,N_17829);
nand U20822 (N_20822,N_17504,N_19183);
nor U20823 (N_20823,N_17779,N_17572);
nand U20824 (N_20824,N_18163,N_19767);
xnor U20825 (N_20825,N_19337,N_19592);
nor U20826 (N_20826,N_18507,N_18805);
or U20827 (N_20827,N_19650,N_18887);
or U20828 (N_20828,N_18201,N_19616);
nand U20829 (N_20829,N_17924,N_18052);
nor U20830 (N_20830,N_18953,N_18635);
or U20831 (N_20831,N_19546,N_17756);
or U20832 (N_20832,N_18585,N_18768);
and U20833 (N_20833,N_17996,N_18336);
xnor U20834 (N_20834,N_18969,N_19772);
xnor U20835 (N_20835,N_17775,N_18965);
nor U20836 (N_20836,N_19121,N_17717);
or U20837 (N_20837,N_18123,N_17623);
nor U20838 (N_20838,N_17955,N_18374);
nor U20839 (N_20839,N_18141,N_18129);
and U20840 (N_20840,N_19134,N_18010);
nand U20841 (N_20841,N_18550,N_17981);
nand U20842 (N_20842,N_18789,N_19271);
nand U20843 (N_20843,N_17789,N_19839);
nand U20844 (N_20844,N_18740,N_19990);
and U20845 (N_20845,N_18311,N_19982);
nor U20846 (N_20846,N_18854,N_17545);
nand U20847 (N_20847,N_19827,N_19305);
xor U20848 (N_20848,N_18009,N_17855);
nand U20849 (N_20849,N_18446,N_18745);
nand U20850 (N_20850,N_17831,N_18004);
and U20851 (N_20851,N_18775,N_19739);
nand U20852 (N_20852,N_18982,N_18566);
or U20853 (N_20853,N_18112,N_18711);
nand U20854 (N_20854,N_19304,N_17638);
and U20855 (N_20855,N_18419,N_19916);
nor U20856 (N_20856,N_19045,N_19311);
nor U20857 (N_20857,N_17896,N_19400);
or U20858 (N_20858,N_19620,N_17739);
or U20859 (N_20859,N_17874,N_19457);
nor U20860 (N_20860,N_19248,N_19615);
nor U20861 (N_20861,N_18757,N_19659);
nor U20862 (N_20862,N_19070,N_18749);
and U20863 (N_20863,N_17757,N_19627);
or U20864 (N_20864,N_17559,N_19512);
or U20865 (N_20865,N_18649,N_18400);
nor U20866 (N_20866,N_19192,N_19630);
nand U20867 (N_20867,N_19315,N_18042);
or U20868 (N_20868,N_19293,N_19913);
nor U20869 (N_20869,N_18804,N_19824);
nor U20870 (N_20870,N_18557,N_19413);
and U20871 (N_20871,N_19220,N_17857);
and U20872 (N_20872,N_19500,N_19547);
or U20873 (N_20873,N_17850,N_19379);
nand U20874 (N_20874,N_18143,N_17733);
or U20875 (N_20875,N_17652,N_18396);
nand U20876 (N_20876,N_19097,N_19120);
and U20877 (N_20877,N_17845,N_19002);
or U20878 (N_20878,N_18320,N_18185);
and U20879 (N_20879,N_19732,N_19360);
and U20880 (N_20880,N_18518,N_19749);
nand U20881 (N_20881,N_17508,N_19822);
nor U20882 (N_20882,N_18630,N_18693);
nand U20883 (N_20883,N_19465,N_17780);
or U20884 (N_20884,N_18559,N_18422);
or U20885 (N_20885,N_17534,N_19888);
nor U20886 (N_20886,N_17635,N_19381);
and U20887 (N_20887,N_19681,N_19705);
nor U20888 (N_20888,N_17880,N_19925);
nand U20889 (N_20889,N_19476,N_19597);
or U20890 (N_20890,N_17916,N_19187);
nand U20891 (N_20891,N_17626,N_19866);
and U20892 (N_20892,N_18072,N_17619);
or U20893 (N_20893,N_18304,N_18364);
xor U20894 (N_20894,N_18168,N_18930);
or U20895 (N_20895,N_18335,N_17758);
or U20896 (N_20896,N_18117,N_17533);
or U20897 (N_20897,N_19745,N_19244);
nand U20898 (N_20898,N_19452,N_18014);
nand U20899 (N_20899,N_19901,N_18562);
xor U20900 (N_20900,N_19286,N_18064);
xnor U20901 (N_20901,N_17937,N_19786);
or U20902 (N_20902,N_18273,N_17697);
nand U20903 (N_20903,N_19917,N_19018);
xnor U20904 (N_20904,N_19673,N_17928);
and U20905 (N_20905,N_18279,N_18079);
nor U20906 (N_20906,N_18896,N_18713);
and U20907 (N_20907,N_19813,N_18354);
nand U20908 (N_20908,N_18196,N_19429);
or U20909 (N_20909,N_18149,N_18097);
xnor U20910 (N_20910,N_17565,N_17561);
and U20911 (N_20911,N_18858,N_18664);
nand U20912 (N_20912,N_17748,N_17863);
nand U20913 (N_20913,N_18509,N_18435);
nand U20914 (N_20914,N_17604,N_17639);
nor U20915 (N_20915,N_17724,N_18115);
nand U20916 (N_20916,N_18043,N_17908);
or U20917 (N_20917,N_19048,N_19418);
and U20918 (N_20918,N_18421,N_17844);
nor U20919 (N_20919,N_17794,N_18869);
xor U20920 (N_20920,N_19490,N_19439);
and U20921 (N_20921,N_18548,N_18476);
nor U20922 (N_20922,N_18065,N_18882);
or U20923 (N_20923,N_17931,N_17966);
and U20924 (N_20924,N_19016,N_17666);
nand U20925 (N_20925,N_18226,N_19734);
and U20926 (N_20926,N_19934,N_18819);
nor U20927 (N_20927,N_19042,N_18627);
or U20928 (N_20928,N_18802,N_17849);
nor U20929 (N_20929,N_18872,N_18806);
or U20930 (N_20930,N_17551,N_19256);
nand U20931 (N_20931,N_18684,N_19151);
nor U20932 (N_20932,N_17838,N_17774);
nand U20933 (N_20933,N_19075,N_19738);
nand U20934 (N_20934,N_17767,N_19111);
and U20935 (N_20935,N_17549,N_18748);
xnor U20936 (N_20936,N_18290,N_18727);
xor U20937 (N_20937,N_19348,N_19840);
nand U20938 (N_20938,N_19717,N_17886);
or U20939 (N_20939,N_18900,N_17846);
nand U20940 (N_20940,N_18431,N_18409);
nand U20941 (N_20941,N_19954,N_18154);
and U20942 (N_20942,N_19437,N_19013);
or U20943 (N_20943,N_19794,N_18092);
and U20944 (N_20944,N_18180,N_19658);
nor U20945 (N_20945,N_17569,N_19633);
and U20946 (N_20946,N_19639,N_18580);
nor U20947 (N_20947,N_18067,N_19729);
and U20948 (N_20948,N_19103,N_18484);
nor U20949 (N_20949,N_18007,N_18472);
and U20950 (N_20950,N_19715,N_19667);
nor U20951 (N_20951,N_18392,N_18379);
nand U20952 (N_20952,N_19536,N_19299);
or U20953 (N_20953,N_17766,N_19986);
xnor U20954 (N_20954,N_17851,N_18631);
nor U20955 (N_20955,N_18785,N_19877);
or U20956 (N_20956,N_19654,N_18565);
nand U20957 (N_20957,N_19728,N_19094);
or U20958 (N_20958,N_19334,N_19243);
or U20959 (N_20959,N_18485,N_19735);
nand U20960 (N_20960,N_19089,N_19323);
nand U20961 (N_20961,N_17869,N_18916);
nand U20962 (N_20962,N_19108,N_19648);
nor U20963 (N_20963,N_17696,N_19801);
and U20964 (N_20964,N_18924,N_18505);
or U20965 (N_20965,N_18261,N_17947);
nand U20966 (N_20966,N_19723,N_19350);
nand U20967 (N_20967,N_18465,N_17971);
nand U20968 (N_20968,N_17612,N_19424);
and U20969 (N_20969,N_18118,N_17825);
nor U20970 (N_20970,N_19902,N_18516);
nor U20971 (N_20971,N_19140,N_19896);
and U20972 (N_20972,N_18521,N_18640);
or U20973 (N_20973,N_18480,N_19803);
or U20974 (N_20974,N_19398,N_18734);
nor U20975 (N_20975,N_19217,N_19502);
nor U20976 (N_20976,N_17878,N_19110);
nor U20977 (N_20977,N_18674,N_18500);
xor U20978 (N_20978,N_19713,N_19218);
nor U20979 (N_20979,N_17702,N_19743);
and U20980 (N_20980,N_18567,N_17877);
or U20981 (N_20981,N_19856,N_18537);
nor U20982 (N_20982,N_17847,N_19586);
or U20983 (N_20983,N_18475,N_19417);
xor U20984 (N_20984,N_18152,N_18853);
nand U20985 (N_20985,N_19928,N_18610);
xnor U20986 (N_20986,N_19516,N_18653);
nand U20987 (N_20987,N_18104,N_19029);
nor U20988 (N_20988,N_19382,N_19911);
nand U20989 (N_20989,N_19335,N_19166);
nor U20990 (N_20990,N_18759,N_19937);
nand U20991 (N_20991,N_18932,N_17997);
nor U20992 (N_20992,N_19073,N_19755);
nand U20993 (N_20993,N_19352,N_19168);
nor U20994 (N_20994,N_19860,N_18979);
and U20995 (N_20995,N_18029,N_18306);
xor U20996 (N_20996,N_17793,N_19768);
nand U20997 (N_20997,N_17515,N_18257);
xor U20998 (N_20998,N_17862,N_17510);
xnor U20999 (N_20999,N_19608,N_18862);
nand U21000 (N_21000,N_17573,N_19653);
nor U21001 (N_21001,N_18918,N_18189);
nor U21002 (N_21002,N_19580,N_19295);
or U21003 (N_21003,N_17842,N_18527);
nor U21004 (N_21004,N_18464,N_18720);
xor U21005 (N_21005,N_19451,N_19059);
nand U21006 (N_21006,N_18083,N_17682);
xnor U21007 (N_21007,N_17641,N_19530);
or U21008 (N_21008,N_18628,N_17500);
nand U21009 (N_21009,N_18483,N_17865);
or U21010 (N_21010,N_19343,N_18231);
xor U21011 (N_21011,N_19477,N_19283);
nand U21012 (N_21012,N_17593,N_18268);
xnor U21013 (N_21013,N_19851,N_19981);
or U21014 (N_21014,N_18986,N_19444);
nand U21015 (N_21015,N_17840,N_19556);
or U21016 (N_21016,N_18233,N_17961);
and U21017 (N_21017,N_19233,N_18264);
and U21018 (N_21018,N_17506,N_18676);
and U21019 (N_21019,N_17792,N_19661);
and U21020 (N_21020,N_18886,N_18594);
nand U21021 (N_21021,N_18801,N_18892);
and U21022 (N_21022,N_18915,N_18050);
and U21023 (N_21023,N_18944,N_19878);
or U21024 (N_21024,N_17768,N_18873);
and U21025 (N_21025,N_18495,N_17770);
or U21026 (N_21026,N_19731,N_18362);
or U21027 (N_21027,N_18248,N_18609);
or U21028 (N_21028,N_18766,N_17803);
nand U21029 (N_21029,N_19493,N_19922);
or U21030 (N_21030,N_17518,N_18022);
or U21031 (N_21031,N_19509,N_18729);
nor U21032 (N_21032,N_19873,N_18156);
nand U21033 (N_21033,N_19053,N_19351);
xnor U21034 (N_21034,N_19216,N_19469);
or U21035 (N_21035,N_19249,N_19837);
nand U21036 (N_21036,N_19907,N_18170);
nand U21037 (N_21037,N_19644,N_18016);
nand U21038 (N_21038,N_17718,N_19542);
nand U21039 (N_21039,N_17817,N_19985);
or U21040 (N_21040,N_19710,N_17952);
nor U21041 (N_21041,N_17932,N_19349);
or U21042 (N_21042,N_18135,N_19280);
nor U21043 (N_21043,N_19391,N_18526);
or U21044 (N_21044,N_19963,N_17591);
and U21045 (N_21045,N_18704,N_18615);
or U21046 (N_21046,N_18415,N_18017);
and U21047 (N_21047,N_18671,N_19665);
xnor U21048 (N_21048,N_19096,N_19206);
nand U21049 (N_21049,N_19405,N_19373);
nand U21050 (N_21050,N_17776,N_19057);
and U21051 (N_21051,N_18110,N_18641);
nand U21052 (N_21052,N_18057,N_18130);
xnor U21053 (N_21053,N_17763,N_17980);
or U21054 (N_21054,N_18758,N_18663);
nand U21055 (N_21055,N_17620,N_19226);
nor U21056 (N_21056,N_19486,N_17527);
and U21057 (N_21057,N_18106,N_18928);
or U21058 (N_21058,N_19080,N_18408);
nor U21059 (N_21059,N_19687,N_19414);
nand U21060 (N_21060,N_19127,N_17968);
or U21061 (N_21061,N_18486,N_17617);
or U21062 (N_21062,N_19520,N_18139);
xnor U21063 (N_21063,N_17746,N_19005);
nor U21064 (N_21064,N_19031,N_19251);
nor U21065 (N_21065,N_18134,N_18338);
or U21066 (N_21066,N_18040,N_18070);
nand U21067 (N_21067,N_17882,N_19320);
or U21068 (N_21068,N_17946,N_18363);
nand U21069 (N_21069,N_18788,N_18442);
and U21070 (N_21070,N_19987,N_18849);
nand U21071 (N_21071,N_18382,N_18060);
nor U21072 (N_21072,N_19240,N_18243);
nand U21073 (N_21073,N_18208,N_19434);
nor U21074 (N_21074,N_17835,N_18589);
and U21075 (N_21075,N_18962,N_17548);
xnor U21076 (N_21076,N_19537,N_18972);
nor U21077 (N_21077,N_18194,N_19730);
nor U21078 (N_21078,N_19043,N_17972);
and U21079 (N_21079,N_19012,N_18515);
xnor U21080 (N_21080,N_19980,N_18453);
nor U21081 (N_21081,N_18884,N_18366);
nor U21082 (N_21082,N_19564,N_17546);
nand U21083 (N_21083,N_18160,N_19632);
or U21084 (N_21084,N_18730,N_19450);
nand U21085 (N_21085,N_19479,N_18834);
xor U21086 (N_21086,N_19802,N_18910);
nand U21087 (N_21087,N_17583,N_18707);
nand U21088 (N_21088,N_18499,N_18774);
nor U21089 (N_21089,N_17742,N_17743);
nor U21090 (N_21090,N_19671,N_17692);
nand U21091 (N_21091,N_19324,N_18159);
and U21092 (N_21092,N_18077,N_17675);
nand U21093 (N_21093,N_18681,N_18912);
and U21094 (N_21094,N_17521,N_19572);
nand U21095 (N_21095,N_18096,N_18316);
and U21096 (N_21096,N_19154,N_17517);
nand U21097 (N_21097,N_19893,N_18645);
and U21098 (N_21098,N_19817,N_18538);
xnor U21099 (N_21099,N_18578,N_19372);
and U21100 (N_21100,N_19055,N_19135);
and U21101 (N_21101,N_19467,N_19364);
or U21102 (N_21102,N_18552,N_19781);
nor U21103 (N_21103,N_19596,N_19410);
nand U21104 (N_21104,N_19306,N_18113);
nor U21105 (N_21105,N_18310,N_17797);
and U21106 (N_21106,N_18384,N_18174);
and U21107 (N_21107,N_18069,N_19898);
nor U21108 (N_21108,N_19989,N_17661);
and U21109 (N_21109,N_19652,N_18041);
and U21110 (N_21110,N_19454,N_19203);
nand U21111 (N_21111,N_18760,N_17601);
or U21112 (N_21112,N_18085,N_19374);
nor U21113 (N_21113,N_18441,N_18947);
or U21114 (N_21114,N_18555,N_18253);
or U21115 (N_21115,N_18901,N_17902);
nor U21116 (N_21116,N_19858,N_18909);
nand U21117 (N_21117,N_19867,N_18256);
and U21118 (N_21118,N_18427,N_19138);
and U21119 (N_21119,N_19504,N_17922);
xor U21120 (N_21120,N_18732,N_19230);
or U21121 (N_21121,N_18596,N_17654);
or U21122 (N_21122,N_19182,N_19407);
nor U21123 (N_21123,N_18114,N_19549);
xnor U21124 (N_21124,N_19330,N_19676);
and U21125 (N_21125,N_18772,N_19076);
nand U21126 (N_21126,N_18688,N_19948);
nand U21127 (N_21127,N_17962,N_18081);
and U21128 (N_21128,N_17975,N_18055);
nor U21129 (N_21129,N_19213,N_19972);
nor U21130 (N_21130,N_19442,N_18428);
nor U21131 (N_21131,N_19595,N_18650);
and U21132 (N_21132,N_19397,N_18414);
nor U21133 (N_21133,N_19680,N_19136);
nor U21134 (N_21134,N_19173,N_19862);
or U21135 (N_21135,N_19185,N_19347);
nand U21136 (N_21136,N_18742,N_18471);
or U21137 (N_21137,N_17771,N_17861);
nor U21138 (N_21138,N_18388,N_17680);
and U21139 (N_21139,N_19997,N_19800);
nand U21140 (N_21140,N_18122,N_18741);
and U21141 (N_21141,N_18219,N_18661);
nor U21142 (N_21142,N_19529,N_19032);
nor U21143 (N_21143,N_18098,N_17618);
nand U21144 (N_21144,N_17563,N_18563);
or U21145 (N_21145,N_18197,N_19393);
nor U21146 (N_21146,N_19276,N_18955);
nand U21147 (N_21147,N_18504,N_19978);
or U21148 (N_21148,N_18218,N_19257);
nand U21149 (N_21149,N_19637,N_17562);
or U21150 (N_21150,N_18217,N_18375);
and U21151 (N_21151,N_19047,N_19881);
and U21152 (N_21152,N_18006,N_18746);
nor U21153 (N_21153,N_18506,N_18857);
nand U21154 (N_21154,N_18333,N_19770);
nor U21155 (N_21155,N_17512,N_18456);
or U21156 (N_21156,N_18403,N_19264);
and U21157 (N_21157,N_19235,N_19678);
nand U21158 (N_21158,N_17974,N_18535);
or U21159 (N_21159,N_19287,N_19314);
nand U21160 (N_21160,N_18249,N_19279);
and U21161 (N_21161,N_17819,N_19977);
or U21162 (N_21162,N_17841,N_18487);
and U21163 (N_21163,N_17726,N_19050);
or U21164 (N_21164,N_18488,N_18968);
or U21165 (N_21165,N_18105,N_18668);
nor U21166 (N_21166,N_19275,N_18951);
or U21167 (N_21167,N_18817,N_19471);
or U21168 (N_21168,N_19082,N_18659);
and U21169 (N_21169,N_19229,N_18314);
nor U21170 (N_21170,N_18056,N_17728);
and U21171 (N_21171,N_17921,N_18059);
or U21172 (N_21172,N_18978,N_18716);
or U21173 (N_21173,N_19870,N_18424);
or U21174 (N_21174,N_19290,N_19889);
nor U21175 (N_21175,N_17891,N_19966);
nor U21176 (N_21176,N_17973,N_18829);
nand U21177 (N_21177,N_19506,N_19962);
and U21178 (N_21178,N_18144,N_19386);
or U21179 (N_21179,N_18177,N_18368);
nor U21180 (N_21180,N_19555,N_17791);
nand U21181 (N_21181,N_19915,N_19625);
nand U21182 (N_21182,N_19838,N_17900);
or U21183 (N_21183,N_17834,N_17644);
or U21184 (N_21184,N_17703,N_18084);
nor U21185 (N_21185,N_18795,N_18034);
and U21186 (N_21186,N_17912,N_17753);
nor U21187 (N_21187,N_19394,N_17629);
nand U21188 (N_21188,N_19399,N_18625);
nor U21189 (N_21189,N_18960,N_18028);
nand U21190 (N_21190,N_18948,N_18705);
or U21191 (N_21191,N_17731,N_18897);
nand U21192 (N_21192,N_17658,N_18432);
nand U21193 (N_21193,N_18818,N_18902);
and U21194 (N_21194,N_19623,N_18108);
or U21195 (N_21195,N_19773,N_19674);
or U21196 (N_21196,N_19604,N_18121);
nor U21197 (N_21197,N_17772,N_17560);
or U21198 (N_21198,N_18855,N_19253);
nand U21199 (N_21199,N_18199,N_17582);
or U21200 (N_21200,N_19498,N_19834);
nand U21201 (N_21201,N_18058,N_18024);
or U21202 (N_21202,N_19577,N_19191);
and U21203 (N_21203,N_18621,N_18221);
and U21204 (N_21204,N_19919,N_19724);
or U21205 (N_21205,N_18131,N_18597);
or U21206 (N_21206,N_18474,N_18044);
nand U21207 (N_21207,N_17824,N_19707);
nor U21208 (N_21208,N_17957,N_19361);
nor U21209 (N_21209,N_19222,N_19430);
and U21210 (N_21210,N_17926,N_19425);
nor U21211 (N_21211,N_18155,N_18303);
and U21212 (N_21212,N_19540,N_18297);
and U21213 (N_21213,N_19624,N_18737);
nand U21214 (N_21214,N_18551,N_19163);
xor U21215 (N_21215,N_18867,N_18491);
and U21216 (N_21216,N_18783,N_19461);
and U21217 (N_21217,N_18975,N_19590);
xor U21218 (N_21218,N_18417,N_18885);
nor U21219 (N_21219,N_18725,N_19921);
and U21220 (N_21220,N_19868,N_19038);
or U21221 (N_21221,N_19046,N_18395);
and U21222 (N_21222,N_18963,N_19716);
nor U21223 (N_21223,N_18449,N_17691);
nor U21224 (N_21224,N_17603,N_17585);
nand U21225 (N_21225,N_18939,N_18206);
nand U21226 (N_21226,N_19511,N_17898);
xor U21227 (N_21227,N_19664,N_17719);
nand U21228 (N_21228,N_19489,N_19239);
nand U21229 (N_21229,N_17713,N_19619);
or U21230 (N_21230,N_19886,N_19876);
nand U21231 (N_21231,N_19527,N_19924);
nand U21232 (N_21232,N_18739,N_19995);
nor U21233 (N_21233,N_18477,N_17765);
or U21234 (N_21234,N_19569,N_18250);
and U21235 (N_21235,N_18581,N_18178);
nor U21236 (N_21236,N_18638,N_18109);
nor U21237 (N_21237,N_18049,N_18988);
xor U21238 (N_21238,N_18529,N_18822);
and U21239 (N_21239,N_17653,N_18200);
nor U21240 (N_21240,N_19201,N_19899);
nand U21241 (N_21241,N_18352,N_19200);
nand U21242 (N_21242,N_19198,N_19058);
nor U21243 (N_21243,N_17785,N_17650);
and U21244 (N_21244,N_17839,N_17879);
nor U21245 (N_21245,N_18712,N_18989);
xor U21246 (N_21246,N_18162,N_18698);
and U21247 (N_21247,N_17986,N_18090);
nand U21248 (N_21248,N_19396,N_18512);
and U21249 (N_21249,N_18577,N_19247);
and U21250 (N_21250,N_19968,N_17770);
or U21251 (N_21251,N_19428,N_19556);
nand U21252 (N_21252,N_19192,N_19163);
nor U21253 (N_21253,N_18219,N_18194);
or U21254 (N_21254,N_18526,N_17633);
nand U21255 (N_21255,N_18600,N_18164);
or U21256 (N_21256,N_19632,N_18364);
or U21257 (N_21257,N_18739,N_18705);
nand U21258 (N_21258,N_19515,N_18956);
and U21259 (N_21259,N_18782,N_17947);
nor U21260 (N_21260,N_18416,N_18335);
nand U21261 (N_21261,N_18003,N_19186);
nand U21262 (N_21262,N_18455,N_18711);
nor U21263 (N_21263,N_17640,N_17899);
and U21264 (N_21264,N_19916,N_18214);
or U21265 (N_21265,N_19366,N_19027);
nand U21266 (N_21266,N_19060,N_19713);
nand U21267 (N_21267,N_19819,N_17930);
xnor U21268 (N_21268,N_18559,N_18920);
nor U21269 (N_21269,N_17945,N_18176);
or U21270 (N_21270,N_17812,N_18362);
nand U21271 (N_21271,N_19554,N_19282);
nand U21272 (N_21272,N_19389,N_18883);
nand U21273 (N_21273,N_19799,N_19271);
nand U21274 (N_21274,N_17521,N_19976);
nand U21275 (N_21275,N_19832,N_19714);
nor U21276 (N_21276,N_18279,N_19206);
xor U21277 (N_21277,N_19403,N_18772);
or U21278 (N_21278,N_18406,N_19056);
and U21279 (N_21279,N_19858,N_19580);
nor U21280 (N_21280,N_19455,N_19078);
nand U21281 (N_21281,N_19355,N_18118);
nor U21282 (N_21282,N_19460,N_19257);
and U21283 (N_21283,N_18398,N_18311);
or U21284 (N_21284,N_18816,N_17739);
or U21285 (N_21285,N_19861,N_18896);
nand U21286 (N_21286,N_19689,N_19153);
or U21287 (N_21287,N_18580,N_19144);
and U21288 (N_21288,N_17681,N_18737);
or U21289 (N_21289,N_19951,N_18536);
nor U21290 (N_21290,N_17580,N_19214);
or U21291 (N_21291,N_19402,N_17789);
xor U21292 (N_21292,N_19320,N_18456);
nand U21293 (N_21293,N_18748,N_18081);
and U21294 (N_21294,N_17941,N_18135);
nand U21295 (N_21295,N_19458,N_19539);
nor U21296 (N_21296,N_19892,N_19209);
nor U21297 (N_21297,N_18373,N_19712);
and U21298 (N_21298,N_19513,N_18480);
or U21299 (N_21299,N_17854,N_18703);
nand U21300 (N_21300,N_17572,N_18674);
nor U21301 (N_21301,N_19646,N_18677);
nand U21302 (N_21302,N_19960,N_19707);
nand U21303 (N_21303,N_18677,N_18746);
nand U21304 (N_21304,N_18480,N_18676);
or U21305 (N_21305,N_18034,N_19915);
or U21306 (N_21306,N_18810,N_19244);
or U21307 (N_21307,N_19539,N_18962);
nor U21308 (N_21308,N_18609,N_19768);
nor U21309 (N_21309,N_18719,N_18955);
and U21310 (N_21310,N_17511,N_19525);
nor U21311 (N_21311,N_17830,N_18943);
nand U21312 (N_21312,N_17625,N_18867);
or U21313 (N_21313,N_19506,N_18858);
and U21314 (N_21314,N_19821,N_19229);
nor U21315 (N_21315,N_19351,N_19038);
and U21316 (N_21316,N_17760,N_19494);
and U21317 (N_21317,N_17716,N_18874);
or U21318 (N_21318,N_18992,N_18095);
and U21319 (N_21319,N_17671,N_19694);
or U21320 (N_21320,N_19963,N_18879);
nor U21321 (N_21321,N_17513,N_19193);
and U21322 (N_21322,N_19431,N_18127);
and U21323 (N_21323,N_18143,N_18477);
and U21324 (N_21324,N_18138,N_19273);
xnor U21325 (N_21325,N_18145,N_19350);
and U21326 (N_21326,N_18186,N_17708);
nand U21327 (N_21327,N_18954,N_18709);
or U21328 (N_21328,N_19584,N_19768);
nor U21329 (N_21329,N_19619,N_18147);
nand U21330 (N_21330,N_18570,N_18646);
nor U21331 (N_21331,N_17816,N_17820);
and U21332 (N_21332,N_18540,N_17819);
or U21333 (N_21333,N_18520,N_18697);
or U21334 (N_21334,N_18627,N_18637);
nor U21335 (N_21335,N_19908,N_17779);
nand U21336 (N_21336,N_19865,N_18111);
nor U21337 (N_21337,N_17730,N_19024);
or U21338 (N_21338,N_19037,N_17806);
and U21339 (N_21339,N_18094,N_18152);
and U21340 (N_21340,N_18026,N_19524);
nor U21341 (N_21341,N_19461,N_19884);
or U21342 (N_21342,N_19948,N_19996);
nor U21343 (N_21343,N_18855,N_19898);
and U21344 (N_21344,N_17965,N_19971);
and U21345 (N_21345,N_18578,N_18576);
or U21346 (N_21346,N_18550,N_17951);
and U21347 (N_21347,N_19218,N_18837);
nand U21348 (N_21348,N_18511,N_19272);
or U21349 (N_21349,N_17635,N_17643);
xor U21350 (N_21350,N_18822,N_19454);
or U21351 (N_21351,N_19237,N_19381);
and U21352 (N_21352,N_19513,N_17830);
and U21353 (N_21353,N_19096,N_17814);
or U21354 (N_21354,N_19567,N_17763);
or U21355 (N_21355,N_18616,N_19565);
or U21356 (N_21356,N_19732,N_19663);
nor U21357 (N_21357,N_18714,N_19702);
and U21358 (N_21358,N_19457,N_18940);
nor U21359 (N_21359,N_19083,N_19348);
or U21360 (N_21360,N_18767,N_17912);
or U21361 (N_21361,N_17828,N_17552);
nand U21362 (N_21362,N_18539,N_18453);
nand U21363 (N_21363,N_17871,N_18687);
xnor U21364 (N_21364,N_19854,N_18978);
or U21365 (N_21365,N_19872,N_17602);
and U21366 (N_21366,N_19408,N_19754);
and U21367 (N_21367,N_18474,N_19942);
or U21368 (N_21368,N_18703,N_19638);
nand U21369 (N_21369,N_18726,N_18079);
and U21370 (N_21370,N_19780,N_18235);
nor U21371 (N_21371,N_18480,N_19705);
and U21372 (N_21372,N_19784,N_19834);
or U21373 (N_21373,N_19778,N_17992);
xnor U21374 (N_21374,N_19327,N_18392);
and U21375 (N_21375,N_19353,N_17705);
nor U21376 (N_21376,N_17757,N_17640);
nand U21377 (N_21377,N_17938,N_18185);
nand U21378 (N_21378,N_19349,N_18895);
nand U21379 (N_21379,N_19702,N_19645);
and U21380 (N_21380,N_19810,N_18479);
and U21381 (N_21381,N_17572,N_19606);
and U21382 (N_21382,N_18433,N_19081);
nand U21383 (N_21383,N_19719,N_18233);
xnor U21384 (N_21384,N_18246,N_17753);
nand U21385 (N_21385,N_19488,N_18303);
or U21386 (N_21386,N_18199,N_17952);
or U21387 (N_21387,N_17978,N_18165);
or U21388 (N_21388,N_19135,N_19968);
or U21389 (N_21389,N_19740,N_18049);
xnor U21390 (N_21390,N_18609,N_18113);
and U21391 (N_21391,N_19665,N_18970);
or U21392 (N_21392,N_18608,N_18233);
xor U21393 (N_21393,N_18561,N_18042);
and U21394 (N_21394,N_18140,N_17915);
nor U21395 (N_21395,N_19774,N_17822);
or U21396 (N_21396,N_19777,N_18343);
nand U21397 (N_21397,N_19961,N_19971);
and U21398 (N_21398,N_18747,N_18050);
nor U21399 (N_21399,N_18370,N_17973);
and U21400 (N_21400,N_17921,N_17756);
xor U21401 (N_21401,N_19228,N_18319);
and U21402 (N_21402,N_19898,N_18784);
or U21403 (N_21403,N_18954,N_17992);
and U21404 (N_21404,N_18826,N_19634);
nor U21405 (N_21405,N_18407,N_19845);
nand U21406 (N_21406,N_18312,N_19763);
nor U21407 (N_21407,N_17678,N_17766);
nand U21408 (N_21408,N_19418,N_18834);
and U21409 (N_21409,N_19816,N_19753);
nand U21410 (N_21410,N_18152,N_17659);
nor U21411 (N_21411,N_17972,N_17515);
and U21412 (N_21412,N_19047,N_18551);
or U21413 (N_21413,N_18786,N_18155);
nor U21414 (N_21414,N_18861,N_18422);
nand U21415 (N_21415,N_19451,N_19330);
and U21416 (N_21416,N_18002,N_19268);
or U21417 (N_21417,N_17940,N_19934);
and U21418 (N_21418,N_18893,N_18925);
and U21419 (N_21419,N_18516,N_18107);
and U21420 (N_21420,N_19044,N_18313);
or U21421 (N_21421,N_19523,N_19975);
nand U21422 (N_21422,N_18605,N_19154);
nor U21423 (N_21423,N_19420,N_18067);
nor U21424 (N_21424,N_18693,N_18258);
or U21425 (N_21425,N_19016,N_18851);
and U21426 (N_21426,N_17512,N_19407);
nand U21427 (N_21427,N_18008,N_19267);
nor U21428 (N_21428,N_18775,N_18257);
or U21429 (N_21429,N_17950,N_19810);
nand U21430 (N_21430,N_19903,N_18158);
and U21431 (N_21431,N_19659,N_18118);
nand U21432 (N_21432,N_18213,N_18993);
nor U21433 (N_21433,N_17809,N_18958);
nor U21434 (N_21434,N_19578,N_18975);
xor U21435 (N_21435,N_19171,N_18023);
and U21436 (N_21436,N_18705,N_19804);
nor U21437 (N_21437,N_19256,N_17535);
nor U21438 (N_21438,N_18857,N_19275);
nor U21439 (N_21439,N_18734,N_18869);
or U21440 (N_21440,N_18796,N_18623);
and U21441 (N_21441,N_18351,N_19941);
and U21442 (N_21442,N_17717,N_18649);
or U21443 (N_21443,N_18511,N_18977);
or U21444 (N_21444,N_18231,N_19813);
xor U21445 (N_21445,N_17572,N_17683);
and U21446 (N_21446,N_19285,N_18586);
nand U21447 (N_21447,N_18662,N_18170);
nand U21448 (N_21448,N_18187,N_19513);
nor U21449 (N_21449,N_17580,N_19914);
or U21450 (N_21450,N_18454,N_17569);
and U21451 (N_21451,N_18542,N_19966);
and U21452 (N_21452,N_17521,N_19761);
or U21453 (N_21453,N_19739,N_19832);
and U21454 (N_21454,N_19045,N_17536);
or U21455 (N_21455,N_17955,N_19354);
or U21456 (N_21456,N_18795,N_19445);
and U21457 (N_21457,N_17712,N_19277);
nor U21458 (N_21458,N_17534,N_18359);
or U21459 (N_21459,N_18407,N_18360);
or U21460 (N_21460,N_19836,N_19567);
or U21461 (N_21461,N_18408,N_19725);
xnor U21462 (N_21462,N_19061,N_19637);
nor U21463 (N_21463,N_19444,N_18909);
nor U21464 (N_21464,N_19021,N_18433);
nand U21465 (N_21465,N_17887,N_18069);
and U21466 (N_21466,N_17903,N_19074);
nand U21467 (N_21467,N_19537,N_17692);
or U21468 (N_21468,N_18662,N_19831);
or U21469 (N_21469,N_19259,N_19444);
or U21470 (N_21470,N_17659,N_17715);
nand U21471 (N_21471,N_19123,N_19423);
nand U21472 (N_21472,N_19344,N_18002);
and U21473 (N_21473,N_18196,N_17904);
or U21474 (N_21474,N_19034,N_19661);
or U21475 (N_21475,N_19641,N_17684);
nand U21476 (N_21476,N_18173,N_19748);
and U21477 (N_21477,N_19131,N_18727);
or U21478 (N_21478,N_19608,N_17784);
nand U21479 (N_21479,N_17668,N_18476);
nor U21480 (N_21480,N_18398,N_18983);
xnor U21481 (N_21481,N_19062,N_19772);
or U21482 (N_21482,N_19275,N_17927);
and U21483 (N_21483,N_18053,N_19336);
nand U21484 (N_21484,N_17700,N_19147);
or U21485 (N_21485,N_18910,N_19829);
nor U21486 (N_21486,N_19448,N_18667);
and U21487 (N_21487,N_19637,N_18404);
xnor U21488 (N_21488,N_17635,N_19776);
nor U21489 (N_21489,N_19884,N_18809);
or U21490 (N_21490,N_18027,N_19675);
nand U21491 (N_21491,N_17679,N_17800);
nor U21492 (N_21492,N_19797,N_19691);
xnor U21493 (N_21493,N_18584,N_18297);
and U21494 (N_21494,N_17894,N_18872);
and U21495 (N_21495,N_19273,N_18561);
nand U21496 (N_21496,N_19885,N_19860);
nor U21497 (N_21497,N_17677,N_18360);
nand U21498 (N_21498,N_19421,N_18537);
or U21499 (N_21499,N_18274,N_19404);
or U21500 (N_21500,N_17875,N_18458);
nor U21501 (N_21501,N_19257,N_19131);
and U21502 (N_21502,N_18573,N_18894);
nor U21503 (N_21503,N_19153,N_19408);
and U21504 (N_21504,N_19635,N_19906);
nor U21505 (N_21505,N_19506,N_19750);
nand U21506 (N_21506,N_18959,N_17946);
or U21507 (N_21507,N_18103,N_19424);
nand U21508 (N_21508,N_19545,N_18380);
or U21509 (N_21509,N_17874,N_18569);
and U21510 (N_21510,N_18428,N_18235);
nand U21511 (N_21511,N_18351,N_18355);
nor U21512 (N_21512,N_19482,N_19739);
or U21513 (N_21513,N_19944,N_18370);
nand U21514 (N_21514,N_17590,N_17868);
and U21515 (N_21515,N_17732,N_17740);
and U21516 (N_21516,N_18975,N_18754);
nor U21517 (N_21517,N_18010,N_19069);
nor U21518 (N_21518,N_19536,N_19749);
nand U21519 (N_21519,N_19328,N_18857);
or U21520 (N_21520,N_17566,N_18216);
nor U21521 (N_21521,N_18905,N_18138);
and U21522 (N_21522,N_17570,N_18192);
or U21523 (N_21523,N_19122,N_18952);
or U21524 (N_21524,N_19341,N_17540);
nand U21525 (N_21525,N_19922,N_18765);
nand U21526 (N_21526,N_19395,N_17715);
or U21527 (N_21527,N_18613,N_18530);
and U21528 (N_21528,N_19656,N_18565);
or U21529 (N_21529,N_18699,N_18753);
xor U21530 (N_21530,N_18391,N_18282);
and U21531 (N_21531,N_19018,N_19480);
or U21532 (N_21532,N_19375,N_19960);
xor U21533 (N_21533,N_17945,N_18337);
and U21534 (N_21534,N_18523,N_19236);
or U21535 (N_21535,N_19431,N_18964);
nand U21536 (N_21536,N_19004,N_18067);
and U21537 (N_21537,N_18169,N_19540);
nor U21538 (N_21538,N_19594,N_18047);
nand U21539 (N_21539,N_18890,N_19956);
or U21540 (N_21540,N_19617,N_18054);
or U21541 (N_21541,N_19075,N_19601);
nor U21542 (N_21542,N_18596,N_17923);
xor U21543 (N_21543,N_19614,N_19758);
nor U21544 (N_21544,N_17581,N_18730);
nor U21545 (N_21545,N_17817,N_18930);
xor U21546 (N_21546,N_19665,N_19672);
nor U21547 (N_21547,N_18827,N_19584);
and U21548 (N_21548,N_18521,N_18969);
nand U21549 (N_21549,N_17557,N_19874);
and U21550 (N_21550,N_18333,N_17719);
xor U21551 (N_21551,N_18626,N_17528);
or U21552 (N_21552,N_17997,N_19587);
and U21553 (N_21553,N_18639,N_19712);
or U21554 (N_21554,N_18541,N_18861);
and U21555 (N_21555,N_19622,N_19944);
nand U21556 (N_21556,N_19967,N_18765);
nand U21557 (N_21557,N_18137,N_19849);
or U21558 (N_21558,N_18980,N_17549);
nor U21559 (N_21559,N_19904,N_17843);
nor U21560 (N_21560,N_18094,N_19522);
nor U21561 (N_21561,N_18170,N_19208);
nand U21562 (N_21562,N_17853,N_19500);
nand U21563 (N_21563,N_19545,N_18500);
xnor U21564 (N_21564,N_18596,N_19567);
nand U21565 (N_21565,N_18390,N_19795);
xnor U21566 (N_21566,N_18812,N_17530);
nand U21567 (N_21567,N_19522,N_17740);
nand U21568 (N_21568,N_18925,N_18123);
nand U21569 (N_21569,N_18359,N_18064);
or U21570 (N_21570,N_19989,N_19985);
nand U21571 (N_21571,N_19971,N_17503);
and U21572 (N_21572,N_18147,N_19987);
nor U21573 (N_21573,N_18406,N_17858);
or U21574 (N_21574,N_19183,N_19606);
or U21575 (N_21575,N_18383,N_19274);
or U21576 (N_21576,N_18315,N_17974);
and U21577 (N_21577,N_19450,N_17623);
and U21578 (N_21578,N_18305,N_18667);
and U21579 (N_21579,N_17962,N_18591);
nand U21580 (N_21580,N_18442,N_18980);
and U21581 (N_21581,N_19835,N_18503);
nor U21582 (N_21582,N_18160,N_18676);
nor U21583 (N_21583,N_18701,N_19936);
nor U21584 (N_21584,N_18020,N_18555);
nand U21585 (N_21585,N_19346,N_18903);
nand U21586 (N_21586,N_19154,N_17825);
nor U21587 (N_21587,N_18280,N_18663);
and U21588 (N_21588,N_17636,N_19272);
and U21589 (N_21589,N_17573,N_18764);
nor U21590 (N_21590,N_19371,N_19512);
nor U21591 (N_21591,N_17984,N_17562);
nor U21592 (N_21592,N_18477,N_17724);
and U21593 (N_21593,N_19086,N_19490);
nand U21594 (N_21594,N_19383,N_17633);
nor U21595 (N_21595,N_18906,N_18229);
and U21596 (N_21596,N_18121,N_17740);
or U21597 (N_21597,N_19312,N_18757);
or U21598 (N_21598,N_18196,N_18954);
and U21599 (N_21599,N_17600,N_19989);
nor U21600 (N_21600,N_17974,N_18712);
nand U21601 (N_21601,N_17865,N_18607);
or U21602 (N_21602,N_19638,N_19403);
nand U21603 (N_21603,N_17723,N_19390);
and U21604 (N_21604,N_17682,N_18569);
nand U21605 (N_21605,N_19320,N_18583);
nand U21606 (N_21606,N_19943,N_19915);
nor U21607 (N_21607,N_17531,N_19502);
nand U21608 (N_21608,N_19294,N_18597);
and U21609 (N_21609,N_17885,N_18975);
nor U21610 (N_21610,N_18611,N_18711);
or U21611 (N_21611,N_19590,N_18103);
or U21612 (N_21612,N_18995,N_17557);
nand U21613 (N_21613,N_18939,N_18174);
and U21614 (N_21614,N_19624,N_19450);
xnor U21615 (N_21615,N_18544,N_19744);
and U21616 (N_21616,N_19288,N_18386);
nor U21617 (N_21617,N_18858,N_18784);
nor U21618 (N_21618,N_17758,N_18437);
and U21619 (N_21619,N_18932,N_17548);
and U21620 (N_21620,N_18144,N_17831);
and U21621 (N_21621,N_17585,N_18303);
nand U21622 (N_21622,N_19237,N_19353);
and U21623 (N_21623,N_18230,N_19664);
nand U21624 (N_21624,N_17547,N_18762);
xnor U21625 (N_21625,N_17792,N_18840);
nor U21626 (N_21626,N_19453,N_17570);
or U21627 (N_21627,N_17832,N_19093);
nand U21628 (N_21628,N_19909,N_18921);
or U21629 (N_21629,N_19056,N_18652);
nand U21630 (N_21630,N_19483,N_18442);
or U21631 (N_21631,N_19129,N_17874);
xnor U21632 (N_21632,N_18772,N_18616);
nor U21633 (N_21633,N_18760,N_18971);
xnor U21634 (N_21634,N_19435,N_17928);
nor U21635 (N_21635,N_19838,N_18630);
nor U21636 (N_21636,N_19035,N_18183);
or U21637 (N_21637,N_18290,N_18740);
nand U21638 (N_21638,N_18259,N_19826);
nor U21639 (N_21639,N_17633,N_18529);
xnor U21640 (N_21640,N_19648,N_19999);
and U21641 (N_21641,N_18507,N_18435);
and U21642 (N_21642,N_19379,N_18848);
nand U21643 (N_21643,N_18445,N_17926);
or U21644 (N_21644,N_18652,N_19295);
and U21645 (N_21645,N_17510,N_18514);
nor U21646 (N_21646,N_17514,N_17706);
nand U21647 (N_21647,N_18726,N_17948);
nor U21648 (N_21648,N_19694,N_19991);
or U21649 (N_21649,N_18900,N_18772);
nor U21650 (N_21650,N_18939,N_18132);
or U21651 (N_21651,N_18037,N_19375);
nand U21652 (N_21652,N_19480,N_18524);
and U21653 (N_21653,N_18330,N_19073);
or U21654 (N_21654,N_17811,N_18458);
or U21655 (N_21655,N_18769,N_19525);
or U21656 (N_21656,N_18378,N_19831);
or U21657 (N_21657,N_19371,N_18583);
or U21658 (N_21658,N_18528,N_19057);
or U21659 (N_21659,N_18549,N_19373);
xnor U21660 (N_21660,N_17992,N_19630);
or U21661 (N_21661,N_19920,N_19002);
and U21662 (N_21662,N_19111,N_19277);
or U21663 (N_21663,N_17837,N_18879);
xnor U21664 (N_21664,N_18057,N_17977);
or U21665 (N_21665,N_18437,N_18148);
nand U21666 (N_21666,N_19450,N_18980);
nor U21667 (N_21667,N_17613,N_18592);
nor U21668 (N_21668,N_19664,N_18700);
and U21669 (N_21669,N_17880,N_17599);
or U21670 (N_21670,N_18428,N_19405);
and U21671 (N_21671,N_19026,N_19343);
or U21672 (N_21672,N_17680,N_19509);
and U21673 (N_21673,N_19104,N_18242);
and U21674 (N_21674,N_17702,N_19583);
nand U21675 (N_21675,N_19950,N_19973);
nand U21676 (N_21676,N_19155,N_18293);
xnor U21677 (N_21677,N_18250,N_17695);
or U21678 (N_21678,N_18561,N_18914);
and U21679 (N_21679,N_17539,N_18058);
or U21680 (N_21680,N_18779,N_19349);
nor U21681 (N_21681,N_19865,N_19110);
nand U21682 (N_21682,N_18321,N_17839);
nor U21683 (N_21683,N_19431,N_19740);
or U21684 (N_21684,N_19015,N_17960);
nor U21685 (N_21685,N_17937,N_18439);
nand U21686 (N_21686,N_19925,N_19341);
nand U21687 (N_21687,N_18572,N_19411);
xnor U21688 (N_21688,N_19653,N_19988);
nor U21689 (N_21689,N_19617,N_19780);
or U21690 (N_21690,N_18716,N_17539);
nand U21691 (N_21691,N_17535,N_17699);
xnor U21692 (N_21692,N_17946,N_18572);
xnor U21693 (N_21693,N_17837,N_19962);
and U21694 (N_21694,N_19794,N_18927);
or U21695 (N_21695,N_18672,N_18198);
nand U21696 (N_21696,N_19536,N_18693);
nand U21697 (N_21697,N_17772,N_18509);
or U21698 (N_21698,N_17629,N_19565);
nand U21699 (N_21699,N_19858,N_19926);
and U21700 (N_21700,N_19687,N_19011);
or U21701 (N_21701,N_19870,N_19192);
nand U21702 (N_21702,N_18375,N_19727);
nor U21703 (N_21703,N_18995,N_18219);
nor U21704 (N_21704,N_19654,N_17651);
or U21705 (N_21705,N_18565,N_19149);
and U21706 (N_21706,N_19347,N_17711);
and U21707 (N_21707,N_18913,N_18348);
and U21708 (N_21708,N_18847,N_18870);
or U21709 (N_21709,N_17661,N_19692);
nor U21710 (N_21710,N_19127,N_19795);
nor U21711 (N_21711,N_18430,N_18867);
nand U21712 (N_21712,N_19796,N_19673);
and U21713 (N_21713,N_18108,N_17733);
and U21714 (N_21714,N_17636,N_19503);
nor U21715 (N_21715,N_17760,N_19030);
nor U21716 (N_21716,N_19644,N_19337);
nand U21717 (N_21717,N_18461,N_19611);
nor U21718 (N_21718,N_18036,N_17993);
or U21719 (N_21719,N_18424,N_18671);
nor U21720 (N_21720,N_19913,N_18661);
nand U21721 (N_21721,N_18502,N_19635);
or U21722 (N_21722,N_18637,N_19067);
and U21723 (N_21723,N_18913,N_19023);
nor U21724 (N_21724,N_19018,N_19558);
xnor U21725 (N_21725,N_17623,N_19490);
nand U21726 (N_21726,N_18970,N_18506);
nor U21727 (N_21727,N_19742,N_17530);
xnor U21728 (N_21728,N_17967,N_18705);
nor U21729 (N_21729,N_17961,N_19910);
xor U21730 (N_21730,N_18951,N_18441);
nor U21731 (N_21731,N_19528,N_17612);
xor U21732 (N_21732,N_18543,N_19300);
or U21733 (N_21733,N_17794,N_17868);
nor U21734 (N_21734,N_17734,N_17750);
xnor U21735 (N_21735,N_19778,N_17563);
or U21736 (N_21736,N_17827,N_17538);
nand U21737 (N_21737,N_17649,N_18523);
nor U21738 (N_21738,N_17744,N_19220);
nor U21739 (N_21739,N_19280,N_18668);
and U21740 (N_21740,N_19411,N_19755);
nand U21741 (N_21741,N_18700,N_19344);
or U21742 (N_21742,N_19335,N_17934);
and U21743 (N_21743,N_19880,N_18723);
xnor U21744 (N_21744,N_18853,N_17825);
nor U21745 (N_21745,N_19547,N_19994);
or U21746 (N_21746,N_19120,N_18830);
nand U21747 (N_21747,N_19128,N_18887);
and U21748 (N_21748,N_19860,N_17561);
or U21749 (N_21749,N_19836,N_18491);
nand U21750 (N_21750,N_19544,N_19313);
nand U21751 (N_21751,N_17865,N_19131);
and U21752 (N_21752,N_18299,N_17972);
xnor U21753 (N_21753,N_18350,N_18497);
xnor U21754 (N_21754,N_18820,N_18133);
and U21755 (N_21755,N_19796,N_18829);
nor U21756 (N_21756,N_17757,N_19623);
or U21757 (N_21757,N_17591,N_18867);
or U21758 (N_21758,N_18655,N_18973);
nor U21759 (N_21759,N_19689,N_19357);
or U21760 (N_21760,N_17503,N_18040);
and U21761 (N_21761,N_19899,N_18171);
xnor U21762 (N_21762,N_19806,N_18783);
nor U21763 (N_21763,N_17661,N_17964);
or U21764 (N_21764,N_17745,N_17648);
nor U21765 (N_21765,N_18554,N_18375);
and U21766 (N_21766,N_18384,N_19564);
nor U21767 (N_21767,N_17939,N_19521);
nor U21768 (N_21768,N_18837,N_18489);
nor U21769 (N_21769,N_18653,N_18949);
or U21770 (N_21770,N_17899,N_18540);
or U21771 (N_21771,N_18075,N_17994);
nor U21772 (N_21772,N_19615,N_18072);
and U21773 (N_21773,N_18809,N_18045);
and U21774 (N_21774,N_17548,N_19687);
nor U21775 (N_21775,N_19199,N_18273);
or U21776 (N_21776,N_18380,N_19326);
and U21777 (N_21777,N_18938,N_19500);
xor U21778 (N_21778,N_19927,N_19938);
or U21779 (N_21779,N_18272,N_18481);
nand U21780 (N_21780,N_17987,N_19547);
xnor U21781 (N_21781,N_19271,N_18112);
or U21782 (N_21782,N_19851,N_19517);
nand U21783 (N_21783,N_19269,N_17860);
nand U21784 (N_21784,N_18194,N_18464);
or U21785 (N_21785,N_19337,N_17944);
nor U21786 (N_21786,N_19835,N_19733);
nand U21787 (N_21787,N_18003,N_18587);
nand U21788 (N_21788,N_19815,N_18903);
and U21789 (N_21789,N_18974,N_19191);
and U21790 (N_21790,N_17866,N_19905);
and U21791 (N_21791,N_19771,N_18112);
nand U21792 (N_21792,N_19092,N_18554);
or U21793 (N_21793,N_18006,N_17642);
nand U21794 (N_21794,N_19552,N_18331);
or U21795 (N_21795,N_18476,N_19462);
nand U21796 (N_21796,N_17823,N_18669);
nor U21797 (N_21797,N_18182,N_19929);
nor U21798 (N_21798,N_17850,N_18246);
or U21799 (N_21799,N_19238,N_19517);
nor U21800 (N_21800,N_17669,N_18533);
nand U21801 (N_21801,N_19622,N_18446);
and U21802 (N_21802,N_19596,N_18979);
or U21803 (N_21803,N_19022,N_19961);
or U21804 (N_21804,N_17540,N_18420);
nor U21805 (N_21805,N_18534,N_17952);
nor U21806 (N_21806,N_18096,N_19890);
xor U21807 (N_21807,N_19881,N_19408);
or U21808 (N_21808,N_19640,N_17826);
nor U21809 (N_21809,N_19243,N_18556);
or U21810 (N_21810,N_19050,N_19189);
or U21811 (N_21811,N_17935,N_19414);
and U21812 (N_21812,N_17704,N_17909);
xnor U21813 (N_21813,N_18880,N_18806);
nor U21814 (N_21814,N_17898,N_18511);
nor U21815 (N_21815,N_17775,N_18387);
and U21816 (N_21816,N_17633,N_17773);
and U21817 (N_21817,N_18536,N_17690);
nand U21818 (N_21818,N_18203,N_18949);
nor U21819 (N_21819,N_17780,N_18205);
and U21820 (N_21820,N_17963,N_19778);
or U21821 (N_21821,N_17618,N_18705);
and U21822 (N_21822,N_19353,N_19046);
nand U21823 (N_21823,N_19653,N_19163);
xnor U21824 (N_21824,N_19985,N_19348);
nor U21825 (N_21825,N_18145,N_18634);
or U21826 (N_21826,N_18179,N_19648);
and U21827 (N_21827,N_18327,N_19195);
and U21828 (N_21828,N_17828,N_19636);
nand U21829 (N_21829,N_18403,N_17763);
and U21830 (N_21830,N_19838,N_18259);
or U21831 (N_21831,N_18014,N_19507);
or U21832 (N_21832,N_18772,N_18520);
nand U21833 (N_21833,N_19720,N_19898);
xnor U21834 (N_21834,N_18847,N_19069);
or U21835 (N_21835,N_19438,N_18486);
and U21836 (N_21836,N_18425,N_19646);
and U21837 (N_21837,N_18922,N_17910);
nor U21838 (N_21838,N_19026,N_17663);
nand U21839 (N_21839,N_18566,N_19615);
nor U21840 (N_21840,N_19757,N_19334);
nor U21841 (N_21841,N_18758,N_19213);
nand U21842 (N_21842,N_19322,N_19672);
nor U21843 (N_21843,N_18529,N_18997);
and U21844 (N_21844,N_19820,N_18041);
and U21845 (N_21845,N_19422,N_18137);
nor U21846 (N_21846,N_17928,N_19503);
and U21847 (N_21847,N_17620,N_19348);
and U21848 (N_21848,N_18607,N_18557);
and U21849 (N_21849,N_19152,N_18594);
xnor U21850 (N_21850,N_17888,N_19602);
nor U21851 (N_21851,N_19893,N_18011);
nor U21852 (N_21852,N_19145,N_18193);
nand U21853 (N_21853,N_18354,N_19369);
and U21854 (N_21854,N_17799,N_19476);
nor U21855 (N_21855,N_18079,N_18958);
or U21856 (N_21856,N_17949,N_19529);
xor U21857 (N_21857,N_17862,N_18381);
xnor U21858 (N_21858,N_19068,N_19327);
nor U21859 (N_21859,N_18788,N_19431);
or U21860 (N_21860,N_18321,N_17537);
nor U21861 (N_21861,N_19956,N_18572);
nor U21862 (N_21862,N_18369,N_17511);
nand U21863 (N_21863,N_18264,N_17913);
and U21864 (N_21864,N_19907,N_17684);
or U21865 (N_21865,N_19918,N_18281);
xor U21866 (N_21866,N_18852,N_18965);
nand U21867 (N_21867,N_18333,N_19154);
and U21868 (N_21868,N_18638,N_17824);
or U21869 (N_21869,N_17888,N_19397);
or U21870 (N_21870,N_17542,N_18399);
or U21871 (N_21871,N_18273,N_18589);
nand U21872 (N_21872,N_18517,N_17806);
nor U21873 (N_21873,N_18996,N_19524);
nor U21874 (N_21874,N_19015,N_18469);
nand U21875 (N_21875,N_18301,N_18810);
or U21876 (N_21876,N_18198,N_18538);
xor U21877 (N_21877,N_19360,N_18430);
xor U21878 (N_21878,N_19297,N_18423);
or U21879 (N_21879,N_18270,N_18090);
or U21880 (N_21880,N_18131,N_19697);
or U21881 (N_21881,N_17906,N_19900);
or U21882 (N_21882,N_17736,N_19850);
and U21883 (N_21883,N_17698,N_17765);
nor U21884 (N_21884,N_17731,N_19376);
and U21885 (N_21885,N_18950,N_18766);
or U21886 (N_21886,N_17789,N_17854);
nand U21887 (N_21887,N_18676,N_18173);
nand U21888 (N_21888,N_18196,N_18458);
and U21889 (N_21889,N_19593,N_18004);
nand U21890 (N_21890,N_18423,N_19479);
nand U21891 (N_21891,N_18287,N_19667);
or U21892 (N_21892,N_19176,N_19682);
xnor U21893 (N_21893,N_18762,N_19880);
or U21894 (N_21894,N_19136,N_18749);
nor U21895 (N_21895,N_19419,N_19007);
nand U21896 (N_21896,N_18173,N_17896);
nand U21897 (N_21897,N_19856,N_17928);
nand U21898 (N_21898,N_18565,N_17722);
or U21899 (N_21899,N_18007,N_18037);
nor U21900 (N_21900,N_17684,N_18839);
nand U21901 (N_21901,N_17917,N_19679);
nor U21902 (N_21902,N_18709,N_19254);
nand U21903 (N_21903,N_18597,N_17584);
or U21904 (N_21904,N_17706,N_19931);
or U21905 (N_21905,N_18162,N_18903);
nor U21906 (N_21906,N_19779,N_17841);
or U21907 (N_21907,N_19546,N_19438);
or U21908 (N_21908,N_18597,N_18474);
nor U21909 (N_21909,N_19113,N_19327);
nor U21910 (N_21910,N_19619,N_17759);
nor U21911 (N_21911,N_19487,N_18578);
nand U21912 (N_21912,N_18319,N_18207);
nand U21913 (N_21913,N_19366,N_17966);
and U21914 (N_21914,N_19321,N_18734);
or U21915 (N_21915,N_18396,N_18780);
xor U21916 (N_21916,N_18540,N_19119);
and U21917 (N_21917,N_19726,N_19985);
nor U21918 (N_21918,N_19845,N_19497);
nor U21919 (N_21919,N_17638,N_18053);
xnor U21920 (N_21920,N_18882,N_19132);
nor U21921 (N_21921,N_19929,N_19425);
nand U21922 (N_21922,N_19991,N_19296);
nand U21923 (N_21923,N_19651,N_19040);
xnor U21924 (N_21924,N_19794,N_18501);
nand U21925 (N_21925,N_19309,N_19946);
or U21926 (N_21926,N_19547,N_19717);
and U21927 (N_21927,N_18759,N_17776);
or U21928 (N_21928,N_18328,N_19196);
or U21929 (N_21929,N_17629,N_19842);
xnor U21930 (N_21930,N_18337,N_17694);
or U21931 (N_21931,N_19220,N_18486);
or U21932 (N_21932,N_19870,N_17928);
or U21933 (N_21933,N_19436,N_18808);
nand U21934 (N_21934,N_17571,N_19646);
or U21935 (N_21935,N_18103,N_19588);
xor U21936 (N_21936,N_19666,N_18425);
nor U21937 (N_21937,N_18415,N_19197);
and U21938 (N_21938,N_18727,N_19156);
nor U21939 (N_21939,N_17547,N_18287);
xnor U21940 (N_21940,N_18518,N_19736);
xor U21941 (N_21941,N_19287,N_18964);
nor U21942 (N_21942,N_19818,N_19341);
xor U21943 (N_21943,N_17834,N_18299);
and U21944 (N_21944,N_18472,N_18159);
nand U21945 (N_21945,N_19496,N_19641);
nor U21946 (N_21946,N_19744,N_17895);
nand U21947 (N_21947,N_17651,N_19946);
or U21948 (N_21948,N_19579,N_18756);
nor U21949 (N_21949,N_17958,N_17780);
nand U21950 (N_21950,N_19618,N_19211);
xor U21951 (N_21951,N_18213,N_19379);
nand U21952 (N_21952,N_18441,N_18086);
or U21953 (N_21953,N_19448,N_18002);
nand U21954 (N_21954,N_18666,N_17504);
and U21955 (N_21955,N_19702,N_19249);
and U21956 (N_21956,N_18996,N_19258);
nand U21957 (N_21957,N_19202,N_17674);
nor U21958 (N_21958,N_19228,N_18310);
nand U21959 (N_21959,N_19187,N_19935);
or U21960 (N_21960,N_19585,N_18983);
and U21961 (N_21961,N_18143,N_19491);
or U21962 (N_21962,N_19376,N_19102);
nand U21963 (N_21963,N_19266,N_18159);
and U21964 (N_21964,N_18712,N_18327);
or U21965 (N_21965,N_19881,N_18021);
nand U21966 (N_21966,N_18296,N_17787);
xnor U21967 (N_21967,N_18547,N_18726);
nor U21968 (N_21968,N_19171,N_17783);
nor U21969 (N_21969,N_19316,N_18837);
nand U21970 (N_21970,N_19743,N_18159);
or U21971 (N_21971,N_18752,N_18959);
nand U21972 (N_21972,N_18548,N_19167);
xor U21973 (N_21973,N_19986,N_18649);
nor U21974 (N_21974,N_19371,N_19276);
nand U21975 (N_21975,N_17947,N_19237);
nor U21976 (N_21976,N_17601,N_18191);
nand U21977 (N_21977,N_19151,N_19892);
xnor U21978 (N_21978,N_18068,N_19596);
xor U21979 (N_21979,N_19125,N_19780);
nor U21980 (N_21980,N_17841,N_19427);
and U21981 (N_21981,N_18943,N_18172);
and U21982 (N_21982,N_19267,N_18414);
nand U21983 (N_21983,N_19408,N_19826);
nand U21984 (N_21984,N_19440,N_18940);
and U21985 (N_21985,N_19788,N_18481);
xnor U21986 (N_21986,N_18926,N_17795);
and U21987 (N_21987,N_18273,N_19523);
and U21988 (N_21988,N_19580,N_19710);
nand U21989 (N_21989,N_19743,N_18523);
nand U21990 (N_21990,N_17558,N_18321);
or U21991 (N_21991,N_17850,N_19695);
nand U21992 (N_21992,N_19957,N_19103);
or U21993 (N_21993,N_18193,N_18296);
and U21994 (N_21994,N_18182,N_18664);
nand U21995 (N_21995,N_18979,N_17702);
nand U21996 (N_21996,N_18516,N_17565);
nand U21997 (N_21997,N_19773,N_18324);
or U21998 (N_21998,N_19917,N_18511);
and U21999 (N_21999,N_19883,N_19018);
nand U22000 (N_22000,N_18125,N_18419);
and U22001 (N_22001,N_17716,N_17518);
and U22002 (N_22002,N_18800,N_18055);
and U22003 (N_22003,N_19841,N_18406);
and U22004 (N_22004,N_17595,N_17764);
and U22005 (N_22005,N_19181,N_19009);
and U22006 (N_22006,N_18660,N_17507);
or U22007 (N_22007,N_19672,N_18770);
xor U22008 (N_22008,N_18709,N_17614);
xnor U22009 (N_22009,N_17951,N_19826);
or U22010 (N_22010,N_18694,N_18924);
nor U22011 (N_22011,N_18730,N_17947);
nand U22012 (N_22012,N_19405,N_19202);
and U22013 (N_22013,N_17711,N_18321);
nand U22014 (N_22014,N_17870,N_19732);
nand U22015 (N_22015,N_17941,N_18710);
or U22016 (N_22016,N_17815,N_19734);
nor U22017 (N_22017,N_19897,N_19937);
and U22018 (N_22018,N_19830,N_19433);
and U22019 (N_22019,N_19612,N_17769);
and U22020 (N_22020,N_18176,N_18936);
or U22021 (N_22021,N_19804,N_18464);
nor U22022 (N_22022,N_18862,N_17807);
nor U22023 (N_22023,N_19533,N_19347);
nor U22024 (N_22024,N_18579,N_18781);
and U22025 (N_22025,N_19076,N_18809);
or U22026 (N_22026,N_18755,N_19980);
nor U22027 (N_22027,N_19497,N_18348);
or U22028 (N_22028,N_19461,N_18355);
or U22029 (N_22029,N_19723,N_18021);
or U22030 (N_22030,N_17916,N_19682);
or U22031 (N_22031,N_18792,N_18093);
or U22032 (N_22032,N_19377,N_17665);
xnor U22033 (N_22033,N_19730,N_18919);
and U22034 (N_22034,N_19036,N_19297);
or U22035 (N_22035,N_18841,N_18555);
nor U22036 (N_22036,N_19669,N_19880);
nor U22037 (N_22037,N_18113,N_18341);
nand U22038 (N_22038,N_19357,N_19941);
or U22039 (N_22039,N_19424,N_19513);
or U22040 (N_22040,N_17742,N_19438);
nor U22041 (N_22041,N_18831,N_17805);
and U22042 (N_22042,N_19411,N_18281);
or U22043 (N_22043,N_17720,N_19183);
nor U22044 (N_22044,N_18218,N_19532);
and U22045 (N_22045,N_18726,N_19372);
or U22046 (N_22046,N_18882,N_18698);
xor U22047 (N_22047,N_19398,N_18990);
xnor U22048 (N_22048,N_18245,N_17533);
or U22049 (N_22049,N_19683,N_19325);
nor U22050 (N_22050,N_17967,N_19884);
nor U22051 (N_22051,N_17830,N_17757);
nand U22052 (N_22052,N_19032,N_18533);
and U22053 (N_22053,N_19213,N_19696);
nand U22054 (N_22054,N_18357,N_18064);
nor U22055 (N_22055,N_18619,N_17658);
nand U22056 (N_22056,N_19666,N_17931);
nor U22057 (N_22057,N_19750,N_17584);
nand U22058 (N_22058,N_19013,N_18373);
nor U22059 (N_22059,N_18229,N_18608);
xor U22060 (N_22060,N_18914,N_19600);
or U22061 (N_22061,N_17658,N_17905);
nor U22062 (N_22062,N_19000,N_19433);
or U22063 (N_22063,N_19993,N_18507);
and U22064 (N_22064,N_18541,N_18192);
or U22065 (N_22065,N_18834,N_17821);
xor U22066 (N_22066,N_18867,N_18513);
or U22067 (N_22067,N_18192,N_17705);
nand U22068 (N_22068,N_17954,N_18194);
or U22069 (N_22069,N_18566,N_18851);
nand U22070 (N_22070,N_17958,N_19200);
and U22071 (N_22071,N_18252,N_18504);
xnor U22072 (N_22072,N_19372,N_18447);
or U22073 (N_22073,N_19907,N_18844);
or U22074 (N_22074,N_19871,N_18681);
or U22075 (N_22075,N_18112,N_17884);
or U22076 (N_22076,N_19775,N_19057);
or U22077 (N_22077,N_19228,N_19961);
nand U22078 (N_22078,N_18429,N_17836);
or U22079 (N_22079,N_19199,N_19335);
nand U22080 (N_22080,N_18194,N_19797);
or U22081 (N_22081,N_17860,N_19498);
nor U22082 (N_22082,N_19177,N_19601);
and U22083 (N_22083,N_18170,N_17804);
or U22084 (N_22084,N_17596,N_18795);
nor U22085 (N_22085,N_17623,N_17877);
nor U22086 (N_22086,N_19186,N_19663);
or U22087 (N_22087,N_18267,N_17723);
and U22088 (N_22088,N_18581,N_17948);
xnor U22089 (N_22089,N_18194,N_17620);
nand U22090 (N_22090,N_17802,N_19546);
or U22091 (N_22091,N_19023,N_17717);
and U22092 (N_22092,N_19693,N_18053);
and U22093 (N_22093,N_18904,N_18300);
and U22094 (N_22094,N_18983,N_19537);
nor U22095 (N_22095,N_19037,N_19532);
and U22096 (N_22096,N_18478,N_18002);
xnor U22097 (N_22097,N_18636,N_18933);
nor U22098 (N_22098,N_19343,N_17993);
nand U22099 (N_22099,N_19858,N_18461);
nand U22100 (N_22100,N_17859,N_18896);
nand U22101 (N_22101,N_18604,N_19563);
nand U22102 (N_22102,N_18849,N_19428);
and U22103 (N_22103,N_19464,N_18788);
xnor U22104 (N_22104,N_17550,N_19414);
or U22105 (N_22105,N_17822,N_18424);
or U22106 (N_22106,N_18346,N_19917);
nand U22107 (N_22107,N_19141,N_17896);
or U22108 (N_22108,N_18502,N_18309);
or U22109 (N_22109,N_19182,N_18673);
and U22110 (N_22110,N_19563,N_18191);
nand U22111 (N_22111,N_19670,N_19159);
or U22112 (N_22112,N_19705,N_18510);
nor U22113 (N_22113,N_17527,N_19228);
nand U22114 (N_22114,N_18036,N_18838);
and U22115 (N_22115,N_18930,N_19676);
nand U22116 (N_22116,N_17866,N_18255);
nor U22117 (N_22117,N_18800,N_17633);
nand U22118 (N_22118,N_19259,N_19291);
nor U22119 (N_22119,N_18155,N_19655);
nor U22120 (N_22120,N_17870,N_18925);
nor U22121 (N_22121,N_18442,N_19240);
or U22122 (N_22122,N_18549,N_19420);
nor U22123 (N_22123,N_18335,N_18778);
nor U22124 (N_22124,N_18129,N_18632);
nor U22125 (N_22125,N_17626,N_19385);
xnor U22126 (N_22126,N_17803,N_18470);
nand U22127 (N_22127,N_17683,N_19741);
nand U22128 (N_22128,N_19397,N_18125);
nand U22129 (N_22129,N_18557,N_18911);
xor U22130 (N_22130,N_18959,N_18243);
nand U22131 (N_22131,N_19005,N_19537);
and U22132 (N_22132,N_19857,N_19415);
nor U22133 (N_22133,N_19710,N_19311);
and U22134 (N_22134,N_19234,N_17931);
and U22135 (N_22135,N_17966,N_19015);
or U22136 (N_22136,N_18875,N_18105);
nor U22137 (N_22137,N_18584,N_19990);
or U22138 (N_22138,N_19548,N_18345);
nor U22139 (N_22139,N_17540,N_19849);
and U22140 (N_22140,N_17778,N_17574);
xnor U22141 (N_22141,N_18975,N_18527);
or U22142 (N_22142,N_18029,N_17711);
nor U22143 (N_22143,N_19958,N_19868);
nor U22144 (N_22144,N_18496,N_18655);
and U22145 (N_22145,N_19935,N_17910);
nand U22146 (N_22146,N_18759,N_19094);
xor U22147 (N_22147,N_18683,N_18644);
or U22148 (N_22148,N_19202,N_19995);
or U22149 (N_22149,N_18938,N_18305);
nor U22150 (N_22150,N_19521,N_19731);
nor U22151 (N_22151,N_18176,N_18312);
nand U22152 (N_22152,N_17975,N_18654);
nand U22153 (N_22153,N_19575,N_18335);
nor U22154 (N_22154,N_18769,N_19076);
and U22155 (N_22155,N_19643,N_19978);
or U22156 (N_22156,N_18086,N_19414);
xnor U22157 (N_22157,N_18925,N_19589);
nand U22158 (N_22158,N_18016,N_19499);
nor U22159 (N_22159,N_17725,N_18108);
xor U22160 (N_22160,N_19046,N_19339);
nor U22161 (N_22161,N_17964,N_18163);
or U22162 (N_22162,N_17652,N_19926);
or U22163 (N_22163,N_19705,N_17901);
nand U22164 (N_22164,N_19446,N_17899);
or U22165 (N_22165,N_19337,N_18759);
xor U22166 (N_22166,N_18444,N_19032);
nand U22167 (N_22167,N_19415,N_19059);
and U22168 (N_22168,N_18664,N_17844);
nor U22169 (N_22169,N_18490,N_17880);
nor U22170 (N_22170,N_19504,N_18436);
nor U22171 (N_22171,N_17619,N_18661);
and U22172 (N_22172,N_17989,N_18686);
and U22173 (N_22173,N_18976,N_19011);
nor U22174 (N_22174,N_19143,N_19158);
nor U22175 (N_22175,N_19456,N_19671);
nand U22176 (N_22176,N_18702,N_17667);
nand U22177 (N_22177,N_19508,N_18370);
xnor U22178 (N_22178,N_18777,N_17529);
nor U22179 (N_22179,N_19700,N_19192);
or U22180 (N_22180,N_18105,N_19968);
or U22181 (N_22181,N_18835,N_17886);
nor U22182 (N_22182,N_18962,N_19757);
and U22183 (N_22183,N_17833,N_19325);
xor U22184 (N_22184,N_18579,N_18371);
or U22185 (N_22185,N_18670,N_19034);
nor U22186 (N_22186,N_17616,N_19284);
xor U22187 (N_22187,N_19576,N_19802);
nand U22188 (N_22188,N_18073,N_18624);
nor U22189 (N_22189,N_18457,N_18915);
or U22190 (N_22190,N_18159,N_19058);
nor U22191 (N_22191,N_18691,N_17943);
xor U22192 (N_22192,N_19239,N_18709);
xor U22193 (N_22193,N_17901,N_19439);
xnor U22194 (N_22194,N_18996,N_18244);
nor U22195 (N_22195,N_18074,N_18918);
nor U22196 (N_22196,N_19143,N_19007);
nor U22197 (N_22197,N_18539,N_19057);
and U22198 (N_22198,N_18289,N_19691);
or U22199 (N_22199,N_18031,N_18409);
and U22200 (N_22200,N_18578,N_19450);
or U22201 (N_22201,N_17902,N_19797);
and U22202 (N_22202,N_19673,N_17717);
and U22203 (N_22203,N_17939,N_18525);
and U22204 (N_22204,N_18953,N_17885);
and U22205 (N_22205,N_18235,N_17595);
nor U22206 (N_22206,N_17600,N_19481);
and U22207 (N_22207,N_18641,N_18118);
xnor U22208 (N_22208,N_17661,N_18859);
xor U22209 (N_22209,N_19003,N_19308);
nand U22210 (N_22210,N_19571,N_17845);
nor U22211 (N_22211,N_19144,N_19465);
nand U22212 (N_22212,N_18795,N_17912);
nand U22213 (N_22213,N_18236,N_19373);
and U22214 (N_22214,N_18685,N_19481);
or U22215 (N_22215,N_18583,N_19662);
xnor U22216 (N_22216,N_18445,N_18308);
nand U22217 (N_22217,N_18132,N_19549);
or U22218 (N_22218,N_18465,N_18953);
or U22219 (N_22219,N_19276,N_18220);
and U22220 (N_22220,N_17668,N_17929);
xor U22221 (N_22221,N_19725,N_17544);
nand U22222 (N_22222,N_19847,N_17765);
nand U22223 (N_22223,N_19132,N_18821);
and U22224 (N_22224,N_18756,N_19591);
and U22225 (N_22225,N_17866,N_17511);
nand U22226 (N_22226,N_19357,N_18525);
and U22227 (N_22227,N_19553,N_19330);
and U22228 (N_22228,N_19564,N_19580);
nand U22229 (N_22229,N_17552,N_17512);
xor U22230 (N_22230,N_19108,N_18110);
or U22231 (N_22231,N_18224,N_18867);
and U22232 (N_22232,N_18025,N_19267);
and U22233 (N_22233,N_18701,N_18321);
or U22234 (N_22234,N_18736,N_19121);
nor U22235 (N_22235,N_18232,N_18045);
nor U22236 (N_22236,N_17644,N_18349);
and U22237 (N_22237,N_18897,N_19392);
nor U22238 (N_22238,N_19328,N_19232);
xor U22239 (N_22239,N_17820,N_18807);
xor U22240 (N_22240,N_17517,N_18754);
xor U22241 (N_22241,N_18210,N_19718);
nor U22242 (N_22242,N_18594,N_18405);
nor U22243 (N_22243,N_19652,N_19627);
or U22244 (N_22244,N_18650,N_19578);
nand U22245 (N_22245,N_17953,N_19622);
or U22246 (N_22246,N_18759,N_17638);
nor U22247 (N_22247,N_19114,N_18494);
and U22248 (N_22248,N_18506,N_17874);
nor U22249 (N_22249,N_17697,N_18464);
and U22250 (N_22250,N_18993,N_18420);
and U22251 (N_22251,N_19349,N_19300);
xnor U22252 (N_22252,N_17611,N_18796);
nor U22253 (N_22253,N_19398,N_18537);
nor U22254 (N_22254,N_19236,N_19199);
nor U22255 (N_22255,N_18358,N_18422);
and U22256 (N_22256,N_17843,N_17994);
nand U22257 (N_22257,N_18510,N_19707);
or U22258 (N_22258,N_17928,N_19380);
xnor U22259 (N_22259,N_19018,N_18935);
nand U22260 (N_22260,N_18208,N_18158);
nor U22261 (N_22261,N_17784,N_18326);
and U22262 (N_22262,N_18750,N_18835);
nand U22263 (N_22263,N_18090,N_19776);
and U22264 (N_22264,N_18995,N_17647);
nand U22265 (N_22265,N_19396,N_19285);
nor U22266 (N_22266,N_18591,N_17744);
nor U22267 (N_22267,N_17972,N_19561);
nor U22268 (N_22268,N_19146,N_19151);
nor U22269 (N_22269,N_18943,N_19834);
nand U22270 (N_22270,N_18488,N_19454);
nand U22271 (N_22271,N_19745,N_19867);
xnor U22272 (N_22272,N_18761,N_19190);
nand U22273 (N_22273,N_19095,N_19047);
or U22274 (N_22274,N_19685,N_18688);
or U22275 (N_22275,N_19411,N_18855);
and U22276 (N_22276,N_18952,N_18391);
nor U22277 (N_22277,N_17910,N_18300);
and U22278 (N_22278,N_18308,N_19433);
xnor U22279 (N_22279,N_19281,N_19312);
xor U22280 (N_22280,N_18251,N_17698);
and U22281 (N_22281,N_19153,N_18547);
nor U22282 (N_22282,N_18476,N_19104);
nor U22283 (N_22283,N_19690,N_18510);
or U22284 (N_22284,N_18391,N_19029);
or U22285 (N_22285,N_17556,N_18173);
xnor U22286 (N_22286,N_19474,N_18686);
nor U22287 (N_22287,N_19835,N_18825);
xor U22288 (N_22288,N_18203,N_18689);
nand U22289 (N_22289,N_19040,N_18068);
or U22290 (N_22290,N_19233,N_18220);
or U22291 (N_22291,N_19787,N_18171);
xor U22292 (N_22292,N_17667,N_18734);
nand U22293 (N_22293,N_18757,N_19570);
or U22294 (N_22294,N_18803,N_17635);
nand U22295 (N_22295,N_19577,N_17665);
and U22296 (N_22296,N_19739,N_18092);
nand U22297 (N_22297,N_17553,N_17904);
nor U22298 (N_22298,N_18673,N_19123);
or U22299 (N_22299,N_18720,N_17920);
xnor U22300 (N_22300,N_19847,N_17873);
or U22301 (N_22301,N_19261,N_17951);
nand U22302 (N_22302,N_18442,N_17901);
or U22303 (N_22303,N_19328,N_18162);
or U22304 (N_22304,N_19814,N_18857);
nor U22305 (N_22305,N_18745,N_18707);
nor U22306 (N_22306,N_18488,N_19481);
and U22307 (N_22307,N_19126,N_19348);
xor U22308 (N_22308,N_19513,N_19138);
nand U22309 (N_22309,N_19250,N_17617);
or U22310 (N_22310,N_19476,N_17923);
nand U22311 (N_22311,N_19167,N_17649);
nor U22312 (N_22312,N_18237,N_18644);
and U22313 (N_22313,N_19670,N_18211);
nor U22314 (N_22314,N_19627,N_19474);
or U22315 (N_22315,N_17544,N_19584);
or U22316 (N_22316,N_17563,N_19577);
xor U22317 (N_22317,N_18949,N_18546);
and U22318 (N_22318,N_18565,N_19164);
or U22319 (N_22319,N_17933,N_19450);
nand U22320 (N_22320,N_18749,N_19839);
or U22321 (N_22321,N_18402,N_17670);
nand U22322 (N_22322,N_18967,N_17771);
or U22323 (N_22323,N_19111,N_18129);
and U22324 (N_22324,N_18189,N_19010);
or U22325 (N_22325,N_18924,N_18730);
or U22326 (N_22326,N_19684,N_19806);
nor U22327 (N_22327,N_18326,N_17927);
and U22328 (N_22328,N_17721,N_18228);
and U22329 (N_22329,N_18084,N_19506);
nand U22330 (N_22330,N_19482,N_18029);
nand U22331 (N_22331,N_18969,N_19060);
and U22332 (N_22332,N_19036,N_18971);
xnor U22333 (N_22333,N_18675,N_19109);
nand U22334 (N_22334,N_19130,N_19517);
nor U22335 (N_22335,N_19373,N_18085);
or U22336 (N_22336,N_18093,N_19802);
nand U22337 (N_22337,N_18979,N_19055);
or U22338 (N_22338,N_17983,N_19354);
nand U22339 (N_22339,N_18616,N_19068);
nor U22340 (N_22340,N_19642,N_18058);
nand U22341 (N_22341,N_18034,N_17990);
or U22342 (N_22342,N_18354,N_18237);
nor U22343 (N_22343,N_18774,N_18200);
nor U22344 (N_22344,N_18798,N_19157);
and U22345 (N_22345,N_17653,N_17905);
nand U22346 (N_22346,N_17993,N_18229);
nand U22347 (N_22347,N_19985,N_18544);
or U22348 (N_22348,N_17602,N_18953);
xnor U22349 (N_22349,N_18594,N_19690);
nor U22350 (N_22350,N_19396,N_18312);
nor U22351 (N_22351,N_17618,N_19399);
or U22352 (N_22352,N_18142,N_19891);
and U22353 (N_22353,N_18634,N_18371);
or U22354 (N_22354,N_18872,N_18460);
or U22355 (N_22355,N_18622,N_17971);
or U22356 (N_22356,N_17645,N_18526);
nor U22357 (N_22357,N_18742,N_18660);
and U22358 (N_22358,N_18885,N_19920);
nor U22359 (N_22359,N_17593,N_19875);
xor U22360 (N_22360,N_19484,N_18565);
nand U22361 (N_22361,N_19464,N_19615);
and U22362 (N_22362,N_17586,N_18560);
and U22363 (N_22363,N_18384,N_17898);
or U22364 (N_22364,N_19771,N_19931);
nand U22365 (N_22365,N_18130,N_19900);
nand U22366 (N_22366,N_18827,N_18039);
and U22367 (N_22367,N_19287,N_18443);
or U22368 (N_22368,N_19535,N_17596);
or U22369 (N_22369,N_19521,N_19225);
and U22370 (N_22370,N_18421,N_18129);
or U22371 (N_22371,N_19900,N_18426);
xor U22372 (N_22372,N_19231,N_18978);
nand U22373 (N_22373,N_19715,N_19011);
and U22374 (N_22374,N_19795,N_17888);
nor U22375 (N_22375,N_19971,N_17999);
and U22376 (N_22376,N_17979,N_19411);
and U22377 (N_22377,N_17998,N_19129);
nand U22378 (N_22378,N_18588,N_17537);
nor U22379 (N_22379,N_19389,N_18235);
xnor U22380 (N_22380,N_18526,N_17511);
nor U22381 (N_22381,N_19675,N_19595);
nor U22382 (N_22382,N_19269,N_19631);
xor U22383 (N_22383,N_18123,N_17581);
nand U22384 (N_22384,N_18633,N_18761);
nor U22385 (N_22385,N_17667,N_18811);
and U22386 (N_22386,N_18137,N_19533);
and U22387 (N_22387,N_18360,N_17899);
nor U22388 (N_22388,N_18536,N_18023);
and U22389 (N_22389,N_18870,N_17932);
or U22390 (N_22390,N_19383,N_18578);
and U22391 (N_22391,N_18961,N_19768);
nand U22392 (N_22392,N_17772,N_18409);
xor U22393 (N_22393,N_17625,N_19610);
nor U22394 (N_22394,N_19294,N_17734);
or U22395 (N_22395,N_19122,N_19089);
xnor U22396 (N_22396,N_18217,N_19975);
nor U22397 (N_22397,N_17990,N_19386);
nand U22398 (N_22398,N_19640,N_17525);
or U22399 (N_22399,N_18995,N_18826);
or U22400 (N_22400,N_18014,N_18050);
nor U22401 (N_22401,N_19315,N_18780);
and U22402 (N_22402,N_18976,N_19224);
and U22403 (N_22403,N_19774,N_18526);
and U22404 (N_22404,N_18837,N_18848);
nand U22405 (N_22405,N_18319,N_17519);
or U22406 (N_22406,N_18114,N_18597);
nor U22407 (N_22407,N_18744,N_19035);
and U22408 (N_22408,N_19305,N_19710);
nor U22409 (N_22409,N_18620,N_17588);
xnor U22410 (N_22410,N_18813,N_18149);
nand U22411 (N_22411,N_18336,N_18162);
nor U22412 (N_22412,N_19372,N_18437);
nor U22413 (N_22413,N_19089,N_18897);
and U22414 (N_22414,N_19837,N_18175);
and U22415 (N_22415,N_19364,N_18932);
nor U22416 (N_22416,N_19786,N_19075);
nand U22417 (N_22417,N_17609,N_18123);
and U22418 (N_22418,N_19372,N_18406);
or U22419 (N_22419,N_19569,N_19004);
nand U22420 (N_22420,N_17751,N_19308);
nand U22421 (N_22421,N_17992,N_19148);
and U22422 (N_22422,N_19582,N_19117);
xnor U22423 (N_22423,N_19829,N_19703);
nor U22424 (N_22424,N_19992,N_17802);
or U22425 (N_22425,N_19504,N_19689);
and U22426 (N_22426,N_17802,N_19335);
or U22427 (N_22427,N_19092,N_18272);
nor U22428 (N_22428,N_18771,N_19731);
and U22429 (N_22429,N_17585,N_19489);
nor U22430 (N_22430,N_17858,N_18513);
nor U22431 (N_22431,N_18499,N_19650);
xor U22432 (N_22432,N_18784,N_19347);
nand U22433 (N_22433,N_18961,N_19709);
and U22434 (N_22434,N_19956,N_18812);
nand U22435 (N_22435,N_19995,N_19619);
xor U22436 (N_22436,N_17868,N_18361);
nand U22437 (N_22437,N_19614,N_19710);
xor U22438 (N_22438,N_18750,N_17992);
xor U22439 (N_22439,N_18246,N_17939);
or U22440 (N_22440,N_18977,N_19989);
nand U22441 (N_22441,N_17758,N_17567);
nor U22442 (N_22442,N_18130,N_17958);
nor U22443 (N_22443,N_19469,N_17873);
xnor U22444 (N_22444,N_19508,N_18524);
nor U22445 (N_22445,N_18296,N_19307);
or U22446 (N_22446,N_17625,N_17836);
or U22447 (N_22447,N_17830,N_18983);
xor U22448 (N_22448,N_19371,N_19429);
or U22449 (N_22449,N_18060,N_18194);
and U22450 (N_22450,N_18243,N_17917);
nand U22451 (N_22451,N_19400,N_19395);
and U22452 (N_22452,N_18092,N_19057);
nor U22453 (N_22453,N_18154,N_19464);
nand U22454 (N_22454,N_19892,N_17991);
or U22455 (N_22455,N_19713,N_19513);
nor U22456 (N_22456,N_18084,N_18616);
nor U22457 (N_22457,N_18540,N_19382);
and U22458 (N_22458,N_19047,N_19634);
nor U22459 (N_22459,N_19787,N_18561);
nand U22460 (N_22460,N_17845,N_18174);
nand U22461 (N_22461,N_19287,N_19637);
nand U22462 (N_22462,N_19952,N_18591);
or U22463 (N_22463,N_19917,N_19750);
nand U22464 (N_22464,N_17662,N_19867);
nor U22465 (N_22465,N_18422,N_18134);
or U22466 (N_22466,N_19467,N_18194);
nand U22467 (N_22467,N_19798,N_19876);
nor U22468 (N_22468,N_17584,N_17842);
or U22469 (N_22469,N_19223,N_19677);
or U22470 (N_22470,N_17787,N_18012);
or U22471 (N_22471,N_19116,N_18052);
nor U22472 (N_22472,N_19318,N_18436);
nor U22473 (N_22473,N_18699,N_18450);
or U22474 (N_22474,N_19702,N_19791);
nand U22475 (N_22475,N_18772,N_17592);
and U22476 (N_22476,N_17851,N_18300);
and U22477 (N_22477,N_18872,N_17962);
and U22478 (N_22478,N_18992,N_17830);
or U22479 (N_22479,N_19762,N_18438);
nor U22480 (N_22480,N_18551,N_19467);
and U22481 (N_22481,N_19092,N_19658);
nand U22482 (N_22482,N_18621,N_17854);
xnor U22483 (N_22483,N_17664,N_19733);
or U22484 (N_22484,N_18060,N_18837);
nand U22485 (N_22485,N_19267,N_18171);
or U22486 (N_22486,N_17890,N_19873);
or U22487 (N_22487,N_19598,N_18415);
nand U22488 (N_22488,N_17642,N_18621);
or U22489 (N_22489,N_19497,N_17550);
nor U22490 (N_22490,N_19010,N_18772);
and U22491 (N_22491,N_18296,N_18759);
nor U22492 (N_22492,N_18563,N_19280);
or U22493 (N_22493,N_19518,N_17642);
nand U22494 (N_22494,N_17704,N_19541);
nor U22495 (N_22495,N_19828,N_19911);
and U22496 (N_22496,N_18111,N_18887);
or U22497 (N_22497,N_19756,N_17637);
and U22498 (N_22498,N_18692,N_18686);
or U22499 (N_22499,N_19648,N_19873);
nand U22500 (N_22500,N_21063,N_20138);
nand U22501 (N_22501,N_20332,N_20403);
nor U22502 (N_22502,N_21901,N_22383);
and U22503 (N_22503,N_20395,N_21095);
nor U22504 (N_22504,N_20312,N_22442);
nand U22505 (N_22505,N_21548,N_21455);
nand U22506 (N_22506,N_22144,N_21560);
or U22507 (N_22507,N_20667,N_20002);
xor U22508 (N_22508,N_21649,N_22438);
and U22509 (N_22509,N_21651,N_20018);
and U22510 (N_22510,N_22317,N_20897);
and U22511 (N_22511,N_20559,N_22499);
and U22512 (N_22512,N_21406,N_20172);
and U22513 (N_22513,N_20646,N_20784);
nand U22514 (N_22514,N_20987,N_21379);
nand U22515 (N_22515,N_22197,N_21249);
nand U22516 (N_22516,N_20668,N_21674);
nor U22517 (N_22517,N_20374,N_20773);
nor U22518 (N_22518,N_21224,N_21290);
nor U22519 (N_22519,N_20610,N_22439);
or U22520 (N_22520,N_20026,N_22325);
nor U22521 (N_22521,N_20641,N_20611);
nand U22522 (N_22522,N_20300,N_21106);
nand U22523 (N_22523,N_21722,N_20745);
or U22524 (N_22524,N_21158,N_21074);
nand U22525 (N_22525,N_20953,N_22463);
nand U22526 (N_22526,N_21351,N_21782);
nor U22527 (N_22527,N_21699,N_22339);
nand U22528 (N_22528,N_21326,N_21539);
and U22529 (N_22529,N_21016,N_21933);
nor U22530 (N_22530,N_21317,N_20583);
nor U22531 (N_22531,N_21680,N_21735);
nor U22532 (N_22532,N_20006,N_20426);
or U22533 (N_22533,N_21545,N_20735);
nor U22534 (N_22534,N_21473,N_20744);
or U22535 (N_22535,N_21426,N_21822);
or U22536 (N_22536,N_22187,N_22465);
and U22537 (N_22537,N_21073,N_21082);
nand U22538 (N_22538,N_22324,N_20356);
and U22539 (N_22539,N_21432,N_22119);
and U22540 (N_22540,N_21508,N_22055);
nand U22541 (N_22541,N_22244,N_22387);
nor U22542 (N_22542,N_22243,N_21839);
nand U22543 (N_22543,N_21123,N_20189);
xnor U22544 (N_22544,N_20813,N_20309);
and U22545 (N_22545,N_20231,N_20588);
nand U22546 (N_22546,N_20830,N_22192);
and U22547 (N_22547,N_21698,N_22448);
or U22548 (N_22548,N_20587,N_20455);
and U22549 (N_22549,N_21739,N_21511);
nand U22550 (N_22550,N_20104,N_21809);
and U22551 (N_22551,N_22043,N_20206);
xnor U22552 (N_22552,N_21859,N_20024);
nor U22553 (N_22553,N_20812,N_21540);
or U22554 (N_22554,N_21000,N_21020);
or U22555 (N_22555,N_21331,N_21741);
nand U22556 (N_22556,N_20107,N_22159);
and U22557 (N_22557,N_20168,N_21627);
nor U22558 (N_22558,N_21576,N_22336);
nand U22559 (N_22559,N_21770,N_21487);
or U22560 (N_22560,N_22136,N_20379);
and U22561 (N_22561,N_20774,N_20730);
or U22562 (N_22562,N_20049,N_20962);
nand U22563 (N_22563,N_20274,N_21213);
nand U22564 (N_22564,N_20153,N_21857);
nor U22565 (N_22565,N_20797,N_21076);
or U22566 (N_22566,N_21585,N_21710);
and U22567 (N_22567,N_22452,N_21816);
nor U22568 (N_22568,N_22231,N_20928);
or U22569 (N_22569,N_21319,N_20530);
and U22570 (N_22570,N_22427,N_20943);
nor U22571 (N_22571,N_22416,N_22108);
or U22572 (N_22572,N_21477,N_20905);
and U22573 (N_22573,N_21926,N_21054);
nand U22574 (N_22574,N_21115,N_21171);
or U22575 (N_22575,N_22316,N_21754);
nor U22576 (N_22576,N_21997,N_22367);
nand U22577 (N_22577,N_20260,N_21228);
or U22578 (N_22578,N_20675,N_20293);
and U22579 (N_22579,N_22314,N_21142);
and U22580 (N_22580,N_21105,N_21904);
nand U22581 (N_22581,N_21053,N_21101);
nand U22582 (N_22582,N_21475,N_22352);
or U22583 (N_22583,N_21506,N_22093);
xor U22584 (N_22584,N_21471,N_21982);
nand U22585 (N_22585,N_20386,N_22412);
nor U22586 (N_22586,N_21701,N_22114);
or U22587 (N_22587,N_21521,N_21097);
nor U22588 (N_22588,N_21441,N_20129);
nand U22589 (N_22589,N_22489,N_20458);
nand U22590 (N_22590,N_21686,N_22125);
and U22591 (N_22591,N_21638,N_22484);
or U22592 (N_22592,N_21631,N_21446);
nand U22593 (N_22593,N_20005,N_21738);
or U22594 (N_22594,N_20051,N_20490);
and U22595 (N_22595,N_20352,N_20564);
nand U22596 (N_22596,N_21443,N_21647);
nor U22597 (N_22597,N_20252,N_21505);
nand U22598 (N_22598,N_21574,N_20299);
nand U22599 (N_22599,N_21294,N_20704);
nor U22600 (N_22600,N_20957,N_20193);
and U22601 (N_22601,N_20636,N_20253);
and U22602 (N_22602,N_21100,N_20476);
nor U22603 (N_22603,N_21579,N_21837);
nand U22604 (N_22604,N_21273,N_21892);
nor U22605 (N_22605,N_21778,N_22293);
nor U22606 (N_22606,N_20048,N_21417);
nand U22607 (N_22607,N_22300,N_22110);
nand U22608 (N_22608,N_22232,N_21241);
nand U22609 (N_22609,N_20012,N_22419);
nor U22610 (N_22610,N_21793,N_21208);
nand U22611 (N_22611,N_21794,N_22353);
or U22612 (N_22612,N_20961,N_21292);
or U22613 (N_22613,N_21977,N_22332);
and U22614 (N_22614,N_20077,N_21120);
or U22615 (N_22615,N_20337,N_20910);
nand U22616 (N_22616,N_20162,N_22425);
or U22617 (N_22617,N_21530,N_20406);
and U22618 (N_22618,N_20810,N_20714);
nor U22619 (N_22619,N_21363,N_20752);
nor U22620 (N_22620,N_20427,N_22259);
xor U22621 (N_22621,N_21360,N_20165);
and U22622 (N_22622,N_22246,N_21994);
and U22623 (N_22623,N_20766,N_20198);
nor U22624 (N_22624,N_21308,N_20452);
nor U22625 (N_22625,N_21881,N_20128);
nand U22626 (N_22626,N_21431,N_20800);
nor U22627 (N_22627,N_21732,N_21595);
and U22628 (N_22628,N_22166,N_21092);
or U22629 (N_22629,N_22486,N_21819);
nand U22630 (N_22630,N_20232,N_22037);
and U22631 (N_22631,N_21993,N_21414);
and U22632 (N_22632,N_21573,N_20184);
xor U22633 (N_22633,N_21399,N_21324);
nor U22634 (N_22634,N_20785,N_22491);
or U22635 (N_22635,N_21225,N_21419);
nand U22636 (N_22636,N_20536,N_21776);
nand U22637 (N_22637,N_21134,N_21329);
nand U22638 (N_22638,N_20974,N_21338);
or U22639 (N_22639,N_21849,N_20862);
nor U22640 (N_22640,N_21872,N_22264);
nand U22641 (N_22641,N_21646,N_21423);
and U22642 (N_22642,N_21131,N_21014);
and U22643 (N_22643,N_20259,N_21744);
and U22644 (N_22644,N_20975,N_20888);
or U22645 (N_22645,N_22320,N_21960);
nand U22646 (N_22646,N_21953,N_21543);
nor U22647 (N_22647,N_20195,N_20575);
nor U22648 (N_22648,N_21855,N_21403);
and U22649 (N_22649,N_20727,N_21510);
nand U22650 (N_22650,N_20434,N_21887);
nor U22651 (N_22651,N_21174,N_22238);
or U22652 (N_22652,N_21719,N_20145);
or U22653 (N_22653,N_21407,N_22292);
nor U22654 (N_22654,N_22370,N_21950);
xor U22655 (N_22655,N_21518,N_21046);
and U22656 (N_22656,N_20676,N_22437);
and U22657 (N_22657,N_21219,N_21884);
nand U22658 (N_22658,N_21517,N_20542);
and U22659 (N_22659,N_21655,N_22441);
nor U22660 (N_22660,N_22393,N_20204);
nand U22661 (N_22661,N_21434,N_22182);
and U22662 (N_22662,N_20461,N_21494);
nand U22663 (N_22663,N_22408,N_21908);
xor U22664 (N_22664,N_20486,N_20729);
nand U22665 (N_22665,N_20709,N_20950);
nand U22666 (N_22666,N_22083,N_20485);
or U22667 (N_22667,N_21026,N_21087);
nor U22668 (N_22668,N_22157,N_21486);
nor U22669 (N_22669,N_21571,N_20852);
nor U22670 (N_22670,N_22302,N_21670);
or U22671 (N_22671,N_20375,N_22457);
or U22672 (N_22672,N_21491,N_21610);
or U22673 (N_22673,N_22013,N_20088);
and U22674 (N_22674,N_20092,N_20883);
and U22675 (N_22675,N_22386,N_22199);
xnor U22676 (N_22676,N_21285,N_20523);
nand U22677 (N_22677,N_21445,N_20424);
nand U22678 (N_22678,N_20146,N_20546);
nand U22679 (N_22679,N_20357,N_22060);
or U22680 (N_22680,N_20914,N_21094);
nand U22681 (N_22681,N_20435,N_21524);
and U22682 (N_22682,N_21564,N_20446);
or U22683 (N_22683,N_21180,N_21798);
nor U22684 (N_22684,N_22440,N_20166);
nor U22685 (N_22685,N_20877,N_22356);
and U22686 (N_22686,N_21626,N_20809);
nand U22687 (N_22687,N_21005,N_20334);
or U22688 (N_22688,N_20670,N_22451);
nand U22689 (N_22689,N_21391,N_20469);
and U22690 (N_22690,N_20865,N_21295);
nand U22691 (N_22691,N_21709,N_20097);
nand U22692 (N_22692,N_20297,N_21973);
nand U22693 (N_22693,N_21863,N_22358);
nor U22694 (N_22694,N_22492,N_21253);
or U22695 (N_22695,N_20893,N_21384);
nand U22696 (N_22696,N_21230,N_22497);
nor U22697 (N_22697,N_21789,N_21847);
xor U22698 (N_22698,N_20903,N_21048);
nand U22699 (N_22699,N_22218,N_20681);
and U22700 (N_22700,N_21736,N_21606);
nor U22701 (N_22701,N_20303,N_20913);
nor U22702 (N_22702,N_22084,N_20388);
nor U22703 (N_22703,N_20907,N_21716);
nand U22704 (N_22704,N_21482,N_21628);
xnor U22705 (N_22705,N_22445,N_20902);
xnor U22706 (N_22706,N_20859,N_20378);
and U22707 (N_22707,N_22458,N_21562);
nand U22708 (N_22708,N_22215,N_20295);
or U22709 (N_22709,N_20529,N_20258);
nand U22710 (N_22710,N_22091,N_20840);
and U22711 (N_22711,N_22444,N_20569);
nor U22712 (N_22712,N_21650,N_21943);
nand U22713 (N_22713,N_21998,N_20108);
or U22714 (N_22714,N_20955,N_21301);
nor U22715 (N_22715,N_21924,N_21935);
and U22716 (N_22716,N_21293,N_21838);
or U22717 (N_22717,N_20627,N_22298);
or U22718 (N_22718,N_20799,N_22434);
xor U22719 (N_22719,N_20023,N_21353);
nand U22720 (N_22720,N_21252,N_20584);
xnor U22721 (N_22721,N_21199,N_21428);
or U22722 (N_22722,N_21765,N_22219);
or U22723 (N_22723,N_22252,N_21611);
nand U22724 (N_22724,N_22122,N_22255);
nor U22725 (N_22725,N_21843,N_21400);
nor U22726 (N_22726,N_20074,N_20246);
nand U22727 (N_22727,N_22056,N_22113);
nand U22728 (N_22728,N_22040,N_20130);
and U22729 (N_22729,N_20043,N_20823);
and U22730 (N_22730,N_20879,N_20020);
nor U22731 (N_22731,N_20599,N_22361);
or U22732 (N_22732,N_20288,N_22277);
or U22733 (N_22733,N_20076,N_20868);
and U22734 (N_22734,N_21251,N_22263);
or U22735 (N_22735,N_22104,N_20158);
or U22736 (N_22736,N_20245,N_20377);
nor U22737 (N_22737,N_22303,N_20554);
nor U22738 (N_22738,N_20571,N_20783);
and U22739 (N_22739,N_21001,N_22435);
nand U22740 (N_22740,N_21247,N_20934);
and U22741 (N_22741,N_22357,N_20718);
xor U22742 (N_22742,N_20963,N_20919);
or U22743 (N_22743,N_20313,N_20413);
and U22744 (N_22744,N_21472,N_20632);
nand U22745 (N_22745,N_20619,N_21879);
or U22746 (N_22746,N_21883,N_21157);
nor U22747 (N_22747,N_21182,N_21612);
xor U22748 (N_22748,N_21978,N_20763);
nor U22749 (N_22749,N_21332,N_21116);
or U22750 (N_22750,N_22268,N_22049);
nand U22751 (N_22751,N_22220,N_22189);
and U22752 (N_22752,N_21086,N_22102);
and U22753 (N_22753,N_20323,N_21167);
and U22754 (N_22754,N_20574,N_21565);
nor U22755 (N_22755,N_20188,N_21282);
nor U22756 (N_22756,N_20392,N_21860);
nand U22757 (N_22757,N_20941,N_20677);
nor U22758 (N_22758,N_21190,N_20824);
or U22759 (N_22759,N_20208,N_21726);
or U22760 (N_22760,N_22158,N_21985);
and U22761 (N_22761,N_20972,N_20673);
nor U22762 (N_22762,N_20789,N_22343);
or U22763 (N_22763,N_21175,N_21844);
nand U22764 (N_22764,N_20110,N_22087);
and U22765 (N_22765,N_20983,N_22363);
and U22766 (N_22766,N_21666,N_21963);
nor U22767 (N_22767,N_20562,N_21525);
and U22768 (N_22768,N_21939,N_21825);
nor U22769 (N_22769,N_20267,N_21952);
or U22770 (N_22770,N_21260,N_20028);
and U22771 (N_22771,N_22063,N_21430);
or U22772 (N_22772,N_22295,N_21512);
nor U22773 (N_22773,N_22217,N_20596);
and U22774 (N_22774,N_20586,N_20421);
and U22775 (N_22775,N_20516,N_21873);
and U22776 (N_22776,N_20102,N_21675);
nand U22777 (N_22777,N_21900,N_21575);
and U22778 (N_22778,N_20346,N_20811);
nand U22779 (N_22779,N_21422,N_21622);
and U22780 (N_22780,N_20924,N_20327);
nor U22781 (N_22781,N_21864,N_21614);
or U22782 (N_22782,N_21316,N_20177);
nand U22783 (N_22783,N_20843,N_20234);
or U22784 (N_22784,N_21932,N_21080);
and U22785 (N_22785,N_22262,N_21918);
or U22786 (N_22786,N_20734,N_21862);
or U22787 (N_22787,N_20923,N_22174);
nor U22788 (N_22788,N_21223,N_22390);
nand U22789 (N_22789,N_20342,N_21922);
and U22790 (N_22790,N_21028,N_20547);
nor U22791 (N_22791,N_21315,N_20242);
nor U22792 (N_22792,N_22072,N_20098);
nand U22793 (N_22793,N_22432,N_21233);
or U22794 (N_22794,N_21246,N_21453);
nor U22795 (N_22795,N_20214,N_22044);
and U22796 (N_22796,N_21243,N_22279);
nor U22797 (N_22797,N_21321,N_21058);
and U22798 (N_22798,N_21708,N_20070);
nand U22799 (N_22799,N_21533,N_20462);
or U22800 (N_22800,N_22034,N_21206);
and U22801 (N_22801,N_20436,N_20060);
xor U22802 (N_22802,N_20444,N_20994);
nor U22803 (N_22803,N_21154,N_20483);
nor U22804 (N_22804,N_21222,N_21038);
or U22805 (N_22805,N_20912,N_20221);
and U22806 (N_22806,N_20200,N_20582);
or U22807 (N_22807,N_21089,N_21577);
and U22808 (N_22808,N_21648,N_22273);
or U22809 (N_22809,N_21619,N_20227);
nand U22810 (N_22810,N_21986,N_20601);
nor U22811 (N_22811,N_21385,N_21415);
or U22812 (N_22812,N_21768,N_20578);
nor U22813 (N_22813,N_22057,N_21383);
and U22814 (N_22814,N_22326,N_22203);
and U22815 (N_22815,N_20999,N_20213);
and U22816 (N_22816,N_20971,N_20143);
nor U22817 (N_22817,N_20011,N_21201);
nand U22818 (N_22818,N_21081,N_21720);
and U22819 (N_22819,N_21919,N_21570);
nand U22820 (N_22820,N_21490,N_20556);
nor U22821 (N_22821,N_21141,N_20411);
or U22822 (N_22822,N_21203,N_20853);
or U22823 (N_22823,N_20541,N_21488);
or U22824 (N_22824,N_22288,N_20515);
and U22825 (N_22825,N_21784,N_20484);
nand U22826 (N_22826,N_21734,N_20030);
nor U22827 (N_22827,N_21874,N_20122);
xnor U22828 (N_22828,N_20197,N_21909);
or U22829 (N_22829,N_22153,N_20353);
and U22830 (N_22830,N_20080,N_20420);
nand U22831 (N_22831,N_20235,N_20320);
and U22832 (N_22832,N_20764,N_22121);
nand U22833 (N_22833,N_21124,N_21609);
xor U22834 (N_22834,N_21418,N_20470);
and U22835 (N_22835,N_20144,N_21774);
nand U22836 (N_22836,N_21071,N_20938);
nand U22837 (N_22837,N_22493,N_20638);
and U22838 (N_22838,N_21663,N_21376);
and U22839 (N_22839,N_21590,N_20655);
or U22840 (N_22840,N_22428,N_20958);
nor U22841 (N_22841,N_20271,N_21745);
or U22842 (N_22842,N_20371,N_21442);
nor U22843 (N_22843,N_22294,N_21546);
nor U22844 (N_22844,N_20058,N_21897);
nor U22845 (N_22845,N_20524,N_22366);
nand U22846 (N_22846,N_21409,N_20393);
nor U22847 (N_22847,N_20114,N_21923);
nor U22848 (N_22848,N_20980,N_22495);
nand U22849 (N_22849,N_20183,N_21931);
or U22850 (N_22850,N_20263,N_20976);
and U22851 (N_22851,N_21394,N_20233);
nor U22852 (N_22852,N_22082,N_22443);
nand U22853 (N_22853,N_21639,N_21211);
nor U22854 (N_22854,N_20453,N_20906);
and U22855 (N_22855,N_20199,N_21484);
xor U22856 (N_22856,N_20939,N_20757);
xor U22857 (N_22857,N_21300,N_22021);
nand U22858 (N_22858,N_20056,N_20580);
and U22859 (N_22859,N_21155,N_20324);
nor U22860 (N_22860,N_22075,N_21370);
nand U22861 (N_22861,N_20926,N_21368);
nand U22862 (N_22862,N_20696,N_22270);
or U22863 (N_22863,N_20385,N_22095);
and U22864 (N_22864,N_21480,N_22151);
nand U22865 (N_22865,N_21150,N_21599);
nand U22866 (N_22866,N_21821,N_20568);
xor U22867 (N_22867,N_21304,N_22156);
nand U22868 (N_22868,N_22397,N_20154);
nor U22869 (N_22869,N_20157,N_21209);
nand U22870 (N_22870,N_21481,N_20133);
and U22871 (N_22871,N_21035,N_21942);
nand U22872 (N_22872,N_21656,N_21737);
or U22873 (N_22873,N_20882,N_20970);
nor U22874 (N_22874,N_22346,N_20846);
and U22875 (N_22875,N_20629,N_21747);
xnor U22876 (N_22876,N_20040,N_21358);
nand U22877 (N_22877,N_21537,N_21306);
or U22878 (N_22878,N_21258,N_21440);
or U22879 (N_22879,N_22436,N_20224);
nor U22880 (N_22880,N_22042,N_20713);
or U22881 (N_22881,N_20397,N_22329);
and U22882 (N_22882,N_21980,N_21526);
and U22883 (N_22883,N_21478,N_20391);
xnor U22884 (N_22884,N_22265,N_21207);
xor U22885 (N_22885,N_22101,N_21658);
or U22886 (N_22886,N_20415,N_21350);
or U22887 (N_22887,N_20590,N_22237);
nor U22888 (N_22888,N_21718,N_21018);
and U22889 (N_22889,N_20750,N_20967);
nand U22890 (N_22890,N_21004,N_20365);
nor U22891 (N_22891,N_21359,N_20935);
xnor U22892 (N_22892,N_20237,N_21163);
and U22893 (N_22893,N_21911,N_21806);
nor U22894 (N_22894,N_21325,N_21657);
nor U22895 (N_22895,N_20850,N_20760);
nand U22896 (N_22896,N_20492,N_20881);
and U22897 (N_22897,N_20333,N_21501);
or U22898 (N_22898,N_20722,N_21580);
and U22899 (N_22899,N_20511,N_20022);
or U22900 (N_22900,N_21547,N_20661);
nand U22901 (N_22901,N_22453,N_20819);
and U22902 (N_22902,N_22485,N_20694);
and U22903 (N_22903,N_20538,N_20027);
nor U22904 (N_22904,N_21591,N_21790);
nand U22905 (N_22905,N_21193,N_20350);
nor U22906 (N_22906,N_20464,N_20858);
nor U22907 (N_22907,N_20500,N_21204);
or U22908 (N_22908,N_20360,N_20545);
and U22909 (N_22909,N_20517,N_20239);
nor U22910 (N_22910,N_20467,N_22011);
nor U22911 (N_22911,N_22400,N_20539);
nand U22912 (N_22912,N_20936,N_20217);
nand U22913 (N_22913,N_21928,N_22322);
nand U22914 (N_22914,N_22046,N_20284);
or U22915 (N_22915,N_20281,N_22376);
nor U22916 (N_22916,N_20419,N_20405);
nand U22917 (N_22917,N_20680,N_21126);
nand U22918 (N_22918,N_20875,N_21156);
or U22919 (N_22919,N_20880,N_20282);
and U22920 (N_22920,N_21678,N_22181);
and U22921 (N_22921,N_21457,N_21069);
nand U22922 (N_22922,N_21369,N_21949);
nand U22923 (N_22923,N_20506,N_21586);
nor U22924 (N_22924,N_20015,N_20720);
and U22925 (N_22925,N_20736,N_22471);
nor U22926 (N_22926,N_21885,N_22476);
and U22927 (N_22927,N_21408,N_21108);
nand U22928 (N_22928,N_20479,N_20156);
and U22929 (N_22929,N_21688,N_21937);
and U22930 (N_22930,N_20771,N_20854);
or U22931 (N_22931,N_21373,N_21955);
nand U22932 (N_22932,N_20649,N_21815);
nor U22933 (N_22933,N_21226,N_20756);
and U22934 (N_22934,N_22379,N_20062);
or U22935 (N_22935,N_21615,N_21060);
or U22936 (N_22936,N_22462,N_22225);
and U22937 (N_22937,N_20042,N_22271);
or U22938 (N_22938,N_21268,N_20528);
or U22939 (N_22939,N_21783,N_22071);
nand U22940 (N_22940,N_20423,N_22172);
nor U22941 (N_22941,N_22132,N_22036);
or U22942 (N_22942,N_21915,N_20451);
or U22943 (N_22943,N_20192,N_20218);
or U22944 (N_22944,N_20016,N_21188);
nand U22945 (N_22945,N_20788,N_21214);
or U22946 (N_22946,N_20430,N_21516);
and U22947 (N_22947,N_21588,N_21396);
nand U22948 (N_22948,N_20466,N_20998);
nand U22949 (N_22949,N_21832,N_22178);
nor U22950 (N_22950,N_22103,N_20244);
nor U22951 (N_22951,N_20780,N_20181);
or U22952 (N_22952,N_22191,N_20116);
nand U22953 (N_22953,N_21200,N_21968);
nor U22954 (N_22954,N_21728,N_22107);
nor U22955 (N_22955,N_21138,N_20032);
nand U22956 (N_22956,N_21807,N_20276);
nand U22957 (N_22957,N_22456,N_20220);
and U22958 (N_22958,N_20152,N_20508);
nand U22959 (N_22959,N_21189,N_21702);
and U22960 (N_22960,N_22168,N_21668);
and U22961 (N_22961,N_20621,N_22235);
or U22962 (N_22962,N_20674,N_20422);
xor U22963 (N_22963,N_22001,N_20702);
xor U22964 (N_22964,N_21593,N_22171);
or U22965 (N_22965,N_20947,N_20577);
nand U22966 (N_22966,N_21769,N_21118);
nor U22967 (N_22967,N_20510,N_21725);
nand U22968 (N_22968,N_20965,N_21781);
xor U22969 (N_22969,N_22318,N_22004);
nor U22970 (N_22970,N_20289,N_21773);
or U22971 (N_22971,N_22184,N_21168);
and U22972 (N_22972,N_22133,N_20398);
nor U22973 (N_22973,N_21818,N_22487);
and U22974 (N_22974,N_21551,N_20141);
xor U22975 (N_22975,N_21137,N_21920);
or U22976 (N_22976,N_22175,N_22478);
nand U22977 (N_22977,N_21042,N_22069);
and U22978 (N_22978,N_21870,N_20657);
nor U22979 (N_22979,N_20683,N_20951);
nand U22980 (N_22980,N_20782,N_20169);
xnor U22981 (N_22981,N_20553,N_20280);
nor U22982 (N_22982,N_21161,N_21436);
xnor U22983 (N_22983,N_21531,N_20639);
or U22984 (N_22984,N_21561,N_21448);
and U22985 (N_22985,N_20954,N_21144);
xnor U22986 (N_22986,N_21298,N_21852);
or U22987 (N_22987,N_21345,N_22481);
and U22988 (N_22988,N_21927,N_20540);
nor U22989 (N_22989,N_21999,N_21502);
nor U22990 (N_22990,N_22145,N_20033);
nand U22991 (N_22991,N_22422,N_20117);
or U22992 (N_22992,N_22315,N_22274);
nor U22993 (N_22993,N_20359,N_20286);
and U22994 (N_22994,N_20272,N_20287);
or U22995 (N_22995,N_22173,N_20857);
or U22996 (N_22996,N_22285,N_21235);
and U22997 (N_22997,N_20869,N_20633);
nand U22998 (N_22998,N_20090,N_21677);
nand U22999 (N_22999,N_21164,N_22234);
and U23000 (N_23000,N_20447,N_20891);
nand U23001 (N_23001,N_22208,N_20089);
nand U23002 (N_23002,N_20025,N_22403);
nor U23003 (N_23003,N_22088,N_20743);
or U23004 (N_23004,N_21660,N_21834);
and U23005 (N_23005,N_20041,N_21504);
nand U23006 (N_23006,N_20831,N_21098);
nor U23007 (N_23007,N_20647,N_21764);
or U23008 (N_23008,N_20180,N_21194);
nand U23009 (N_23009,N_20179,N_20139);
nand U23010 (N_23010,N_20842,N_21397);
and U23011 (N_23011,N_21681,N_21342);
nor U23012 (N_23012,N_20050,N_21280);
nand U23013 (N_23013,N_21538,N_20255);
and U23014 (N_23014,N_20805,N_21704);
and U23015 (N_23015,N_22020,N_21854);
or U23016 (N_23016,N_21791,N_20990);
nor U23017 (N_23017,N_20806,N_21404);
nand U23018 (N_23018,N_20296,N_20477);
or U23019 (N_23019,N_21947,N_21731);
nor U23020 (N_23020,N_21542,N_21582);
or U23021 (N_23021,N_21851,N_21869);
or U23022 (N_23022,N_21387,N_22068);
nand U23023 (N_23023,N_21813,N_21826);
and U23024 (N_23024,N_21177,N_20591);
nand U23025 (N_23025,N_20078,N_21210);
or U23026 (N_23026,N_21043,N_20326);
nand U23027 (N_23027,N_22143,N_20440);
nand U23028 (N_23028,N_20821,N_22460);
or U23029 (N_23029,N_20608,N_22029);
nor U23030 (N_23030,N_22468,N_20396);
nor U23031 (N_23031,N_21799,N_20841);
nor U23032 (N_23032,N_20003,N_21972);
and U23033 (N_23033,N_22052,N_21500);
xor U23034 (N_23034,N_21692,N_22027);
nor U23035 (N_23035,N_20298,N_20631);
nor U23036 (N_23036,N_21967,N_22409);
and U23037 (N_23037,N_20010,N_22105);
xor U23038 (N_23038,N_21858,N_21632);
nor U23039 (N_23039,N_21812,N_20534);
or U23040 (N_23040,N_21483,N_20463);
and U23041 (N_23041,N_21589,N_20343);
or U23042 (N_23042,N_21659,N_20732);
and U23043 (N_23043,N_20790,N_21617);
or U23044 (N_23044,N_21954,N_20278);
or U23045 (N_23045,N_21803,N_20021);
and U23046 (N_23046,N_20978,N_20243);
or U23047 (N_23047,N_20147,N_21696);
nand U23048 (N_23048,N_22449,N_20723);
nor U23049 (N_23049,N_20895,N_22321);
xnor U23050 (N_23050,N_20543,N_20505);
nand U23051 (N_23051,N_21114,N_20454);
nor U23052 (N_23052,N_21683,N_21398);
and U23053 (N_23053,N_21254,N_21075);
and U23054 (N_23054,N_20828,N_20262);
nor U23055 (N_23055,N_21061,N_21039);
xor U23056 (N_23056,N_21479,N_21969);
xor U23057 (N_23057,N_20460,N_22109);
or U23058 (N_23058,N_21067,N_20093);
or U23059 (N_23059,N_20796,N_21762);
and U23060 (N_23060,N_20336,N_22258);
nand U23061 (N_23061,N_21775,N_22365);
nand U23062 (N_23062,N_20698,N_21202);
and U23063 (N_23063,N_20725,N_21066);
nor U23064 (N_23064,N_21705,N_20899);
or U23065 (N_23065,N_21152,N_22212);
or U23066 (N_23066,N_22359,N_20124);
nor U23067 (N_23067,N_20959,N_21421);
or U23068 (N_23068,N_20065,N_22450);
or U23069 (N_23069,N_21476,N_21880);
nor U23070 (N_23070,N_21673,N_21085);
or U23071 (N_23071,N_21380,N_20091);
nor U23072 (N_23072,N_21381,N_21051);
xnor U23073 (N_23073,N_22388,N_20901);
nand U23074 (N_23074,N_22140,N_21914);
or U23075 (N_23075,N_21341,N_22312);
or U23076 (N_23076,N_21310,N_20160);
or U23077 (N_23077,N_20429,N_21305);
and U23078 (N_23078,N_20710,N_20878);
nor U23079 (N_23079,N_21003,N_22307);
xor U23080 (N_23080,N_20678,N_20509);
or U23081 (N_23081,N_21340,N_21093);
or U23082 (N_23082,N_22026,N_20776);
xnor U23083 (N_23083,N_22227,N_20911);
and U23084 (N_23084,N_21685,N_20019);
nor U23085 (N_23085,N_22483,N_20733);
xnor U23086 (N_23086,N_20101,N_22129);
and U23087 (N_23087,N_20219,N_22030);
nand U23088 (N_23088,N_21096,N_22354);
and U23089 (N_23089,N_22065,N_22276);
nor U23090 (N_23090,N_21653,N_20123);
nand U23091 (N_23091,N_21742,N_20835);
nand U23092 (N_23092,N_21264,N_21466);
and U23093 (N_23093,N_22423,N_20087);
nor U23094 (N_23094,N_20770,N_20798);
nand U23095 (N_23095,N_20570,N_22417);
nand U23096 (N_23096,N_20844,N_21604);
nand U23097 (N_23097,N_21642,N_20561);
or U23098 (N_23098,N_20659,N_21796);
or U23099 (N_23099,N_20920,N_21644);
and U23100 (N_23100,N_21169,N_21029);
or U23101 (N_23101,N_20075,N_21410);
nor U23102 (N_23102,N_22002,N_21232);
or U23103 (N_23103,N_22134,N_20417);
and U23104 (N_23104,N_21009,N_21987);
nor U23105 (N_23105,N_21621,N_20407);
nand U23106 (N_23106,N_20996,N_21119);
nand U23107 (N_23107,N_20307,N_20155);
or U23108 (N_23108,N_21088,N_20416);
nand U23109 (N_23109,N_22341,N_20383);
nor U23110 (N_23110,N_20277,N_21755);
or U23111 (N_23111,N_22385,N_21853);
nand U23112 (N_23112,N_20600,N_21983);
nand U23113 (N_23113,N_20185,N_20348);
and U23114 (N_23114,N_21749,N_20594);
or U23115 (N_23115,N_22205,N_21198);
nor U23116 (N_23116,N_20013,N_21671);
or U23117 (N_23117,N_21756,N_20956);
nand U23118 (N_23118,N_21684,N_21536);
and U23119 (N_23119,N_20471,N_22411);
or U23120 (N_23120,N_22062,N_22216);
or U23121 (N_23121,N_21296,N_21700);
and U23122 (N_23122,N_20264,N_21474);
nand U23123 (N_23123,N_21040,N_20236);
nand U23124 (N_23124,N_21139,N_21541);
nor U23125 (N_23125,N_20609,N_22176);
and U23126 (N_23126,N_21495,N_21509);
and U23127 (N_23127,N_21669,N_20031);
or U23128 (N_23128,N_20045,N_21068);
or U23129 (N_23129,N_20112,N_22032);
xnor U23130 (N_23130,N_20247,N_20717);
and U23131 (N_23131,N_21992,N_22424);
xnor U23132 (N_23132,N_20294,N_22048);
xor U23133 (N_23133,N_22459,N_21411);
nand U23134 (N_23134,N_22045,N_21289);
nand U23135 (N_23135,N_21147,N_20731);
nand U23136 (N_23136,N_21205,N_21382);
and U23137 (N_23137,N_20491,N_22054);
and U23138 (N_23138,N_20697,N_21979);
nor U23139 (N_23139,N_22399,N_20459);
and U23140 (N_23140,N_21975,N_20503);
nand U23141 (N_23141,N_22214,N_20456);
and U23142 (N_23142,N_20354,N_22410);
nand U23143 (N_23143,N_20993,N_20754);
or U23144 (N_23144,N_22233,N_21748);
or U23145 (N_23145,N_21011,N_20741);
and U23146 (N_23146,N_20952,N_20178);
nand U23147 (N_23147,N_21450,N_21777);
and U23148 (N_23148,N_20644,N_22050);
and U23149 (N_23149,N_22240,N_22488);
nor U23150 (N_23150,N_21633,N_21336);
nand U23151 (N_23151,N_20986,N_20249);
nor U23152 (N_23152,N_20890,N_21420);
nand U23153 (N_23153,N_20579,N_21277);
nor U23154 (N_23154,N_20628,N_20566);
and U23155 (N_23155,N_21216,N_20820);
nand U23156 (N_23156,N_21497,N_20175);
nor U23157 (N_23157,N_20624,N_21062);
nand U23158 (N_23158,N_21787,N_21730);
xnor U23159 (N_23159,N_21601,N_21449);
nor U23160 (N_23160,N_22142,N_22195);
nand U23161 (N_23161,N_22099,N_20894);
and U23162 (N_23162,N_20266,N_22418);
and U23163 (N_23163,N_21903,N_21695);
nor U23164 (N_23164,N_21959,N_21895);
nand U23165 (N_23165,N_22179,N_21971);
or U23166 (N_23166,N_20616,N_20635);
nor U23167 (N_23167,N_22395,N_20475);
or U23168 (N_23168,N_21578,N_21652);
nor U23169 (N_23169,N_22382,N_22275);
or U23170 (N_23170,N_21459,N_22194);
nor U23171 (N_23171,N_20966,N_22127);
nand U23172 (N_23172,N_20685,N_20069);
nand U23173 (N_23173,N_21751,N_21229);
and U23174 (N_23174,N_21461,N_21499);
and U23175 (N_23175,N_22310,N_20052);
and U23176 (N_23176,N_21598,N_20855);
or U23177 (N_23177,N_20482,N_21613);
and U23178 (N_23178,N_21362,N_20612);
and U23179 (N_23179,N_20167,N_22000);
nor U23180 (N_23180,N_20664,N_21636);
nor U23181 (N_23181,N_21103,N_21513);
nor U23182 (N_23182,N_21283,N_22330);
nand U23183 (N_23183,N_21527,N_21314);
xnor U23184 (N_23184,N_20120,N_20283);
and U23185 (N_23185,N_20254,N_22368);
and U23186 (N_23186,N_21957,N_21532);
or U23187 (N_23187,N_20306,N_21600);
nor U23188 (N_23188,N_20291,N_20656);
xnor U23189 (N_23189,N_20606,N_20308);
or U23190 (N_23190,N_20728,N_22380);
or U23191 (N_23191,N_22338,N_20186);
nor U23192 (N_23192,N_22147,N_20328);
nor U23193 (N_23193,N_21464,N_20039);
or U23194 (N_23194,N_22028,N_21311);
nor U23195 (N_23195,N_21438,N_22290);
or U23196 (N_23196,N_21554,N_21550);
nor U23197 (N_23197,N_20645,N_21890);
or U23198 (N_23198,N_20908,N_20273);
nor U23199 (N_23199,N_22017,N_20513);
and U23200 (N_23200,N_22169,N_21587);
or U23201 (N_23201,N_22394,N_20035);
nand U23202 (N_23202,N_20182,N_22498);
and U23203 (N_23203,N_22213,N_20372);
nand U23204 (N_23204,N_21616,N_21836);
xor U23205 (N_23205,N_22335,N_20769);
and U23206 (N_23206,N_20968,N_21786);
xnor U23207 (N_23207,N_21912,N_21492);
or U23208 (N_23208,N_20140,N_21172);
and U23209 (N_23209,N_21007,N_20250);
and U23210 (N_23210,N_20414,N_20366);
nand U23211 (N_23211,N_22247,N_22185);
xnor U23212 (N_23212,N_20988,N_22306);
or U23213 (N_23213,N_22389,N_20497);
and U23214 (N_23214,N_20814,N_21425);
and U23215 (N_23215,N_20325,N_22031);
or U23216 (N_23216,N_20595,N_22070);
or U23217 (N_23217,N_20063,N_20099);
or U23218 (N_23218,N_22420,N_22466);
or U23219 (N_23219,N_20418,N_21330);
nor U23220 (N_23220,N_21757,N_20514);
or U23221 (N_23221,N_20448,N_21733);
nor U23222 (N_23222,N_21217,N_22333);
or U23223 (N_23223,N_20593,N_20948);
or U23224 (N_23224,N_22007,N_20765);
nand U23225 (N_23225,N_20480,N_20061);
or U23226 (N_23226,N_20652,N_21711);
nor U23227 (N_23227,N_21019,N_22479);
or U23228 (N_23228,N_20654,N_20532);
or U23229 (N_23229,N_21458,N_21183);
xor U23230 (N_23230,N_21256,N_22230);
nand U23231 (N_23231,N_21489,N_22291);
xnor U23232 (N_23232,N_21218,N_21637);
nor U23233 (N_23233,N_22005,N_20364);
nor U23234 (N_23234,N_21309,N_21145);
nor U23235 (N_23235,N_21493,N_20176);
or U23236 (N_23236,N_22297,N_21930);
nor U23237 (N_23237,N_21706,N_20519);
nand U23238 (N_23238,N_21452,N_21469);
nor U23239 (N_23239,N_21125,N_22204);
or U23240 (N_23240,N_22461,N_20630);
or U23241 (N_23241,N_22490,N_21645);
nand U23242 (N_23242,N_21566,N_21375);
or U23243 (N_23243,N_20351,N_20522);
nor U23244 (N_23244,N_20302,N_22115);
xnor U23245 (N_23245,N_20761,N_22038);
nor U23246 (N_23246,N_22257,N_21916);
and U23247 (N_23247,N_21620,N_22112);
nand U23248 (N_23248,N_21447,N_22128);
or U23249 (N_23249,N_22373,N_21297);
nand U23250 (N_23250,N_20119,N_21878);
nor U23251 (N_23251,N_21242,N_21934);
nand U23252 (N_23252,N_21248,N_21898);
and U23253 (N_23253,N_20535,N_21597);
and U23254 (N_23254,N_21629,N_20946);
nor U23255 (N_23255,N_22469,N_20465);
nand U23256 (N_23256,N_20339,N_20057);
and U23257 (N_23257,N_20240,N_20793);
nor U23258 (N_23258,N_21128,N_20256);
nor U23259 (N_23259,N_22131,N_21693);
or U23260 (N_23260,N_20103,N_22146);
nand U23261 (N_23261,N_22010,N_20439);
and U23262 (N_23262,N_21965,N_21689);
or U23263 (N_23263,N_21347,N_20585);
xnor U23264 (N_23264,N_22480,N_22089);
and U23265 (N_23265,N_20148,N_22241);
nand U23266 (N_23266,N_20173,N_21654);
nor U23267 (N_23267,N_21760,N_20808);
and U23268 (N_23268,N_22473,N_21635);
nand U23269 (N_23269,N_20640,N_21804);
xnor U23270 (N_23270,N_21023,N_21031);
nand U23271 (N_23271,N_21792,N_21366);
nor U23272 (N_23272,N_21416,N_22165);
and U23273 (N_23273,N_21823,N_21995);
nor U23274 (N_23274,N_20170,N_21034);
or U23275 (N_23275,N_21344,N_22008);
and U23276 (N_23276,N_20716,N_21797);
nor U23277 (N_23277,N_22012,N_21703);
xnor U23278 (N_23278,N_21033,N_22016);
nand U23279 (N_23279,N_21412,N_22281);
or U23280 (N_23280,N_21166,N_21866);
and U23281 (N_23281,N_21808,N_21135);
or U23282 (N_23282,N_20861,N_21195);
or U23283 (N_23283,N_21281,N_20642);
and U23284 (N_23284,N_21130,N_21667);
or U23285 (N_23285,N_21801,N_21187);
nor U23286 (N_23286,N_21259,N_20121);
or U23287 (N_23287,N_20816,N_22378);
xnor U23288 (N_23288,N_20331,N_20550);
or U23289 (N_23289,N_20408,N_20682);
xnor U23290 (N_23290,N_20560,N_22405);
nand U23291 (N_23291,N_20643,N_21944);
or U23292 (N_23292,N_22077,N_20567);
and U23293 (N_23293,N_20555,N_20073);
or U23294 (N_23294,N_21221,N_21393);
and U23295 (N_23295,N_22116,N_20775);
and U23296 (N_23296,N_20742,N_22496);
or U23297 (N_23297,N_20748,N_21752);
nor U23298 (N_23298,N_22344,N_21267);
and U23299 (N_23299,N_21640,N_21022);
xor U23300 (N_23300,N_21318,N_20887);
xor U23301 (N_23301,N_22429,N_21286);
and U23302 (N_23302,N_21723,N_21850);
nand U23303 (N_23303,N_21618,N_22066);
xor U23304 (N_23304,N_21958,N_21078);
nand U23305 (N_23305,N_20533,N_20053);
nor U23306 (N_23306,N_21159,N_22340);
or U23307 (N_23307,N_21996,N_22254);
nand U23308 (N_23308,N_21845,N_20488);
nor U23309 (N_23309,N_22304,N_22073);
nand U23310 (N_23310,N_20985,N_21906);
nor U23311 (N_23311,N_21602,N_20301);
xor U23312 (N_23312,N_20521,N_21049);
xnor U23313 (N_23313,N_21743,N_20401);
and U23314 (N_23314,N_21624,N_21842);
or U23315 (N_23315,N_21148,N_20746);
nand U23316 (N_23316,N_20791,N_22152);
and U23317 (N_23317,N_22482,N_21829);
nand U23318 (N_23318,N_21966,N_22170);
xnor U23319 (N_23319,N_20201,N_20449);
and U23320 (N_23320,N_21761,N_22014);
or U23321 (N_23321,N_20651,N_20856);
or U23322 (N_23322,N_21800,N_20394);
nand U23323 (N_23323,N_21165,N_21921);
and U23324 (N_23324,N_20792,N_20229);
or U23325 (N_23325,N_20740,N_20340);
nand U23326 (N_23326,N_20067,N_22033);
nand U23327 (N_23327,N_20563,N_21288);
and U23328 (N_23328,N_20072,N_20445);
xor U23329 (N_23329,N_21237,N_21771);
nor U23330 (N_23330,N_20305,N_21323);
nand U23331 (N_23331,N_20711,N_21938);
xnor U23332 (N_23332,N_22123,N_20402);
xor U23333 (N_23333,N_21444,N_21848);
nor U23334 (N_23334,N_20008,N_20134);
nand U23335 (N_23335,N_20269,N_20344);
and U23336 (N_23336,N_21463,N_21274);
xor U23337 (N_23337,N_22475,N_21584);
and U23338 (N_23338,N_20916,N_22161);
xnor U23339 (N_23339,N_22006,N_21549);
and U23340 (N_23340,N_20190,N_21010);
nand U23341 (N_23341,N_20607,N_20549);
xor U23342 (N_23342,N_21713,N_21810);
nor U23343 (N_23343,N_22406,N_21630);
and U23344 (N_23344,N_21255,N_21535);
and U23345 (N_23345,N_20241,N_21084);
nand U23346 (N_23346,N_22280,N_21262);
nand U23347 (N_23347,N_21817,N_22167);
nor U23348 (N_23348,N_20111,N_21465);
or U23349 (N_23349,N_20795,N_21581);
xnor U23350 (N_23350,N_20548,N_21875);
xnor U23351 (N_23351,N_20589,N_20494);
and U23352 (N_23352,N_20940,N_21772);
nand U23353 (N_23353,N_20507,N_22155);
nand U23354 (N_23354,N_20450,N_20662);
xnor U23355 (N_23355,N_20755,N_20767);
and U23356 (N_23356,N_21178,N_20358);
nand U23357 (N_23357,N_20832,N_20376);
or U23358 (N_23358,N_20672,N_21970);
or U23359 (N_23359,N_21690,N_21896);
and U23360 (N_23360,N_20687,N_20876);
nor U23361 (N_23361,N_22261,N_21717);
nor U23362 (N_23362,N_21056,N_20979);
nand U23363 (N_23363,N_21231,N_21021);
nor U23364 (N_23364,N_20316,N_20794);
nand U23365 (N_23365,N_22494,N_22305);
nand U23366 (N_23366,N_21435,N_21805);
nor U23367 (N_23367,N_20699,N_21715);
or U23368 (N_23368,N_21913,N_21354);
xnor U23369 (N_23369,N_21454,N_20228);
and U23370 (N_23370,N_20037,N_20265);
nor U23371 (N_23371,N_22433,N_21239);
nand U23372 (N_23372,N_20428,N_21894);
nand U23373 (N_23373,N_21941,N_21867);
nor U23374 (N_23374,N_21811,N_20817);
nor U23375 (N_23375,N_20251,N_21889);
xnor U23376 (N_23376,N_20552,N_21643);
xor U23377 (N_23377,N_20174,N_20285);
nor U23378 (N_23378,N_21109,N_21045);
or U23379 (N_23379,N_22200,N_20690);
nor U23380 (N_23380,N_21865,N_20442);
nor U23381 (N_23381,N_21037,N_21047);
nor U23382 (N_23382,N_21557,N_20314);
xnor U23383 (N_23383,N_21841,N_20724);
nor U23384 (N_23384,N_21820,N_20311);
and U23385 (N_23385,N_22162,N_20373);
or U23386 (N_23386,N_22347,N_20848);
and U23387 (N_23387,N_20238,N_20432);
xnor U23388 (N_23388,N_20889,N_20867);
or U23389 (N_23389,N_21238,N_20845);
xnor U23390 (N_23390,N_22025,N_20658);
or U23391 (N_23391,N_21988,N_21153);
nor U23392 (N_23392,N_21529,N_20487);
nand U23393 (N_23393,N_20836,N_22039);
nor U23394 (N_23394,N_22059,N_21871);
or U23395 (N_23395,N_22150,N_20038);
xnor U23396 (N_23396,N_21149,N_22223);
nand U23397 (N_23397,N_21623,N_22319);
or U23398 (N_23398,N_20410,N_22323);
or U23399 (N_23399,N_21041,N_20034);
nor U23400 (N_23400,N_22282,N_21824);
nand U23401 (N_23401,N_21013,N_22313);
and U23402 (N_23402,N_20151,N_22080);
nand U23403 (N_23403,N_20787,N_21910);
and U23404 (N_23404,N_21608,N_20838);
or U23405 (N_23405,N_21523,N_20203);
and U23406 (N_23406,N_21945,N_21050);
and U23407 (N_23407,N_21917,N_22327);
or U23408 (N_23408,N_21307,N_21552);
nor U23409 (N_23409,N_20701,N_22349);
nand U23410 (N_23410,N_20520,N_20614);
nand U23411 (N_23411,N_20225,N_21117);
and U23412 (N_23412,N_21121,N_20581);
and U23413 (N_23413,N_21846,N_20164);
and U23414 (N_23414,N_21868,N_21275);
and U23415 (N_23415,N_21215,N_21055);
nor U23416 (N_23416,N_20933,N_21185);
or U23417 (N_23417,N_21687,N_21572);
xnor U23418 (N_23418,N_21451,N_20526);
and U23419 (N_23419,N_21496,N_20115);
and U23420 (N_23420,N_20707,N_21991);
nor U23421 (N_23421,N_20136,N_22272);
or U23422 (N_23422,N_20338,N_20279);
nor U23423 (N_23423,N_21312,N_21899);
nand U23424 (N_23424,N_20969,N_21559);
nand U23425 (N_23425,N_22078,N_20572);
nor U23426 (N_23426,N_20347,N_21374);
nor U23427 (N_23427,N_21556,N_20925);
nor U23428 (N_23428,N_21044,N_20973);
or U23429 (N_23429,N_20094,N_20753);
xnor U23430 (N_23430,N_20142,N_20896);
or U23431 (N_23431,N_21367,N_20318);
nand U23432 (N_23432,N_21429,N_22251);
xnor U23433 (N_23433,N_20196,N_22198);
nand U23434 (N_23434,N_21104,N_22260);
nand U23435 (N_23435,N_22236,N_20669);
and U23436 (N_23436,N_21856,N_22398);
nor U23437 (N_23437,N_20558,N_20495);
or U23438 (N_23438,N_22351,N_20786);
nand U23439 (N_23439,N_21099,N_21257);
and U23440 (N_23440,N_21027,N_22160);
nand U23441 (N_23441,N_21515,N_21940);
nand U23442 (N_23442,N_21017,N_22051);
and U23443 (N_23443,N_20623,N_20995);
or U23444 (N_23444,N_21395,N_20726);
or U23445 (N_23445,N_22149,N_21664);
and U23446 (N_23446,N_22209,N_22067);
nor U23447 (N_23447,N_22064,N_20319);
nor U23448 (N_23448,N_20330,N_20489);
and U23449 (N_23449,N_20839,N_21349);
and U23450 (N_23450,N_20991,N_20759);
and U23451 (N_23451,N_20501,N_21245);
nand U23452 (N_23452,N_20149,N_22296);
nor U23453 (N_23453,N_20369,N_21827);
or U23454 (N_23454,N_20257,N_22148);
xnor U23455 (N_23455,N_20425,N_21840);
nand U23456 (N_23456,N_22228,N_20671);
and U23457 (N_23457,N_20871,N_20977);
or U23458 (N_23458,N_20860,N_20504);
xor U23459 (N_23459,N_20712,N_20310);
or U23460 (N_23460,N_21830,N_20409);
nand U23461 (N_23461,N_22372,N_21059);
xnor U23462 (N_23462,N_21176,N_22047);
nor U23463 (N_23463,N_20126,N_21763);
nor U23464 (N_23464,N_21191,N_20207);
nand U23465 (N_23465,N_20762,N_22210);
nand U23466 (N_23466,N_21759,N_22138);
nor U23467 (N_23467,N_21694,N_21456);
or U23468 (N_23468,N_21372,N_22311);
and U23469 (N_23469,N_20749,N_21090);
nand U23470 (N_23470,N_22202,N_21008);
nor U23471 (N_23471,N_20650,N_21102);
nand U23472 (N_23472,N_21976,N_20863);
xnor U23473 (N_23473,N_20437,N_22183);
or U23474 (N_23474,N_22024,N_21192);
nand U23475 (N_23475,N_21364,N_21320);
nor U23476 (N_23476,N_20209,N_20004);
nor U23477 (N_23477,N_22221,N_21951);
and U23478 (N_23478,N_21327,N_22301);
and U23479 (N_23479,N_20036,N_22396);
nand U23480 (N_23480,N_22309,N_20909);
nor U23481 (N_23481,N_20322,N_21514);
or U23482 (N_23482,N_21503,N_20017);
and U23483 (N_23483,N_20949,N_21625);
nor U23484 (N_23484,N_20997,N_20127);
and U23485 (N_23485,N_20131,N_20807);
nor U23486 (N_23486,N_20937,N_22308);
nor U23487 (N_23487,N_20345,N_20803);
nor U23488 (N_23488,N_21140,N_21729);
or U23489 (N_23489,N_20833,N_21250);
or U23490 (N_23490,N_22407,N_21468);
and U23491 (N_23491,N_22222,N_20095);
or U23492 (N_23492,N_22269,N_20399);
xor U23493 (N_23493,N_21460,N_20739);
or U23494 (N_23494,N_22364,N_21377);
nand U23495 (N_23495,N_21424,N_20537);
nand U23496 (N_23496,N_22100,N_22287);
and U23497 (N_23497,N_21989,N_21553);
nor U23498 (N_23498,N_21641,N_22242);
nor U23499 (N_23499,N_20068,N_21227);
nand U23500 (N_23500,N_21032,N_20705);
nor U23501 (N_23501,N_20692,N_21132);
or U23502 (N_23502,N_21413,N_21064);
nor U23503 (N_23503,N_20826,N_20390);
nor U23504 (N_23504,N_22470,N_20125);
xnor U23505 (N_23505,N_20758,N_20215);
nor U23506 (N_23506,N_22266,N_21785);
nor U23507 (N_23507,N_20132,N_21136);
and U23508 (N_23508,N_20118,N_22413);
xnor U23509 (N_23509,N_21981,N_20597);
xnor U23510 (N_23510,N_20615,N_21196);
and U23511 (N_23511,N_20380,N_21179);
nor U23512 (N_23512,N_22081,N_20989);
and U23513 (N_23513,N_22207,N_21386);
nor U23514 (N_23514,N_21888,N_20202);
nor U23515 (N_23515,N_20499,N_21672);
nand U23516 (N_23516,N_20226,N_20290);
and U23517 (N_23517,N_20163,N_22076);
and U23518 (N_23518,N_20665,N_21278);
nand U23519 (N_23519,N_21437,N_22426);
and U23520 (N_23520,N_21439,N_22118);
or U23521 (N_23521,N_20866,N_20942);
nor U23522 (N_23522,N_20109,N_21302);
and U23523 (N_23523,N_20412,N_22190);
nand U23524 (N_23524,N_21605,N_20029);
and U23525 (N_23525,N_21365,N_20747);
xor U23526 (N_23526,N_22278,N_20622);
or U23527 (N_23527,N_21946,N_22180);
nand U23528 (N_23528,N_21236,N_21592);
or U23529 (N_23529,N_20892,N_21212);
nor U23530 (N_23530,N_21181,N_20438);
nor U23531 (N_23531,N_21893,N_22392);
and U23532 (N_23532,N_21766,N_20468);
xor U23533 (N_23533,N_22193,N_20381);
and U23534 (N_23534,N_21544,N_22085);
nor U23535 (N_23535,N_22331,N_20653);
and U23536 (N_23536,N_20472,N_20960);
or U23537 (N_23537,N_20557,N_22348);
nor U23538 (N_23538,N_20135,N_21112);
xor U23539 (N_23539,N_21015,N_21802);
or U23540 (N_23540,N_22284,N_20929);
nor U23541 (N_23541,N_22137,N_20047);
xnor U23542 (N_23542,N_22337,N_20706);
and U23543 (N_23543,N_21470,N_20054);
and U23544 (N_23544,N_20066,N_22377);
nand U23545 (N_23545,N_21962,N_20981);
nor U23546 (N_23546,N_21269,N_20834);
nand U23547 (N_23547,N_20205,N_21303);
nor U23548 (N_23548,N_20161,N_22455);
nand U23549 (N_23549,N_20009,N_22267);
or U23550 (N_23550,N_21244,N_20603);
or U23551 (N_23551,N_20370,N_22239);
and U23552 (N_23552,N_21519,N_22256);
nand U23553 (N_23553,N_21990,N_20512);
or U23554 (N_23554,N_21507,N_22250);
nor U23555 (N_23555,N_20825,N_20064);
nor U23556 (N_23556,N_20626,N_21170);
nor U23557 (N_23557,N_20804,N_21220);
nand U23558 (N_23558,N_21714,N_20930);
or U23559 (N_23559,N_21528,N_20248);
nor U23560 (N_23560,N_21272,N_20270);
nand U23561 (N_23561,N_22079,N_21348);
and U23562 (N_23562,N_22224,N_20898);
or U23563 (N_23563,N_20473,N_22421);
and U23564 (N_23564,N_20917,N_20014);
nor U23565 (N_23565,N_22248,N_21079);
xnor U23566 (N_23566,N_20605,N_21984);
nand U23567 (N_23567,N_20772,N_21002);
nand U23568 (N_23568,N_21758,N_22141);
and U23569 (N_23569,N_21746,N_20544);
xnor U23570 (N_23570,N_21877,N_22355);
nand U23571 (N_23571,N_20329,N_21902);
nand U23572 (N_23572,N_20904,N_20222);
nand U23573 (N_23573,N_20084,N_22035);
and U23574 (N_23574,N_22111,N_21122);
nor U23575 (N_23575,N_20551,N_21065);
or U23576 (N_23576,N_21133,N_22090);
and U23577 (N_23577,N_20531,N_22369);
nor U23578 (N_23578,N_22286,N_20815);
and U23579 (N_23579,N_20261,N_20708);
xor U23580 (N_23580,N_20518,N_20900);
or U23581 (N_23581,N_21961,N_20085);
nand U23582 (N_23582,N_20847,N_20105);
xor U23583 (N_23583,N_21313,N_22430);
nand U23584 (N_23584,N_21024,N_20945);
nand U23585 (N_23585,N_21160,N_22362);
xor U23586 (N_23586,N_21355,N_21143);
nor U23587 (N_23587,N_21265,N_20349);
or U23588 (N_23588,N_21343,N_22375);
or U23589 (N_23589,N_21929,N_22384);
nand U23590 (N_23590,N_21882,N_22106);
nand U23591 (N_23591,N_20666,N_20625);
and U23592 (N_23592,N_22342,N_21779);
and U23593 (N_23593,N_20693,N_21886);
and U23594 (N_23594,N_22206,N_20481);
or U23595 (N_23595,N_20082,N_22053);
nor U23596 (N_23596,N_22086,N_22096);
or U23597 (N_23597,N_20317,N_22446);
nor U23598 (N_23598,N_21750,N_21052);
nor U23599 (N_23599,N_22401,N_22472);
nor U23600 (N_23600,N_21263,N_21270);
and U23601 (N_23601,N_22474,N_22454);
or U23602 (N_23602,N_21146,N_20443);
and U23603 (N_23603,N_21113,N_20618);
and U23604 (N_23604,N_21831,N_22126);
nand U23605 (N_23605,N_21401,N_20191);
nand U23606 (N_23606,N_22074,N_20837);
nor U23607 (N_23607,N_21184,N_20781);
or U23608 (N_23608,N_21974,N_21780);
or U23609 (N_23609,N_22245,N_20944);
xor U23610 (N_23610,N_20502,N_20389);
nand U23611 (N_23611,N_21724,N_21025);
and U23612 (N_23612,N_20044,N_22009);
nor U23613 (N_23613,N_21814,N_21405);
or U23614 (N_23614,N_20620,N_21392);
nand U23615 (N_23615,N_21299,N_21679);
nand U23616 (N_23616,N_20361,N_22177);
or U23617 (N_23617,N_20387,N_20171);
nor U23618 (N_23618,N_22098,N_20721);
or U23619 (N_23619,N_21665,N_21036);
nand U23620 (N_23620,N_20691,N_21891);
or U23621 (N_23621,N_21691,N_21427);
xor U23622 (N_23622,N_21335,N_20404);
and U23623 (N_23623,N_20660,N_21828);
nor U23624 (N_23624,N_20096,N_21697);
nand U23625 (N_23625,N_22201,N_20870);
or U23626 (N_23626,N_22328,N_21388);
nand U23627 (N_23627,N_21129,N_22124);
or U23628 (N_23628,N_20738,N_21186);
xnor U23629 (N_23629,N_21662,N_22299);
nand U23630 (N_23630,N_20777,N_22464);
or U23631 (N_23631,N_20400,N_21083);
or U23632 (N_23632,N_21569,N_22211);
or U23633 (N_23633,N_20083,N_20335);
and U23634 (N_23634,N_20496,N_21110);
nand U23635 (N_23635,N_21433,N_20059);
or U23636 (N_23636,N_22117,N_22019);
and U23637 (N_23637,N_21107,N_20525);
nand U23638 (N_23638,N_20604,N_21328);
nand U23639 (N_23639,N_20684,N_20368);
and U23640 (N_23640,N_20431,N_20703);
nand U23641 (N_23641,N_20573,N_21271);
nor U23642 (N_23642,N_20055,N_20802);
nand U23643 (N_23643,N_21876,N_20700);
nor U23644 (N_23644,N_20187,N_20362);
or U23645 (N_23645,N_22135,N_20778);
nor U23646 (N_23646,N_21006,N_22139);
and U23647 (N_23647,N_21534,N_20915);
or U23648 (N_23648,N_21389,N_22345);
nor U23649 (N_23649,N_21485,N_22350);
and U23650 (N_23650,N_20565,N_21197);
nor U23651 (N_23651,N_20000,N_22196);
and U23652 (N_23652,N_20210,N_22154);
or U23653 (N_23653,N_22402,N_22371);
xnor U23654 (N_23654,N_20864,N_20932);
and U23655 (N_23655,N_21520,N_20688);
nor U23656 (N_23656,N_22018,N_21740);
or U23657 (N_23657,N_21833,N_21127);
or U23658 (N_23658,N_21682,N_20964);
nand U23659 (N_23659,N_21948,N_20292);
nor U23660 (N_23660,N_22188,N_20751);
nor U23661 (N_23661,N_21240,N_21563);
nor U23662 (N_23662,N_21956,N_22186);
nand U23663 (N_23663,N_21287,N_21070);
nand U23664 (N_23664,N_21712,N_21402);
nand U23665 (N_23665,N_20433,N_22015);
or U23666 (N_23666,N_21936,N_21594);
and U23667 (N_23667,N_22467,N_20927);
and U23668 (N_23668,N_22022,N_21964);
nand U23669 (N_23669,N_21337,N_20984);
xor U23670 (N_23670,N_20079,N_21788);
and U23671 (N_23671,N_21276,N_21861);
and U23672 (N_23672,N_20211,N_20689);
nor U23673 (N_23673,N_20827,N_21558);
or U23674 (N_23674,N_20872,N_21339);
nand U23675 (N_23675,N_20321,N_20801);
nand U23676 (N_23676,N_21352,N_21072);
nand U23677 (N_23677,N_22431,N_21077);
and U23678 (N_23678,N_21173,N_20046);
or U23679 (N_23679,N_20874,N_21603);
xnor U23680 (N_23680,N_22404,N_21467);
and U23681 (N_23681,N_20715,N_21284);
nor U23682 (N_23682,N_21334,N_20576);
and U23683 (N_23683,N_20931,N_20001);
nand U23684 (N_23684,N_20212,N_20886);
or U23685 (N_23685,N_20478,N_20150);
xor U23686 (N_23686,N_21462,N_20695);
nor U23687 (N_23687,N_22130,N_22163);
xor U23688 (N_23688,N_20648,N_21634);
xnor U23689 (N_23689,N_21567,N_20086);
nand U23690 (N_23690,N_21767,N_22253);
nand U23691 (N_23691,N_21291,N_21753);
or U23692 (N_23692,N_20873,N_21346);
or U23693 (N_23693,N_21162,N_21707);
nand U23694 (N_23694,N_21596,N_20230);
and U23695 (N_23695,N_22023,N_20592);
nand U23696 (N_23696,N_21030,N_20779);
xor U23697 (N_23697,N_20275,N_20223);
nand U23698 (N_23698,N_20982,N_20341);
xor U23699 (N_23699,N_22164,N_22447);
and U23700 (N_23700,N_20918,N_20849);
xor U23701 (N_23701,N_22094,N_20384);
xnor U23702 (N_23702,N_22391,N_21905);
and U23703 (N_23703,N_22374,N_21371);
nand U23704 (N_23704,N_20686,N_20598);
nand U23705 (N_23705,N_22415,N_20818);
nand U23706 (N_23706,N_21498,N_20884);
nor U23707 (N_23707,N_22414,N_20885);
or U23708 (N_23708,N_21835,N_20922);
or U23709 (N_23709,N_20382,N_20851);
or U23710 (N_23710,N_21012,N_20367);
or U23711 (N_23711,N_21607,N_21727);
nand U23712 (N_23712,N_21522,N_20613);
nor U23713 (N_23713,N_22289,N_20829);
or U23714 (N_23714,N_21378,N_21279);
nand U23715 (N_23715,N_20355,N_21333);
and U23716 (N_23716,N_21925,N_20268);
and U23717 (N_23717,N_22283,N_20081);
and U23718 (N_23718,N_21676,N_20719);
nand U23719 (N_23719,N_22226,N_20679);
nand U23720 (N_23720,N_20216,N_22097);
xor U23721 (N_23721,N_21234,N_20498);
nand U23722 (N_23722,N_20663,N_22061);
and U23723 (N_23723,N_20159,N_21266);
nand U23724 (N_23724,N_22092,N_22229);
and U23725 (N_23725,N_21568,N_20634);
nand U23726 (N_23726,N_22477,N_21356);
nor U23727 (N_23727,N_20315,N_20106);
and U23728 (N_23728,N_20441,N_22003);
or U23729 (N_23729,N_21151,N_21361);
nand U23730 (N_23730,N_20100,N_21555);
nor U23731 (N_23731,N_20457,N_20363);
nand U23732 (N_23732,N_21583,N_21721);
nor U23733 (N_23733,N_22058,N_20007);
or U23734 (N_23734,N_20637,N_22041);
and U23735 (N_23735,N_20527,N_20737);
nand U23736 (N_23736,N_21795,N_20822);
nand U23737 (N_23737,N_21661,N_21111);
or U23738 (N_23738,N_21907,N_20194);
or U23739 (N_23739,N_20113,N_20474);
or U23740 (N_23740,N_20921,N_21390);
nor U23741 (N_23741,N_22381,N_21091);
nand U23742 (N_23742,N_21261,N_21322);
xnor U23743 (N_23743,N_21057,N_22360);
and U23744 (N_23744,N_22334,N_20137);
nand U23745 (N_23745,N_21357,N_20493);
and U23746 (N_23746,N_20768,N_20617);
and U23747 (N_23747,N_20992,N_20304);
or U23748 (N_23748,N_20602,N_22249);
or U23749 (N_23749,N_22120,N_20071);
or U23750 (N_23750,N_22108,N_20351);
nor U23751 (N_23751,N_21842,N_20527);
nor U23752 (N_23752,N_22042,N_21678);
xor U23753 (N_23753,N_20757,N_22150);
and U23754 (N_23754,N_20519,N_21337);
and U23755 (N_23755,N_21398,N_22398);
or U23756 (N_23756,N_21167,N_21747);
nand U23757 (N_23757,N_22315,N_20167);
or U23758 (N_23758,N_21344,N_21453);
or U23759 (N_23759,N_22374,N_20540);
nor U23760 (N_23760,N_20594,N_21142);
xor U23761 (N_23761,N_20060,N_20644);
and U23762 (N_23762,N_20132,N_22050);
and U23763 (N_23763,N_21257,N_21806);
nor U23764 (N_23764,N_21757,N_21131);
nand U23765 (N_23765,N_20922,N_22488);
and U23766 (N_23766,N_21586,N_22227);
xor U23767 (N_23767,N_20909,N_20359);
or U23768 (N_23768,N_20987,N_22234);
and U23769 (N_23769,N_20098,N_20585);
and U23770 (N_23770,N_21185,N_20303);
nand U23771 (N_23771,N_20091,N_22173);
nand U23772 (N_23772,N_22249,N_21984);
nand U23773 (N_23773,N_21185,N_22065);
or U23774 (N_23774,N_21630,N_21896);
and U23775 (N_23775,N_20487,N_21980);
or U23776 (N_23776,N_21869,N_20892);
and U23777 (N_23777,N_21407,N_21457);
nor U23778 (N_23778,N_21718,N_22343);
xor U23779 (N_23779,N_21167,N_21171);
nor U23780 (N_23780,N_21899,N_21418);
or U23781 (N_23781,N_20342,N_21996);
nand U23782 (N_23782,N_21133,N_20128);
nand U23783 (N_23783,N_21314,N_22066);
nand U23784 (N_23784,N_20636,N_21926);
and U23785 (N_23785,N_21485,N_20894);
or U23786 (N_23786,N_20009,N_21635);
nand U23787 (N_23787,N_20553,N_20977);
nor U23788 (N_23788,N_21140,N_21645);
nor U23789 (N_23789,N_20116,N_22104);
nand U23790 (N_23790,N_20854,N_21842);
nand U23791 (N_23791,N_20749,N_21249);
nor U23792 (N_23792,N_20393,N_22181);
xnor U23793 (N_23793,N_21441,N_21573);
nor U23794 (N_23794,N_21513,N_21453);
nor U23795 (N_23795,N_22099,N_21696);
nand U23796 (N_23796,N_20017,N_22225);
and U23797 (N_23797,N_21068,N_21681);
or U23798 (N_23798,N_21970,N_20452);
and U23799 (N_23799,N_21672,N_21562);
xor U23800 (N_23800,N_21297,N_20648);
and U23801 (N_23801,N_22060,N_21600);
or U23802 (N_23802,N_21605,N_21457);
nor U23803 (N_23803,N_21946,N_20706);
and U23804 (N_23804,N_20557,N_21066);
nor U23805 (N_23805,N_22399,N_20921);
and U23806 (N_23806,N_20494,N_22096);
nand U23807 (N_23807,N_21831,N_22487);
or U23808 (N_23808,N_20789,N_21161);
nor U23809 (N_23809,N_21448,N_21357);
nand U23810 (N_23810,N_20701,N_20625);
nor U23811 (N_23811,N_20579,N_20067);
nand U23812 (N_23812,N_21917,N_21827);
nor U23813 (N_23813,N_21414,N_20964);
or U23814 (N_23814,N_22117,N_20816);
nand U23815 (N_23815,N_21572,N_20751);
or U23816 (N_23816,N_22276,N_22278);
nand U23817 (N_23817,N_21982,N_21533);
nand U23818 (N_23818,N_20317,N_21483);
nor U23819 (N_23819,N_20547,N_20966);
nand U23820 (N_23820,N_21822,N_21337);
or U23821 (N_23821,N_22250,N_22481);
and U23822 (N_23822,N_21630,N_20850);
or U23823 (N_23823,N_20472,N_21608);
or U23824 (N_23824,N_20087,N_21725);
xor U23825 (N_23825,N_20737,N_22424);
nor U23826 (N_23826,N_20775,N_22488);
nor U23827 (N_23827,N_20852,N_21563);
nand U23828 (N_23828,N_21343,N_20426);
and U23829 (N_23829,N_20541,N_21897);
xnor U23830 (N_23830,N_20411,N_20537);
or U23831 (N_23831,N_21200,N_20546);
nor U23832 (N_23832,N_22331,N_22240);
nand U23833 (N_23833,N_21184,N_21780);
nand U23834 (N_23834,N_21320,N_22370);
or U23835 (N_23835,N_20156,N_20170);
xnor U23836 (N_23836,N_20821,N_21683);
and U23837 (N_23837,N_22105,N_20409);
xnor U23838 (N_23838,N_21462,N_22148);
or U23839 (N_23839,N_22474,N_20311);
and U23840 (N_23840,N_22380,N_22434);
nor U23841 (N_23841,N_20795,N_21559);
or U23842 (N_23842,N_21318,N_20334);
nor U23843 (N_23843,N_21013,N_20439);
nor U23844 (N_23844,N_21275,N_20319);
or U23845 (N_23845,N_21983,N_20329);
or U23846 (N_23846,N_22369,N_20988);
nor U23847 (N_23847,N_20725,N_20475);
or U23848 (N_23848,N_21367,N_20899);
xor U23849 (N_23849,N_21034,N_21783);
nor U23850 (N_23850,N_22350,N_21478);
nand U23851 (N_23851,N_21870,N_20754);
nor U23852 (N_23852,N_20616,N_20322);
or U23853 (N_23853,N_20140,N_22178);
nand U23854 (N_23854,N_22430,N_21674);
and U23855 (N_23855,N_20414,N_21473);
nand U23856 (N_23856,N_20657,N_21026);
nand U23857 (N_23857,N_21642,N_21925);
nand U23858 (N_23858,N_21990,N_20733);
nor U23859 (N_23859,N_21186,N_21391);
nand U23860 (N_23860,N_21119,N_21934);
or U23861 (N_23861,N_21885,N_20369);
or U23862 (N_23862,N_21446,N_21138);
or U23863 (N_23863,N_20154,N_21065);
or U23864 (N_23864,N_20207,N_21102);
nor U23865 (N_23865,N_21349,N_21649);
xor U23866 (N_23866,N_21211,N_22461);
and U23867 (N_23867,N_21255,N_21498);
nor U23868 (N_23868,N_21775,N_20285);
nor U23869 (N_23869,N_21117,N_21899);
nand U23870 (N_23870,N_20673,N_22010);
nor U23871 (N_23871,N_21029,N_22193);
or U23872 (N_23872,N_20811,N_20460);
or U23873 (N_23873,N_22000,N_20277);
nand U23874 (N_23874,N_20334,N_20264);
nand U23875 (N_23875,N_21211,N_21173);
nor U23876 (N_23876,N_22145,N_20800);
nand U23877 (N_23877,N_22153,N_21889);
nand U23878 (N_23878,N_22428,N_22277);
or U23879 (N_23879,N_21745,N_20125);
nor U23880 (N_23880,N_21842,N_21000);
nand U23881 (N_23881,N_22375,N_20044);
xor U23882 (N_23882,N_21218,N_22259);
nand U23883 (N_23883,N_21128,N_21055);
nor U23884 (N_23884,N_20141,N_21974);
or U23885 (N_23885,N_21209,N_22384);
or U23886 (N_23886,N_20848,N_22332);
and U23887 (N_23887,N_22012,N_21864);
and U23888 (N_23888,N_21388,N_21936);
and U23889 (N_23889,N_20566,N_20363);
xnor U23890 (N_23890,N_22116,N_20642);
and U23891 (N_23891,N_22447,N_21096);
or U23892 (N_23892,N_22221,N_20641);
xor U23893 (N_23893,N_22238,N_21582);
or U23894 (N_23894,N_21309,N_21488);
xor U23895 (N_23895,N_21297,N_21430);
or U23896 (N_23896,N_20659,N_21420);
nand U23897 (N_23897,N_20237,N_21096);
xnor U23898 (N_23898,N_21407,N_20363);
and U23899 (N_23899,N_21075,N_20049);
nor U23900 (N_23900,N_21321,N_21580);
nand U23901 (N_23901,N_21389,N_20553);
nand U23902 (N_23902,N_21032,N_20083);
nor U23903 (N_23903,N_21951,N_20996);
nand U23904 (N_23904,N_21528,N_20458);
nand U23905 (N_23905,N_22176,N_20130);
or U23906 (N_23906,N_20419,N_20443);
and U23907 (N_23907,N_22497,N_20952);
xor U23908 (N_23908,N_21291,N_22294);
and U23909 (N_23909,N_21147,N_20193);
or U23910 (N_23910,N_20796,N_22049);
or U23911 (N_23911,N_22102,N_21719);
or U23912 (N_23912,N_22349,N_21346);
and U23913 (N_23913,N_21495,N_22052);
and U23914 (N_23914,N_22206,N_21894);
nor U23915 (N_23915,N_20684,N_21372);
and U23916 (N_23916,N_21327,N_21002);
or U23917 (N_23917,N_22335,N_20212);
nand U23918 (N_23918,N_20774,N_21811);
nor U23919 (N_23919,N_20979,N_20384);
and U23920 (N_23920,N_20306,N_22302);
and U23921 (N_23921,N_20257,N_20905);
and U23922 (N_23922,N_20576,N_20001);
and U23923 (N_23923,N_22220,N_21317);
nand U23924 (N_23924,N_21899,N_21509);
or U23925 (N_23925,N_21262,N_20257);
or U23926 (N_23926,N_20582,N_20342);
nor U23927 (N_23927,N_21718,N_20184);
and U23928 (N_23928,N_22385,N_20373);
or U23929 (N_23929,N_22346,N_20970);
or U23930 (N_23930,N_20686,N_20878);
or U23931 (N_23931,N_22332,N_20032);
nor U23932 (N_23932,N_20168,N_21002);
nor U23933 (N_23933,N_21204,N_20464);
or U23934 (N_23934,N_21559,N_20445);
nor U23935 (N_23935,N_21734,N_22021);
or U23936 (N_23936,N_20073,N_21544);
xnor U23937 (N_23937,N_22024,N_20221);
xor U23938 (N_23938,N_22479,N_21881);
nor U23939 (N_23939,N_21597,N_20941);
and U23940 (N_23940,N_20405,N_21924);
nor U23941 (N_23941,N_21543,N_20632);
nor U23942 (N_23942,N_20997,N_21960);
and U23943 (N_23943,N_20895,N_20478);
nor U23944 (N_23944,N_20867,N_22319);
nand U23945 (N_23945,N_21348,N_21835);
or U23946 (N_23946,N_21691,N_21876);
nor U23947 (N_23947,N_20199,N_22357);
nor U23948 (N_23948,N_21466,N_21709);
nand U23949 (N_23949,N_20916,N_22453);
or U23950 (N_23950,N_20633,N_20783);
and U23951 (N_23951,N_21954,N_20724);
nor U23952 (N_23952,N_22420,N_20441);
or U23953 (N_23953,N_21333,N_21000);
nand U23954 (N_23954,N_21457,N_20986);
nand U23955 (N_23955,N_20074,N_20124);
or U23956 (N_23956,N_22080,N_22217);
nor U23957 (N_23957,N_21280,N_22248);
or U23958 (N_23958,N_22466,N_20191);
nand U23959 (N_23959,N_20496,N_20853);
or U23960 (N_23960,N_20872,N_20432);
nand U23961 (N_23961,N_21538,N_22066);
and U23962 (N_23962,N_20094,N_22224);
or U23963 (N_23963,N_21561,N_22240);
or U23964 (N_23964,N_20584,N_20271);
nor U23965 (N_23965,N_22130,N_20631);
nor U23966 (N_23966,N_20440,N_21483);
nand U23967 (N_23967,N_21699,N_21702);
nor U23968 (N_23968,N_20871,N_21776);
xnor U23969 (N_23969,N_21222,N_20184);
xor U23970 (N_23970,N_22014,N_21826);
nand U23971 (N_23971,N_20376,N_20168);
or U23972 (N_23972,N_21581,N_20719);
xor U23973 (N_23973,N_20780,N_22044);
nand U23974 (N_23974,N_20381,N_22274);
or U23975 (N_23975,N_22143,N_22086);
nand U23976 (N_23976,N_21725,N_22163);
or U23977 (N_23977,N_20452,N_21106);
xnor U23978 (N_23978,N_20305,N_21706);
nor U23979 (N_23979,N_20551,N_21143);
or U23980 (N_23980,N_20821,N_20718);
xor U23981 (N_23981,N_20710,N_20800);
and U23982 (N_23982,N_20645,N_20715);
nand U23983 (N_23983,N_21434,N_22409);
xnor U23984 (N_23984,N_22066,N_20062);
nor U23985 (N_23985,N_22140,N_21821);
or U23986 (N_23986,N_22321,N_20772);
or U23987 (N_23987,N_20375,N_21914);
nor U23988 (N_23988,N_21465,N_20875);
nand U23989 (N_23989,N_20601,N_21239);
nor U23990 (N_23990,N_20618,N_20654);
nor U23991 (N_23991,N_20864,N_20920);
nor U23992 (N_23992,N_21109,N_21479);
nor U23993 (N_23993,N_21598,N_20267);
and U23994 (N_23994,N_21069,N_22231);
nand U23995 (N_23995,N_22470,N_21783);
nand U23996 (N_23996,N_22421,N_21080);
and U23997 (N_23997,N_21022,N_22137);
nor U23998 (N_23998,N_20185,N_21028);
nor U23999 (N_23999,N_21296,N_21200);
nand U24000 (N_24000,N_22276,N_20315);
nand U24001 (N_24001,N_20672,N_21620);
nand U24002 (N_24002,N_22129,N_20163);
and U24003 (N_24003,N_20687,N_22013);
and U24004 (N_24004,N_21659,N_20557);
or U24005 (N_24005,N_22270,N_21337);
or U24006 (N_24006,N_22220,N_20853);
nand U24007 (N_24007,N_22174,N_22382);
and U24008 (N_24008,N_20352,N_21117);
nand U24009 (N_24009,N_21025,N_20950);
nor U24010 (N_24010,N_21708,N_20106);
xnor U24011 (N_24011,N_21147,N_22447);
nand U24012 (N_24012,N_21990,N_21027);
xor U24013 (N_24013,N_21582,N_20993);
nand U24014 (N_24014,N_21376,N_21503);
nand U24015 (N_24015,N_20564,N_21199);
nor U24016 (N_24016,N_20612,N_21331);
or U24017 (N_24017,N_20532,N_21438);
and U24018 (N_24018,N_21018,N_22371);
and U24019 (N_24019,N_20062,N_21764);
or U24020 (N_24020,N_20791,N_20048);
nand U24021 (N_24021,N_21688,N_20387);
nor U24022 (N_24022,N_21478,N_21382);
nor U24023 (N_24023,N_20732,N_21623);
nand U24024 (N_24024,N_21011,N_21095);
nor U24025 (N_24025,N_21923,N_21245);
or U24026 (N_24026,N_21443,N_20511);
and U24027 (N_24027,N_20542,N_21482);
nand U24028 (N_24028,N_20073,N_20263);
and U24029 (N_24029,N_21965,N_21410);
or U24030 (N_24030,N_22492,N_21248);
and U24031 (N_24031,N_21724,N_21798);
nand U24032 (N_24032,N_21059,N_21982);
xnor U24033 (N_24033,N_21343,N_22073);
nand U24034 (N_24034,N_22427,N_20064);
or U24035 (N_24035,N_20687,N_20917);
or U24036 (N_24036,N_20810,N_21678);
or U24037 (N_24037,N_22256,N_20056);
nand U24038 (N_24038,N_22351,N_21316);
xnor U24039 (N_24039,N_22339,N_22420);
or U24040 (N_24040,N_21522,N_20271);
nor U24041 (N_24041,N_20773,N_20788);
and U24042 (N_24042,N_21841,N_20129);
nand U24043 (N_24043,N_20914,N_22344);
and U24044 (N_24044,N_20145,N_21228);
nor U24045 (N_24045,N_22037,N_21892);
nor U24046 (N_24046,N_20485,N_22005);
and U24047 (N_24047,N_20220,N_21508);
and U24048 (N_24048,N_20686,N_20776);
and U24049 (N_24049,N_21578,N_20061);
and U24050 (N_24050,N_21341,N_20334);
and U24051 (N_24051,N_20506,N_20143);
nand U24052 (N_24052,N_20519,N_21431);
and U24053 (N_24053,N_21304,N_20390);
and U24054 (N_24054,N_22016,N_21261);
nor U24055 (N_24055,N_22310,N_21619);
and U24056 (N_24056,N_22012,N_21769);
or U24057 (N_24057,N_22347,N_20826);
nor U24058 (N_24058,N_21593,N_20663);
and U24059 (N_24059,N_22314,N_20388);
or U24060 (N_24060,N_20583,N_20464);
nor U24061 (N_24061,N_21517,N_21669);
or U24062 (N_24062,N_21492,N_20573);
nor U24063 (N_24063,N_21843,N_20832);
and U24064 (N_24064,N_21056,N_22150);
or U24065 (N_24065,N_20670,N_20616);
or U24066 (N_24066,N_22479,N_20758);
nand U24067 (N_24067,N_21780,N_20678);
nand U24068 (N_24068,N_22451,N_20214);
nor U24069 (N_24069,N_21471,N_20580);
nor U24070 (N_24070,N_21481,N_22097);
nor U24071 (N_24071,N_21451,N_20762);
and U24072 (N_24072,N_22004,N_22080);
nor U24073 (N_24073,N_20482,N_20626);
nor U24074 (N_24074,N_21894,N_20170);
nor U24075 (N_24075,N_21559,N_22409);
nand U24076 (N_24076,N_21421,N_20535);
nand U24077 (N_24077,N_21033,N_21535);
nor U24078 (N_24078,N_21642,N_21961);
nand U24079 (N_24079,N_21362,N_20616);
and U24080 (N_24080,N_22019,N_20935);
and U24081 (N_24081,N_21828,N_20187);
and U24082 (N_24082,N_20693,N_21371);
and U24083 (N_24083,N_21104,N_21261);
nand U24084 (N_24084,N_22285,N_21206);
and U24085 (N_24085,N_21286,N_21134);
nand U24086 (N_24086,N_21296,N_21842);
nand U24087 (N_24087,N_20861,N_22140);
nor U24088 (N_24088,N_20532,N_21380);
nor U24089 (N_24089,N_21525,N_20985);
xor U24090 (N_24090,N_20137,N_21228);
nand U24091 (N_24091,N_21993,N_22257);
and U24092 (N_24092,N_21033,N_21272);
nor U24093 (N_24093,N_22140,N_20543);
nand U24094 (N_24094,N_21379,N_21178);
nand U24095 (N_24095,N_22091,N_21908);
nand U24096 (N_24096,N_20495,N_21689);
and U24097 (N_24097,N_20184,N_22268);
and U24098 (N_24098,N_20226,N_21849);
or U24099 (N_24099,N_21425,N_20878);
xor U24100 (N_24100,N_21118,N_21946);
nand U24101 (N_24101,N_22014,N_20962);
xnor U24102 (N_24102,N_21878,N_21716);
or U24103 (N_24103,N_21978,N_21640);
and U24104 (N_24104,N_21520,N_22226);
xnor U24105 (N_24105,N_20993,N_20530);
nand U24106 (N_24106,N_20604,N_22305);
xnor U24107 (N_24107,N_20594,N_21758);
and U24108 (N_24108,N_20437,N_22200);
xnor U24109 (N_24109,N_20146,N_22070);
or U24110 (N_24110,N_20495,N_22358);
nor U24111 (N_24111,N_20710,N_22115);
nand U24112 (N_24112,N_22034,N_21071);
and U24113 (N_24113,N_21720,N_20777);
and U24114 (N_24114,N_20957,N_20831);
nor U24115 (N_24115,N_21609,N_21787);
nand U24116 (N_24116,N_21587,N_21565);
nor U24117 (N_24117,N_20252,N_20057);
or U24118 (N_24118,N_21067,N_20840);
or U24119 (N_24119,N_22203,N_20896);
nand U24120 (N_24120,N_20498,N_22135);
and U24121 (N_24121,N_20500,N_22061);
and U24122 (N_24122,N_20894,N_20749);
or U24123 (N_24123,N_21214,N_22102);
nand U24124 (N_24124,N_21760,N_20452);
nand U24125 (N_24125,N_21666,N_20483);
nor U24126 (N_24126,N_22162,N_20144);
nand U24127 (N_24127,N_20323,N_21816);
or U24128 (N_24128,N_21910,N_22090);
nand U24129 (N_24129,N_22158,N_20812);
nand U24130 (N_24130,N_22116,N_21828);
nor U24131 (N_24131,N_20602,N_21239);
nand U24132 (N_24132,N_21000,N_20698);
and U24133 (N_24133,N_20292,N_21523);
or U24134 (N_24134,N_21134,N_20016);
nand U24135 (N_24135,N_20978,N_20900);
or U24136 (N_24136,N_22174,N_20324);
nor U24137 (N_24137,N_20031,N_22442);
and U24138 (N_24138,N_22363,N_21037);
or U24139 (N_24139,N_21873,N_20314);
nor U24140 (N_24140,N_22025,N_20677);
nand U24141 (N_24141,N_21304,N_20582);
nor U24142 (N_24142,N_20437,N_22275);
or U24143 (N_24143,N_22277,N_21712);
nor U24144 (N_24144,N_20410,N_22374);
and U24145 (N_24145,N_20051,N_20764);
and U24146 (N_24146,N_20157,N_22377);
nor U24147 (N_24147,N_21415,N_20545);
and U24148 (N_24148,N_21234,N_20080);
and U24149 (N_24149,N_21641,N_22096);
xnor U24150 (N_24150,N_22436,N_21980);
and U24151 (N_24151,N_21210,N_21094);
and U24152 (N_24152,N_22173,N_20348);
nor U24153 (N_24153,N_22216,N_21176);
nand U24154 (N_24154,N_20381,N_21166);
and U24155 (N_24155,N_20032,N_20966);
or U24156 (N_24156,N_20267,N_22151);
and U24157 (N_24157,N_21449,N_21030);
nor U24158 (N_24158,N_20469,N_21586);
or U24159 (N_24159,N_20277,N_21352);
xnor U24160 (N_24160,N_21354,N_22253);
nand U24161 (N_24161,N_21844,N_21964);
or U24162 (N_24162,N_21422,N_22261);
or U24163 (N_24163,N_21785,N_20507);
and U24164 (N_24164,N_21066,N_20691);
and U24165 (N_24165,N_22221,N_20978);
nand U24166 (N_24166,N_20327,N_20691);
and U24167 (N_24167,N_21219,N_22150);
or U24168 (N_24168,N_21390,N_20096);
nand U24169 (N_24169,N_21213,N_20672);
nor U24170 (N_24170,N_20609,N_20009);
or U24171 (N_24171,N_21268,N_22458);
nor U24172 (N_24172,N_21220,N_21084);
and U24173 (N_24173,N_20141,N_20130);
xor U24174 (N_24174,N_20354,N_21873);
or U24175 (N_24175,N_21655,N_22467);
xor U24176 (N_24176,N_20443,N_20923);
nand U24177 (N_24177,N_22314,N_21596);
or U24178 (N_24178,N_20048,N_21557);
and U24179 (N_24179,N_21697,N_21827);
nor U24180 (N_24180,N_22440,N_20579);
xor U24181 (N_24181,N_20317,N_20453);
or U24182 (N_24182,N_22069,N_21676);
or U24183 (N_24183,N_21616,N_20022);
nor U24184 (N_24184,N_21807,N_21368);
nor U24185 (N_24185,N_20698,N_21108);
nand U24186 (N_24186,N_20886,N_21027);
nand U24187 (N_24187,N_21030,N_20466);
nand U24188 (N_24188,N_22008,N_20468);
or U24189 (N_24189,N_21707,N_22088);
and U24190 (N_24190,N_21960,N_21939);
and U24191 (N_24191,N_20902,N_21099);
nor U24192 (N_24192,N_22296,N_20450);
nor U24193 (N_24193,N_20373,N_20559);
nor U24194 (N_24194,N_21040,N_20279);
and U24195 (N_24195,N_21594,N_22498);
and U24196 (N_24196,N_21107,N_22393);
and U24197 (N_24197,N_20609,N_20994);
and U24198 (N_24198,N_21355,N_21346);
and U24199 (N_24199,N_21735,N_20188);
and U24200 (N_24200,N_20834,N_22186);
or U24201 (N_24201,N_22318,N_21186);
nand U24202 (N_24202,N_21097,N_21758);
or U24203 (N_24203,N_22467,N_21705);
nor U24204 (N_24204,N_20617,N_22433);
nand U24205 (N_24205,N_22127,N_22326);
nand U24206 (N_24206,N_20715,N_21153);
or U24207 (N_24207,N_21280,N_21253);
nand U24208 (N_24208,N_21777,N_22244);
nor U24209 (N_24209,N_22097,N_20390);
xor U24210 (N_24210,N_21310,N_21753);
xnor U24211 (N_24211,N_22317,N_20226);
and U24212 (N_24212,N_20424,N_22261);
and U24213 (N_24213,N_21249,N_21801);
nor U24214 (N_24214,N_22232,N_20715);
and U24215 (N_24215,N_20013,N_20345);
or U24216 (N_24216,N_21837,N_21015);
xnor U24217 (N_24217,N_21152,N_20447);
or U24218 (N_24218,N_21166,N_21119);
and U24219 (N_24219,N_22495,N_22100);
and U24220 (N_24220,N_21698,N_22428);
nand U24221 (N_24221,N_22446,N_20603);
nand U24222 (N_24222,N_22032,N_21533);
nor U24223 (N_24223,N_21561,N_21925);
xnor U24224 (N_24224,N_20849,N_20706);
nand U24225 (N_24225,N_21069,N_20201);
and U24226 (N_24226,N_21000,N_20431);
xnor U24227 (N_24227,N_21533,N_21869);
nor U24228 (N_24228,N_20291,N_20331);
or U24229 (N_24229,N_22317,N_20345);
nand U24230 (N_24230,N_20644,N_21741);
nor U24231 (N_24231,N_21431,N_20154);
xor U24232 (N_24232,N_21406,N_22452);
nand U24233 (N_24233,N_22078,N_21837);
and U24234 (N_24234,N_21412,N_21621);
xnor U24235 (N_24235,N_21370,N_20025);
nor U24236 (N_24236,N_20556,N_22399);
or U24237 (N_24237,N_20525,N_21453);
xnor U24238 (N_24238,N_22392,N_20039);
xor U24239 (N_24239,N_21471,N_22439);
and U24240 (N_24240,N_21053,N_21287);
nor U24241 (N_24241,N_20414,N_20056);
and U24242 (N_24242,N_21128,N_21513);
or U24243 (N_24243,N_20101,N_20887);
nand U24244 (N_24244,N_20952,N_21454);
nand U24245 (N_24245,N_22264,N_20392);
xnor U24246 (N_24246,N_21228,N_21341);
and U24247 (N_24247,N_20270,N_20668);
xor U24248 (N_24248,N_20266,N_21736);
nor U24249 (N_24249,N_21712,N_20524);
nand U24250 (N_24250,N_20258,N_21053);
and U24251 (N_24251,N_20586,N_20476);
nor U24252 (N_24252,N_20982,N_20101);
nand U24253 (N_24253,N_21482,N_20648);
xor U24254 (N_24254,N_21708,N_22400);
and U24255 (N_24255,N_21750,N_20004);
xnor U24256 (N_24256,N_21340,N_20522);
nand U24257 (N_24257,N_20473,N_20705);
or U24258 (N_24258,N_21900,N_20493);
nand U24259 (N_24259,N_21040,N_21873);
nand U24260 (N_24260,N_22051,N_21200);
nand U24261 (N_24261,N_20191,N_22087);
or U24262 (N_24262,N_21422,N_21928);
nor U24263 (N_24263,N_21455,N_22317);
nand U24264 (N_24264,N_20414,N_20432);
nor U24265 (N_24265,N_21532,N_22236);
nor U24266 (N_24266,N_21268,N_20471);
or U24267 (N_24267,N_22301,N_20778);
xnor U24268 (N_24268,N_20565,N_21029);
or U24269 (N_24269,N_22359,N_22363);
or U24270 (N_24270,N_21202,N_20214);
or U24271 (N_24271,N_20196,N_20667);
nand U24272 (N_24272,N_21571,N_20493);
and U24273 (N_24273,N_20235,N_20918);
nor U24274 (N_24274,N_21283,N_20334);
nand U24275 (N_24275,N_22418,N_21433);
or U24276 (N_24276,N_20990,N_21836);
nor U24277 (N_24277,N_21584,N_20235);
nor U24278 (N_24278,N_21707,N_20637);
nor U24279 (N_24279,N_22146,N_20480);
nor U24280 (N_24280,N_20850,N_20759);
and U24281 (N_24281,N_20563,N_21899);
or U24282 (N_24282,N_22154,N_22438);
and U24283 (N_24283,N_20541,N_21295);
or U24284 (N_24284,N_21338,N_21500);
xnor U24285 (N_24285,N_20987,N_21181);
or U24286 (N_24286,N_21251,N_21565);
xnor U24287 (N_24287,N_21025,N_21123);
or U24288 (N_24288,N_20327,N_20504);
or U24289 (N_24289,N_21031,N_22194);
nand U24290 (N_24290,N_20761,N_20268);
or U24291 (N_24291,N_20015,N_21249);
nor U24292 (N_24292,N_21666,N_22405);
nand U24293 (N_24293,N_21538,N_20838);
nand U24294 (N_24294,N_20804,N_21267);
and U24295 (N_24295,N_21851,N_21746);
xnor U24296 (N_24296,N_20419,N_21272);
xnor U24297 (N_24297,N_21777,N_20675);
nor U24298 (N_24298,N_22164,N_21426);
and U24299 (N_24299,N_20734,N_20762);
nand U24300 (N_24300,N_20004,N_21489);
or U24301 (N_24301,N_20425,N_22372);
xor U24302 (N_24302,N_21909,N_20845);
and U24303 (N_24303,N_21411,N_20970);
and U24304 (N_24304,N_22039,N_22160);
nor U24305 (N_24305,N_22477,N_21131);
nor U24306 (N_24306,N_21977,N_21473);
nor U24307 (N_24307,N_21157,N_20637);
or U24308 (N_24308,N_21692,N_20827);
nand U24309 (N_24309,N_20199,N_20772);
nor U24310 (N_24310,N_21009,N_21031);
xnor U24311 (N_24311,N_22382,N_21387);
nor U24312 (N_24312,N_21936,N_22191);
xor U24313 (N_24313,N_20046,N_21234);
and U24314 (N_24314,N_22451,N_21692);
xnor U24315 (N_24315,N_20625,N_20268);
nand U24316 (N_24316,N_21486,N_21498);
or U24317 (N_24317,N_21469,N_21352);
or U24318 (N_24318,N_20381,N_22445);
nor U24319 (N_24319,N_20403,N_20846);
nand U24320 (N_24320,N_20822,N_22095);
or U24321 (N_24321,N_20236,N_20972);
nor U24322 (N_24322,N_20674,N_22270);
or U24323 (N_24323,N_20551,N_21859);
nand U24324 (N_24324,N_21750,N_20773);
or U24325 (N_24325,N_21709,N_22263);
and U24326 (N_24326,N_20964,N_22480);
nor U24327 (N_24327,N_21896,N_21732);
or U24328 (N_24328,N_20687,N_22199);
and U24329 (N_24329,N_22231,N_20180);
nand U24330 (N_24330,N_20526,N_21138);
and U24331 (N_24331,N_21399,N_20896);
xnor U24332 (N_24332,N_21889,N_21932);
or U24333 (N_24333,N_22315,N_20392);
nand U24334 (N_24334,N_20645,N_20854);
xor U24335 (N_24335,N_21616,N_21449);
or U24336 (N_24336,N_21634,N_20372);
and U24337 (N_24337,N_20180,N_20574);
nand U24338 (N_24338,N_22440,N_21487);
or U24339 (N_24339,N_20119,N_20885);
and U24340 (N_24340,N_20602,N_22282);
nor U24341 (N_24341,N_20499,N_20772);
and U24342 (N_24342,N_21948,N_21999);
nand U24343 (N_24343,N_20009,N_21911);
or U24344 (N_24344,N_21415,N_20011);
and U24345 (N_24345,N_21215,N_20103);
nor U24346 (N_24346,N_20647,N_22316);
nor U24347 (N_24347,N_22246,N_21647);
and U24348 (N_24348,N_22464,N_20404);
or U24349 (N_24349,N_22249,N_20479);
or U24350 (N_24350,N_20233,N_20850);
nor U24351 (N_24351,N_21524,N_21427);
nand U24352 (N_24352,N_22311,N_20689);
or U24353 (N_24353,N_22109,N_21348);
xor U24354 (N_24354,N_21502,N_20700);
nand U24355 (N_24355,N_21515,N_20954);
nand U24356 (N_24356,N_21876,N_21620);
xor U24357 (N_24357,N_22187,N_20764);
and U24358 (N_24358,N_21254,N_20666);
nor U24359 (N_24359,N_21358,N_20673);
and U24360 (N_24360,N_22311,N_21803);
nand U24361 (N_24361,N_20571,N_20351);
or U24362 (N_24362,N_22223,N_22185);
xor U24363 (N_24363,N_20316,N_20011);
or U24364 (N_24364,N_22495,N_21148);
nand U24365 (N_24365,N_20286,N_21052);
and U24366 (N_24366,N_22224,N_21794);
xor U24367 (N_24367,N_21161,N_20887);
nor U24368 (N_24368,N_21731,N_20567);
or U24369 (N_24369,N_21237,N_20245);
nand U24370 (N_24370,N_21400,N_20936);
nand U24371 (N_24371,N_20593,N_21343);
nand U24372 (N_24372,N_21030,N_21052);
nor U24373 (N_24373,N_21517,N_21435);
or U24374 (N_24374,N_22461,N_21515);
xnor U24375 (N_24375,N_22169,N_21073);
nor U24376 (N_24376,N_21493,N_21431);
or U24377 (N_24377,N_21736,N_20170);
nor U24378 (N_24378,N_20300,N_20230);
nor U24379 (N_24379,N_20723,N_20824);
nand U24380 (N_24380,N_21295,N_20982);
nand U24381 (N_24381,N_21699,N_21416);
nor U24382 (N_24382,N_22052,N_21829);
nand U24383 (N_24383,N_20339,N_21598);
nor U24384 (N_24384,N_20132,N_21453);
xor U24385 (N_24385,N_20914,N_22394);
xnor U24386 (N_24386,N_21646,N_20823);
and U24387 (N_24387,N_21234,N_20217);
nor U24388 (N_24388,N_20484,N_22285);
nor U24389 (N_24389,N_22207,N_21687);
nand U24390 (N_24390,N_22117,N_21154);
nor U24391 (N_24391,N_20402,N_21009);
and U24392 (N_24392,N_20187,N_22142);
xnor U24393 (N_24393,N_20434,N_20864);
or U24394 (N_24394,N_21108,N_20192);
and U24395 (N_24395,N_21415,N_21813);
nor U24396 (N_24396,N_22030,N_20256);
and U24397 (N_24397,N_21799,N_20120);
or U24398 (N_24398,N_20973,N_22271);
nand U24399 (N_24399,N_22138,N_22340);
xnor U24400 (N_24400,N_21129,N_20021);
nand U24401 (N_24401,N_20706,N_20000);
nor U24402 (N_24402,N_21039,N_20845);
and U24403 (N_24403,N_22345,N_22097);
nand U24404 (N_24404,N_20948,N_22313);
nor U24405 (N_24405,N_22204,N_20703);
xnor U24406 (N_24406,N_21459,N_22042);
nor U24407 (N_24407,N_22247,N_20560);
nor U24408 (N_24408,N_20798,N_21628);
xor U24409 (N_24409,N_21889,N_21840);
nand U24410 (N_24410,N_21807,N_20970);
nand U24411 (N_24411,N_21474,N_20419);
nand U24412 (N_24412,N_21590,N_20068);
or U24413 (N_24413,N_20619,N_20386);
xor U24414 (N_24414,N_20321,N_21948);
or U24415 (N_24415,N_20654,N_20949);
or U24416 (N_24416,N_21408,N_20716);
nor U24417 (N_24417,N_21170,N_20689);
and U24418 (N_24418,N_21194,N_21999);
or U24419 (N_24419,N_21894,N_21071);
and U24420 (N_24420,N_20194,N_21892);
nand U24421 (N_24421,N_21036,N_21489);
xor U24422 (N_24422,N_21728,N_22064);
nor U24423 (N_24423,N_20897,N_20220);
or U24424 (N_24424,N_20093,N_21718);
and U24425 (N_24425,N_21960,N_20606);
nand U24426 (N_24426,N_20980,N_21982);
nand U24427 (N_24427,N_20347,N_22211);
nand U24428 (N_24428,N_20769,N_21329);
or U24429 (N_24429,N_21159,N_21243);
or U24430 (N_24430,N_20230,N_21043);
xor U24431 (N_24431,N_21048,N_21479);
or U24432 (N_24432,N_21568,N_20762);
or U24433 (N_24433,N_21396,N_20125);
or U24434 (N_24434,N_22020,N_22379);
or U24435 (N_24435,N_20545,N_20690);
nand U24436 (N_24436,N_21866,N_22409);
nor U24437 (N_24437,N_20559,N_20003);
nand U24438 (N_24438,N_21407,N_20074);
nor U24439 (N_24439,N_21120,N_22059);
nand U24440 (N_24440,N_20618,N_22070);
nor U24441 (N_24441,N_21723,N_21167);
xnor U24442 (N_24442,N_22048,N_22487);
nand U24443 (N_24443,N_20725,N_20573);
nand U24444 (N_24444,N_20474,N_21415);
nand U24445 (N_24445,N_21297,N_20641);
nand U24446 (N_24446,N_22290,N_22468);
and U24447 (N_24447,N_21061,N_20879);
nand U24448 (N_24448,N_21076,N_20497);
nor U24449 (N_24449,N_21692,N_20349);
xor U24450 (N_24450,N_20422,N_22372);
nand U24451 (N_24451,N_22062,N_22149);
or U24452 (N_24452,N_20527,N_21189);
nand U24453 (N_24453,N_21790,N_20473);
and U24454 (N_24454,N_21532,N_20837);
nand U24455 (N_24455,N_22019,N_22094);
or U24456 (N_24456,N_20148,N_20725);
or U24457 (N_24457,N_22137,N_21762);
nor U24458 (N_24458,N_20168,N_21347);
nor U24459 (N_24459,N_21348,N_21579);
and U24460 (N_24460,N_21262,N_22409);
or U24461 (N_24461,N_21804,N_21392);
or U24462 (N_24462,N_20445,N_22034);
nand U24463 (N_24463,N_20292,N_20601);
or U24464 (N_24464,N_21657,N_20214);
nor U24465 (N_24465,N_20733,N_20402);
nand U24466 (N_24466,N_22085,N_20493);
xor U24467 (N_24467,N_22251,N_20236);
nor U24468 (N_24468,N_20307,N_22465);
xnor U24469 (N_24469,N_21145,N_21845);
and U24470 (N_24470,N_22216,N_21251);
and U24471 (N_24471,N_21626,N_21551);
xnor U24472 (N_24472,N_20548,N_22005);
nor U24473 (N_24473,N_21253,N_22369);
nor U24474 (N_24474,N_21642,N_21621);
nand U24475 (N_24475,N_21022,N_21600);
and U24476 (N_24476,N_22112,N_21784);
nand U24477 (N_24477,N_20670,N_20149);
nand U24478 (N_24478,N_20352,N_21866);
or U24479 (N_24479,N_22356,N_21522);
nor U24480 (N_24480,N_22122,N_21237);
nor U24481 (N_24481,N_21615,N_21819);
and U24482 (N_24482,N_22458,N_22050);
xor U24483 (N_24483,N_20798,N_21372);
or U24484 (N_24484,N_22476,N_20173);
or U24485 (N_24485,N_21277,N_21549);
and U24486 (N_24486,N_21633,N_21837);
or U24487 (N_24487,N_20907,N_21596);
nor U24488 (N_24488,N_21070,N_20986);
nand U24489 (N_24489,N_21654,N_22073);
and U24490 (N_24490,N_21300,N_20159);
nand U24491 (N_24491,N_21797,N_20804);
and U24492 (N_24492,N_20087,N_21332);
nor U24493 (N_24493,N_22452,N_20968);
nor U24494 (N_24494,N_22377,N_21282);
nor U24495 (N_24495,N_21557,N_20520);
or U24496 (N_24496,N_22320,N_20283);
nand U24497 (N_24497,N_21553,N_21693);
nand U24498 (N_24498,N_22242,N_20183);
nor U24499 (N_24499,N_20077,N_20736);
or U24500 (N_24500,N_21051,N_20083);
nand U24501 (N_24501,N_22369,N_22461);
and U24502 (N_24502,N_20233,N_20200);
nor U24503 (N_24503,N_21940,N_20696);
nor U24504 (N_24504,N_22456,N_22060);
nand U24505 (N_24505,N_20496,N_20271);
nor U24506 (N_24506,N_21402,N_21377);
and U24507 (N_24507,N_21970,N_21744);
nand U24508 (N_24508,N_20295,N_21636);
or U24509 (N_24509,N_21499,N_20737);
nand U24510 (N_24510,N_20842,N_20076);
nand U24511 (N_24511,N_21433,N_22053);
nor U24512 (N_24512,N_20463,N_20457);
xor U24513 (N_24513,N_20142,N_21566);
xnor U24514 (N_24514,N_20785,N_21087);
and U24515 (N_24515,N_20541,N_20851);
nand U24516 (N_24516,N_22075,N_22030);
nand U24517 (N_24517,N_20147,N_21262);
or U24518 (N_24518,N_21041,N_20547);
nor U24519 (N_24519,N_21638,N_21255);
and U24520 (N_24520,N_20088,N_21011);
or U24521 (N_24521,N_20642,N_20393);
and U24522 (N_24522,N_20180,N_21542);
nor U24523 (N_24523,N_20340,N_20658);
nand U24524 (N_24524,N_22334,N_21796);
and U24525 (N_24525,N_21439,N_20913);
xnor U24526 (N_24526,N_21375,N_20838);
or U24527 (N_24527,N_20919,N_21310);
xor U24528 (N_24528,N_21211,N_20005);
nor U24529 (N_24529,N_20440,N_22430);
nor U24530 (N_24530,N_20150,N_22228);
nor U24531 (N_24531,N_21653,N_20748);
or U24532 (N_24532,N_20640,N_20676);
nor U24533 (N_24533,N_21795,N_20798);
nand U24534 (N_24534,N_22458,N_20434);
xor U24535 (N_24535,N_21775,N_22223);
and U24536 (N_24536,N_21837,N_21256);
nor U24537 (N_24537,N_21814,N_21388);
or U24538 (N_24538,N_20359,N_20885);
nor U24539 (N_24539,N_20535,N_20856);
nor U24540 (N_24540,N_21869,N_20504);
nand U24541 (N_24541,N_22479,N_21896);
and U24542 (N_24542,N_22171,N_20833);
and U24543 (N_24543,N_20100,N_21658);
nand U24544 (N_24544,N_22079,N_21157);
xnor U24545 (N_24545,N_21437,N_20628);
and U24546 (N_24546,N_20339,N_20706);
nor U24547 (N_24547,N_21873,N_20700);
and U24548 (N_24548,N_20375,N_22450);
nor U24549 (N_24549,N_21940,N_20878);
xnor U24550 (N_24550,N_21617,N_22348);
xor U24551 (N_24551,N_22140,N_21141);
nor U24552 (N_24552,N_21753,N_22324);
or U24553 (N_24553,N_21957,N_21260);
and U24554 (N_24554,N_22133,N_21630);
and U24555 (N_24555,N_20892,N_20062);
and U24556 (N_24556,N_20190,N_22487);
and U24557 (N_24557,N_21774,N_20145);
nand U24558 (N_24558,N_22133,N_22033);
and U24559 (N_24559,N_21415,N_20128);
nor U24560 (N_24560,N_21318,N_21063);
or U24561 (N_24561,N_21375,N_21569);
nand U24562 (N_24562,N_21816,N_22246);
xor U24563 (N_24563,N_21758,N_22177);
nand U24564 (N_24564,N_20910,N_20863);
nand U24565 (N_24565,N_20196,N_21898);
and U24566 (N_24566,N_22292,N_20006);
nand U24567 (N_24567,N_21051,N_20704);
nor U24568 (N_24568,N_21669,N_20370);
nand U24569 (N_24569,N_20390,N_21717);
and U24570 (N_24570,N_22188,N_20075);
or U24571 (N_24571,N_21384,N_21381);
and U24572 (N_24572,N_20466,N_21439);
and U24573 (N_24573,N_21104,N_21224);
nor U24574 (N_24574,N_20986,N_21053);
nor U24575 (N_24575,N_20800,N_22111);
nor U24576 (N_24576,N_20237,N_21894);
and U24577 (N_24577,N_22406,N_21995);
and U24578 (N_24578,N_21049,N_21265);
and U24579 (N_24579,N_21951,N_22446);
nor U24580 (N_24580,N_20287,N_20166);
nand U24581 (N_24581,N_22153,N_21550);
nand U24582 (N_24582,N_21595,N_21089);
xnor U24583 (N_24583,N_21691,N_21466);
nand U24584 (N_24584,N_21520,N_22257);
or U24585 (N_24585,N_20067,N_21710);
and U24586 (N_24586,N_21709,N_20662);
or U24587 (N_24587,N_21108,N_21984);
nor U24588 (N_24588,N_20663,N_20514);
or U24589 (N_24589,N_20172,N_20407);
or U24590 (N_24590,N_22119,N_21051);
and U24591 (N_24591,N_21365,N_20339);
and U24592 (N_24592,N_22300,N_20209);
nor U24593 (N_24593,N_22479,N_21020);
and U24594 (N_24594,N_21254,N_22304);
xnor U24595 (N_24595,N_21437,N_20596);
and U24596 (N_24596,N_20767,N_21695);
and U24597 (N_24597,N_20058,N_21676);
or U24598 (N_24598,N_21297,N_20402);
xnor U24599 (N_24599,N_20414,N_21986);
nand U24600 (N_24600,N_22303,N_22041);
nand U24601 (N_24601,N_22247,N_22264);
and U24602 (N_24602,N_20821,N_20136);
nor U24603 (N_24603,N_21652,N_22138);
or U24604 (N_24604,N_20850,N_21133);
xnor U24605 (N_24605,N_21452,N_22489);
and U24606 (N_24606,N_20705,N_20079);
xor U24607 (N_24607,N_20248,N_21282);
or U24608 (N_24608,N_20325,N_20567);
nand U24609 (N_24609,N_21036,N_21577);
or U24610 (N_24610,N_22153,N_21509);
nand U24611 (N_24611,N_20877,N_20799);
or U24612 (N_24612,N_21996,N_22266);
and U24613 (N_24613,N_21480,N_21140);
or U24614 (N_24614,N_20344,N_20710);
nand U24615 (N_24615,N_20541,N_20697);
nand U24616 (N_24616,N_20595,N_20997);
and U24617 (N_24617,N_22251,N_20875);
and U24618 (N_24618,N_21483,N_21639);
nand U24619 (N_24619,N_21382,N_20782);
or U24620 (N_24620,N_20545,N_21766);
nor U24621 (N_24621,N_21622,N_20249);
or U24622 (N_24622,N_20498,N_22003);
nor U24623 (N_24623,N_22111,N_21741);
and U24624 (N_24624,N_21570,N_20004);
nor U24625 (N_24625,N_20235,N_21955);
nor U24626 (N_24626,N_20954,N_21752);
nor U24627 (N_24627,N_20693,N_22431);
or U24628 (N_24628,N_20644,N_21413);
nor U24629 (N_24629,N_20757,N_22355);
and U24630 (N_24630,N_22484,N_22218);
nor U24631 (N_24631,N_21159,N_20961);
and U24632 (N_24632,N_20791,N_20587);
and U24633 (N_24633,N_22266,N_20019);
or U24634 (N_24634,N_21031,N_20780);
and U24635 (N_24635,N_20170,N_22302);
or U24636 (N_24636,N_20307,N_22029);
nand U24637 (N_24637,N_20066,N_21812);
nor U24638 (N_24638,N_21598,N_21649);
xor U24639 (N_24639,N_22002,N_21729);
nand U24640 (N_24640,N_21683,N_22443);
xnor U24641 (N_24641,N_20493,N_21721);
and U24642 (N_24642,N_22278,N_20708);
xor U24643 (N_24643,N_20693,N_20542);
nor U24644 (N_24644,N_20986,N_21031);
nor U24645 (N_24645,N_20662,N_21146);
nand U24646 (N_24646,N_22290,N_21401);
nor U24647 (N_24647,N_21610,N_22115);
nand U24648 (N_24648,N_20799,N_21371);
and U24649 (N_24649,N_22220,N_22471);
or U24650 (N_24650,N_20561,N_21945);
nand U24651 (N_24651,N_21725,N_22242);
xor U24652 (N_24652,N_22319,N_21504);
nand U24653 (N_24653,N_21210,N_21273);
nand U24654 (N_24654,N_21078,N_21537);
xor U24655 (N_24655,N_20063,N_21039);
nand U24656 (N_24656,N_21539,N_21928);
or U24657 (N_24657,N_22425,N_22139);
nor U24658 (N_24658,N_21723,N_20700);
or U24659 (N_24659,N_22376,N_20429);
or U24660 (N_24660,N_22098,N_20310);
nand U24661 (N_24661,N_21576,N_21810);
and U24662 (N_24662,N_21575,N_20948);
nand U24663 (N_24663,N_20262,N_21370);
or U24664 (N_24664,N_20703,N_21030);
or U24665 (N_24665,N_22302,N_21687);
nand U24666 (N_24666,N_21185,N_21903);
nor U24667 (N_24667,N_21913,N_20408);
nand U24668 (N_24668,N_21452,N_21592);
nor U24669 (N_24669,N_21065,N_20532);
or U24670 (N_24670,N_21296,N_20255);
or U24671 (N_24671,N_21450,N_20600);
xnor U24672 (N_24672,N_21847,N_20559);
and U24673 (N_24673,N_20674,N_20385);
nand U24674 (N_24674,N_21643,N_21339);
and U24675 (N_24675,N_22062,N_22247);
nand U24676 (N_24676,N_21542,N_20596);
nor U24677 (N_24677,N_21278,N_21356);
or U24678 (N_24678,N_21274,N_22460);
and U24679 (N_24679,N_20921,N_21161);
and U24680 (N_24680,N_20345,N_21729);
or U24681 (N_24681,N_22229,N_21285);
or U24682 (N_24682,N_20405,N_20282);
and U24683 (N_24683,N_21230,N_21086);
nand U24684 (N_24684,N_21947,N_21629);
nand U24685 (N_24685,N_20689,N_21677);
xor U24686 (N_24686,N_21637,N_20979);
xnor U24687 (N_24687,N_20896,N_21594);
nand U24688 (N_24688,N_22326,N_22379);
nand U24689 (N_24689,N_20288,N_20069);
or U24690 (N_24690,N_20929,N_20139);
nor U24691 (N_24691,N_21612,N_20678);
xnor U24692 (N_24692,N_20682,N_20113);
nor U24693 (N_24693,N_22109,N_21909);
nand U24694 (N_24694,N_21400,N_20911);
or U24695 (N_24695,N_21160,N_22106);
and U24696 (N_24696,N_22327,N_22259);
nand U24697 (N_24697,N_22143,N_21754);
and U24698 (N_24698,N_20791,N_21388);
nor U24699 (N_24699,N_22481,N_22072);
nand U24700 (N_24700,N_20187,N_20509);
nor U24701 (N_24701,N_20950,N_21279);
nand U24702 (N_24702,N_21543,N_21559);
or U24703 (N_24703,N_21151,N_21338);
or U24704 (N_24704,N_22121,N_20209);
nand U24705 (N_24705,N_22463,N_22143);
nor U24706 (N_24706,N_21177,N_20662);
nor U24707 (N_24707,N_20323,N_22081);
or U24708 (N_24708,N_21408,N_20106);
or U24709 (N_24709,N_20064,N_21708);
nand U24710 (N_24710,N_21214,N_20038);
or U24711 (N_24711,N_21964,N_22411);
or U24712 (N_24712,N_22217,N_20998);
nand U24713 (N_24713,N_20571,N_21950);
and U24714 (N_24714,N_20824,N_21499);
nor U24715 (N_24715,N_21323,N_21414);
nor U24716 (N_24716,N_21520,N_21086);
and U24717 (N_24717,N_22199,N_22038);
and U24718 (N_24718,N_22212,N_22480);
xor U24719 (N_24719,N_20919,N_21915);
or U24720 (N_24720,N_21820,N_21258);
and U24721 (N_24721,N_21781,N_20446);
and U24722 (N_24722,N_22158,N_20004);
and U24723 (N_24723,N_21882,N_21952);
nor U24724 (N_24724,N_21839,N_21158);
nor U24725 (N_24725,N_21980,N_22255);
nor U24726 (N_24726,N_20726,N_21113);
nor U24727 (N_24727,N_21734,N_22461);
nor U24728 (N_24728,N_22002,N_21373);
nand U24729 (N_24729,N_20605,N_21306);
or U24730 (N_24730,N_21546,N_20638);
nor U24731 (N_24731,N_21333,N_21211);
or U24732 (N_24732,N_22180,N_20628);
nor U24733 (N_24733,N_21787,N_21351);
nand U24734 (N_24734,N_20453,N_21307);
nand U24735 (N_24735,N_20773,N_21936);
nor U24736 (N_24736,N_21554,N_21563);
nor U24737 (N_24737,N_20472,N_21282);
and U24738 (N_24738,N_20320,N_20772);
and U24739 (N_24739,N_20574,N_20278);
nor U24740 (N_24740,N_20829,N_20166);
nor U24741 (N_24741,N_21805,N_20241);
and U24742 (N_24742,N_21723,N_21350);
and U24743 (N_24743,N_20136,N_20589);
nand U24744 (N_24744,N_20504,N_20887);
nand U24745 (N_24745,N_22293,N_21831);
and U24746 (N_24746,N_20391,N_21334);
nand U24747 (N_24747,N_20517,N_22323);
and U24748 (N_24748,N_20867,N_20289);
nand U24749 (N_24749,N_21705,N_20796);
and U24750 (N_24750,N_22480,N_21969);
nor U24751 (N_24751,N_20940,N_20727);
nand U24752 (N_24752,N_20092,N_21861);
or U24753 (N_24753,N_21020,N_21196);
nor U24754 (N_24754,N_20426,N_22390);
or U24755 (N_24755,N_21144,N_22082);
or U24756 (N_24756,N_20713,N_20544);
or U24757 (N_24757,N_20100,N_20271);
and U24758 (N_24758,N_21404,N_20866);
and U24759 (N_24759,N_21353,N_21282);
or U24760 (N_24760,N_20926,N_20542);
or U24761 (N_24761,N_21966,N_20206);
and U24762 (N_24762,N_20637,N_22130);
xnor U24763 (N_24763,N_20783,N_21422);
and U24764 (N_24764,N_21317,N_20994);
or U24765 (N_24765,N_22359,N_22479);
or U24766 (N_24766,N_21265,N_21065);
and U24767 (N_24767,N_20449,N_20921);
and U24768 (N_24768,N_22301,N_21283);
or U24769 (N_24769,N_21344,N_22289);
nor U24770 (N_24770,N_20472,N_21939);
nor U24771 (N_24771,N_21822,N_20657);
xnor U24772 (N_24772,N_21434,N_22169);
or U24773 (N_24773,N_21613,N_22005);
or U24774 (N_24774,N_22423,N_22072);
or U24775 (N_24775,N_21578,N_20825);
and U24776 (N_24776,N_20592,N_21896);
nand U24777 (N_24777,N_21841,N_21579);
nor U24778 (N_24778,N_20976,N_20958);
and U24779 (N_24779,N_21556,N_21005);
nand U24780 (N_24780,N_22185,N_22491);
nor U24781 (N_24781,N_21081,N_21102);
nand U24782 (N_24782,N_21465,N_20973);
nor U24783 (N_24783,N_21753,N_21325);
or U24784 (N_24784,N_21889,N_20579);
or U24785 (N_24785,N_21494,N_21165);
nor U24786 (N_24786,N_21163,N_20728);
nor U24787 (N_24787,N_22457,N_20236);
and U24788 (N_24788,N_21032,N_20184);
or U24789 (N_24789,N_22354,N_20777);
and U24790 (N_24790,N_21064,N_22186);
nand U24791 (N_24791,N_20934,N_20307);
or U24792 (N_24792,N_20418,N_22047);
nand U24793 (N_24793,N_21732,N_21388);
nand U24794 (N_24794,N_20551,N_20801);
or U24795 (N_24795,N_21207,N_21018);
xnor U24796 (N_24796,N_20897,N_20370);
nand U24797 (N_24797,N_20298,N_21290);
nand U24798 (N_24798,N_22487,N_21617);
nand U24799 (N_24799,N_21361,N_21419);
or U24800 (N_24800,N_22329,N_22019);
nor U24801 (N_24801,N_20950,N_22363);
and U24802 (N_24802,N_20804,N_21349);
nand U24803 (N_24803,N_22142,N_22342);
nor U24804 (N_24804,N_20585,N_21972);
nor U24805 (N_24805,N_21614,N_22289);
and U24806 (N_24806,N_20118,N_20904);
nand U24807 (N_24807,N_22252,N_21669);
and U24808 (N_24808,N_20566,N_21899);
and U24809 (N_24809,N_22417,N_20721);
xor U24810 (N_24810,N_21044,N_21258);
nor U24811 (N_24811,N_20744,N_22427);
nand U24812 (N_24812,N_20870,N_22389);
nand U24813 (N_24813,N_21185,N_20228);
nor U24814 (N_24814,N_20367,N_20045);
nand U24815 (N_24815,N_22340,N_20963);
and U24816 (N_24816,N_20303,N_21969);
nand U24817 (N_24817,N_21017,N_20521);
nor U24818 (N_24818,N_20685,N_22052);
or U24819 (N_24819,N_20552,N_21672);
nand U24820 (N_24820,N_21541,N_22338);
nor U24821 (N_24821,N_22000,N_20683);
and U24822 (N_24822,N_20598,N_22482);
and U24823 (N_24823,N_21848,N_21682);
and U24824 (N_24824,N_21645,N_21799);
nand U24825 (N_24825,N_21824,N_21783);
nor U24826 (N_24826,N_21188,N_20053);
and U24827 (N_24827,N_20497,N_20905);
or U24828 (N_24828,N_20225,N_22002);
nor U24829 (N_24829,N_22078,N_20713);
or U24830 (N_24830,N_21279,N_20283);
and U24831 (N_24831,N_20112,N_21925);
xnor U24832 (N_24832,N_22115,N_21315);
nand U24833 (N_24833,N_20289,N_21259);
and U24834 (N_24834,N_21809,N_21521);
nand U24835 (N_24835,N_20672,N_20291);
nand U24836 (N_24836,N_21539,N_21672);
and U24837 (N_24837,N_22056,N_20244);
nand U24838 (N_24838,N_21639,N_22034);
nand U24839 (N_24839,N_20239,N_20616);
xor U24840 (N_24840,N_20799,N_21919);
nand U24841 (N_24841,N_20993,N_22174);
and U24842 (N_24842,N_20357,N_22421);
and U24843 (N_24843,N_20837,N_22331);
nand U24844 (N_24844,N_20586,N_20838);
or U24845 (N_24845,N_22389,N_21020);
and U24846 (N_24846,N_22259,N_21917);
or U24847 (N_24847,N_20067,N_21087);
or U24848 (N_24848,N_20895,N_20110);
nor U24849 (N_24849,N_22115,N_21185);
and U24850 (N_24850,N_20482,N_20916);
or U24851 (N_24851,N_22195,N_20586);
nor U24852 (N_24852,N_20869,N_20830);
and U24853 (N_24853,N_21620,N_20303);
nand U24854 (N_24854,N_21343,N_21059);
nand U24855 (N_24855,N_20350,N_21127);
nand U24856 (N_24856,N_21375,N_22284);
and U24857 (N_24857,N_21956,N_21026);
or U24858 (N_24858,N_21236,N_20353);
and U24859 (N_24859,N_21280,N_22337);
nor U24860 (N_24860,N_21001,N_21833);
nor U24861 (N_24861,N_20296,N_21269);
xnor U24862 (N_24862,N_20767,N_21518);
nand U24863 (N_24863,N_22118,N_20864);
nor U24864 (N_24864,N_20072,N_20600);
nor U24865 (N_24865,N_21175,N_20266);
and U24866 (N_24866,N_21169,N_22260);
xnor U24867 (N_24867,N_20372,N_21191);
nor U24868 (N_24868,N_21582,N_20676);
nor U24869 (N_24869,N_22015,N_20590);
or U24870 (N_24870,N_20195,N_21747);
nor U24871 (N_24871,N_21354,N_21537);
or U24872 (N_24872,N_21058,N_21625);
and U24873 (N_24873,N_20837,N_20801);
nand U24874 (N_24874,N_22210,N_21555);
nand U24875 (N_24875,N_20915,N_22297);
nand U24876 (N_24876,N_20221,N_22031);
xor U24877 (N_24877,N_22338,N_20777);
nor U24878 (N_24878,N_21457,N_20363);
nor U24879 (N_24879,N_20985,N_20285);
or U24880 (N_24880,N_21398,N_22352);
and U24881 (N_24881,N_20937,N_20410);
nor U24882 (N_24882,N_21713,N_22488);
nor U24883 (N_24883,N_21958,N_21760);
or U24884 (N_24884,N_21237,N_20449);
nand U24885 (N_24885,N_20888,N_22069);
nand U24886 (N_24886,N_21802,N_22430);
and U24887 (N_24887,N_21228,N_22008);
and U24888 (N_24888,N_20492,N_21166);
or U24889 (N_24889,N_20635,N_20577);
and U24890 (N_24890,N_22122,N_21295);
nand U24891 (N_24891,N_21906,N_22072);
or U24892 (N_24892,N_21443,N_21427);
and U24893 (N_24893,N_22457,N_20094);
nand U24894 (N_24894,N_20620,N_22008);
and U24895 (N_24895,N_21029,N_21128);
nand U24896 (N_24896,N_20078,N_20204);
nor U24897 (N_24897,N_20647,N_22198);
or U24898 (N_24898,N_20063,N_21673);
or U24899 (N_24899,N_20193,N_20708);
and U24900 (N_24900,N_20006,N_21771);
nor U24901 (N_24901,N_22259,N_20346);
nor U24902 (N_24902,N_20525,N_20629);
or U24903 (N_24903,N_20344,N_21978);
xor U24904 (N_24904,N_22034,N_21687);
or U24905 (N_24905,N_21834,N_20015);
nor U24906 (N_24906,N_20665,N_21755);
and U24907 (N_24907,N_21673,N_22030);
or U24908 (N_24908,N_20631,N_20186);
or U24909 (N_24909,N_20450,N_21020);
or U24910 (N_24910,N_21887,N_22457);
and U24911 (N_24911,N_21837,N_20358);
nand U24912 (N_24912,N_21534,N_20527);
nand U24913 (N_24913,N_20086,N_22362);
and U24914 (N_24914,N_21956,N_21498);
and U24915 (N_24915,N_22004,N_22260);
and U24916 (N_24916,N_21226,N_21794);
and U24917 (N_24917,N_21585,N_20398);
and U24918 (N_24918,N_20010,N_22198);
or U24919 (N_24919,N_20259,N_20643);
or U24920 (N_24920,N_20012,N_20658);
nor U24921 (N_24921,N_20995,N_21088);
nor U24922 (N_24922,N_20084,N_20169);
xor U24923 (N_24923,N_20432,N_22192);
or U24924 (N_24924,N_21039,N_21653);
and U24925 (N_24925,N_20229,N_21001);
nand U24926 (N_24926,N_21242,N_20981);
and U24927 (N_24927,N_22013,N_21268);
nor U24928 (N_24928,N_20446,N_20726);
and U24929 (N_24929,N_21189,N_22146);
xnor U24930 (N_24930,N_22217,N_21107);
nor U24931 (N_24931,N_22499,N_20668);
and U24932 (N_24932,N_20166,N_20709);
nand U24933 (N_24933,N_22444,N_22272);
nor U24934 (N_24934,N_20311,N_20727);
nand U24935 (N_24935,N_22202,N_20421);
nand U24936 (N_24936,N_21951,N_21572);
nor U24937 (N_24937,N_20141,N_22452);
nor U24938 (N_24938,N_20233,N_21917);
nand U24939 (N_24939,N_20292,N_20939);
and U24940 (N_24940,N_21331,N_20472);
nor U24941 (N_24941,N_22228,N_22137);
and U24942 (N_24942,N_21166,N_21302);
nand U24943 (N_24943,N_20891,N_22474);
and U24944 (N_24944,N_21323,N_22283);
or U24945 (N_24945,N_22473,N_21628);
xnor U24946 (N_24946,N_22263,N_20792);
nand U24947 (N_24947,N_22218,N_20451);
nor U24948 (N_24948,N_20237,N_21969);
nand U24949 (N_24949,N_21453,N_20710);
and U24950 (N_24950,N_20272,N_22461);
nand U24951 (N_24951,N_22467,N_20111);
or U24952 (N_24952,N_22197,N_21580);
nor U24953 (N_24953,N_21843,N_21491);
and U24954 (N_24954,N_21465,N_21738);
and U24955 (N_24955,N_20120,N_20625);
nand U24956 (N_24956,N_20398,N_21212);
or U24957 (N_24957,N_21878,N_21629);
xnor U24958 (N_24958,N_20680,N_20133);
and U24959 (N_24959,N_21842,N_21232);
or U24960 (N_24960,N_21492,N_22434);
and U24961 (N_24961,N_20972,N_20230);
nor U24962 (N_24962,N_21536,N_22333);
nor U24963 (N_24963,N_20194,N_22111);
and U24964 (N_24964,N_20765,N_21504);
nand U24965 (N_24965,N_22279,N_20094);
nor U24966 (N_24966,N_20009,N_21041);
nor U24967 (N_24967,N_20295,N_21006);
nand U24968 (N_24968,N_21415,N_20477);
nor U24969 (N_24969,N_21594,N_21426);
and U24970 (N_24970,N_20735,N_21131);
nand U24971 (N_24971,N_21160,N_22168);
nand U24972 (N_24972,N_21596,N_21736);
nor U24973 (N_24973,N_21162,N_20455);
nor U24974 (N_24974,N_21430,N_21493);
and U24975 (N_24975,N_21438,N_20475);
xor U24976 (N_24976,N_21020,N_21682);
nand U24977 (N_24977,N_20292,N_20570);
or U24978 (N_24978,N_21554,N_21704);
or U24979 (N_24979,N_20293,N_20796);
nand U24980 (N_24980,N_20611,N_20503);
or U24981 (N_24981,N_20788,N_21154);
or U24982 (N_24982,N_21866,N_22158);
nor U24983 (N_24983,N_20998,N_21569);
nor U24984 (N_24984,N_20195,N_20891);
or U24985 (N_24985,N_21678,N_20379);
and U24986 (N_24986,N_21979,N_22041);
or U24987 (N_24987,N_20313,N_21817);
nor U24988 (N_24988,N_20303,N_20252);
and U24989 (N_24989,N_21387,N_20878);
nand U24990 (N_24990,N_21101,N_21348);
nor U24991 (N_24991,N_20499,N_22430);
nand U24992 (N_24992,N_20861,N_21569);
xnor U24993 (N_24993,N_20508,N_21813);
and U24994 (N_24994,N_21923,N_21410);
nand U24995 (N_24995,N_22328,N_20242);
nor U24996 (N_24996,N_20100,N_21878);
nor U24997 (N_24997,N_21579,N_22430);
or U24998 (N_24998,N_20796,N_21865);
or U24999 (N_24999,N_22127,N_22061);
and U25000 (N_25000,N_23897,N_22870);
xor U25001 (N_25001,N_24546,N_23637);
or U25002 (N_25002,N_24632,N_24949);
xnor U25003 (N_25003,N_22612,N_24526);
nand U25004 (N_25004,N_22843,N_24338);
and U25005 (N_25005,N_24838,N_24140);
nor U25006 (N_25006,N_23295,N_24030);
nand U25007 (N_25007,N_23900,N_24864);
or U25008 (N_25008,N_24499,N_22754);
nand U25009 (N_25009,N_24688,N_22519);
nor U25010 (N_25010,N_22602,N_23397);
nor U25011 (N_25011,N_23902,N_24899);
and U25012 (N_25012,N_24804,N_23879);
nand U25013 (N_25013,N_24407,N_24649);
or U25014 (N_25014,N_24141,N_24859);
or U25015 (N_25015,N_23182,N_23613);
nand U25016 (N_25016,N_22712,N_23574);
nand U25017 (N_25017,N_24081,N_22962);
or U25018 (N_25018,N_23602,N_24795);
nor U25019 (N_25019,N_22773,N_22595);
nand U25020 (N_25020,N_23297,N_24462);
nand U25021 (N_25021,N_24591,N_22846);
nor U25022 (N_25022,N_23786,N_23199);
or U25023 (N_25023,N_24988,N_23383);
nand U25024 (N_25024,N_24729,N_23288);
or U25025 (N_25025,N_23649,N_23190);
or U25026 (N_25026,N_24093,N_22573);
and U25027 (N_25027,N_24353,N_24370);
and U25028 (N_25028,N_23329,N_23831);
xor U25029 (N_25029,N_24938,N_23527);
or U25030 (N_25030,N_24722,N_23091);
and U25031 (N_25031,N_24398,N_23701);
nand U25032 (N_25032,N_23954,N_23474);
xnor U25033 (N_25033,N_23721,N_23193);
or U25034 (N_25034,N_23100,N_22639);
nand U25035 (N_25035,N_23445,N_23338);
nor U25036 (N_25036,N_24281,N_22828);
xor U25037 (N_25037,N_23848,N_23370);
and U25038 (N_25038,N_23979,N_24461);
nand U25039 (N_25039,N_23884,N_24516);
nor U25040 (N_25040,N_23990,N_23513);
nand U25041 (N_25041,N_24507,N_23268);
and U25042 (N_25042,N_22837,N_24505);
or U25043 (N_25043,N_22545,N_23547);
nand U25044 (N_25044,N_24702,N_22874);
nand U25045 (N_25045,N_24563,N_23195);
nand U25046 (N_25046,N_22983,N_23022);
nor U25047 (N_25047,N_24612,N_23846);
and U25048 (N_25048,N_22804,N_22640);
xnor U25049 (N_25049,N_24029,N_23673);
or U25050 (N_25050,N_22501,N_23108);
or U25051 (N_25051,N_23362,N_24378);
nor U25052 (N_25052,N_22878,N_24173);
nor U25053 (N_25053,N_24144,N_23286);
or U25054 (N_25054,N_22582,N_24038);
xor U25055 (N_25055,N_23192,N_23728);
or U25056 (N_25056,N_22950,N_24900);
nor U25057 (N_25057,N_23388,N_24249);
and U25058 (N_25058,N_23097,N_23250);
or U25059 (N_25059,N_23978,N_24169);
nor U25060 (N_25060,N_23194,N_24957);
nor U25061 (N_25061,N_23044,N_24276);
xnor U25062 (N_25062,N_24786,N_23891);
or U25063 (N_25063,N_23928,N_24282);
nand U25064 (N_25064,N_24262,N_24316);
or U25065 (N_25065,N_24655,N_22802);
and U25066 (N_25066,N_22757,N_24454);
or U25067 (N_25067,N_23207,N_24801);
or U25068 (N_25068,N_24617,N_24481);
nor U25069 (N_25069,N_24349,N_23791);
nand U25070 (N_25070,N_22761,N_24968);
and U25071 (N_25071,N_24569,N_22951);
and U25072 (N_25072,N_23985,N_23430);
or U25073 (N_25073,N_23001,N_22551);
nand U25074 (N_25074,N_23943,N_23890);
or U25075 (N_25075,N_22738,N_22644);
xnor U25076 (N_25076,N_24672,N_24757);
nand U25077 (N_25077,N_24313,N_24011);
or U25078 (N_25078,N_22570,N_24912);
nand U25079 (N_25079,N_24978,N_23627);
or U25080 (N_25080,N_22966,N_24741);
or U25081 (N_25081,N_23765,N_22641);
nor U25082 (N_25082,N_23959,N_24180);
or U25083 (N_25083,N_23582,N_24130);
or U25084 (N_25084,N_23224,N_24844);
and U25085 (N_25085,N_23921,N_23096);
nor U25086 (N_25086,N_23013,N_22515);
xnor U25087 (N_25087,N_23822,N_24871);
or U25088 (N_25088,N_24597,N_23155);
nand U25089 (N_25089,N_24643,N_24965);
and U25090 (N_25090,N_23568,N_23368);
or U25091 (N_25091,N_23622,N_24110);
and U25092 (N_25092,N_22805,N_23534);
nand U25093 (N_25093,N_23107,N_23748);
nand U25094 (N_25094,N_24113,N_22981);
and U25095 (N_25095,N_22745,N_24626);
or U25096 (N_25096,N_24363,N_24682);
nor U25097 (N_25097,N_24830,N_24824);
nand U25098 (N_25098,N_22936,N_23781);
nand U25099 (N_25099,N_24645,N_24136);
and U25100 (N_25100,N_23188,N_22677);
or U25101 (N_25101,N_22642,N_23744);
or U25102 (N_25102,N_24556,N_23485);
nand U25103 (N_25103,N_23783,N_24037);
nand U25104 (N_25104,N_22539,N_22880);
nor U25105 (N_25105,N_24847,N_23840);
or U25106 (N_25106,N_24685,N_23023);
and U25107 (N_25107,N_23467,N_23006);
and U25108 (N_25108,N_23905,N_24399);
nand U25109 (N_25109,N_22584,N_24325);
and U25110 (N_25110,N_24427,N_23931);
xnor U25111 (N_25111,N_22635,N_24434);
nor U25112 (N_25112,N_23175,N_22540);
and U25113 (N_25113,N_23166,N_24792);
nor U25114 (N_25114,N_24204,N_23417);
or U25115 (N_25115,N_23715,N_23420);
and U25116 (N_25116,N_24225,N_24915);
nor U25117 (N_25117,N_24101,N_24855);
and U25118 (N_25118,N_24761,N_24480);
xnor U25119 (N_25119,N_24845,N_24028);
and U25120 (N_25120,N_23641,N_24634);
xor U25121 (N_25121,N_22624,N_23165);
nor U25122 (N_25122,N_23685,N_24456);
and U25123 (N_25123,N_24721,N_24740);
or U25124 (N_25124,N_23306,N_23614);
nand U25125 (N_25125,N_23148,N_23153);
nor U25126 (N_25126,N_24298,N_22935);
xnor U25127 (N_25127,N_23694,N_22796);
nand U25128 (N_25128,N_23828,N_24587);
and U25129 (N_25129,N_24050,N_22821);
or U25130 (N_25130,N_22788,N_24687);
or U25131 (N_25131,N_22800,N_24942);
or U25132 (N_25132,N_23291,N_24537);
or U25133 (N_25133,N_24941,N_22562);
nand U25134 (N_25134,N_23626,N_24084);
and U25135 (N_25135,N_23593,N_24498);
nand U25136 (N_25136,N_23855,N_24438);
and U25137 (N_25137,N_23010,N_24483);
nand U25138 (N_25138,N_24976,N_24263);
nor U25139 (N_25139,N_23341,N_24317);
or U25140 (N_25140,N_23633,N_23551);
nor U25141 (N_25141,N_24787,N_24286);
or U25142 (N_25142,N_23779,N_23259);
and U25143 (N_25143,N_24016,N_23907);
xor U25144 (N_25144,N_23745,N_23693);
or U25145 (N_25145,N_23455,N_22702);
nand U25146 (N_25146,N_22939,N_24035);
or U25147 (N_25147,N_23965,N_24337);
or U25148 (N_25148,N_22986,N_23560);
nand U25149 (N_25149,N_22668,N_23039);
nand U25150 (N_25150,N_24832,N_24633);
nor U25151 (N_25151,N_23048,N_24416);
and U25152 (N_25152,N_24272,N_24239);
nor U25153 (N_25153,N_23367,N_22662);
nand U25154 (N_25154,N_24241,N_23147);
nand U25155 (N_25155,N_24319,N_24202);
nand U25156 (N_25156,N_23599,N_24040);
and U25157 (N_25157,N_23081,N_24376);
or U25158 (N_25158,N_23734,N_23677);
or U25159 (N_25159,N_23285,N_23646);
nand U25160 (N_25160,N_24385,N_23282);
and U25161 (N_25161,N_23446,N_23760);
nor U25162 (N_25162,N_24441,N_22947);
nor U25163 (N_25163,N_24259,N_24477);
and U25164 (N_25164,N_24760,N_23323);
xnor U25165 (N_25165,N_24223,N_24958);
nand U25166 (N_25166,N_24921,N_23178);
and U25167 (N_25167,N_24464,N_23079);
nand U25168 (N_25168,N_22603,N_24167);
and U25169 (N_25169,N_23032,N_24161);
or U25170 (N_25170,N_23443,N_24548);
nand U25171 (N_25171,N_24079,N_23804);
or U25172 (N_25172,N_22750,N_23955);
nor U25173 (N_25173,N_24125,N_24596);
and U25174 (N_25174,N_22681,N_22513);
or U25175 (N_25175,N_23495,N_23055);
nand U25176 (N_25176,N_23517,N_24908);
and U25177 (N_25177,N_24022,N_23819);
and U25178 (N_25178,N_23761,N_23428);
nand U25179 (N_25179,N_22553,N_22849);
and U25180 (N_25180,N_24100,N_24087);
xnor U25181 (N_25181,N_24493,N_23380);
nand U25182 (N_25182,N_23720,N_23016);
xnor U25183 (N_25183,N_23137,N_23336);
and U25184 (N_25184,N_23363,N_23413);
or U25185 (N_25185,N_22675,N_24515);
and U25186 (N_25186,N_23398,N_24390);
nor U25187 (N_25187,N_23895,N_23688);
and U25188 (N_25188,N_22608,N_23557);
nand U25189 (N_25189,N_24068,N_24867);
or U25190 (N_25190,N_23575,N_23117);
nand U25191 (N_25191,N_22910,N_22543);
xnor U25192 (N_25192,N_22799,N_23466);
and U25193 (N_25193,N_24163,N_24767);
nor U25194 (N_25194,N_24391,N_23631);
nor U25195 (N_25195,N_23735,N_24102);
xor U25196 (N_25196,N_23678,N_23986);
xor U25197 (N_25197,N_23403,N_24166);
nand U25198 (N_25198,N_24153,N_23957);
nor U25199 (N_25199,N_22974,N_24913);
xnor U25200 (N_25200,N_23841,N_24808);
and U25201 (N_25201,N_23115,N_22779);
or U25202 (N_25202,N_22721,N_24265);
nor U25203 (N_25203,N_22833,N_23885);
or U25204 (N_25204,N_23670,N_24268);
and U25205 (N_25205,N_23703,N_23431);
nor U25206 (N_25206,N_24120,N_23519);
nand U25207 (N_25207,N_23658,N_23508);
xor U25208 (N_25208,N_23040,N_23889);
or U25209 (N_25209,N_24952,N_24565);
and U25210 (N_25210,N_23852,N_23909);
or U25211 (N_25211,N_23078,N_22782);
nor U25212 (N_25212,N_22891,N_22563);
xor U25213 (N_25213,N_22917,N_22905);
xor U25214 (N_25214,N_24288,N_23283);
or U25215 (N_25215,N_24646,N_24670);
or U25216 (N_25216,N_23812,N_24254);
nand U25217 (N_25217,N_23656,N_22520);
or U25218 (N_25218,N_22998,N_24625);
nand U25219 (N_25219,N_24692,N_22708);
or U25220 (N_25220,N_23869,N_22728);
xor U25221 (N_25221,N_22847,N_23315);
and U25222 (N_25222,N_24051,N_22529);
and U25223 (N_25223,N_23103,N_24200);
nor U25224 (N_25224,N_24024,N_23436);
xnor U25225 (N_25225,N_23186,N_23334);
nand U25226 (N_25226,N_22895,N_23011);
xor U25227 (N_25227,N_24583,N_24196);
xnor U25228 (N_25228,N_23709,N_23950);
and U25229 (N_25229,N_24064,N_24007);
or U25230 (N_25230,N_23857,N_24530);
or U25231 (N_25231,N_23144,N_23083);
nor U25232 (N_25232,N_24137,N_23882);
nand U25233 (N_25233,N_24106,N_22673);
xor U25234 (N_25234,N_23507,N_23316);
xor U25235 (N_25235,N_24994,N_23922);
and U25236 (N_25236,N_23887,N_22541);
xnor U25237 (N_25237,N_23894,N_24224);
and U25238 (N_25238,N_24457,N_24212);
xor U25239 (N_25239,N_24570,N_24524);
nand U25240 (N_25240,N_24798,N_22789);
nand U25241 (N_25241,N_23939,N_23768);
nor U25242 (N_25242,N_23934,N_24598);
or U25243 (N_25243,N_24105,N_23465);
nor U25244 (N_25244,N_24594,N_24025);
nand U25245 (N_25245,N_23941,N_23350);
or U25246 (N_25246,N_22868,N_24920);
nor U25247 (N_25247,N_24049,N_24227);
or U25248 (N_25248,N_22625,N_24631);
nor U25249 (N_25249,N_24420,N_24255);
nand U25250 (N_25250,N_24812,N_23667);
nand U25251 (N_25251,N_24473,N_24532);
xor U25252 (N_25252,N_24359,N_24763);
nand U25253 (N_25253,N_23300,N_22948);
or U25254 (N_25254,N_24788,N_23378);
nand U25255 (N_25255,N_23643,N_24094);
nand U25256 (N_25256,N_23699,N_24898);
nand U25257 (N_25257,N_22767,N_23002);
and U25258 (N_25258,N_23874,N_23152);
or U25259 (N_25259,N_23080,N_22652);
nor U25260 (N_25260,N_23119,N_23415);
nand U25261 (N_25261,N_24246,N_22622);
or U25262 (N_25262,N_22588,N_23865);
nand U25263 (N_25263,N_23844,N_22954);
xnor U25264 (N_25264,N_22985,N_24863);
and U25265 (N_25265,N_24836,N_23470);
nand U25266 (N_25266,N_23414,N_22806);
nand U25267 (N_25267,N_23104,N_23948);
and U25268 (N_25268,N_23966,N_23516);
nor U25269 (N_25269,N_22872,N_24573);
and U25270 (N_25270,N_23974,N_24593);
xor U25271 (N_25271,N_23390,N_22912);
and U25272 (N_25272,N_23893,N_23871);
nor U25273 (N_25273,N_24476,N_22734);
and U25274 (N_25274,N_22812,N_23838);
nand U25275 (N_25275,N_22686,N_24356);
and U25276 (N_25276,N_22975,N_22537);
nor U25277 (N_25277,N_23354,N_24116);
and U25278 (N_25278,N_23468,N_23662);
xor U25279 (N_25279,N_23377,N_24509);
and U25280 (N_25280,N_23025,N_24642);
nor U25281 (N_25281,N_23784,N_23853);
nor U25282 (N_25282,N_23037,N_24354);
nor U25283 (N_25283,N_23294,N_23142);
xor U25284 (N_25284,N_23384,N_22690);
or U25285 (N_25285,N_23053,N_24709);
and U25286 (N_25286,N_22502,N_23442);
nor U25287 (N_25287,N_22506,N_24868);
xor U25288 (N_25288,N_24243,N_24768);
or U25289 (N_25289,N_22769,N_24175);
or U25290 (N_25290,N_23070,N_23608);
or U25291 (N_25291,N_24096,N_24168);
nand U25292 (N_25292,N_24292,N_22660);
xor U25293 (N_25293,N_24848,N_24214);
and U25294 (N_25294,N_24657,N_24531);
or U25295 (N_25295,N_24665,N_24036);
and U25296 (N_25296,N_23548,N_24566);
nand U25297 (N_25297,N_23752,N_22887);
xor U25298 (N_25298,N_24628,N_22760);
nor U25299 (N_25299,N_24061,N_23753);
or U25300 (N_25300,N_24329,N_22959);
or U25301 (N_25301,N_22654,N_22546);
and U25302 (N_25302,N_23481,N_24793);
nand U25303 (N_25303,N_22834,N_24162);
nand U25304 (N_25304,N_23727,N_23603);
nor U25305 (N_25305,N_24108,N_24380);
nor U25306 (N_25306,N_23041,N_23122);
or U25307 (N_25307,N_24675,N_23059);
xnor U25308 (N_25308,N_23569,N_23225);
nand U25309 (N_25309,N_23652,N_22973);
or U25310 (N_25310,N_22523,N_22946);
nor U25311 (N_25311,N_22739,N_24719);
or U25312 (N_25312,N_24327,N_24652);
nand U25313 (N_25313,N_24584,N_22964);
nor U25314 (N_25314,N_23689,N_23346);
nand U25315 (N_25315,N_22809,N_23851);
nor U25316 (N_25316,N_23510,N_24235);
nor U25317 (N_25317,N_22671,N_24790);
nor U25318 (N_25318,N_24659,N_24261);
and U25319 (N_25319,N_22934,N_24662);
nor U25320 (N_25320,N_22763,N_23679);
or U25321 (N_25321,N_24910,N_24890);
or U25322 (N_25322,N_24295,N_23644);
nand U25323 (N_25323,N_23988,N_24766);
or U25324 (N_25324,N_23014,N_23837);
or U25325 (N_25325,N_23374,N_23591);
and U25326 (N_25326,N_24046,N_22617);
and U25327 (N_25327,N_24070,N_24318);
nor U25328 (N_25328,N_23043,N_22716);
and U25329 (N_25329,N_24197,N_23161);
nor U25330 (N_25330,N_23307,N_24213);
and U25331 (N_25331,N_23254,N_22882);
xor U25332 (N_25332,N_23475,N_24529);
nor U25333 (N_25333,N_23304,N_24321);
nand U25334 (N_25334,N_23808,N_23769);
and U25335 (N_25335,N_24660,N_24220);
nor U25336 (N_25336,N_24901,N_22748);
or U25337 (N_25337,N_23234,N_24063);
nor U25338 (N_25338,N_23886,N_23056);
and U25339 (N_25339,N_23977,N_24310);
nor U25340 (N_25340,N_24723,N_24334);
or U25341 (N_25341,N_23826,N_22719);
nor U25342 (N_25342,N_23425,N_24572);
xnor U25343 (N_25343,N_23924,N_23916);
nor U25344 (N_25344,N_24713,N_22718);
nor U25345 (N_25345,N_23129,N_23710);
nand U25346 (N_25346,N_24240,N_23324);
xor U25347 (N_25347,N_24852,N_24605);
nand U25348 (N_25348,N_23372,N_24242);
nand U25349 (N_25349,N_23141,N_23550);
nand U25350 (N_25350,N_23127,N_22587);
xor U25351 (N_25351,N_22791,N_22916);
nor U25352 (N_25352,N_23167,N_22700);
nand U25353 (N_25353,N_24060,N_23584);
nand U25354 (N_25354,N_23628,N_24020);
nor U25355 (N_25355,N_23086,N_24624);
and U25356 (N_25356,N_23275,N_22670);
nor U25357 (N_25357,N_23337,N_23116);
xor U25358 (N_25358,N_23859,N_23320);
nor U25359 (N_25359,N_23231,N_23706);
or U25360 (N_25360,N_22938,N_23702);
nor U25361 (N_25361,N_23946,N_24730);
and U25362 (N_25362,N_22967,N_24411);
nor U25363 (N_25363,N_22830,N_22751);
or U25364 (N_25364,N_24034,N_22982);
xor U25365 (N_25365,N_23008,N_24233);
nor U25366 (N_25366,N_23064,N_22928);
and U25367 (N_25367,N_22899,N_22811);
or U25368 (N_25368,N_23424,N_24485);
and U25369 (N_25369,N_23272,N_24728);
nor U25370 (N_25370,N_22886,N_23215);
nor U25371 (N_25371,N_23034,N_23312);
and U25372 (N_25372,N_22988,N_23197);
and U25373 (N_25373,N_24925,N_23191);
and U25374 (N_25374,N_23716,N_23118);
and U25375 (N_25375,N_23801,N_22643);
or U25376 (N_25376,N_24135,N_22869);
nand U25377 (N_25377,N_23502,N_22577);
nor U25378 (N_25378,N_24751,N_23766);
nor U25379 (N_25379,N_23252,N_24897);
or U25380 (N_25380,N_23732,N_24075);
or U25381 (N_25381,N_23065,N_22691);
nand U25382 (N_25382,N_24271,N_24950);
nand U25383 (N_25383,N_24935,N_23409);
xnor U25384 (N_25384,N_24273,N_24746);
nand U25385 (N_25385,N_23206,N_24216);
or U25386 (N_25386,N_23563,N_22535);
xnor U25387 (N_25387,N_22667,N_23311);
nand U25388 (N_25388,N_22558,N_23705);
nor U25389 (N_25389,N_24508,N_22787);
nor U25390 (N_25390,N_24208,N_22579);
and U25391 (N_25391,N_23216,N_22969);
nor U25392 (N_25392,N_24071,N_24082);
or U25393 (N_25393,N_24171,N_23963);
nand U25394 (N_25394,N_22932,N_24850);
and U25395 (N_25395,N_23149,N_22924);
nand U25396 (N_25396,N_22857,N_22749);
or U25397 (N_25397,N_24823,N_23305);
nor U25398 (N_25398,N_23723,N_22785);
or U25399 (N_25399,N_23799,N_23491);
xnor U25400 (N_25400,N_23429,N_22632);
and U25401 (N_25401,N_24033,N_24504);
nor U25402 (N_25402,N_24435,N_24205);
nor U25403 (N_25403,N_23531,N_24145);
and U25404 (N_25404,N_23395,N_24371);
nand U25405 (N_25405,N_23621,N_23993);
nor U25406 (N_25406,N_23412,N_24959);
and U25407 (N_25407,N_23578,N_22972);
and U25408 (N_25408,N_23625,N_24917);
and U25409 (N_25409,N_24000,N_24443);
nand U25410 (N_25410,N_24817,N_24496);
or U25411 (N_25411,N_22596,N_24486);
or U25412 (N_25412,N_24849,N_24335);
and U25413 (N_25413,N_24977,N_22518);
nand U25414 (N_25414,N_24820,N_22914);
and U25415 (N_25415,N_22547,N_23497);
nor U25416 (N_25416,N_22621,N_24139);
xnor U25417 (N_25417,N_24275,N_22999);
nor U25418 (N_25418,N_22875,N_23824);
xor U25419 (N_25419,N_24933,N_24878);
and U25420 (N_25420,N_24708,N_24403);
nor U25421 (N_25421,N_24858,N_24637);
xor U25422 (N_25422,N_22979,N_22774);
nor U25423 (N_25423,N_23751,N_23883);
nor U25424 (N_25424,N_24344,N_23746);
xnor U25425 (N_25425,N_24001,N_24718);
xor U25426 (N_25426,N_24734,N_24127);
xor U25427 (N_25427,N_24112,N_24129);
nand U25428 (N_25428,N_22861,N_22729);
nor U25429 (N_25429,N_22560,N_22710);
nor U25430 (N_25430,N_24773,N_23636);
nand U25431 (N_25431,N_23787,N_24973);
nor U25432 (N_25432,N_24415,N_23146);
or U25433 (N_25433,N_24562,N_22957);
xnor U25434 (N_25434,N_22693,N_24111);
or U25435 (N_25435,N_24188,N_22770);
and U25436 (N_25436,N_23061,N_23998);
or U25437 (N_25437,N_24339,N_23313);
nand U25438 (N_25438,N_23333,N_22548);
nor U25439 (N_25439,N_23763,N_24707);
and U25440 (N_25440,N_23717,N_24043);
nor U25441 (N_25441,N_24154,N_22853);
or U25442 (N_25442,N_23968,N_24807);
nor U25443 (N_25443,N_24870,N_24876);
or U25444 (N_25444,N_24495,N_22568);
or U25445 (N_25445,N_23351,N_23618);
xor U25446 (N_25446,N_22601,N_24929);
nor U25447 (N_25447,N_23901,N_24635);
and U25448 (N_25448,N_23066,N_23668);
nand U25449 (N_25449,N_23981,N_24669);
or U25450 (N_25450,N_22589,N_23795);
nand U25451 (N_25451,N_22695,N_23686);
nor U25452 (N_25452,N_24698,N_22715);
nand U25453 (N_25453,N_22552,N_23947);
and U25454 (N_25454,N_23898,N_24712);
or U25455 (N_25455,N_23406,N_24658);
nor U25456 (N_25456,N_24873,N_24616);
nor U25457 (N_25457,N_24187,N_22741);
xnor U25458 (N_25458,N_23579,N_23482);
nor U25459 (N_25459,N_24742,N_23340);
and U25460 (N_25460,N_24437,N_23394);
or U25461 (N_25461,N_24361,N_23964);
nand U25462 (N_25462,N_24326,N_22942);
nor U25463 (N_25463,N_22663,N_22937);
and U25464 (N_25464,N_22883,N_22755);
nor U25465 (N_25465,N_24877,N_22585);
nor U25466 (N_25466,N_24641,N_23980);
nor U25467 (N_25467,N_23743,N_24078);
nor U25468 (N_25468,N_23084,N_24544);
or U25469 (N_25469,N_23544,N_23332);
or U25470 (N_25470,N_23208,N_23456);
or U25471 (N_25471,N_23348,N_24303);
and U25472 (N_25472,N_23211,N_23233);
and U25473 (N_25473,N_23049,N_24442);
and U25474 (N_25474,N_22978,N_23847);
nor U25475 (N_25475,N_24745,N_22907);
or U25476 (N_25476,N_24513,N_24375);
nand U25477 (N_25477,N_23526,N_24693);
nor U25478 (N_25478,N_23484,N_22709);
or U25479 (N_25479,N_23441,N_23450);
nand U25480 (N_25480,N_22664,N_22628);
xnor U25481 (N_25481,N_24600,N_23663);
nor U25482 (N_25482,N_23512,N_23447);
or U25483 (N_25483,N_24727,N_23310);
nand U25484 (N_25484,N_24814,N_22864);
and U25485 (N_25485,N_23212,N_24260);
nor U25486 (N_25486,N_24117,N_22680);
xnor U25487 (N_25487,N_23472,N_23226);
nand U25488 (N_25488,N_23094,N_24603);
and U25489 (N_25489,N_24460,N_22897);
nor U25490 (N_25490,N_24664,N_23642);
or U25491 (N_25491,N_24512,N_22658);
xnor U25492 (N_25492,N_24392,N_24463);
xnor U25493 (N_25493,N_23892,N_24429);
nand U25494 (N_25494,N_23558,N_23160);
and U25495 (N_25495,N_24618,N_24575);
nand U25496 (N_25496,N_23478,N_24066);
nor U25497 (N_25497,N_23085,N_23845);
and U25498 (N_25498,N_22871,N_24553);
nor U25499 (N_25499,N_22555,N_24433);
nor U25500 (N_25500,N_22775,N_24369);
and U25501 (N_25501,N_22724,N_22820);
or U25502 (N_25502,N_24322,N_23878);
nand U25503 (N_25503,N_24244,N_23407);
nor U25504 (N_25504,N_24384,N_24903);
or U25505 (N_25505,N_22704,N_23553);
nor U25506 (N_25506,N_23913,N_22534);
nand U25507 (N_25507,N_24995,N_24882);
xnor U25508 (N_25508,N_24484,N_23776);
or U25509 (N_25509,N_24615,N_24955);
nor U25510 (N_25510,N_23274,N_22778);
and U25511 (N_25511,N_23532,N_24654);
nand U25512 (N_25512,N_23994,N_24364);
nand U25513 (N_25513,N_24157,N_24866);
nand U25514 (N_25514,N_23873,N_24301);
nand U25515 (N_25515,N_24835,N_23598);
and U25516 (N_25516,N_24956,N_23210);
nor U25517 (N_25517,N_23772,N_23266);
nor U25518 (N_25518,N_22503,N_23279);
and U25519 (N_25519,N_23352,N_24092);
or U25520 (N_25520,N_24183,N_23205);
or U25521 (N_25521,N_23690,N_24520);
and U25522 (N_25522,N_22958,N_24452);
or U25523 (N_25523,N_23358,N_24198);
nor U25524 (N_25524,N_24843,N_23322);
or U25525 (N_25525,N_24440,N_24684);
and U25526 (N_25526,N_23671,N_24518);
and U25527 (N_25527,N_24706,N_23523);
xor U25528 (N_25528,N_23648,N_22593);
and U25529 (N_25529,N_23219,N_24019);
nor U25530 (N_25530,N_22851,N_23536);
or U25531 (N_25531,N_23817,N_24737);
nand U25532 (N_25532,N_22881,N_23836);
nand U25533 (N_25533,N_23396,N_23938);
nand U25534 (N_25534,N_24571,N_24347);
and U25535 (N_25535,N_22747,N_24796);
xor U25536 (N_25536,N_24426,N_24311);
and U25537 (N_25537,N_23543,N_22634);
nor U25538 (N_25538,N_23169,N_23493);
nor U25539 (N_25539,N_22933,N_24342);
nand U25540 (N_25540,N_23401,N_24896);
and U25541 (N_25541,N_24138,N_23704);
or U25542 (N_25542,N_23251,N_23058);
and U25543 (N_25543,N_22971,N_22713);
nor U25544 (N_25544,N_23780,N_22829);
or U25545 (N_25545,N_24217,N_24080);
and U25546 (N_25546,N_23615,N_23028);
nand U25547 (N_25547,N_24422,N_24164);
xnor U25548 (N_25548,N_24536,N_23045);
or U25549 (N_25549,N_23114,N_24229);
and U25550 (N_25550,N_24372,N_23856);
or U25551 (N_25551,N_23927,N_24891);
nand U25552 (N_25552,N_24122,N_22701);
nand U25553 (N_25553,N_22901,N_24013);
or U25554 (N_25554,N_24045,N_24880);
nor U25555 (N_25555,N_23570,N_24232);
or U25556 (N_25556,N_23778,N_24054);
nand U25557 (N_25557,N_22583,N_23459);
and U25558 (N_25558,N_23733,N_22525);
and U25559 (N_25559,N_22530,N_23075);
or U25560 (N_25560,N_23835,N_24449);
and U25561 (N_25561,N_24827,N_23290);
and U25562 (N_25562,N_23138,N_22841);
and U25563 (N_25563,N_24888,N_24750);
nor U25564 (N_25564,N_24699,N_22599);
nand U25565 (N_25565,N_23842,N_23669);
nand U25566 (N_25566,N_22963,N_24165);
and U25567 (N_25567,N_24404,N_23174);
xor U25568 (N_25568,N_24410,N_24602);
or U25569 (N_25569,N_23019,N_24041);
nand U25570 (N_25570,N_24018,N_23680);
nand U25571 (N_25571,N_23738,N_22554);
nand U25572 (N_25572,N_23418,N_22819);
and U25573 (N_25573,N_24279,N_23026);
nor U25574 (N_25574,N_22771,N_22844);
and U25575 (N_25575,N_22666,N_23009);
xor U25576 (N_25576,N_22656,N_22561);
or U25577 (N_25577,N_23814,N_23408);
xor U25578 (N_25578,N_24985,N_24002);
nand U25579 (N_25579,N_24776,N_23235);
and U25580 (N_25580,N_22703,N_22890);
or U25581 (N_25581,N_23213,N_23712);
or U25582 (N_25582,N_23095,N_24436);
xor U25583 (N_25583,N_24775,N_24991);
and U25584 (N_25584,N_24738,N_24307);
and U25585 (N_25585,N_24393,N_24674);
or U25586 (N_25586,N_24613,N_23592);
and U25587 (N_25587,N_24283,N_23344);
or U25588 (N_25588,N_22996,N_22609);
nand U25589 (N_25589,N_23506,N_23287);
nand U25590 (N_25590,N_24234,N_24032);
xor U25591 (N_25591,N_24131,N_22648);
nor U25592 (N_25592,N_23449,N_24609);
nor U25593 (N_25593,N_24510,N_22618);
nor U25594 (N_25594,N_24954,N_23452);
or U25595 (N_25595,N_23379,N_24539);
nand U25596 (N_25596,N_22835,N_23426);
nor U25597 (N_25597,N_24931,N_23912);
nand U25598 (N_25598,N_24946,N_23432);
xnor U25599 (N_25599,N_23217,N_24606);
or U25600 (N_25600,N_22682,N_24521);
or U25601 (N_25601,N_22765,N_22813);
nand U25602 (N_25602,N_22904,N_23807);
and U25603 (N_25603,N_24382,N_24986);
nor U25604 (N_25604,N_24599,N_24661);
nor U25605 (N_25605,N_23469,N_22736);
or U25606 (N_25606,N_23479,N_24758);
or U25607 (N_25607,N_24947,N_23330);
and U25608 (N_25608,N_23820,N_24818);
and U25609 (N_25609,N_22902,N_23528);
xor U25610 (N_25610,N_23764,N_23813);
or U25611 (N_25611,N_23278,N_24846);
or U25612 (N_25612,N_24277,N_24340);
or U25613 (N_25613,N_23184,N_24549);
nand U25614 (N_25614,N_22696,N_24015);
nor U25615 (N_25615,N_24269,N_23750);
nand U25616 (N_25616,N_22892,N_24782);
nand U25617 (N_25617,N_24860,N_24455);
xor U25618 (N_25618,N_23908,N_22792);
or U25619 (N_25619,N_23872,N_24251);
or U25620 (N_25620,N_24417,N_23533);
or U25621 (N_25621,N_24803,N_23573);
nor U25622 (N_25622,N_22722,N_23438);
nor U25623 (N_25623,N_23404,N_23936);
or U25624 (N_25624,N_23619,N_22688);
or U25625 (N_25625,N_24176,N_24009);
nand U25626 (N_25626,N_23421,N_23089);
or U25627 (N_25627,N_24621,N_23419);
or U25628 (N_25628,N_23494,N_23803);
xnor U25629 (N_25629,N_24577,N_22645);
or U25630 (N_25630,N_24258,N_23366);
nor U25631 (N_25631,N_23566,N_22885);
nor U25632 (N_25632,N_24911,N_24736);
nor U25633 (N_25633,N_24614,N_22840);
xnor U25634 (N_25634,N_23223,N_23969);
nor U25635 (N_25635,N_22706,N_24474);
nand U25636 (N_25636,N_23681,N_24373);
and U25637 (N_25637,N_24151,N_23503);
nor U25638 (N_25638,N_24379,N_24012);
or U25639 (N_25639,N_23018,N_22814);
xnor U25640 (N_25640,N_24466,N_23995);
nand U25641 (N_25641,N_22542,N_23247);
xnor U25642 (N_25642,N_24695,N_24749);
xnor U25643 (N_25643,N_23610,N_24568);
and U25644 (N_25644,N_23371,N_24190);
nor U25645 (N_25645,N_24813,N_24998);
or U25646 (N_25646,N_24124,N_22517);
and U25647 (N_25647,N_24185,N_24350);
nor U25648 (N_25648,N_22649,N_24589);
nor U25649 (N_25649,N_23017,N_23711);
and U25650 (N_25650,N_24252,N_24388);
or U25651 (N_25651,N_24178,N_24926);
and U25652 (N_25652,N_24547,N_24627);
nor U25653 (N_25653,N_24089,N_24097);
nand U25654 (N_25654,N_24648,N_22915);
nand U25655 (N_25655,N_23168,N_24039);
nand U25656 (N_25656,N_23477,N_22610);
xnor U25657 (N_25657,N_23522,N_23027);
or U25658 (N_25658,N_24971,N_24152);
or U25659 (N_25659,N_24759,N_23657);
nor U25660 (N_25660,N_24330,N_24799);
nor U25661 (N_25661,N_22726,N_22918);
nor U25662 (N_25662,N_24992,N_23473);
nand U25663 (N_25663,N_24647,N_23674);
and U25664 (N_25664,N_22858,N_22822);
nor U25665 (N_25665,N_23942,N_23806);
nand U25666 (N_25666,N_23758,N_22731);
nand U25667 (N_25667,N_23640,N_23464);
nor U25668 (N_25668,N_24290,N_24472);
and U25669 (N_25669,N_24756,N_22557);
nor U25670 (N_25670,N_24748,N_24927);
nand U25671 (N_25671,N_23248,N_24439);
and U25672 (N_25672,N_24245,N_24887);
or U25673 (N_25673,N_22629,N_23318);
xor U25674 (N_25674,N_22659,N_22862);
nor U25675 (N_25675,N_24305,N_23020);
or U25676 (N_25676,N_22637,N_24837);
and U25677 (N_25677,N_22961,N_24228);
nor U25678 (N_25678,N_24128,N_23770);
and U25679 (N_25679,N_22679,N_23364);
or U25680 (N_25680,N_23754,N_22859);
nor U25681 (N_25681,N_23971,N_22574);
nor U25682 (N_25682,N_24052,N_22894);
or U25683 (N_25683,N_24148,N_23243);
nand U25684 (N_25684,N_24491,N_24826);
nand U25685 (N_25685,N_24236,N_24511);
nor U25686 (N_25686,N_23308,N_24656);
and U25687 (N_25687,N_23005,N_22909);
and U25688 (N_25688,N_22650,N_23896);
nor U25689 (N_25689,N_23539,N_22965);
and U25690 (N_25690,N_23914,N_24085);
nor U25691 (N_25691,N_23911,N_23373);
nor U25692 (N_25692,N_22927,N_24360);
and U25693 (N_25693,N_23740,N_23792);
or U25694 (N_25694,N_22735,N_23376);
nand U25695 (N_25695,N_23177,N_24851);
and U25696 (N_25696,N_24253,N_24405);
nand U25697 (N_25697,N_23264,N_24557);
or U25698 (N_25698,N_22759,N_22943);
nor U25699 (N_25699,N_23940,N_24678);
xor U25700 (N_25700,N_24006,N_24266);
nor U25701 (N_25701,N_24753,N_22565);
and U25702 (N_25702,N_24964,N_24471);
nor U25703 (N_25703,N_24209,N_23256);
or U25704 (N_25704,N_22955,N_23183);
and U25705 (N_25705,N_23355,N_23258);
nand U25706 (N_25706,N_23860,N_23876);
nand U25707 (N_25707,N_22879,N_23833);
or U25708 (N_25708,N_24755,N_24989);
and U25709 (N_25709,N_24284,N_24972);
nor U25710 (N_25710,N_23777,N_23269);
and U25711 (N_25711,N_23796,N_24104);
nand U25712 (N_25712,N_23695,N_24943);
and U25713 (N_25713,N_22991,N_23024);
and U25714 (N_25714,N_24922,N_23236);
nand U25715 (N_25715,N_24555,N_22606);
nand U25716 (N_25716,N_24783,N_22810);
nand U25717 (N_25717,N_24107,N_24700);
and U25718 (N_25718,N_24770,N_23088);
or U25719 (N_25719,N_22997,N_24819);
nor U25720 (N_25720,N_22674,N_22922);
or U25721 (N_25721,N_22944,N_24211);
or U25722 (N_25722,N_24720,N_22926);
nor U25723 (N_25723,N_23265,N_23292);
and U25724 (N_25724,N_22505,N_24506);
or U25725 (N_25725,N_23124,N_23492);
nor U25726 (N_25726,N_22598,N_24579);
nor U25727 (N_25727,N_24743,N_23173);
or U25728 (N_25728,N_24014,N_24809);
nand U25729 (N_25729,N_24825,N_22818);
and U25730 (N_25730,N_22794,N_24975);
nand U25731 (N_25731,N_23697,N_22615);
and U25732 (N_25732,N_22500,N_22684);
or U25733 (N_25733,N_24541,N_24469);
nand U25734 (N_25734,N_23427,N_23071);
and U25735 (N_25735,N_22544,N_23815);
nand U25736 (N_25736,N_23755,N_24250);
and U25737 (N_25737,N_23672,N_23162);
or U25738 (N_25738,N_23970,N_23782);
nor U25739 (N_25739,N_24711,N_22953);
nor U25740 (N_25740,N_24822,N_24053);
nand U25741 (N_25741,N_24237,N_24862);
or U25742 (N_25742,N_23093,N_23767);
xor U25743 (N_25743,N_24098,N_23864);
and U25744 (N_25744,N_22678,N_22631);
or U25745 (N_25745,N_23480,N_22549);
nor U25746 (N_25746,N_23331,N_24629);
xor U25747 (N_25747,N_24121,N_23325);
nor U25748 (N_25748,N_23171,N_24856);
nor U25749 (N_25749,N_23899,N_24296);
and U25750 (N_25750,N_24077,N_23069);
and U25751 (N_25751,N_23929,N_24406);
and U25752 (N_25752,N_24044,N_23052);
and U25753 (N_25753,N_22581,N_23958);
and U25754 (N_25754,N_22533,N_22923);
or U25755 (N_25755,N_24432,N_24478);
or U25756 (N_25756,N_23661,N_23245);
and U25757 (N_25757,N_23257,N_24774);
nand U25758 (N_25758,N_23724,N_24083);
or U25759 (N_25759,N_22848,N_23821);
nand U25760 (N_25760,N_23389,N_24923);
or U25761 (N_25761,N_23090,N_23956);
nor U25762 (N_25762,N_23410,N_23158);
nand U25763 (N_25763,N_22919,N_22575);
and U25764 (N_25764,N_23774,N_24869);
and U25765 (N_25765,N_24487,N_23630);
and U25766 (N_25766,N_22737,N_24401);
nand U25767 (N_25767,N_22753,N_24677);
or U25768 (N_25768,N_24802,N_23267);
nand U25769 (N_25769,N_22877,N_24534);
nor U25770 (N_25770,N_23220,N_22762);
and U25771 (N_25771,N_24280,N_24595);
or U25772 (N_25772,N_24062,N_24008);
nand U25773 (N_25773,N_24667,N_24503);
nor U25774 (N_25774,N_22968,N_23588);
xor U25775 (N_25775,N_24744,N_22685);
nor U25776 (N_25776,N_23402,N_23616);
xor U25777 (N_25777,N_23237,N_24114);
and U25778 (N_25778,N_24201,N_23932);
nand U25779 (N_25779,N_23387,N_24924);
nor U25780 (N_25780,N_24834,N_24983);
nor U25781 (N_25781,N_24186,N_24785);
or U25782 (N_25782,N_23982,N_24314);
nand U25783 (N_25783,N_24256,N_23623);
and U25784 (N_25784,N_24058,N_23453);
nor U25785 (N_25785,N_23937,N_24247);
nor U25786 (N_25786,N_24226,N_23339);
or U25787 (N_25787,N_24936,N_23156);
or U25788 (N_25788,N_24294,N_23576);
and U25789 (N_25789,N_23021,N_22522);
nor U25790 (N_25790,N_24932,N_24608);
xor U25791 (N_25791,N_23607,N_23298);
or U25792 (N_25792,N_24690,N_23303);
or U25793 (N_25793,N_23866,N_23529);
and U25794 (N_25794,N_22528,N_23203);
and U25795 (N_25795,N_24365,N_24358);
xnor U25796 (N_25796,N_23951,N_23038);
nand U25797 (N_25797,N_22865,N_22732);
and U25798 (N_25798,N_24651,N_23989);
nand U25799 (N_25799,N_23742,N_23345);
and U25800 (N_25800,N_24828,N_23189);
xor U25801 (N_25801,N_24945,N_23594);
nor U25802 (N_25802,N_23460,N_23567);
nand U25803 (N_25803,N_23365,N_24918);
or U25804 (N_25804,N_24806,N_23262);
or U25805 (N_25805,N_22993,N_23263);
nand U25806 (N_25806,N_22698,N_24320);
and U25807 (N_25807,N_23369,N_23204);
and U25808 (N_25808,N_23121,N_23087);
and U25809 (N_25809,N_24095,N_23829);
nand U25810 (N_25810,N_23255,N_23057);
nor U25811 (N_25811,N_22611,N_22795);
nor U25812 (N_25812,N_22727,N_24703);
nor U25813 (N_25813,N_24323,N_23535);
nor U25814 (N_25814,N_23923,N_22908);
nand U25815 (N_25815,N_24545,N_24780);
nor U25816 (N_25816,N_24291,N_24332);
nor U25817 (N_25817,N_23953,N_23284);
or U25818 (N_25818,N_24351,N_23487);
nor U25819 (N_25819,N_23157,N_23839);
nand U25820 (N_25820,N_22852,N_24146);
nand U25821 (N_25821,N_22825,N_23854);
or U25822 (N_25822,N_22532,N_24428);
or U25823 (N_25823,N_23561,N_23877);
nand U25824 (N_25824,N_23827,N_23606);
nor U25825 (N_25825,N_24059,N_23682);
nor U25826 (N_25826,N_24207,N_24465);
nand U25827 (N_25827,N_22591,N_24468);
and U25828 (N_25828,N_23961,N_24668);
nor U25829 (N_25829,N_23196,N_22556);
and U25830 (N_25830,N_22766,N_23098);
nand U25831 (N_25831,N_22854,N_23511);
nor U25832 (N_25832,N_22945,N_23521);
nand U25833 (N_25833,N_24564,N_24997);
and U25834 (N_25834,N_24300,N_22994);
nor U25835 (N_25835,N_23545,N_24993);
or U25836 (N_25836,N_22860,N_24960);
nor U25837 (N_25837,N_24816,N_22600);
or U25838 (N_25838,N_22989,N_23476);
or U25839 (N_25839,N_22913,N_22956);
nor U25840 (N_25840,N_23489,N_23007);
nor U25841 (N_25841,N_24184,N_24969);
nand U25842 (N_25842,N_23382,N_23151);
and U25843 (N_25843,N_24528,N_23150);
or U25844 (N_25844,N_24492,N_24811);
nor U25845 (N_25845,N_22616,N_23850);
nand U25846 (N_25846,N_24073,N_24861);
and U25847 (N_25847,N_24333,N_22992);
nand U25848 (N_25848,N_22842,N_24331);
or U25849 (N_25849,N_24535,N_24554);
and U25850 (N_25850,N_23972,N_23099);
and U25851 (N_25851,N_24308,N_22776);
xor U25852 (N_25852,N_24650,N_23843);
and U25853 (N_25853,N_22839,N_23747);
nand U25854 (N_25854,N_24815,N_24752);
and U25855 (N_25855,N_24710,N_23202);
or U25856 (N_25856,N_22823,N_23072);
nor U25857 (N_25857,N_22733,N_22571);
nand U25858 (N_25858,N_23659,N_24413);
nand U25859 (N_25859,N_22661,N_23246);
nand U25860 (N_25860,N_22507,N_23604);
nand U25861 (N_25861,N_23054,N_24377);
and U25862 (N_25862,N_24987,N_23868);
xnor U25863 (N_25863,N_24951,N_23185);
and U25864 (N_25864,N_24689,N_23296);
nand U25865 (N_25865,N_23875,N_22740);
nor U25866 (N_25866,N_23131,N_24810);
nand U25867 (N_25867,N_22723,N_22619);
or U25868 (N_25868,N_22580,N_22845);
nor U25869 (N_25869,N_23004,N_23437);
nor U25870 (N_25870,N_23164,N_22653);
nor U25871 (N_25871,N_23101,N_22578);
nor U25872 (N_25872,N_24047,N_24026);
xor U25873 (N_25873,N_24394,N_24467);
nand U25874 (N_25874,N_24490,N_24027);
nor U25875 (N_25875,N_24109,N_23577);
and U25876 (N_25876,N_24902,N_22586);
xor U25877 (N_25877,N_24914,N_23861);
and U25878 (N_25878,N_23172,N_23309);
and U25879 (N_25879,N_24076,N_24754);
nor U25880 (N_25880,N_23076,N_23917);
xnor U25881 (N_25881,N_22508,N_23832);
nand U25882 (N_25882,N_22655,N_24270);
and U25883 (N_25883,N_24423,N_24502);
nor U25884 (N_25884,N_22672,N_23241);
and U25885 (N_25885,N_22889,N_23229);
or U25886 (N_25886,N_22536,N_24150);
nor U25887 (N_25887,N_24716,N_24765);
nand U25888 (N_25888,N_23249,N_23983);
xor U25889 (N_25889,N_24875,N_23488);
nand U25890 (N_25890,N_23068,N_23227);
and U25891 (N_25891,N_24414,N_24381);
or U25892 (N_25892,N_24396,N_22783);
xnor U25893 (N_25893,N_24086,N_22597);
xor U25894 (N_25894,N_23042,N_23356);
or U25895 (N_25895,N_22786,N_24663);
xnor U25896 (N_25896,N_24343,N_23440);
or U25897 (N_25897,N_23600,N_22717);
nor U25898 (N_25898,N_24696,N_22884);
or U25899 (N_25899,N_22607,N_24889);
and U25900 (N_25900,N_22676,N_23261);
nor U25901 (N_25901,N_24293,N_24257);
and U25902 (N_25902,N_22784,N_23790);
nor U25903 (N_25903,N_22592,N_24797);
or U25904 (N_25904,N_22925,N_22873);
nor U25905 (N_25905,N_23700,N_24179);
and U25906 (N_25906,N_24218,N_23063);
or U25907 (N_25907,N_23714,N_23154);
nor U25908 (N_25908,N_24324,N_24928);
xnor U25909 (N_25909,N_23609,N_24299);
nor U25910 (N_25910,N_24091,N_24939);
nor U25911 (N_25911,N_24355,N_23299);
and U25912 (N_25912,N_23074,N_24673);
nor U25913 (N_25913,N_22863,N_22758);
and U25914 (N_25914,N_23504,N_24907);
and U25915 (N_25915,N_22960,N_23918);
xnor U25916 (N_25916,N_24691,N_23973);
xor U25917 (N_25917,N_24031,N_23862);
or U25918 (N_25918,N_22832,N_23919);
and U25919 (N_25919,N_22743,N_24297);
or U25920 (N_25920,N_23109,N_24408);
nor U25921 (N_25921,N_22720,N_23741);
nand U25922 (N_25922,N_22777,N_24961);
and U25923 (N_25923,N_23239,N_23134);
xor U25924 (N_25924,N_23240,N_23785);
and U25925 (N_25925,N_23718,N_24771);
nor U25926 (N_25926,N_24362,N_23825);
nand U25927 (N_25927,N_24784,N_23771);
or U25928 (N_25928,N_24522,N_23811);
nor U25929 (N_25929,N_23416,N_23620);
and U25930 (N_25930,N_24445,N_23949);
nor U25931 (N_25931,N_23130,N_24368);
or U25932 (N_25932,N_22538,N_23126);
xor U25933 (N_25933,N_23556,N_22630);
or U25934 (N_25934,N_24453,N_23562);
nor U25935 (N_25935,N_23816,N_22831);
and U25936 (N_25936,N_24944,N_23029);
xnor U25937 (N_25937,N_23933,N_22817);
and U25938 (N_25938,N_23737,N_24206);
or U25939 (N_25939,N_23392,N_22793);
nand U25940 (N_25940,N_24412,N_22512);
and U25941 (N_25941,N_22856,N_23209);
nand U25942 (N_25942,N_24431,N_23458);
and U25943 (N_25943,N_23462,N_24447);
xnor U25944 (N_25944,N_23498,N_23361);
and U25945 (N_25945,N_24666,N_24425);
nand U25946 (N_25946,N_23794,N_22801);
and U25947 (N_25947,N_24514,N_24586);
nor U25948 (N_25948,N_23015,N_22576);
xor U25949 (N_25949,N_24764,N_24620);
nand U25950 (N_25950,N_23228,N_23984);
or U25951 (N_25951,N_22707,N_24733);
or U25952 (N_25952,N_23434,N_24588);
or U25953 (N_25953,N_23775,N_24934);
and U25954 (N_25954,N_24984,N_22633);
nor U25955 (N_25955,N_24402,N_24967);
nand U25956 (N_25956,N_24341,N_22514);
or U25957 (N_25957,N_22527,N_24287);
nand U25958 (N_25958,N_24424,N_23326);
or U25959 (N_25959,N_23139,N_23991);
nand U25960 (N_25960,N_23572,N_23435);
or U25961 (N_25961,N_23242,N_22987);
nor U25962 (N_25962,N_24578,N_23359);
nand U25963 (N_25963,N_22888,N_24383);
nand U25964 (N_25964,N_24488,N_24494);
or U25965 (N_25965,N_22626,N_23719);
and U25966 (N_25966,N_23232,N_23800);
and U25967 (N_25967,N_24328,N_23834);
xor U25968 (N_25968,N_24470,N_23439);
or U25969 (N_25969,N_22906,N_23143);
nor U25970 (N_25970,N_24559,N_24735);
nand U25971 (N_25971,N_22764,N_24074);
nor U25972 (N_25972,N_23666,N_23525);
nand U25973 (N_25973,N_23586,N_24374);
and U25974 (N_25974,N_24306,N_23035);
nor U25975 (N_25975,N_24777,N_24772);
xor U25976 (N_25976,N_23062,N_23270);
nor U25977 (N_25977,N_22646,N_24221);
xnor U25978 (N_25978,N_24230,N_23036);
xor U25979 (N_25979,N_24348,N_22550);
or U25980 (N_25980,N_23399,N_23000);
nor U25981 (N_25981,N_24248,N_23293);
or U25982 (N_25982,N_23360,N_23818);
nand U25983 (N_25983,N_24193,N_24916);
and U25984 (N_25984,N_22531,N_23423);
nand U25985 (N_25985,N_23335,N_23967);
nand U25986 (N_25986,N_23422,N_22694);
and U25987 (N_25987,N_23756,N_23589);
xnor U25988 (N_25988,N_23112,N_24879);
xor U25989 (N_25989,N_22620,N_23353);
xnor U25990 (N_25990,N_23327,N_23632);
or U25991 (N_25991,N_23645,N_24400);
nor U25992 (N_25992,N_24215,N_24088);
nor U25993 (N_25993,N_24567,N_24289);
and U25994 (N_25994,N_24450,N_24865);
or U25995 (N_25995,N_23880,N_24724);
xnor U25996 (N_25996,N_23571,N_24679);
and U25997 (N_25997,N_23483,N_24199);
nand U25998 (N_25998,N_24585,N_24714);
nand U25999 (N_25999,N_24839,N_23962);
and U26000 (N_26000,N_22613,N_24103);
nand U26001 (N_26001,N_24930,N_24893);
and U26002 (N_26002,N_23524,N_22952);
nor U26003 (N_26003,N_24739,N_23163);
and U26004 (N_26004,N_24558,N_24715);
nor U26005 (N_26005,N_23580,N_23102);
and U26006 (N_26006,N_23906,N_22504);
or U26007 (N_26007,N_23647,N_23903);
nand U26008 (N_26008,N_24519,N_22711);
and U26009 (N_26009,N_23319,N_23597);
nand U26010 (N_26010,N_22572,N_23135);
and U26011 (N_26011,N_24747,N_23696);
or U26012 (N_26012,N_23617,N_24090);
or U26013 (N_26013,N_24794,N_22594);
nand U26014 (N_26014,N_24805,N_23945);
and U26015 (N_26015,N_23629,N_24459);
or U26016 (N_26016,N_24854,N_24446);
nor U26017 (N_26017,N_24561,N_23385);
nand U26018 (N_26018,N_23925,N_24181);
nor U26019 (N_26019,N_23461,N_22941);
and U26020 (N_26020,N_24336,N_22816);
nor U26021 (N_26021,N_24979,N_22559);
nor U26022 (N_26022,N_23140,N_24762);
nand U26023 (N_26023,N_24542,N_24982);
and U26024 (N_26024,N_24312,N_22797);
and U26025 (N_26025,N_24636,N_22808);
xnor U26026 (N_26026,N_23301,N_24905);
and U26027 (N_26027,N_23555,N_23505);
and U26028 (N_26028,N_24919,N_23106);
and U26029 (N_26029,N_22665,N_23201);
or U26030 (N_26030,N_24386,N_24966);
xor U26031 (N_26031,N_24791,N_24142);
nand U26032 (N_26032,N_24126,N_24886);
xnor U26033 (N_26033,N_23012,N_22984);
nand U26034 (N_26034,N_24883,N_23996);
nand U26035 (N_26035,N_24203,N_23200);
and U26036 (N_26036,N_23321,N_23520);
or U26037 (N_26037,N_24638,N_24681);
xnor U26038 (N_26038,N_24133,N_22697);
nor U26039 (N_26039,N_22604,N_23514);
or U26040 (N_26040,N_24172,N_24781);
and U26041 (N_26041,N_23133,N_24210);
nand U26042 (N_26042,N_23542,N_23793);
or U26043 (N_26043,N_24683,N_22995);
and U26044 (N_26044,N_23726,N_24999);
nand U26045 (N_26045,N_23451,N_24981);
xnor U26046 (N_26046,N_24623,N_23650);
and U26047 (N_26047,N_22900,N_22638);
nor U26048 (N_26048,N_22911,N_23581);
nand U26049 (N_26049,N_23960,N_24147);
and U26050 (N_26050,N_23501,N_23731);
or U26051 (N_26051,N_24551,N_24676);
or U26052 (N_26052,N_23713,N_23448);
xnor U26053 (N_26053,N_24500,N_24304);
xor U26054 (N_26054,N_23707,N_24704);
or U26055 (N_26055,N_24489,N_23221);
nor U26056 (N_26056,N_24686,N_23349);
or U26057 (N_26057,N_24264,N_23725);
and U26058 (N_26058,N_23411,N_24592);
nor U26059 (N_26059,N_23518,N_24065);
nor U26060 (N_26060,N_22511,N_23665);
xor U26061 (N_26061,N_23391,N_22614);
nor U26062 (N_26062,N_22929,N_22516);
and U26063 (N_26063,N_23433,N_24523);
nor U26064 (N_26064,N_22756,N_23585);
and U26065 (N_26065,N_24630,N_24527);
and U26066 (N_26066,N_23179,N_23244);
nor U26067 (N_26067,N_24222,N_23537);
and U26068 (N_26068,N_24345,N_22826);
nor U26069 (N_26069,N_24143,N_22940);
or U26070 (N_26070,N_23082,N_22807);
or U26071 (N_26071,N_23277,N_24560);
or U26072 (N_26072,N_24948,N_23976);
and U26073 (N_26073,N_24048,N_24894);
nand U26074 (N_26074,N_23187,N_24601);
or U26075 (N_26075,N_23654,N_24067);
nor U26076 (N_26076,N_23809,N_24974);
and U26077 (N_26077,N_23587,N_24874);
or U26078 (N_26078,N_23271,N_24552);
nor U26079 (N_26079,N_22564,N_23357);
and U26080 (N_26080,N_23867,N_22980);
xnor U26081 (N_26081,N_23559,N_23050);
nand U26082 (N_26082,N_23067,N_24238);
nor U26083 (N_26083,N_22567,N_23736);
nor U26084 (N_26084,N_24497,N_24680);
nand U26085 (N_26085,N_24800,N_24857);
and U26086 (N_26086,N_24619,N_22590);
xor U26087 (N_26087,N_23047,N_24302);
nand U26088 (N_26088,N_23997,N_22898);
and U26089 (N_26089,N_23749,N_23238);
or U26090 (N_26090,N_24149,N_24725);
and U26091 (N_26091,N_24192,N_23253);
and U26092 (N_26092,N_24779,N_24004);
or U26093 (N_26093,N_24069,N_23930);
nor U26094 (N_26094,N_22866,N_24732);
nor U26095 (N_26095,N_23798,N_24005);
nand U26096 (N_26096,N_22623,N_23046);
nor U26097 (N_26097,N_24278,N_24458);
xnor U26098 (N_26098,N_24581,N_22725);
and U26099 (N_26099,N_23471,N_24158);
nor U26100 (N_26100,N_23280,N_23624);
nor U26101 (N_26101,N_23683,N_24444);
and U26102 (N_26102,N_24482,N_23281);
or U26103 (N_26103,N_22687,N_23992);
nand U26104 (N_26104,N_24023,N_23915);
xnor U26105 (N_26105,N_22798,N_24639);
nor U26106 (N_26106,N_23444,N_23676);
xnor U26107 (N_26107,N_24895,N_23722);
or U26108 (N_26108,N_22657,N_24829);
and U26109 (N_26109,N_23375,N_22920);
nand U26110 (N_26110,N_23920,N_24543);
nand U26111 (N_26111,N_24219,N_23222);
and U26112 (N_26112,N_23692,N_22876);
or U26113 (N_26113,N_22867,N_23031);
xor U26114 (N_26114,N_24366,N_23214);
nand U26115 (N_26115,N_22692,N_23999);
and U26116 (N_26116,N_24904,N_23500);
xnor U26117 (N_26117,N_23454,N_23823);
nand U26118 (N_26118,N_24099,N_23128);
nand U26119 (N_26119,N_24622,N_24395);
nor U26120 (N_26120,N_22921,N_24182);
nand U26121 (N_26121,N_24389,N_23759);
or U26122 (N_26122,N_24778,N_22714);
or U26123 (N_26123,N_23651,N_23698);
nor U26124 (N_26124,N_22636,N_24357);
nor U26125 (N_26125,N_24705,N_24448);
xor U26126 (N_26126,N_23757,N_23596);
and U26127 (N_26127,N_24421,N_24159);
and U26128 (N_26128,N_23564,N_24155);
nor U26129 (N_26129,N_24418,N_23111);
nor U26130 (N_26130,N_24021,N_23490);
nor U26131 (N_26131,N_23073,N_22699);
or U26132 (N_26132,N_23541,N_24194);
nand U26133 (N_26133,N_24352,N_22855);
and U26134 (N_26134,N_23730,N_23077);
and U26135 (N_26135,N_24517,N_24170);
nand U26136 (N_26136,N_24134,N_24057);
nand U26137 (N_26137,N_23314,N_24831);
nor U26138 (N_26138,N_24409,N_24177);
xor U26139 (N_26139,N_24833,N_23789);
or U26140 (N_26140,N_24156,N_22781);
nor U26141 (N_26141,N_22689,N_24644);
and U26142 (N_26142,N_24538,N_23145);
and U26143 (N_26143,N_24962,N_22526);
and U26144 (N_26144,N_24990,N_23797);
nor U26145 (N_26145,N_23664,N_24906);
nand U26146 (N_26146,N_23583,N_24611);
nand U26147 (N_26147,N_23639,N_22742);
nor U26148 (N_26148,N_23530,N_23605);
and U26149 (N_26149,N_24576,N_24610);
xnor U26150 (N_26150,N_24640,N_24115);
nand U26151 (N_26151,N_23276,N_23538);
or U26152 (N_26152,N_24892,N_24160);
xnor U26153 (N_26153,N_23400,N_23830);
and U26154 (N_26154,N_23565,N_23463);
nor U26155 (N_26155,N_23863,N_23198);
and U26156 (N_26156,N_24346,N_23849);
nor U26157 (N_26157,N_23675,N_24881);
nand U26158 (N_26158,N_24937,N_24479);
and U26159 (N_26159,N_23176,N_24540);
nor U26160 (N_26160,N_23858,N_22815);
nand U26161 (N_26161,N_24872,N_23457);
nor U26162 (N_26162,N_22903,N_23260);
or U26163 (N_26163,N_23328,N_22931);
or U26164 (N_26164,N_24042,N_24501);
and U26165 (N_26165,N_24118,N_23805);
and U26166 (N_26166,N_22730,N_23552);
or U26167 (N_26167,N_24970,N_24821);
nor U26168 (N_26168,N_23003,N_23888);
nor U26169 (N_26169,N_24963,N_23870);
or U26170 (N_26170,N_23499,N_23590);
or U26171 (N_26171,N_23110,N_23729);
nor U26172 (N_26172,N_24010,N_22705);
nand U26173 (N_26173,N_22976,N_23317);
or U26174 (N_26174,N_23810,N_24191);
xor U26175 (N_26175,N_23687,N_23881);
or U26176 (N_26176,N_23612,N_24055);
nand U26177 (N_26177,N_23926,N_24174);
or U26178 (N_26178,N_24430,N_23405);
or U26179 (N_26179,N_23509,N_23170);
nor U26180 (N_26180,N_23132,N_24717);
nor U26181 (N_26181,N_23105,N_23092);
or U26182 (N_26182,N_22744,N_23123);
nand U26183 (N_26183,N_24056,N_22521);
xnor U26184 (N_26184,N_24451,N_23381);
and U26185 (N_26185,N_24697,N_23635);
nor U26186 (N_26186,N_24653,N_22510);
and U26187 (N_26187,N_24315,N_22772);
and U26188 (N_26188,N_23180,N_23910);
and U26189 (N_26189,N_23611,N_23595);
nand U26190 (N_26190,N_24072,N_23218);
nand U26191 (N_26191,N_23987,N_22569);
nand U26192 (N_26192,N_22669,N_23343);
xnor U26193 (N_26193,N_24195,N_23546);
xnor U26194 (N_26194,N_24189,N_23773);
nand U26195 (N_26195,N_23515,N_23060);
nand U26196 (N_26196,N_24123,N_23347);
and U26197 (N_26197,N_23708,N_23496);
or U26198 (N_26198,N_23952,N_23684);
nor U26199 (N_26199,N_24309,N_24525);
nor U26200 (N_26200,N_22990,N_22970);
xnor U26201 (N_26201,N_24397,N_24789);
and U26202 (N_26202,N_24574,N_24731);
and U26203 (N_26203,N_22850,N_24671);
or U26204 (N_26204,N_23033,N_23386);
or U26205 (N_26205,N_23554,N_23655);
nor U26206 (N_26206,N_24953,N_22746);
and U26207 (N_26207,N_23393,N_24017);
and U26208 (N_26208,N_22896,N_23634);
or U26209 (N_26209,N_24419,N_23975);
nor U26210 (N_26210,N_23638,N_23944);
and U26211 (N_26211,N_22752,N_23549);
nor U26212 (N_26212,N_22893,N_24996);
or U26213 (N_26213,N_24726,N_23289);
nor U26214 (N_26214,N_24550,N_23113);
xor U26215 (N_26215,N_23030,N_24119);
and U26216 (N_26216,N_22827,N_22824);
and U26217 (N_26217,N_24909,N_22780);
or U26218 (N_26218,N_24604,N_24590);
and U26219 (N_26219,N_22977,N_22651);
nor U26220 (N_26220,N_22790,N_24980);
nand U26221 (N_26221,N_24387,N_23762);
nor U26222 (N_26222,N_24580,N_24475);
xnor U26223 (N_26223,N_22836,N_24367);
nor U26224 (N_26224,N_22566,N_23788);
nor U26225 (N_26225,N_23051,N_23486);
nand U26226 (N_26226,N_23660,N_24267);
nand U26227 (N_26227,N_22803,N_23691);
nand U26228 (N_26228,N_23136,N_23230);
or U26229 (N_26229,N_22683,N_22768);
or U26230 (N_26230,N_22605,N_24274);
nand U26231 (N_26231,N_23935,N_24701);
nor U26232 (N_26232,N_23739,N_24285);
nor U26233 (N_26233,N_22647,N_24853);
and U26234 (N_26234,N_22524,N_22509);
or U26235 (N_26235,N_24840,N_23273);
or U26236 (N_26236,N_23125,N_24940);
or U26237 (N_26237,N_24607,N_24533);
and U26238 (N_26238,N_24694,N_23904);
nor U26239 (N_26239,N_23540,N_24769);
nor U26240 (N_26240,N_24582,N_23601);
or U26241 (N_26241,N_23653,N_22627);
or U26242 (N_26242,N_24841,N_24885);
nor U26243 (N_26243,N_22838,N_23342);
or U26244 (N_26244,N_23181,N_23120);
xnor U26245 (N_26245,N_22949,N_23159);
nand U26246 (N_26246,N_24884,N_23802);
or U26247 (N_26247,N_24003,N_24132);
or U26248 (N_26248,N_22930,N_23302);
xnor U26249 (N_26249,N_24842,N_24231);
and U26250 (N_26250,N_23688,N_22990);
nand U26251 (N_26251,N_23124,N_23070);
xnor U26252 (N_26252,N_23478,N_24131);
xor U26253 (N_26253,N_23073,N_22618);
nand U26254 (N_26254,N_24089,N_23950);
nor U26255 (N_26255,N_22960,N_24488);
xnor U26256 (N_26256,N_23765,N_24796);
nor U26257 (N_26257,N_24762,N_23006);
and U26258 (N_26258,N_24480,N_24309);
nand U26259 (N_26259,N_24811,N_23271);
or U26260 (N_26260,N_23729,N_23454);
or U26261 (N_26261,N_24441,N_23500);
and U26262 (N_26262,N_23826,N_24065);
or U26263 (N_26263,N_23420,N_23179);
or U26264 (N_26264,N_22640,N_24521);
and U26265 (N_26265,N_23923,N_24620);
nand U26266 (N_26266,N_24828,N_23097);
nand U26267 (N_26267,N_22751,N_22692);
or U26268 (N_26268,N_22946,N_24267);
and U26269 (N_26269,N_24834,N_24114);
or U26270 (N_26270,N_24096,N_23374);
and U26271 (N_26271,N_23584,N_23390);
and U26272 (N_26272,N_24128,N_24353);
nor U26273 (N_26273,N_23524,N_22756);
nor U26274 (N_26274,N_23705,N_24463);
nor U26275 (N_26275,N_23581,N_24581);
nand U26276 (N_26276,N_22922,N_22576);
nor U26277 (N_26277,N_24210,N_22846);
nor U26278 (N_26278,N_24965,N_23869);
or U26279 (N_26279,N_24170,N_23531);
nor U26280 (N_26280,N_24271,N_24719);
or U26281 (N_26281,N_24001,N_24899);
nand U26282 (N_26282,N_24894,N_24297);
nand U26283 (N_26283,N_23061,N_24139);
and U26284 (N_26284,N_23063,N_24906);
nor U26285 (N_26285,N_24320,N_24166);
nor U26286 (N_26286,N_23177,N_22823);
nand U26287 (N_26287,N_24892,N_24345);
nor U26288 (N_26288,N_23535,N_24085);
or U26289 (N_26289,N_22536,N_24793);
xor U26290 (N_26290,N_24504,N_24164);
nand U26291 (N_26291,N_24645,N_23702);
nand U26292 (N_26292,N_23444,N_24804);
and U26293 (N_26293,N_24634,N_23313);
or U26294 (N_26294,N_23585,N_22945);
xor U26295 (N_26295,N_23357,N_24193);
nand U26296 (N_26296,N_24609,N_22673);
nand U26297 (N_26297,N_24685,N_24185);
and U26298 (N_26298,N_24521,N_22989);
and U26299 (N_26299,N_23655,N_24346);
nand U26300 (N_26300,N_24641,N_24156);
nor U26301 (N_26301,N_24002,N_24058);
and U26302 (N_26302,N_23453,N_24757);
and U26303 (N_26303,N_23763,N_24694);
xnor U26304 (N_26304,N_23663,N_23999);
nand U26305 (N_26305,N_24624,N_24571);
or U26306 (N_26306,N_24076,N_23356);
nor U26307 (N_26307,N_23035,N_22928);
or U26308 (N_26308,N_23913,N_23686);
or U26309 (N_26309,N_22771,N_23014);
nand U26310 (N_26310,N_23222,N_23959);
xnor U26311 (N_26311,N_23742,N_24029);
nor U26312 (N_26312,N_23825,N_23642);
xor U26313 (N_26313,N_22956,N_23617);
or U26314 (N_26314,N_23938,N_23473);
and U26315 (N_26315,N_22851,N_24132);
nor U26316 (N_26316,N_24102,N_24440);
and U26317 (N_26317,N_24487,N_24017);
and U26318 (N_26318,N_23937,N_22784);
nand U26319 (N_26319,N_22789,N_23709);
nor U26320 (N_26320,N_24969,N_24690);
nor U26321 (N_26321,N_23910,N_24846);
and U26322 (N_26322,N_24240,N_23332);
nand U26323 (N_26323,N_24261,N_23988);
and U26324 (N_26324,N_23945,N_24335);
and U26325 (N_26325,N_23894,N_22842);
nand U26326 (N_26326,N_22806,N_22900);
nor U26327 (N_26327,N_23635,N_22629);
or U26328 (N_26328,N_23995,N_23723);
or U26329 (N_26329,N_23159,N_22681);
xor U26330 (N_26330,N_22701,N_24200);
or U26331 (N_26331,N_24374,N_24268);
nand U26332 (N_26332,N_23496,N_22783);
nor U26333 (N_26333,N_23935,N_24375);
and U26334 (N_26334,N_22579,N_22898);
and U26335 (N_26335,N_24763,N_22671);
nand U26336 (N_26336,N_24464,N_24328);
and U26337 (N_26337,N_22509,N_23102);
nor U26338 (N_26338,N_24093,N_24076);
nand U26339 (N_26339,N_24477,N_24027);
nor U26340 (N_26340,N_23648,N_24220);
nor U26341 (N_26341,N_22853,N_23546);
nand U26342 (N_26342,N_23435,N_23108);
nand U26343 (N_26343,N_23529,N_22748);
or U26344 (N_26344,N_23359,N_22750);
nor U26345 (N_26345,N_23278,N_24464);
nand U26346 (N_26346,N_24647,N_24048);
xor U26347 (N_26347,N_23777,N_24743);
xnor U26348 (N_26348,N_22850,N_24059);
and U26349 (N_26349,N_22630,N_23651);
and U26350 (N_26350,N_24956,N_24290);
or U26351 (N_26351,N_23050,N_22804);
or U26352 (N_26352,N_24032,N_23312);
or U26353 (N_26353,N_23569,N_23346);
or U26354 (N_26354,N_23828,N_23097);
and U26355 (N_26355,N_23769,N_24119);
nand U26356 (N_26356,N_22930,N_24454);
or U26357 (N_26357,N_24749,N_24371);
and U26358 (N_26358,N_24839,N_23979);
and U26359 (N_26359,N_24792,N_23204);
and U26360 (N_26360,N_23368,N_24902);
and U26361 (N_26361,N_22893,N_23328);
nand U26362 (N_26362,N_23197,N_23774);
nand U26363 (N_26363,N_23694,N_22894);
xnor U26364 (N_26364,N_24659,N_24306);
and U26365 (N_26365,N_23109,N_23706);
xnor U26366 (N_26366,N_23040,N_24051);
nand U26367 (N_26367,N_24859,N_22737);
and U26368 (N_26368,N_24739,N_24305);
and U26369 (N_26369,N_23568,N_23858);
nor U26370 (N_26370,N_23093,N_24844);
and U26371 (N_26371,N_24478,N_22508);
nor U26372 (N_26372,N_24620,N_22661);
or U26373 (N_26373,N_24834,N_22683);
and U26374 (N_26374,N_23504,N_24913);
xnor U26375 (N_26375,N_24098,N_24872);
nand U26376 (N_26376,N_22667,N_23684);
nand U26377 (N_26377,N_23071,N_23352);
nand U26378 (N_26378,N_23503,N_24915);
or U26379 (N_26379,N_22652,N_24728);
or U26380 (N_26380,N_24550,N_22758);
xnor U26381 (N_26381,N_22997,N_23161);
nand U26382 (N_26382,N_23161,N_23369);
nand U26383 (N_26383,N_24930,N_24085);
nor U26384 (N_26384,N_22559,N_24997);
nor U26385 (N_26385,N_22609,N_23806);
nor U26386 (N_26386,N_23645,N_23047);
xor U26387 (N_26387,N_24116,N_24832);
nand U26388 (N_26388,N_24108,N_23436);
nor U26389 (N_26389,N_24052,N_23595);
nor U26390 (N_26390,N_24351,N_23843);
nand U26391 (N_26391,N_23823,N_24186);
nor U26392 (N_26392,N_23653,N_24732);
and U26393 (N_26393,N_23326,N_24451);
or U26394 (N_26394,N_23008,N_24440);
nand U26395 (N_26395,N_24344,N_23210);
and U26396 (N_26396,N_23119,N_22858);
nand U26397 (N_26397,N_23760,N_24592);
and U26398 (N_26398,N_24933,N_24557);
and U26399 (N_26399,N_22606,N_23086);
xnor U26400 (N_26400,N_24883,N_23192);
or U26401 (N_26401,N_23173,N_22674);
nor U26402 (N_26402,N_23575,N_23793);
or U26403 (N_26403,N_23628,N_24849);
or U26404 (N_26404,N_24974,N_22598);
xnor U26405 (N_26405,N_24932,N_24584);
or U26406 (N_26406,N_22792,N_22796);
or U26407 (N_26407,N_23622,N_24220);
nand U26408 (N_26408,N_24907,N_22853);
nand U26409 (N_26409,N_24439,N_23481);
or U26410 (N_26410,N_23062,N_22556);
and U26411 (N_26411,N_23862,N_23980);
xor U26412 (N_26412,N_24334,N_23069);
and U26413 (N_26413,N_23030,N_23070);
and U26414 (N_26414,N_24588,N_24741);
and U26415 (N_26415,N_22754,N_23349);
and U26416 (N_26416,N_24548,N_22946);
nor U26417 (N_26417,N_23460,N_22754);
nor U26418 (N_26418,N_24860,N_22728);
xor U26419 (N_26419,N_23723,N_24598);
or U26420 (N_26420,N_24417,N_23981);
nand U26421 (N_26421,N_22755,N_24662);
xor U26422 (N_26422,N_24955,N_24583);
and U26423 (N_26423,N_22629,N_24029);
or U26424 (N_26424,N_23300,N_23431);
and U26425 (N_26425,N_24911,N_23939);
nand U26426 (N_26426,N_23741,N_24142);
nand U26427 (N_26427,N_24396,N_22815);
nand U26428 (N_26428,N_24994,N_23950);
nor U26429 (N_26429,N_24889,N_23477);
and U26430 (N_26430,N_23370,N_23900);
or U26431 (N_26431,N_23220,N_24488);
nand U26432 (N_26432,N_24039,N_24645);
xnor U26433 (N_26433,N_23919,N_22651);
nor U26434 (N_26434,N_23043,N_22907);
nand U26435 (N_26435,N_23229,N_22959);
xnor U26436 (N_26436,N_24891,N_23770);
and U26437 (N_26437,N_23457,N_23140);
or U26438 (N_26438,N_23511,N_22546);
nand U26439 (N_26439,N_23339,N_24522);
nand U26440 (N_26440,N_23792,N_22575);
xnor U26441 (N_26441,N_22978,N_24868);
nor U26442 (N_26442,N_24281,N_24366);
nand U26443 (N_26443,N_24647,N_22997);
nor U26444 (N_26444,N_23541,N_23768);
and U26445 (N_26445,N_23654,N_23753);
xor U26446 (N_26446,N_23896,N_23937);
nor U26447 (N_26447,N_22512,N_22569);
and U26448 (N_26448,N_24293,N_23377);
nor U26449 (N_26449,N_23076,N_23483);
nor U26450 (N_26450,N_24731,N_24036);
or U26451 (N_26451,N_23833,N_23515);
xnor U26452 (N_26452,N_23526,N_24429);
nand U26453 (N_26453,N_23312,N_24659);
or U26454 (N_26454,N_24353,N_24627);
nor U26455 (N_26455,N_24621,N_23372);
or U26456 (N_26456,N_23206,N_24174);
or U26457 (N_26457,N_23332,N_23228);
xor U26458 (N_26458,N_24284,N_22757);
xnor U26459 (N_26459,N_24357,N_23188);
nor U26460 (N_26460,N_24737,N_23443);
nor U26461 (N_26461,N_24096,N_23733);
or U26462 (N_26462,N_24403,N_24723);
and U26463 (N_26463,N_23473,N_23073);
nand U26464 (N_26464,N_24098,N_22951);
or U26465 (N_26465,N_23877,N_24665);
and U26466 (N_26466,N_24097,N_24092);
or U26467 (N_26467,N_23464,N_23401);
or U26468 (N_26468,N_23442,N_24641);
nor U26469 (N_26469,N_22757,N_22606);
nand U26470 (N_26470,N_24625,N_23678);
nand U26471 (N_26471,N_24440,N_23699);
nor U26472 (N_26472,N_22630,N_23207);
nand U26473 (N_26473,N_24022,N_24351);
or U26474 (N_26474,N_23641,N_24238);
nor U26475 (N_26475,N_24558,N_23898);
nor U26476 (N_26476,N_23645,N_23723);
and U26477 (N_26477,N_22707,N_23852);
nor U26478 (N_26478,N_23506,N_24129);
nand U26479 (N_26479,N_23080,N_24719);
nor U26480 (N_26480,N_24800,N_23224);
or U26481 (N_26481,N_23104,N_22846);
or U26482 (N_26482,N_22917,N_24213);
nand U26483 (N_26483,N_23644,N_24451);
nor U26484 (N_26484,N_24856,N_23497);
or U26485 (N_26485,N_23749,N_24928);
nand U26486 (N_26486,N_24159,N_24962);
and U26487 (N_26487,N_22653,N_24246);
or U26488 (N_26488,N_23487,N_24421);
and U26489 (N_26489,N_23307,N_24800);
and U26490 (N_26490,N_23826,N_23995);
or U26491 (N_26491,N_24350,N_24396);
or U26492 (N_26492,N_24441,N_23138);
nor U26493 (N_26493,N_24478,N_24991);
nor U26494 (N_26494,N_23024,N_24854);
or U26495 (N_26495,N_24998,N_22741);
and U26496 (N_26496,N_22629,N_22627);
xnor U26497 (N_26497,N_22861,N_22579);
nor U26498 (N_26498,N_23854,N_24079);
or U26499 (N_26499,N_24694,N_24277);
or U26500 (N_26500,N_22819,N_24640);
and U26501 (N_26501,N_24881,N_23647);
nand U26502 (N_26502,N_23957,N_23899);
or U26503 (N_26503,N_24290,N_24378);
xor U26504 (N_26504,N_24291,N_23672);
nor U26505 (N_26505,N_23394,N_23393);
or U26506 (N_26506,N_23908,N_24908);
nand U26507 (N_26507,N_22858,N_23926);
nor U26508 (N_26508,N_24997,N_23952);
nand U26509 (N_26509,N_23471,N_22885);
and U26510 (N_26510,N_24563,N_23124);
or U26511 (N_26511,N_24610,N_23209);
nand U26512 (N_26512,N_23026,N_24505);
nor U26513 (N_26513,N_22887,N_24076);
nand U26514 (N_26514,N_24607,N_22945);
xor U26515 (N_26515,N_23332,N_23909);
nor U26516 (N_26516,N_22899,N_24446);
and U26517 (N_26517,N_24814,N_24119);
nand U26518 (N_26518,N_23788,N_24696);
nand U26519 (N_26519,N_22886,N_23855);
nor U26520 (N_26520,N_22620,N_23575);
and U26521 (N_26521,N_22527,N_23844);
or U26522 (N_26522,N_23265,N_24532);
nor U26523 (N_26523,N_23606,N_23430);
nand U26524 (N_26524,N_24928,N_24348);
and U26525 (N_26525,N_22862,N_23878);
and U26526 (N_26526,N_23372,N_24799);
or U26527 (N_26527,N_22681,N_23117);
and U26528 (N_26528,N_22868,N_22982);
xor U26529 (N_26529,N_23693,N_24769);
or U26530 (N_26530,N_24011,N_23149);
or U26531 (N_26531,N_24053,N_23991);
nor U26532 (N_26532,N_24012,N_24617);
nor U26533 (N_26533,N_24289,N_22740);
nand U26534 (N_26534,N_22752,N_24694);
nor U26535 (N_26535,N_24160,N_22980);
and U26536 (N_26536,N_23037,N_24261);
or U26537 (N_26537,N_24213,N_23203);
or U26538 (N_26538,N_24972,N_24740);
nand U26539 (N_26539,N_23521,N_24669);
nor U26540 (N_26540,N_24233,N_22817);
or U26541 (N_26541,N_24941,N_23849);
or U26542 (N_26542,N_24795,N_22574);
or U26543 (N_26543,N_24048,N_23437);
or U26544 (N_26544,N_23144,N_24123);
nand U26545 (N_26545,N_24348,N_23892);
nand U26546 (N_26546,N_22556,N_22991);
and U26547 (N_26547,N_24375,N_23751);
or U26548 (N_26548,N_23035,N_24328);
or U26549 (N_26549,N_23481,N_24839);
xor U26550 (N_26550,N_24892,N_23754);
or U26551 (N_26551,N_24000,N_24076);
xnor U26552 (N_26552,N_23185,N_23371);
or U26553 (N_26553,N_24107,N_23365);
xnor U26554 (N_26554,N_22973,N_24244);
nand U26555 (N_26555,N_23632,N_23206);
and U26556 (N_26556,N_23444,N_24997);
or U26557 (N_26557,N_24260,N_23544);
or U26558 (N_26558,N_22611,N_23519);
nor U26559 (N_26559,N_23410,N_24887);
xnor U26560 (N_26560,N_22700,N_22671);
nor U26561 (N_26561,N_24287,N_24610);
nand U26562 (N_26562,N_24608,N_22757);
nor U26563 (N_26563,N_22617,N_22699);
xnor U26564 (N_26564,N_23743,N_24610);
and U26565 (N_26565,N_24270,N_23123);
xnor U26566 (N_26566,N_23997,N_23869);
nor U26567 (N_26567,N_22884,N_23010);
or U26568 (N_26568,N_23221,N_22736);
nand U26569 (N_26569,N_23824,N_23978);
or U26570 (N_26570,N_22532,N_23859);
xnor U26571 (N_26571,N_24422,N_24640);
xnor U26572 (N_26572,N_22603,N_24770);
nor U26573 (N_26573,N_24711,N_24182);
nand U26574 (N_26574,N_23933,N_23755);
and U26575 (N_26575,N_22693,N_22986);
nor U26576 (N_26576,N_24177,N_23327);
nand U26577 (N_26577,N_24119,N_23434);
nor U26578 (N_26578,N_22974,N_22526);
xor U26579 (N_26579,N_24474,N_23548);
or U26580 (N_26580,N_23164,N_24467);
and U26581 (N_26581,N_22643,N_23101);
xnor U26582 (N_26582,N_22780,N_23679);
xor U26583 (N_26583,N_22713,N_23042);
nor U26584 (N_26584,N_24463,N_24083);
nand U26585 (N_26585,N_23010,N_22787);
nor U26586 (N_26586,N_24291,N_23525);
xor U26587 (N_26587,N_24060,N_23126);
nand U26588 (N_26588,N_24114,N_23419);
and U26589 (N_26589,N_23211,N_24277);
xnor U26590 (N_26590,N_24533,N_23145);
or U26591 (N_26591,N_23574,N_24153);
and U26592 (N_26592,N_22805,N_22641);
or U26593 (N_26593,N_24550,N_23768);
and U26594 (N_26594,N_24701,N_24873);
and U26595 (N_26595,N_24714,N_23025);
nor U26596 (N_26596,N_22819,N_22707);
nor U26597 (N_26597,N_22549,N_24190);
xnor U26598 (N_26598,N_24139,N_22871);
xor U26599 (N_26599,N_23149,N_24120);
and U26600 (N_26600,N_23832,N_22929);
and U26601 (N_26601,N_24229,N_24776);
nand U26602 (N_26602,N_24933,N_24190);
or U26603 (N_26603,N_22683,N_24020);
and U26604 (N_26604,N_23069,N_24572);
nor U26605 (N_26605,N_24268,N_24814);
nor U26606 (N_26606,N_23415,N_24256);
xor U26607 (N_26607,N_23275,N_23534);
or U26608 (N_26608,N_24410,N_23571);
nor U26609 (N_26609,N_23768,N_24724);
and U26610 (N_26610,N_22532,N_23667);
nand U26611 (N_26611,N_23734,N_24529);
and U26612 (N_26612,N_22660,N_24910);
or U26613 (N_26613,N_23490,N_23058);
nor U26614 (N_26614,N_24133,N_22961);
or U26615 (N_26615,N_22887,N_23770);
and U26616 (N_26616,N_24338,N_23928);
or U26617 (N_26617,N_23149,N_24012);
or U26618 (N_26618,N_23561,N_23850);
nor U26619 (N_26619,N_23064,N_24139);
nand U26620 (N_26620,N_24706,N_24400);
nor U26621 (N_26621,N_24961,N_24411);
and U26622 (N_26622,N_22740,N_23410);
nor U26623 (N_26623,N_23395,N_24328);
and U26624 (N_26624,N_24778,N_23687);
nor U26625 (N_26625,N_24663,N_24135);
nand U26626 (N_26626,N_24959,N_23870);
or U26627 (N_26627,N_23131,N_24019);
and U26628 (N_26628,N_23771,N_24062);
nor U26629 (N_26629,N_24098,N_24532);
nand U26630 (N_26630,N_22819,N_23086);
nand U26631 (N_26631,N_24886,N_23518);
nor U26632 (N_26632,N_23064,N_24650);
and U26633 (N_26633,N_24213,N_23556);
nand U26634 (N_26634,N_24684,N_22975);
or U26635 (N_26635,N_22506,N_23074);
xor U26636 (N_26636,N_22797,N_22882);
nand U26637 (N_26637,N_23922,N_24013);
nand U26638 (N_26638,N_23992,N_22962);
nor U26639 (N_26639,N_22771,N_22879);
nand U26640 (N_26640,N_24297,N_23963);
xor U26641 (N_26641,N_23926,N_23067);
or U26642 (N_26642,N_22981,N_23172);
nand U26643 (N_26643,N_24958,N_22642);
xor U26644 (N_26644,N_23565,N_23802);
nand U26645 (N_26645,N_22675,N_22514);
or U26646 (N_26646,N_24522,N_24009);
nand U26647 (N_26647,N_22543,N_23501);
nor U26648 (N_26648,N_24705,N_23406);
nor U26649 (N_26649,N_24294,N_23705);
or U26650 (N_26650,N_24620,N_23822);
nand U26651 (N_26651,N_24961,N_24113);
nand U26652 (N_26652,N_24448,N_24594);
nand U26653 (N_26653,N_23827,N_23359);
and U26654 (N_26654,N_23553,N_22631);
and U26655 (N_26655,N_24372,N_24595);
or U26656 (N_26656,N_23165,N_22523);
nand U26657 (N_26657,N_22570,N_24070);
nor U26658 (N_26658,N_24716,N_22684);
xor U26659 (N_26659,N_22654,N_23053);
nand U26660 (N_26660,N_22577,N_22967);
nor U26661 (N_26661,N_24317,N_22743);
nor U26662 (N_26662,N_22720,N_23478);
or U26663 (N_26663,N_24511,N_22744);
or U26664 (N_26664,N_23759,N_22844);
nor U26665 (N_26665,N_23097,N_22975);
xor U26666 (N_26666,N_23853,N_22780);
nand U26667 (N_26667,N_24739,N_23123);
nand U26668 (N_26668,N_23361,N_24989);
and U26669 (N_26669,N_23359,N_24864);
or U26670 (N_26670,N_24787,N_23292);
and U26671 (N_26671,N_22633,N_23545);
xor U26672 (N_26672,N_23615,N_24336);
nand U26673 (N_26673,N_24249,N_24029);
nor U26674 (N_26674,N_23924,N_24813);
nor U26675 (N_26675,N_23999,N_24595);
nor U26676 (N_26676,N_23778,N_24082);
or U26677 (N_26677,N_23558,N_23024);
and U26678 (N_26678,N_24076,N_24871);
nor U26679 (N_26679,N_22918,N_24629);
or U26680 (N_26680,N_23580,N_24073);
xnor U26681 (N_26681,N_24318,N_24697);
xor U26682 (N_26682,N_24732,N_24411);
or U26683 (N_26683,N_22764,N_24612);
xnor U26684 (N_26684,N_24754,N_23754);
or U26685 (N_26685,N_24922,N_24422);
and U26686 (N_26686,N_24875,N_22804);
and U26687 (N_26687,N_24005,N_23391);
or U26688 (N_26688,N_22832,N_22946);
nor U26689 (N_26689,N_24967,N_23079);
nor U26690 (N_26690,N_24718,N_22509);
nor U26691 (N_26691,N_22588,N_22627);
nor U26692 (N_26692,N_22514,N_24207);
or U26693 (N_26693,N_24548,N_22562);
or U26694 (N_26694,N_23114,N_23001);
or U26695 (N_26695,N_23738,N_24831);
and U26696 (N_26696,N_22701,N_24409);
nand U26697 (N_26697,N_24972,N_24230);
or U26698 (N_26698,N_23544,N_23729);
and U26699 (N_26699,N_23714,N_24857);
or U26700 (N_26700,N_22815,N_23288);
nand U26701 (N_26701,N_24199,N_22998);
nor U26702 (N_26702,N_24159,N_23389);
nand U26703 (N_26703,N_24323,N_24853);
or U26704 (N_26704,N_23863,N_24974);
and U26705 (N_26705,N_22993,N_24999);
and U26706 (N_26706,N_23590,N_22672);
nor U26707 (N_26707,N_23677,N_24732);
and U26708 (N_26708,N_22837,N_23278);
or U26709 (N_26709,N_24827,N_22700);
nor U26710 (N_26710,N_23262,N_23036);
or U26711 (N_26711,N_23666,N_24706);
nand U26712 (N_26712,N_24570,N_23153);
and U26713 (N_26713,N_22745,N_23076);
xnor U26714 (N_26714,N_23193,N_24532);
or U26715 (N_26715,N_24810,N_24728);
nand U26716 (N_26716,N_23016,N_22504);
and U26717 (N_26717,N_24994,N_22761);
nor U26718 (N_26718,N_23035,N_22563);
or U26719 (N_26719,N_24873,N_24981);
nor U26720 (N_26720,N_23482,N_23091);
nand U26721 (N_26721,N_23834,N_23198);
and U26722 (N_26722,N_24988,N_22665);
or U26723 (N_26723,N_22718,N_24014);
or U26724 (N_26724,N_24320,N_24413);
and U26725 (N_26725,N_22811,N_23673);
nor U26726 (N_26726,N_22658,N_23336);
and U26727 (N_26727,N_22983,N_23052);
nor U26728 (N_26728,N_23504,N_24925);
nor U26729 (N_26729,N_23340,N_22770);
and U26730 (N_26730,N_23216,N_24257);
and U26731 (N_26731,N_22828,N_23001);
xnor U26732 (N_26732,N_24595,N_24853);
xnor U26733 (N_26733,N_24513,N_22615);
nand U26734 (N_26734,N_23177,N_24846);
nor U26735 (N_26735,N_23263,N_22965);
or U26736 (N_26736,N_23029,N_24574);
and U26737 (N_26737,N_24186,N_23948);
nor U26738 (N_26738,N_22660,N_23651);
nor U26739 (N_26739,N_24251,N_23926);
or U26740 (N_26740,N_22992,N_24115);
nand U26741 (N_26741,N_23863,N_22726);
nand U26742 (N_26742,N_23653,N_24823);
nand U26743 (N_26743,N_24617,N_24725);
or U26744 (N_26744,N_22789,N_23636);
nor U26745 (N_26745,N_24185,N_22655);
or U26746 (N_26746,N_24473,N_23598);
and U26747 (N_26747,N_22578,N_23850);
nand U26748 (N_26748,N_23833,N_24114);
xnor U26749 (N_26749,N_24976,N_24430);
nor U26750 (N_26750,N_22593,N_23922);
nand U26751 (N_26751,N_23276,N_22524);
xnor U26752 (N_26752,N_23255,N_23022);
and U26753 (N_26753,N_24082,N_23432);
and U26754 (N_26754,N_24233,N_24595);
nand U26755 (N_26755,N_23272,N_24115);
or U26756 (N_26756,N_24981,N_24825);
or U26757 (N_26757,N_24100,N_22571);
or U26758 (N_26758,N_23837,N_24489);
or U26759 (N_26759,N_24571,N_24663);
nand U26760 (N_26760,N_23492,N_23719);
or U26761 (N_26761,N_22719,N_22841);
nand U26762 (N_26762,N_22879,N_23322);
or U26763 (N_26763,N_23469,N_23534);
or U26764 (N_26764,N_23281,N_24355);
or U26765 (N_26765,N_24410,N_24058);
or U26766 (N_26766,N_23806,N_23008);
nand U26767 (N_26767,N_24644,N_24936);
nand U26768 (N_26768,N_23296,N_24892);
xnor U26769 (N_26769,N_22849,N_24296);
or U26770 (N_26770,N_23968,N_23304);
nand U26771 (N_26771,N_24263,N_24526);
xor U26772 (N_26772,N_23463,N_24906);
nor U26773 (N_26773,N_24283,N_23810);
or U26774 (N_26774,N_24394,N_24471);
nand U26775 (N_26775,N_24932,N_22655);
nor U26776 (N_26776,N_24771,N_24222);
nand U26777 (N_26777,N_23049,N_24363);
and U26778 (N_26778,N_22635,N_24841);
and U26779 (N_26779,N_22900,N_24525);
or U26780 (N_26780,N_24739,N_23735);
nand U26781 (N_26781,N_24466,N_24715);
nor U26782 (N_26782,N_23481,N_23534);
nor U26783 (N_26783,N_22607,N_23577);
and U26784 (N_26784,N_24521,N_22542);
and U26785 (N_26785,N_24026,N_23847);
nand U26786 (N_26786,N_22688,N_24333);
and U26787 (N_26787,N_22733,N_24791);
nor U26788 (N_26788,N_23456,N_24211);
nand U26789 (N_26789,N_22783,N_22546);
xnor U26790 (N_26790,N_23321,N_23565);
nor U26791 (N_26791,N_22788,N_24714);
and U26792 (N_26792,N_22635,N_24861);
nand U26793 (N_26793,N_24202,N_23554);
xor U26794 (N_26794,N_23374,N_23828);
or U26795 (N_26795,N_24878,N_24568);
and U26796 (N_26796,N_23071,N_23850);
nor U26797 (N_26797,N_23563,N_23962);
or U26798 (N_26798,N_23839,N_22992);
xnor U26799 (N_26799,N_24411,N_24117);
nor U26800 (N_26800,N_24774,N_24756);
nor U26801 (N_26801,N_23416,N_23698);
nand U26802 (N_26802,N_23824,N_24387);
xnor U26803 (N_26803,N_24830,N_24163);
nand U26804 (N_26804,N_22929,N_23910);
nand U26805 (N_26805,N_22512,N_23969);
or U26806 (N_26806,N_24007,N_23036);
or U26807 (N_26807,N_24445,N_23342);
nand U26808 (N_26808,N_22804,N_23186);
xor U26809 (N_26809,N_23733,N_23451);
nor U26810 (N_26810,N_22884,N_23599);
nor U26811 (N_26811,N_24079,N_22560);
and U26812 (N_26812,N_23852,N_24251);
nor U26813 (N_26813,N_23997,N_24138);
and U26814 (N_26814,N_23943,N_23594);
xnor U26815 (N_26815,N_24355,N_24582);
nor U26816 (N_26816,N_23467,N_23492);
nor U26817 (N_26817,N_24639,N_24233);
and U26818 (N_26818,N_22854,N_24048);
nand U26819 (N_26819,N_24400,N_23171);
nand U26820 (N_26820,N_22546,N_23208);
nand U26821 (N_26821,N_24804,N_23833);
and U26822 (N_26822,N_24405,N_23494);
xnor U26823 (N_26823,N_23183,N_22869);
nor U26824 (N_26824,N_23489,N_24359);
and U26825 (N_26825,N_24875,N_23802);
nand U26826 (N_26826,N_24197,N_24137);
nand U26827 (N_26827,N_23117,N_24868);
nor U26828 (N_26828,N_22918,N_24426);
nand U26829 (N_26829,N_23875,N_24234);
nand U26830 (N_26830,N_24861,N_24207);
or U26831 (N_26831,N_23640,N_23490);
nor U26832 (N_26832,N_22760,N_24979);
or U26833 (N_26833,N_23627,N_24812);
nor U26834 (N_26834,N_22897,N_24287);
nor U26835 (N_26835,N_24974,N_22934);
nor U26836 (N_26836,N_23549,N_22609);
and U26837 (N_26837,N_24894,N_23654);
and U26838 (N_26838,N_24771,N_22801);
and U26839 (N_26839,N_23082,N_23175);
and U26840 (N_26840,N_22756,N_23363);
nand U26841 (N_26841,N_23384,N_23357);
nor U26842 (N_26842,N_24783,N_24163);
xnor U26843 (N_26843,N_23365,N_24905);
or U26844 (N_26844,N_23528,N_23482);
or U26845 (N_26845,N_23256,N_23985);
nor U26846 (N_26846,N_24234,N_23444);
or U26847 (N_26847,N_24779,N_23029);
and U26848 (N_26848,N_24732,N_23718);
and U26849 (N_26849,N_23777,N_24650);
or U26850 (N_26850,N_22646,N_23232);
nand U26851 (N_26851,N_22828,N_23031);
and U26852 (N_26852,N_22641,N_24688);
and U26853 (N_26853,N_24740,N_23354);
and U26854 (N_26854,N_23053,N_24052);
nor U26855 (N_26855,N_23487,N_24985);
and U26856 (N_26856,N_23932,N_23516);
nor U26857 (N_26857,N_22720,N_22579);
or U26858 (N_26858,N_23715,N_24257);
nand U26859 (N_26859,N_24109,N_22542);
and U26860 (N_26860,N_23373,N_23328);
nor U26861 (N_26861,N_24273,N_24397);
nand U26862 (N_26862,N_23629,N_22608);
or U26863 (N_26863,N_23117,N_24224);
or U26864 (N_26864,N_24541,N_24733);
or U26865 (N_26865,N_24339,N_23474);
xnor U26866 (N_26866,N_23621,N_23082);
and U26867 (N_26867,N_24889,N_22781);
and U26868 (N_26868,N_23430,N_23174);
nor U26869 (N_26869,N_22618,N_24574);
nor U26870 (N_26870,N_23501,N_23099);
nand U26871 (N_26871,N_24781,N_24855);
nand U26872 (N_26872,N_24103,N_24112);
and U26873 (N_26873,N_23807,N_23575);
nand U26874 (N_26874,N_24971,N_22983);
nand U26875 (N_26875,N_24009,N_22840);
nand U26876 (N_26876,N_24242,N_24770);
or U26877 (N_26877,N_24356,N_24272);
and U26878 (N_26878,N_22968,N_24482);
nor U26879 (N_26879,N_22867,N_23606);
nor U26880 (N_26880,N_23709,N_24854);
nand U26881 (N_26881,N_22521,N_23670);
nor U26882 (N_26882,N_24424,N_24933);
or U26883 (N_26883,N_22589,N_22803);
nand U26884 (N_26884,N_24642,N_24928);
nand U26885 (N_26885,N_22871,N_23104);
nand U26886 (N_26886,N_24118,N_24015);
nor U26887 (N_26887,N_24850,N_24362);
xor U26888 (N_26888,N_23084,N_24782);
and U26889 (N_26889,N_24618,N_23074);
and U26890 (N_26890,N_23645,N_22706);
or U26891 (N_26891,N_24429,N_24519);
nor U26892 (N_26892,N_23411,N_22642);
and U26893 (N_26893,N_23471,N_24463);
or U26894 (N_26894,N_23093,N_24151);
nand U26895 (N_26895,N_24998,N_24741);
or U26896 (N_26896,N_22683,N_24812);
xnor U26897 (N_26897,N_23479,N_23541);
nand U26898 (N_26898,N_23425,N_24250);
and U26899 (N_26899,N_24678,N_23845);
nor U26900 (N_26900,N_24728,N_24915);
nand U26901 (N_26901,N_22638,N_22844);
nor U26902 (N_26902,N_24386,N_22744);
and U26903 (N_26903,N_24699,N_23148);
or U26904 (N_26904,N_24348,N_24552);
and U26905 (N_26905,N_24248,N_22771);
nor U26906 (N_26906,N_23762,N_23067);
nor U26907 (N_26907,N_23794,N_23748);
nand U26908 (N_26908,N_23456,N_23534);
nand U26909 (N_26909,N_23698,N_23002);
nor U26910 (N_26910,N_23084,N_24029);
nand U26911 (N_26911,N_23397,N_23515);
nor U26912 (N_26912,N_22957,N_22582);
nand U26913 (N_26913,N_24436,N_23926);
nand U26914 (N_26914,N_23036,N_23549);
or U26915 (N_26915,N_23928,N_24985);
nand U26916 (N_26916,N_23032,N_24505);
xnor U26917 (N_26917,N_22754,N_24537);
nand U26918 (N_26918,N_23579,N_23288);
or U26919 (N_26919,N_22783,N_24059);
and U26920 (N_26920,N_24948,N_24877);
and U26921 (N_26921,N_23807,N_24436);
and U26922 (N_26922,N_23874,N_24964);
xor U26923 (N_26923,N_24961,N_23617);
nor U26924 (N_26924,N_24067,N_23285);
nor U26925 (N_26925,N_23775,N_22652);
xor U26926 (N_26926,N_23666,N_23348);
xor U26927 (N_26927,N_23158,N_24435);
or U26928 (N_26928,N_23253,N_22940);
nor U26929 (N_26929,N_24742,N_24315);
or U26930 (N_26930,N_24187,N_24026);
nand U26931 (N_26931,N_23419,N_24746);
and U26932 (N_26932,N_24372,N_22614);
or U26933 (N_26933,N_24501,N_22618);
nand U26934 (N_26934,N_22936,N_23711);
xnor U26935 (N_26935,N_24917,N_23385);
and U26936 (N_26936,N_23936,N_23095);
and U26937 (N_26937,N_24300,N_24078);
nand U26938 (N_26938,N_23509,N_22966);
or U26939 (N_26939,N_22525,N_24373);
nor U26940 (N_26940,N_24895,N_22593);
nor U26941 (N_26941,N_24053,N_22524);
or U26942 (N_26942,N_23776,N_22543);
nor U26943 (N_26943,N_24196,N_23492);
or U26944 (N_26944,N_24760,N_24823);
or U26945 (N_26945,N_23023,N_24861);
nor U26946 (N_26946,N_24291,N_22574);
nor U26947 (N_26947,N_24699,N_22914);
and U26948 (N_26948,N_24486,N_23624);
or U26949 (N_26949,N_23355,N_24058);
nand U26950 (N_26950,N_22684,N_23144);
nor U26951 (N_26951,N_23096,N_23283);
or U26952 (N_26952,N_24707,N_24886);
nand U26953 (N_26953,N_23139,N_24636);
nand U26954 (N_26954,N_23798,N_23097);
nand U26955 (N_26955,N_24311,N_24524);
or U26956 (N_26956,N_24019,N_22707);
nor U26957 (N_26957,N_24132,N_22960);
or U26958 (N_26958,N_24498,N_23415);
and U26959 (N_26959,N_23880,N_22714);
and U26960 (N_26960,N_23105,N_24948);
or U26961 (N_26961,N_23668,N_23102);
nor U26962 (N_26962,N_23859,N_24073);
nand U26963 (N_26963,N_24836,N_22922);
and U26964 (N_26964,N_24923,N_23268);
or U26965 (N_26965,N_23688,N_23767);
nand U26966 (N_26966,N_23921,N_23133);
nand U26967 (N_26967,N_24459,N_24122);
nor U26968 (N_26968,N_23622,N_22620);
or U26969 (N_26969,N_24798,N_22786);
nand U26970 (N_26970,N_22929,N_22864);
nor U26971 (N_26971,N_23171,N_23521);
or U26972 (N_26972,N_24526,N_24979);
xor U26973 (N_26973,N_23955,N_24614);
nand U26974 (N_26974,N_22825,N_23925);
nor U26975 (N_26975,N_23917,N_22874);
and U26976 (N_26976,N_23197,N_24575);
xnor U26977 (N_26977,N_22714,N_24923);
nor U26978 (N_26978,N_24058,N_24897);
nand U26979 (N_26979,N_22580,N_24530);
nand U26980 (N_26980,N_24542,N_22501);
xnor U26981 (N_26981,N_23699,N_22692);
and U26982 (N_26982,N_23195,N_24501);
and U26983 (N_26983,N_22980,N_24369);
nor U26984 (N_26984,N_22559,N_24182);
nand U26985 (N_26985,N_23268,N_24408);
nand U26986 (N_26986,N_22586,N_24215);
nand U26987 (N_26987,N_24653,N_22558);
or U26988 (N_26988,N_23891,N_23553);
or U26989 (N_26989,N_22914,N_23828);
nand U26990 (N_26990,N_24937,N_24467);
and U26991 (N_26991,N_23527,N_23434);
and U26992 (N_26992,N_23797,N_24364);
and U26993 (N_26993,N_24016,N_23588);
nor U26994 (N_26994,N_22670,N_24389);
or U26995 (N_26995,N_23018,N_23539);
or U26996 (N_26996,N_24158,N_24406);
xor U26997 (N_26997,N_23668,N_24536);
xnor U26998 (N_26998,N_24897,N_23695);
nand U26999 (N_26999,N_23464,N_23590);
or U27000 (N_27000,N_23684,N_22683);
and U27001 (N_27001,N_24328,N_23839);
nor U27002 (N_27002,N_24181,N_23911);
nor U27003 (N_27003,N_23790,N_23398);
or U27004 (N_27004,N_24113,N_22646);
or U27005 (N_27005,N_23743,N_24726);
or U27006 (N_27006,N_22686,N_24959);
and U27007 (N_27007,N_23993,N_24398);
or U27008 (N_27008,N_23221,N_22884);
or U27009 (N_27009,N_22672,N_23449);
or U27010 (N_27010,N_24981,N_22611);
nor U27011 (N_27011,N_23368,N_23349);
nor U27012 (N_27012,N_22723,N_23908);
nor U27013 (N_27013,N_22809,N_24109);
nor U27014 (N_27014,N_22552,N_23359);
and U27015 (N_27015,N_22979,N_24556);
nor U27016 (N_27016,N_23742,N_23567);
nand U27017 (N_27017,N_22972,N_23484);
nor U27018 (N_27018,N_22714,N_24334);
xnor U27019 (N_27019,N_23935,N_22647);
or U27020 (N_27020,N_23681,N_24444);
xnor U27021 (N_27021,N_24374,N_24172);
nand U27022 (N_27022,N_23918,N_23151);
and U27023 (N_27023,N_23394,N_22702);
nor U27024 (N_27024,N_23261,N_22755);
nand U27025 (N_27025,N_23247,N_24400);
nor U27026 (N_27026,N_23457,N_23513);
nand U27027 (N_27027,N_24283,N_24739);
nand U27028 (N_27028,N_22557,N_23676);
nand U27029 (N_27029,N_23054,N_24515);
nand U27030 (N_27030,N_23174,N_23302);
nor U27031 (N_27031,N_23526,N_23316);
or U27032 (N_27032,N_24063,N_24006);
and U27033 (N_27033,N_23159,N_23821);
nor U27034 (N_27034,N_24898,N_23304);
nand U27035 (N_27035,N_24094,N_23748);
and U27036 (N_27036,N_23187,N_22979);
nand U27037 (N_27037,N_23115,N_23683);
and U27038 (N_27038,N_23323,N_24876);
nor U27039 (N_27039,N_24268,N_22501);
or U27040 (N_27040,N_24816,N_22932);
or U27041 (N_27041,N_24006,N_24076);
nor U27042 (N_27042,N_24384,N_22693);
nor U27043 (N_27043,N_22941,N_23751);
nor U27044 (N_27044,N_22792,N_23656);
nor U27045 (N_27045,N_23580,N_23776);
nand U27046 (N_27046,N_24016,N_24320);
and U27047 (N_27047,N_22514,N_24583);
nand U27048 (N_27048,N_23590,N_24287);
nand U27049 (N_27049,N_23149,N_23299);
nand U27050 (N_27050,N_23072,N_23453);
nand U27051 (N_27051,N_22726,N_23996);
nand U27052 (N_27052,N_23404,N_22869);
nand U27053 (N_27053,N_22979,N_24606);
xnor U27054 (N_27054,N_23275,N_24872);
nor U27055 (N_27055,N_23195,N_22732);
nand U27056 (N_27056,N_24543,N_23919);
and U27057 (N_27057,N_24139,N_24545);
nor U27058 (N_27058,N_24958,N_23960);
nand U27059 (N_27059,N_24212,N_23182);
or U27060 (N_27060,N_24608,N_24142);
or U27061 (N_27061,N_23584,N_22664);
nor U27062 (N_27062,N_23081,N_24460);
nor U27063 (N_27063,N_23233,N_23728);
nand U27064 (N_27064,N_22950,N_22548);
xnor U27065 (N_27065,N_23968,N_22531);
nor U27066 (N_27066,N_23620,N_23091);
and U27067 (N_27067,N_22878,N_23478);
or U27068 (N_27068,N_22941,N_24068);
and U27069 (N_27069,N_23576,N_23075);
and U27070 (N_27070,N_23458,N_23794);
nor U27071 (N_27071,N_22925,N_24770);
and U27072 (N_27072,N_23729,N_23453);
xnor U27073 (N_27073,N_23959,N_24838);
and U27074 (N_27074,N_23781,N_22524);
nand U27075 (N_27075,N_23684,N_23279);
nor U27076 (N_27076,N_24946,N_23319);
xor U27077 (N_27077,N_24055,N_23488);
nor U27078 (N_27078,N_22639,N_23283);
xor U27079 (N_27079,N_24881,N_23243);
nor U27080 (N_27080,N_23641,N_24328);
and U27081 (N_27081,N_23819,N_24453);
nand U27082 (N_27082,N_22731,N_23653);
and U27083 (N_27083,N_23342,N_22509);
nand U27084 (N_27084,N_23870,N_23885);
or U27085 (N_27085,N_23735,N_23690);
nor U27086 (N_27086,N_24318,N_24933);
xnor U27087 (N_27087,N_24629,N_23753);
and U27088 (N_27088,N_23708,N_24580);
and U27089 (N_27089,N_23619,N_24811);
nor U27090 (N_27090,N_24520,N_24551);
xor U27091 (N_27091,N_24883,N_23668);
nand U27092 (N_27092,N_23218,N_24964);
nor U27093 (N_27093,N_24936,N_24938);
xnor U27094 (N_27094,N_23164,N_23227);
nor U27095 (N_27095,N_22700,N_24815);
and U27096 (N_27096,N_23783,N_23626);
xnor U27097 (N_27097,N_23241,N_24737);
or U27098 (N_27098,N_24271,N_24234);
xor U27099 (N_27099,N_22618,N_22578);
nor U27100 (N_27100,N_24379,N_23456);
nand U27101 (N_27101,N_22873,N_24112);
nand U27102 (N_27102,N_24820,N_23407);
and U27103 (N_27103,N_24565,N_22673);
or U27104 (N_27104,N_24449,N_24189);
nor U27105 (N_27105,N_23057,N_23222);
and U27106 (N_27106,N_24469,N_24359);
xnor U27107 (N_27107,N_24463,N_23825);
nor U27108 (N_27108,N_24126,N_24876);
nor U27109 (N_27109,N_24501,N_24697);
nand U27110 (N_27110,N_24005,N_23894);
and U27111 (N_27111,N_24044,N_23224);
nor U27112 (N_27112,N_23184,N_23062);
nor U27113 (N_27113,N_23171,N_23653);
nor U27114 (N_27114,N_22835,N_23107);
or U27115 (N_27115,N_24434,N_22604);
nor U27116 (N_27116,N_23855,N_24269);
or U27117 (N_27117,N_22559,N_22567);
nor U27118 (N_27118,N_23914,N_23491);
and U27119 (N_27119,N_23118,N_24031);
nor U27120 (N_27120,N_24485,N_23781);
nand U27121 (N_27121,N_23764,N_23788);
nand U27122 (N_27122,N_23409,N_22573);
nand U27123 (N_27123,N_22708,N_24385);
nand U27124 (N_27124,N_23979,N_23330);
nor U27125 (N_27125,N_23210,N_24184);
or U27126 (N_27126,N_24485,N_23436);
or U27127 (N_27127,N_22649,N_23592);
nand U27128 (N_27128,N_23414,N_22576);
or U27129 (N_27129,N_23294,N_24534);
and U27130 (N_27130,N_24209,N_23820);
or U27131 (N_27131,N_22708,N_22844);
nor U27132 (N_27132,N_22786,N_23277);
nor U27133 (N_27133,N_23279,N_22985);
nor U27134 (N_27134,N_23143,N_22921);
nor U27135 (N_27135,N_22827,N_24702);
nand U27136 (N_27136,N_23923,N_24893);
and U27137 (N_27137,N_24873,N_23866);
or U27138 (N_27138,N_22653,N_24509);
and U27139 (N_27139,N_24741,N_24696);
nor U27140 (N_27140,N_24825,N_23023);
or U27141 (N_27141,N_23598,N_22889);
and U27142 (N_27142,N_22852,N_23768);
nand U27143 (N_27143,N_22913,N_23535);
nand U27144 (N_27144,N_24533,N_24408);
nor U27145 (N_27145,N_23221,N_24196);
or U27146 (N_27146,N_22888,N_23849);
or U27147 (N_27147,N_23656,N_24105);
or U27148 (N_27148,N_24671,N_24055);
and U27149 (N_27149,N_23556,N_23567);
nor U27150 (N_27150,N_24188,N_24212);
and U27151 (N_27151,N_22505,N_24476);
nor U27152 (N_27152,N_23577,N_23999);
and U27153 (N_27153,N_24649,N_24528);
or U27154 (N_27154,N_24910,N_22709);
nor U27155 (N_27155,N_24320,N_24003);
nand U27156 (N_27156,N_22979,N_23084);
nor U27157 (N_27157,N_24189,N_24544);
and U27158 (N_27158,N_22777,N_23541);
or U27159 (N_27159,N_23710,N_24656);
and U27160 (N_27160,N_22880,N_23241);
xnor U27161 (N_27161,N_22713,N_23893);
nand U27162 (N_27162,N_23839,N_24990);
or U27163 (N_27163,N_23591,N_24645);
nor U27164 (N_27164,N_24726,N_24021);
or U27165 (N_27165,N_24868,N_23268);
nand U27166 (N_27166,N_24361,N_23556);
nand U27167 (N_27167,N_23945,N_24837);
nor U27168 (N_27168,N_22820,N_24889);
or U27169 (N_27169,N_22730,N_24181);
or U27170 (N_27170,N_23039,N_24520);
nand U27171 (N_27171,N_23631,N_23259);
nand U27172 (N_27172,N_23029,N_24984);
nand U27173 (N_27173,N_24391,N_24826);
nand U27174 (N_27174,N_23297,N_22735);
nand U27175 (N_27175,N_22657,N_24722);
and U27176 (N_27176,N_22814,N_24458);
and U27177 (N_27177,N_24354,N_24430);
and U27178 (N_27178,N_24786,N_23902);
xor U27179 (N_27179,N_24878,N_24966);
nand U27180 (N_27180,N_22685,N_24541);
or U27181 (N_27181,N_23860,N_22973);
nand U27182 (N_27182,N_24051,N_22875);
nand U27183 (N_27183,N_24937,N_23028);
or U27184 (N_27184,N_24186,N_22922);
nor U27185 (N_27185,N_23713,N_23113);
and U27186 (N_27186,N_23663,N_22806);
and U27187 (N_27187,N_22744,N_23740);
nand U27188 (N_27188,N_23922,N_23993);
or U27189 (N_27189,N_23673,N_23342);
nor U27190 (N_27190,N_23982,N_22945);
nor U27191 (N_27191,N_23861,N_24611);
nor U27192 (N_27192,N_24487,N_23169);
and U27193 (N_27193,N_24705,N_23695);
nand U27194 (N_27194,N_24922,N_23537);
and U27195 (N_27195,N_23146,N_24618);
nand U27196 (N_27196,N_24563,N_23411);
and U27197 (N_27197,N_24301,N_24464);
xor U27198 (N_27198,N_24078,N_24174);
or U27199 (N_27199,N_23240,N_23370);
nor U27200 (N_27200,N_23821,N_23066);
nor U27201 (N_27201,N_23841,N_22923);
and U27202 (N_27202,N_24419,N_23424);
nor U27203 (N_27203,N_24534,N_23600);
nand U27204 (N_27204,N_24078,N_22839);
and U27205 (N_27205,N_24056,N_22550);
or U27206 (N_27206,N_23597,N_24861);
nor U27207 (N_27207,N_24120,N_23874);
and U27208 (N_27208,N_23673,N_22904);
and U27209 (N_27209,N_24393,N_24404);
nand U27210 (N_27210,N_24503,N_22587);
nor U27211 (N_27211,N_24646,N_23125);
xnor U27212 (N_27212,N_23564,N_22964);
xor U27213 (N_27213,N_24122,N_23313);
and U27214 (N_27214,N_22706,N_24318);
and U27215 (N_27215,N_23534,N_24958);
or U27216 (N_27216,N_24663,N_23043);
nand U27217 (N_27217,N_23392,N_23474);
nor U27218 (N_27218,N_24280,N_22504);
or U27219 (N_27219,N_23948,N_24378);
xnor U27220 (N_27220,N_24797,N_24862);
and U27221 (N_27221,N_22916,N_22666);
nor U27222 (N_27222,N_22850,N_22728);
nand U27223 (N_27223,N_22670,N_23656);
nor U27224 (N_27224,N_23399,N_23484);
and U27225 (N_27225,N_22730,N_23885);
and U27226 (N_27226,N_23922,N_24417);
nor U27227 (N_27227,N_24913,N_22668);
or U27228 (N_27228,N_24013,N_23545);
or U27229 (N_27229,N_23930,N_23897);
and U27230 (N_27230,N_24806,N_24642);
nor U27231 (N_27231,N_22700,N_23226);
nand U27232 (N_27232,N_24925,N_22682);
nor U27233 (N_27233,N_24338,N_23537);
or U27234 (N_27234,N_23660,N_24675);
xor U27235 (N_27235,N_23642,N_24455);
nor U27236 (N_27236,N_23377,N_24073);
nand U27237 (N_27237,N_23883,N_24358);
nor U27238 (N_27238,N_24907,N_23304);
or U27239 (N_27239,N_24469,N_24749);
nand U27240 (N_27240,N_24235,N_23773);
and U27241 (N_27241,N_23723,N_22958);
nor U27242 (N_27242,N_24120,N_24596);
nor U27243 (N_27243,N_23183,N_24139);
xnor U27244 (N_27244,N_24052,N_22512);
or U27245 (N_27245,N_23348,N_23017);
nor U27246 (N_27246,N_23785,N_24088);
nand U27247 (N_27247,N_22764,N_24036);
or U27248 (N_27248,N_23343,N_23933);
or U27249 (N_27249,N_23525,N_22691);
nor U27250 (N_27250,N_24433,N_23501);
xor U27251 (N_27251,N_24692,N_24500);
and U27252 (N_27252,N_24480,N_23889);
and U27253 (N_27253,N_24587,N_24924);
nand U27254 (N_27254,N_23856,N_23408);
nor U27255 (N_27255,N_24358,N_22518);
and U27256 (N_27256,N_24866,N_24321);
and U27257 (N_27257,N_24598,N_24658);
nor U27258 (N_27258,N_24272,N_23630);
nor U27259 (N_27259,N_24389,N_24432);
nand U27260 (N_27260,N_22722,N_23238);
xnor U27261 (N_27261,N_24763,N_24980);
nand U27262 (N_27262,N_22670,N_23879);
nor U27263 (N_27263,N_22616,N_24292);
or U27264 (N_27264,N_24807,N_24516);
nand U27265 (N_27265,N_23171,N_23677);
xnor U27266 (N_27266,N_24608,N_22545);
nor U27267 (N_27267,N_24073,N_24740);
and U27268 (N_27268,N_23579,N_22934);
xnor U27269 (N_27269,N_22927,N_23109);
and U27270 (N_27270,N_24515,N_23991);
nand U27271 (N_27271,N_24952,N_24360);
nand U27272 (N_27272,N_24944,N_23466);
nor U27273 (N_27273,N_23127,N_22905);
nor U27274 (N_27274,N_24777,N_24751);
nand U27275 (N_27275,N_24190,N_24889);
and U27276 (N_27276,N_24171,N_23542);
nor U27277 (N_27277,N_22862,N_23651);
and U27278 (N_27278,N_22883,N_22531);
and U27279 (N_27279,N_24111,N_22524);
or U27280 (N_27280,N_22841,N_23319);
nand U27281 (N_27281,N_24954,N_23294);
nor U27282 (N_27282,N_22788,N_23188);
nor U27283 (N_27283,N_23519,N_23354);
and U27284 (N_27284,N_23498,N_23491);
nand U27285 (N_27285,N_23227,N_23811);
and U27286 (N_27286,N_24143,N_24772);
nand U27287 (N_27287,N_22921,N_24087);
or U27288 (N_27288,N_23850,N_24109);
nor U27289 (N_27289,N_23495,N_23747);
xor U27290 (N_27290,N_24833,N_24794);
nand U27291 (N_27291,N_24847,N_23072);
and U27292 (N_27292,N_24424,N_24667);
and U27293 (N_27293,N_23990,N_24354);
or U27294 (N_27294,N_24776,N_22830);
and U27295 (N_27295,N_23233,N_24645);
nor U27296 (N_27296,N_22589,N_23830);
and U27297 (N_27297,N_22747,N_23539);
xnor U27298 (N_27298,N_22711,N_23573);
and U27299 (N_27299,N_23062,N_24205);
nand U27300 (N_27300,N_24127,N_22891);
nand U27301 (N_27301,N_22704,N_24854);
nor U27302 (N_27302,N_24732,N_24930);
nor U27303 (N_27303,N_24835,N_24586);
nor U27304 (N_27304,N_24828,N_22620);
nand U27305 (N_27305,N_23448,N_24720);
nor U27306 (N_27306,N_22838,N_23971);
nor U27307 (N_27307,N_23049,N_22751);
and U27308 (N_27308,N_24628,N_24711);
and U27309 (N_27309,N_23806,N_23913);
nand U27310 (N_27310,N_24492,N_23383);
or U27311 (N_27311,N_23587,N_22709);
nor U27312 (N_27312,N_23941,N_23083);
or U27313 (N_27313,N_23659,N_22762);
nand U27314 (N_27314,N_22567,N_23078);
xnor U27315 (N_27315,N_23772,N_22761);
and U27316 (N_27316,N_22832,N_24025);
nor U27317 (N_27317,N_24964,N_23238);
nor U27318 (N_27318,N_22824,N_24678);
or U27319 (N_27319,N_24249,N_23773);
and U27320 (N_27320,N_22541,N_23305);
and U27321 (N_27321,N_23626,N_23649);
and U27322 (N_27322,N_24291,N_23105);
nor U27323 (N_27323,N_23356,N_23570);
nor U27324 (N_27324,N_23021,N_24671);
and U27325 (N_27325,N_22705,N_23305);
and U27326 (N_27326,N_22601,N_23240);
nand U27327 (N_27327,N_23363,N_23477);
or U27328 (N_27328,N_22975,N_22988);
or U27329 (N_27329,N_24400,N_23624);
or U27330 (N_27330,N_23691,N_23718);
or U27331 (N_27331,N_24192,N_23358);
and U27332 (N_27332,N_23672,N_23651);
nor U27333 (N_27333,N_22963,N_23408);
and U27334 (N_27334,N_24898,N_23105);
nand U27335 (N_27335,N_24378,N_22636);
or U27336 (N_27336,N_23599,N_23764);
or U27337 (N_27337,N_24173,N_24297);
or U27338 (N_27338,N_24320,N_22578);
nand U27339 (N_27339,N_24306,N_22817);
nor U27340 (N_27340,N_24246,N_22524);
and U27341 (N_27341,N_23762,N_23058);
and U27342 (N_27342,N_24603,N_24800);
and U27343 (N_27343,N_24829,N_22782);
nor U27344 (N_27344,N_24616,N_23317);
or U27345 (N_27345,N_23587,N_24062);
nand U27346 (N_27346,N_23002,N_23901);
and U27347 (N_27347,N_23148,N_24801);
or U27348 (N_27348,N_24946,N_23793);
nor U27349 (N_27349,N_23126,N_24992);
xnor U27350 (N_27350,N_22989,N_23660);
and U27351 (N_27351,N_23594,N_24765);
and U27352 (N_27352,N_24368,N_23198);
nor U27353 (N_27353,N_22561,N_22917);
nor U27354 (N_27354,N_24498,N_23644);
nor U27355 (N_27355,N_23638,N_24223);
nor U27356 (N_27356,N_23575,N_24523);
and U27357 (N_27357,N_23454,N_22761);
nand U27358 (N_27358,N_23297,N_24290);
nor U27359 (N_27359,N_23159,N_23005);
and U27360 (N_27360,N_23160,N_24799);
nor U27361 (N_27361,N_22503,N_23062);
nor U27362 (N_27362,N_23886,N_24455);
nor U27363 (N_27363,N_23595,N_23163);
nand U27364 (N_27364,N_24130,N_22830);
or U27365 (N_27365,N_24374,N_24017);
and U27366 (N_27366,N_23074,N_23039);
or U27367 (N_27367,N_22833,N_23749);
nand U27368 (N_27368,N_22992,N_22671);
nor U27369 (N_27369,N_23116,N_22596);
and U27370 (N_27370,N_24875,N_23217);
or U27371 (N_27371,N_24266,N_22912);
nand U27372 (N_27372,N_23491,N_23020);
nor U27373 (N_27373,N_24895,N_23080);
nand U27374 (N_27374,N_22624,N_24634);
nand U27375 (N_27375,N_23760,N_24582);
xor U27376 (N_27376,N_24534,N_23132);
or U27377 (N_27377,N_24010,N_23595);
and U27378 (N_27378,N_23679,N_22502);
or U27379 (N_27379,N_23973,N_23393);
nor U27380 (N_27380,N_24109,N_22556);
and U27381 (N_27381,N_23009,N_23232);
or U27382 (N_27382,N_23095,N_23814);
nor U27383 (N_27383,N_22736,N_24303);
nor U27384 (N_27384,N_23284,N_23890);
nand U27385 (N_27385,N_22817,N_24010);
or U27386 (N_27386,N_22581,N_24009);
nor U27387 (N_27387,N_23729,N_23566);
or U27388 (N_27388,N_24308,N_24488);
or U27389 (N_27389,N_23863,N_24414);
or U27390 (N_27390,N_22797,N_24175);
nor U27391 (N_27391,N_23289,N_24754);
nand U27392 (N_27392,N_24779,N_24416);
nor U27393 (N_27393,N_24347,N_24773);
or U27394 (N_27394,N_23503,N_24144);
or U27395 (N_27395,N_24510,N_22871);
or U27396 (N_27396,N_24649,N_23001);
nand U27397 (N_27397,N_22931,N_22961);
xor U27398 (N_27398,N_23914,N_24358);
or U27399 (N_27399,N_23646,N_23036);
and U27400 (N_27400,N_22737,N_23526);
nor U27401 (N_27401,N_23160,N_24285);
nand U27402 (N_27402,N_24791,N_22714);
or U27403 (N_27403,N_24276,N_24734);
nor U27404 (N_27404,N_23582,N_24351);
and U27405 (N_27405,N_24157,N_24156);
or U27406 (N_27406,N_24607,N_23647);
nand U27407 (N_27407,N_22663,N_22551);
or U27408 (N_27408,N_23900,N_24270);
nand U27409 (N_27409,N_24212,N_23815);
nand U27410 (N_27410,N_22952,N_23155);
and U27411 (N_27411,N_24778,N_22531);
or U27412 (N_27412,N_24672,N_24220);
xnor U27413 (N_27413,N_24987,N_23305);
or U27414 (N_27414,N_23070,N_24820);
nand U27415 (N_27415,N_22556,N_23507);
nor U27416 (N_27416,N_24767,N_23134);
nand U27417 (N_27417,N_22649,N_23447);
or U27418 (N_27418,N_23873,N_23974);
nor U27419 (N_27419,N_22794,N_23063);
nand U27420 (N_27420,N_23433,N_23454);
and U27421 (N_27421,N_22535,N_24911);
xor U27422 (N_27422,N_22511,N_24287);
or U27423 (N_27423,N_23850,N_23932);
nand U27424 (N_27424,N_24010,N_22578);
nand U27425 (N_27425,N_24564,N_24290);
nand U27426 (N_27426,N_22822,N_22837);
and U27427 (N_27427,N_22739,N_23671);
nor U27428 (N_27428,N_23937,N_22779);
xnor U27429 (N_27429,N_23317,N_23516);
or U27430 (N_27430,N_24632,N_22886);
and U27431 (N_27431,N_23660,N_24754);
xor U27432 (N_27432,N_24134,N_22925);
nor U27433 (N_27433,N_23753,N_24265);
nand U27434 (N_27434,N_24035,N_22851);
and U27435 (N_27435,N_24024,N_23275);
and U27436 (N_27436,N_24806,N_24490);
nand U27437 (N_27437,N_24971,N_22685);
or U27438 (N_27438,N_22739,N_23916);
or U27439 (N_27439,N_24799,N_23693);
nor U27440 (N_27440,N_22657,N_23104);
or U27441 (N_27441,N_22603,N_23193);
nor U27442 (N_27442,N_24799,N_23905);
nand U27443 (N_27443,N_22549,N_22915);
and U27444 (N_27444,N_23560,N_23826);
nor U27445 (N_27445,N_22573,N_22905);
nor U27446 (N_27446,N_23845,N_24797);
or U27447 (N_27447,N_24849,N_24448);
and U27448 (N_27448,N_23717,N_22840);
nor U27449 (N_27449,N_23885,N_24285);
nor U27450 (N_27450,N_24971,N_23250);
nor U27451 (N_27451,N_23583,N_24635);
nor U27452 (N_27452,N_24951,N_22959);
nor U27453 (N_27453,N_24894,N_23661);
nor U27454 (N_27454,N_22839,N_23844);
nand U27455 (N_27455,N_23405,N_23606);
or U27456 (N_27456,N_24862,N_22929);
nand U27457 (N_27457,N_22912,N_23491);
nor U27458 (N_27458,N_22918,N_23297);
or U27459 (N_27459,N_24704,N_23091);
nand U27460 (N_27460,N_22627,N_23227);
nor U27461 (N_27461,N_24726,N_24651);
nor U27462 (N_27462,N_24635,N_23326);
or U27463 (N_27463,N_24459,N_23421);
or U27464 (N_27464,N_24798,N_24301);
or U27465 (N_27465,N_24801,N_22646);
and U27466 (N_27466,N_24576,N_24843);
or U27467 (N_27467,N_23131,N_23953);
xor U27468 (N_27468,N_22554,N_24739);
and U27469 (N_27469,N_24040,N_23254);
nand U27470 (N_27470,N_24934,N_23856);
and U27471 (N_27471,N_24161,N_24148);
nand U27472 (N_27472,N_24346,N_24679);
nor U27473 (N_27473,N_23457,N_24235);
or U27474 (N_27474,N_24688,N_22760);
nand U27475 (N_27475,N_24437,N_22968);
and U27476 (N_27476,N_22548,N_24622);
nand U27477 (N_27477,N_22594,N_24869);
xor U27478 (N_27478,N_23325,N_22625);
and U27479 (N_27479,N_23305,N_23558);
nor U27480 (N_27480,N_23207,N_24272);
and U27481 (N_27481,N_23679,N_22747);
nor U27482 (N_27482,N_24750,N_23256);
nor U27483 (N_27483,N_23233,N_22960);
nor U27484 (N_27484,N_23148,N_23538);
nor U27485 (N_27485,N_23877,N_23186);
and U27486 (N_27486,N_24502,N_22657);
and U27487 (N_27487,N_23814,N_23722);
nor U27488 (N_27488,N_23888,N_24741);
nor U27489 (N_27489,N_23145,N_24313);
nor U27490 (N_27490,N_24092,N_24332);
or U27491 (N_27491,N_22631,N_24712);
nor U27492 (N_27492,N_23918,N_24526);
nor U27493 (N_27493,N_23178,N_23409);
and U27494 (N_27494,N_23262,N_23705);
and U27495 (N_27495,N_24369,N_23181);
or U27496 (N_27496,N_24418,N_23536);
nor U27497 (N_27497,N_22563,N_24698);
nand U27498 (N_27498,N_23129,N_23669);
nor U27499 (N_27499,N_22540,N_24147);
or U27500 (N_27500,N_26320,N_26384);
and U27501 (N_27501,N_27038,N_25735);
nor U27502 (N_27502,N_26364,N_26629);
nand U27503 (N_27503,N_26668,N_26980);
and U27504 (N_27504,N_27467,N_27353);
and U27505 (N_27505,N_25654,N_26662);
and U27506 (N_27506,N_26479,N_25430);
nor U27507 (N_27507,N_25083,N_26904);
nor U27508 (N_27508,N_25760,N_27156);
nor U27509 (N_27509,N_25614,N_25959);
or U27510 (N_27510,N_27194,N_25167);
nand U27511 (N_27511,N_25973,N_25867);
or U27512 (N_27512,N_26601,N_25473);
or U27513 (N_27513,N_26416,N_25633);
and U27514 (N_27514,N_25099,N_25953);
nand U27515 (N_27515,N_27248,N_25252);
and U27516 (N_27516,N_25608,N_25024);
nor U27517 (N_27517,N_26190,N_26971);
or U27518 (N_27518,N_26068,N_26071);
or U27519 (N_27519,N_27050,N_26468);
or U27520 (N_27520,N_25928,N_25085);
nor U27521 (N_27521,N_25896,N_26221);
xnor U27522 (N_27522,N_26218,N_25849);
nor U27523 (N_27523,N_26721,N_25926);
and U27524 (N_27524,N_26767,N_26982);
and U27525 (N_27525,N_25979,N_25182);
or U27526 (N_27526,N_26185,N_26739);
or U27527 (N_27527,N_26509,N_26446);
and U27528 (N_27528,N_26057,N_26812);
nand U27529 (N_27529,N_26089,N_25870);
nand U27530 (N_27530,N_27040,N_27497);
nor U27531 (N_27531,N_27259,N_25732);
and U27532 (N_27532,N_25217,N_27073);
xor U27533 (N_27533,N_27010,N_25147);
nor U27534 (N_27534,N_27075,N_26209);
nand U27535 (N_27535,N_25353,N_26162);
nor U27536 (N_27536,N_26444,N_27455);
and U27537 (N_27537,N_27071,N_26451);
nor U27538 (N_27538,N_27111,N_25306);
nand U27539 (N_27539,N_26230,N_26074);
nand U27540 (N_27540,N_25558,N_27325);
xnor U27541 (N_27541,N_25802,N_25390);
nor U27542 (N_27542,N_26537,N_26039);
nand U27543 (N_27543,N_25609,N_25058);
and U27544 (N_27544,N_26019,N_26711);
and U27545 (N_27545,N_26883,N_25179);
nor U27546 (N_27546,N_25133,N_27413);
nand U27547 (N_27547,N_26674,N_26925);
nor U27548 (N_27548,N_26053,N_25559);
nor U27549 (N_27549,N_26679,N_26440);
nand U27550 (N_27550,N_25830,N_25241);
nor U27551 (N_27551,N_25383,N_25520);
nand U27552 (N_27552,N_26646,N_25750);
and U27553 (N_27553,N_25478,N_25098);
and U27554 (N_27554,N_25529,N_27190);
and U27555 (N_27555,N_26953,N_26398);
or U27556 (N_27556,N_25017,N_25131);
nor U27557 (N_27557,N_26870,N_26041);
nor U27558 (N_27558,N_26803,N_25259);
or U27559 (N_27559,N_26058,N_26558);
nor U27560 (N_27560,N_26078,N_25978);
nand U27561 (N_27561,N_26347,N_27496);
nand U27562 (N_27562,N_25866,N_26849);
and U27563 (N_27563,N_26880,N_27238);
nand U27564 (N_27564,N_27202,N_25455);
nor U27565 (N_27565,N_25221,N_27113);
or U27566 (N_27566,N_26075,N_25984);
nor U27567 (N_27567,N_26283,N_25066);
or U27568 (N_27568,N_25186,N_25004);
nand U27569 (N_27569,N_26649,N_27285);
nand U27570 (N_27570,N_25521,N_26609);
nand U27571 (N_27571,N_26457,N_25351);
nor U27572 (N_27572,N_25144,N_25827);
or U27573 (N_27573,N_26865,N_26226);
and U27574 (N_27574,N_25785,N_26889);
and U27575 (N_27575,N_25352,N_26085);
or U27576 (N_27576,N_25676,N_26860);
nand U27577 (N_27577,N_26306,N_26102);
and U27578 (N_27578,N_26709,N_26343);
nand U27579 (N_27579,N_27481,N_26148);
nor U27580 (N_27580,N_26867,N_27335);
nand U27581 (N_27581,N_26521,N_27043);
nand U27582 (N_27582,N_26139,N_25831);
xnor U27583 (N_27583,N_27064,N_25825);
nand U27584 (N_27584,N_26678,N_25403);
nor U27585 (N_27585,N_26536,N_26620);
and U27586 (N_27586,N_26869,N_27129);
nand U27587 (N_27587,N_26023,N_26790);
and U27588 (N_27588,N_27205,N_26008);
or U27589 (N_27589,N_26723,N_27381);
or U27590 (N_27590,N_25591,N_27167);
xnor U27591 (N_27591,N_25649,N_25685);
nand U27592 (N_27592,N_27363,N_25770);
or U27593 (N_27593,N_27005,N_27119);
or U27594 (N_27594,N_25122,N_25929);
and U27595 (N_27595,N_26831,N_26055);
or U27596 (N_27596,N_25104,N_26696);
nand U27597 (N_27597,N_26730,N_25662);
and U27598 (N_27598,N_25965,N_25700);
nand U27599 (N_27599,N_26981,N_27244);
nor U27600 (N_27600,N_25300,N_26694);
or U27601 (N_27601,N_27240,N_25804);
nor U27602 (N_27602,N_27147,N_26338);
nor U27603 (N_27603,N_26616,N_25015);
nand U27604 (N_27604,N_25009,N_25795);
xnor U27605 (N_27605,N_25360,N_26836);
nor U27606 (N_27606,N_26647,N_26143);
nand U27607 (N_27607,N_26969,N_26888);
nor U27608 (N_27608,N_25669,N_25696);
or U27609 (N_27609,N_26610,N_25041);
nand U27610 (N_27610,N_25899,N_25222);
nor U27611 (N_27611,N_26847,N_26665);
or U27612 (N_27612,N_27380,N_26675);
nand U27613 (N_27613,N_25239,N_27269);
and U27614 (N_27614,N_27412,N_27107);
or U27615 (N_27615,N_26020,N_26307);
and U27616 (N_27616,N_27337,N_27112);
and U27617 (N_27617,N_25783,N_25923);
nand U27618 (N_27618,N_26123,N_25328);
nor U27619 (N_27619,N_26851,N_25840);
and U27620 (N_27620,N_25684,N_26204);
and U27621 (N_27621,N_25916,N_26192);
and U27622 (N_27622,N_26002,N_25069);
or U27623 (N_27623,N_26699,N_25173);
nand U27624 (N_27624,N_25742,N_25565);
and U27625 (N_27625,N_25140,N_27401);
or U27626 (N_27626,N_26517,N_25918);
xor U27627 (N_27627,N_25367,N_25238);
and U27628 (N_27628,N_26210,N_26167);
or U27629 (N_27629,N_26681,N_25093);
nor U27630 (N_27630,N_26223,N_25219);
nor U27631 (N_27631,N_27076,N_25100);
nor U27632 (N_27632,N_25151,N_25970);
and U27633 (N_27633,N_27477,N_25014);
xnor U27634 (N_27634,N_26030,N_26378);
nor U27635 (N_27635,N_25574,N_27308);
nand U27636 (N_27636,N_26915,N_26477);
or U27637 (N_27637,N_27025,N_27378);
nor U27638 (N_27638,N_25949,N_26467);
xor U27639 (N_27639,N_26268,N_26375);
nor U27640 (N_27640,N_26096,N_25698);
or U27641 (N_27641,N_26590,N_26025);
xor U27642 (N_27642,N_26181,N_26511);
nand U27643 (N_27643,N_26466,N_26939);
nor U27644 (N_27644,N_26919,N_27416);
nor U27645 (N_27645,N_25214,N_27163);
and U27646 (N_27646,N_26994,N_25958);
and U27647 (N_27647,N_27395,N_27011);
nand U27648 (N_27648,N_26772,N_27106);
nand U27649 (N_27649,N_27439,N_26195);
nand U27650 (N_27650,N_27144,N_26563);
or U27651 (N_27651,N_27003,N_26692);
nor U27652 (N_27652,N_26103,N_25052);
xnor U27653 (N_27653,N_25192,N_27309);
and U27654 (N_27654,N_25416,N_27383);
or U27655 (N_27655,N_25376,N_25717);
nand U27656 (N_27656,N_25769,N_26186);
nor U27657 (N_27657,N_26406,N_25433);
or U27658 (N_27658,N_25692,N_25070);
or U27659 (N_27659,N_26825,N_26234);
and U27660 (N_27660,N_25553,N_25767);
or U27661 (N_27661,N_26224,N_25138);
and U27662 (N_27662,N_26695,N_25939);
and U27663 (N_27663,N_27438,N_25975);
or U27664 (N_27664,N_26383,N_27022);
and U27665 (N_27665,N_26855,N_26056);
and U27666 (N_27666,N_25354,N_26534);
nand U27667 (N_27667,N_26505,N_26997);
and U27668 (N_27668,N_26069,N_25508);
or U27669 (N_27669,N_26878,N_25026);
nor U27670 (N_27670,N_26155,N_27149);
nand U27671 (N_27671,N_26449,N_25678);
or U27672 (N_27672,N_27448,N_25243);
and U27673 (N_27673,N_26564,N_27220);
and U27674 (N_27674,N_27152,N_26152);
or U27675 (N_27675,N_26807,N_25375);
nand U27676 (N_27676,N_26233,N_26542);
nor U27677 (N_27677,N_27387,N_27384);
and U27678 (N_27678,N_26009,N_25905);
and U27679 (N_27679,N_25385,N_27195);
and U27680 (N_27680,N_25321,N_25150);
nand U27681 (N_27681,N_26028,N_25666);
nor U27682 (N_27682,N_27030,N_27365);
or U27683 (N_27683,N_26172,N_25940);
nand U27684 (N_27684,N_26463,N_26781);
nor U27685 (N_27685,N_25183,N_25601);
nand U27686 (N_27686,N_26508,N_25090);
xor U27687 (N_27687,N_26729,N_25618);
and U27688 (N_27688,N_27334,N_26553);
nand U27689 (N_27689,N_27424,N_25616);
nor U27690 (N_27690,N_26461,N_25149);
nand U27691 (N_27691,N_26633,N_27026);
or U27692 (N_27692,N_26175,N_26635);
or U27693 (N_27693,N_25189,N_27160);
and U27694 (N_27694,N_27016,N_26289);
nor U27695 (N_27695,N_26297,N_26432);
nand U27696 (N_27696,N_25305,N_25648);
nand U27697 (N_27697,N_25109,N_25605);
or U27698 (N_27698,N_26965,N_26555);
nor U27699 (N_27699,N_27227,N_26073);
or U27700 (N_27700,N_26519,N_25155);
nand U27701 (N_27701,N_26125,N_27488);
nand U27702 (N_27702,N_26052,N_26854);
or U27703 (N_27703,N_26399,N_25293);
and U27704 (N_27704,N_26832,N_27045);
and U27705 (N_27705,N_25900,N_25278);
nand U27706 (N_27706,N_26197,N_26524);
nand U27707 (N_27707,N_26983,N_26876);
nand U27708 (N_27708,N_26262,N_26690);
nand U27709 (N_27709,N_25229,N_26967);
or U27710 (N_27710,N_26487,N_26607);
and U27711 (N_27711,N_26345,N_25382);
nor U27712 (N_27712,N_25462,N_27229);
nor U27713 (N_27713,N_25855,N_25668);
nand U27714 (N_27714,N_25702,N_27018);
nor U27715 (N_27715,N_27493,N_26473);
and U27716 (N_27716,N_27246,N_27223);
or U27717 (N_27717,N_26944,N_25612);
nand U27718 (N_27718,N_25693,N_26964);
nand U27719 (N_27719,N_25996,N_26042);
nand U27720 (N_27720,N_25697,N_25065);
and U27721 (N_27721,N_26650,N_27153);
or U27722 (N_27722,N_26110,N_26786);
or U27723 (N_27723,N_26744,N_25049);
or U27724 (N_27724,N_25937,N_25631);
nor U27725 (N_27725,N_26626,N_27459);
xor U27726 (N_27726,N_26095,N_25748);
and U27727 (N_27727,N_26159,N_25081);
or U27728 (N_27728,N_25424,N_27457);
nor U27729 (N_27729,N_25790,N_25022);
and U27730 (N_27730,N_26193,N_25835);
nor U27731 (N_27731,N_25661,N_26659);
and U27732 (N_27732,N_26957,N_27362);
or U27733 (N_27733,N_26951,N_27186);
nor U27734 (N_27734,N_26992,N_25195);
nand U27735 (N_27735,N_25772,N_26504);
nand U27736 (N_27736,N_26066,N_26545);
or U27737 (N_27737,N_26546,N_25288);
and U27738 (N_27738,N_26923,N_27339);
or U27739 (N_27739,N_26707,N_27065);
and U27740 (N_27740,N_25055,N_25722);
nor U27741 (N_27741,N_25613,N_25419);
nand U27742 (N_27742,N_25818,N_26294);
nor U27743 (N_27743,N_25815,N_25811);
nor U27744 (N_27744,N_25469,N_25549);
nor U27745 (N_27745,N_25610,N_26111);
nand U27746 (N_27746,N_25792,N_25522);
or U27747 (N_27747,N_25340,N_26092);
and U27748 (N_27748,N_25747,N_26879);
xor U27749 (N_27749,N_25930,N_26421);
nor U27750 (N_27750,N_26845,N_27456);
or U27751 (N_27751,N_26079,N_25161);
nand U27752 (N_27752,N_26701,N_25977);
and U27753 (N_27753,N_25944,N_25429);
and U27754 (N_27754,N_27303,N_25235);
or U27755 (N_27755,N_26912,N_25551);
or U27756 (N_27756,N_27352,N_27399);
or U27757 (N_27757,N_25757,N_26672);
nand U27758 (N_27758,N_26483,N_27330);
nand U27759 (N_27759,N_25345,N_25743);
xor U27760 (N_27760,N_25226,N_27272);
or U27761 (N_27761,N_25181,N_25881);
nand U27762 (N_27762,N_27027,N_25803);
nor U27763 (N_27763,N_27080,N_25600);
or U27764 (N_27764,N_25200,N_26918);
nor U27765 (N_27765,N_25868,N_25848);
xor U27766 (N_27766,N_26570,N_26379);
nand U27767 (N_27767,N_27154,N_27141);
and U27768 (N_27768,N_27475,N_26410);
nor U27769 (N_27769,N_27197,N_26308);
nor U27770 (N_27770,N_26285,N_25483);
nor U27771 (N_27771,N_25983,N_26314);
nor U27772 (N_27772,N_25587,N_27126);
nand U27773 (N_27773,N_27097,N_26251);
nand U27774 (N_27774,N_26751,N_25725);
xnor U27775 (N_27775,N_26207,N_27023);
nand U27776 (N_27776,N_25639,N_27069);
and U27777 (N_27777,N_25184,N_27077);
nor U27778 (N_27778,N_26720,N_25442);
and U27779 (N_27779,N_26991,N_26010);
or U27780 (N_27780,N_26084,N_25799);
xor U27781 (N_27781,N_27495,N_26503);
nand U27782 (N_27782,N_26911,N_26902);
nor U27783 (N_27783,N_25249,N_26284);
nor U27784 (N_27784,N_26179,N_25525);
and U27785 (N_27785,N_25957,N_25490);
or U27786 (N_27786,N_26012,N_26921);
and U27787 (N_27787,N_27301,N_26138);
xor U27788 (N_27788,N_26376,N_26974);
nor U27789 (N_27789,N_26024,N_25879);
nand U27790 (N_27790,N_26280,N_27172);
and U27791 (N_27791,N_26121,N_26022);
xnor U27792 (N_27792,N_26459,N_27458);
nor U27793 (N_27793,N_27215,N_25486);
and U27794 (N_27794,N_27464,N_27222);
xor U27795 (N_27795,N_25739,N_25458);
and U27796 (N_27796,N_26506,N_25117);
or U27797 (N_27797,N_25793,N_27212);
nor U27798 (N_27798,N_27135,N_26360);
nand U27799 (N_27799,N_26330,N_26083);
nor U27800 (N_27800,N_26265,N_27347);
or U27801 (N_27801,N_25808,N_25006);
xnor U27802 (N_27802,N_25956,N_25637);
nor U27803 (N_27803,N_27425,N_25524);
and U27804 (N_27804,N_27288,N_25324);
xor U27805 (N_27805,N_25244,N_26702);
nor U27806 (N_27806,N_25057,N_27148);
nor U27807 (N_27807,N_25401,N_25096);
nand U27808 (N_27808,N_27157,N_25079);
nand U27809 (N_27809,N_26060,N_26898);
nor U27810 (N_27810,N_26061,N_27391);
and U27811 (N_27811,N_27093,N_27376);
nand U27812 (N_27812,N_26541,N_26523);
nor U27813 (N_27813,N_25755,N_26780);
nand U27814 (N_27814,N_25913,N_25400);
xor U27815 (N_27815,N_26250,N_25987);
nor U27816 (N_27816,N_27498,N_25745);
nor U27817 (N_27817,N_25157,N_25498);
or U27818 (N_27818,N_26049,N_26894);
or U27819 (N_27819,N_25509,N_26628);
xnor U27820 (N_27820,N_26493,N_26557);
xor U27821 (N_27821,N_27235,N_25168);
and U27822 (N_27822,N_26201,N_26257);
nand U27823 (N_27823,N_26496,N_25846);
and U27824 (N_27824,N_25332,N_25990);
nor U27825 (N_27825,N_26312,N_27367);
or U27826 (N_27826,N_25634,N_27290);
nand U27827 (N_27827,N_26819,N_25664);
nand U27828 (N_27828,N_25263,N_26995);
and U27829 (N_27829,N_25331,N_26782);
nand U27830 (N_27830,N_25407,N_26535);
or U27831 (N_27831,N_25906,N_26458);
nor U27832 (N_27832,N_25843,N_26352);
nand U27833 (N_27833,N_27315,N_26722);
xor U27834 (N_27834,N_25450,N_25223);
nand U27835 (N_27835,N_25550,N_27209);
xor U27836 (N_27836,N_26342,N_25632);
nor U27837 (N_27837,N_25643,N_26666);
nand U27838 (N_27838,N_26403,N_27258);
nand U27839 (N_27839,N_26673,N_26853);
xor U27840 (N_27840,N_27094,N_25125);
nand U27841 (N_27841,N_27241,N_25689);
or U27842 (N_27842,N_25933,N_26724);
and U27843 (N_27843,N_27444,N_25560);
nor U27844 (N_27844,N_26833,N_26104);
or U27845 (N_27845,N_27369,N_25210);
and U27846 (N_27846,N_26177,N_25164);
or U27847 (N_27847,N_25051,N_25557);
or U27848 (N_27848,N_26326,N_25464);
and U27849 (N_27849,N_27035,N_25163);
and U27850 (N_27850,N_25256,N_25935);
and U27851 (N_27851,N_27017,N_25660);
nor U27852 (N_27852,N_25021,N_26048);
or U27853 (N_27853,N_27121,N_25343);
and U27854 (N_27854,N_27450,N_25277);
or U27855 (N_27855,N_25736,N_27390);
nor U27856 (N_27856,N_27115,N_26425);
nor U27857 (N_27857,N_27291,N_26683);
and U27858 (N_27858,N_26435,N_25650);
nor U27859 (N_27859,N_27392,N_25759);
or U27860 (N_27860,N_25279,N_26515);
and U27861 (N_27861,N_26336,N_26282);
and U27862 (N_27862,N_25703,N_26742);
nor U27863 (N_27863,N_25665,N_25007);
and U27864 (N_27864,N_25396,N_25744);
and U27865 (N_27865,N_25280,N_25493);
and U27866 (N_27866,N_25175,N_26968);
or U27867 (N_27867,N_26036,N_26154);
xnor U27868 (N_27868,N_25567,N_26706);
or U27869 (N_27869,N_25115,N_25029);
or U27870 (N_27870,N_27299,N_26811);
nand U27871 (N_27871,N_25129,N_25726);
nand U27872 (N_27872,N_27417,N_25106);
nand U27873 (N_27873,N_27029,N_25680);
nor U27874 (N_27874,N_25365,N_25907);
or U27875 (N_27875,N_27004,N_27155);
and U27876 (N_27876,N_25771,N_26959);
or U27877 (N_27877,N_25452,N_26934);
nor U27878 (N_27878,N_26164,N_25814);
nand U27879 (N_27879,N_25422,N_25585);
and U27880 (N_27880,N_26237,N_25655);
nand U27881 (N_27881,N_25874,N_27254);
nor U27882 (N_27882,N_26941,N_25152);
nor U27883 (N_27883,N_26745,N_25087);
and U27884 (N_27884,N_27333,N_26478);
and U27885 (N_27885,N_25046,N_26612);
nand U27886 (N_27886,N_27159,N_25399);
nand U27887 (N_27887,N_26916,N_25976);
nand U27888 (N_27888,N_26333,N_27312);
nor U27889 (N_27889,N_27420,N_27371);
or U27890 (N_27890,N_25054,N_25539);
nor U27891 (N_27891,N_27445,N_26598);
or U27892 (N_27892,N_25145,N_25171);
nor U27893 (N_27893,N_25974,N_27046);
xor U27894 (N_27894,N_25690,N_25528);
or U27895 (N_27895,N_27386,N_25798);
nand U27896 (N_27896,N_25889,N_25341);
and U27897 (N_27897,N_25311,N_25962);
or U27898 (N_27898,N_26676,N_26584);
and U27899 (N_27899,N_27338,N_27364);
or U27900 (N_27900,N_25800,N_25507);
nor U27901 (N_27901,N_27421,N_26595);
nor U27902 (N_27902,N_25089,N_26267);
nor U27903 (N_27903,N_26931,N_25543);
nor U27904 (N_27904,N_27185,N_25912);
or U27905 (N_27905,N_27418,N_27104);
and U27906 (N_27906,N_25356,N_26539);
nor U27907 (N_27907,N_26947,N_27377);
nor U27908 (N_27908,N_26486,N_26212);
nand U27909 (N_27909,N_25651,N_27060);
and U27910 (N_27910,N_25854,N_26391);
or U27911 (N_27911,N_26263,N_26047);
or U27912 (N_27912,N_26452,N_26928);
or U27913 (N_27913,N_26339,N_25514);
nor U27914 (N_27914,N_26805,N_26731);
or U27915 (N_27915,N_26841,N_25768);
nor U27916 (N_27916,N_27317,N_26591);
xnor U27917 (N_27917,N_27012,N_26369);
or U27918 (N_27918,N_26313,N_25126);
or U27919 (N_27919,N_25130,N_25578);
and U27920 (N_27920,N_25882,N_25418);
nand U27921 (N_27921,N_25720,N_27368);
nand U27922 (N_27922,N_25504,N_26160);
nand U27923 (N_27923,N_26644,N_26188);
xor U27924 (N_27924,N_26604,N_27174);
nor U27925 (N_27925,N_26147,N_26419);
nand U27926 (N_27926,N_25146,N_25707);
nand U27927 (N_27927,N_27162,N_25833);
and U27928 (N_27928,N_26259,N_27085);
and U27929 (N_27929,N_27008,N_26013);
nand U27930 (N_27930,N_26641,N_25968);
or U27931 (N_27931,N_27007,N_25517);
and U27932 (N_27932,N_26126,N_27454);
xor U27933 (N_27933,N_27161,N_26499);
nand U27934 (N_27934,N_26543,N_26815);
nand U27935 (N_27935,N_26623,N_25586);
and U27936 (N_27936,N_26163,N_25209);
nor U27937 (N_27937,N_27319,N_25713);
and U27938 (N_27938,N_27471,N_25705);
nand U27939 (N_27939,N_26926,N_27078);
and U27940 (N_27940,N_27137,N_27382);
nand U27941 (N_27941,N_25158,N_27201);
or U27942 (N_27942,N_25088,N_25516);
or U27943 (N_27943,N_25512,N_26323);
and U27944 (N_27944,N_25193,N_26838);
xor U27945 (N_27945,N_25472,N_26725);
or U27946 (N_27946,N_26513,N_26475);
nor U27947 (N_27947,N_25487,N_26642);
xnor U27948 (N_27948,N_25315,N_25494);
nand U27949 (N_27949,N_27116,N_25723);
or U27950 (N_27950,N_26462,N_25875);
and U27951 (N_27951,N_25606,N_25495);
and U27952 (N_27952,N_25603,N_25503);
nor U27953 (N_27953,N_25820,N_25178);
or U27954 (N_27954,N_25894,N_27452);
nand U27955 (N_27955,N_26287,N_26861);
and U27956 (N_27956,N_27021,N_26528);
or U27957 (N_27957,N_27020,N_25828);
or U27958 (N_27958,N_25880,N_26003);
nor U27959 (N_27959,N_26990,N_27388);
nand U27960 (N_27960,N_26761,N_26043);
and U27961 (N_27961,N_26522,N_27287);
nor U27962 (N_27962,N_25640,N_27210);
nand U27963 (N_27963,N_25290,N_25064);
xor U27964 (N_27964,N_26905,N_25479);
nor U27965 (N_27965,N_25296,N_25947);
nand U27966 (N_27966,N_27143,N_27292);
or U27967 (N_27967,N_26773,N_27042);
xnor U27968 (N_27968,N_26859,N_26655);
and U27969 (N_27969,N_26949,N_27427);
nor U27970 (N_27970,N_27203,N_26520);
xor U27971 (N_27971,N_27298,N_25439);
xor U27972 (N_27972,N_27015,N_25220);
xor U27973 (N_27973,N_27407,N_27473);
and U27974 (N_27974,N_26667,N_26796);
or U27975 (N_27975,N_27499,N_27358);
or U27976 (N_27976,N_25991,N_26261);
xor U27977 (N_27977,N_26622,N_27440);
and U27978 (N_27978,N_26489,N_25656);
nand U27979 (N_27979,N_26100,N_25903);
and U27980 (N_27980,N_26789,N_26600);
and U27981 (N_27981,N_25188,N_25839);
or U27982 (N_27982,N_27239,N_25056);
and U27983 (N_27983,N_26914,N_25727);
nand U27984 (N_27984,N_26472,N_27173);
nand U27985 (N_27985,N_26442,N_25541);
or U27986 (N_27986,N_27127,N_26388);
nor U27987 (N_27987,N_26910,N_25598);
or U27988 (N_27988,N_25538,N_26412);
or U27989 (N_27989,N_25368,N_26245);
and U27990 (N_27990,N_26718,N_27177);
or U27991 (N_27991,N_27273,N_26443);
nand U27992 (N_27992,N_25646,N_26029);
xor U27993 (N_27993,N_27446,N_27221);
nor U27994 (N_27994,N_26937,N_25819);
xnor U27995 (N_27995,N_26275,N_25813);
or U27996 (N_27996,N_25001,N_26743);
or U27997 (N_27997,N_25294,N_26279);
nand U27998 (N_27998,N_25170,N_26037);
or U27999 (N_27999,N_26407,N_25533);
nand U28000 (N_28000,N_25682,N_26728);
nor U28001 (N_28001,N_25670,N_25201);
xnor U28002 (N_28002,N_27125,N_25316);
nor U28003 (N_28003,N_26206,N_25274);
nand U28004 (N_28004,N_25505,N_25110);
nand U28005 (N_28005,N_26219,N_25691);
or U28006 (N_28006,N_25092,N_25298);
and U28007 (N_28007,N_25071,N_25863);
or U28008 (N_28008,N_26437,N_26404);
or U28009 (N_28009,N_25295,N_27207);
or U28010 (N_28010,N_27271,N_27061);
or U28011 (N_28011,N_27048,N_27468);
nand U28012 (N_28012,N_25791,N_26215);
nand U28013 (N_28013,N_25053,N_26005);
nand U28014 (N_28014,N_26018,N_26180);
nand U28015 (N_28015,N_25208,N_26844);
or U28016 (N_28016,N_25677,N_25191);
nor U28017 (N_28017,N_27281,N_25236);
xor U28018 (N_28018,N_25806,N_26054);
and U28019 (N_28019,N_26300,N_26821);
or U28020 (N_28020,N_25420,N_25451);
nor U28021 (N_28021,N_26813,N_27492);
nor U28022 (N_28022,N_25108,N_27245);
nor U28023 (N_28023,N_27411,N_25265);
xnor U28024 (N_28024,N_25169,N_26006);
or U28025 (N_28025,N_25119,N_27136);
nor U28026 (N_28026,N_26611,N_25363);
and U28027 (N_28027,N_26903,N_26448);
and U28028 (N_28028,N_25925,N_26824);
nor U28029 (N_28029,N_26027,N_27057);
or U28030 (N_28030,N_26454,N_26579);
and U28031 (N_28031,N_27140,N_26080);
or U28032 (N_28032,N_26606,N_26450);
nor U28033 (N_28033,N_26225,N_27165);
and U28034 (N_28034,N_25604,N_26183);
and U28035 (N_28035,N_25728,N_26804);
or U28036 (N_28036,N_26808,N_25091);
or U28037 (N_28037,N_25409,N_26229);
nor U28038 (N_28038,N_25499,N_26277);
nor U28039 (N_28039,N_25101,N_26319);
nand U28040 (N_28040,N_26630,N_25000);
or U28041 (N_28041,N_27443,N_27479);
or U28042 (N_28042,N_25834,N_25774);
xnor U28043 (N_28043,N_27171,N_27070);
nor U28044 (N_28044,N_27139,N_27489);
and U28045 (N_28045,N_27176,N_25386);
or U28046 (N_28046,N_26090,N_27250);
nor U28047 (N_28047,N_27055,N_25877);
nor U28048 (N_28048,N_26787,N_25132);
and U28049 (N_28049,N_26405,N_25459);
nor U28050 (N_28050,N_25961,N_25061);
or U28051 (N_28051,N_26132,N_26114);
nand U28052 (N_28052,N_26059,N_27187);
or U28053 (N_28053,N_26216,N_26569);
nor U28054 (N_28054,N_26989,N_26507);
nand U28055 (N_28055,N_27311,N_26136);
xor U28056 (N_28056,N_25438,N_25440);
nand U28057 (N_28057,N_27437,N_25596);
nand U28058 (N_28058,N_26045,N_27354);
or U28059 (N_28059,N_26906,N_27214);
or U28060 (N_28060,N_25540,N_27253);
and U28061 (N_28061,N_26882,N_27331);
nand U28062 (N_28062,N_27019,N_25919);
xor U28063 (N_28063,N_26411,N_27435);
xnor U28064 (N_28064,N_26488,N_27058);
nor U28065 (N_28065,N_26638,N_26762);
and U28066 (N_28066,N_26331,N_25952);
and U28067 (N_28067,N_26007,N_25807);
nor U28068 (N_28068,N_25625,N_25139);
or U28069 (N_28069,N_26434,N_26748);
nand U28070 (N_28070,N_26130,N_25456);
nand U28071 (N_28071,N_27083,N_25635);
and U28072 (N_28072,N_25207,N_26298);
or U28073 (N_28073,N_26252,N_27373);
or U28074 (N_28074,N_26619,N_25788);
or U28075 (N_28075,N_27079,N_25060);
and U28076 (N_28076,N_27101,N_25932);
nand U28077 (N_28077,N_25724,N_26149);
or U28078 (N_28078,N_25485,N_26198);
or U28079 (N_28079,N_27396,N_27249);
or U28080 (N_28080,N_25273,N_25018);
and U28081 (N_28081,N_26337,N_26169);
nor U28082 (N_28082,N_26494,N_27423);
or U28083 (N_28083,N_25915,N_26241);
nor U28084 (N_28084,N_26389,N_27326);
xnor U28085 (N_28085,N_26247,N_25911);
xnor U28086 (N_28086,N_27039,N_26754);
nor U28087 (N_28087,N_26671,N_26658);
and U28088 (N_28088,N_26397,N_27252);
and U28089 (N_28089,N_26617,N_25909);
nand U28090 (N_28090,N_27138,N_26712);
nand U28091 (N_28091,N_26884,N_27179);
and U28092 (N_28092,N_26791,N_26713);
or U28093 (N_28093,N_26386,N_26862);
xnor U28094 (N_28094,N_25715,N_25850);
or U28095 (N_28095,N_25513,N_26354);
nor U28096 (N_28096,N_26952,N_26122);
and U28097 (N_28097,N_25302,N_26295);
and U28098 (N_28098,N_27117,N_26415);
or U28099 (N_28099,N_26174,N_26943);
or U28100 (N_28100,N_25237,N_26350);
nor U28101 (N_28101,N_25372,N_26064);
xnor U28102 (N_28102,N_25449,N_26501);
and U28103 (N_28103,N_27120,N_25257);
nor U28104 (N_28104,N_25297,N_26698);
nand U28105 (N_28105,N_27404,N_26240);
xor U28106 (N_28106,N_25730,N_26829);
nor U28107 (N_28107,N_25039,N_26909);
xor U28108 (N_28108,N_25829,N_25240);
or U28109 (N_28109,N_27282,N_26986);
xor U28110 (N_28110,N_25753,N_25474);
nand U28111 (N_28111,N_25627,N_25571);
xnor U28112 (N_28112,N_25213,N_25920);
or U28113 (N_28113,N_26191,N_25355);
nor U28114 (N_28114,N_25225,N_25335);
and U28115 (N_28115,N_26077,N_25897);
or U28116 (N_28116,N_26236,N_25534);
and U28117 (N_28117,N_25361,N_25251);
and U28118 (N_28118,N_26286,N_26260);
nor U28119 (N_28119,N_27099,N_25142);
nor U28120 (N_28120,N_27297,N_25285);
and U28121 (N_28121,N_25038,N_26317);
nand U28122 (N_28122,N_26438,N_25579);
xnor U28123 (N_28123,N_25624,N_25358);
and U28124 (N_28124,N_25476,N_25084);
nor U28125 (N_28125,N_25141,N_25037);
and U28126 (N_28126,N_27068,N_25763);
or U28127 (N_28127,N_25137,N_27268);
xnor U28128 (N_28128,N_25105,N_27262);
nand U28129 (N_28129,N_26278,N_25518);
xor U28130 (N_28130,N_27118,N_27478);
nand U28131 (N_28131,N_25412,N_26227);
and U28132 (N_28132,N_25761,N_25841);
nand U28133 (N_28133,N_26429,N_27402);
nor U28134 (N_28134,N_25346,N_25135);
and U28135 (N_28135,N_26341,N_27289);
nor U28136 (N_28136,N_25766,N_25542);
and U28137 (N_28137,N_26106,N_26817);
and U28138 (N_28138,N_26777,N_25687);
nand U28139 (N_28139,N_25711,N_26474);
xor U28140 (N_28140,N_26857,N_27049);
and U28141 (N_28141,N_26645,N_25357);
xnor U28142 (N_28142,N_26608,N_26750);
and U28143 (N_28143,N_25599,N_26827);
and U28144 (N_28144,N_26717,N_25568);
and U28145 (N_28145,N_25369,N_26495);
nor U28146 (N_28146,N_25989,N_27211);
nand U28147 (N_28147,N_25094,N_25709);
or U28148 (N_28148,N_26481,N_26413);
nor U28149 (N_28149,N_25746,N_27096);
nor U28150 (N_28150,N_26086,N_25716);
and U28151 (N_28151,N_25113,N_25447);
and U28152 (N_28152,N_27277,N_25547);
and U28153 (N_28153,N_27409,N_26779);
nand U28154 (N_28154,N_26356,N_25269);
and U28155 (N_28155,N_25307,N_25589);
nand U28156 (N_28156,N_26291,N_26213);
and U28157 (N_28157,N_25338,N_25837);
and U28158 (N_28158,N_25378,N_25329);
nand U28159 (N_28159,N_26116,N_27466);
nand U28160 (N_28160,N_25555,N_26361);
and U28161 (N_28161,N_25569,N_26254);
xor U28162 (N_28162,N_25394,N_26714);
and U28163 (N_28163,N_26828,N_25496);
nand U28164 (N_28164,N_25805,N_26150);
xnor U28165 (N_28165,N_25592,N_25588);
nor U28166 (N_28166,N_27002,N_27188);
xnor U28167 (N_28167,N_27124,N_26776);
nand U28168 (N_28168,N_26741,N_26593);
nand U28169 (N_28169,N_25410,N_25878);
and U28170 (N_28170,N_27230,N_25924);
or U28171 (N_28171,N_27491,N_27310);
nand U28172 (N_28172,N_27359,N_26559);
nor U28173 (N_28173,N_27196,N_26001);
nor U28174 (N_28174,N_26476,N_27305);
nand U28175 (N_28175,N_26357,N_26614);
and U28176 (N_28176,N_26460,N_25373);
nor U28177 (N_28177,N_27433,N_25914);
nand U28178 (N_28178,N_25276,N_25426);
and U28179 (N_28179,N_25941,N_26134);
nor U28180 (N_28180,N_25180,N_26296);
nor U28181 (N_28181,N_26266,N_26580);
nand U28182 (N_28182,N_27322,N_27072);
and U28183 (N_28183,N_25809,N_25245);
nor U28184 (N_28184,N_25844,N_25659);
and U28185 (N_28185,N_27164,N_25415);
and U28186 (N_28186,N_25461,N_26321);
nor U28187 (N_28187,N_25873,N_26141);
nand U28188 (N_28188,N_26129,N_25333);
or U28189 (N_28189,N_25786,N_26705);
xor U28190 (N_28190,N_27342,N_26070);
nand U28191 (N_28191,N_25118,N_25515);
nand U28192 (N_28192,N_26034,N_26881);
and U28193 (N_28193,N_26984,N_27430);
nor U28194 (N_28194,N_26492,N_26453);
xnor U28195 (N_28195,N_25030,N_26302);
nand U28196 (N_28196,N_26663,N_26011);
nor U28197 (N_28197,N_25816,N_26325);
xnor U28198 (N_28198,N_25537,N_26830);
xnor U28199 (N_28199,N_27441,N_27200);
nand U28200 (N_28200,N_25773,N_26999);
or U28201 (N_28201,N_25563,N_26098);
nor U28202 (N_28202,N_27357,N_25154);
xnor U28203 (N_28203,N_26834,N_25040);
xor U28204 (N_28204,N_25619,N_27356);
or U28205 (N_28205,N_27476,N_27234);
and U28206 (N_28206,N_26072,N_25938);
nor U28207 (N_28207,N_25561,N_25582);
and U28208 (N_28208,N_26768,N_26715);
nor U28209 (N_28209,N_26568,N_25886);
or U28210 (N_28210,N_25999,N_27132);
nor U28211 (N_28211,N_25111,N_25421);
or U28212 (N_28212,N_26238,N_27224);
or U28213 (N_28213,N_25362,N_26792);
nand U28214 (N_28214,N_25308,N_25359);
or U28215 (N_28215,N_25570,N_26640);
xnor U28216 (N_28216,N_26549,N_25206);
nand U28217 (N_28217,N_25644,N_25615);
and U28218 (N_28218,N_26581,N_26566);
nor U28219 (N_28219,N_26890,N_26362);
or U28220 (N_28220,N_27095,N_25019);
nand U28221 (N_28221,N_25871,N_26954);
xnor U28222 (N_28222,N_27329,N_26170);
nor U28223 (N_28223,N_26107,N_25260);
or U28224 (N_28224,N_25381,N_25950);
xor U28225 (N_28225,N_27434,N_25630);
nand U28226 (N_28226,N_26794,N_26372);
nor U28227 (N_28227,N_26371,N_25322);
and U28228 (N_28228,N_25859,N_25044);
and U28229 (N_28229,N_27263,N_26797);
and U28230 (N_28230,N_26735,N_26178);
and U28231 (N_28231,N_25752,N_25951);
and U28232 (N_28232,N_25224,N_27323);
xnor U28233 (N_28233,N_27090,N_25282);
or U28234 (N_28234,N_25035,N_27324);
nor U28235 (N_28235,N_26394,N_25674);
nand U28236 (N_28236,N_25325,N_25284);
xnor U28237 (N_28237,N_26863,N_25444);
xnor U28238 (N_28238,N_26597,N_25888);
or U28239 (N_28239,N_25162,N_26571);
nand U28240 (N_28240,N_26746,N_25303);
and U28241 (N_28241,N_25212,N_26526);
nand U28242 (N_28242,N_25211,N_25202);
or U28243 (N_28243,N_27130,N_27264);
or U28244 (N_28244,N_27379,N_25901);
nor U28245 (N_28245,N_27472,N_25074);
or U28246 (N_28246,N_25153,N_26393);
and U28247 (N_28247,N_26774,N_27100);
nor U28248 (N_28248,N_25165,N_27054);
and U28249 (N_28249,N_25733,N_25320);
or U28250 (N_28250,N_26756,N_27302);
or U28251 (N_28251,N_25611,N_27108);
nor U28252 (N_28252,N_25121,N_25836);
or U28253 (N_28253,N_26367,N_26359);
nor U28254 (N_28254,N_27233,N_26166);
nor U28255 (N_28255,N_26482,N_26933);
and U28256 (N_28256,N_25286,N_25706);
and U28257 (N_28257,N_27320,N_25292);
nor U28258 (N_28258,N_25718,N_25291);
and U28259 (N_28259,N_25077,N_26977);
xor U28260 (N_28260,N_26242,N_27088);
nand U28261 (N_28261,N_26349,N_26806);
and U28262 (N_28262,N_27484,N_26544);
and U28263 (N_28263,N_25960,N_26763);
nor U28264 (N_28264,N_27236,N_26930);
nand U28265 (N_28265,N_26929,N_26118);
or U28266 (N_28266,N_26648,N_25337);
and U28267 (N_28267,N_26874,N_25327);
nand U28268 (N_28268,N_26087,N_27442);
nor U28269 (N_28269,N_26875,N_25156);
nor U28270 (N_28270,N_25010,N_25782);
nor U28271 (N_28271,N_26396,N_26015);
or U28272 (N_28272,N_25166,N_25258);
and U28273 (N_28273,N_25086,N_25016);
nand U28274 (N_28274,N_26334,N_27405);
nand U28275 (N_28275,N_25980,N_26439);
or U28276 (N_28276,N_26866,N_26993);
nor U28277 (N_28277,N_26305,N_26656);
nand U28278 (N_28278,N_25027,N_26533);
xor U28279 (N_28279,N_26365,N_25261);
and U28280 (N_28280,N_27133,N_25872);
nand U28281 (N_28281,N_27218,N_27013);
nand U28282 (N_28282,N_27490,N_25078);
or U28283 (N_28283,N_25134,N_27066);
nand U28284 (N_28284,N_26137,N_25764);
nor U28285 (N_28285,N_25842,N_26747);
or U28286 (N_28286,N_25176,N_25203);
nand U28287 (N_28287,N_27461,N_25642);
nand U28288 (N_28288,N_26004,N_27170);
or U28289 (N_28289,N_26316,N_25740);
nor U28290 (N_28290,N_27295,N_26689);
or U28291 (N_28291,N_26471,N_25546);
xor U28292 (N_28292,N_26366,N_25481);
nor U28293 (N_28293,N_27082,N_25851);
or U28294 (N_28294,N_26063,N_26998);
nand U28295 (N_28295,N_25366,N_25187);
or U28296 (N_28296,N_27184,N_25460);
and U28297 (N_28297,N_27494,N_26823);
nor U28298 (N_28298,N_25266,N_25112);
nand U28299 (N_28299,N_26738,N_27074);
or U28300 (N_28300,N_26962,N_26900);
or U28301 (N_28301,N_25160,N_26465);
and U28302 (N_28302,N_25034,N_26531);
or U28303 (N_28303,N_25020,N_27198);
or U28304 (N_28304,N_26344,N_25227);
nand U28305 (N_28305,N_27463,N_26670);
or U28306 (N_28306,N_25675,N_25969);
or U28307 (N_28307,N_27398,N_27276);
xnor U28308 (N_28308,N_25233,N_26502);
and U28309 (N_28309,N_26329,N_26382);
xor U28310 (N_28310,N_26202,N_26956);
nor U28311 (N_28311,N_26826,N_25908);
and U28312 (N_28312,N_26311,N_25673);
and U28313 (N_28313,N_26627,N_27428);
nand U28314 (N_28314,N_26044,N_25847);
nor U28315 (N_28315,N_25527,N_26335);
nor U28316 (N_28316,N_27260,N_27346);
nand U28317 (N_28317,N_26661,N_26755);
and U28318 (N_28318,N_27123,N_26117);
nor U28319 (N_28319,N_26554,N_25701);
and U28320 (N_28320,N_26920,N_26127);
and U28321 (N_28321,N_26271,N_25392);
nor U28322 (N_28322,N_25047,N_26583);
nand U28323 (N_28323,N_26447,N_26892);
and U28324 (N_28324,N_26248,N_25002);
and U28325 (N_28325,N_25347,N_25653);
and U28326 (N_28326,N_27178,N_27393);
or U28327 (N_28327,N_26436,N_25411);
xor U28328 (N_28328,N_25636,N_26408);
or U28329 (N_28329,N_26693,N_25580);
or U28330 (N_28330,N_26605,N_25986);
xor U28331 (N_28331,N_26076,N_27014);
nor U28332 (N_28332,N_27348,N_26189);
or U28333 (N_28333,N_26514,N_25120);
nand U28334 (N_28334,N_26769,N_25003);
nor U28335 (N_28335,N_26046,N_26799);
or U28336 (N_28336,N_25095,N_26491);
nor U28337 (N_28337,N_25681,N_27208);
xor U28338 (N_28338,N_26120,N_26196);
nor U28339 (N_28339,N_26101,N_26686);
xor U28340 (N_28340,N_25955,N_27314);
or U28341 (N_28341,N_25910,N_26156);
nand U28342 (N_28342,N_27375,N_25374);
and U28343 (N_28343,N_27266,N_27256);
or U28344 (N_28344,N_26837,N_26340);
or U28345 (N_28345,N_27336,N_25314);
nor U28346 (N_28346,N_26239,N_25342);
and U28347 (N_28347,N_25641,N_26441);
or U28348 (N_28348,N_27327,N_25398);
nand U28349 (N_28349,N_26573,N_26199);
and U28350 (N_28350,N_26691,N_25289);
nor U28351 (N_28351,N_27483,N_25556);
xnor U28352 (N_28352,N_26708,N_26348);
nor U28353 (N_28353,N_26846,N_26140);
nand U28354 (N_28354,N_26802,N_25622);
nor U28355 (N_28355,N_26128,N_25234);
and U28356 (N_28356,N_26414,N_26232);
nor U28357 (N_28357,N_27032,N_25988);
nand U28358 (N_28358,N_26540,N_25349);
nor U28359 (N_28359,N_26469,N_25593);
nand U28360 (N_28360,N_26732,N_27086);
or U28361 (N_28361,N_25059,N_25794);
or U28362 (N_28362,N_27316,N_25845);
nand U28363 (N_28363,N_26327,N_26822);
or U28364 (N_28364,N_25796,N_25312);
or U28365 (N_28365,N_26653,N_26293);
or U28366 (N_28366,N_27033,N_25050);
nand U28367 (N_28367,N_25067,N_26498);
and U28368 (N_28368,N_25789,N_25934);
xnor U28369 (N_28369,N_25127,N_26778);
nor U28370 (N_28370,N_25575,N_25511);
nand U28371 (N_28371,N_26108,N_25397);
nor U28372 (N_28372,N_27414,N_25250);
nand U28373 (N_28373,N_26624,N_26917);
nor U28374 (N_28374,N_25694,N_25590);
or U28375 (N_28375,N_25281,N_27374);
or U28376 (N_28376,N_27361,N_27265);
and U28377 (N_28377,N_26538,N_25484);
and U28378 (N_28378,N_26757,N_26244);
xor U28379 (N_28379,N_25272,N_26996);
nor U28380 (N_28380,N_25942,N_26637);
nand U28381 (N_28381,N_25552,N_25425);
and U28382 (N_28382,N_25594,N_26530);
or U28383 (N_28383,N_26556,N_26801);
nor U28384 (N_28384,N_26795,N_25645);
nand U28385 (N_28385,N_25391,N_26840);
and U28386 (N_28386,N_26592,N_25028);
nor U28387 (N_28387,N_26470,N_26016);
and U28388 (N_28388,N_27408,N_25762);
xnor U28389 (N_28389,N_26243,N_26490);
nand U28390 (N_28390,N_26987,N_26328);
nand U28391 (N_28391,N_27394,N_25023);
and U28392 (N_28392,N_26272,N_27300);
nor U28393 (N_28393,N_25012,N_27403);
nor U28394 (N_28394,N_26680,N_26766);
nand U28395 (N_28395,N_25262,N_26292);
nand U28396 (N_28396,N_26818,N_27056);
or U28397 (N_28397,N_25993,N_25196);
or U28398 (N_28398,N_25657,N_25228);
nand U28399 (N_28399,N_27397,N_25042);
and U28400 (N_28400,N_26835,N_26173);
nand U28401 (N_28401,N_25780,N_26235);
and U28402 (N_28402,N_26373,N_26281);
and U28403 (N_28403,N_27432,N_25544);
or U28404 (N_28404,N_25492,N_26793);
nor U28405 (N_28405,N_26788,N_25985);
and U28406 (N_28406,N_25128,N_27306);
or U28407 (N_28407,N_27332,N_26255);
or U28408 (N_28408,N_25963,N_26800);
nand U28409 (N_28409,N_25068,N_25199);
nor U28410 (N_28410,N_26927,N_25045);
nand U28411 (N_28411,N_26551,N_25787);
nand U28412 (N_28412,N_26784,N_26753);
nand U28413 (N_28413,N_25247,N_27480);
nor U28414 (N_28414,N_26760,N_27087);
nand U28415 (N_28415,N_25441,N_25032);
and U28416 (N_28416,N_25597,N_25749);
or U28417 (N_28417,N_27355,N_27009);
or U28418 (N_28418,N_25758,N_26021);
and U28419 (N_28419,N_25982,N_25434);
nor U28420 (N_28420,N_26200,N_26783);
nor U28421 (N_28421,N_25695,N_25402);
or U28422 (N_28422,N_25688,N_25777);
or U28423 (N_28423,N_25082,N_27385);
and U28424 (N_28424,N_25470,N_25617);
nor U28425 (N_28425,N_25435,N_25454);
and U28426 (N_28426,N_25671,N_26577);
and U28427 (N_28427,N_26726,N_25573);
nand U28428 (N_28428,N_25801,N_26400);
nor U28429 (N_28429,N_25185,N_26144);
and U28430 (N_28430,N_25995,N_25853);
nand U28431 (N_28431,N_26422,N_27278);
nor U28432 (N_28432,N_26856,N_27284);
or U28433 (N_28433,N_25393,N_25075);
and U28434 (N_28434,N_26643,N_25216);
or U28435 (N_28435,N_26142,N_26816);
or U28436 (N_28436,N_27128,N_26682);
or U28437 (N_28437,N_27351,N_26430);
nor U28438 (N_28438,N_26716,N_25721);
nor U28439 (N_28439,N_25319,N_27270);
and U28440 (N_28440,N_26850,N_26370);
nor U28441 (N_28441,N_27460,N_26031);
or U28442 (N_28442,N_26820,N_26332);
and U28443 (N_28443,N_26770,N_25865);
nand U28444 (N_28444,N_25738,N_27150);
nor U28445 (N_28445,N_25025,N_26222);
nand U28446 (N_28446,N_26594,N_25043);
and U28447 (N_28447,N_27145,N_25647);
nor U28448 (N_28448,N_27447,N_27122);
or U28449 (N_28449,N_27183,N_25756);
and U28450 (N_28450,N_25204,N_26214);
or U28451 (N_28451,N_26727,N_25194);
or U28452 (N_28452,N_26588,N_26290);
xor U28453 (N_28453,N_26764,N_26704);
nand U28454 (N_28454,N_26703,N_26368);
and U28455 (N_28455,N_25895,N_26161);
or U28456 (N_28456,N_26963,N_25971);
xor U28457 (N_28457,N_25488,N_26589);
xor U28458 (N_28458,N_26050,N_27181);
and U28459 (N_28459,N_26978,N_25658);
and U28460 (N_28460,N_25902,N_26970);
xnor U28461 (N_28461,N_25884,N_26893);
and U28462 (N_28462,N_26082,N_26035);
or U28463 (N_28463,N_27360,N_25936);
or U28464 (N_28464,N_27340,N_26088);
and U28465 (N_28465,N_26759,N_26417);
and U28466 (N_28466,N_26017,N_25497);
or U28467 (N_28467,N_25945,N_25861);
and U28468 (N_28468,N_26431,N_26205);
or U28469 (N_28469,N_26099,N_27474);
or U28470 (N_28470,N_25304,N_26809);
nand U28471 (N_28471,N_25779,N_25500);
nor U28472 (N_28472,N_25948,N_27225);
nor U28473 (N_28473,N_25116,N_26877);
nand U28474 (N_28474,N_26562,N_27226);
and U28475 (N_28475,N_26377,N_25883);
nand U28476 (N_28476,N_26380,N_25370);
nand U28477 (N_28477,N_26258,N_26385);
nand U28478 (N_28478,N_26596,N_26897);
nand U28479 (N_28479,N_25299,N_25287);
xnor U28480 (N_28480,N_25822,N_26392);
nor U28481 (N_28481,N_26940,N_25904);
or U28482 (N_28482,N_26785,N_26864);
or U28483 (N_28483,N_25595,N_25114);
and U28484 (N_28484,N_25123,N_25344);
nand U28485 (N_28485,N_26958,N_26587);
or U28486 (N_28486,N_25893,N_27091);
and U28487 (N_28487,N_25823,N_26288);
and U28488 (N_28488,N_26631,N_25530);
nor U28489 (N_28489,N_27110,N_25255);
xor U28490 (N_28490,N_25443,N_26324);
nand U28491 (N_28491,N_26985,N_26062);
nand U28492 (N_28492,N_25177,N_27169);
nand U28493 (N_28493,N_26895,N_25917);
or U28494 (N_28494,N_26363,N_27175);
xor U28495 (N_28495,N_26165,N_26358);
nor U28496 (N_28496,N_25858,N_25781);
nor U28497 (N_28497,N_26409,N_25063);
or U28498 (N_28498,N_26151,N_26576);
nor U28499 (N_28499,N_25405,N_25817);
nor U28500 (N_28500,N_27313,N_26171);
nor U28501 (N_28501,N_27426,N_26560);
or U28502 (N_28502,N_26961,N_27247);
and U28503 (N_28503,N_25519,N_26208);
and U28504 (N_28504,N_26652,N_25446);
xnor U28505 (N_28505,N_26901,N_25428);
nand U28506 (N_28506,N_26625,N_26896);
nor U28507 (N_28507,N_25532,N_27453);
nand U28508 (N_28508,N_25268,N_26124);
and U28509 (N_28509,N_27307,N_26578);
nor U28510 (N_28510,N_26651,N_27114);
nor U28511 (N_28511,N_26907,N_25330);
or U28512 (N_28512,N_26734,N_26852);
and U28513 (N_28513,N_27193,N_25395);
nor U28514 (N_28514,N_26113,N_26532);
nor U28515 (N_28515,N_27098,N_27231);
nand U28516 (N_28516,N_26885,N_25810);
and U28517 (N_28517,N_25334,N_26387);
and U28518 (N_28518,N_26942,N_25501);
or U28519 (N_28519,N_25413,N_25445);
nor U28520 (N_28520,N_25097,N_25310);
nor U28521 (N_28521,N_26374,N_25242);
or U28522 (N_28522,N_26839,N_26872);
nor U28523 (N_28523,N_27255,N_26932);
and U28524 (N_28524,N_25623,N_25013);
and U28525 (N_28525,N_25062,N_26868);
nor U28526 (N_28526,N_27293,N_26572);
and U28527 (N_28527,N_25921,N_26184);
and U28528 (N_28528,N_26182,N_26873);
and U28529 (N_28529,N_27406,N_26935);
nor U28530 (N_28530,N_27001,N_26246);
and U28531 (N_28531,N_27415,N_26700);
or U28532 (N_28532,N_26972,N_26135);
nor U28533 (N_28533,N_25436,N_26480);
xor U28534 (N_28534,N_26664,N_26615);
nand U28535 (N_28535,N_26456,N_25741);
and U28536 (N_28536,N_25467,N_25710);
nor U28537 (N_28537,N_26273,N_25554);
or U28538 (N_28538,N_26685,N_26032);
nand U28539 (N_28539,N_26960,N_26264);
or U28540 (N_28540,N_26687,N_25629);
nor U28541 (N_28541,N_27024,N_26303);
or U28542 (N_28542,N_25033,N_26948);
nor U28543 (N_28543,N_26871,N_27419);
nor U28544 (N_28544,N_26322,N_26582);
and U28545 (N_28545,N_27041,N_26220);
or U28546 (N_28546,N_27199,N_25406);
nor U28547 (N_28547,N_26660,N_25708);
or U28548 (N_28548,N_25502,N_26274);
and U28549 (N_28549,N_25864,N_26891);
nand U28550 (N_28550,N_26145,N_26810);
nand U28551 (N_28551,N_27142,N_25389);
nor U28552 (N_28552,N_26115,N_26758);
and U28553 (N_28553,N_25535,N_25775);
xnor U28554 (N_28554,N_25326,N_25964);
or U28555 (N_28555,N_26688,N_27431);
xor U28556 (N_28556,N_25427,N_25048);
nor U28557 (N_28557,N_25143,N_25927);
and U28558 (N_28558,N_25080,N_26381);
nor U28559 (N_28559,N_26428,N_27053);
or U28560 (N_28560,N_25136,N_27341);
nand U28561 (N_28561,N_25566,N_26550);
and U28562 (N_28562,N_27449,N_25339);
and U28563 (N_28563,N_25318,N_26585);
xnor U28564 (N_28564,N_25253,N_25408);
nor U28565 (N_28565,N_26433,N_26632);
or U28566 (N_28566,N_27062,N_26081);
nand U28567 (N_28567,N_26858,N_26304);
nand U28568 (N_28568,N_27000,N_25826);
nor U28569 (N_28569,N_27280,N_25966);
and U28570 (N_28570,N_25463,N_26253);
nor U28571 (N_28571,N_26599,N_25536);
or U28572 (N_28572,N_26131,N_25190);
nand U28573 (N_28573,N_27034,N_26908);
xnor U28574 (N_28574,N_26922,N_25417);
nand U28575 (N_28575,N_27422,N_27151);
nor U28576 (N_28576,N_25754,N_25387);
nand U28577 (N_28577,N_27103,N_26346);
nand U28578 (N_28578,N_26565,N_25994);
and U28579 (N_28579,N_26105,N_25943);
and U28580 (N_28580,N_25679,N_25008);
xnor U28581 (N_28581,N_26657,N_27191);
nand U28582 (N_28582,N_25453,N_26217);
nor U28583 (N_28583,N_26091,N_26051);
nand U28584 (N_28584,N_26310,N_25477);
xnor U28585 (N_28585,N_25432,N_26710);
or U28586 (N_28586,N_27059,N_25954);
and U28587 (N_28587,N_26798,N_25626);
or U28588 (N_28588,N_26737,N_27037);
nand U28589 (N_28589,N_26924,N_25283);
xor U28590 (N_28590,N_27166,N_25124);
nand U28591 (N_28591,N_26575,N_27084);
and U28592 (N_28592,N_25526,N_25548);
nand U28593 (N_28593,N_25270,N_25482);
nand U28594 (N_28594,N_25457,N_27370);
and U28595 (N_28595,N_25506,N_27067);
nand U28596 (N_28596,N_25384,N_27296);
nand U28597 (N_28597,N_27349,N_26026);
or U28598 (N_28598,N_26157,N_25148);
xor U28599 (N_28599,N_25107,N_26843);
nand U28600 (N_28600,N_26684,N_26719);
and U28601 (N_28601,N_27436,N_26950);
and U28602 (N_28602,N_25704,N_25103);
nor U28603 (N_28603,N_26979,N_25672);
or U28604 (N_28604,N_26946,N_25892);
and U28605 (N_28605,N_26228,N_26561);
and U28606 (N_28606,N_25998,N_25275);
and U28607 (N_28607,N_25667,N_26749);
and U28608 (N_28608,N_27217,N_26814);
or U28609 (N_28609,N_26395,N_27063);
and U28610 (N_28610,N_25336,N_27092);
or U28611 (N_28611,N_25857,N_25663);
or U28612 (N_28612,N_25404,N_27274);
and U28613 (N_28613,N_25737,N_25620);
and U28614 (N_28614,N_26094,N_25475);
or U28615 (N_28615,N_25607,N_27131);
and U28616 (N_28616,N_26351,N_27006);
nor U28617 (N_28617,N_26355,N_26176);
or U28618 (N_28618,N_25576,N_25812);
nor U28619 (N_28619,N_26736,N_26146);
nand U28620 (N_28620,N_25480,N_25267);
nand U28621 (N_28621,N_26153,N_26636);
nor U28622 (N_28622,N_25471,N_25734);
xor U28623 (N_28623,N_26040,N_25323);
nor U28624 (N_28624,N_27047,N_25072);
xor U28625 (N_28625,N_26315,N_26133);
or U28626 (N_28626,N_25652,N_25377);
nor U28627 (N_28627,N_26067,N_25581);
nor U28628 (N_28628,N_26014,N_27189);
and U28629 (N_28629,N_26158,N_25562);
xnor U28630 (N_28630,N_26299,N_25876);
and U28631 (N_28631,N_26613,N_27036);
nand U28632 (N_28632,N_25545,N_25005);
nor U28633 (N_28633,N_26418,N_26842);
or U28634 (N_28634,N_27213,N_26552);
and U28635 (N_28635,N_26603,N_25301);
and U28636 (N_28636,N_25862,N_25602);
and U28637 (N_28637,N_26586,N_26574);
nor U28638 (N_28638,N_27470,N_26512);
nor U28639 (N_28639,N_26249,N_25491);
and U28640 (N_28640,N_26187,N_27168);
and U28641 (N_28641,N_25431,N_27286);
or U28642 (N_28642,N_26567,N_25364);
and U28643 (N_28643,N_25686,N_25838);
nand U28644 (N_28644,N_25317,N_27134);
and U28645 (N_28645,N_25931,N_26955);
or U28646 (N_28646,N_25076,N_27182);
nand U28647 (N_28647,N_27344,N_25638);
xnor U28648 (N_28648,N_26426,N_26445);
nor U28649 (N_28649,N_27389,N_25437);
and U28650 (N_28650,N_25584,N_25981);
and U28651 (N_28651,N_26966,N_26464);
nor U28652 (N_28652,N_25465,N_25852);
nor U28653 (N_28653,N_26194,N_25073);
xnor U28654 (N_28654,N_25683,N_27343);
or U28655 (N_28655,N_27051,N_27462);
nor U28656 (N_28656,N_26270,N_26423);
xor U28657 (N_28657,N_25232,N_26775);
nand U28658 (N_28658,N_26269,N_25572);
nor U28659 (N_28659,N_27031,N_25348);
and U28660 (N_28660,N_27102,N_26276);
and U28661 (N_28661,N_26309,N_26109);
or U28662 (N_28662,N_27372,N_25248);
or U28663 (N_28663,N_26093,N_27482);
and U28664 (N_28664,N_26390,N_25031);
xnor U28665 (N_28665,N_26231,N_26733);
nand U28666 (N_28666,N_25309,N_27345);
nor U28667 (N_28667,N_26510,N_26500);
or U28668 (N_28668,N_26256,N_25890);
nand U28669 (N_28669,N_27451,N_25350);
nor U28670 (N_28670,N_26548,N_27158);
and U28671 (N_28671,N_27410,N_27487);
and U28672 (N_28672,N_27237,N_26887);
and U28673 (N_28673,N_25628,N_25821);
or U28674 (N_28674,N_26973,N_27089);
or U28675 (N_28675,N_25776,N_25102);
nor U28676 (N_28676,N_27251,N_27465);
nor U28677 (N_28677,N_25885,N_26938);
nor U28678 (N_28678,N_26618,N_26353);
and U28679 (N_28679,N_25778,N_26886);
nand U28680 (N_28680,N_25784,N_25712);
and U28681 (N_28681,N_27146,N_25824);
nand U28682 (N_28682,N_25231,N_25797);
or U28683 (N_28683,N_25468,N_25972);
nor U28684 (N_28684,N_26497,N_25246);
nand U28685 (N_28685,N_27486,N_26669);
or U28686 (N_28686,N_25271,N_26455);
and U28687 (N_28687,N_26602,N_26621);
xnor U28688 (N_28688,N_27267,N_25380);
nand U28689 (N_28689,N_26527,N_25531);
and U28690 (N_28690,N_25011,N_26697);
nor U28691 (N_28691,N_26547,N_27204);
or U28692 (N_28692,N_25510,N_26936);
and U28693 (N_28693,N_25159,N_25466);
xnor U28694 (N_28694,N_27328,N_26639);
nand U28695 (N_28695,N_25765,N_27243);
and U28696 (N_28696,N_26033,N_27429);
nor U28697 (N_28697,N_27232,N_26097);
nand U28698 (N_28698,N_26913,N_26988);
xnor U28699 (N_28699,N_25371,N_26301);
xnor U28700 (N_28700,N_27242,N_25489);
nand U28701 (N_28701,N_25197,N_25230);
xor U28702 (N_28702,N_26634,N_26484);
or U28703 (N_28703,N_25254,N_26529);
xor U28704 (N_28704,N_26525,N_27216);
nor U28705 (N_28705,N_25564,N_26485);
nand U28706 (N_28706,N_27044,N_26516);
nor U28707 (N_28707,N_25036,N_25313);
xor U28708 (N_28708,N_25922,N_27192);
nor U28709 (N_28709,N_25423,N_27350);
or U28710 (N_28710,N_26427,N_27485);
nand U28711 (N_28711,N_27318,N_27105);
nor U28712 (N_28712,N_25198,N_26848);
and U28713 (N_28713,N_26203,N_27275);
nand U28714 (N_28714,N_26765,N_26899);
nand U28715 (N_28715,N_26211,N_27028);
nand U28716 (N_28716,N_25174,N_26168);
nor U28717 (N_28717,N_26677,N_25751);
nand U28718 (N_28718,N_26420,N_25448);
nor U28719 (N_28719,N_25832,N_25898);
and U28720 (N_28720,N_25388,N_25218);
nor U28721 (N_28721,N_27081,N_27180);
nor U28722 (N_28722,N_25205,N_27257);
and U28723 (N_28723,N_26740,N_27109);
and U28724 (N_28724,N_25860,N_25523);
nor U28725 (N_28725,N_26402,N_25891);
nor U28726 (N_28726,N_25414,N_27321);
xnor U28727 (N_28727,N_27228,N_27052);
nand U28728 (N_28728,N_26401,N_26654);
or U28729 (N_28729,N_25172,N_25731);
nand U28730 (N_28730,N_25967,N_27366);
and U28731 (N_28731,N_26771,N_25621);
or U28732 (N_28732,N_25997,N_26945);
or U28733 (N_28733,N_26038,N_26518);
or U28734 (N_28734,N_25856,N_27400);
nor U28735 (N_28735,N_26065,N_25264);
and U28736 (N_28736,N_25699,N_25992);
nor U28737 (N_28737,N_25719,N_26000);
nor U28738 (N_28738,N_25379,N_26752);
or U28739 (N_28739,N_25577,N_25729);
and U28740 (N_28740,N_26975,N_27283);
nor U28741 (N_28741,N_25887,N_27279);
nand U28742 (N_28742,N_25215,N_25946);
or U28743 (N_28743,N_26424,N_25714);
nand U28744 (N_28744,N_25869,N_26112);
nor U28745 (N_28745,N_26318,N_27206);
nor U28746 (N_28746,N_27294,N_27304);
xor U28747 (N_28747,N_25583,N_27219);
and U28748 (N_28748,N_27261,N_27469);
or U28749 (N_28749,N_26976,N_26119);
nand U28750 (N_28750,N_26236,N_25344);
nor U28751 (N_28751,N_25105,N_26435);
nand U28752 (N_28752,N_26826,N_26073);
and U28753 (N_28753,N_26127,N_26882);
xnor U28754 (N_28754,N_27087,N_27142);
xor U28755 (N_28755,N_25721,N_26731);
nor U28756 (N_28756,N_26729,N_27066);
nand U28757 (N_28757,N_26865,N_25722);
and U28758 (N_28758,N_25859,N_25507);
and U28759 (N_28759,N_27145,N_25092);
xor U28760 (N_28760,N_26612,N_27476);
nor U28761 (N_28761,N_25948,N_26422);
xor U28762 (N_28762,N_27484,N_27400);
nor U28763 (N_28763,N_27028,N_25788);
nand U28764 (N_28764,N_27058,N_25279);
xor U28765 (N_28765,N_27308,N_26283);
nor U28766 (N_28766,N_25157,N_27239);
nor U28767 (N_28767,N_26314,N_27383);
or U28768 (N_28768,N_26707,N_26482);
nor U28769 (N_28769,N_25622,N_25101);
nand U28770 (N_28770,N_27378,N_26595);
or U28771 (N_28771,N_26802,N_25216);
or U28772 (N_28772,N_26528,N_26314);
or U28773 (N_28773,N_27171,N_26087);
and U28774 (N_28774,N_26337,N_27334);
or U28775 (N_28775,N_26338,N_26540);
nor U28776 (N_28776,N_25525,N_25502);
xnor U28777 (N_28777,N_27344,N_27398);
nand U28778 (N_28778,N_27191,N_26422);
nor U28779 (N_28779,N_27472,N_25929);
and U28780 (N_28780,N_25002,N_25515);
and U28781 (N_28781,N_26832,N_26127);
nand U28782 (N_28782,N_25197,N_26436);
or U28783 (N_28783,N_25052,N_25868);
or U28784 (N_28784,N_26506,N_26659);
xnor U28785 (N_28785,N_25948,N_25270);
or U28786 (N_28786,N_27339,N_27493);
and U28787 (N_28787,N_25244,N_26449);
nor U28788 (N_28788,N_26994,N_25895);
and U28789 (N_28789,N_25464,N_25888);
nor U28790 (N_28790,N_25051,N_25232);
nand U28791 (N_28791,N_25488,N_25440);
nand U28792 (N_28792,N_26873,N_27414);
or U28793 (N_28793,N_25698,N_25361);
nand U28794 (N_28794,N_25906,N_26979);
xnor U28795 (N_28795,N_25253,N_25141);
nand U28796 (N_28796,N_26940,N_26545);
or U28797 (N_28797,N_27030,N_25778);
and U28798 (N_28798,N_25915,N_25062);
and U28799 (N_28799,N_26250,N_27003);
or U28800 (N_28800,N_27157,N_27021);
and U28801 (N_28801,N_27421,N_25084);
nand U28802 (N_28802,N_27068,N_26665);
or U28803 (N_28803,N_26654,N_27366);
nor U28804 (N_28804,N_27325,N_25751);
nand U28805 (N_28805,N_26444,N_26768);
nand U28806 (N_28806,N_25952,N_27220);
xnor U28807 (N_28807,N_27088,N_27205);
nand U28808 (N_28808,N_27338,N_27230);
or U28809 (N_28809,N_27206,N_25727);
and U28810 (N_28810,N_25690,N_27427);
nor U28811 (N_28811,N_25108,N_26562);
nor U28812 (N_28812,N_25105,N_25893);
xor U28813 (N_28813,N_26262,N_26410);
or U28814 (N_28814,N_26732,N_27136);
and U28815 (N_28815,N_25451,N_25179);
and U28816 (N_28816,N_27373,N_27274);
nand U28817 (N_28817,N_25862,N_27199);
nand U28818 (N_28818,N_25606,N_27154);
and U28819 (N_28819,N_25639,N_25047);
and U28820 (N_28820,N_27017,N_25562);
xnor U28821 (N_28821,N_27439,N_26799);
nor U28822 (N_28822,N_25729,N_25538);
or U28823 (N_28823,N_26282,N_27102);
or U28824 (N_28824,N_27388,N_25617);
or U28825 (N_28825,N_26441,N_26910);
nor U28826 (N_28826,N_27406,N_27047);
or U28827 (N_28827,N_27366,N_26200);
nand U28828 (N_28828,N_26468,N_25025);
or U28829 (N_28829,N_25442,N_25162);
or U28830 (N_28830,N_27303,N_25811);
and U28831 (N_28831,N_25590,N_27361);
nor U28832 (N_28832,N_26872,N_26895);
xor U28833 (N_28833,N_27217,N_25289);
and U28834 (N_28834,N_25247,N_25972);
nor U28835 (N_28835,N_25970,N_26974);
nor U28836 (N_28836,N_26541,N_26893);
and U28837 (N_28837,N_25985,N_25952);
xor U28838 (N_28838,N_27096,N_26120);
xor U28839 (N_28839,N_25743,N_26607);
or U28840 (N_28840,N_25645,N_25967);
or U28841 (N_28841,N_26390,N_27075);
or U28842 (N_28842,N_27149,N_25636);
or U28843 (N_28843,N_26559,N_27377);
and U28844 (N_28844,N_26191,N_26627);
or U28845 (N_28845,N_26315,N_26654);
and U28846 (N_28846,N_26860,N_26991);
nand U28847 (N_28847,N_25672,N_26025);
nand U28848 (N_28848,N_25032,N_25074);
nor U28849 (N_28849,N_26390,N_26457);
or U28850 (N_28850,N_25623,N_25610);
xnor U28851 (N_28851,N_26848,N_26290);
and U28852 (N_28852,N_26384,N_27114);
and U28853 (N_28853,N_26920,N_25592);
and U28854 (N_28854,N_25166,N_27009);
xnor U28855 (N_28855,N_26384,N_27038);
nand U28856 (N_28856,N_25256,N_26754);
and U28857 (N_28857,N_25641,N_27261);
nor U28858 (N_28858,N_27447,N_25398);
and U28859 (N_28859,N_25708,N_25672);
or U28860 (N_28860,N_26420,N_26391);
nor U28861 (N_28861,N_26106,N_26409);
nand U28862 (N_28862,N_25290,N_26051);
and U28863 (N_28863,N_26850,N_26506);
and U28864 (N_28864,N_25186,N_26196);
and U28865 (N_28865,N_25431,N_26431);
nor U28866 (N_28866,N_27353,N_26645);
nor U28867 (N_28867,N_26360,N_25201);
nand U28868 (N_28868,N_26049,N_26420);
nand U28869 (N_28869,N_26174,N_27021);
nor U28870 (N_28870,N_26277,N_26742);
nor U28871 (N_28871,N_25705,N_27230);
or U28872 (N_28872,N_25270,N_26784);
nor U28873 (N_28873,N_25273,N_26737);
nor U28874 (N_28874,N_27131,N_26313);
nor U28875 (N_28875,N_26254,N_26893);
nor U28876 (N_28876,N_25919,N_25871);
and U28877 (N_28877,N_25432,N_25387);
or U28878 (N_28878,N_26621,N_25160);
and U28879 (N_28879,N_25919,N_26381);
nand U28880 (N_28880,N_26832,N_26521);
nand U28881 (N_28881,N_25994,N_25703);
and U28882 (N_28882,N_26015,N_25706);
nor U28883 (N_28883,N_26107,N_25608);
nor U28884 (N_28884,N_25857,N_25390);
nor U28885 (N_28885,N_27318,N_26492);
nor U28886 (N_28886,N_25634,N_26951);
and U28887 (N_28887,N_27481,N_25173);
nand U28888 (N_28888,N_25792,N_27202);
nand U28889 (N_28889,N_27429,N_26357);
nand U28890 (N_28890,N_26175,N_25406);
and U28891 (N_28891,N_25978,N_25738);
xnor U28892 (N_28892,N_26979,N_27299);
nand U28893 (N_28893,N_26658,N_26569);
and U28894 (N_28894,N_27466,N_26388);
or U28895 (N_28895,N_26260,N_26130);
and U28896 (N_28896,N_26356,N_27082);
or U28897 (N_28897,N_26491,N_27086);
nor U28898 (N_28898,N_26149,N_26814);
nor U28899 (N_28899,N_25471,N_26628);
and U28900 (N_28900,N_26111,N_26008);
nand U28901 (N_28901,N_26001,N_26460);
and U28902 (N_28902,N_26668,N_25783);
or U28903 (N_28903,N_25065,N_27031);
and U28904 (N_28904,N_26446,N_27434);
and U28905 (N_28905,N_27000,N_27239);
or U28906 (N_28906,N_25981,N_25276);
nand U28907 (N_28907,N_26871,N_25842);
and U28908 (N_28908,N_26559,N_26856);
nand U28909 (N_28909,N_27104,N_26823);
nor U28910 (N_28910,N_26449,N_26188);
or U28911 (N_28911,N_27455,N_27289);
xnor U28912 (N_28912,N_26950,N_27484);
nand U28913 (N_28913,N_25017,N_27198);
and U28914 (N_28914,N_26959,N_25615);
nand U28915 (N_28915,N_27413,N_26938);
and U28916 (N_28916,N_27040,N_25631);
and U28917 (N_28917,N_25827,N_26754);
and U28918 (N_28918,N_25036,N_25564);
nand U28919 (N_28919,N_25314,N_25110);
nand U28920 (N_28920,N_27101,N_26169);
and U28921 (N_28921,N_25221,N_26932);
nor U28922 (N_28922,N_26835,N_25721);
nor U28923 (N_28923,N_25471,N_25434);
nor U28924 (N_28924,N_25689,N_25124);
nor U28925 (N_28925,N_26659,N_25831);
and U28926 (N_28926,N_26202,N_26383);
and U28927 (N_28927,N_25997,N_25291);
or U28928 (N_28928,N_26511,N_26072);
nand U28929 (N_28929,N_26549,N_27295);
or U28930 (N_28930,N_26017,N_26782);
or U28931 (N_28931,N_27187,N_25078);
nand U28932 (N_28932,N_26635,N_26288);
nand U28933 (N_28933,N_25163,N_25760);
nand U28934 (N_28934,N_27409,N_26170);
or U28935 (N_28935,N_27207,N_25686);
nor U28936 (N_28936,N_27032,N_26833);
or U28937 (N_28937,N_26171,N_27377);
or U28938 (N_28938,N_26847,N_25975);
nand U28939 (N_28939,N_25609,N_27007);
nand U28940 (N_28940,N_26582,N_26757);
and U28941 (N_28941,N_25427,N_25667);
or U28942 (N_28942,N_27338,N_27213);
xnor U28943 (N_28943,N_26868,N_26778);
and U28944 (N_28944,N_26917,N_25829);
or U28945 (N_28945,N_27009,N_27498);
xor U28946 (N_28946,N_26470,N_25470);
and U28947 (N_28947,N_27038,N_25788);
nand U28948 (N_28948,N_26852,N_27407);
nor U28949 (N_28949,N_25349,N_27212);
nand U28950 (N_28950,N_26954,N_25994);
or U28951 (N_28951,N_27087,N_27369);
or U28952 (N_28952,N_26033,N_26902);
nand U28953 (N_28953,N_27483,N_25932);
and U28954 (N_28954,N_26047,N_26375);
or U28955 (N_28955,N_26630,N_26190);
or U28956 (N_28956,N_25713,N_27496);
and U28957 (N_28957,N_26502,N_27421);
nor U28958 (N_28958,N_27249,N_27135);
xnor U28959 (N_28959,N_25963,N_25324);
xnor U28960 (N_28960,N_27408,N_27266);
nand U28961 (N_28961,N_25074,N_26689);
or U28962 (N_28962,N_25845,N_26295);
nor U28963 (N_28963,N_25190,N_26602);
nand U28964 (N_28964,N_27174,N_26959);
or U28965 (N_28965,N_26373,N_27244);
or U28966 (N_28966,N_27141,N_25110);
or U28967 (N_28967,N_25983,N_27200);
and U28968 (N_28968,N_25443,N_26049);
nand U28969 (N_28969,N_26588,N_25667);
and U28970 (N_28970,N_26097,N_27171);
nor U28971 (N_28971,N_25585,N_27176);
nand U28972 (N_28972,N_26872,N_26533);
nand U28973 (N_28973,N_25996,N_26149);
nand U28974 (N_28974,N_26998,N_26699);
and U28975 (N_28975,N_25888,N_25674);
xor U28976 (N_28976,N_25310,N_25093);
nand U28977 (N_28977,N_26417,N_26328);
nand U28978 (N_28978,N_27207,N_26935);
nor U28979 (N_28979,N_26385,N_25483);
xnor U28980 (N_28980,N_27171,N_26232);
nand U28981 (N_28981,N_26310,N_27429);
nand U28982 (N_28982,N_26040,N_25335);
nor U28983 (N_28983,N_27252,N_27236);
or U28984 (N_28984,N_25217,N_27164);
nand U28985 (N_28985,N_27166,N_25538);
nand U28986 (N_28986,N_26260,N_25159);
and U28987 (N_28987,N_26036,N_25437);
and U28988 (N_28988,N_25572,N_25426);
nor U28989 (N_28989,N_26225,N_26955);
nand U28990 (N_28990,N_25859,N_25355);
xor U28991 (N_28991,N_26903,N_25753);
nor U28992 (N_28992,N_26403,N_26350);
nand U28993 (N_28993,N_27201,N_27251);
and U28994 (N_28994,N_26462,N_25153);
and U28995 (N_28995,N_25933,N_27030);
xnor U28996 (N_28996,N_27123,N_26655);
or U28997 (N_28997,N_25228,N_25538);
nor U28998 (N_28998,N_25664,N_27337);
or U28999 (N_28999,N_25696,N_26105);
nand U29000 (N_29000,N_26289,N_26267);
or U29001 (N_29001,N_27245,N_25380);
nand U29002 (N_29002,N_25340,N_25717);
xor U29003 (N_29003,N_25022,N_25363);
or U29004 (N_29004,N_25542,N_26180);
nand U29005 (N_29005,N_26510,N_25833);
or U29006 (N_29006,N_26604,N_25567);
or U29007 (N_29007,N_27287,N_25014);
and U29008 (N_29008,N_26648,N_25523);
nor U29009 (N_29009,N_27134,N_26014);
nor U29010 (N_29010,N_26692,N_25716);
xnor U29011 (N_29011,N_25085,N_26822);
or U29012 (N_29012,N_27456,N_25302);
nor U29013 (N_29013,N_26194,N_25921);
nor U29014 (N_29014,N_25852,N_27193);
or U29015 (N_29015,N_25073,N_25601);
nor U29016 (N_29016,N_26665,N_25749);
or U29017 (N_29017,N_25416,N_27005);
nor U29018 (N_29018,N_27484,N_26521);
nand U29019 (N_29019,N_27295,N_25538);
and U29020 (N_29020,N_25513,N_25848);
xor U29021 (N_29021,N_26140,N_27125);
nand U29022 (N_29022,N_27125,N_26887);
nand U29023 (N_29023,N_26618,N_26953);
and U29024 (N_29024,N_25000,N_25485);
or U29025 (N_29025,N_25081,N_27391);
nand U29026 (N_29026,N_27495,N_26650);
and U29027 (N_29027,N_26989,N_25784);
nand U29028 (N_29028,N_25294,N_26124);
and U29029 (N_29029,N_26762,N_26040);
and U29030 (N_29030,N_25490,N_27400);
or U29031 (N_29031,N_26209,N_26769);
nand U29032 (N_29032,N_26587,N_27431);
or U29033 (N_29033,N_27340,N_26163);
nor U29034 (N_29034,N_25160,N_26165);
and U29035 (N_29035,N_26454,N_25052);
nand U29036 (N_29036,N_26106,N_26791);
and U29037 (N_29037,N_27027,N_25931);
nor U29038 (N_29038,N_25806,N_26164);
and U29039 (N_29039,N_26718,N_26058);
nor U29040 (N_29040,N_26338,N_27493);
nor U29041 (N_29041,N_26588,N_26027);
nand U29042 (N_29042,N_26874,N_27456);
nor U29043 (N_29043,N_25004,N_26816);
and U29044 (N_29044,N_26858,N_25614);
nor U29045 (N_29045,N_25301,N_27438);
xnor U29046 (N_29046,N_26065,N_25474);
and U29047 (N_29047,N_25324,N_26638);
nor U29048 (N_29048,N_25524,N_25461);
nor U29049 (N_29049,N_26884,N_25712);
or U29050 (N_29050,N_26084,N_25256);
xnor U29051 (N_29051,N_26297,N_27138);
or U29052 (N_29052,N_27404,N_25686);
and U29053 (N_29053,N_26636,N_26576);
nand U29054 (N_29054,N_27107,N_26668);
nand U29055 (N_29055,N_26571,N_27288);
nor U29056 (N_29056,N_25109,N_26772);
or U29057 (N_29057,N_27106,N_26736);
nand U29058 (N_29058,N_26775,N_26026);
nand U29059 (N_29059,N_26621,N_27420);
nor U29060 (N_29060,N_25248,N_25776);
and U29061 (N_29061,N_26101,N_27197);
or U29062 (N_29062,N_25814,N_25807);
nand U29063 (N_29063,N_27026,N_27410);
nor U29064 (N_29064,N_26450,N_27425);
nor U29065 (N_29065,N_26947,N_25916);
nor U29066 (N_29066,N_26121,N_25479);
and U29067 (N_29067,N_25757,N_26090);
nand U29068 (N_29068,N_25311,N_25754);
and U29069 (N_29069,N_26432,N_27025);
nand U29070 (N_29070,N_25351,N_26222);
or U29071 (N_29071,N_26317,N_25950);
nand U29072 (N_29072,N_26862,N_26175);
and U29073 (N_29073,N_27308,N_25377);
or U29074 (N_29074,N_26982,N_25659);
or U29075 (N_29075,N_26331,N_25432);
or U29076 (N_29076,N_26889,N_26183);
and U29077 (N_29077,N_26438,N_26183);
xnor U29078 (N_29078,N_25917,N_26136);
and U29079 (N_29079,N_25376,N_27372);
xor U29080 (N_29080,N_25728,N_27229);
nand U29081 (N_29081,N_26617,N_26624);
or U29082 (N_29082,N_25376,N_27483);
nand U29083 (N_29083,N_25613,N_27484);
and U29084 (N_29084,N_25196,N_25384);
nor U29085 (N_29085,N_26027,N_26315);
nor U29086 (N_29086,N_27465,N_26201);
and U29087 (N_29087,N_26494,N_25818);
and U29088 (N_29088,N_26311,N_26456);
and U29089 (N_29089,N_25738,N_26372);
and U29090 (N_29090,N_27042,N_25073);
nand U29091 (N_29091,N_27266,N_25081);
and U29092 (N_29092,N_27046,N_26564);
xnor U29093 (N_29093,N_26266,N_26613);
and U29094 (N_29094,N_26230,N_27367);
nand U29095 (N_29095,N_25206,N_27083);
or U29096 (N_29096,N_27015,N_27251);
nor U29097 (N_29097,N_26931,N_27445);
nand U29098 (N_29098,N_25154,N_26244);
nand U29099 (N_29099,N_25142,N_26400);
and U29100 (N_29100,N_26164,N_26069);
nand U29101 (N_29101,N_25968,N_26310);
or U29102 (N_29102,N_26709,N_25937);
nand U29103 (N_29103,N_25470,N_26646);
or U29104 (N_29104,N_25363,N_27491);
or U29105 (N_29105,N_25580,N_25224);
xnor U29106 (N_29106,N_25987,N_26713);
or U29107 (N_29107,N_26730,N_26063);
nand U29108 (N_29108,N_26894,N_26457);
xnor U29109 (N_29109,N_25852,N_25413);
nand U29110 (N_29110,N_27387,N_26538);
or U29111 (N_29111,N_26164,N_26915);
nand U29112 (N_29112,N_26744,N_26999);
nand U29113 (N_29113,N_26016,N_27368);
xnor U29114 (N_29114,N_26158,N_27059);
or U29115 (N_29115,N_26021,N_25917);
or U29116 (N_29116,N_26491,N_25123);
nor U29117 (N_29117,N_25109,N_26504);
nand U29118 (N_29118,N_27241,N_25016);
nor U29119 (N_29119,N_25322,N_27359);
or U29120 (N_29120,N_26696,N_27313);
nand U29121 (N_29121,N_26595,N_25474);
or U29122 (N_29122,N_25651,N_25204);
and U29123 (N_29123,N_27026,N_25227);
and U29124 (N_29124,N_26116,N_27014);
and U29125 (N_29125,N_25173,N_26244);
xor U29126 (N_29126,N_25126,N_27149);
or U29127 (N_29127,N_25406,N_25189);
and U29128 (N_29128,N_26145,N_27152);
and U29129 (N_29129,N_25618,N_25449);
or U29130 (N_29130,N_25332,N_25570);
or U29131 (N_29131,N_27290,N_25648);
nand U29132 (N_29132,N_27272,N_25486);
xnor U29133 (N_29133,N_27021,N_25730);
xnor U29134 (N_29134,N_25457,N_25749);
nand U29135 (N_29135,N_26514,N_26304);
and U29136 (N_29136,N_27372,N_27153);
or U29137 (N_29137,N_26920,N_27468);
xnor U29138 (N_29138,N_26326,N_25868);
xnor U29139 (N_29139,N_26407,N_26380);
xnor U29140 (N_29140,N_27071,N_25927);
and U29141 (N_29141,N_25664,N_26615);
or U29142 (N_29142,N_26045,N_26006);
nand U29143 (N_29143,N_25458,N_27131);
nand U29144 (N_29144,N_26007,N_26824);
nor U29145 (N_29145,N_25546,N_27286);
nor U29146 (N_29146,N_25958,N_25388);
xor U29147 (N_29147,N_26541,N_27199);
or U29148 (N_29148,N_26240,N_25449);
or U29149 (N_29149,N_26164,N_25035);
or U29150 (N_29150,N_26891,N_27137);
nor U29151 (N_29151,N_25946,N_25872);
and U29152 (N_29152,N_25053,N_25858);
and U29153 (N_29153,N_25333,N_26558);
nand U29154 (N_29154,N_25883,N_26246);
nor U29155 (N_29155,N_25741,N_25742);
or U29156 (N_29156,N_25085,N_26888);
nor U29157 (N_29157,N_27358,N_27402);
and U29158 (N_29158,N_25757,N_26129);
and U29159 (N_29159,N_25609,N_27020);
nand U29160 (N_29160,N_26830,N_26359);
or U29161 (N_29161,N_26020,N_26749);
nand U29162 (N_29162,N_26234,N_27183);
nand U29163 (N_29163,N_26699,N_25803);
or U29164 (N_29164,N_26541,N_26912);
and U29165 (N_29165,N_26543,N_26401);
or U29166 (N_29166,N_26366,N_27217);
nand U29167 (N_29167,N_25335,N_26763);
nor U29168 (N_29168,N_26849,N_26564);
and U29169 (N_29169,N_25931,N_25593);
nor U29170 (N_29170,N_26260,N_26587);
nand U29171 (N_29171,N_25904,N_25773);
nand U29172 (N_29172,N_26218,N_27279);
nor U29173 (N_29173,N_25991,N_27499);
nor U29174 (N_29174,N_26224,N_25453);
nor U29175 (N_29175,N_27109,N_26208);
and U29176 (N_29176,N_25883,N_25991);
nor U29177 (N_29177,N_26450,N_25362);
nand U29178 (N_29178,N_25522,N_25397);
nand U29179 (N_29179,N_26622,N_26991);
and U29180 (N_29180,N_26257,N_25800);
and U29181 (N_29181,N_26638,N_26097);
and U29182 (N_29182,N_27089,N_25518);
nor U29183 (N_29183,N_25873,N_27278);
or U29184 (N_29184,N_25717,N_27153);
nand U29185 (N_29185,N_25751,N_26472);
nand U29186 (N_29186,N_25689,N_26481);
nor U29187 (N_29187,N_26839,N_25276);
nor U29188 (N_29188,N_25703,N_26922);
or U29189 (N_29189,N_26043,N_25330);
nand U29190 (N_29190,N_27357,N_25951);
or U29191 (N_29191,N_26597,N_26238);
nand U29192 (N_29192,N_25420,N_25954);
or U29193 (N_29193,N_27474,N_27258);
nand U29194 (N_29194,N_25095,N_26711);
xor U29195 (N_29195,N_25867,N_27366);
nand U29196 (N_29196,N_26396,N_26276);
nor U29197 (N_29197,N_27081,N_26347);
xor U29198 (N_29198,N_26765,N_26047);
xor U29199 (N_29199,N_27180,N_27092);
xor U29200 (N_29200,N_25071,N_25906);
nor U29201 (N_29201,N_27138,N_26834);
nand U29202 (N_29202,N_25897,N_27273);
nand U29203 (N_29203,N_25896,N_25694);
nor U29204 (N_29204,N_26896,N_26772);
nand U29205 (N_29205,N_27343,N_26090);
nand U29206 (N_29206,N_27441,N_26641);
or U29207 (N_29207,N_25305,N_26587);
nor U29208 (N_29208,N_25624,N_26678);
nand U29209 (N_29209,N_26242,N_25092);
nand U29210 (N_29210,N_26324,N_26815);
and U29211 (N_29211,N_26782,N_26112);
nand U29212 (N_29212,N_26724,N_26615);
or U29213 (N_29213,N_25895,N_25405);
nand U29214 (N_29214,N_26530,N_26332);
xnor U29215 (N_29215,N_27064,N_26735);
and U29216 (N_29216,N_25138,N_25889);
or U29217 (N_29217,N_26636,N_25212);
and U29218 (N_29218,N_25243,N_25708);
and U29219 (N_29219,N_27476,N_26909);
and U29220 (N_29220,N_27343,N_26101);
nand U29221 (N_29221,N_25632,N_25897);
and U29222 (N_29222,N_26436,N_27158);
and U29223 (N_29223,N_25010,N_25075);
nor U29224 (N_29224,N_26947,N_26641);
and U29225 (N_29225,N_27408,N_26788);
nor U29226 (N_29226,N_25009,N_25242);
xor U29227 (N_29227,N_26860,N_26205);
nor U29228 (N_29228,N_26775,N_26975);
nand U29229 (N_29229,N_25472,N_25805);
nand U29230 (N_29230,N_27169,N_27423);
and U29231 (N_29231,N_26297,N_25180);
xnor U29232 (N_29232,N_25885,N_26912);
nand U29233 (N_29233,N_25834,N_26863);
or U29234 (N_29234,N_27232,N_25702);
or U29235 (N_29235,N_25303,N_27264);
or U29236 (N_29236,N_27407,N_27328);
and U29237 (N_29237,N_25497,N_25585);
nor U29238 (N_29238,N_25048,N_26240);
and U29239 (N_29239,N_27253,N_26712);
and U29240 (N_29240,N_26677,N_26006);
nor U29241 (N_29241,N_26883,N_25784);
or U29242 (N_29242,N_25564,N_25587);
or U29243 (N_29243,N_25496,N_25045);
or U29244 (N_29244,N_27293,N_26600);
nor U29245 (N_29245,N_26603,N_27055);
and U29246 (N_29246,N_26273,N_25062);
nor U29247 (N_29247,N_27279,N_25220);
nand U29248 (N_29248,N_26867,N_25692);
and U29249 (N_29249,N_26303,N_26563);
xnor U29250 (N_29250,N_27372,N_26463);
nor U29251 (N_29251,N_27089,N_26746);
xnor U29252 (N_29252,N_25704,N_25688);
nand U29253 (N_29253,N_25177,N_27295);
nand U29254 (N_29254,N_25916,N_27436);
xnor U29255 (N_29255,N_25078,N_26864);
xor U29256 (N_29256,N_27368,N_27438);
nand U29257 (N_29257,N_26476,N_27385);
nor U29258 (N_29258,N_26250,N_25004);
and U29259 (N_29259,N_25901,N_25465);
xnor U29260 (N_29260,N_26342,N_26458);
nor U29261 (N_29261,N_26268,N_27181);
nor U29262 (N_29262,N_25199,N_26384);
nor U29263 (N_29263,N_26523,N_26525);
and U29264 (N_29264,N_27379,N_25798);
or U29265 (N_29265,N_25794,N_26921);
nor U29266 (N_29266,N_25346,N_26102);
or U29267 (N_29267,N_26207,N_27148);
nor U29268 (N_29268,N_26175,N_25570);
or U29269 (N_29269,N_25709,N_27332);
nor U29270 (N_29270,N_25958,N_26145);
and U29271 (N_29271,N_26316,N_25096);
and U29272 (N_29272,N_26796,N_26560);
and U29273 (N_29273,N_26258,N_25531);
nor U29274 (N_29274,N_27024,N_25177);
nor U29275 (N_29275,N_26070,N_25354);
and U29276 (N_29276,N_27202,N_26372);
nand U29277 (N_29277,N_26707,N_25576);
nand U29278 (N_29278,N_25664,N_25397);
xor U29279 (N_29279,N_25865,N_26855);
nand U29280 (N_29280,N_25260,N_27280);
and U29281 (N_29281,N_26579,N_26032);
nor U29282 (N_29282,N_26162,N_27460);
nor U29283 (N_29283,N_27222,N_27347);
and U29284 (N_29284,N_26415,N_26234);
or U29285 (N_29285,N_25596,N_26701);
xnor U29286 (N_29286,N_26140,N_27077);
nor U29287 (N_29287,N_25156,N_26536);
and U29288 (N_29288,N_26999,N_25466);
nor U29289 (N_29289,N_27081,N_26643);
and U29290 (N_29290,N_25423,N_26857);
and U29291 (N_29291,N_26922,N_27091);
and U29292 (N_29292,N_25335,N_26710);
or U29293 (N_29293,N_26760,N_26276);
nand U29294 (N_29294,N_26686,N_26496);
nand U29295 (N_29295,N_26704,N_25997);
nand U29296 (N_29296,N_25890,N_27060);
and U29297 (N_29297,N_26858,N_27049);
nand U29298 (N_29298,N_26042,N_25414);
nor U29299 (N_29299,N_27229,N_26627);
and U29300 (N_29300,N_27230,N_27401);
and U29301 (N_29301,N_25552,N_25471);
or U29302 (N_29302,N_26047,N_27375);
or U29303 (N_29303,N_27359,N_26298);
nand U29304 (N_29304,N_25347,N_27302);
nand U29305 (N_29305,N_25046,N_25016);
nand U29306 (N_29306,N_25929,N_25091);
nor U29307 (N_29307,N_25115,N_25140);
and U29308 (N_29308,N_26867,N_26264);
nor U29309 (N_29309,N_27147,N_26049);
or U29310 (N_29310,N_25710,N_27319);
nor U29311 (N_29311,N_27177,N_27336);
nand U29312 (N_29312,N_27220,N_26802);
nand U29313 (N_29313,N_26080,N_26515);
or U29314 (N_29314,N_27370,N_26904);
nand U29315 (N_29315,N_26256,N_27193);
nand U29316 (N_29316,N_27306,N_26901);
xor U29317 (N_29317,N_26680,N_25788);
or U29318 (N_29318,N_26228,N_26601);
and U29319 (N_29319,N_26464,N_26158);
nor U29320 (N_29320,N_27297,N_27315);
and U29321 (N_29321,N_26124,N_27406);
or U29322 (N_29322,N_26055,N_25701);
and U29323 (N_29323,N_26374,N_25001);
and U29324 (N_29324,N_26134,N_26816);
and U29325 (N_29325,N_26475,N_26601);
or U29326 (N_29326,N_25726,N_25503);
and U29327 (N_29327,N_27303,N_25998);
nand U29328 (N_29328,N_27448,N_27333);
nand U29329 (N_29329,N_25044,N_26637);
nand U29330 (N_29330,N_25482,N_27487);
xnor U29331 (N_29331,N_25918,N_26975);
nand U29332 (N_29332,N_27014,N_26902);
or U29333 (N_29333,N_25763,N_27157);
or U29334 (N_29334,N_26786,N_26255);
and U29335 (N_29335,N_25670,N_26842);
xor U29336 (N_29336,N_27099,N_25502);
nand U29337 (N_29337,N_27177,N_25431);
nor U29338 (N_29338,N_25454,N_25159);
nor U29339 (N_29339,N_27015,N_25245);
nor U29340 (N_29340,N_27457,N_26175);
nand U29341 (N_29341,N_26536,N_27072);
or U29342 (N_29342,N_25639,N_25431);
or U29343 (N_29343,N_26991,N_25214);
xnor U29344 (N_29344,N_25385,N_27316);
nor U29345 (N_29345,N_25902,N_26397);
or U29346 (N_29346,N_26550,N_26587);
nand U29347 (N_29347,N_26712,N_25296);
nand U29348 (N_29348,N_25963,N_26451);
and U29349 (N_29349,N_26553,N_26363);
nand U29350 (N_29350,N_25468,N_27459);
xor U29351 (N_29351,N_27054,N_25174);
nor U29352 (N_29352,N_27215,N_25757);
nand U29353 (N_29353,N_27117,N_26027);
and U29354 (N_29354,N_26893,N_25051);
nor U29355 (N_29355,N_26661,N_25690);
and U29356 (N_29356,N_25775,N_27310);
nor U29357 (N_29357,N_25696,N_26533);
nand U29358 (N_29358,N_26632,N_26742);
or U29359 (N_29359,N_26929,N_26374);
nor U29360 (N_29360,N_25136,N_25431);
or U29361 (N_29361,N_25343,N_25586);
nor U29362 (N_29362,N_25142,N_26383);
nand U29363 (N_29363,N_26056,N_26789);
nor U29364 (N_29364,N_25109,N_26586);
nand U29365 (N_29365,N_26678,N_26188);
nand U29366 (N_29366,N_25921,N_25025);
nor U29367 (N_29367,N_25852,N_26238);
and U29368 (N_29368,N_25412,N_26394);
nor U29369 (N_29369,N_27288,N_26143);
nand U29370 (N_29370,N_27260,N_26206);
or U29371 (N_29371,N_27179,N_26152);
and U29372 (N_29372,N_25418,N_27147);
nor U29373 (N_29373,N_25142,N_26037);
or U29374 (N_29374,N_25577,N_26105);
or U29375 (N_29375,N_26707,N_26637);
xnor U29376 (N_29376,N_26034,N_26971);
nor U29377 (N_29377,N_25950,N_25354);
nor U29378 (N_29378,N_25439,N_25519);
xnor U29379 (N_29379,N_25701,N_25931);
or U29380 (N_29380,N_26828,N_25889);
nand U29381 (N_29381,N_27221,N_26941);
nor U29382 (N_29382,N_25278,N_25997);
and U29383 (N_29383,N_25886,N_26574);
and U29384 (N_29384,N_26595,N_26400);
or U29385 (N_29385,N_26234,N_27487);
and U29386 (N_29386,N_26643,N_26375);
nor U29387 (N_29387,N_27354,N_25423);
nor U29388 (N_29388,N_25898,N_26610);
nor U29389 (N_29389,N_25305,N_26672);
nand U29390 (N_29390,N_25403,N_25852);
nor U29391 (N_29391,N_25222,N_25849);
and U29392 (N_29392,N_26351,N_25669);
or U29393 (N_29393,N_26184,N_25756);
nand U29394 (N_29394,N_25752,N_27439);
nand U29395 (N_29395,N_26778,N_27399);
or U29396 (N_29396,N_26827,N_27432);
nand U29397 (N_29397,N_26867,N_26246);
xnor U29398 (N_29398,N_26719,N_26887);
nand U29399 (N_29399,N_25979,N_25694);
and U29400 (N_29400,N_27308,N_27321);
and U29401 (N_29401,N_25034,N_25537);
xnor U29402 (N_29402,N_25746,N_26503);
nor U29403 (N_29403,N_27311,N_26744);
nand U29404 (N_29404,N_26281,N_25875);
xnor U29405 (N_29405,N_25978,N_27453);
or U29406 (N_29406,N_26194,N_27243);
nor U29407 (N_29407,N_25816,N_27491);
or U29408 (N_29408,N_27179,N_27437);
or U29409 (N_29409,N_26054,N_27138);
or U29410 (N_29410,N_26728,N_25641);
nor U29411 (N_29411,N_26190,N_25942);
and U29412 (N_29412,N_25017,N_26467);
nor U29413 (N_29413,N_25006,N_25754);
nor U29414 (N_29414,N_25425,N_25416);
nor U29415 (N_29415,N_26919,N_25570);
and U29416 (N_29416,N_27241,N_27042);
nand U29417 (N_29417,N_26046,N_25738);
and U29418 (N_29418,N_26157,N_26093);
and U29419 (N_29419,N_26756,N_26303);
nor U29420 (N_29420,N_27040,N_27498);
and U29421 (N_29421,N_25761,N_27293);
nor U29422 (N_29422,N_26579,N_25809);
or U29423 (N_29423,N_27324,N_26079);
or U29424 (N_29424,N_26847,N_26099);
or U29425 (N_29425,N_25884,N_25881);
xnor U29426 (N_29426,N_25665,N_26178);
or U29427 (N_29427,N_27228,N_25788);
nor U29428 (N_29428,N_25162,N_26986);
or U29429 (N_29429,N_27184,N_25831);
or U29430 (N_29430,N_27344,N_26154);
and U29431 (N_29431,N_26031,N_26315);
nor U29432 (N_29432,N_26674,N_25830);
nand U29433 (N_29433,N_26717,N_25515);
and U29434 (N_29434,N_26465,N_25756);
nand U29435 (N_29435,N_25934,N_26766);
and U29436 (N_29436,N_25410,N_25323);
xnor U29437 (N_29437,N_25435,N_25309);
or U29438 (N_29438,N_25842,N_26957);
nand U29439 (N_29439,N_26447,N_25012);
or U29440 (N_29440,N_25701,N_25874);
or U29441 (N_29441,N_25633,N_25714);
nand U29442 (N_29442,N_25887,N_26815);
and U29443 (N_29443,N_26761,N_25763);
and U29444 (N_29444,N_27181,N_25059);
nand U29445 (N_29445,N_25691,N_26077);
nand U29446 (N_29446,N_26935,N_25266);
xor U29447 (N_29447,N_26358,N_26018);
and U29448 (N_29448,N_25585,N_25251);
or U29449 (N_29449,N_26286,N_26229);
and U29450 (N_29450,N_26890,N_26490);
xnor U29451 (N_29451,N_26380,N_27221);
or U29452 (N_29452,N_25268,N_27412);
nand U29453 (N_29453,N_25837,N_26588);
nand U29454 (N_29454,N_27308,N_26812);
nand U29455 (N_29455,N_25218,N_26285);
nor U29456 (N_29456,N_26357,N_26957);
or U29457 (N_29457,N_25688,N_26610);
or U29458 (N_29458,N_26874,N_26632);
nand U29459 (N_29459,N_25405,N_26265);
or U29460 (N_29460,N_25941,N_25538);
nor U29461 (N_29461,N_26205,N_25390);
nor U29462 (N_29462,N_26964,N_27231);
or U29463 (N_29463,N_25863,N_25355);
and U29464 (N_29464,N_26812,N_26421);
or U29465 (N_29465,N_25957,N_26622);
nand U29466 (N_29466,N_26477,N_25367);
and U29467 (N_29467,N_27051,N_26061);
nand U29468 (N_29468,N_25814,N_25533);
and U29469 (N_29469,N_25419,N_27062);
or U29470 (N_29470,N_26812,N_25008);
nor U29471 (N_29471,N_25200,N_26894);
and U29472 (N_29472,N_25129,N_26232);
and U29473 (N_29473,N_26209,N_27140);
xnor U29474 (N_29474,N_26068,N_25945);
or U29475 (N_29475,N_26902,N_25578);
nand U29476 (N_29476,N_26191,N_26789);
nor U29477 (N_29477,N_25700,N_27044);
or U29478 (N_29478,N_26871,N_25973);
and U29479 (N_29479,N_25038,N_25716);
nand U29480 (N_29480,N_25205,N_27437);
or U29481 (N_29481,N_25995,N_27268);
or U29482 (N_29482,N_27175,N_26192);
nand U29483 (N_29483,N_26472,N_27201);
and U29484 (N_29484,N_25473,N_26945);
nor U29485 (N_29485,N_26091,N_26311);
or U29486 (N_29486,N_25553,N_25126);
and U29487 (N_29487,N_26160,N_26655);
nand U29488 (N_29488,N_25996,N_26824);
and U29489 (N_29489,N_26464,N_26833);
and U29490 (N_29490,N_26155,N_26498);
nor U29491 (N_29491,N_26173,N_26878);
xnor U29492 (N_29492,N_25040,N_25660);
nand U29493 (N_29493,N_25559,N_26695);
and U29494 (N_29494,N_26109,N_25857);
and U29495 (N_29495,N_27046,N_25677);
and U29496 (N_29496,N_27310,N_25186);
xnor U29497 (N_29497,N_26003,N_25215);
nand U29498 (N_29498,N_25718,N_25857);
or U29499 (N_29499,N_27163,N_27377);
and U29500 (N_29500,N_25701,N_27411);
and U29501 (N_29501,N_26000,N_26614);
nand U29502 (N_29502,N_26585,N_27313);
or U29503 (N_29503,N_25643,N_25732);
and U29504 (N_29504,N_26087,N_25005);
and U29505 (N_29505,N_26625,N_25316);
nand U29506 (N_29506,N_25073,N_25929);
and U29507 (N_29507,N_26007,N_26122);
and U29508 (N_29508,N_25239,N_25579);
nand U29509 (N_29509,N_25128,N_26829);
or U29510 (N_29510,N_26400,N_25527);
nor U29511 (N_29511,N_26552,N_25817);
or U29512 (N_29512,N_26546,N_26333);
xnor U29513 (N_29513,N_25113,N_27382);
nor U29514 (N_29514,N_26159,N_25722);
and U29515 (N_29515,N_26125,N_26990);
and U29516 (N_29516,N_27318,N_25277);
nand U29517 (N_29517,N_26769,N_26246);
nand U29518 (N_29518,N_25707,N_25161);
nor U29519 (N_29519,N_25135,N_26616);
nand U29520 (N_29520,N_27483,N_25255);
nand U29521 (N_29521,N_26136,N_26617);
nor U29522 (N_29522,N_26990,N_25343);
nor U29523 (N_29523,N_26691,N_25571);
or U29524 (N_29524,N_25051,N_25740);
nand U29525 (N_29525,N_26360,N_27099);
and U29526 (N_29526,N_26807,N_26254);
or U29527 (N_29527,N_27163,N_25997);
nor U29528 (N_29528,N_26645,N_27067);
nand U29529 (N_29529,N_27197,N_26859);
and U29530 (N_29530,N_26855,N_26360);
nor U29531 (N_29531,N_25493,N_25934);
or U29532 (N_29532,N_25163,N_25408);
nor U29533 (N_29533,N_25863,N_25955);
or U29534 (N_29534,N_27096,N_25729);
nor U29535 (N_29535,N_25965,N_27146);
nand U29536 (N_29536,N_25814,N_27140);
or U29537 (N_29537,N_25890,N_26053);
and U29538 (N_29538,N_25124,N_26601);
and U29539 (N_29539,N_25247,N_27451);
or U29540 (N_29540,N_26641,N_26460);
nor U29541 (N_29541,N_27118,N_26158);
or U29542 (N_29542,N_25799,N_26008);
nor U29543 (N_29543,N_26287,N_25677);
nor U29544 (N_29544,N_26231,N_27421);
nor U29545 (N_29545,N_27480,N_25620);
xor U29546 (N_29546,N_26051,N_25504);
or U29547 (N_29547,N_26544,N_25536);
or U29548 (N_29548,N_27486,N_25190);
and U29549 (N_29549,N_25686,N_25042);
and U29550 (N_29550,N_25780,N_27070);
nor U29551 (N_29551,N_26846,N_25772);
or U29552 (N_29552,N_27338,N_27312);
or U29553 (N_29553,N_25775,N_26073);
nand U29554 (N_29554,N_25210,N_25645);
nor U29555 (N_29555,N_25681,N_27273);
and U29556 (N_29556,N_25008,N_25670);
or U29557 (N_29557,N_26307,N_25681);
nor U29558 (N_29558,N_27491,N_26378);
nand U29559 (N_29559,N_25435,N_26353);
nor U29560 (N_29560,N_26522,N_27421);
nand U29561 (N_29561,N_26882,N_25332);
or U29562 (N_29562,N_27061,N_27153);
nor U29563 (N_29563,N_27485,N_26464);
or U29564 (N_29564,N_26567,N_26972);
nor U29565 (N_29565,N_27108,N_25214);
nor U29566 (N_29566,N_26822,N_27102);
nor U29567 (N_29567,N_26342,N_26675);
and U29568 (N_29568,N_25510,N_26640);
xnor U29569 (N_29569,N_25680,N_26750);
nand U29570 (N_29570,N_27287,N_25013);
nand U29571 (N_29571,N_26263,N_27228);
nand U29572 (N_29572,N_25283,N_26558);
and U29573 (N_29573,N_26279,N_25204);
nand U29574 (N_29574,N_26977,N_25125);
nor U29575 (N_29575,N_25371,N_26974);
nand U29576 (N_29576,N_26544,N_25027);
nor U29577 (N_29577,N_26753,N_25534);
or U29578 (N_29578,N_27241,N_27063);
nor U29579 (N_29579,N_26125,N_25609);
or U29580 (N_29580,N_25647,N_25571);
nor U29581 (N_29581,N_26840,N_27266);
or U29582 (N_29582,N_26668,N_25109);
nor U29583 (N_29583,N_26608,N_25003);
nand U29584 (N_29584,N_26332,N_25624);
or U29585 (N_29585,N_27304,N_27258);
or U29586 (N_29586,N_25442,N_25797);
nor U29587 (N_29587,N_26191,N_27221);
or U29588 (N_29588,N_25305,N_27329);
nor U29589 (N_29589,N_25503,N_26792);
nand U29590 (N_29590,N_25694,N_27422);
nor U29591 (N_29591,N_26548,N_25943);
nand U29592 (N_29592,N_25537,N_27044);
and U29593 (N_29593,N_25099,N_26299);
nor U29594 (N_29594,N_27400,N_25268);
nand U29595 (N_29595,N_26424,N_26921);
nand U29596 (N_29596,N_26794,N_26759);
and U29597 (N_29597,N_25234,N_25084);
xnor U29598 (N_29598,N_27213,N_25503);
nand U29599 (N_29599,N_26243,N_27371);
nor U29600 (N_29600,N_27272,N_25279);
nand U29601 (N_29601,N_25282,N_25214);
nand U29602 (N_29602,N_26188,N_25125);
and U29603 (N_29603,N_26811,N_25736);
nor U29604 (N_29604,N_25733,N_26002);
and U29605 (N_29605,N_26484,N_25528);
xor U29606 (N_29606,N_26442,N_25751);
or U29607 (N_29607,N_25564,N_25235);
nand U29608 (N_29608,N_25195,N_25280);
nand U29609 (N_29609,N_25027,N_26802);
nor U29610 (N_29610,N_25216,N_25720);
and U29611 (N_29611,N_26557,N_27008);
and U29612 (N_29612,N_26370,N_27336);
nand U29613 (N_29613,N_26436,N_25177);
and U29614 (N_29614,N_26861,N_26534);
and U29615 (N_29615,N_27132,N_26589);
and U29616 (N_29616,N_27173,N_25581);
and U29617 (N_29617,N_25656,N_27071);
nand U29618 (N_29618,N_25751,N_25967);
xnor U29619 (N_29619,N_26673,N_25539);
or U29620 (N_29620,N_27078,N_26496);
xnor U29621 (N_29621,N_25316,N_25473);
nand U29622 (N_29622,N_25773,N_25671);
or U29623 (N_29623,N_26691,N_26346);
nor U29624 (N_29624,N_27125,N_25700);
xor U29625 (N_29625,N_25438,N_26902);
and U29626 (N_29626,N_25569,N_26973);
nor U29627 (N_29627,N_25274,N_25429);
or U29628 (N_29628,N_26564,N_27098);
nand U29629 (N_29629,N_25748,N_25141);
xor U29630 (N_29630,N_25303,N_26795);
nor U29631 (N_29631,N_26144,N_25953);
and U29632 (N_29632,N_25470,N_25018);
or U29633 (N_29633,N_25740,N_26256);
nand U29634 (N_29634,N_27185,N_26115);
nand U29635 (N_29635,N_26858,N_26987);
nor U29636 (N_29636,N_27024,N_27353);
and U29637 (N_29637,N_26548,N_25848);
nor U29638 (N_29638,N_27205,N_27317);
nand U29639 (N_29639,N_26694,N_27070);
and U29640 (N_29640,N_26664,N_27378);
or U29641 (N_29641,N_25118,N_25399);
or U29642 (N_29642,N_25072,N_25170);
nand U29643 (N_29643,N_27406,N_26011);
or U29644 (N_29644,N_26221,N_26568);
or U29645 (N_29645,N_25265,N_25596);
or U29646 (N_29646,N_25515,N_27364);
and U29647 (N_29647,N_27414,N_27271);
or U29648 (N_29648,N_26461,N_25357);
or U29649 (N_29649,N_25645,N_25354);
nand U29650 (N_29650,N_25590,N_25380);
or U29651 (N_29651,N_25707,N_27279);
nor U29652 (N_29652,N_25282,N_25314);
or U29653 (N_29653,N_25086,N_26573);
nand U29654 (N_29654,N_25267,N_25762);
nor U29655 (N_29655,N_27115,N_26645);
or U29656 (N_29656,N_25554,N_27450);
nand U29657 (N_29657,N_25083,N_26197);
xor U29658 (N_29658,N_26186,N_25421);
nand U29659 (N_29659,N_25512,N_26948);
or U29660 (N_29660,N_25318,N_26107);
nor U29661 (N_29661,N_26492,N_25488);
nor U29662 (N_29662,N_26293,N_26696);
nor U29663 (N_29663,N_25525,N_26416);
and U29664 (N_29664,N_25259,N_26744);
and U29665 (N_29665,N_26266,N_26792);
nand U29666 (N_29666,N_26870,N_25938);
or U29667 (N_29667,N_26070,N_27341);
nand U29668 (N_29668,N_26912,N_27467);
and U29669 (N_29669,N_25877,N_25831);
nand U29670 (N_29670,N_25770,N_27308);
and U29671 (N_29671,N_26513,N_26504);
nand U29672 (N_29672,N_27497,N_26684);
and U29673 (N_29673,N_26134,N_26659);
nand U29674 (N_29674,N_27237,N_26804);
nand U29675 (N_29675,N_25175,N_25727);
or U29676 (N_29676,N_26643,N_25273);
nand U29677 (N_29677,N_26454,N_26498);
nor U29678 (N_29678,N_26039,N_26712);
nor U29679 (N_29679,N_27459,N_26017);
or U29680 (N_29680,N_26421,N_27366);
nor U29681 (N_29681,N_25591,N_25220);
nor U29682 (N_29682,N_25522,N_25984);
xor U29683 (N_29683,N_26682,N_25726);
nand U29684 (N_29684,N_26563,N_25471);
nor U29685 (N_29685,N_27099,N_25657);
or U29686 (N_29686,N_25736,N_26128);
and U29687 (N_29687,N_26577,N_26370);
nor U29688 (N_29688,N_26571,N_26289);
nor U29689 (N_29689,N_25337,N_27134);
nand U29690 (N_29690,N_26341,N_25156);
and U29691 (N_29691,N_25826,N_26430);
or U29692 (N_29692,N_26444,N_27012);
and U29693 (N_29693,N_25404,N_27322);
nand U29694 (N_29694,N_27307,N_26057);
nand U29695 (N_29695,N_25630,N_25158);
nand U29696 (N_29696,N_25592,N_26708);
xor U29697 (N_29697,N_25596,N_25494);
or U29698 (N_29698,N_26636,N_25641);
or U29699 (N_29699,N_25580,N_26780);
nor U29700 (N_29700,N_26317,N_27175);
or U29701 (N_29701,N_26923,N_26138);
nand U29702 (N_29702,N_25912,N_26489);
nand U29703 (N_29703,N_25914,N_27291);
nor U29704 (N_29704,N_27071,N_27253);
and U29705 (N_29705,N_25042,N_26826);
nor U29706 (N_29706,N_27468,N_25455);
xor U29707 (N_29707,N_25699,N_26347);
or U29708 (N_29708,N_26232,N_27456);
nor U29709 (N_29709,N_26150,N_27172);
nand U29710 (N_29710,N_26996,N_26875);
nor U29711 (N_29711,N_26756,N_25364);
and U29712 (N_29712,N_26910,N_26487);
xor U29713 (N_29713,N_26481,N_27200);
nand U29714 (N_29714,N_27384,N_26607);
and U29715 (N_29715,N_26799,N_25854);
xor U29716 (N_29716,N_26571,N_25608);
nand U29717 (N_29717,N_25109,N_27277);
nor U29718 (N_29718,N_25669,N_26362);
nor U29719 (N_29719,N_26319,N_26282);
nand U29720 (N_29720,N_25554,N_27229);
and U29721 (N_29721,N_25093,N_27358);
nor U29722 (N_29722,N_27354,N_25362);
or U29723 (N_29723,N_25091,N_26101);
nor U29724 (N_29724,N_26355,N_25111);
nand U29725 (N_29725,N_27033,N_25356);
nor U29726 (N_29726,N_26410,N_26111);
or U29727 (N_29727,N_25455,N_27196);
nor U29728 (N_29728,N_26287,N_25525);
and U29729 (N_29729,N_26819,N_26006);
xnor U29730 (N_29730,N_25178,N_25501);
nor U29731 (N_29731,N_26872,N_27396);
nand U29732 (N_29732,N_25517,N_25957);
or U29733 (N_29733,N_26738,N_25211);
nor U29734 (N_29734,N_26967,N_26653);
and U29735 (N_29735,N_25125,N_26044);
nor U29736 (N_29736,N_27224,N_26236);
nand U29737 (N_29737,N_25879,N_26747);
nor U29738 (N_29738,N_26196,N_25077);
nand U29739 (N_29739,N_26865,N_26100);
or U29740 (N_29740,N_26419,N_25908);
nor U29741 (N_29741,N_27323,N_25172);
nand U29742 (N_29742,N_26015,N_26268);
or U29743 (N_29743,N_27082,N_25640);
nand U29744 (N_29744,N_26408,N_26943);
or U29745 (N_29745,N_27421,N_26987);
nor U29746 (N_29746,N_25990,N_26954);
nand U29747 (N_29747,N_26580,N_25364);
nand U29748 (N_29748,N_27205,N_25291);
nand U29749 (N_29749,N_26688,N_27389);
and U29750 (N_29750,N_25292,N_27216);
nand U29751 (N_29751,N_25327,N_26012);
or U29752 (N_29752,N_25254,N_26596);
or U29753 (N_29753,N_25644,N_27452);
and U29754 (N_29754,N_25735,N_27146);
or U29755 (N_29755,N_25108,N_25762);
and U29756 (N_29756,N_26215,N_26950);
and U29757 (N_29757,N_25436,N_25443);
or U29758 (N_29758,N_26531,N_26378);
or U29759 (N_29759,N_26824,N_25319);
nand U29760 (N_29760,N_27326,N_26899);
nor U29761 (N_29761,N_27006,N_27012);
xnor U29762 (N_29762,N_26905,N_26270);
nor U29763 (N_29763,N_26727,N_26634);
and U29764 (N_29764,N_26633,N_27292);
nor U29765 (N_29765,N_26860,N_25622);
xor U29766 (N_29766,N_25286,N_26192);
nor U29767 (N_29767,N_26581,N_25662);
nor U29768 (N_29768,N_26067,N_26151);
nor U29769 (N_29769,N_26123,N_26315);
and U29770 (N_29770,N_26565,N_25631);
or U29771 (N_29771,N_26585,N_25601);
nand U29772 (N_29772,N_26181,N_26571);
nor U29773 (N_29773,N_26968,N_25730);
nand U29774 (N_29774,N_25347,N_25014);
nand U29775 (N_29775,N_26790,N_25331);
or U29776 (N_29776,N_26292,N_27121);
and U29777 (N_29777,N_25436,N_25039);
and U29778 (N_29778,N_25346,N_26572);
nand U29779 (N_29779,N_26662,N_27004);
or U29780 (N_29780,N_25606,N_27247);
nand U29781 (N_29781,N_26947,N_26301);
xor U29782 (N_29782,N_25899,N_25235);
nor U29783 (N_29783,N_25969,N_26622);
and U29784 (N_29784,N_26613,N_27091);
xor U29785 (N_29785,N_26205,N_26053);
or U29786 (N_29786,N_26190,N_26631);
nand U29787 (N_29787,N_27281,N_25008);
nor U29788 (N_29788,N_26836,N_27199);
nor U29789 (N_29789,N_27282,N_25643);
or U29790 (N_29790,N_26137,N_25462);
or U29791 (N_29791,N_27355,N_27144);
or U29792 (N_29792,N_26017,N_25173);
nor U29793 (N_29793,N_25550,N_26892);
nor U29794 (N_29794,N_25894,N_26238);
and U29795 (N_29795,N_26747,N_25858);
xnor U29796 (N_29796,N_25602,N_26099);
or U29797 (N_29797,N_26362,N_26218);
xnor U29798 (N_29798,N_25344,N_25384);
or U29799 (N_29799,N_27180,N_25869);
nor U29800 (N_29800,N_26590,N_26960);
xor U29801 (N_29801,N_27255,N_26643);
nor U29802 (N_29802,N_25413,N_27136);
nand U29803 (N_29803,N_25953,N_26982);
and U29804 (N_29804,N_27135,N_27018);
nor U29805 (N_29805,N_27299,N_26012);
nand U29806 (N_29806,N_25466,N_26036);
or U29807 (N_29807,N_26486,N_27161);
and U29808 (N_29808,N_25897,N_26791);
nand U29809 (N_29809,N_27097,N_27166);
and U29810 (N_29810,N_26203,N_27412);
xor U29811 (N_29811,N_26523,N_27205);
nand U29812 (N_29812,N_26501,N_25033);
nand U29813 (N_29813,N_26033,N_26953);
or U29814 (N_29814,N_26923,N_25617);
nor U29815 (N_29815,N_25711,N_27241);
nand U29816 (N_29816,N_27348,N_25252);
nor U29817 (N_29817,N_27444,N_27341);
or U29818 (N_29818,N_25275,N_26220);
or U29819 (N_29819,N_25476,N_26566);
nand U29820 (N_29820,N_25652,N_26136);
or U29821 (N_29821,N_27328,N_26292);
and U29822 (N_29822,N_26463,N_26725);
or U29823 (N_29823,N_25250,N_25252);
nand U29824 (N_29824,N_26547,N_25664);
nand U29825 (N_29825,N_26646,N_25098);
nor U29826 (N_29826,N_26211,N_26835);
and U29827 (N_29827,N_26003,N_27393);
xnor U29828 (N_29828,N_26381,N_25511);
nand U29829 (N_29829,N_27233,N_27239);
or U29830 (N_29830,N_25415,N_25526);
xor U29831 (N_29831,N_27218,N_25967);
and U29832 (N_29832,N_26584,N_26758);
nand U29833 (N_29833,N_25852,N_27445);
or U29834 (N_29834,N_26984,N_26134);
nand U29835 (N_29835,N_26772,N_27195);
xor U29836 (N_29836,N_27072,N_25399);
xnor U29837 (N_29837,N_26514,N_27323);
nand U29838 (N_29838,N_27391,N_26084);
or U29839 (N_29839,N_27293,N_26936);
xor U29840 (N_29840,N_26161,N_25820);
nor U29841 (N_29841,N_25793,N_26410);
and U29842 (N_29842,N_25324,N_25711);
and U29843 (N_29843,N_26450,N_25958);
nand U29844 (N_29844,N_25376,N_26112);
and U29845 (N_29845,N_25029,N_27260);
nand U29846 (N_29846,N_25332,N_26960);
or U29847 (N_29847,N_26100,N_25455);
and U29848 (N_29848,N_27379,N_26381);
nor U29849 (N_29849,N_26504,N_25485);
nor U29850 (N_29850,N_27399,N_26070);
or U29851 (N_29851,N_27221,N_25050);
nor U29852 (N_29852,N_26625,N_25461);
and U29853 (N_29853,N_25622,N_27377);
nor U29854 (N_29854,N_27481,N_27289);
xnor U29855 (N_29855,N_26192,N_25992);
nor U29856 (N_29856,N_26247,N_27404);
or U29857 (N_29857,N_27098,N_26087);
nand U29858 (N_29858,N_25557,N_26811);
or U29859 (N_29859,N_25133,N_25401);
nand U29860 (N_29860,N_26582,N_27172);
or U29861 (N_29861,N_27287,N_26676);
nand U29862 (N_29862,N_26549,N_26535);
nand U29863 (N_29863,N_25321,N_25948);
nor U29864 (N_29864,N_25160,N_27027);
nor U29865 (N_29865,N_25478,N_25152);
nor U29866 (N_29866,N_26856,N_27121);
nor U29867 (N_29867,N_25901,N_27414);
xnor U29868 (N_29868,N_25264,N_26847);
xnor U29869 (N_29869,N_26569,N_25152);
and U29870 (N_29870,N_25715,N_25975);
nor U29871 (N_29871,N_26126,N_26818);
or U29872 (N_29872,N_25569,N_26713);
and U29873 (N_29873,N_25887,N_26347);
and U29874 (N_29874,N_26703,N_25748);
or U29875 (N_29875,N_25376,N_26434);
nor U29876 (N_29876,N_25343,N_26506);
xnor U29877 (N_29877,N_25005,N_27372);
or U29878 (N_29878,N_26152,N_25064);
nor U29879 (N_29879,N_25238,N_26219);
xor U29880 (N_29880,N_26384,N_25698);
nand U29881 (N_29881,N_25506,N_25498);
nor U29882 (N_29882,N_26759,N_25741);
or U29883 (N_29883,N_25240,N_26185);
nand U29884 (N_29884,N_25487,N_26223);
nand U29885 (N_29885,N_27098,N_25189);
and U29886 (N_29886,N_26878,N_25434);
nor U29887 (N_29887,N_25366,N_27325);
nor U29888 (N_29888,N_27137,N_27227);
nor U29889 (N_29889,N_25499,N_25208);
and U29890 (N_29890,N_26539,N_26294);
or U29891 (N_29891,N_25100,N_27307);
or U29892 (N_29892,N_26782,N_25770);
nor U29893 (N_29893,N_25879,N_27498);
nor U29894 (N_29894,N_27050,N_25832);
or U29895 (N_29895,N_25474,N_25084);
and U29896 (N_29896,N_27457,N_26085);
nand U29897 (N_29897,N_25534,N_25986);
or U29898 (N_29898,N_27378,N_26097);
nor U29899 (N_29899,N_26178,N_25719);
and U29900 (N_29900,N_25662,N_25877);
or U29901 (N_29901,N_25419,N_26649);
nor U29902 (N_29902,N_26208,N_25335);
nor U29903 (N_29903,N_26698,N_27066);
or U29904 (N_29904,N_25588,N_26137);
nand U29905 (N_29905,N_27403,N_26161);
nor U29906 (N_29906,N_25836,N_25335);
or U29907 (N_29907,N_26062,N_26956);
nor U29908 (N_29908,N_26718,N_26952);
nor U29909 (N_29909,N_25386,N_26710);
or U29910 (N_29910,N_25305,N_27122);
xor U29911 (N_29911,N_25238,N_27094);
xor U29912 (N_29912,N_27484,N_27080);
nand U29913 (N_29913,N_27122,N_26126);
nor U29914 (N_29914,N_26909,N_27024);
nand U29915 (N_29915,N_26063,N_25548);
or U29916 (N_29916,N_25442,N_26220);
or U29917 (N_29917,N_27367,N_25181);
xor U29918 (N_29918,N_25762,N_27152);
and U29919 (N_29919,N_27004,N_25719);
nor U29920 (N_29920,N_25088,N_27158);
and U29921 (N_29921,N_25795,N_25851);
or U29922 (N_29922,N_25756,N_25652);
and U29923 (N_29923,N_26496,N_25501);
or U29924 (N_29924,N_26635,N_26436);
or U29925 (N_29925,N_26098,N_25777);
nor U29926 (N_29926,N_25159,N_26623);
or U29927 (N_29927,N_27302,N_26080);
or U29928 (N_29928,N_26597,N_25314);
nor U29929 (N_29929,N_27130,N_26479);
nand U29930 (N_29930,N_25172,N_25781);
nand U29931 (N_29931,N_26202,N_26026);
and U29932 (N_29932,N_27252,N_26831);
and U29933 (N_29933,N_26936,N_25282);
and U29934 (N_29934,N_26686,N_26269);
nand U29935 (N_29935,N_27047,N_27017);
nor U29936 (N_29936,N_25746,N_26607);
nor U29937 (N_29937,N_25158,N_27235);
nor U29938 (N_29938,N_27288,N_27470);
xnor U29939 (N_29939,N_26493,N_26081);
or U29940 (N_29940,N_26567,N_26069);
xor U29941 (N_29941,N_27203,N_25090);
nand U29942 (N_29942,N_26414,N_26745);
nor U29943 (N_29943,N_27338,N_25336);
nand U29944 (N_29944,N_27419,N_25050);
or U29945 (N_29945,N_25440,N_27037);
or U29946 (N_29946,N_27240,N_27460);
or U29947 (N_29947,N_26808,N_26966);
nor U29948 (N_29948,N_27276,N_25809);
nand U29949 (N_29949,N_26833,N_27411);
or U29950 (N_29950,N_26830,N_26782);
or U29951 (N_29951,N_27238,N_26611);
and U29952 (N_29952,N_25035,N_26114);
or U29953 (N_29953,N_25186,N_26627);
or U29954 (N_29954,N_26897,N_27466);
or U29955 (N_29955,N_26150,N_26989);
nand U29956 (N_29956,N_26695,N_26123);
nor U29957 (N_29957,N_25665,N_27419);
xnor U29958 (N_29958,N_27137,N_26966);
nand U29959 (N_29959,N_27272,N_27367);
nor U29960 (N_29960,N_26670,N_26517);
nor U29961 (N_29961,N_27160,N_25951);
or U29962 (N_29962,N_26887,N_27350);
nor U29963 (N_29963,N_26574,N_26718);
nor U29964 (N_29964,N_26600,N_25446);
or U29965 (N_29965,N_26151,N_26618);
or U29966 (N_29966,N_26183,N_27298);
and U29967 (N_29967,N_25573,N_26852);
nor U29968 (N_29968,N_25522,N_25979);
nand U29969 (N_29969,N_26191,N_27111);
and U29970 (N_29970,N_25199,N_26740);
or U29971 (N_29971,N_27493,N_25456);
and U29972 (N_29972,N_25022,N_27178);
nand U29973 (N_29973,N_26434,N_27273);
or U29974 (N_29974,N_26949,N_25682);
nand U29975 (N_29975,N_25503,N_27370);
nor U29976 (N_29976,N_26595,N_25022);
and U29977 (N_29977,N_25162,N_25987);
nor U29978 (N_29978,N_25085,N_27318);
nand U29979 (N_29979,N_27405,N_25008);
or U29980 (N_29980,N_25736,N_27371);
nor U29981 (N_29981,N_26276,N_25646);
xor U29982 (N_29982,N_26876,N_25603);
nand U29983 (N_29983,N_26132,N_26347);
and U29984 (N_29984,N_25971,N_25922);
nand U29985 (N_29985,N_27350,N_25198);
and U29986 (N_29986,N_26855,N_25182);
and U29987 (N_29987,N_25837,N_26318);
or U29988 (N_29988,N_26191,N_26784);
and U29989 (N_29989,N_26456,N_25596);
and U29990 (N_29990,N_26742,N_26467);
nor U29991 (N_29991,N_25879,N_27388);
or U29992 (N_29992,N_25944,N_26526);
nand U29993 (N_29993,N_27372,N_27321);
nand U29994 (N_29994,N_26546,N_25321);
nor U29995 (N_29995,N_25389,N_25836);
and U29996 (N_29996,N_25670,N_25939);
and U29997 (N_29997,N_26310,N_25096);
or U29998 (N_29998,N_27362,N_27026);
or U29999 (N_29999,N_25721,N_27265);
nor U30000 (N_30000,N_28379,N_29990);
and U30001 (N_30001,N_29168,N_28195);
nor U30002 (N_30002,N_28920,N_28155);
nor U30003 (N_30003,N_28216,N_28338);
and U30004 (N_30004,N_29665,N_27509);
or U30005 (N_30005,N_28954,N_29087);
and U30006 (N_30006,N_27659,N_29238);
and U30007 (N_30007,N_27913,N_29541);
nand U30008 (N_30008,N_28905,N_29848);
or U30009 (N_30009,N_29020,N_29799);
nor U30010 (N_30010,N_28450,N_29893);
or U30011 (N_30011,N_29525,N_27822);
or U30012 (N_30012,N_29490,N_29842);
and U30013 (N_30013,N_29270,N_29171);
and U30014 (N_30014,N_29948,N_28213);
and U30015 (N_30015,N_29755,N_29573);
nand U30016 (N_30016,N_29607,N_29539);
and U30017 (N_30017,N_28381,N_29899);
nor U30018 (N_30018,N_28826,N_29666);
or U30019 (N_30019,N_29350,N_29521);
and U30020 (N_30020,N_28491,N_29392);
xor U30021 (N_30021,N_29152,N_28459);
or U30022 (N_30022,N_29697,N_28031);
nand U30023 (N_30023,N_29069,N_28192);
or U30024 (N_30024,N_29526,N_27943);
and U30025 (N_30025,N_28142,N_29482);
and U30026 (N_30026,N_28964,N_28750);
nand U30027 (N_30027,N_29940,N_28460);
and U30028 (N_30028,N_29113,N_27647);
nor U30029 (N_30029,N_29636,N_29680);
and U30030 (N_30030,N_29324,N_27761);
nand U30031 (N_30031,N_29244,N_28711);
nor U30032 (N_30032,N_29172,N_29655);
and U30033 (N_30033,N_28896,N_29742);
nand U30034 (N_30034,N_29690,N_29094);
or U30035 (N_30035,N_28997,N_28669);
xnor U30036 (N_30036,N_28691,N_27724);
xnor U30037 (N_30037,N_28341,N_28180);
or U30038 (N_30038,N_29040,N_27637);
and U30039 (N_30039,N_29519,N_28360);
and U30040 (N_30040,N_27734,N_28435);
or U30041 (N_30041,N_28787,N_27903);
xnor U30042 (N_30042,N_29207,N_28891);
and U30043 (N_30043,N_28495,N_29986);
nand U30044 (N_30044,N_29248,N_28919);
nand U30045 (N_30045,N_28267,N_28064);
nand U30046 (N_30046,N_28694,N_28413);
or U30047 (N_30047,N_28453,N_28193);
and U30048 (N_30048,N_28825,N_28373);
nor U30049 (N_30049,N_27936,N_29272);
nand U30050 (N_30050,N_28377,N_28113);
nor U30051 (N_30051,N_28148,N_28418);
and U30052 (N_30052,N_28440,N_27571);
or U30053 (N_30053,N_27881,N_28152);
nand U30054 (N_30054,N_27671,N_28956);
nor U30055 (N_30055,N_29016,N_27833);
nor U30056 (N_30056,N_28422,N_29089);
nor U30057 (N_30057,N_29782,N_29922);
or U30058 (N_30058,N_28281,N_27969);
or U30059 (N_30059,N_27544,N_28108);
nand U30060 (N_30060,N_28587,N_27521);
or U30061 (N_30061,N_29745,N_28976);
nor U30062 (N_30062,N_29117,N_29076);
or U30063 (N_30063,N_27743,N_28814);
nand U30064 (N_30064,N_28786,N_27829);
nor U30065 (N_30065,N_27744,N_29875);
or U30066 (N_30066,N_28952,N_29748);
or U30067 (N_30067,N_29141,N_29304);
nor U30068 (N_30068,N_29174,N_28176);
nand U30069 (N_30069,N_29714,N_28808);
or U30070 (N_30070,N_28465,N_28716);
and U30071 (N_30071,N_28126,N_27918);
nor U30072 (N_30072,N_29378,N_27548);
nand U30073 (N_30073,N_27774,N_29488);
nor U30074 (N_30074,N_28878,N_29780);
nor U30075 (N_30075,N_29105,N_29943);
or U30076 (N_30076,N_28145,N_27512);
nand U30077 (N_30077,N_28405,N_27648);
nor U30078 (N_30078,N_27631,N_27565);
nand U30079 (N_30079,N_29630,N_27755);
or U30080 (N_30080,N_28452,N_27554);
nor U30081 (N_30081,N_29142,N_29375);
nor U30082 (N_30082,N_29284,N_29215);
or U30083 (N_30083,N_27530,N_29370);
and U30084 (N_30084,N_27793,N_27590);
and U30085 (N_30085,N_29546,N_29312);
nor U30086 (N_30086,N_27987,N_28348);
nand U30087 (N_30087,N_28770,N_28498);
or U30088 (N_30088,N_29461,N_28873);
nand U30089 (N_30089,N_28563,N_29717);
nor U30090 (N_30090,N_29879,N_29432);
or U30091 (N_30091,N_29837,N_27906);
or U30092 (N_30092,N_29014,N_27666);
nand U30093 (N_30093,N_27777,N_28950);
nand U30094 (N_30094,N_28749,N_27873);
nand U30095 (N_30095,N_29718,N_29416);
nand U30096 (N_30096,N_28758,N_28048);
nand U30097 (N_30097,N_27775,N_28332);
nand U30098 (N_30098,N_29715,N_29209);
nand U30099 (N_30099,N_28067,N_28893);
and U30100 (N_30100,N_28911,N_28886);
or U30101 (N_30101,N_29464,N_28904);
and U30102 (N_30102,N_28899,N_27596);
nor U30103 (N_30103,N_28778,N_28820);
or U30104 (N_30104,N_27961,N_28625);
xor U30105 (N_30105,N_28722,N_28871);
nor U30106 (N_30106,N_27668,N_27947);
nor U30107 (N_30107,N_29769,N_29423);
xnor U30108 (N_30108,N_27506,N_29812);
or U30109 (N_30109,N_29388,N_28185);
and U30110 (N_30110,N_29263,N_29682);
or U30111 (N_30111,N_28471,N_29628);
nand U30112 (N_30112,N_27963,N_29779);
xnor U30113 (N_30113,N_28647,N_28224);
nor U30114 (N_30114,N_28497,N_28368);
nand U30115 (N_30115,N_27799,N_28071);
xor U30116 (N_30116,N_28649,N_27992);
xnor U30117 (N_30117,N_28564,N_29027);
or U30118 (N_30118,N_28857,N_28507);
nand U30119 (N_30119,N_29055,N_28553);
nor U30120 (N_30120,N_27713,N_27900);
and U30121 (N_30121,N_28828,N_29723);
and U30122 (N_30122,N_29686,N_29993);
nor U30123 (N_30123,N_28310,N_27733);
nand U30124 (N_30124,N_29951,N_29969);
nand U30125 (N_30125,N_27818,N_29957);
nand U30126 (N_30126,N_29889,N_27875);
nand U30127 (N_30127,N_28057,N_29906);
and U30128 (N_30128,N_29140,N_29491);
and U30129 (N_30129,N_27846,N_28539);
or U30130 (N_30130,N_29753,N_28854);
xor U30131 (N_30131,N_28050,N_28325);
nor U30132 (N_30132,N_27682,N_28755);
nor U30133 (N_30133,N_28703,N_28385);
nand U30134 (N_30134,N_27798,N_29676);
nor U30135 (N_30135,N_28592,N_28922);
and U30136 (N_30136,N_29472,N_28081);
nor U30137 (N_30137,N_28033,N_28679);
and U30138 (N_30138,N_28913,N_28095);
or U30139 (N_30139,N_28372,N_29874);
nand U30140 (N_30140,N_28622,N_28469);
nand U30141 (N_30141,N_27670,N_29817);
nand U30142 (N_30142,N_29162,N_28846);
and U30143 (N_30143,N_27819,N_29219);
and U30144 (N_30144,N_28906,N_27675);
xor U30145 (N_30145,N_29947,N_27653);
or U30146 (N_30146,N_29414,N_29732);
nor U30147 (N_30147,N_29281,N_29905);
nor U30148 (N_30148,N_28365,N_27534);
or U30149 (N_30149,N_29548,N_27619);
or U30150 (N_30150,N_28544,N_27537);
nand U30151 (N_30151,N_29394,N_29708);
and U30152 (N_30152,N_28877,N_29317);
or U30153 (N_30153,N_28968,N_29157);
xnor U30154 (N_30154,N_28702,N_28209);
xnor U30155 (N_30155,N_28322,N_29413);
xnor U30156 (N_30156,N_28079,N_29200);
xnor U30157 (N_30157,N_27696,N_28311);
nand U30158 (N_30158,N_27518,N_29455);
or U30159 (N_30159,N_29385,N_29793);
nor U30160 (N_30160,N_27754,N_29195);
and U30161 (N_30161,N_29529,N_27826);
and U30162 (N_30162,N_29599,N_28608);
nand U30163 (N_30163,N_29576,N_29705);
nor U30164 (N_30164,N_29661,N_29012);
nand U30165 (N_30165,N_29685,N_28009);
or U30166 (N_30166,N_28895,N_27885);
xor U30167 (N_30167,N_28940,N_27676);
and U30168 (N_30168,N_28189,N_27847);
nand U30169 (N_30169,N_29329,N_28859);
xnor U30170 (N_30170,N_28797,N_29193);
and U30171 (N_30171,N_28754,N_29429);
and U30172 (N_30172,N_29005,N_29315);
nand U30173 (N_30173,N_28907,N_29347);
and U30174 (N_30174,N_29167,N_27879);
nor U30175 (N_30175,N_27658,N_28593);
or U30176 (N_30176,N_28077,N_27709);
and U30177 (N_30177,N_27551,N_29731);
nand U30178 (N_30178,N_28502,N_29953);
nand U30179 (N_30179,N_27574,N_29321);
or U30180 (N_30180,N_29850,N_28757);
or U30181 (N_30181,N_29306,N_28663);
or U30182 (N_30182,N_29921,N_28936);
and U30183 (N_30183,N_28414,N_28961);
xnor U30184 (N_30184,N_29343,N_29971);
or U30185 (N_30185,N_27964,N_29199);
or U30186 (N_30186,N_27550,N_28784);
xor U30187 (N_30187,N_29447,N_29107);
and U30188 (N_30188,N_28687,N_29448);
or U30189 (N_30189,N_27657,N_27556);
nor U30190 (N_30190,N_29147,N_29358);
or U30191 (N_30191,N_29620,N_29398);
and U30192 (N_30192,N_29866,N_29439);
nor U30193 (N_30193,N_29647,N_27928);
and U30194 (N_30194,N_28041,N_28437);
nor U30195 (N_30195,N_29767,N_28590);
or U30196 (N_30196,N_29043,N_29991);
nor U30197 (N_30197,N_27699,N_29608);
and U30198 (N_30198,N_29499,N_28549);
nor U30199 (N_30199,N_28179,N_28276);
or U30200 (N_30200,N_28366,N_28137);
or U30201 (N_30201,N_29202,N_29417);
xor U30202 (N_30202,N_28205,N_28078);
nand U30203 (N_30203,N_28642,N_28136);
or U30204 (N_30204,N_28163,N_29015);
and U30205 (N_30205,N_27629,N_29872);
nor U30206 (N_30206,N_29565,N_29006);
xor U30207 (N_30207,N_28406,N_29211);
xnor U30208 (N_30208,N_29078,N_29130);
or U30209 (N_30209,N_27684,N_28550);
and U30210 (N_30210,N_29104,N_27807);
or U30211 (N_30211,N_28083,N_27522);
and U30212 (N_30212,N_28329,N_27805);
nand U30213 (N_30213,N_29713,N_27573);
and U30214 (N_30214,N_27971,N_28146);
or U30215 (N_30215,N_27828,N_28287);
xor U30216 (N_30216,N_29273,N_29917);
or U30217 (N_30217,N_27994,N_27929);
or U30218 (N_30218,N_29404,N_27862);
or U30219 (N_30219,N_28259,N_29789);
nor U30220 (N_30220,N_28548,N_29096);
nand U30221 (N_30221,N_27806,N_29696);
xnor U30222 (N_30222,N_28938,N_28234);
nand U30223 (N_30223,N_28845,N_29907);
nor U30224 (N_30224,N_29515,N_27804);
nand U30225 (N_30225,N_27500,N_28352);
nand U30226 (N_30226,N_28164,N_28280);
nand U30227 (N_30227,N_29856,N_29532);
nand U30228 (N_30228,N_29537,N_29367);
xor U30229 (N_30229,N_28836,N_29783);
or U30230 (N_30230,N_28204,N_29758);
and U30231 (N_30231,N_28515,N_28745);
nor U30232 (N_30232,N_29619,N_27718);
xnor U30233 (N_30233,N_29048,N_29438);
and U30234 (N_30234,N_29477,N_28850);
and U30235 (N_30235,N_29282,N_29934);
or U30236 (N_30236,N_28616,N_28959);
xnor U30237 (N_30237,N_28069,N_28951);
nand U30238 (N_30238,N_28229,N_27516);
nor U30239 (N_30239,N_28586,N_28074);
and U30240 (N_30240,N_28781,N_27614);
nor U30241 (N_30241,N_29065,N_28733);
nor U30242 (N_30242,N_28159,N_28852);
nand U30243 (N_30243,N_28288,N_28239);
or U30244 (N_30244,N_28093,N_29924);
or U30245 (N_30245,N_28779,N_29258);
or U30246 (N_30246,N_29859,N_28606);
xnor U30247 (N_30247,N_28504,N_29536);
nor U30248 (N_30248,N_28614,N_28666);
nor U30249 (N_30249,N_27716,N_29695);
nand U30250 (N_30250,N_28926,N_28613);
xor U30251 (N_30251,N_29233,N_27887);
xnor U30252 (N_30252,N_29938,N_29387);
nor U30253 (N_30253,N_27702,N_29977);
or U30254 (N_30254,N_27841,N_27753);
and U30255 (N_30255,N_28639,N_28867);
xor U30256 (N_30256,N_29846,N_28816);
and U30257 (N_30257,N_28979,N_29054);
xnor U30258 (N_30258,N_28034,N_29738);
nor U30259 (N_30259,N_28300,N_29556);
or U30260 (N_30260,N_29833,N_29319);
or U30261 (N_30261,N_28272,N_29929);
nand U30262 (N_30262,N_28402,N_28092);
or U30263 (N_30263,N_29386,N_28110);
nand U30264 (N_30264,N_29442,N_29979);
xor U30265 (N_30265,N_27557,N_28173);
or U30266 (N_30266,N_29898,N_29345);
nand U30267 (N_30267,N_27858,N_29928);
xnor U30268 (N_30268,N_29505,N_27834);
and U30269 (N_30269,N_28753,N_29246);
xor U30270 (N_30270,N_27925,N_29843);
nor U30271 (N_30271,N_29841,N_29533);
nand U30272 (N_30272,N_28088,N_29111);
nor U30273 (N_30273,N_28923,N_27649);
and U30274 (N_30274,N_28391,N_28971);
nor U30275 (N_30275,N_29606,N_28600);
and U30276 (N_30276,N_28449,N_28201);
nand U30277 (N_30277,N_28133,N_28645);
nand U30278 (N_30278,N_28742,N_28432);
nor U30279 (N_30279,N_28257,N_27732);
and U30280 (N_30280,N_27937,N_28851);
nor U30281 (N_30281,N_28350,N_28569);
and U30282 (N_30282,N_29474,N_29310);
nor U30283 (N_30283,N_29108,N_27844);
nor U30284 (N_30284,N_28627,N_28732);
nor U30285 (N_30285,N_29173,N_29585);
nor U30286 (N_30286,N_28918,N_27762);
or U30287 (N_30287,N_29511,N_28063);
or U30288 (N_30288,N_28506,N_28861);
nand U30289 (N_30289,N_27635,N_29944);
or U30290 (N_30290,N_29466,N_27856);
nand U30291 (N_30291,N_29610,N_29641);
nor U30292 (N_30292,N_29545,N_28116);
or U30293 (N_30293,N_28894,N_28783);
and U30294 (N_30294,N_29517,N_27582);
or U30295 (N_30295,N_29510,N_29074);
nor U30296 (N_30296,N_27617,N_27627);
or U30297 (N_30297,N_29895,N_28383);
and U30298 (N_30298,N_27831,N_28358);
nand U30299 (N_30299,N_27687,N_29316);
xor U30300 (N_30300,N_29904,N_28244);
or U30301 (N_30301,N_29425,N_28208);
and U30302 (N_30302,N_28171,N_29884);
nand U30303 (N_30303,N_28611,N_28933);
xnor U30304 (N_30304,N_28010,N_28412);
nor U30305 (N_30305,N_29290,N_29299);
and U30306 (N_30306,N_28865,N_29967);
and U30307 (N_30307,N_29952,N_28874);
nor U30308 (N_30308,N_28141,N_29937);
nor U30309 (N_30309,N_29465,N_28494);
and U30310 (N_30310,N_29954,N_27584);
or U30311 (N_30311,N_27997,N_28935);
and U30312 (N_30312,N_28118,N_28228);
xor U30313 (N_30313,N_28135,N_28247);
nand U30314 (N_30314,N_28217,N_28774);
nand U30315 (N_30315,N_27532,N_29459);
nand U30316 (N_30316,N_28819,N_27698);
nor U30317 (N_30317,N_29145,N_29064);
and U30318 (N_30318,N_28046,N_29662);
nand U30319 (N_30319,N_29920,N_27664);
nor U30320 (N_30320,N_27707,N_28296);
and U30321 (N_30321,N_28393,N_27974);
xor U30322 (N_30322,N_28132,N_29964);
nand U30323 (N_30323,N_28099,N_29287);
and U30324 (N_30324,N_29498,N_28995);
xor U30325 (N_30325,N_28168,N_28517);
or U30326 (N_30326,N_28012,N_29596);
xor U30327 (N_30327,N_28963,N_27673);
nand U30328 (N_30328,N_28076,N_29987);
nand U30329 (N_30329,N_29734,N_28712);
or U30330 (N_30330,N_29419,N_28479);
and U30331 (N_30331,N_27908,N_29369);
nor U30332 (N_30332,N_28104,N_29025);
and U30333 (N_30333,N_29547,N_28640);
or U30334 (N_30334,N_28025,N_27944);
nand U30335 (N_30335,N_29470,N_27787);
nor U30336 (N_30336,N_27926,N_28945);
nor U30337 (N_30337,N_29509,N_29955);
or U30338 (N_30338,N_28051,N_29400);
nand U30339 (N_30339,N_28795,N_29433);
and U30340 (N_30340,N_28170,N_27502);
and U30341 (N_30341,N_28986,N_27514);
nand U30342 (N_30342,N_28085,N_29201);
nand U30343 (N_30343,N_28289,N_29729);
nor U30344 (N_30344,N_27932,N_28036);
and U30345 (N_30345,N_28708,N_29560);
xnor U30346 (N_30346,N_28028,N_28988);
nor U30347 (N_30347,N_28697,N_29518);
nand U30348 (N_30348,N_28771,N_29431);
nor U30349 (N_30349,N_27643,N_27545);
nor U30350 (N_30350,N_29139,N_29513);
and U30351 (N_30351,N_29437,N_29058);
nand U30352 (N_30352,N_28818,N_27977);
xnor U30353 (N_30353,N_27525,N_29935);
nand U30354 (N_30354,N_27857,N_29462);
xor U30355 (N_30355,N_28477,N_27711);
xnor U30356 (N_30356,N_29654,N_29257);
xor U30357 (N_30357,N_29237,N_27731);
xnor U30358 (N_30358,N_27546,N_27622);
and U30359 (N_30359,N_27912,N_28378);
nor U30360 (N_30360,N_27957,N_29653);
nand U30361 (N_30361,N_29741,N_29544);
and U30362 (N_30362,N_28617,N_29503);
xor U30363 (N_30363,N_28880,N_27758);
nor U30364 (N_30364,N_28039,N_27864);
and U30365 (N_30365,N_27983,N_27956);
and U30366 (N_30366,N_28340,N_29227);
nand U30367 (N_30367,N_28603,N_27835);
nor U30368 (N_30368,N_29373,N_28537);
nor U30369 (N_30369,N_28513,N_29881);
or U30370 (N_30370,N_28751,N_28551);
nand U30371 (N_30371,N_27837,N_28618);
xnor U30372 (N_30372,N_28181,N_28972);
xnor U30373 (N_30373,N_28015,N_28572);
xnor U30374 (N_30374,N_28326,N_29134);
xnor U30375 (N_30375,N_27816,N_28261);
or U30376 (N_30376,N_29349,N_28026);
and U30377 (N_30377,N_28726,N_28250);
xor U30378 (N_30378,N_29692,N_28467);
and U30379 (N_30379,N_27786,N_29956);
or U30380 (N_30380,N_27780,N_29452);
nor U30381 (N_30381,N_29053,N_27868);
xor U30382 (N_30382,N_29088,N_27642);
and U30383 (N_30383,N_28804,N_28944);
and U30384 (N_30384,N_28410,N_29249);
and U30385 (N_30385,N_29933,N_28022);
or U30386 (N_30386,N_28652,N_28884);
and U30387 (N_30387,N_29531,N_29289);
or U30388 (N_30388,N_28937,N_27889);
nand U30389 (N_30389,N_28233,N_29808);
nor U30390 (N_30390,N_28474,N_29709);
or U30391 (N_30391,N_28897,N_29426);
xnor U30392 (N_30392,N_28809,N_29985);
nor U30393 (N_30393,N_27503,N_29973);
xnor U30394 (N_30394,N_28457,N_29009);
nor U30395 (N_30395,N_28955,N_29612);
or U30396 (N_30396,N_29232,N_29828);
xnor U30397 (N_30397,N_29772,N_29106);
or U30398 (N_30398,N_27559,N_28243);
nor U30399 (N_30399,N_28002,N_28843);
nor U30400 (N_30400,N_28690,N_28187);
or U30401 (N_30401,N_28744,N_28656);
nor U30402 (N_30402,N_27749,N_28903);
nor U30403 (N_30403,N_27859,N_27691);
nand U30404 (N_30404,N_29327,N_27938);
and U30405 (N_30405,N_28120,N_27638);
nor U30406 (N_30406,N_29376,N_28908);
or U30407 (N_30407,N_29642,N_28473);
and U30408 (N_30408,N_28109,N_29389);
nor U30409 (N_30409,N_29568,N_27549);
or U30410 (N_30410,N_29790,N_29136);
xnor U30411 (N_30411,N_28785,N_28456);
nor U30412 (N_30412,N_29471,N_27511);
or U30413 (N_30413,N_29864,N_28980);
nand U30414 (N_30414,N_27941,N_28594);
or U30415 (N_30415,N_27767,N_28401);
and U30416 (N_30416,N_27730,N_29572);
and U30417 (N_30417,N_29984,N_27607);
and U30418 (N_30418,N_28395,N_28914);
nor U30419 (N_30419,N_28178,N_28314);
nand U30420 (N_30420,N_28162,N_29514);
and U30421 (N_30421,N_28860,N_29150);
nor U30422 (N_30422,N_28212,N_27832);
nor U30423 (N_30423,N_28169,N_27569);
nand U30424 (N_30424,N_28191,N_28580);
nor U30425 (N_30425,N_28442,N_29269);
or U30426 (N_30426,N_29821,N_29352);
xnor U30427 (N_30427,N_29188,N_27851);
nand U30428 (N_30428,N_28431,N_28571);
and U30429 (N_30429,N_29976,N_29579);
or U30430 (N_30430,N_29410,N_28998);
nand U30431 (N_30431,N_28388,N_29046);
or U30432 (N_30432,N_28374,N_29224);
xnor U30433 (N_30433,N_28890,N_29604);
nand U30434 (N_30434,N_27727,N_29775);
and U30435 (N_30435,N_29070,N_29720);
nand U30436 (N_30436,N_28480,N_29516);
nor U30437 (N_30437,N_27870,N_29190);
or U30438 (N_30438,N_29119,N_29341);
nand U30439 (N_30439,N_28514,N_28793);
xnor U30440 (N_30440,N_29176,N_29786);
or U30441 (N_30441,N_27692,N_28470);
and U30442 (N_30442,N_29077,N_27904);
and U30443 (N_30443,N_29165,N_29570);
nand U30444 (N_30444,N_29302,N_29357);
nor U30445 (N_30445,N_29855,N_28837);
or U30446 (N_30446,N_28319,N_29222);
nor U30447 (N_30447,N_28264,N_29399);
nand U30448 (N_30448,N_28686,N_29406);
nand U30449 (N_30449,N_28800,N_28008);
nor U30450 (N_30450,N_28870,N_28006);
xor U30451 (N_30451,N_27924,N_27628);
nor U30452 (N_30452,N_29885,N_28541);
and U30453 (N_30453,N_28235,N_29485);
xor U30454 (N_30454,N_28577,N_27843);
or U30455 (N_30455,N_27842,N_27935);
or U30456 (N_30456,N_27770,N_28464);
or U30457 (N_30457,N_29274,N_27588);
nand U30458 (N_30458,N_27539,N_29340);
nand U30459 (N_30459,N_28803,N_27869);
nor U30460 (N_30460,N_28558,N_29970);
xor U30461 (N_30461,N_27616,N_27872);
nor U30462 (N_30462,N_29247,N_29080);
or U30463 (N_30463,N_29230,N_29041);
nor U30464 (N_30464,N_27955,N_27880);
xor U30465 (N_30465,N_29339,N_29868);
nand U30466 (N_30466,N_29355,N_28721);
nand U30467 (N_30467,N_27945,N_27940);
and U30468 (N_30468,N_29445,N_28720);
or U30469 (N_30469,N_27771,N_27954);
or U30470 (N_30470,N_28538,N_28285);
or U30471 (N_30471,N_27921,N_28570);
nand U30472 (N_30472,N_29225,N_28766);
nor U30473 (N_30473,N_28994,N_28121);
xnor U30474 (N_30474,N_27568,N_28723);
nand U30475 (N_30475,N_28024,N_28518);
or U30476 (N_30476,N_28194,N_29283);
or U30477 (N_30477,N_27636,N_29795);
or U30478 (N_30478,N_28305,N_28375);
nor U30479 (N_30479,N_28419,N_27876);
and U30480 (N_30480,N_27905,N_27815);
nand U30481 (N_30481,N_29589,N_29722);
and U30482 (N_30482,N_29361,N_29693);
xor U30483 (N_30483,N_29422,N_28096);
or U30484 (N_30484,N_28634,N_27669);
and U30485 (N_30485,N_29084,N_29684);
xnor U30486 (N_30486,N_28901,N_29298);
nand U30487 (N_30487,N_29085,N_27610);
nor U30488 (N_30488,N_28328,N_28227);
xor U30489 (N_30489,N_29750,N_29643);
nand U30490 (N_30490,N_27633,N_29260);
nor U30491 (N_30491,N_29687,N_28202);
and U30492 (N_30492,N_27660,N_29549);
nor U30493 (N_30493,N_27860,N_28977);
or U30494 (N_30494,N_29022,N_27751);
or U30495 (N_30495,N_27874,N_28728);
nor U30496 (N_30496,N_29632,N_28761);
or U30497 (N_30497,N_29348,N_29980);
or U30498 (N_30498,N_29508,N_29184);
and U30499 (N_30499,N_27555,N_27579);
nor U30500 (N_30500,N_27714,N_27848);
nand U30501 (N_30501,N_29900,N_27645);
nand U30502 (N_30502,N_27795,N_29667);
nor U30503 (N_30503,N_29807,N_28601);
or U30504 (N_30504,N_28397,N_29144);
xor U30505 (N_30505,N_27540,N_29453);
nor U30506 (N_30506,N_27854,N_27896);
or U30507 (N_30507,N_29194,N_29183);
nand U30508 (N_30508,N_29743,N_28505);
nor U30509 (N_30509,N_28693,N_29434);
and U30510 (N_30510,N_28623,N_29469);
and U30511 (N_30511,N_28660,N_28312);
or U30512 (N_30512,N_28632,N_28916);
nor U30513 (N_30513,N_29280,N_28543);
or U30514 (N_30514,N_27504,N_29800);
or U30515 (N_30515,N_29458,N_28646);
xor U30516 (N_30516,N_28889,N_28166);
nand U30517 (N_30517,N_28503,N_29163);
nand U30518 (N_30518,N_28361,N_28719);
or U30519 (N_30519,N_28394,N_28355);
xor U30520 (N_30520,N_28434,N_28705);
xnor U30521 (N_30521,N_29402,N_27722);
nor U30522 (N_30522,N_27981,N_28527);
and U30523 (N_30523,N_29191,N_27517);
xor U30524 (N_30524,N_28628,N_29467);
and U30525 (N_30525,N_29028,N_28773);
nor U30526 (N_30526,N_29186,N_28461);
nor U30527 (N_30527,N_29801,N_29983);
or U30528 (N_30528,N_28536,N_29300);
or U30529 (N_30529,N_27853,N_29865);
xor U30530 (N_30530,N_28509,N_29411);
nand U30531 (N_30531,N_28876,N_28604);
xnor U30532 (N_30532,N_28673,N_29861);
nand U30533 (N_30533,N_28512,N_27611);
xor U30534 (N_30534,N_29332,N_28130);
nor U30535 (N_30535,N_28425,N_28983);
and U30536 (N_30536,N_29945,N_29564);
nand U30537 (N_30537,N_29034,N_28421);
or U30538 (N_30538,N_29823,N_29441);
and U30539 (N_30539,N_29982,N_29587);
and U30540 (N_30540,N_29366,N_27705);
nand U30541 (N_30541,N_27897,N_29480);
nor U30542 (N_30542,N_27759,N_29994);
and U30543 (N_30543,N_28294,N_28999);
and U30544 (N_30544,N_28684,N_29902);
or U30545 (N_30545,N_27942,N_29594);
and U30546 (N_30546,N_28855,N_29562);
or U30547 (N_30547,N_27953,N_29791);
or U30548 (N_30548,N_29153,N_28717);
nor U30549 (N_30549,N_27650,N_27855);
nor U30550 (N_30550,N_27970,N_28398);
nor U30551 (N_30551,N_27952,N_27883);
and U30552 (N_30552,N_29245,N_28984);
nand U30553 (N_30553,N_27776,N_28094);
xor U30554 (N_30554,N_29652,N_29220);
and U30555 (N_30555,N_27677,N_28759);
nand U30556 (N_30556,N_29659,N_28718);
and U30557 (N_30557,N_29346,N_29129);
nor U30558 (N_30558,N_28790,N_27746);
nand U30559 (N_30559,N_28225,N_29524);
nor U30560 (N_30560,N_29305,N_29362);
nand U30561 (N_30561,N_29939,N_28864);
nor U30562 (N_30562,N_28508,N_28528);
or U30563 (N_30563,N_28698,N_29903);
or U30564 (N_30564,N_28967,N_28334);
nand U30565 (N_30565,N_29114,N_28842);
nor U30566 (N_30566,N_29778,N_27695);
xnor U30567 (N_30567,N_29645,N_27562);
xnor U30568 (N_30568,N_28297,N_28380);
nor U30569 (N_30569,N_28829,N_28872);
nand U30570 (N_30570,N_29322,N_29733);
xor U30571 (N_30571,N_29262,N_29688);
nand U30572 (N_30572,N_29824,N_28122);
and U30573 (N_30573,N_28633,N_27578);
or U30574 (N_30574,N_29216,N_29037);
or U30575 (N_30575,N_29910,N_28306);
nor U30576 (N_30576,N_28399,N_28458);
or U30577 (N_30577,N_28451,N_28727);
nand U30578 (N_30578,N_28404,N_29835);
and U30579 (N_30579,N_27922,N_28265);
or U30580 (N_30580,N_29479,N_27741);
nand U30581 (N_30581,N_29013,N_27823);
nand U30582 (N_30582,N_29932,N_29242);
nor U30583 (N_30583,N_28567,N_29271);
or U30584 (N_30584,N_27973,N_28147);
nand U30585 (N_30585,N_28042,N_29633);
or U30586 (N_30586,N_28330,N_28928);
nand U30587 (N_30587,N_29719,N_27934);
nand U30588 (N_30588,N_28966,N_27552);
nor U30589 (N_30589,N_29701,N_28969);
nand U30590 (N_30590,N_27779,N_27890);
xor U30591 (N_30591,N_29815,N_29456);
nand U30592 (N_30592,N_28248,N_29840);
xor U30593 (N_30593,N_28282,N_29658);
xor U30594 (N_30594,N_28965,N_28098);
nor U30595 (N_30595,N_28219,N_28794);
and U30596 (N_30596,N_28620,N_29487);
nor U30597 (N_30597,N_29727,N_28254);
nand U30598 (N_30598,N_29639,N_27693);
xor U30599 (N_30599,N_28186,N_28791);
nand U30600 (N_30600,N_28102,N_29056);
nor U30601 (N_30601,N_27686,N_29081);
nor U30602 (N_30602,N_27756,N_29409);
nor U30603 (N_30603,N_29038,N_28535);
and U30604 (N_30604,N_28483,N_27782);
and U30605 (N_30605,N_27808,N_28915);
nor U30606 (N_30606,N_27593,N_28409);
or U30607 (N_30607,N_29454,N_28696);
nor U30608 (N_30608,N_29888,N_28802);
or U30609 (N_30609,N_28765,N_29451);
nand U30610 (N_30610,N_27572,N_27989);
nor U30611 (N_30611,N_29083,N_29540);
xor U30612 (N_30612,N_28462,N_27735);
or U30613 (N_30613,N_28056,N_27979);
or U30614 (N_30614,N_29486,N_28581);
or U30615 (N_30615,N_28887,N_28356);
nor U30616 (N_30616,N_28080,N_29179);
nand U30617 (N_30617,N_29133,N_28704);
and U30618 (N_30618,N_29353,N_29047);
and U30619 (N_30619,N_29811,N_28607);
or U30620 (N_30620,N_29143,N_28384);
or U30621 (N_30621,N_28321,N_28824);
nand U30622 (N_30622,N_29635,N_28061);
nand U30623 (N_30623,N_29071,N_28011);
and U30624 (N_30624,N_28838,N_27697);
and U30625 (N_30625,N_28767,N_28062);
or U30626 (N_30626,N_28475,N_27606);
nor U30627 (N_30627,N_28129,N_29806);
xor U30628 (N_30628,N_29039,N_29699);
nand U30629 (N_30629,N_28683,N_29878);
and U30630 (N_30630,N_28030,N_28561);
nand U30631 (N_30631,N_28258,N_29814);
or U30632 (N_30632,N_28001,N_29288);
nand U30633 (N_30633,N_29158,N_27769);
nor U30634 (N_30634,N_28830,N_29736);
nand U30635 (N_30635,N_27958,N_28293);
nor U30636 (N_30636,N_28929,N_29961);
nand U30637 (N_30637,N_29591,N_28598);
nor U30638 (N_30638,N_29975,N_27533);
or U30639 (N_30639,N_29418,N_29810);
nand U30640 (N_30640,N_28382,N_28107);
and U30641 (N_30641,N_27968,N_29716);
nand U30642 (N_30642,N_28273,N_29035);
and U30643 (N_30643,N_27586,N_28659);
nor U30644 (N_30644,N_29605,N_29236);
or U30645 (N_30645,N_28602,N_28788);
xor U30646 (N_30646,N_28655,N_28831);
or U30647 (N_30647,N_27515,N_29877);
or U30648 (N_30648,N_27923,N_28441);
or U30649 (N_30649,N_27513,N_29492);
and U30650 (N_30650,N_27639,N_27688);
and U30651 (N_30651,N_28534,N_29614);
and U30652 (N_30652,N_28308,N_29000);
or U30653 (N_30653,N_28301,N_27700);
and U30654 (N_30654,N_29704,N_29440);
nor U30655 (N_30655,N_27612,N_29534);
and U30656 (N_30656,N_28307,N_29555);
or U30657 (N_30657,N_29916,N_28575);
nor U30658 (N_30658,N_29813,N_27543);
and U30659 (N_30659,N_28973,N_28978);
and U30660 (N_30660,N_27694,N_28128);
and U30661 (N_30661,N_28174,N_28671);
xor U30662 (N_30662,N_29067,N_29725);
nand U30663 (N_30663,N_28554,N_29571);
or U30664 (N_30664,N_27839,N_27930);
and U30665 (N_30665,N_28752,N_29024);
nand U30666 (N_30666,N_28863,N_28263);
nor U30667 (N_30667,N_29627,N_28127);
nor U30668 (N_30668,N_28941,N_29170);
nand U30669 (N_30669,N_27920,N_29328);
and U30670 (N_30670,N_29776,N_28084);
xor U30671 (N_30671,N_28685,N_27520);
or U30672 (N_30672,N_29010,N_27747);
nand U30673 (N_30673,N_29891,N_29177);
nor U30674 (N_30674,N_27946,N_27867);
nand U30675 (N_30675,N_29155,N_28501);
nand U30676 (N_30676,N_28900,N_29847);
nor U30677 (N_30677,N_28251,N_28638);
nand U30678 (N_30678,N_29896,N_27728);
nand U30679 (N_30679,N_29196,N_28533);
nor U30680 (N_30680,N_27919,N_28161);
and U30681 (N_30681,N_29256,N_27538);
nor U30682 (N_30682,N_29189,N_29763);
or U30683 (N_30683,N_28737,N_27877);
nand U30684 (N_30684,N_29239,N_29583);
nand U30685 (N_30685,N_27809,N_29208);
nor U30686 (N_30686,N_28493,N_28242);
nand U30687 (N_30687,N_28531,N_29435);
nand U30688 (N_30688,N_27640,N_29703);
nor U30689 (N_30689,N_28268,N_29062);
nand U30690 (N_30690,N_29029,N_29582);
nand U30691 (N_30691,N_28677,N_27899);
nor U30692 (N_30692,N_28675,N_29326);
nor U30693 (N_30693,N_27763,N_29334);
nor U30694 (N_30694,N_29552,N_28123);
or U30695 (N_30695,N_29131,N_29212);
xnor U30696 (N_30696,N_28546,N_29128);
or U30697 (N_30697,N_28032,N_28525);
nor U30698 (N_30698,N_28156,N_29648);
and U30699 (N_30699,N_29377,N_28392);
or U30700 (N_30700,N_29770,N_29001);
xnor U30701 (N_30701,N_29235,N_27662);
or U30702 (N_30702,N_29834,N_29761);
nor U30703 (N_30703,N_27665,N_28424);
and U30704 (N_30704,N_29784,N_29363);
nor U30705 (N_30705,N_28369,N_28167);
nand U30706 (N_30706,N_27772,N_28482);
nor U30707 (N_30707,N_29829,N_28560);
nand U30708 (N_30708,N_28200,N_27738);
and U30709 (N_30709,N_28680,N_28302);
nor U30710 (N_30710,N_28207,N_27577);
or U30711 (N_30711,N_27797,N_28805);
and U30712 (N_30712,N_29575,N_28740);
nand U30713 (N_30713,N_28681,N_27901);
and U30714 (N_30714,N_28055,N_29749);
nor U30715 (N_30715,N_29592,N_29651);
nor U30716 (N_30716,N_29681,N_28706);
nand U30717 (N_30717,N_29057,N_28446);
and U30718 (N_30718,N_27982,N_29138);
nor U30719 (N_30719,N_29593,N_27865);
and U30720 (N_30720,N_27681,N_29691);
and U30721 (N_30721,N_27814,N_27541);
nor U30722 (N_30722,N_28729,N_29318);
nand U30723 (N_30723,N_29379,N_29463);
nor U30724 (N_30724,N_29042,N_29751);
nor U30725 (N_30725,N_27721,N_28134);
nand U30726 (N_30726,N_28143,N_28832);
and U30727 (N_30727,N_28653,N_29936);
nand U30728 (N_30728,N_27850,N_29059);
or U30729 (N_30729,N_27740,N_28565);
or U30730 (N_30730,N_29468,N_27861);
nor U30731 (N_30731,N_29963,N_29876);
nand U30732 (N_30732,N_28286,N_28018);
and U30733 (N_30733,N_27547,N_29901);
nor U30734 (N_30734,N_28875,N_28932);
nor U30735 (N_30735,N_29551,N_27656);
nand U30736 (N_30736,N_29372,N_28579);
nor U30737 (N_30737,N_27651,N_27984);
nor U30738 (N_30738,N_29182,N_28768);
nand U30739 (N_30739,N_27674,N_29380);
xnor U30740 (N_30740,N_28417,N_28357);
nor U30741 (N_30741,N_27501,N_28278);
or U30742 (N_30742,N_27838,N_27725);
nor U30743 (N_30743,N_28866,N_28364);
nor U30744 (N_30744,N_29566,N_27620);
nor U30745 (N_30745,N_29359,N_29735);
nor U30746 (N_30746,N_28833,N_28255);
or U30747 (N_30747,N_29036,N_29997);
and U30748 (N_30748,N_28665,N_29586);
nor U30749 (N_30749,N_29839,N_27766);
and U30750 (N_30750,N_29950,N_28658);
xnor U30751 (N_30751,N_27884,N_28931);
nand U30752 (N_30752,N_28230,N_29887);
or U30753 (N_30753,N_27603,N_27528);
xnor U30754 (N_30754,N_29689,N_29637);
nand U30755 (N_30755,N_29360,N_29797);
nor U30756 (N_30756,N_28354,N_28160);
nand U30757 (N_30757,N_29060,N_29598);
or U30758 (N_30758,N_29045,N_29495);
nand U30759 (N_30759,N_28466,N_28333);
or U30760 (N_30760,N_27915,N_28345);
and U30761 (N_30761,N_27561,N_27991);
and U30762 (N_30762,N_29095,N_28237);
nor U30763 (N_30763,N_29112,N_28610);
xor U30764 (N_30764,N_29925,N_29915);
nand U30765 (N_30765,N_28436,N_27773);
or U30766 (N_30766,N_29251,N_29126);
or U30767 (N_30767,N_27710,N_29146);
nand U30768 (N_30768,N_29068,N_29781);
nand U30769 (N_30769,N_29099,N_29668);
xnor U30770 (N_30770,N_29217,N_27712);
and U30771 (N_30771,N_29444,N_29031);
nand U30772 (N_30772,N_28668,N_29670);
or U30773 (N_30773,N_27599,N_29981);
nor U30774 (N_30774,N_28555,N_29602);
or U30775 (N_30775,N_29710,N_28519);
nand U30776 (N_30776,N_29618,N_29240);
nor U30777 (N_30777,N_29989,N_28676);
and U30778 (N_30778,N_27742,N_28540);
nand U30779 (N_30779,N_29018,N_29023);
nand U30780 (N_30780,N_29580,N_29169);
and U30781 (N_30781,N_28769,N_29051);
and U30782 (N_30782,N_29481,N_29886);
xor U30783 (N_30783,N_28981,N_28946);
nor U30784 (N_30784,N_29122,N_28747);
xnor U30785 (N_30785,N_27962,N_28521);
and U30786 (N_30786,N_27560,N_28196);
and U30787 (N_30787,N_28689,N_27708);
or U30788 (N_30788,N_28454,N_27654);
nor U30789 (N_30789,N_27542,N_28947);
xnor U30790 (N_30790,N_29794,N_29805);
or U30791 (N_30791,N_28220,N_28106);
or U30792 (N_30792,N_29871,N_27966);
nor U30793 (N_30793,N_29543,N_29873);
nor U30794 (N_30794,N_29923,N_29996);
nand U30795 (N_30795,N_28992,N_27892);
nor U30796 (N_30796,N_29883,N_28343);
nand U30797 (N_30797,N_28112,N_28934);
nor U30798 (N_30798,N_28103,N_28428);
nand U30799 (N_30799,N_28739,N_28060);
and U30800 (N_30800,N_27706,N_29966);
and U30801 (N_30801,N_29102,N_28840);
nor U30802 (N_30802,N_28037,N_29754);
or U30803 (N_30803,N_28157,N_29002);
or U30804 (N_30804,N_28782,N_29926);
and U30805 (N_30805,N_27778,N_28439);
or U30806 (N_30806,N_28574,N_29650);
and U30807 (N_30807,N_28316,N_29286);
nand U30808 (N_30808,N_29275,N_28303);
nand U30809 (N_30809,N_29611,N_27580);
nand U30810 (N_30810,N_28007,N_28930);
or U30811 (N_30811,N_29671,N_27576);
nand U30812 (N_30812,N_28151,N_29857);
and U30813 (N_30813,N_28921,N_29497);
nor U30814 (N_30814,N_29506,N_29912);
xnor U30815 (N_30815,N_28500,N_29382);
or U30816 (N_30816,N_29862,N_27893);
and U30817 (N_30817,N_29226,N_29476);
nor U30818 (N_30818,N_28725,N_29296);
nor U30819 (N_30819,N_28017,N_28626);
nand U30820 (N_30820,N_28047,N_29792);
and U30821 (N_30821,N_28637,N_29221);
nor U30822 (N_30822,N_29785,N_27529);
or U30823 (N_30823,N_28688,N_28014);
and U30824 (N_30824,N_28882,N_29771);
and U30825 (N_30825,N_28262,N_28823);
and U30826 (N_30826,N_29550,N_28481);
nand U30827 (N_30827,N_29802,N_29197);
and U30828 (N_30828,N_28478,N_28584);
or U30829 (N_30829,N_28315,N_29079);
nand U30830 (N_30830,N_29528,N_29325);
nor U30831 (N_30831,N_27535,N_28924);
and U30832 (N_30832,N_28426,N_28596);
nor U30833 (N_30833,N_28035,N_29777);
or U30834 (N_30834,N_29712,N_28898);
and U30835 (N_30835,N_28070,N_29747);
or U30836 (N_30836,N_29285,N_28568);
and U30837 (N_30837,N_28089,N_27939);
and U30838 (N_30838,N_29622,N_29804);
nor U30839 (N_30839,N_27729,N_28420);
nand U30840 (N_30840,N_28231,N_29092);
nor U30841 (N_30841,N_27604,N_29223);
and U30842 (N_30842,N_29185,N_28043);
or U30843 (N_30843,N_29436,N_28430);
and U30844 (N_30844,N_29115,N_27951);
or U30845 (N_30845,N_28636,N_29756);
nor U30846 (N_30846,N_29867,N_28370);
nor U30847 (N_30847,N_29853,N_28714);
or U30848 (N_30848,N_29228,N_29567);
nand U30849 (N_30849,N_29757,N_28582);
nor U30850 (N_30850,N_29374,N_29818);
xor U30851 (N_30851,N_29427,N_29276);
and U30852 (N_30852,N_28524,N_29003);
or U30853 (N_30853,N_27790,N_29890);
nand U30854 (N_30854,N_29253,N_29768);
nand U30855 (N_30855,N_28522,N_29457);
or U30856 (N_30856,N_28741,N_28566);
or U30857 (N_30857,N_27726,N_28695);
or U30858 (N_30858,N_28124,N_28588);
xor U30859 (N_30859,N_27813,N_29726);
or U30860 (N_30860,N_29803,N_27600);
and U30861 (N_30861,N_29116,N_27679);
and U30862 (N_30862,N_28682,N_29962);
or U30863 (N_30863,N_27783,N_27715);
and U30864 (N_30864,N_29093,N_27882);
nor U30865 (N_30865,N_29946,N_27752);
or U30866 (N_30866,N_27661,N_29588);
or U30867 (N_30867,N_29277,N_27788);
nand U30868 (N_30868,N_29744,N_27737);
nor U30869 (N_30869,N_27626,N_29301);
or U30870 (N_30870,N_29880,N_28796);
nand U30871 (N_30871,N_28105,N_28892);
xor U30872 (N_30872,N_28817,N_28827);
xnor U30873 (N_30873,N_29309,N_29677);
nand U30874 (N_30874,N_29259,N_29826);
xnor U30875 (N_30875,N_29819,N_29336);
or U30876 (N_30876,N_28190,N_28004);
nand U30877 (N_30877,N_28885,N_27581);
nand U30878 (N_30878,N_28295,N_28068);
nor U30879 (N_30879,N_28799,N_29897);
nand U30880 (N_30880,N_28175,N_29581);
xnor U30881 (N_30881,N_29640,N_28433);
or U30882 (N_30882,N_29314,N_29942);
nor U30883 (N_30883,N_29557,N_29397);
nor U30884 (N_30884,N_29073,N_27996);
nor U30885 (N_30885,N_29132,N_29827);
xor U30886 (N_30886,N_27959,N_28743);
or U30887 (N_30887,N_29634,N_28117);
and U30888 (N_30888,N_29473,N_29086);
nand U30889 (N_30889,N_28114,N_29210);
and U30890 (N_30890,N_29965,N_28337);
nand U30891 (N_30891,N_28621,N_29851);
and U30892 (N_30892,N_29992,N_27570);
nor U30893 (N_30893,N_29011,N_27824);
or U30894 (N_30894,N_28848,N_27701);
and U30895 (N_30895,N_27985,N_27689);
nor U30896 (N_30896,N_29203,N_29395);
xor U30897 (N_30897,N_29520,N_28445);
or U30898 (N_30898,N_28547,N_28853);
and U30899 (N_30899,N_29121,N_29295);
or U30900 (N_30900,N_28701,N_29631);
nand U30901 (N_30901,N_27685,N_27898);
and U30902 (N_30902,N_28650,N_29523);
xor U30903 (N_30903,N_28962,N_29844);
nand U30904 (N_30904,N_27888,N_28327);
nand U30905 (N_30905,N_27602,N_29330);
nand U30906 (N_30906,N_27812,N_28353);
nand U30907 (N_30907,N_28991,N_28082);
or U30908 (N_30908,N_28738,N_28279);
nor U30909 (N_30909,N_29323,N_28086);
nand U30910 (N_30910,N_28985,N_28232);
xor U30911 (N_30911,N_28844,N_27605);
and U30912 (N_30912,N_29090,N_28489);
and U30913 (N_30913,N_29908,N_27632);
or U30914 (N_30914,N_28925,N_28670);
or U30915 (N_30915,N_27592,N_28780);
xor U30916 (N_30916,N_29569,N_27948);
and U30917 (N_30917,N_29489,N_29484);
nand U30918 (N_30918,N_28111,N_28427);
or U30919 (N_30919,N_28299,N_28021);
and U30920 (N_30920,N_28777,N_28849);
and U30921 (N_30921,N_29008,N_28746);
nand U30922 (N_30922,N_29266,N_28710);
xor U30923 (N_30923,N_29100,N_28943);
nor U30924 (N_30924,N_29421,N_28290);
and U30925 (N_30925,N_29052,N_27972);
nand U30926 (N_30926,N_29390,N_28188);
xor U30927 (N_30927,N_29759,N_28269);
or U30928 (N_30928,N_29530,N_29135);
or U30929 (N_30929,N_29825,N_28530);
nor U30930 (N_30930,N_28256,N_28054);
nand U30931 (N_30931,N_28756,N_29033);
and U30932 (N_30932,N_28949,N_28249);
nand U30933 (N_30933,N_28005,N_28764);
nand U30934 (N_30934,N_29773,N_29218);
nor U30935 (N_30935,N_28651,N_29007);
and U30936 (N_30936,N_29333,N_29307);
and U30937 (N_30937,N_28003,N_29254);
or U30938 (N_30938,N_28556,N_29075);
or U30939 (N_30939,N_27796,N_27820);
or U30940 (N_30940,N_28841,N_29313);
nor U30941 (N_30941,N_29617,N_29494);
nor U30942 (N_30942,N_28221,N_29860);
and U30943 (N_30943,N_28724,N_27863);
and U30944 (N_30944,N_29595,N_27736);
nor U30945 (N_30945,N_28331,N_29774);
and U30946 (N_30946,N_28748,N_29600);
xnor U30947 (N_30947,N_28763,N_27519);
and U30948 (N_30948,N_29721,N_27785);
nor U30949 (N_30949,N_29660,N_29160);
nand U30950 (N_30950,N_27615,N_28444);
nor U30951 (N_30951,N_29496,N_29892);
nand U30952 (N_30952,N_28073,N_28359);
nor U30953 (N_30953,N_28313,N_27871);
and U30954 (N_30954,N_28423,N_27553);
nor U30955 (N_30955,N_29344,N_27986);
and U30956 (N_30956,N_29294,N_28144);
and U30957 (N_30957,N_27825,N_28990);
and U30958 (N_30958,N_29430,N_28700);
or U30959 (N_30959,N_29292,N_28709);
nand U30960 (N_30960,N_28045,N_28591);
or U30961 (N_30961,N_28993,N_29017);
or U30962 (N_30962,N_28862,N_29443);
nor U30963 (N_30963,N_27609,N_27811);
or U30964 (N_30964,N_28776,N_29672);
xnor U30965 (N_30965,N_28266,N_27830);
nand U30966 (N_30966,N_28529,N_28813);
nor U30967 (N_30967,N_29542,N_27597);
and U30968 (N_30968,N_27613,N_28654);
and U30969 (N_30969,N_29164,N_29408);
nand U30970 (N_30970,N_29512,N_27523);
and U30971 (N_30971,N_27914,N_28792);
or U30972 (N_30972,N_27585,N_27840);
and U30973 (N_30973,N_28040,N_29683);
nor U30974 (N_30974,N_27672,N_29091);
and U30975 (N_30975,N_29446,N_27866);
or U30976 (N_30976,N_29331,N_29626);
xor U30977 (N_30977,N_29724,N_29291);
nand U30978 (N_30978,N_29120,N_29674);
nand U30979 (N_30979,N_27927,N_27817);
xnor U30980 (N_30980,N_28736,N_28821);
nand U30981 (N_30981,N_27507,N_29664);
and U30982 (N_30982,N_28499,N_28214);
or U30983 (N_30983,N_28798,N_28641);
nand U30984 (N_30984,N_28879,N_29148);
and U30985 (N_30985,N_27827,N_29988);
or U30986 (N_30986,N_29737,N_29616);
nor U30987 (N_30987,N_29175,N_28447);
and U30988 (N_30988,N_29050,N_29103);
and U30989 (N_30989,N_28542,N_28038);
and U30990 (N_30990,N_27510,N_29629);
or U30991 (N_30991,N_27967,N_27646);
or U30992 (N_30992,N_28526,N_27949);
nand U30993 (N_30993,N_28942,N_27976);
or U30994 (N_30994,N_28346,N_28635);
or U30995 (N_30995,N_28390,N_29261);
xor U30996 (N_30996,N_29609,N_27836);
nand U30997 (N_30997,N_28492,N_27587);
nor U30998 (N_30998,N_29198,N_28667);
and U30999 (N_30999,N_27644,N_29460);
and U31000 (N_31000,N_27630,N_28119);
and U31001 (N_31001,N_29424,N_28835);
nand U31002 (N_31002,N_29553,N_27566);
nand U31003 (N_31003,N_27641,N_29911);
nor U31004 (N_31004,N_29021,N_29475);
nor U31005 (N_31005,N_28730,N_29371);
or U31006 (N_31006,N_29338,N_29205);
nor U31007 (N_31007,N_27849,N_27886);
nand U31008 (N_31008,N_28615,N_29836);
or U31009 (N_31009,N_27717,N_29124);
and U31010 (N_31010,N_29368,N_28443);
nor U31011 (N_31011,N_27558,N_29563);
nand U31012 (N_31012,N_28198,N_29384);
and U31013 (N_31013,N_27719,N_28253);
or U31014 (N_31014,N_28274,N_28463);
nor U31015 (N_31015,N_29700,N_27608);
nor U31016 (N_31016,N_28416,N_27595);
nand U31017 (N_31017,N_28090,N_29854);
or U31018 (N_31018,N_29268,N_29252);
and U31019 (N_31019,N_29097,N_28583);
and U31020 (N_31020,N_28883,N_28511);
or U31021 (N_31021,N_28974,N_28881);
nor U31022 (N_31022,N_28206,N_29809);
nand U31023 (N_31023,N_28484,N_29365);
nor U31024 (N_31024,N_29746,N_28363);
and U31025 (N_31025,N_29383,N_27810);
nand U31026 (N_31026,N_29830,N_28989);
nand U31027 (N_31027,N_27690,N_29978);
and U31028 (N_31028,N_29279,N_29415);
nand U31029 (N_31029,N_27821,N_29393);
xor U31030 (N_31030,N_28595,N_29788);
and U31031 (N_31031,N_27508,N_27999);
or U31032 (N_31032,N_27784,N_27995);
and U31033 (N_31033,N_29858,N_28339);
nand U31034 (N_31034,N_28516,N_28211);
and U31035 (N_31035,N_27768,N_28429);
and U31036 (N_31036,N_29822,N_27988);
and U31037 (N_31037,N_28415,N_28801);
or U31038 (N_31038,N_28858,N_27667);
or U31039 (N_31039,N_29845,N_28557);
xnor U31040 (N_31040,N_27739,N_28888);
nor U31041 (N_31041,N_28713,N_28624);
or U31042 (N_31042,N_28183,N_27634);
or U31043 (N_31043,N_28177,N_29192);
nand U31044 (N_31044,N_28939,N_28087);
nor U31045 (N_31045,N_28455,N_28948);
and U31046 (N_31046,N_28957,N_28223);
or U31047 (N_31047,N_28072,N_28058);
or U31048 (N_31048,N_28403,N_28912);
nand U31049 (N_31049,N_29657,N_29231);
nor U31050 (N_31050,N_29762,N_28016);
nand U31051 (N_31051,N_28662,N_29852);
nor U31052 (N_31052,N_28648,N_27594);
and U31053 (N_31053,N_29449,N_29396);
nor U31054 (N_31054,N_29999,N_29403);
nor U31055 (N_31055,N_29538,N_29838);
nand U31056 (N_31056,N_29764,N_28772);
nor U31057 (N_31057,N_27683,N_28182);
nor U31058 (N_31058,N_29909,N_28323);
or U31059 (N_31059,N_29137,N_28812);
xor U31060 (N_31060,N_28245,N_28097);
nor U31061 (N_31061,N_28674,N_28775);
and U31062 (N_31062,N_28044,N_28241);
nand U31063 (N_31063,N_28407,N_28902);
nand U31064 (N_31064,N_28910,N_29234);
nand U31065 (N_31065,N_28578,N_27878);
nand U31066 (N_31066,N_29849,N_28573);
nor U31067 (N_31067,N_28490,N_29584);
or U31068 (N_31068,N_28309,N_29213);
or U31069 (N_31069,N_29870,N_28387);
and U31070 (N_31070,N_29798,N_27891);
or U31071 (N_31071,N_29728,N_29351);
xor U31072 (N_31072,N_29646,N_28917);
nand U31073 (N_31073,N_29354,N_28734);
and U31074 (N_31074,N_28020,N_28839);
nand U31075 (N_31075,N_29381,N_28631);
or U31076 (N_31076,N_29420,N_28485);
nand U31077 (N_31077,N_28270,N_29214);
nand U31078 (N_31078,N_28545,N_29320);
or U31079 (N_31079,N_27575,N_29061);
xor U31080 (N_31080,N_28612,N_29577);
and U31081 (N_31081,N_29229,N_27894);
nor U31082 (N_31082,N_28856,N_27960);
nor U31083 (N_31083,N_28304,N_28927);
nand U31084 (N_31084,N_28488,N_27583);
and U31085 (N_31085,N_29405,N_28351);
nand U31086 (N_31086,N_27527,N_29675);
nand U31087 (N_31087,N_29149,N_28222);
nand U31088 (N_31088,N_29894,N_29972);
and U31089 (N_31089,N_29356,N_27895);
nand U31090 (N_31090,N_27950,N_29559);
and U31091 (N_31091,N_28815,N_29154);
nand U31092 (N_31092,N_28210,N_28807);
and U31093 (N_31093,N_29613,N_29156);
nor U31094 (N_31094,N_28342,N_28605);
xor U31095 (N_31095,N_27764,N_27917);
or U31096 (N_31096,N_27845,N_28960);
nor U31097 (N_31097,N_29178,N_27624);
and U31098 (N_31098,N_29765,N_27526);
nor U31099 (N_31099,N_28731,N_29026);
nor U31100 (N_31100,N_28408,N_29739);
and U31101 (N_31101,N_29590,N_27625);
nand U31102 (N_31102,N_29679,N_29958);
or U31103 (N_31103,N_28362,N_29049);
or U31104 (N_31104,N_28271,N_29578);
and U31105 (N_31105,N_29930,N_28140);
and U31106 (N_31106,N_29278,N_28661);
or U31107 (N_31107,N_29303,N_29206);
or U31108 (N_31108,N_28532,N_29623);
nand U31109 (N_31109,N_27621,N_27531);
nand U31110 (N_31110,N_28298,N_29098);
and U31111 (N_31111,N_27678,N_29502);
or U31112 (N_31112,N_28523,N_28052);
nor U31113 (N_31113,N_29123,N_28158);
nor U31114 (N_31114,N_29558,N_29927);
nand U31115 (N_31115,N_28059,N_29918);
or U31116 (N_31116,N_28335,N_29342);
or U31117 (N_31117,N_29364,N_27910);
and U31118 (N_31118,N_28371,N_28252);
xor U31119 (N_31119,N_28320,N_28240);
xor U31120 (N_31120,N_28496,N_28619);
nor U31121 (N_31121,N_28760,N_29638);
nand U31122 (N_31122,N_28472,N_29044);
or U31123 (N_31123,N_28349,N_27623);
nor U31124 (N_31124,N_28344,N_28115);
and U31125 (N_31125,N_28153,N_29110);
or U31126 (N_31126,N_28317,N_27852);
nor U31127 (N_31127,N_29391,N_29250);
xor U31128 (N_31128,N_28975,N_29787);
and U31129 (N_31129,N_29669,N_28643);
or U31130 (N_31130,N_27704,N_28789);
or U31131 (N_31131,N_29656,N_28847);
or U31132 (N_31132,N_27803,N_27965);
and U31133 (N_31133,N_27978,N_27655);
xnor U31134 (N_31134,N_29968,N_28982);
or U31135 (N_31135,N_28199,N_28822);
or U31136 (N_31136,N_29161,N_28707);
and U31137 (N_31137,N_28138,N_28762);
and U31138 (N_31138,N_29101,N_27524);
nor U31139 (N_31139,N_28715,N_28476);
nand U31140 (N_31140,N_27911,N_29032);
and U31141 (N_31141,N_27931,N_29663);
or U31142 (N_31142,N_27564,N_29428);
nand U31143 (N_31143,N_27902,N_29621);
nor U31144 (N_31144,N_29554,N_27652);
nand U31145 (N_31145,N_29995,N_29151);
and U31146 (N_31146,N_29109,N_28487);
nand U31147 (N_31147,N_28609,N_28589);
and U31148 (N_31148,N_28909,N_29267);
or U31149 (N_31149,N_29412,N_29311);
nand U31150 (N_31150,N_28629,N_28970);
and U31151 (N_31151,N_29931,N_29863);
nor U31152 (N_31152,N_27601,N_28953);
xnor U31153 (N_31153,N_28027,N_28336);
and U31154 (N_31154,N_29308,N_27745);
nand U31155 (N_31155,N_27760,N_28868);
nor U31156 (N_31156,N_28576,N_28238);
nor U31157 (N_31157,N_28075,N_27563);
nand U31158 (N_31158,N_29522,N_27505);
nor U31159 (N_31159,N_27794,N_27789);
xor U31160 (N_31160,N_28389,N_28091);
nor U31161 (N_31161,N_28165,N_28154);
nand U31162 (N_31162,N_28101,N_29919);
or U31163 (N_31163,N_28411,N_29960);
nor U31164 (N_31164,N_28284,N_28664);
nand U31165 (N_31165,N_29166,N_29625);
xor U31166 (N_31166,N_28131,N_27598);
nand U31167 (N_31167,N_29913,N_28065);
or U31168 (N_31168,N_29949,N_29941);
and U31169 (N_31169,N_29574,N_28277);
and U31170 (N_31170,N_27591,N_29127);
nor U31171 (N_31171,N_27907,N_28283);
and U31172 (N_31172,N_29914,N_29478);
or U31173 (N_31173,N_28066,N_27909);
and U31174 (N_31174,N_28559,N_29293);
or U31175 (N_31175,N_29974,N_27801);
nand U31176 (N_31176,N_28347,N_29820);
nand U31177 (N_31177,N_28552,N_27589);
nor U31178 (N_31178,N_29831,N_27980);
nor U31179 (N_31179,N_29082,N_28448);
and U31180 (N_31180,N_29483,N_28486);
or U31181 (N_31181,N_28510,N_29243);
nor U31182 (N_31182,N_28692,N_28468);
or U31183 (N_31183,N_29624,N_28246);
nor U31184 (N_31184,N_28811,N_29959);
and U31185 (N_31185,N_29241,N_29561);
and U31186 (N_31186,N_29072,N_28438);
or U31187 (N_31187,N_29796,N_29694);
nor U31188 (N_31188,N_29601,N_29597);
and U31189 (N_31189,N_29063,N_29766);
and U31190 (N_31190,N_28029,N_28260);
nand U31191 (N_31191,N_27720,N_29066);
xor U31192 (N_31192,N_27800,N_28562);
nand U31193 (N_31193,N_27993,N_29159);
and U31194 (N_31194,N_29707,N_28806);
and U31195 (N_31195,N_28996,N_28013);
and U31196 (N_31196,N_28585,N_29297);
xor U31197 (N_31197,N_27618,N_27723);
xnor U31198 (N_31198,N_29882,N_28810);
nor U31199 (N_31199,N_28125,N_28000);
nor U31200 (N_31200,N_29752,N_27680);
and U31201 (N_31201,N_27663,N_29603);
or U31202 (N_31202,N_29730,N_29706);
nand U31203 (N_31203,N_27536,N_29493);
or U31204 (N_31204,N_28672,N_28215);
or U31205 (N_31205,N_28644,N_28292);
or U31206 (N_31206,N_28291,N_29869);
xnor U31207 (N_31207,N_28735,N_29698);
nor U31208 (N_31208,N_27933,N_29030);
xor U31209 (N_31209,N_29507,N_29673);
or U31210 (N_31210,N_28400,N_29118);
nand U31211 (N_31211,N_29004,N_28987);
nand U31212 (N_31212,N_28049,N_29181);
nor U31213 (N_31213,N_28184,N_29527);
nor U31214 (N_31214,N_28678,N_27916);
and U31215 (N_31215,N_28386,N_28139);
nor U31216 (N_31216,N_29649,N_29019);
and U31217 (N_31217,N_28520,N_28275);
nor U31218 (N_31218,N_28699,N_28149);
nand U31219 (N_31219,N_29740,N_28019);
xnor U31220 (N_31220,N_29255,N_28367);
nor U31221 (N_31221,N_28236,N_27792);
and U31222 (N_31222,N_29401,N_28023);
or U31223 (N_31223,N_29500,N_28226);
and U31224 (N_31224,N_28197,N_28869);
xnor U31225 (N_31225,N_29504,N_28630);
nor U31226 (N_31226,N_29832,N_29125);
or U31227 (N_31227,N_27998,N_29337);
nand U31228 (N_31228,N_29450,N_29187);
and U31229 (N_31229,N_29644,N_29180);
xor U31230 (N_31230,N_29678,N_27791);
and U31231 (N_31231,N_27765,N_28150);
nand U31232 (N_31232,N_29760,N_29998);
and U31233 (N_31233,N_27750,N_29204);
nor U31234 (N_31234,N_29407,N_29265);
nand U31235 (N_31235,N_28100,N_28657);
nand U31236 (N_31236,N_28958,N_28396);
nand U31237 (N_31237,N_28599,N_27781);
nand U31238 (N_31238,N_28318,N_27748);
xnor U31239 (N_31239,N_29816,N_29615);
nand U31240 (N_31240,N_29702,N_28218);
and U31241 (N_31241,N_27990,N_27567);
or U31242 (N_31242,N_28597,N_28203);
nor U31243 (N_31243,N_27757,N_28834);
and U31244 (N_31244,N_28053,N_29711);
nor U31245 (N_31245,N_27703,N_29335);
nor U31246 (N_31246,N_27975,N_29264);
and U31247 (N_31247,N_28172,N_27802);
or U31248 (N_31248,N_28324,N_29501);
or U31249 (N_31249,N_29535,N_28376);
nand U31250 (N_31250,N_27702,N_29585);
xor U31251 (N_31251,N_28480,N_29510);
or U31252 (N_31252,N_27644,N_27601);
xnor U31253 (N_31253,N_29839,N_29872);
and U31254 (N_31254,N_27601,N_29966);
nor U31255 (N_31255,N_28456,N_29705);
nand U31256 (N_31256,N_28743,N_27599);
and U31257 (N_31257,N_28545,N_27941);
or U31258 (N_31258,N_28250,N_28785);
xnor U31259 (N_31259,N_29464,N_29702);
xnor U31260 (N_31260,N_28545,N_28533);
or U31261 (N_31261,N_27928,N_28391);
nor U31262 (N_31262,N_28838,N_29920);
and U31263 (N_31263,N_27760,N_27590);
or U31264 (N_31264,N_28673,N_29703);
and U31265 (N_31265,N_29876,N_28287);
xnor U31266 (N_31266,N_28162,N_29652);
nand U31267 (N_31267,N_29418,N_28187);
nand U31268 (N_31268,N_27847,N_29693);
or U31269 (N_31269,N_28911,N_29488);
nand U31270 (N_31270,N_29435,N_28056);
nor U31271 (N_31271,N_29113,N_28849);
nand U31272 (N_31272,N_27515,N_29624);
nand U31273 (N_31273,N_28734,N_28237);
nor U31274 (N_31274,N_29070,N_29141);
and U31275 (N_31275,N_27903,N_28181);
or U31276 (N_31276,N_29250,N_29620);
or U31277 (N_31277,N_28121,N_29155);
xor U31278 (N_31278,N_28887,N_29106);
or U31279 (N_31279,N_29620,N_29000);
nor U31280 (N_31280,N_27893,N_29732);
nor U31281 (N_31281,N_28851,N_28990);
and U31282 (N_31282,N_29558,N_29768);
or U31283 (N_31283,N_27918,N_29536);
nand U31284 (N_31284,N_29808,N_28471);
or U31285 (N_31285,N_27602,N_28112);
nand U31286 (N_31286,N_28691,N_28594);
nor U31287 (N_31287,N_29365,N_29229);
or U31288 (N_31288,N_28811,N_28669);
nor U31289 (N_31289,N_28837,N_28982);
nand U31290 (N_31290,N_29808,N_29497);
or U31291 (N_31291,N_27902,N_29118);
nor U31292 (N_31292,N_28673,N_29994);
and U31293 (N_31293,N_28681,N_29385);
xnor U31294 (N_31294,N_28433,N_29383);
or U31295 (N_31295,N_29521,N_29248);
nor U31296 (N_31296,N_29131,N_29782);
and U31297 (N_31297,N_29573,N_29842);
nand U31298 (N_31298,N_29621,N_29419);
or U31299 (N_31299,N_29200,N_28766);
or U31300 (N_31300,N_28010,N_29412);
nand U31301 (N_31301,N_27907,N_27583);
or U31302 (N_31302,N_28025,N_28925);
and U31303 (N_31303,N_27585,N_28174);
and U31304 (N_31304,N_27882,N_28960);
nand U31305 (N_31305,N_28373,N_28804);
xnor U31306 (N_31306,N_28109,N_29160);
nand U31307 (N_31307,N_27507,N_29984);
nor U31308 (N_31308,N_29977,N_29774);
xor U31309 (N_31309,N_28849,N_29988);
and U31310 (N_31310,N_28092,N_29821);
or U31311 (N_31311,N_28671,N_28834);
or U31312 (N_31312,N_27960,N_28855);
nor U31313 (N_31313,N_29316,N_29466);
nand U31314 (N_31314,N_28208,N_28090);
and U31315 (N_31315,N_28169,N_29381);
and U31316 (N_31316,N_28909,N_28356);
or U31317 (N_31317,N_29103,N_28548);
nor U31318 (N_31318,N_27856,N_28438);
nor U31319 (N_31319,N_29961,N_29287);
nand U31320 (N_31320,N_28679,N_28566);
nand U31321 (N_31321,N_29546,N_28825);
nor U31322 (N_31322,N_28564,N_29717);
nor U31323 (N_31323,N_28061,N_27616);
nor U31324 (N_31324,N_29650,N_27939);
nand U31325 (N_31325,N_29915,N_27684);
and U31326 (N_31326,N_29550,N_28853);
nand U31327 (N_31327,N_27579,N_29567);
nand U31328 (N_31328,N_28418,N_29493);
nor U31329 (N_31329,N_28431,N_28870);
xor U31330 (N_31330,N_29814,N_28817);
nand U31331 (N_31331,N_27937,N_28860);
or U31332 (N_31332,N_28013,N_27758);
nand U31333 (N_31333,N_27913,N_28989);
xor U31334 (N_31334,N_27604,N_27626);
nand U31335 (N_31335,N_28587,N_29653);
nand U31336 (N_31336,N_28892,N_28395);
nand U31337 (N_31337,N_29390,N_28992);
nor U31338 (N_31338,N_29758,N_27929);
nand U31339 (N_31339,N_28082,N_27924);
or U31340 (N_31340,N_28104,N_27824);
nor U31341 (N_31341,N_28599,N_27500);
and U31342 (N_31342,N_28112,N_29364);
nor U31343 (N_31343,N_29977,N_29449);
xor U31344 (N_31344,N_29900,N_28310);
xnor U31345 (N_31345,N_29227,N_27688);
or U31346 (N_31346,N_29730,N_28816);
and U31347 (N_31347,N_29003,N_28435);
nand U31348 (N_31348,N_29518,N_29245);
and U31349 (N_31349,N_27584,N_28128);
and U31350 (N_31350,N_27801,N_28872);
and U31351 (N_31351,N_29503,N_29142);
xnor U31352 (N_31352,N_29519,N_28163);
and U31353 (N_31353,N_28640,N_29280);
and U31354 (N_31354,N_28745,N_29897);
and U31355 (N_31355,N_28653,N_29451);
nand U31356 (N_31356,N_29760,N_29347);
nand U31357 (N_31357,N_29971,N_29361);
or U31358 (N_31358,N_27986,N_29019);
nand U31359 (N_31359,N_29636,N_28601);
xnor U31360 (N_31360,N_27536,N_28654);
or U31361 (N_31361,N_27793,N_27959);
or U31362 (N_31362,N_29533,N_28822);
nor U31363 (N_31363,N_27710,N_29991);
nor U31364 (N_31364,N_28336,N_29466);
nor U31365 (N_31365,N_29919,N_27871);
or U31366 (N_31366,N_29877,N_29550);
nand U31367 (N_31367,N_28474,N_27933);
or U31368 (N_31368,N_27877,N_29478);
nor U31369 (N_31369,N_28308,N_29059);
nor U31370 (N_31370,N_27730,N_29843);
and U31371 (N_31371,N_28980,N_28684);
nor U31372 (N_31372,N_28843,N_29562);
nor U31373 (N_31373,N_27839,N_29318);
nand U31374 (N_31374,N_27698,N_28784);
or U31375 (N_31375,N_27585,N_29430);
and U31376 (N_31376,N_27923,N_28477);
nand U31377 (N_31377,N_29873,N_28248);
and U31378 (N_31378,N_28890,N_28959);
nand U31379 (N_31379,N_29110,N_29886);
nand U31380 (N_31380,N_29884,N_28371);
nor U31381 (N_31381,N_28470,N_28341);
or U31382 (N_31382,N_27706,N_28543);
or U31383 (N_31383,N_28115,N_29087);
or U31384 (N_31384,N_28094,N_29285);
and U31385 (N_31385,N_28067,N_29810);
and U31386 (N_31386,N_27637,N_29539);
nand U31387 (N_31387,N_29573,N_27723);
nand U31388 (N_31388,N_27504,N_27567);
nor U31389 (N_31389,N_29926,N_29044);
or U31390 (N_31390,N_29762,N_28767);
or U31391 (N_31391,N_27675,N_28234);
xnor U31392 (N_31392,N_28765,N_29703);
xnor U31393 (N_31393,N_29180,N_27770);
or U31394 (N_31394,N_29066,N_29254);
and U31395 (N_31395,N_29924,N_28870);
or U31396 (N_31396,N_28784,N_29059);
or U31397 (N_31397,N_28601,N_28847);
or U31398 (N_31398,N_29976,N_28707);
nand U31399 (N_31399,N_27695,N_29831);
or U31400 (N_31400,N_29215,N_29539);
or U31401 (N_31401,N_28472,N_28019);
nand U31402 (N_31402,N_28278,N_29655);
nor U31403 (N_31403,N_29351,N_29291);
nor U31404 (N_31404,N_27587,N_29393);
or U31405 (N_31405,N_27587,N_29099);
and U31406 (N_31406,N_29806,N_28186);
and U31407 (N_31407,N_28333,N_28065);
nand U31408 (N_31408,N_28226,N_29403);
or U31409 (N_31409,N_27642,N_29073);
nor U31410 (N_31410,N_29897,N_29529);
and U31411 (N_31411,N_29310,N_27718);
nor U31412 (N_31412,N_28634,N_27943);
nor U31413 (N_31413,N_28650,N_28818);
or U31414 (N_31414,N_29478,N_27615);
or U31415 (N_31415,N_27530,N_29215);
or U31416 (N_31416,N_29343,N_29233);
nand U31417 (N_31417,N_28263,N_29194);
nor U31418 (N_31418,N_27644,N_29328);
nand U31419 (N_31419,N_29813,N_29009);
nand U31420 (N_31420,N_28182,N_28798);
nor U31421 (N_31421,N_28586,N_29938);
xor U31422 (N_31422,N_28406,N_27579);
nand U31423 (N_31423,N_29916,N_28706);
or U31424 (N_31424,N_29218,N_29347);
nor U31425 (N_31425,N_27970,N_27555);
xnor U31426 (N_31426,N_28445,N_29210);
nand U31427 (N_31427,N_29670,N_28113);
and U31428 (N_31428,N_28928,N_28876);
nor U31429 (N_31429,N_27934,N_28127);
nor U31430 (N_31430,N_29057,N_28172);
nand U31431 (N_31431,N_29169,N_27745);
or U31432 (N_31432,N_29978,N_28043);
and U31433 (N_31433,N_29531,N_29595);
and U31434 (N_31434,N_29007,N_28267);
and U31435 (N_31435,N_29270,N_29485);
xnor U31436 (N_31436,N_29498,N_28805);
nor U31437 (N_31437,N_29613,N_29243);
nor U31438 (N_31438,N_27979,N_28852);
xor U31439 (N_31439,N_27993,N_28880);
nand U31440 (N_31440,N_28324,N_29458);
nor U31441 (N_31441,N_29948,N_28402);
xnor U31442 (N_31442,N_29264,N_27985);
or U31443 (N_31443,N_27818,N_29495);
or U31444 (N_31444,N_27990,N_28830);
nor U31445 (N_31445,N_28479,N_28013);
nand U31446 (N_31446,N_27773,N_29072);
nand U31447 (N_31447,N_28240,N_28633);
nand U31448 (N_31448,N_28825,N_29009);
and U31449 (N_31449,N_28669,N_28654);
and U31450 (N_31450,N_28767,N_28880);
xor U31451 (N_31451,N_29129,N_27845);
nor U31452 (N_31452,N_27672,N_28802);
nor U31453 (N_31453,N_28994,N_28651);
and U31454 (N_31454,N_28802,N_27915);
or U31455 (N_31455,N_28048,N_29871);
nor U31456 (N_31456,N_29201,N_27502);
or U31457 (N_31457,N_28476,N_28975);
or U31458 (N_31458,N_29147,N_28700);
nor U31459 (N_31459,N_28788,N_27556);
nor U31460 (N_31460,N_29448,N_29774);
nor U31461 (N_31461,N_29253,N_29386);
or U31462 (N_31462,N_27876,N_29642);
or U31463 (N_31463,N_29168,N_29854);
or U31464 (N_31464,N_28298,N_29555);
or U31465 (N_31465,N_27848,N_29622);
or U31466 (N_31466,N_29127,N_27512);
or U31467 (N_31467,N_29117,N_29008);
nand U31468 (N_31468,N_27671,N_29961);
nor U31469 (N_31469,N_29230,N_29906);
or U31470 (N_31470,N_28509,N_29834);
and U31471 (N_31471,N_28716,N_29185);
nand U31472 (N_31472,N_29100,N_28513);
and U31473 (N_31473,N_27664,N_28638);
nor U31474 (N_31474,N_27614,N_29631);
or U31475 (N_31475,N_27867,N_28868);
or U31476 (N_31476,N_29499,N_27669);
and U31477 (N_31477,N_28847,N_28229);
and U31478 (N_31478,N_27707,N_29247);
nand U31479 (N_31479,N_28229,N_28667);
xnor U31480 (N_31480,N_28733,N_29267);
and U31481 (N_31481,N_29869,N_29195);
or U31482 (N_31482,N_29598,N_28526);
and U31483 (N_31483,N_27667,N_29724);
nand U31484 (N_31484,N_28624,N_28108);
xnor U31485 (N_31485,N_29606,N_29234);
nand U31486 (N_31486,N_27770,N_29454);
nand U31487 (N_31487,N_28126,N_29959);
and U31488 (N_31488,N_28699,N_27890);
nand U31489 (N_31489,N_28484,N_27780);
and U31490 (N_31490,N_27834,N_27977);
or U31491 (N_31491,N_29491,N_28299);
and U31492 (N_31492,N_27776,N_29057);
xnor U31493 (N_31493,N_29233,N_28695);
nand U31494 (N_31494,N_29970,N_27757);
and U31495 (N_31495,N_29044,N_28327);
nor U31496 (N_31496,N_29488,N_29286);
nor U31497 (N_31497,N_29565,N_28410);
xor U31498 (N_31498,N_28308,N_29237);
or U31499 (N_31499,N_29388,N_27507);
xor U31500 (N_31500,N_28296,N_29766);
nand U31501 (N_31501,N_29977,N_28670);
and U31502 (N_31502,N_28549,N_28842);
nand U31503 (N_31503,N_28096,N_27594);
nand U31504 (N_31504,N_27691,N_27960);
nor U31505 (N_31505,N_28969,N_27730);
nor U31506 (N_31506,N_29441,N_29258);
and U31507 (N_31507,N_27781,N_29803);
nor U31508 (N_31508,N_29526,N_29985);
nor U31509 (N_31509,N_29284,N_29665);
nand U31510 (N_31510,N_27511,N_29602);
or U31511 (N_31511,N_27549,N_29754);
nor U31512 (N_31512,N_29556,N_29362);
nand U31513 (N_31513,N_28894,N_28881);
nand U31514 (N_31514,N_29641,N_29319);
nand U31515 (N_31515,N_28065,N_27701);
nand U31516 (N_31516,N_28723,N_29519);
nor U31517 (N_31517,N_29583,N_28008);
nor U31518 (N_31518,N_29357,N_29516);
and U31519 (N_31519,N_28223,N_28164);
or U31520 (N_31520,N_29195,N_27507);
xnor U31521 (N_31521,N_29562,N_28623);
and U31522 (N_31522,N_28848,N_28430);
nand U31523 (N_31523,N_27578,N_29093);
nand U31524 (N_31524,N_29989,N_28768);
nor U31525 (N_31525,N_28860,N_28010);
nand U31526 (N_31526,N_28615,N_29536);
and U31527 (N_31527,N_28903,N_28233);
nor U31528 (N_31528,N_29380,N_28505);
or U31529 (N_31529,N_28848,N_29348);
nor U31530 (N_31530,N_28971,N_29312);
or U31531 (N_31531,N_27635,N_28965);
nor U31532 (N_31532,N_29634,N_28018);
and U31533 (N_31533,N_28811,N_27705);
nor U31534 (N_31534,N_28861,N_27857);
and U31535 (N_31535,N_27844,N_27829);
or U31536 (N_31536,N_28093,N_27573);
or U31537 (N_31537,N_27914,N_29670);
or U31538 (N_31538,N_29178,N_29309);
xnor U31539 (N_31539,N_28619,N_28238);
nor U31540 (N_31540,N_28720,N_29218);
nor U31541 (N_31541,N_27849,N_29679);
nor U31542 (N_31542,N_29682,N_28335);
xor U31543 (N_31543,N_27566,N_29284);
nor U31544 (N_31544,N_28012,N_28769);
and U31545 (N_31545,N_29339,N_29572);
nor U31546 (N_31546,N_28953,N_27947);
nand U31547 (N_31547,N_28548,N_29333);
xor U31548 (N_31548,N_27505,N_28934);
xnor U31549 (N_31549,N_29412,N_29729);
or U31550 (N_31550,N_28912,N_29061);
nor U31551 (N_31551,N_27911,N_28893);
nand U31552 (N_31552,N_28734,N_29847);
and U31553 (N_31553,N_28402,N_29401);
xor U31554 (N_31554,N_28047,N_28163);
nor U31555 (N_31555,N_28546,N_28366);
and U31556 (N_31556,N_27536,N_28593);
and U31557 (N_31557,N_29460,N_28241);
and U31558 (N_31558,N_27666,N_27537);
nor U31559 (N_31559,N_28624,N_28990);
nand U31560 (N_31560,N_28331,N_29040);
nor U31561 (N_31561,N_29939,N_28567);
nand U31562 (N_31562,N_28558,N_28779);
and U31563 (N_31563,N_29794,N_28491);
and U31564 (N_31564,N_29582,N_28932);
nand U31565 (N_31565,N_28582,N_29484);
nor U31566 (N_31566,N_27743,N_29021);
nor U31567 (N_31567,N_29829,N_28427);
and U31568 (N_31568,N_28102,N_28794);
and U31569 (N_31569,N_28622,N_28515);
or U31570 (N_31570,N_29212,N_29670);
nor U31571 (N_31571,N_28126,N_29153);
nand U31572 (N_31572,N_27855,N_28383);
or U31573 (N_31573,N_27993,N_28312);
or U31574 (N_31574,N_28797,N_27688);
or U31575 (N_31575,N_29406,N_29003);
xnor U31576 (N_31576,N_28970,N_28273);
or U31577 (N_31577,N_28869,N_28596);
or U31578 (N_31578,N_28077,N_28114);
nand U31579 (N_31579,N_27895,N_29186);
nor U31580 (N_31580,N_28824,N_27538);
and U31581 (N_31581,N_27786,N_28351);
xnor U31582 (N_31582,N_27699,N_27894);
nand U31583 (N_31583,N_27980,N_28459);
nand U31584 (N_31584,N_29432,N_28693);
xnor U31585 (N_31585,N_28034,N_29669);
nor U31586 (N_31586,N_29519,N_29692);
or U31587 (N_31587,N_28336,N_28957);
or U31588 (N_31588,N_29599,N_28001);
or U31589 (N_31589,N_29582,N_28177);
or U31590 (N_31590,N_28621,N_29049);
xor U31591 (N_31591,N_28846,N_27623);
or U31592 (N_31592,N_29510,N_27872);
or U31593 (N_31593,N_29143,N_27623);
and U31594 (N_31594,N_28763,N_28185);
nand U31595 (N_31595,N_28550,N_27892);
and U31596 (N_31596,N_29269,N_28944);
nand U31597 (N_31597,N_29852,N_29919);
nor U31598 (N_31598,N_27588,N_27556);
and U31599 (N_31599,N_28875,N_29077);
nand U31600 (N_31600,N_28591,N_28089);
xor U31601 (N_31601,N_27679,N_28186);
nor U31602 (N_31602,N_29273,N_27546);
or U31603 (N_31603,N_28982,N_29096);
xor U31604 (N_31604,N_27563,N_28671);
or U31605 (N_31605,N_29165,N_28921);
nand U31606 (N_31606,N_29822,N_29618);
or U31607 (N_31607,N_28938,N_27513);
nand U31608 (N_31608,N_28120,N_28152);
or U31609 (N_31609,N_28665,N_28806);
nor U31610 (N_31610,N_27996,N_29314);
nand U31611 (N_31611,N_27595,N_28785);
or U31612 (N_31612,N_29035,N_29348);
nor U31613 (N_31613,N_28668,N_28837);
and U31614 (N_31614,N_27539,N_28036);
nor U31615 (N_31615,N_27598,N_29226);
or U31616 (N_31616,N_27586,N_28476);
or U31617 (N_31617,N_27858,N_29109);
and U31618 (N_31618,N_29232,N_27975);
nor U31619 (N_31619,N_29136,N_29345);
xor U31620 (N_31620,N_29179,N_29200);
nor U31621 (N_31621,N_27894,N_28371);
nor U31622 (N_31622,N_29754,N_28797);
nor U31623 (N_31623,N_29276,N_28201);
nand U31624 (N_31624,N_27753,N_28763);
or U31625 (N_31625,N_27565,N_29847);
and U31626 (N_31626,N_28876,N_28729);
nor U31627 (N_31627,N_28906,N_28758);
nand U31628 (N_31628,N_29001,N_28629);
nand U31629 (N_31629,N_28312,N_28119);
and U31630 (N_31630,N_29633,N_29293);
or U31631 (N_31631,N_28794,N_28817);
or U31632 (N_31632,N_27872,N_28446);
nor U31633 (N_31633,N_29412,N_29138);
xor U31634 (N_31634,N_28867,N_29135);
xor U31635 (N_31635,N_28153,N_28203);
nor U31636 (N_31636,N_29029,N_29564);
nand U31637 (N_31637,N_28993,N_28645);
xnor U31638 (N_31638,N_28703,N_28953);
nor U31639 (N_31639,N_29987,N_28742);
and U31640 (N_31640,N_28119,N_28457);
and U31641 (N_31641,N_29999,N_28756);
nor U31642 (N_31642,N_28443,N_29049);
or U31643 (N_31643,N_28335,N_29330);
nor U31644 (N_31644,N_27846,N_28200);
nand U31645 (N_31645,N_28446,N_29231);
nor U31646 (N_31646,N_28219,N_28568);
nand U31647 (N_31647,N_27630,N_27755);
nand U31648 (N_31648,N_28976,N_28704);
nor U31649 (N_31649,N_28900,N_28582);
nand U31650 (N_31650,N_28121,N_28265);
nor U31651 (N_31651,N_29674,N_29024);
nand U31652 (N_31652,N_28552,N_29816);
and U31653 (N_31653,N_28345,N_28307);
xnor U31654 (N_31654,N_27974,N_29814);
xor U31655 (N_31655,N_28714,N_28337);
nand U31656 (N_31656,N_29403,N_28261);
nor U31657 (N_31657,N_27900,N_28086);
nor U31658 (N_31658,N_27911,N_28720);
xor U31659 (N_31659,N_28497,N_27558);
or U31660 (N_31660,N_29021,N_29534);
or U31661 (N_31661,N_29980,N_27626);
nand U31662 (N_31662,N_29751,N_27757);
nand U31663 (N_31663,N_28753,N_29588);
nor U31664 (N_31664,N_27692,N_29215);
nand U31665 (N_31665,N_29192,N_29013);
xnor U31666 (N_31666,N_27811,N_29785);
nor U31667 (N_31667,N_27684,N_29118);
and U31668 (N_31668,N_28846,N_28577);
and U31669 (N_31669,N_29873,N_27859);
nand U31670 (N_31670,N_28956,N_29656);
xnor U31671 (N_31671,N_28141,N_27683);
or U31672 (N_31672,N_29901,N_29845);
nand U31673 (N_31673,N_27987,N_29702);
or U31674 (N_31674,N_27765,N_27992);
nand U31675 (N_31675,N_29080,N_28975);
nor U31676 (N_31676,N_28014,N_27925);
nand U31677 (N_31677,N_28295,N_27688);
xor U31678 (N_31678,N_28599,N_29653);
and U31679 (N_31679,N_29881,N_29268);
and U31680 (N_31680,N_29474,N_28843);
nor U31681 (N_31681,N_28602,N_28021);
or U31682 (N_31682,N_29194,N_29400);
and U31683 (N_31683,N_28237,N_29532);
nor U31684 (N_31684,N_29283,N_28180);
nand U31685 (N_31685,N_28332,N_28222);
xor U31686 (N_31686,N_28189,N_29458);
xor U31687 (N_31687,N_28460,N_28571);
and U31688 (N_31688,N_27993,N_29748);
nor U31689 (N_31689,N_27602,N_29295);
or U31690 (N_31690,N_27735,N_27903);
nand U31691 (N_31691,N_28475,N_29286);
nor U31692 (N_31692,N_27634,N_29285);
nand U31693 (N_31693,N_29579,N_29590);
xnor U31694 (N_31694,N_28241,N_27931);
or U31695 (N_31695,N_28588,N_29376);
nand U31696 (N_31696,N_28305,N_27985);
nor U31697 (N_31697,N_27851,N_29865);
nand U31698 (N_31698,N_28944,N_29645);
nor U31699 (N_31699,N_29021,N_27930);
and U31700 (N_31700,N_29087,N_28045);
and U31701 (N_31701,N_29577,N_28646);
xnor U31702 (N_31702,N_29689,N_29246);
and U31703 (N_31703,N_27693,N_29779);
or U31704 (N_31704,N_29743,N_28739);
or U31705 (N_31705,N_27962,N_29583);
xnor U31706 (N_31706,N_29845,N_29127);
and U31707 (N_31707,N_29461,N_28820);
or U31708 (N_31708,N_28803,N_29162);
or U31709 (N_31709,N_28708,N_29878);
xor U31710 (N_31710,N_28665,N_29651);
xor U31711 (N_31711,N_28218,N_29840);
and U31712 (N_31712,N_29119,N_29574);
nor U31713 (N_31713,N_27926,N_28732);
nand U31714 (N_31714,N_28030,N_29123);
or U31715 (N_31715,N_28468,N_28204);
or U31716 (N_31716,N_28864,N_27978);
or U31717 (N_31717,N_28831,N_29483);
and U31718 (N_31718,N_28101,N_29232);
nor U31719 (N_31719,N_28515,N_29253);
and U31720 (N_31720,N_28799,N_29456);
xor U31721 (N_31721,N_28904,N_29269);
nor U31722 (N_31722,N_29523,N_29498);
xnor U31723 (N_31723,N_29062,N_29419);
or U31724 (N_31724,N_27529,N_29949);
and U31725 (N_31725,N_29891,N_29588);
and U31726 (N_31726,N_29530,N_28040);
nand U31727 (N_31727,N_29543,N_29501);
xnor U31728 (N_31728,N_27698,N_29687);
or U31729 (N_31729,N_29197,N_29668);
or U31730 (N_31730,N_29937,N_28097);
xor U31731 (N_31731,N_29197,N_29957);
xnor U31732 (N_31732,N_29453,N_28897);
xnor U31733 (N_31733,N_29711,N_29351);
xor U31734 (N_31734,N_27973,N_28803);
or U31735 (N_31735,N_28482,N_29779);
and U31736 (N_31736,N_29852,N_29101);
nand U31737 (N_31737,N_29155,N_29746);
or U31738 (N_31738,N_29961,N_27903);
xnor U31739 (N_31739,N_29885,N_29562);
or U31740 (N_31740,N_28591,N_27527);
nor U31741 (N_31741,N_29188,N_29270);
xor U31742 (N_31742,N_28650,N_29516);
nor U31743 (N_31743,N_28579,N_27981);
and U31744 (N_31744,N_28076,N_28673);
or U31745 (N_31745,N_29536,N_28888);
nor U31746 (N_31746,N_28515,N_29286);
nand U31747 (N_31747,N_28203,N_28480);
and U31748 (N_31748,N_27720,N_28751);
xor U31749 (N_31749,N_29195,N_28822);
or U31750 (N_31750,N_29392,N_29431);
or U31751 (N_31751,N_29168,N_28147);
and U31752 (N_31752,N_29903,N_28024);
xnor U31753 (N_31753,N_29898,N_29109);
nor U31754 (N_31754,N_29515,N_28339);
and U31755 (N_31755,N_29105,N_28241);
xor U31756 (N_31756,N_28283,N_29858);
nand U31757 (N_31757,N_29140,N_29531);
or U31758 (N_31758,N_28266,N_28728);
xor U31759 (N_31759,N_29566,N_27889);
and U31760 (N_31760,N_28997,N_28041);
and U31761 (N_31761,N_28109,N_27982);
or U31762 (N_31762,N_27783,N_29155);
or U31763 (N_31763,N_29336,N_29302);
xnor U31764 (N_31764,N_27883,N_28100);
nand U31765 (N_31765,N_27589,N_29945);
and U31766 (N_31766,N_28069,N_29019);
and U31767 (N_31767,N_29535,N_27948);
nand U31768 (N_31768,N_27846,N_29687);
or U31769 (N_31769,N_28785,N_29058);
and U31770 (N_31770,N_29649,N_27972);
nor U31771 (N_31771,N_27564,N_28492);
nor U31772 (N_31772,N_27890,N_28797);
xor U31773 (N_31773,N_28423,N_29042);
or U31774 (N_31774,N_28266,N_27681);
nand U31775 (N_31775,N_29712,N_28865);
xnor U31776 (N_31776,N_27969,N_28946);
nand U31777 (N_31777,N_29570,N_28943);
and U31778 (N_31778,N_29912,N_29787);
or U31779 (N_31779,N_29626,N_28864);
nor U31780 (N_31780,N_29294,N_28332);
and U31781 (N_31781,N_27847,N_29794);
nand U31782 (N_31782,N_27970,N_29833);
or U31783 (N_31783,N_28302,N_28189);
nand U31784 (N_31784,N_29712,N_28355);
and U31785 (N_31785,N_28351,N_28074);
and U31786 (N_31786,N_29981,N_29496);
nand U31787 (N_31787,N_28084,N_28576);
or U31788 (N_31788,N_29505,N_28542);
xnor U31789 (N_31789,N_28402,N_28378);
and U31790 (N_31790,N_29483,N_28420);
or U31791 (N_31791,N_27645,N_28934);
and U31792 (N_31792,N_29269,N_27979);
or U31793 (N_31793,N_28209,N_28072);
nor U31794 (N_31794,N_28464,N_28617);
and U31795 (N_31795,N_28981,N_29967);
nand U31796 (N_31796,N_28993,N_28971);
or U31797 (N_31797,N_28823,N_29183);
xnor U31798 (N_31798,N_27693,N_28535);
nand U31799 (N_31799,N_29553,N_29930);
or U31800 (N_31800,N_29539,N_28835);
nand U31801 (N_31801,N_29635,N_28761);
and U31802 (N_31802,N_28130,N_28028);
or U31803 (N_31803,N_29804,N_27599);
nand U31804 (N_31804,N_27829,N_27898);
xor U31805 (N_31805,N_28372,N_28627);
nand U31806 (N_31806,N_27762,N_27582);
xnor U31807 (N_31807,N_27540,N_28801);
xnor U31808 (N_31808,N_29767,N_28349);
and U31809 (N_31809,N_29415,N_29676);
or U31810 (N_31810,N_28730,N_29129);
xnor U31811 (N_31811,N_27880,N_29717);
or U31812 (N_31812,N_28605,N_28953);
or U31813 (N_31813,N_28837,N_29294);
nor U31814 (N_31814,N_28735,N_29499);
nand U31815 (N_31815,N_29922,N_29984);
nor U31816 (N_31816,N_29811,N_29013);
nand U31817 (N_31817,N_29854,N_28544);
and U31818 (N_31818,N_29606,N_27559);
and U31819 (N_31819,N_29562,N_28229);
or U31820 (N_31820,N_28612,N_28175);
and U31821 (N_31821,N_27554,N_29525);
nor U31822 (N_31822,N_29783,N_27845);
nand U31823 (N_31823,N_29492,N_29260);
and U31824 (N_31824,N_27744,N_28060);
and U31825 (N_31825,N_28639,N_27753);
or U31826 (N_31826,N_28859,N_28544);
nor U31827 (N_31827,N_28150,N_27706);
nor U31828 (N_31828,N_27618,N_28311);
or U31829 (N_31829,N_28222,N_29561);
nor U31830 (N_31830,N_29755,N_27879);
nand U31831 (N_31831,N_28258,N_27649);
nor U31832 (N_31832,N_28622,N_29137);
nor U31833 (N_31833,N_28857,N_28155);
nor U31834 (N_31834,N_27640,N_29113);
nand U31835 (N_31835,N_28620,N_29374);
or U31836 (N_31836,N_28546,N_28115);
nor U31837 (N_31837,N_29786,N_28318);
nand U31838 (N_31838,N_29200,N_28907);
nand U31839 (N_31839,N_29571,N_29959);
nor U31840 (N_31840,N_28395,N_28659);
or U31841 (N_31841,N_28223,N_29885);
nor U31842 (N_31842,N_27960,N_28263);
and U31843 (N_31843,N_29907,N_29642);
or U31844 (N_31844,N_28747,N_29244);
nor U31845 (N_31845,N_29256,N_28069);
and U31846 (N_31846,N_28000,N_28883);
or U31847 (N_31847,N_27708,N_27632);
or U31848 (N_31848,N_29970,N_29775);
or U31849 (N_31849,N_29773,N_29537);
or U31850 (N_31850,N_28097,N_29035);
and U31851 (N_31851,N_27995,N_28253);
xnor U31852 (N_31852,N_29305,N_29903);
nand U31853 (N_31853,N_28251,N_29791);
or U31854 (N_31854,N_28857,N_29718);
nand U31855 (N_31855,N_27916,N_28229);
or U31856 (N_31856,N_29766,N_28135);
or U31857 (N_31857,N_29934,N_29553);
nand U31858 (N_31858,N_29642,N_29778);
nor U31859 (N_31859,N_29172,N_28172);
or U31860 (N_31860,N_29358,N_29764);
nand U31861 (N_31861,N_27839,N_28711);
and U31862 (N_31862,N_28820,N_28212);
nor U31863 (N_31863,N_28453,N_27753);
nand U31864 (N_31864,N_27679,N_29051);
xor U31865 (N_31865,N_28121,N_28570);
or U31866 (N_31866,N_29765,N_28556);
nand U31867 (N_31867,N_29083,N_28384);
nor U31868 (N_31868,N_29293,N_28324);
nor U31869 (N_31869,N_28230,N_29723);
nand U31870 (N_31870,N_29061,N_29799);
nand U31871 (N_31871,N_29734,N_29446);
xor U31872 (N_31872,N_27692,N_28389);
and U31873 (N_31873,N_29316,N_27647);
and U31874 (N_31874,N_27832,N_29181);
xor U31875 (N_31875,N_29603,N_28388);
nand U31876 (N_31876,N_27693,N_28544);
nand U31877 (N_31877,N_27538,N_29870);
or U31878 (N_31878,N_28794,N_29853);
and U31879 (N_31879,N_28725,N_29848);
or U31880 (N_31880,N_29472,N_28853);
nand U31881 (N_31881,N_27544,N_28099);
nor U31882 (N_31882,N_29128,N_29687);
nand U31883 (N_31883,N_29942,N_29797);
nor U31884 (N_31884,N_28168,N_27788);
or U31885 (N_31885,N_29945,N_29460);
or U31886 (N_31886,N_28203,N_28687);
or U31887 (N_31887,N_29919,N_27565);
xor U31888 (N_31888,N_28425,N_28004);
or U31889 (N_31889,N_27882,N_28144);
nand U31890 (N_31890,N_29842,N_28718);
nand U31891 (N_31891,N_29955,N_28594);
nor U31892 (N_31892,N_28247,N_28225);
xnor U31893 (N_31893,N_29598,N_27770);
nand U31894 (N_31894,N_28318,N_29774);
nand U31895 (N_31895,N_27672,N_27524);
or U31896 (N_31896,N_29003,N_27912);
nand U31897 (N_31897,N_28863,N_28258);
or U31898 (N_31898,N_28343,N_29399);
and U31899 (N_31899,N_29066,N_28692);
nand U31900 (N_31900,N_28596,N_29954);
nand U31901 (N_31901,N_27741,N_29411);
xor U31902 (N_31902,N_28789,N_27640);
nor U31903 (N_31903,N_27896,N_28367);
or U31904 (N_31904,N_29519,N_28606);
or U31905 (N_31905,N_28430,N_29685);
xor U31906 (N_31906,N_29910,N_29446);
xor U31907 (N_31907,N_29812,N_29881);
nand U31908 (N_31908,N_28406,N_28479);
nand U31909 (N_31909,N_28046,N_28831);
or U31910 (N_31910,N_28948,N_29384);
nor U31911 (N_31911,N_27804,N_28046);
and U31912 (N_31912,N_28634,N_27570);
and U31913 (N_31913,N_28101,N_29431);
nand U31914 (N_31914,N_29984,N_29227);
and U31915 (N_31915,N_27939,N_28547);
nor U31916 (N_31916,N_27737,N_27798);
nand U31917 (N_31917,N_29054,N_27914);
xor U31918 (N_31918,N_28303,N_28219);
nor U31919 (N_31919,N_28458,N_29910);
xnor U31920 (N_31920,N_29159,N_29065);
or U31921 (N_31921,N_27938,N_28495);
or U31922 (N_31922,N_29817,N_29055);
or U31923 (N_31923,N_29462,N_29750);
nand U31924 (N_31924,N_28444,N_29731);
nor U31925 (N_31925,N_29073,N_27939);
xnor U31926 (N_31926,N_29330,N_28482);
nand U31927 (N_31927,N_29650,N_29893);
and U31928 (N_31928,N_29918,N_29198);
nor U31929 (N_31929,N_29172,N_28921);
nor U31930 (N_31930,N_28428,N_28945);
nor U31931 (N_31931,N_28724,N_28328);
or U31932 (N_31932,N_28313,N_27923);
or U31933 (N_31933,N_27920,N_28995);
nand U31934 (N_31934,N_29317,N_27791);
nor U31935 (N_31935,N_29134,N_27984);
or U31936 (N_31936,N_28184,N_28138);
and U31937 (N_31937,N_28811,N_28705);
and U31938 (N_31938,N_29385,N_29597);
nor U31939 (N_31939,N_29891,N_29932);
or U31940 (N_31940,N_29317,N_29047);
nand U31941 (N_31941,N_27826,N_27725);
or U31942 (N_31942,N_27695,N_28591);
nand U31943 (N_31943,N_29636,N_27693);
nor U31944 (N_31944,N_28157,N_29711);
xnor U31945 (N_31945,N_28443,N_29598);
nand U31946 (N_31946,N_28109,N_27609);
nand U31947 (N_31947,N_29803,N_28039);
or U31948 (N_31948,N_29691,N_27621);
nand U31949 (N_31949,N_28873,N_29934);
nand U31950 (N_31950,N_29847,N_29412);
nor U31951 (N_31951,N_29247,N_27562);
nor U31952 (N_31952,N_29157,N_28124);
xnor U31953 (N_31953,N_27852,N_29080);
and U31954 (N_31954,N_29434,N_29932);
or U31955 (N_31955,N_28660,N_29457);
or U31956 (N_31956,N_28567,N_28616);
or U31957 (N_31957,N_27683,N_29491);
and U31958 (N_31958,N_28591,N_27540);
or U31959 (N_31959,N_28622,N_29734);
and U31960 (N_31960,N_29750,N_28637);
and U31961 (N_31961,N_27571,N_29347);
xnor U31962 (N_31962,N_27937,N_27748);
nor U31963 (N_31963,N_28915,N_28465);
nor U31964 (N_31964,N_27678,N_29021);
xor U31965 (N_31965,N_29932,N_28223);
and U31966 (N_31966,N_27735,N_29979);
or U31967 (N_31967,N_29023,N_27565);
xor U31968 (N_31968,N_29214,N_28727);
or U31969 (N_31969,N_28560,N_28101);
nor U31970 (N_31970,N_29527,N_28948);
nor U31971 (N_31971,N_28799,N_27716);
nand U31972 (N_31972,N_29567,N_28842);
or U31973 (N_31973,N_28957,N_28448);
or U31974 (N_31974,N_28976,N_28119);
or U31975 (N_31975,N_28257,N_28900);
xor U31976 (N_31976,N_27883,N_28303);
nand U31977 (N_31977,N_29101,N_29513);
and U31978 (N_31978,N_27858,N_27927);
or U31979 (N_31979,N_27835,N_28204);
xor U31980 (N_31980,N_28646,N_29259);
nand U31981 (N_31981,N_27509,N_27796);
xor U31982 (N_31982,N_28700,N_28296);
xor U31983 (N_31983,N_27526,N_29175);
xnor U31984 (N_31984,N_29520,N_28719);
or U31985 (N_31985,N_28151,N_29691);
or U31986 (N_31986,N_27711,N_28913);
nor U31987 (N_31987,N_27964,N_29809);
nor U31988 (N_31988,N_28555,N_29184);
and U31989 (N_31989,N_28026,N_29963);
and U31990 (N_31990,N_28747,N_29861);
or U31991 (N_31991,N_27702,N_28507);
nand U31992 (N_31992,N_29063,N_27535);
and U31993 (N_31993,N_28152,N_29674);
nor U31994 (N_31994,N_29629,N_28137);
or U31995 (N_31995,N_28625,N_27758);
nor U31996 (N_31996,N_29043,N_28561);
nor U31997 (N_31997,N_29352,N_29405);
or U31998 (N_31998,N_28348,N_28498);
and U31999 (N_31999,N_27677,N_29455);
xor U32000 (N_32000,N_28566,N_29706);
and U32001 (N_32001,N_28128,N_28649);
nor U32002 (N_32002,N_29415,N_27820);
nor U32003 (N_32003,N_27557,N_29424);
or U32004 (N_32004,N_29591,N_29331);
nand U32005 (N_32005,N_29243,N_28238);
nor U32006 (N_32006,N_27635,N_27571);
xnor U32007 (N_32007,N_28390,N_29283);
or U32008 (N_32008,N_27981,N_27741);
nor U32009 (N_32009,N_29705,N_29017);
and U32010 (N_32010,N_28492,N_29423);
and U32011 (N_32011,N_29537,N_28973);
or U32012 (N_32012,N_28633,N_29304);
xnor U32013 (N_32013,N_27644,N_29208);
or U32014 (N_32014,N_28797,N_29309);
and U32015 (N_32015,N_27754,N_29872);
and U32016 (N_32016,N_27806,N_29223);
and U32017 (N_32017,N_29724,N_29195);
xor U32018 (N_32018,N_28860,N_28106);
nor U32019 (N_32019,N_28399,N_28234);
or U32020 (N_32020,N_28556,N_28006);
nand U32021 (N_32021,N_27568,N_28869);
nand U32022 (N_32022,N_29166,N_29151);
nand U32023 (N_32023,N_28433,N_28431);
xor U32024 (N_32024,N_29499,N_29544);
nor U32025 (N_32025,N_28315,N_28995);
nor U32026 (N_32026,N_28416,N_29261);
nor U32027 (N_32027,N_27807,N_28732);
xnor U32028 (N_32028,N_28441,N_29854);
nand U32029 (N_32029,N_28864,N_29434);
or U32030 (N_32030,N_29223,N_29566);
or U32031 (N_32031,N_28971,N_29831);
or U32032 (N_32032,N_29441,N_28144);
nor U32033 (N_32033,N_27809,N_27692);
nand U32034 (N_32034,N_27776,N_28815);
xor U32035 (N_32035,N_28476,N_29552);
nand U32036 (N_32036,N_29693,N_28367);
and U32037 (N_32037,N_28225,N_29914);
and U32038 (N_32038,N_28543,N_28918);
xor U32039 (N_32039,N_27843,N_29445);
nor U32040 (N_32040,N_28707,N_28677);
nand U32041 (N_32041,N_28908,N_29692);
nand U32042 (N_32042,N_29802,N_29326);
xnor U32043 (N_32043,N_29025,N_28612);
xor U32044 (N_32044,N_28848,N_28004);
and U32045 (N_32045,N_28063,N_28670);
and U32046 (N_32046,N_27969,N_27762);
nor U32047 (N_32047,N_28783,N_29478);
nor U32048 (N_32048,N_27777,N_28782);
nor U32049 (N_32049,N_29921,N_29941);
nand U32050 (N_32050,N_27610,N_27564);
nor U32051 (N_32051,N_29287,N_28085);
xor U32052 (N_32052,N_28604,N_28316);
nor U32053 (N_32053,N_28599,N_29234);
and U32054 (N_32054,N_27605,N_29187);
nand U32055 (N_32055,N_29541,N_29746);
nand U32056 (N_32056,N_28069,N_28459);
nand U32057 (N_32057,N_29057,N_28923);
nand U32058 (N_32058,N_27972,N_28521);
nand U32059 (N_32059,N_29924,N_28373);
and U32060 (N_32060,N_28267,N_28906);
nor U32061 (N_32061,N_28548,N_28290);
or U32062 (N_32062,N_28066,N_29401);
and U32063 (N_32063,N_28916,N_27529);
nor U32064 (N_32064,N_29617,N_29038);
and U32065 (N_32065,N_27560,N_27887);
and U32066 (N_32066,N_27983,N_28932);
and U32067 (N_32067,N_27812,N_27503);
nor U32068 (N_32068,N_29143,N_29361);
xnor U32069 (N_32069,N_28221,N_28231);
xnor U32070 (N_32070,N_29739,N_28770);
or U32071 (N_32071,N_29513,N_28965);
nor U32072 (N_32072,N_29740,N_29906);
and U32073 (N_32073,N_27521,N_29062);
nor U32074 (N_32074,N_28024,N_29606);
nand U32075 (N_32075,N_28703,N_27887);
and U32076 (N_32076,N_29452,N_29124);
and U32077 (N_32077,N_29459,N_28310);
or U32078 (N_32078,N_29584,N_29062);
nor U32079 (N_32079,N_29615,N_27505);
nor U32080 (N_32080,N_28037,N_29601);
nand U32081 (N_32081,N_27526,N_28011);
and U32082 (N_32082,N_29733,N_29953);
nand U32083 (N_32083,N_27614,N_28680);
nor U32084 (N_32084,N_29844,N_28173);
nor U32085 (N_32085,N_28387,N_29470);
nor U32086 (N_32086,N_27515,N_29406);
nand U32087 (N_32087,N_29785,N_27918);
nor U32088 (N_32088,N_28346,N_29186);
and U32089 (N_32089,N_28449,N_29396);
or U32090 (N_32090,N_28380,N_29495);
or U32091 (N_32091,N_28601,N_29540);
and U32092 (N_32092,N_28083,N_29982);
nand U32093 (N_32093,N_28553,N_28379);
nand U32094 (N_32094,N_28773,N_29895);
and U32095 (N_32095,N_27536,N_28558);
xor U32096 (N_32096,N_28594,N_28230);
nor U32097 (N_32097,N_29293,N_29942);
nand U32098 (N_32098,N_28124,N_29042);
and U32099 (N_32099,N_28219,N_28980);
or U32100 (N_32100,N_29686,N_29627);
and U32101 (N_32101,N_27585,N_28637);
xnor U32102 (N_32102,N_28928,N_27731);
nand U32103 (N_32103,N_29178,N_28020);
nand U32104 (N_32104,N_27976,N_29202);
and U32105 (N_32105,N_29129,N_29002);
nor U32106 (N_32106,N_29226,N_28847);
nand U32107 (N_32107,N_27648,N_29788);
and U32108 (N_32108,N_28163,N_28765);
nor U32109 (N_32109,N_27540,N_28902);
and U32110 (N_32110,N_29779,N_29975);
or U32111 (N_32111,N_27990,N_27920);
and U32112 (N_32112,N_29037,N_28385);
or U32113 (N_32113,N_28011,N_28627);
or U32114 (N_32114,N_28420,N_29485);
and U32115 (N_32115,N_27604,N_28042);
nor U32116 (N_32116,N_27623,N_29507);
or U32117 (N_32117,N_28758,N_29433);
nand U32118 (N_32118,N_28931,N_29639);
and U32119 (N_32119,N_28205,N_29929);
nand U32120 (N_32120,N_27754,N_29480);
nand U32121 (N_32121,N_27992,N_28849);
or U32122 (N_32122,N_29487,N_27673);
or U32123 (N_32123,N_28017,N_27835);
nor U32124 (N_32124,N_28953,N_29810);
xnor U32125 (N_32125,N_29508,N_28822);
or U32126 (N_32126,N_28417,N_28328);
xnor U32127 (N_32127,N_29381,N_27689);
nand U32128 (N_32128,N_27538,N_29270);
nand U32129 (N_32129,N_29951,N_29188);
nor U32130 (N_32130,N_28227,N_27791);
and U32131 (N_32131,N_28491,N_27749);
nor U32132 (N_32132,N_28402,N_29642);
nor U32133 (N_32133,N_27821,N_27969);
nand U32134 (N_32134,N_29655,N_29698);
nor U32135 (N_32135,N_27751,N_28282);
or U32136 (N_32136,N_29507,N_28666);
and U32137 (N_32137,N_28355,N_27537);
and U32138 (N_32138,N_28250,N_28341);
xor U32139 (N_32139,N_27802,N_29804);
nand U32140 (N_32140,N_27528,N_29008);
and U32141 (N_32141,N_28941,N_27593);
and U32142 (N_32142,N_29171,N_28247);
and U32143 (N_32143,N_28310,N_29358);
nand U32144 (N_32144,N_29998,N_27671);
and U32145 (N_32145,N_28436,N_28708);
xnor U32146 (N_32146,N_28267,N_29646);
nor U32147 (N_32147,N_29177,N_28742);
nand U32148 (N_32148,N_28048,N_29226);
and U32149 (N_32149,N_28828,N_29419);
nor U32150 (N_32150,N_28210,N_29341);
nor U32151 (N_32151,N_28477,N_29308);
xnor U32152 (N_32152,N_28338,N_27930);
nor U32153 (N_32153,N_29986,N_29006);
nand U32154 (N_32154,N_29325,N_28041);
and U32155 (N_32155,N_29575,N_29256);
nor U32156 (N_32156,N_29556,N_29383);
nand U32157 (N_32157,N_29918,N_27689);
xor U32158 (N_32158,N_29537,N_29983);
nand U32159 (N_32159,N_28481,N_29017);
nor U32160 (N_32160,N_28818,N_28712);
nor U32161 (N_32161,N_29567,N_28741);
xnor U32162 (N_32162,N_28854,N_28506);
or U32163 (N_32163,N_27869,N_29657);
and U32164 (N_32164,N_28356,N_28877);
xor U32165 (N_32165,N_28825,N_27613);
nor U32166 (N_32166,N_29020,N_27819);
or U32167 (N_32167,N_28310,N_29052);
nand U32168 (N_32168,N_29311,N_29275);
and U32169 (N_32169,N_29287,N_28841);
or U32170 (N_32170,N_28706,N_27685);
nand U32171 (N_32171,N_27609,N_27905);
nor U32172 (N_32172,N_28183,N_29133);
nor U32173 (N_32173,N_29459,N_28662);
or U32174 (N_32174,N_27858,N_27527);
nor U32175 (N_32175,N_28162,N_29483);
nand U32176 (N_32176,N_28252,N_27637);
xor U32177 (N_32177,N_28848,N_28471);
nor U32178 (N_32178,N_28313,N_28762);
nand U32179 (N_32179,N_28870,N_27573);
or U32180 (N_32180,N_28479,N_29902);
nand U32181 (N_32181,N_27895,N_29471);
and U32182 (N_32182,N_29941,N_29901);
xnor U32183 (N_32183,N_29417,N_27675);
and U32184 (N_32184,N_29771,N_29136);
and U32185 (N_32185,N_28116,N_28552);
and U32186 (N_32186,N_29505,N_29620);
and U32187 (N_32187,N_29868,N_29800);
nand U32188 (N_32188,N_29820,N_27532);
and U32189 (N_32189,N_29409,N_29144);
and U32190 (N_32190,N_27800,N_27626);
nand U32191 (N_32191,N_29615,N_28053);
and U32192 (N_32192,N_27685,N_29265);
or U32193 (N_32193,N_29272,N_28877);
and U32194 (N_32194,N_29298,N_29214);
and U32195 (N_32195,N_28669,N_28106);
nor U32196 (N_32196,N_27642,N_29275);
or U32197 (N_32197,N_29818,N_28339);
nand U32198 (N_32198,N_28646,N_28701);
and U32199 (N_32199,N_29315,N_29052);
nor U32200 (N_32200,N_28407,N_28358);
or U32201 (N_32201,N_29541,N_27871);
and U32202 (N_32202,N_27691,N_29397);
or U32203 (N_32203,N_29714,N_28156);
xnor U32204 (N_32204,N_27751,N_29455);
nand U32205 (N_32205,N_27713,N_29252);
nor U32206 (N_32206,N_27653,N_28704);
nor U32207 (N_32207,N_27967,N_27884);
and U32208 (N_32208,N_28968,N_28148);
nand U32209 (N_32209,N_27826,N_29894);
and U32210 (N_32210,N_29973,N_27738);
nor U32211 (N_32211,N_29149,N_29882);
nor U32212 (N_32212,N_27906,N_28927);
xor U32213 (N_32213,N_29213,N_29660);
or U32214 (N_32214,N_28314,N_28110);
and U32215 (N_32215,N_28444,N_27609);
and U32216 (N_32216,N_29375,N_27719);
xor U32217 (N_32217,N_29495,N_28213);
or U32218 (N_32218,N_27651,N_27835);
and U32219 (N_32219,N_29483,N_28546);
or U32220 (N_32220,N_28608,N_29683);
and U32221 (N_32221,N_28225,N_29443);
and U32222 (N_32222,N_29863,N_29423);
or U32223 (N_32223,N_28062,N_29510);
nor U32224 (N_32224,N_28023,N_28766);
or U32225 (N_32225,N_27696,N_29543);
and U32226 (N_32226,N_29265,N_29458);
or U32227 (N_32227,N_29803,N_28489);
nor U32228 (N_32228,N_27576,N_29557);
or U32229 (N_32229,N_27576,N_29525);
xnor U32230 (N_32230,N_28867,N_28208);
and U32231 (N_32231,N_29773,N_27545);
nor U32232 (N_32232,N_27607,N_28686);
and U32233 (N_32233,N_28558,N_29051);
nand U32234 (N_32234,N_27999,N_28148);
nand U32235 (N_32235,N_28313,N_29558);
xnor U32236 (N_32236,N_29227,N_28570);
xor U32237 (N_32237,N_28046,N_29218);
nor U32238 (N_32238,N_28852,N_29184);
or U32239 (N_32239,N_29791,N_27659);
nor U32240 (N_32240,N_29904,N_28588);
nand U32241 (N_32241,N_29748,N_29326);
or U32242 (N_32242,N_27731,N_29771);
or U32243 (N_32243,N_29589,N_27790);
or U32244 (N_32244,N_28547,N_27549);
xor U32245 (N_32245,N_28105,N_29693);
or U32246 (N_32246,N_28341,N_28185);
nor U32247 (N_32247,N_27856,N_29128);
xnor U32248 (N_32248,N_29861,N_29727);
or U32249 (N_32249,N_29629,N_29684);
nor U32250 (N_32250,N_28146,N_27868);
xor U32251 (N_32251,N_28435,N_28591);
nor U32252 (N_32252,N_28927,N_29506);
nor U32253 (N_32253,N_28533,N_29290);
and U32254 (N_32254,N_29253,N_27761);
nor U32255 (N_32255,N_29998,N_28628);
and U32256 (N_32256,N_28683,N_29661);
or U32257 (N_32257,N_29935,N_27542);
or U32258 (N_32258,N_28305,N_28114);
xor U32259 (N_32259,N_28455,N_28800);
nand U32260 (N_32260,N_28334,N_27888);
and U32261 (N_32261,N_27705,N_28868);
or U32262 (N_32262,N_28464,N_28996);
or U32263 (N_32263,N_28211,N_28123);
or U32264 (N_32264,N_27941,N_28048);
nand U32265 (N_32265,N_29397,N_29836);
nor U32266 (N_32266,N_27588,N_27926);
or U32267 (N_32267,N_29776,N_28522);
nand U32268 (N_32268,N_29971,N_28021);
nor U32269 (N_32269,N_29224,N_29968);
nand U32270 (N_32270,N_29113,N_28274);
or U32271 (N_32271,N_28677,N_29760);
and U32272 (N_32272,N_29191,N_29451);
nor U32273 (N_32273,N_29761,N_28465);
nor U32274 (N_32274,N_28773,N_27824);
nor U32275 (N_32275,N_27915,N_27989);
or U32276 (N_32276,N_28739,N_27623);
and U32277 (N_32277,N_28812,N_29634);
nand U32278 (N_32278,N_28736,N_28614);
or U32279 (N_32279,N_29365,N_28928);
and U32280 (N_32280,N_28439,N_27593);
and U32281 (N_32281,N_28584,N_27674);
nand U32282 (N_32282,N_29777,N_28372);
nor U32283 (N_32283,N_29321,N_29717);
nand U32284 (N_32284,N_28557,N_28647);
nor U32285 (N_32285,N_29460,N_29599);
nand U32286 (N_32286,N_29020,N_29651);
or U32287 (N_32287,N_27907,N_29142);
xor U32288 (N_32288,N_29352,N_27631);
nand U32289 (N_32289,N_27946,N_28141);
nand U32290 (N_32290,N_28005,N_29534);
nand U32291 (N_32291,N_29059,N_29734);
or U32292 (N_32292,N_28699,N_29360);
nand U32293 (N_32293,N_28979,N_29435);
nor U32294 (N_32294,N_27574,N_28756);
nor U32295 (N_32295,N_29588,N_27822);
nand U32296 (N_32296,N_28182,N_28080);
nand U32297 (N_32297,N_28465,N_29869);
nor U32298 (N_32298,N_27872,N_28576);
and U32299 (N_32299,N_29383,N_27638);
and U32300 (N_32300,N_29859,N_29231);
xnor U32301 (N_32301,N_27703,N_28569);
nor U32302 (N_32302,N_29452,N_29464);
nor U32303 (N_32303,N_29338,N_29555);
and U32304 (N_32304,N_27984,N_29011);
or U32305 (N_32305,N_29723,N_29645);
xor U32306 (N_32306,N_29804,N_28583);
and U32307 (N_32307,N_29475,N_29686);
nor U32308 (N_32308,N_29846,N_28465);
nor U32309 (N_32309,N_27892,N_29171);
and U32310 (N_32310,N_27746,N_29594);
or U32311 (N_32311,N_27881,N_29385);
xor U32312 (N_32312,N_29019,N_27937);
and U32313 (N_32313,N_29861,N_29184);
and U32314 (N_32314,N_29328,N_28303);
or U32315 (N_32315,N_28084,N_27608);
nand U32316 (N_32316,N_28593,N_28425);
and U32317 (N_32317,N_27925,N_29097);
and U32318 (N_32318,N_28094,N_27804);
and U32319 (N_32319,N_28205,N_29108);
or U32320 (N_32320,N_29982,N_27751);
nand U32321 (N_32321,N_28224,N_28455);
and U32322 (N_32322,N_29654,N_29163);
nand U32323 (N_32323,N_27828,N_27719);
nand U32324 (N_32324,N_28554,N_29586);
and U32325 (N_32325,N_27880,N_27741);
nor U32326 (N_32326,N_29026,N_29039);
nor U32327 (N_32327,N_27642,N_27937);
nand U32328 (N_32328,N_29688,N_29821);
or U32329 (N_32329,N_29286,N_28276);
or U32330 (N_32330,N_28624,N_28850);
nand U32331 (N_32331,N_27596,N_29005);
and U32332 (N_32332,N_29603,N_29372);
and U32333 (N_32333,N_28005,N_28485);
nand U32334 (N_32334,N_28455,N_29044);
nor U32335 (N_32335,N_29155,N_28393);
and U32336 (N_32336,N_28688,N_29811);
or U32337 (N_32337,N_27575,N_27913);
or U32338 (N_32338,N_29372,N_28411);
nor U32339 (N_32339,N_29545,N_28179);
nand U32340 (N_32340,N_28745,N_28489);
nand U32341 (N_32341,N_28791,N_29675);
or U32342 (N_32342,N_28657,N_29804);
nand U32343 (N_32343,N_28991,N_28596);
nand U32344 (N_32344,N_29246,N_27996);
nand U32345 (N_32345,N_28331,N_29910);
nand U32346 (N_32346,N_28873,N_29984);
and U32347 (N_32347,N_28774,N_29291);
or U32348 (N_32348,N_28860,N_28358);
and U32349 (N_32349,N_28992,N_27506);
or U32350 (N_32350,N_28897,N_29921);
nor U32351 (N_32351,N_28233,N_27900);
nor U32352 (N_32352,N_28166,N_27602);
nor U32353 (N_32353,N_28372,N_28916);
nand U32354 (N_32354,N_28897,N_28257);
or U32355 (N_32355,N_29346,N_29516);
nor U32356 (N_32356,N_29339,N_28790);
or U32357 (N_32357,N_28095,N_28560);
or U32358 (N_32358,N_29359,N_28062);
and U32359 (N_32359,N_28818,N_29514);
nand U32360 (N_32360,N_28619,N_28857);
and U32361 (N_32361,N_28988,N_29589);
and U32362 (N_32362,N_27610,N_29579);
nand U32363 (N_32363,N_28829,N_27523);
or U32364 (N_32364,N_28222,N_29416);
nand U32365 (N_32365,N_29466,N_29396);
nor U32366 (N_32366,N_28963,N_28064);
nand U32367 (N_32367,N_29139,N_29935);
nand U32368 (N_32368,N_29477,N_29920);
nor U32369 (N_32369,N_27657,N_29120);
and U32370 (N_32370,N_28500,N_27953);
nor U32371 (N_32371,N_29013,N_28388);
and U32372 (N_32372,N_28042,N_28758);
or U32373 (N_32373,N_28331,N_28929);
or U32374 (N_32374,N_28140,N_29991);
nor U32375 (N_32375,N_29700,N_29707);
and U32376 (N_32376,N_28648,N_29657);
or U32377 (N_32377,N_29264,N_28483);
nor U32378 (N_32378,N_28345,N_29936);
xnor U32379 (N_32379,N_29778,N_28681);
nand U32380 (N_32380,N_28987,N_28766);
and U32381 (N_32381,N_29113,N_29653);
nand U32382 (N_32382,N_29692,N_28576);
and U32383 (N_32383,N_29474,N_28651);
xnor U32384 (N_32384,N_29151,N_27743);
nand U32385 (N_32385,N_28759,N_29674);
and U32386 (N_32386,N_29181,N_29130);
nor U32387 (N_32387,N_27556,N_29855);
nand U32388 (N_32388,N_29454,N_28361);
nor U32389 (N_32389,N_27819,N_29509);
nand U32390 (N_32390,N_28934,N_28669);
nand U32391 (N_32391,N_29963,N_29314);
nor U32392 (N_32392,N_28209,N_28329);
or U32393 (N_32393,N_28941,N_28748);
nor U32394 (N_32394,N_27714,N_28992);
and U32395 (N_32395,N_29882,N_27552);
xor U32396 (N_32396,N_28791,N_29393);
or U32397 (N_32397,N_29076,N_29287);
and U32398 (N_32398,N_29352,N_28024);
and U32399 (N_32399,N_27669,N_28907);
and U32400 (N_32400,N_29506,N_27560);
nor U32401 (N_32401,N_28982,N_29831);
and U32402 (N_32402,N_28959,N_27653);
nand U32403 (N_32403,N_28970,N_28337);
nand U32404 (N_32404,N_29913,N_29207);
nand U32405 (N_32405,N_29660,N_29210);
nor U32406 (N_32406,N_27781,N_28058);
or U32407 (N_32407,N_27947,N_28369);
or U32408 (N_32408,N_29947,N_29946);
and U32409 (N_32409,N_28431,N_28165);
and U32410 (N_32410,N_28877,N_27723);
nor U32411 (N_32411,N_28685,N_29194);
and U32412 (N_32412,N_28067,N_27547);
and U32413 (N_32413,N_29554,N_29459);
nand U32414 (N_32414,N_29152,N_28232);
and U32415 (N_32415,N_27701,N_28900);
and U32416 (N_32416,N_28732,N_27552);
and U32417 (N_32417,N_28420,N_28856);
nand U32418 (N_32418,N_28423,N_28392);
nor U32419 (N_32419,N_28908,N_29953);
and U32420 (N_32420,N_27686,N_29646);
nor U32421 (N_32421,N_27625,N_27773);
or U32422 (N_32422,N_29305,N_29020);
nor U32423 (N_32423,N_27995,N_29244);
nor U32424 (N_32424,N_29847,N_27915);
nand U32425 (N_32425,N_27709,N_29087);
xor U32426 (N_32426,N_28539,N_29971);
nor U32427 (N_32427,N_28117,N_27556);
and U32428 (N_32428,N_28140,N_27625);
and U32429 (N_32429,N_28179,N_28421);
xnor U32430 (N_32430,N_28100,N_28843);
nor U32431 (N_32431,N_28414,N_29032);
nor U32432 (N_32432,N_28190,N_28666);
and U32433 (N_32433,N_29898,N_29408);
and U32434 (N_32434,N_28952,N_28657);
and U32435 (N_32435,N_29835,N_29826);
and U32436 (N_32436,N_29313,N_28710);
or U32437 (N_32437,N_28831,N_28744);
and U32438 (N_32438,N_27917,N_29005);
and U32439 (N_32439,N_28299,N_29156);
nor U32440 (N_32440,N_29215,N_29420);
xnor U32441 (N_32441,N_28984,N_29268);
or U32442 (N_32442,N_27716,N_29869);
nand U32443 (N_32443,N_28906,N_28444);
nand U32444 (N_32444,N_27613,N_28351);
nor U32445 (N_32445,N_28508,N_28432);
nor U32446 (N_32446,N_28889,N_27742);
nor U32447 (N_32447,N_29511,N_29086);
nor U32448 (N_32448,N_28498,N_28643);
xnor U32449 (N_32449,N_29422,N_28267);
nor U32450 (N_32450,N_29577,N_27879);
and U32451 (N_32451,N_29275,N_28616);
or U32452 (N_32452,N_28794,N_29932);
and U32453 (N_32453,N_29419,N_27984);
nor U32454 (N_32454,N_28286,N_27988);
or U32455 (N_32455,N_27541,N_28019);
nand U32456 (N_32456,N_29953,N_27660);
and U32457 (N_32457,N_28783,N_28291);
xnor U32458 (N_32458,N_28321,N_29235);
or U32459 (N_32459,N_28339,N_29223);
xnor U32460 (N_32460,N_27550,N_29818);
or U32461 (N_32461,N_29194,N_29950);
nor U32462 (N_32462,N_29303,N_28526);
nand U32463 (N_32463,N_27855,N_29329);
xnor U32464 (N_32464,N_29698,N_29396);
and U32465 (N_32465,N_28476,N_29715);
or U32466 (N_32466,N_27565,N_28234);
or U32467 (N_32467,N_29025,N_29860);
nor U32468 (N_32468,N_29350,N_27539);
nor U32469 (N_32469,N_29390,N_28733);
xor U32470 (N_32470,N_29791,N_29954);
or U32471 (N_32471,N_28161,N_29489);
nor U32472 (N_32472,N_27527,N_29534);
and U32473 (N_32473,N_28262,N_29146);
or U32474 (N_32474,N_28660,N_28226);
or U32475 (N_32475,N_28174,N_29191);
or U32476 (N_32476,N_28717,N_27766);
nor U32477 (N_32477,N_28998,N_27987);
or U32478 (N_32478,N_29980,N_28170);
nand U32479 (N_32479,N_29850,N_27856);
xor U32480 (N_32480,N_27721,N_29876);
nor U32481 (N_32481,N_28509,N_27941);
or U32482 (N_32482,N_27923,N_28944);
and U32483 (N_32483,N_29133,N_27592);
or U32484 (N_32484,N_28439,N_29884);
or U32485 (N_32485,N_28256,N_28414);
or U32486 (N_32486,N_28383,N_28793);
or U32487 (N_32487,N_29898,N_28107);
or U32488 (N_32488,N_28400,N_29584);
xor U32489 (N_32489,N_29269,N_28629);
and U32490 (N_32490,N_29688,N_28334);
nand U32491 (N_32491,N_28854,N_29292);
xor U32492 (N_32492,N_29160,N_29036);
nand U32493 (N_32493,N_28911,N_28883);
xor U32494 (N_32494,N_28406,N_28397);
and U32495 (N_32495,N_29442,N_27883);
or U32496 (N_32496,N_29314,N_27716);
or U32497 (N_32497,N_29765,N_29641);
nand U32498 (N_32498,N_27767,N_28213);
nor U32499 (N_32499,N_29124,N_28700);
nor U32500 (N_32500,N_32200,N_32072);
nand U32501 (N_32501,N_31602,N_31424);
nand U32502 (N_32502,N_31068,N_32291);
and U32503 (N_32503,N_31684,N_30867);
nor U32504 (N_32504,N_31638,N_31323);
and U32505 (N_32505,N_30789,N_31896);
nor U32506 (N_32506,N_30513,N_30319);
nand U32507 (N_32507,N_30022,N_31038);
nor U32508 (N_32508,N_31186,N_31527);
nand U32509 (N_32509,N_30247,N_32151);
nand U32510 (N_32510,N_32315,N_32280);
or U32511 (N_32511,N_31918,N_30184);
nor U32512 (N_32512,N_30044,N_31506);
nor U32513 (N_32513,N_31137,N_30428);
nor U32514 (N_32514,N_30514,N_30765);
or U32515 (N_32515,N_30379,N_31912);
or U32516 (N_32516,N_30078,N_31787);
or U32517 (N_32517,N_31035,N_31046);
xnor U32518 (N_32518,N_31840,N_30463);
and U32519 (N_32519,N_30502,N_32090);
and U32520 (N_32520,N_31683,N_31389);
nand U32521 (N_32521,N_31198,N_32243);
nand U32522 (N_32522,N_30220,N_31493);
nand U32523 (N_32523,N_30777,N_30903);
nand U32524 (N_32524,N_31436,N_32462);
nor U32525 (N_32525,N_31981,N_30877);
and U32526 (N_32526,N_32460,N_31783);
nor U32527 (N_32527,N_31055,N_32353);
nand U32528 (N_32528,N_31997,N_32437);
or U32529 (N_32529,N_31970,N_31969);
and U32530 (N_32530,N_30511,N_30103);
nor U32531 (N_32531,N_31777,N_30760);
and U32532 (N_32532,N_30161,N_30870);
and U32533 (N_32533,N_30456,N_30941);
and U32534 (N_32534,N_30522,N_32366);
and U32535 (N_32535,N_31722,N_30085);
nor U32536 (N_32536,N_31448,N_30214);
nand U32537 (N_32537,N_31491,N_32050);
or U32538 (N_32538,N_30454,N_30628);
or U32539 (N_32539,N_30614,N_32038);
nand U32540 (N_32540,N_32195,N_31181);
nand U32541 (N_32541,N_30178,N_32154);
nand U32542 (N_32542,N_31397,N_31639);
nor U32543 (N_32543,N_32069,N_30027);
nand U32544 (N_32544,N_30776,N_31362);
nor U32545 (N_32545,N_30238,N_30665);
nand U32546 (N_32546,N_30258,N_31563);
and U32547 (N_32547,N_32428,N_30248);
or U32548 (N_32548,N_31763,N_30586);
or U32549 (N_32549,N_32040,N_32438);
or U32550 (N_32550,N_32492,N_30748);
xor U32551 (N_32551,N_32276,N_31309);
and U32552 (N_32552,N_31614,N_32468);
and U32553 (N_32553,N_31232,N_30151);
or U32554 (N_32554,N_31607,N_32019);
nand U32555 (N_32555,N_31347,N_30501);
nand U32556 (N_32556,N_30858,N_32032);
and U32557 (N_32557,N_31419,N_30003);
nand U32558 (N_32558,N_32237,N_31123);
nor U32559 (N_32559,N_30953,N_32312);
nand U32560 (N_32560,N_32373,N_31313);
and U32561 (N_32561,N_30123,N_30942);
nor U32562 (N_32562,N_31327,N_32397);
nand U32563 (N_32563,N_32281,N_32006);
nand U32564 (N_32564,N_32254,N_31630);
xnor U32565 (N_32565,N_31672,N_30605);
or U32566 (N_32566,N_30599,N_32402);
and U32567 (N_32567,N_32263,N_32126);
and U32568 (N_32568,N_30126,N_30958);
xnor U32569 (N_32569,N_30210,N_32333);
xor U32570 (N_32570,N_30312,N_31950);
and U32571 (N_32571,N_30466,N_31246);
nor U32572 (N_32572,N_32020,N_31132);
xnor U32573 (N_32573,N_31281,N_30965);
or U32574 (N_32574,N_30332,N_31008);
nand U32575 (N_32575,N_31268,N_31119);
nor U32576 (N_32576,N_30250,N_31219);
nor U32577 (N_32577,N_30472,N_31386);
or U32578 (N_32578,N_31533,N_31361);
xnor U32579 (N_32579,N_30730,N_32095);
and U32580 (N_32580,N_30735,N_30913);
nand U32581 (N_32581,N_30716,N_31189);
or U32582 (N_32582,N_30484,N_31465);
and U32583 (N_32583,N_31815,N_31336);
nand U32584 (N_32584,N_30695,N_32235);
and U32585 (N_32585,N_30598,N_32015);
nand U32586 (N_32586,N_31736,N_31501);
or U32587 (N_32587,N_30260,N_31260);
nand U32588 (N_32588,N_31050,N_32433);
nand U32589 (N_32589,N_31959,N_32142);
nor U32590 (N_32590,N_30759,N_30545);
or U32591 (N_32591,N_32357,N_31565);
nand U32592 (N_32592,N_31779,N_30970);
and U32593 (N_32593,N_31377,N_32182);
nand U32594 (N_32594,N_30234,N_32201);
or U32595 (N_32595,N_30441,N_31828);
nor U32596 (N_32596,N_31460,N_32171);
nor U32597 (N_32597,N_31932,N_30021);
or U32598 (N_32598,N_30782,N_31299);
nand U32599 (N_32599,N_31228,N_30120);
nor U32600 (N_32600,N_30621,N_31590);
nand U32601 (N_32601,N_31117,N_31519);
nand U32602 (N_32602,N_31091,N_31234);
nor U32603 (N_32603,N_30311,N_32054);
or U32604 (N_32604,N_31149,N_31171);
and U32605 (N_32605,N_31188,N_30082);
or U32606 (N_32606,N_30711,N_30575);
xnor U32607 (N_32607,N_30807,N_31656);
or U32608 (N_32608,N_30757,N_31223);
nor U32609 (N_32609,N_31028,N_32136);
and U32610 (N_32610,N_31109,N_30920);
or U32611 (N_32611,N_30147,N_31670);
or U32612 (N_32612,N_32396,N_32094);
nand U32613 (N_32613,N_31151,N_31387);
xor U32614 (N_32614,N_31252,N_32239);
or U32615 (N_32615,N_31720,N_31578);
nand U32616 (N_32616,N_30440,N_31306);
and U32617 (N_32617,N_30866,N_31690);
xor U32618 (N_32618,N_30849,N_31699);
nand U32619 (N_32619,N_30774,N_30862);
nand U32620 (N_32620,N_31017,N_30356);
nor U32621 (N_32621,N_32422,N_31985);
or U32622 (N_32622,N_30682,N_30904);
or U32623 (N_32623,N_31741,N_31201);
or U32624 (N_32624,N_30141,N_32056);
nand U32625 (N_32625,N_30833,N_32170);
xnor U32626 (N_32626,N_31834,N_31712);
nand U32627 (N_32627,N_30616,N_32247);
or U32628 (N_32628,N_30015,N_30612);
nand U32629 (N_32629,N_31438,N_30887);
nand U32630 (N_32630,N_30198,N_30232);
nand U32631 (N_32631,N_30462,N_30416);
nand U32632 (N_32632,N_31325,N_32003);
and U32633 (N_32633,N_30421,N_32296);
and U32634 (N_32634,N_31090,N_31818);
and U32635 (N_32635,N_31956,N_32259);
nand U32636 (N_32636,N_31030,N_31660);
and U32637 (N_32637,N_32073,N_31671);
xor U32638 (N_32638,N_31431,N_32068);
or U32639 (N_32639,N_30893,N_30909);
or U32640 (N_32640,N_30381,N_31802);
xnor U32641 (N_32641,N_30772,N_30115);
nor U32642 (N_32642,N_30073,N_30275);
nor U32643 (N_32643,N_30798,N_31958);
nor U32644 (N_32644,N_32447,N_30725);
nand U32645 (N_32645,N_32378,N_31897);
or U32646 (N_32646,N_32481,N_30324);
and U32647 (N_32647,N_30487,N_31618);
nor U32648 (N_32648,N_30281,N_31473);
nor U32649 (N_32649,N_32332,N_31576);
nor U32650 (N_32650,N_30921,N_30876);
nand U32651 (N_32651,N_30063,N_31497);
or U32652 (N_32652,N_31128,N_31014);
nand U32653 (N_32653,N_30802,N_31365);
and U32654 (N_32654,N_30996,N_32217);
xnor U32655 (N_32655,N_31575,N_30938);
nand U32656 (N_32656,N_31946,N_30212);
nand U32657 (N_32657,N_31000,N_30329);
nor U32658 (N_32658,N_31675,N_31271);
and U32659 (N_32659,N_30559,N_32035);
and U32660 (N_32660,N_31928,N_30737);
nor U32661 (N_32661,N_31564,N_30933);
nor U32662 (N_32662,N_31237,N_30295);
and U32663 (N_32663,N_32388,N_30129);
nor U32664 (N_32664,N_32342,N_30578);
or U32665 (N_32665,N_31645,N_31835);
nor U32666 (N_32666,N_32081,N_30345);
nor U32667 (N_32667,N_30592,N_30959);
and U32668 (N_32668,N_31369,N_30786);
and U32669 (N_32669,N_32351,N_32377);
or U32670 (N_32670,N_30203,N_32343);
nand U32671 (N_32671,N_32087,N_31755);
nor U32672 (N_32672,N_32328,N_31865);
nor U32673 (N_32673,N_30733,N_31513);
or U32674 (N_32674,N_31734,N_31713);
or U32675 (N_32675,N_30955,N_31678);
and U32676 (N_32676,N_31303,N_31544);
nand U32677 (N_32677,N_31455,N_32426);
or U32678 (N_32678,N_31374,N_31382);
xnor U32679 (N_32679,N_31087,N_31516);
xnor U32680 (N_32680,N_31425,N_31085);
or U32681 (N_32681,N_31278,N_31013);
and U32682 (N_32682,N_31767,N_30464);
and U32683 (N_32683,N_32246,N_30901);
xnor U32684 (N_32684,N_30678,N_30080);
and U32685 (N_32685,N_30093,N_30179);
nor U32686 (N_32686,N_32309,N_32461);
nor U32687 (N_32687,N_30148,N_30000);
and U32688 (N_32688,N_30417,N_31975);
xnor U32689 (N_32689,N_31284,N_31968);
and U32690 (N_32690,N_32103,N_31941);
or U32691 (N_32691,N_31541,N_30404);
nand U32692 (N_32692,N_30527,N_30927);
or U32693 (N_32693,N_32042,N_30001);
nand U32694 (N_32694,N_31737,N_31852);
and U32695 (N_32695,N_30461,N_32355);
nor U32696 (N_32696,N_32197,N_32029);
nand U32697 (N_32697,N_30626,N_30425);
xor U32698 (N_32698,N_31372,N_31290);
nand U32699 (N_32699,N_31040,N_31923);
or U32700 (N_32700,N_30651,N_31523);
and U32701 (N_32701,N_30071,N_32334);
nand U32702 (N_32702,N_32091,N_30205);
nand U32703 (N_32703,N_30674,N_30564);
and U32704 (N_32704,N_30687,N_32250);
nor U32705 (N_32705,N_32302,N_31937);
xor U32706 (N_32706,N_31052,N_32406);
or U32707 (N_32707,N_31376,N_31832);
xor U32708 (N_32708,N_30305,N_31826);
xnor U32709 (N_32709,N_32215,N_31384);
nand U32710 (N_32710,N_31170,N_30675);
nand U32711 (N_32711,N_31654,N_30851);
nor U32712 (N_32712,N_30335,N_30552);
nand U32713 (N_32713,N_32112,N_31153);
or U32714 (N_32714,N_32016,N_30816);
or U32715 (N_32715,N_30197,N_31514);
or U32716 (N_32716,N_30004,N_31892);
and U32717 (N_32717,N_32297,N_32439);
or U32718 (N_32718,N_30981,N_32004);
nor U32719 (N_32719,N_31502,N_31124);
nand U32720 (N_32720,N_31581,N_32471);
nand U32721 (N_32721,N_31948,N_30821);
and U32722 (N_32722,N_31995,N_31820);
nand U32723 (N_32723,N_30536,N_31939);
nor U32724 (N_32724,N_30768,N_30935);
nor U32725 (N_32725,N_32206,N_32470);
nand U32726 (N_32726,N_31688,N_30011);
or U32727 (N_32727,N_32390,N_31193);
nand U32728 (N_32728,N_30583,N_30283);
or U32729 (N_32729,N_32435,N_30924);
nand U32730 (N_32730,N_30221,N_31164);
nor U32731 (N_32731,N_30029,N_30540);
nor U32732 (N_32732,N_31595,N_30882);
or U32733 (N_32733,N_31215,N_31305);
and U32734 (N_32734,N_31626,N_31803);
or U32735 (N_32735,N_30482,N_31813);
and U32736 (N_32736,N_31543,N_32172);
and U32737 (N_32737,N_30727,N_31531);
and U32738 (N_32738,N_31135,N_31337);
and U32739 (N_32739,N_32371,N_32000);
and U32740 (N_32740,N_30788,N_30244);
nand U32741 (N_32741,N_30330,N_30173);
and U32742 (N_32742,N_30167,N_30715);
and U32743 (N_32743,N_30743,N_31287);
and U32744 (N_32744,N_30287,N_30124);
xor U32745 (N_32745,N_31805,N_31668);
nor U32746 (N_32746,N_32420,N_31343);
nand U32747 (N_32747,N_30369,N_30347);
xor U32748 (N_32748,N_31752,N_30784);
or U32749 (N_32749,N_30274,N_32213);
nor U32750 (N_32750,N_31204,N_30794);
or U32751 (N_32751,N_32132,N_31944);
or U32752 (N_32752,N_30262,N_30191);
nand U32753 (N_32753,N_32374,N_30642);
or U32754 (N_32754,N_31251,N_30321);
or U32755 (N_32755,N_30383,N_31549);
nand U32756 (N_32756,N_30257,N_32381);
nor U32757 (N_32757,N_32146,N_30973);
nand U32758 (N_32758,N_30848,N_31603);
and U32759 (N_32759,N_31742,N_30145);
nor U32760 (N_32760,N_31358,N_31141);
nor U32761 (N_32761,N_30622,N_30714);
and U32762 (N_32762,N_32221,N_31480);
and U32763 (N_32763,N_31854,N_30939);
nand U32764 (N_32764,N_30566,N_31462);
and U32765 (N_32765,N_31872,N_30346);
nor U32766 (N_32766,N_31583,N_31799);
xor U32767 (N_32767,N_31746,N_30518);
or U32768 (N_32768,N_31966,N_30246);
nand U32769 (N_32769,N_30470,N_30493);
nand U32770 (N_32770,N_30864,N_30731);
or U32771 (N_32771,N_30139,N_30850);
nand U32772 (N_32772,N_32293,N_30426);
or U32773 (N_32773,N_30204,N_30652);
and U32774 (N_32774,N_30562,N_30506);
nor U32775 (N_32775,N_32079,N_30698);
or U32776 (N_32776,N_30991,N_30497);
nand U32777 (N_32777,N_32064,N_32419);
nor U32778 (N_32778,N_30028,N_31833);
xor U32779 (N_32779,N_31196,N_31443);
and U32780 (N_32780,N_30138,N_31613);
xor U32781 (N_32781,N_31812,N_30363);
xor U32782 (N_32782,N_30570,N_31391);
nand U32783 (N_32783,N_31875,N_31963);
and U32784 (N_32784,N_32028,N_30684);
xnor U32785 (N_32785,N_31096,N_31029);
nand U32786 (N_32786,N_31836,N_30932);
nand U32787 (N_32787,N_30677,N_31640);
nor U32788 (N_32788,N_30127,N_30433);
nand U32789 (N_32789,N_31267,N_30524);
nor U32790 (N_32790,N_31914,N_30136);
nor U32791 (N_32791,N_30300,N_31240);
nor U32792 (N_32792,N_30199,N_31866);
xnor U32793 (N_32793,N_31871,N_31316);
and U32794 (N_32794,N_32036,N_30606);
nor U32795 (N_32795,N_31609,N_31167);
nor U32796 (N_32796,N_30106,N_31441);
or U32797 (N_32797,N_31230,N_31134);
nand U32798 (N_32798,N_31274,N_31743);
nor U32799 (N_32799,N_30801,N_31723);
or U32800 (N_32800,N_32034,N_31483);
nand U32801 (N_32801,N_31778,N_30081);
nand U32802 (N_32802,N_30696,N_31573);
and U32803 (N_32803,N_31711,N_30193);
nor U32804 (N_32804,N_31718,N_30888);
and U32805 (N_32805,N_31403,N_31445);
or U32806 (N_32806,N_31587,N_31469);
or U32807 (N_32807,N_32025,N_32314);
and U32808 (N_32808,N_30307,N_30704);
and U32809 (N_32809,N_31423,N_31676);
and U32810 (N_32810,N_31227,N_30945);
nor U32811 (N_32811,N_30646,N_30961);
or U32812 (N_32812,N_31404,N_32260);
or U32813 (N_32813,N_31520,N_30783);
and U32814 (N_32814,N_30722,N_31851);
and U32815 (N_32815,N_32441,N_31457);
nor U32816 (N_32816,N_30393,N_32156);
nand U32817 (N_32817,N_31398,N_31036);
nor U32818 (N_32818,N_30243,N_30133);
and U32819 (N_32819,N_32349,N_30899);
or U32820 (N_32820,N_32454,N_30742);
nand U32821 (N_32821,N_31144,N_30037);
or U32822 (N_32822,N_31115,N_32498);
or U32823 (N_32823,N_30846,N_31666);
and U32824 (N_32824,N_31857,N_31916);
or U32825 (N_32825,N_30349,N_31704);
nand U32826 (N_32826,N_30019,N_32191);
and U32827 (N_32827,N_30405,N_30668);
nand U32828 (N_32828,N_31716,N_31118);
and U32829 (N_32829,N_32078,N_32053);
and U32830 (N_32830,N_30038,N_30091);
nand U32831 (N_32831,N_30892,N_31293);
nand U32832 (N_32832,N_31474,N_30940);
or U32833 (N_32833,N_30581,N_31371);
or U32834 (N_32834,N_31827,N_31102);
nand U32835 (N_32835,N_31558,N_32337);
and U32836 (N_32836,N_30089,N_30611);
and U32837 (N_32837,N_31070,N_30597);
nor U32838 (N_32838,N_30676,N_32340);
nor U32839 (N_32839,N_31314,N_32128);
or U32840 (N_32840,N_30620,N_32173);
or U32841 (N_32841,N_32188,N_30496);
and U32842 (N_32842,N_30439,N_30800);
nor U32843 (N_32843,N_32356,N_32354);
nor U32844 (N_32844,N_31951,N_31121);
nand U32845 (N_32845,N_31468,N_30617);
and U32846 (N_32846,N_32131,N_31194);
nand U32847 (N_32847,N_32076,N_30042);
nor U32848 (N_32848,N_30432,N_30529);
or U32849 (N_32849,N_31360,N_31733);
nand U32850 (N_32850,N_30658,N_31911);
nand U32851 (N_32851,N_31136,N_30568);
or U32852 (N_32852,N_30012,N_31789);
and U32853 (N_32853,N_32062,N_32089);
and U32854 (N_32854,N_31147,N_30697);
nor U32855 (N_32855,N_31582,N_30930);
or U32856 (N_32856,N_31632,N_30014);
nor U32857 (N_32857,N_31453,N_31208);
and U32858 (N_32858,N_30006,N_30931);
and U32859 (N_32859,N_30749,N_30934);
or U32860 (N_32860,N_31127,N_30579);
nor U32861 (N_32861,N_31620,N_31600);
nand U32862 (N_32862,N_32024,N_31884);
or U32863 (N_32863,N_31021,N_31524);
or U32864 (N_32864,N_30070,N_32185);
xor U32865 (N_32865,N_30431,N_31681);
nand U32866 (N_32866,N_30724,N_32486);
and U32867 (N_32867,N_30160,N_30686);
nand U32868 (N_32868,N_30631,N_32127);
nand U32869 (N_32869,N_30539,N_32379);
nand U32870 (N_32870,N_31992,N_31988);
nor U32871 (N_32871,N_32408,N_31172);
nand U32872 (N_32872,N_30710,N_31971);
nor U32873 (N_32873,N_30072,N_31781);
nor U32874 (N_32874,N_31550,N_31103);
xnor U32875 (N_32875,N_32140,N_32484);
nand U32876 (N_32876,N_31224,N_30845);
and U32877 (N_32877,N_31760,N_32262);
and U32878 (N_32878,N_31929,N_31610);
or U32879 (N_32879,N_31870,N_30902);
nand U32880 (N_32880,N_31798,N_32412);
nand U32881 (N_32881,N_30008,N_30131);
and U32882 (N_32882,N_30637,N_32469);
xor U32883 (N_32883,N_32229,N_30744);
nand U32884 (N_32884,N_32018,N_30897);
or U32885 (N_32885,N_32096,N_30746);
or U32886 (N_32886,N_31098,N_31659);
nor U32887 (N_32887,N_31526,N_31867);
nand U32888 (N_32888,N_30976,N_31579);
nor U32889 (N_32889,N_31811,N_31308);
and U32890 (N_32890,N_30031,N_32008);
nand U32891 (N_32891,N_30033,N_32395);
nor U32892 (N_32892,N_31176,N_30299);
or U32893 (N_32893,N_30298,N_30251);
nor U32894 (N_32894,N_30092,N_30956);
nand U32895 (N_32895,N_30364,N_31726);
nor U32896 (N_32896,N_30526,N_31146);
and U32897 (N_32897,N_30812,N_32212);
nand U32898 (N_32898,N_30256,N_30608);
nand U32899 (N_32899,N_31059,N_31965);
nand U32900 (N_32900,N_30105,N_31079);
nand U32901 (N_32901,N_30362,N_32456);
or U32902 (N_32902,N_30987,N_30130);
and U32903 (N_32903,N_31764,N_32306);
and U32904 (N_32904,N_31795,N_30587);
or U32905 (N_32905,N_30806,N_32181);
nor U32906 (N_32906,N_30672,N_31860);
xor U32907 (N_32907,N_31433,N_31221);
nor U32908 (N_32908,N_31326,N_30825);
or U32909 (N_32909,N_30692,N_31275);
and U32910 (N_32910,N_32101,N_30435);
and U32911 (N_32911,N_30679,N_30745);
nor U32912 (N_32912,N_30708,N_30860);
and U32913 (N_32913,N_31285,N_31288);
or U32914 (N_32914,N_32049,N_30781);
nand U32915 (N_32915,N_31508,N_30555);
or U32916 (N_32916,N_32478,N_32288);
and U32917 (N_32917,N_31140,N_30448);
nor U32918 (N_32918,N_30153,N_31740);
or U32919 (N_32919,N_30169,N_30842);
or U32920 (N_32920,N_31589,N_31922);
or U32921 (N_32921,N_32031,N_32123);
or U32922 (N_32922,N_31310,N_31381);
and U32923 (N_32923,N_30271,N_30810);
nor U32924 (N_32924,N_31105,N_31301);
and U32925 (N_32925,N_31001,N_31191);
nand U32926 (N_32926,N_30367,N_32279);
nor U32927 (N_32927,N_30861,N_32178);
or U32928 (N_32928,N_31168,N_30325);
nand U32929 (N_32929,N_31318,N_31031);
or U32930 (N_32930,N_30998,N_31364);
nor U32931 (N_32931,N_30360,N_31321);
and U32932 (N_32932,N_32483,N_30847);
nand U32933 (N_32933,N_32234,N_30828);
nor U32934 (N_32934,N_30521,N_31955);
or U32935 (N_32935,N_30655,N_31804);
or U32936 (N_32936,N_31496,N_30331);
nand U32937 (N_32937,N_30074,N_30202);
nor U32938 (N_32938,N_30490,N_30310);
and U32939 (N_32939,N_30398,N_31470);
and U32940 (N_32940,N_30334,N_30891);
nor U32941 (N_32941,N_30712,N_31300);
nand U32942 (N_32942,N_32467,N_31463);
xnor U32943 (N_32943,N_31529,N_32167);
and U32944 (N_32944,N_31915,N_30154);
nand U32945 (N_32945,N_31138,N_31745);
and U32946 (N_32946,N_30728,N_30430);
or U32947 (N_32947,N_32219,N_30185);
nor U32948 (N_32948,N_31159,N_32488);
nand U32949 (N_32949,N_31207,N_32313);
or U32950 (N_32950,N_32386,N_31270);
or U32951 (N_32951,N_31466,N_31253);
nor U32952 (N_32952,N_32199,N_30445);
xor U32953 (N_32953,N_32046,N_30064);
and U32954 (N_32954,N_31071,N_30832);
nand U32955 (N_32955,N_30415,N_30403);
nor U32956 (N_32956,N_32252,N_31706);
and U32957 (N_32957,N_30503,N_31330);
nor U32958 (N_32958,N_31572,N_30101);
nor U32959 (N_32959,N_31155,N_31003);
nor U32960 (N_32960,N_30457,N_31165);
nand U32961 (N_32961,N_31351,N_31476);
nor U32962 (N_32962,N_31856,N_31701);
and U32963 (N_32963,N_30297,N_31503);
xor U32964 (N_32964,N_32137,N_31909);
nor U32965 (N_32965,N_30495,N_30799);
nor U32966 (N_32966,N_32256,N_32100);
xor U32967 (N_32967,N_32176,N_30055);
xnor U32968 (N_32968,N_31107,N_30424);
nor U32969 (N_32969,N_31846,N_30766);
or U32970 (N_32970,N_30750,N_31843);
or U32971 (N_32971,N_31673,N_32407);
xnor U32972 (N_32972,N_30485,N_30067);
xor U32973 (N_32973,N_31642,N_31788);
and U32974 (N_32974,N_31749,N_31202);
or U32975 (N_32975,N_30572,N_30925);
nor U32976 (N_32976,N_30420,N_31636);
nand U32977 (N_32977,N_30165,N_30437);
or U32978 (N_32978,N_30778,N_32310);
and U32979 (N_32979,N_32232,N_31027);
xnor U32980 (N_32980,N_32230,N_31719);
and U32981 (N_32981,N_31751,N_30928);
nor U32982 (N_32982,N_32060,N_32013);
nand U32983 (N_32983,N_31294,N_32113);
nand U32984 (N_32984,N_31150,N_31577);
nand U32985 (N_32985,N_31414,N_31877);
nor U32986 (N_32986,N_30112,N_31821);
or U32987 (N_32987,N_31489,N_31819);
or U32988 (N_32988,N_31899,N_31131);
xor U32989 (N_32989,N_30168,N_31408);
and U32990 (N_32990,N_31823,N_30320);
and U32991 (N_32991,N_31346,N_32475);
and U32992 (N_32992,N_31368,N_30183);
or U32993 (N_32993,N_32301,N_31487);
nor U32994 (N_32994,N_30779,N_31509);
or U32995 (N_32995,N_30787,N_31890);
nor U32996 (N_32996,N_31032,N_31903);
or U32997 (N_32997,N_31461,N_31498);
nor U32998 (N_32998,N_31080,N_30670);
and U32999 (N_32999,N_31005,N_30336);
nor U33000 (N_33000,N_31195,N_30831);
nand U33001 (N_33001,N_32319,N_32166);
nand U33002 (N_33002,N_30459,N_30289);
and U33003 (N_33003,N_32411,N_31822);
nor U33004 (N_33004,N_32347,N_30609);
nand U33005 (N_33005,N_31717,N_31900);
and U33006 (N_33006,N_30792,N_31212);
and U33007 (N_33007,N_31435,N_31794);
nand U33008 (N_33008,N_31979,N_31947);
xnor U33009 (N_33009,N_31551,N_32465);
and U33010 (N_33010,N_30556,N_30150);
or U33011 (N_33011,N_32214,N_31904);
nand U33012 (N_33012,N_31101,N_31536);
nor U33013 (N_33013,N_31366,N_30914);
nand U33014 (N_33014,N_31383,N_31009);
and U33015 (N_33015,N_32352,N_30738);
xor U33016 (N_33016,N_31905,N_31731);
xor U33017 (N_33017,N_31927,N_30411);
nor U33018 (N_33018,N_32086,N_30255);
and U33019 (N_33019,N_31616,N_32216);
nor U33020 (N_33020,N_31824,N_31456);
and U33021 (N_33021,N_30446,N_31729);
xor U33022 (N_33022,N_30837,N_32318);
or U33023 (N_33023,N_31738,N_32300);
or U33024 (N_33024,N_30318,N_31604);
or U33025 (N_33025,N_31652,N_30900);
and U33026 (N_33026,N_32344,N_30465);
nand U33027 (N_33027,N_32289,N_30290);
nand U33028 (N_33028,N_30100,N_30666);
xor U33029 (N_33029,N_32331,N_30873);
nand U33030 (N_33030,N_30650,N_31385);
and U33031 (N_33031,N_31883,N_30943);
and U33032 (N_33032,N_31292,N_30264);
nand U33033 (N_33033,N_30689,N_31845);
or U33034 (N_33034,N_30230,N_31593);
nor U33035 (N_33035,N_30280,N_30580);
nor U33036 (N_33036,N_30990,N_31108);
nand U33037 (N_33037,N_30875,N_30211);
and U33038 (N_33038,N_32434,N_30648);
nor U33039 (N_33039,N_32414,N_30844);
and U33040 (N_33040,N_30829,N_30315);
or U33041 (N_33041,N_31559,N_31505);
nand U33042 (N_33042,N_31791,N_30390);
or U33043 (N_33043,N_30795,N_31961);
or U33044 (N_33044,N_31236,N_31169);
xor U33045 (N_33045,N_30690,N_32322);
nor U33046 (N_33046,N_31409,N_31214);
nor U33047 (N_33047,N_32294,N_31047);
nor U33048 (N_33048,N_31211,N_30890);
nor U33049 (N_33049,N_30240,N_31444);
nand U33050 (N_33050,N_31279,N_30159);
and U33051 (N_33051,N_30149,N_31881);
and U33052 (N_33052,N_30296,N_30673);
xor U33053 (N_33053,N_30016,N_30507);
nand U33054 (N_33054,N_31554,N_30929);
and U33055 (N_33055,N_30039,N_31104);
nor U33056 (N_33056,N_31319,N_31721);
nand U33057 (N_33057,N_31154,N_30217);
nand U33058 (N_33058,N_31174,N_30375);
nor U33059 (N_33059,N_32376,N_30979);
or U33060 (N_33060,N_31679,N_31682);
and U33061 (N_33061,N_31507,N_31410);
and U33062 (N_33062,N_31627,N_31472);
nand U33063 (N_33063,N_30543,N_31247);
or U33064 (N_33064,N_32403,N_31982);
nor U33065 (N_33065,N_31567,N_30333);
nand U33066 (N_33066,N_31769,N_32149);
nand U33067 (N_33067,N_31143,N_31901);
nor U33068 (N_33068,N_31065,N_32385);
and U33069 (N_33069,N_30654,N_30102);
nor U33070 (N_33070,N_30434,N_30239);
nand U33071 (N_33071,N_30563,N_32431);
or U33072 (N_33072,N_30879,N_32320);
or U33073 (N_33073,N_32299,N_31855);
xnor U33074 (N_33074,N_31847,N_30999);
and U33075 (N_33075,N_30116,N_30357);
or U33076 (N_33076,N_32104,N_31077);
nand U33077 (N_33077,N_30739,N_31210);
and U33078 (N_33078,N_30685,N_31621);
nand U33079 (N_33079,N_32159,N_30371);
nor U33080 (N_33080,N_30041,N_32277);
and U33081 (N_33081,N_31333,N_31762);
nand U33082 (N_33082,N_30259,N_30249);
nor U33083 (N_33083,N_32175,N_31060);
xor U33084 (N_33084,N_30734,N_31691);
nor U33085 (N_33085,N_30499,N_30468);
xor U33086 (N_33086,N_32490,N_30964);
nand U33087 (N_33087,N_30024,N_32043);
or U33088 (N_33088,N_30550,N_32324);
nand U33089 (N_33089,N_30986,N_32359);
nand U33090 (N_33090,N_32361,N_32122);
and U33091 (N_33091,N_32233,N_30627);
nand U33092 (N_33092,N_31999,N_31917);
nor U33093 (N_33093,N_32241,N_30721);
and U33094 (N_33094,N_32440,N_31488);
nand U33095 (N_33095,N_30368,N_30076);
or U33096 (N_33096,N_30661,N_30773);
nand U33097 (N_33097,N_31588,N_30479);
and U33098 (N_33098,N_31148,N_30822);
nand U33099 (N_33099,N_30741,N_31283);
or U33100 (N_33100,N_32463,N_31315);
or U33101 (N_33101,N_30740,N_32098);
nand U33102 (N_33102,N_31882,N_32161);
nor U33103 (N_33103,N_32202,N_31667);
and U33104 (N_33104,N_31611,N_32047);
nor U33105 (N_33105,N_31353,N_30060);
or U33106 (N_33106,N_31317,N_32265);
or U33107 (N_33107,N_30010,N_31933);
nand U33108 (N_33108,N_30498,N_30549);
and U33109 (N_33109,N_30302,N_32144);
nand U33110 (N_33110,N_30868,N_30163);
or U33111 (N_33111,N_31429,N_30649);
and U33112 (N_33112,N_31166,N_32455);
and U33113 (N_33113,N_30206,N_32417);
and U33114 (N_33114,N_30767,N_30128);
or U33115 (N_33115,N_30056,N_30277);
or U33116 (N_33116,N_30265,N_31597);
nand U33117 (N_33117,N_32245,N_31838);
nor U33118 (N_33118,N_30337,N_30201);
nor U33119 (N_33119,N_31532,N_31859);
xnor U33120 (N_33120,N_30489,N_30050);
or U33121 (N_33121,N_32399,N_31139);
and U33122 (N_33122,N_30922,N_30699);
nor U33123 (N_33123,N_31095,N_31535);
xnor U33124 (N_33124,N_32066,N_31924);
xnor U33125 (N_33125,N_32092,N_30591);
nand U33126 (N_33126,N_30156,N_31048);
or U33127 (N_33127,N_31413,N_32135);
nand U33128 (N_33128,N_30374,N_31266);
or U33129 (N_33129,N_30896,N_30057);
and U33130 (N_33130,N_31585,N_32187);
and U33131 (N_33131,N_32041,N_30835);
nand U33132 (N_33132,N_31698,N_30190);
xor U33133 (N_33133,N_30576,N_31390);
and U33134 (N_33134,N_31510,N_32039);
nand U33135 (N_33135,N_30088,N_30585);
and U33136 (N_33136,N_30408,N_30820);
nor U33137 (N_33137,N_30808,N_31669);
or U33138 (N_33138,N_30378,N_30702);
xor U33139 (N_33139,N_31991,N_32152);
or U33140 (N_33140,N_32278,N_32400);
nor U33141 (N_33141,N_30451,N_30515);
and U33142 (N_33142,N_30036,N_31853);
and U33143 (N_33143,N_31156,N_30372);
or U33144 (N_33144,N_30984,N_30442);
or U33145 (N_33145,N_31727,N_30803);
or U33146 (N_33146,N_32453,N_30162);
nand U33147 (N_33147,N_32269,N_30110);
and U33148 (N_33148,N_30219,N_30595);
nand U33149 (N_33149,N_31229,N_30397);
nor U33150 (N_33150,N_31686,N_31580);
and U33151 (N_33151,N_31797,N_31296);
or U33152 (N_33152,N_30978,N_32238);
xor U33153 (N_33153,N_32147,N_31484);
xor U33154 (N_33154,N_30736,N_31786);
nand U33155 (N_33155,N_31254,N_30342);
nor U33156 (N_33156,N_31873,N_31495);
and U33157 (N_33157,N_31311,N_31687);
or U33158 (N_33158,N_31482,N_32346);
or U33159 (N_33159,N_32295,N_31930);
nor U33160 (N_33160,N_31657,N_31935);
and U33161 (N_33161,N_31225,N_30269);
and U33162 (N_33162,N_30355,N_31863);
xnor U33163 (N_33163,N_30977,N_32075);
and U33164 (N_33164,N_31412,N_30883);
nor U33165 (N_33165,N_30948,N_32111);
xor U33166 (N_33166,N_31714,N_31428);
or U33167 (N_33167,N_30134,N_31710);
and U33168 (N_33168,N_32327,N_32286);
or U33169 (N_33169,N_32317,N_30636);
nor U33170 (N_33170,N_32114,N_30632);
xnor U33171 (N_33171,N_30359,N_31399);
xor U33172 (N_33172,N_30284,N_30796);
nor U33173 (N_33173,N_31486,N_30152);
nor U33174 (N_33174,N_30122,N_30213);
or U33175 (N_33175,N_32208,N_30032);
nor U33176 (N_33176,N_31192,N_30603);
nand U33177 (N_33177,N_32336,N_32223);
nor U33178 (N_33178,N_32077,N_31477);
xnor U33179 (N_33179,N_31257,N_31018);
nand U33180 (N_33180,N_30365,N_31735);
nand U33181 (N_33181,N_32134,N_30483);
nand U33182 (N_33182,N_30653,N_30993);
nor U33183 (N_33183,N_31571,N_32421);
or U33184 (N_33184,N_31338,N_32458);
nand U33185 (N_33185,N_31990,N_32474);
or U33186 (N_33186,N_32443,N_30815);
nand U33187 (N_33187,N_31878,N_31297);
xor U33188 (N_33188,N_31076,N_31530);
and U33189 (N_33189,N_32168,N_31471);
nand U33190 (N_33190,N_31850,N_30252);
nand U33191 (N_33191,N_30533,N_32473);
xnor U33192 (N_33192,N_31931,N_31983);
and U33193 (N_33193,N_31183,N_32052);
nand U33194 (N_33194,N_31635,N_31481);
or U33195 (N_33195,N_31747,N_30528);
and U33196 (N_33196,N_32393,N_32255);
nor U33197 (N_33197,N_32364,N_31392);
and U33198 (N_33198,N_32249,N_31907);
nor U33199 (N_33199,N_32416,N_31622);
nor U33200 (N_33200,N_32404,N_32097);
or U33201 (N_33201,N_31887,N_30554);
nand U33202 (N_33202,N_30640,N_30775);
nor U33203 (N_33203,N_31099,N_31072);
nor U33204 (N_33204,N_32192,N_30601);
nand U33205 (N_33205,N_30481,N_30293);
nor U33206 (N_33206,N_32198,N_31647);
nor U33207 (N_33207,N_30664,N_30657);
nor U33208 (N_33208,N_31596,N_32496);
xor U33209 (N_33209,N_30659,N_30361);
xnor U33210 (N_33210,N_30557,N_32472);
and U33211 (N_33211,N_31058,N_30035);
and U33212 (N_33212,N_31898,N_32445);
and U33213 (N_33213,N_31708,N_30351);
or U33214 (N_33214,N_31891,N_30048);
or U33215 (N_33215,N_32099,N_30177);
and U33216 (N_33216,N_30962,N_30582);
or U33217 (N_33217,N_31500,N_31421);
xor U33218 (N_33218,N_31357,N_31396);
and U33219 (N_33219,N_30309,N_32164);
nor U33220 (N_33220,N_30223,N_31973);
or U33221 (N_33221,N_31010,N_31940);
nor U33222 (N_33222,N_30558,N_30826);
nor U33223 (N_33223,N_31653,N_30957);
or U33224 (N_33224,N_31161,N_31242);
nor U33225 (N_33225,N_30253,N_30994);
nor U33226 (N_33226,N_31092,N_31025);
and U33227 (N_33227,N_31960,N_30969);
xor U33228 (N_33228,N_31816,N_30532);
nor U33229 (N_33229,N_31644,N_32345);
or U33230 (N_33230,N_31039,N_30017);
nand U33231 (N_33231,N_31938,N_30771);
nand U33232 (N_33232,N_31231,N_32011);
and U33233 (N_33233,N_30317,N_31546);
nor U33234 (N_33234,N_32367,N_30805);
nand U33235 (N_33235,N_32466,N_31440);
nand U33236 (N_33236,N_31542,N_31920);
or U33237 (N_33237,N_30195,N_31015);
and U33238 (N_33238,N_30625,N_32117);
nand U33239 (N_33239,N_31034,N_30713);
or U33240 (N_33240,N_30841,N_32372);
nor U33241 (N_33241,N_31776,N_31839);
and U33242 (N_33242,N_30376,N_32449);
nor U33243 (N_33243,N_30273,N_30705);
nor U33244 (N_33244,N_32368,N_30394);
or U33245 (N_33245,N_30449,N_30607);
or U33246 (N_33246,N_32027,N_31379);
nor U33247 (N_33247,N_30752,N_31693);
nand U33248 (N_33248,N_30874,N_30377);
or U33249 (N_33249,N_31265,N_30971);
or U33250 (N_33250,N_31954,N_30937);
and U33251 (N_33251,N_31272,N_31407);
nor U33252 (N_33252,N_31049,N_32358);
and U33253 (N_33253,N_32105,N_30588);
and U33254 (N_33254,N_30980,N_32326);
and U33255 (N_33255,N_31395,N_31163);
and U33256 (N_33256,N_31753,N_31561);
or U33257 (N_33257,N_30797,N_30700);
or U33258 (N_33258,N_30517,N_31641);
nor U33259 (N_33259,N_31088,N_31261);
nand U33260 (N_33260,N_31750,N_30989);
nand U33261 (N_33261,N_31598,N_32348);
nor U33262 (N_33262,N_31646,N_31044);
nand U33263 (N_33263,N_32258,N_30002);
nor U33264 (N_33264,N_30303,N_31538);
or U33265 (N_33265,N_32284,N_31926);
or U33266 (N_33266,N_30043,N_31792);
nand U33267 (N_33267,N_31051,N_31370);
or U33268 (N_33268,N_30030,N_31348);
or U33269 (N_33269,N_31511,N_30083);
and U33270 (N_33270,N_30228,N_31250);
and U33271 (N_33271,N_32329,N_30146);
nor U33272 (N_33272,N_31876,N_30188);
nand U33273 (N_33273,N_31492,N_30898);
or U33274 (N_33274,N_31175,N_32055);
and U33275 (N_33275,N_31548,N_30751);
and U33276 (N_33276,N_31817,N_32093);
nand U33277 (N_33277,N_30551,N_30117);
and U33278 (N_33278,N_30669,N_32163);
and U33279 (N_33279,N_31499,N_32325);
and U33280 (N_33280,N_30753,N_31053);
nor U33281 (N_33281,N_31993,N_31262);
nand U33282 (N_33282,N_30094,N_30096);
nand U33283 (N_33283,N_30018,N_30143);
nand U33284 (N_33284,N_30282,N_31744);
or U33285 (N_33285,N_30755,N_32457);
or U33286 (N_33286,N_31724,N_31352);
or U33287 (N_33287,N_31574,N_31125);
nor U33288 (N_33288,N_31774,N_32160);
or U33289 (N_33289,N_30401,N_30200);
nor U33290 (N_33290,N_31355,N_30843);
or U33291 (N_33291,N_30859,N_32248);
xor U33292 (N_33292,N_30869,N_31634);
nor U33293 (N_33293,N_31962,N_32120);
nand U33294 (N_33294,N_30473,N_30504);
and U33295 (N_33295,N_31113,N_31619);
or U33296 (N_33296,N_32387,N_31402);
nor U33297 (N_33297,N_30406,N_31280);
nor U33298 (N_33298,N_30460,N_31631);
xnor U33299 (N_33299,N_32451,N_32001);
and U33300 (N_33300,N_30171,N_32063);
and U33301 (N_33301,N_32065,N_30639);
nor U33302 (N_33302,N_31556,N_32021);
nand U33303 (N_33303,N_32067,N_30791);
nor U33304 (N_33304,N_31213,N_30350);
or U33305 (N_33305,N_30052,N_31393);
nand U33306 (N_33306,N_31158,N_31793);
and U33307 (N_33307,N_30429,N_30066);
nor U33308 (N_33308,N_30471,N_30121);
and U33309 (N_33309,N_30509,N_32209);
or U33310 (N_33310,N_30453,N_30099);
nand U33311 (N_33311,N_31073,N_31083);
nor U33312 (N_33312,N_30619,N_32218);
or U33313 (N_33313,N_30985,N_30491);
xor U33314 (N_33314,N_31235,N_32145);
nand U33315 (N_33315,N_30380,N_31322);
nand U33316 (N_33316,N_32222,N_32133);
nand U33317 (N_33317,N_32023,N_32082);
and U33318 (N_33318,N_30339,N_32158);
nand U33319 (N_33319,N_32316,N_31152);
or U33320 (N_33320,N_30291,N_32186);
nand U33321 (N_33321,N_31986,N_30720);
or U33322 (N_33322,N_32010,N_30109);
nor U33323 (N_33323,N_30013,N_32303);
xnor U33324 (N_33324,N_30316,N_30571);
or U33325 (N_33325,N_32177,N_32125);
nor U33326 (N_33326,N_31528,N_31515);
nand U33327 (N_33327,N_31697,N_31332);
and U33328 (N_33328,N_31324,N_32138);
nand U33329 (N_33329,N_31002,N_30158);
nand U33330 (N_33330,N_31298,N_30602);
nor U33331 (N_33331,N_32184,N_32189);
xnor U33332 (N_33332,N_30075,N_31592);
nor U33333 (N_33333,N_30754,N_31081);
nor U33334 (N_33334,N_32143,N_32391);
nand U33335 (N_33335,N_32257,N_30387);
nor U33336 (N_33336,N_30967,N_30344);
or U33337 (N_33337,N_31785,N_31540);
nand U33338 (N_33338,N_31606,N_30327);
xnor U33339 (N_33339,N_30553,N_31608);
nand U33340 (N_33340,N_30407,N_31570);
and U33341 (N_33341,N_31952,N_32383);
and U33342 (N_33342,N_30905,N_30354);
nand U33343 (N_33343,N_30049,N_30726);
or U33344 (N_33344,N_30189,N_32489);
or U33345 (N_33345,N_31662,N_30412);
xor U33346 (N_33346,N_32476,N_32494);
or U33347 (N_33347,N_31004,N_30992);
nand U33348 (N_33348,N_31187,N_32026);
or U33349 (N_33349,N_30386,N_32264);
nor U33350 (N_33350,N_31972,N_31605);
or U33351 (N_33351,N_30908,N_31800);
or U33352 (N_33352,N_31043,N_32491);
nand U33353 (N_33353,N_31807,N_30438);
nor U33354 (N_33354,N_30569,N_30288);
nand U33355 (N_33355,N_30995,N_30104);
nand U33356 (N_33356,N_30233,N_31555);
and U33357 (N_33357,N_31459,N_30155);
nand U33358 (N_33358,N_31354,N_30227);
nor U33359 (N_33359,N_32446,N_31977);
nand U33360 (N_33360,N_32285,N_30077);
and U33361 (N_33361,N_31525,N_32225);
and U33362 (N_33362,N_32074,N_32401);
nor U33363 (N_33363,N_30594,N_30034);
nand U33364 (N_33364,N_32030,N_30338);
nor U33365 (N_33365,N_31451,N_30758);
xnor U33366 (N_33366,N_30975,N_30391);
nor U33367 (N_33367,N_32150,N_32014);
or U33368 (N_33368,N_30756,N_30192);
nor U33369 (N_33369,N_31075,N_30196);
xnor U33370 (N_33370,N_32058,N_31730);
nand U33371 (N_33371,N_30618,N_30906);
nor U33372 (N_33372,N_30061,N_30747);
nand U33373 (N_33373,N_31566,N_30340);
or U33374 (N_33374,N_32009,N_31702);
nor U33375 (N_33375,N_31624,N_31485);
nand U33376 (N_33376,N_31184,N_32362);
and U33377 (N_33377,N_30894,N_32179);
nor U33378 (N_33378,N_30414,N_31715);
nand U33379 (N_33379,N_31913,N_30194);
nor U33380 (N_33380,N_30172,N_30486);
and U33381 (N_33381,N_31648,N_30561);
nor U33382 (N_33382,N_31022,N_31732);
and U33383 (N_33383,N_32339,N_30308);
or U33384 (N_33384,N_30884,N_31766);
or U33385 (N_33385,N_30423,N_31910);
and U33386 (N_33386,N_32290,N_30137);
nor U33387 (N_33387,N_30254,N_31356);
and U33388 (N_33388,N_31868,N_30589);
nor U33389 (N_33389,N_32141,N_31069);
nand U33390 (N_33390,N_32017,N_30936);
and U33391 (N_33391,N_32061,N_31655);
and U33392 (N_33392,N_30187,N_31378);
and U33393 (N_33393,N_31380,N_32242);
or U33394 (N_33394,N_30114,N_31637);
nor U33395 (N_33395,N_31016,N_31061);
nor U33396 (N_33396,N_31949,N_31562);
and U33397 (N_33397,N_31199,N_30285);
nor U33398 (N_33398,N_30634,N_30025);
or U33399 (N_33399,N_31844,N_31394);
nand U33400 (N_33400,N_32118,N_32287);
and U33401 (N_33401,N_32244,N_30764);
and U33402 (N_33402,N_30400,N_31238);
or U33403 (N_33403,N_30040,N_31490);
nor U33404 (N_33404,N_32380,N_32330);
nand U33405 (N_33405,N_30836,N_30638);
nor U33406 (N_33406,N_31919,N_30476);
nor U33407 (N_33407,N_31056,N_31661);
nand U33408 (N_33408,N_30494,N_32305);
and U33409 (N_33409,N_32227,N_31373);
or U33410 (N_33410,N_31895,N_30671);
or U33411 (N_33411,N_31367,N_30348);
nor U33412 (N_33412,N_31906,N_31801);
and U33413 (N_33413,N_31943,N_31458);
and U33414 (N_33414,N_31967,N_31097);
or U33415 (N_33415,N_30709,N_32477);
nor U33416 (N_33416,N_30630,N_31200);
nand U33417 (N_33417,N_30729,N_32119);
and U33418 (N_33418,N_30790,N_30087);
or U33419 (N_33419,N_30079,N_30680);
or U33420 (N_33420,N_31422,N_32005);
or U33421 (N_33421,N_30814,N_31978);
nand U33422 (N_33422,N_31651,N_30447);
nand U33423 (N_33423,N_31757,N_31276);
and U33424 (N_33424,N_30827,N_30236);
nand U33425 (N_33425,N_30343,N_30098);
xnor U33426 (N_33426,N_30216,N_30097);
nand U33427 (N_33427,N_31831,N_31584);
nor U33428 (N_33428,N_31849,N_30118);
or U33429 (N_33429,N_31244,N_30604);
and U33430 (N_33430,N_31674,N_31291);
xnor U33431 (N_33431,N_31705,N_30523);
nor U33432 (N_33432,N_31114,N_31569);
and U33433 (N_33433,N_30395,N_32190);
nor U33434 (N_33434,N_32338,N_30278);
and U33435 (N_33435,N_30313,N_30301);
nor U33436 (N_33436,N_31335,N_31130);
nor U33437 (N_33437,N_31226,N_31934);
xnor U33438 (N_33438,N_31837,N_30144);
nand U33439 (N_33439,N_30306,N_30918);
nor U33440 (N_33440,N_31007,N_30525);
xor U33441 (N_33441,N_31420,N_31885);
or U33442 (N_33442,N_31886,N_31206);
or U33443 (N_33443,N_30629,N_30950);
or U33444 (N_33444,N_32169,N_32282);
nor U33445 (N_33445,N_30174,N_31825);
or U33446 (N_33446,N_30974,N_31725);
and U33447 (N_33447,N_30926,N_30886);
and U33448 (N_33448,N_30422,N_31464);
or U33449 (N_33449,N_32444,N_31259);
and U33450 (N_33450,N_30853,N_31539);
nand U33451 (N_33451,N_32211,N_30688);
nand U33452 (N_33452,N_30656,N_32124);
xnor U33453 (N_33453,N_30450,N_30023);
and U33454 (N_33454,N_32253,N_30681);
xor U33455 (N_33455,N_30694,N_32193);
nor U33456 (N_33456,N_30341,N_31331);
and U33457 (N_33457,N_31594,N_32044);
nand U33458 (N_33458,N_31964,N_31078);
nor U33459 (N_33459,N_32442,N_30500);
nand U33460 (N_33460,N_31880,N_31633);
nand U33461 (N_33461,N_30181,N_30142);
or U33462 (N_33462,N_30209,N_32273);
nand U33463 (N_33463,N_32485,N_30531);
nor U33464 (N_33464,N_31249,N_32180);
nor U33465 (N_33465,N_31829,N_32405);
nor U33466 (N_33466,N_30402,N_32430);
nand U33467 (N_33467,N_31782,N_31342);
and U33468 (N_33468,N_32012,N_30548);
or U33469 (N_33469,N_32071,N_30005);
or U33470 (N_33470,N_30488,N_31177);
and U33471 (N_33471,N_31696,N_30577);
and U33472 (N_33472,N_31100,N_31808);
or U33473 (N_33473,N_30399,N_30322);
xor U33474 (N_33474,N_30157,N_30567);
nor U33475 (N_33475,N_30600,N_32059);
and U33476 (N_33476,N_32382,N_32107);
or U33477 (N_33477,N_30610,N_32384);
or U33478 (N_33478,N_31765,N_31302);
and U33479 (N_33479,N_30095,N_30263);
and U33480 (N_33480,N_31442,N_31334);
nand U33481 (N_33481,N_30058,N_30267);
and U33482 (N_33482,N_31248,N_31976);
nor U33483 (N_33483,N_30270,N_32499);
and U33484 (N_33484,N_31263,N_32084);
and U33485 (N_33485,N_32240,N_30384);
nor U33486 (N_33486,N_30917,N_32196);
or U33487 (N_33487,N_30857,N_31568);
or U33488 (N_33488,N_31989,N_30427);
and U33489 (N_33489,N_32418,N_30852);
or U33490 (N_33490,N_30225,N_30009);
or U33491 (N_33491,N_30966,N_30769);
or U33492 (N_33492,N_31806,N_30910);
nor U33493 (N_33493,N_32370,N_30780);
nand U33494 (N_33494,N_30701,N_31994);
nand U33495 (N_33495,N_31612,N_30125);
and U33496 (N_33496,N_30762,N_30065);
nor U33497 (N_33497,N_31980,N_31110);
xor U33498 (N_33498,N_30108,N_31479);
and U33499 (N_33499,N_32308,N_30051);
and U33500 (N_33500,N_32464,N_32495);
nand U33501 (N_33501,N_32261,N_32033);
xor U33502 (N_33502,N_31289,N_32110);
or U33503 (N_33503,N_32432,N_30323);
and U33504 (N_33504,N_32236,N_30276);
nand U33505 (N_33505,N_30516,N_30419);
nand U33506 (N_33506,N_31649,N_30045);
xor U33507 (N_33507,N_30180,N_31145);
nand U33508 (N_33508,N_30132,N_30723);
or U33509 (N_33509,N_30294,N_31416);
nor U33510 (N_33510,N_30389,N_31925);
and U33511 (N_33511,N_31478,N_30916);
and U33512 (N_33512,N_32392,N_31350);
and U33513 (N_33513,N_32413,N_32283);
nor U33514 (N_33514,N_30455,N_30838);
and U33515 (N_33515,N_30467,N_30912);
and U33516 (N_33516,N_32394,N_30855);
xnor U33517 (N_33517,N_30111,N_30809);
and U33518 (N_33518,N_31830,N_31434);
nand U33519 (N_33519,N_31756,N_30215);
and U33520 (N_33520,N_31809,N_30624);
or U33521 (N_33521,N_31328,N_32363);
and U33522 (N_33522,N_31771,N_32109);
nand U33523 (N_33523,N_30068,N_32002);
nor U33524 (N_33524,N_31344,N_31677);
nand U33525 (N_33525,N_31475,N_32231);
nor U33526 (N_33526,N_32450,N_31012);
and U33527 (N_33527,N_31277,N_31245);
nor U33528 (N_33528,N_31106,N_30328);
or U33529 (N_33529,N_30268,N_30565);
nand U33530 (N_33530,N_32341,N_31133);
nor U33531 (N_33531,N_31658,N_32048);
xnor U33532 (N_33532,N_30761,N_31185);
and U33533 (N_33533,N_31197,N_30410);
nand U33534 (N_33534,N_30053,N_31264);
or U33535 (N_33535,N_30830,N_31045);
and U33536 (N_33536,N_32070,N_30046);
nor U33537 (N_33537,N_30373,N_32121);
nor U33538 (N_33538,N_30972,N_30633);
nand U33539 (N_33539,N_31157,N_30519);
and U33540 (N_33540,N_31447,N_30613);
nor U33541 (N_33541,N_32272,N_31586);
or U33542 (N_33542,N_32224,N_31282);
or U33543 (N_33543,N_30480,N_30647);
nor U33544 (N_33544,N_31233,N_32116);
nor U33545 (N_33545,N_30719,N_31178);
nor U33546 (N_33546,N_30535,N_30542);
and U33547 (N_33547,N_32425,N_31874);
nor U33548 (N_33548,N_30660,N_30615);
or U33549 (N_33549,N_31748,N_31273);
nor U33550 (N_33550,N_30541,N_30880);
nor U33551 (N_33551,N_30895,N_31057);
nor U33552 (N_33552,N_30413,N_30218);
nor U33553 (N_33553,N_31841,N_30889);
or U33554 (N_33554,N_31216,N_31758);
nor U33555 (N_33555,N_31112,N_32080);
nor U33556 (N_33556,N_30706,N_31220);
nand U33557 (N_33557,N_31093,N_31996);
nand U33558 (N_33558,N_30683,N_31066);
nor U33559 (N_33559,N_30878,N_31773);
nand U33560 (N_33560,N_31663,N_30988);
nor U33561 (N_33561,N_31615,N_31430);
and U33562 (N_33562,N_32153,N_30635);
or U33563 (N_33563,N_32497,N_30436);
or U33564 (N_33564,N_31650,N_30643);
xnor U33565 (N_33565,N_30949,N_30915);
xor U33566 (N_33566,N_31494,N_31450);
or U33567 (N_33567,N_32375,N_31142);
and U33568 (N_33568,N_31862,N_30823);
nand U33569 (N_33569,N_30396,N_32452);
nand U33570 (N_33570,N_31908,N_30007);
xor U33571 (N_33571,N_31452,N_32174);
nor U33572 (N_33572,N_31426,N_31415);
or U33573 (N_33573,N_30475,N_31709);
or U33574 (N_33574,N_31796,N_31728);
and U33575 (N_33575,N_31120,N_32088);
xor U33576 (N_33576,N_32335,N_31401);
and U33577 (N_33577,N_30353,N_31341);
or U33578 (N_33578,N_31388,N_31218);
nand U33579 (N_33579,N_30596,N_30286);
nand U33580 (N_33580,N_30547,N_32108);
nor U33581 (N_33581,N_31084,N_31547);
or U33582 (N_33582,N_31534,N_31754);
nor U33583 (N_33583,N_30119,N_30245);
and U33584 (N_33584,N_31617,N_31902);
nor U33585 (N_33585,N_31557,N_30919);
and U33586 (N_33586,N_30366,N_30944);
or U33587 (N_33587,N_32228,N_31241);
and U33588 (N_33588,N_32251,N_31848);
or U33589 (N_33589,N_30785,N_30663);
or U33590 (N_33590,N_31623,N_30458);
nor U33591 (N_33591,N_30644,N_30314);
nor U33592 (N_33592,N_32323,N_31790);
nor U33593 (N_33593,N_31162,N_30952);
xor U33594 (N_33594,N_30590,N_30140);
nor U33595 (N_33595,N_30242,N_31063);
xor U33596 (N_33596,N_30793,N_31094);
or U33597 (N_33597,N_30084,N_30304);
nor U33598 (N_33598,N_31089,N_31439);
xnor U33599 (N_33599,N_30231,N_31775);
and U33600 (N_33600,N_30175,N_31984);
and U33601 (N_33601,N_31942,N_32051);
and U33602 (N_33602,N_31116,N_30272);
nor U33603 (N_33603,N_32037,N_32083);
nor U33604 (N_33604,N_32268,N_30443);
or U33605 (N_33605,N_31217,N_30865);
and U33606 (N_33606,N_30505,N_31255);
nor U33607 (N_33607,N_30718,N_30069);
nor U33608 (N_33608,N_31329,N_31375);
xnor U33609 (N_33609,N_30090,N_30047);
xnor U33610 (N_33610,N_31814,N_32480);
and U33611 (N_33611,N_31418,N_30834);
xor U33612 (N_33612,N_32203,N_32007);
nand U33613 (N_33613,N_30279,N_32226);
and U33614 (N_33614,N_30584,N_31953);
nor U33615 (N_33615,N_32220,N_31205);
nand U33616 (N_33616,N_31518,N_31180);
nor U33617 (N_33617,N_30261,N_30770);
or U33618 (N_33618,N_31861,N_30054);
and U33619 (N_33619,N_31643,N_30534);
nor U33620 (N_33620,N_31768,N_31400);
and U33621 (N_33621,N_31256,N_30352);
and U33622 (N_33622,N_30520,N_30241);
xor U33623 (N_33623,N_32487,N_31692);
and U33624 (N_33624,N_31694,N_30020);
xor U33625 (N_33625,N_32106,N_31179);
and U33626 (N_33626,N_31062,N_32115);
nand U33627 (N_33627,N_31869,N_30732);
nor U33628 (N_33628,N_30418,N_31067);
nor U33629 (N_33629,N_31888,N_31894);
and U33630 (N_33630,N_32270,N_30623);
and U33631 (N_33631,N_30546,N_31449);
nor U33632 (N_33632,N_32398,N_30818);
or U33633 (N_33633,N_31041,N_32365);
or U33634 (N_33634,N_30854,N_30946);
nand U33635 (N_33635,N_30947,N_31552);
nor U33636 (N_33636,N_30982,N_30824);
nand U33637 (N_33637,N_30186,N_31243);
nand U33638 (N_33638,N_31664,N_31553);
or U33639 (N_33639,N_31054,N_30813);
and U33640 (N_33640,N_30871,N_32194);
and U33641 (N_33641,N_30222,N_30226);
and U33642 (N_33642,N_32267,N_31082);
nor U33643 (N_33643,N_30292,N_31680);
nand U33644 (N_33644,N_30452,N_30817);
xnor U33645 (N_33645,N_30804,N_30530);
or U33646 (N_33646,N_31599,N_30409);
and U33647 (N_33647,N_31417,N_31628);
and U33648 (N_33648,N_32045,N_31560);
nand U33649 (N_33649,N_30538,N_32204);
and U33650 (N_33650,N_30811,N_32448);
and U33651 (N_33651,N_32205,N_30478);
or U33652 (N_33652,N_31889,N_31998);
nand U33653 (N_33653,N_30182,N_31893);
nand U33654 (N_33654,N_30963,N_30382);
nor U33655 (N_33655,N_32369,N_31405);
or U33656 (N_33656,N_31020,N_30856);
or U33657 (N_33657,N_30326,N_31784);
nand U33658 (N_33658,N_31312,N_31437);
nand U33659 (N_33659,N_32130,N_32307);
and U33660 (N_33660,N_32129,N_31239);
nor U33661 (N_33661,N_31601,N_30107);
and U33662 (N_33662,N_31340,N_30358);
nor U33663 (N_33663,N_31629,N_32162);
and U33664 (N_33664,N_31665,N_31359);
nor U33665 (N_33665,N_31454,N_32424);
and U33666 (N_33666,N_30537,N_31160);
or U33667 (N_33667,N_30164,N_31307);
nand U33668 (N_33668,N_31987,N_30881);
and U33669 (N_33669,N_30983,N_31695);
nor U33670 (N_33670,N_30667,N_31411);
nor U33671 (N_33671,N_31545,N_30229);
and U33672 (N_33672,N_30385,N_31945);
nor U33673 (N_33673,N_31304,N_30763);
nor U33674 (N_33674,N_30997,N_31772);
or U33675 (N_33675,N_30968,N_30208);
nor U33676 (N_33676,N_31446,N_32057);
nand U33677 (N_33677,N_31625,N_32479);
nor U33678 (N_33678,N_32423,N_32292);
or U33679 (N_33679,N_32165,N_31086);
nor U33680 (N_33680,N_31759,N_30266);
and U33681 (N_33681,N_30224,N_32155);
nand U33682 (N_33682,N_31521,N_30176);
xor U33683 (N_33683,N_32304,N_32311);
nand U33684 (N_33684,N_31345,N_32409);
nand U33685 (N_33685,N_31770,N_30923);
or U33686 (N_33686,N_30885,N_31703);
or U33687 (N_33687,N_31258,N_30717);
nor U33688 (N_33688,N_31006,N_31203);
and U33689 (N_33689,N_31182,N_30707);
nand U33690 (N_33690,N_30872,N_31111);
and U33691 (N_33691,N_31363,N_31190);
and U33692 (N_33692,N_31936,N_30510);
and U33693 (N_33693,N_30059,N_30086);
and U33694 (N_33694,N_32207,N_30474);
or U33695 (N_33695,N_32459,N_31537);
nor U33696 (N_33696,N_30508,N_31467);
or U33697 (N_33697,N_30573,N_32183);
nor U33698 (N_33698,N_30207,N_30560);
and U33699 (N_33699,N_30544,N_30370);
nand U33700 (N_33700,N_32274,N_31427);
nand U33701 (N_33701,N_31064,N_31074);
xnor U33702 (N_33702,N_31286,N_31023);
nor U33703 (N_33703,N_31512,N_32493);
nor U33704 (N_33704,N_32139,N_30469);
and U33705 (N_33705,N_31026,N_30492);
nor U33706 (N_33706,N_30839,N_30237);
or U33707 (N_33707,N_32482,N_31858);
and U33708 (N_33708,N_31129,N_30235);
nor U33709 (N_33709,N_31504,N_32350);
nand U33710 (N_33710,N_32360,N_31810);
nand U33711 (N_33711,N_30135,N_30911);
or U33712 (N_33712,N_30593,N_31209);
xnor U33713 (N_33713,N_30863,N_30951);
xor U33714 (N_33714,N_30444,N_31320);
or U33715 (N_33715,N_31339,N_32022);
and U33716 (N_33716,N_31864,N_31522);
or U33717 (N_33717,N_31406,N_31295);
nor U33718 (N_33718,N_31222,N_32102);
and U33719 (N_33719,N_31432,N_31019);
and U33720 (N_33720,N_32436,N_32321);
nand U33721 (N_33721,N_30512,N_32298);
xor U33722 (N_33722,N_30840,N_31879);
nand U33723 (N_33723,N_31780,N_30907);
or U33724 (N_33724,N_32210,N_31739);
or U33725 (N_33725,N_30170,N_31517);
nand U33726 (N_33726,N_31173,N_30703);
or U33727 (N_33727,N_32415,N_31974);
nand U33728 (N_33728,N_30691,N_30113);
nor U33729 (N_33729,N_30392,N_31126);
and U33730 (N_33730,N_32157,N_30645);
and U33731 (N_33731,N_31957,N_31033);
xnor U33732 (N_33732,N_32429,N_30641);
or U33733 (N_33733,N_30062,N_31122);
nor U33734 (N_33734,N_32266,N_31761);
and U33735 (N_33735,N_30574,N_30693);
or U33736 (N_33736,N_31921,N_30026);
and U33737 (N_33737,N_31842,N_32085);
nor U33738 (N_33738,N_30388,N_30960);
and U33739 (N_33739,N_31037,N_31685);
xor U33740 (N_33740,N_32148,N_30662);
xor U33741 (N_33741,N_31011,N_30954);
and U33742 (N_33742,N_32275,N_32410);
or U33743 (N_33743,N_31024,N_31700);
nor U33744 (N_33744,N_32427,N_31591);
nor U33745 (N_33745,N_30819,N_31349);
or U33746 (N_33746,N_30166,N_31042);
nor U33747 (N_33747,N_30477,N_32389);
and U33748 (N_33748,N_31707,N_31689);
and U33749 (N_33749,N_31269,N_32271);
xnor U33750 (N_33750,N_31584,N_30218);
nor U33751 (N_33751,N_30861,N_31535);
nand U33752 (N_33752,N_31688,N_32198);
or U33753 (N_33753,N_31240,N_30602);
and U33754 (N_33754,N_30437,N_31342);
and U33755 (N_33755,N_32087,N_31817);
and U33756 (N_33756,N_31471,N_31744);
nor U33757 (N_33757,N_30124,N_31391);
xor U33758 (N_33758,N_30930,N_30378);
nand U33759 (N_33759,N_32410,N_31999);
and U33760 (N_33760,N_31667,N_31178);
and U33761 (N_33761,N_31507,N_30276);
nand U33762 (N_33762,N_31897,N_30497);
nor U33763 (N_33763,N_31660,N_31588);
nand U33764 (N_33764,N_31093,N_30510);
nor U33765 (N_33765,N_30271,N_30240);
and U33766 (N_33766,N_30005,N_31843);
nand U33767 (N_33767,N_30272,N_31037);
nor U33768 (N_33768,N_32236,N_31710);
nor U33769 (N_33769,N_31553,N_30061);
nor U33770 (N_33770,N_31925,N_31943);
and U33771 (N_33771,N_32090,N_31125);
nand U33772 (N_33772,N_32316,N_32229);
xor U33773 (N_33773,N_31868,N_31524);
nand U33774 (N_33774,N_32348,N_31008);
xnor U33775 (N_33775,N_31173,N_30193);
or U33776 (N_33776,N_31911,N_30225);
and U33777 (N_33777,N_31694,N_31286);
nor U33778 (N_33778,N_31317,N_30893);
and U33779 (N_33779,N_30783,N_31613);
and U33780 (N_33780,N_31549,N_30867);
nor U33781 (N_33781,N_32237,N_30332);
nand U33782 (N_33782,N_30177,N_30656);
xnor U33783 (N_33783,N_32491,N_30377);
and U33784 (N_33784,N_30305,N_30763);
or U33785 (N_33785,N_31210,N_30060);
nand U33786 (N_33786,N_32424,N_31317);
nor U33787 (N_33787,N_32454,N_30783);
nand U33788 (N_33788,N_30620,N_31923);
or U33789 (N_33789,N_30069,N_32312);
nand U33790 (N_33790,N_30392,N_31566);
nor U33791 (N_33791,N_31346,N_30643);
or U33792 (N_33792,N_30407,N_30191);
xor U33793 (N_33793,N_31418,N_30827);
and U33794 (N_33794,N_30888,N_30461);
nor U33795 (N_33795,N_32090,N_31487);
or U33796 (N_33796,N_30121,N_30032);
and U33797 (N_33797,N_31444,N_30890);
nand U33798 (N_33798,N_30393,N_31372);
nor U33799 (N_33799,N_31002,N_31921);
and U33800 (N_33800,N_30195,N_30493);
nand U33801 (N_33801,N_31403,N_32387);
and U33802 (N_33802,N_30367,N_30710);
and U33803 (N_33803,N_31408,N_30692);
and U33804 (N_33804,N_32192,N_32386);
xnor U33805 (N_33805,N_32430,N_30660);
or U33806 (N_33806,N_31990,N_32269);
nor U33807 (N_33807,N_32422,N_30150);
or U33808 (N_33808,N_30087,N_30386);
nand U33809 (N_33809,N_32303,N_30650);
nor U33810 (N_33810,N_30254,N_32400);
or U33811 (N_33811,N_31169,N_30920);
nand U33812 (N_33812,N_32353,N_31757);
xor U33813 (N_33813,N_30604,N_30136);
and U33814 (N_33814,N_30463,N_32157);
nor U33815 (N_33815,N_31804,N_32251);
or U33816 (N_33816,N_30141,N_30218);
and U33817 (N_33817,N_31037,N_31448);
nand U33818 (N_33818,N_31948,N_32421);
nand U33819 (N_33819,N_30628,N_31364);
and U33820 (N_33820,N_30453,N_32055);
nand U33821 (N_33821,N_30418,N_31634);
nand U33822 (N_33822,N_32314,N_30210);
nand U33823 (N_33823,N_31762,N_32289);
and U33824 (N_33824,N_30906,N_31661);
or U33825 (N_33825,N_31792,N_30686);
nor U33826 (N_33826,N_31105,N_32449);
nor U33827 (N_33827,N_31825,N_32284);
nor U33828 (N_33828,N_30872,N_32013);
nor U33829 (N_33829,N_32095,N_31300);
nor U33830 (N_33830,N_31139,N_31355);
xor U33831 (N_33831,N_31386,N_31004);
xnor U33832 (N_33832,N_31739,N_32361);
and U33833 (N_33833,N_32221,N_31086);
nor U33834 (N_33834,N_30361,N_32052);
nand U33835 (N_33835,N_32178,N_31507);
nor U33836 (N_33836,N_32052,N_31728);
and U33837 (N_33837,N_31520,N_32243);
nor U33838 (N_33838,N_30662,N_31975);
or U33839 (N_33839,N_31874,N_32160);
nor U33840 (N_33840,N_30160,N_31524);
xor U33841 (N_33841,N_32411,N_30902);
nand U33842 (N_33842,N_30980,N_30717);
or U33843 (N_33843,N_31458,N_32409);
nor U33844 (N_33844,N_31014,N_30634);
or U33845 (N_33845,N_30892,N_32277);
nor U33846 (N_33846,N_30325,N_31031);
or U33847 (N_33847,N_31164,N_31561);
and U33848 (N_33848,N_32473,N_31895);
nand U33849 (N_33849,N_30725,N_32017);
nor U33850 (N_33850,N_31986,N_31188);
nand U33851 (N_33851,N_31832,N_31597);
nand U33852 (N_33852,N_32483,N_31876);
or U33853 (N_33853,N_31474,N_32012);
or U33854 (N_33854,N_31149,N_30543);
or U33855 (N_33855,N_30745,N_31429);
nor U33856 (N_33856,N_30895,N_31726);
nor U33857 (N_33857,N_31684,N_30322);
or U33858 (N_33858,N_32051,N_31227);
xnor U33859 (N_33859,N_30484,N_30246);
or U33860 (N_33860,N_30069,N_31742);
nand U33861 (N_33861,N_31790,N_30272);
and U33862 (N_33862,N_31636,N_32043);
and U33863 (N_33863,N_30416,N_30738);
nand U33864 (N_33864,N_30447,N_32437);
or U33865 (N_33865,N_31594,N_30908);
or U33866 (N_33866,N_31473,N_31837);
nand U33867 (N_33867,N_31432,N_30494);
and U33868 (N_33868,N_31003,N_31992);
or U33869 (N_33869,N_31403,N_30524);
and U33870 (N_33870,N_31242,N_30986);
nand U33871 (N_33871,N_31418,N_31780);
or U33872 (N_33872,N_31279,N_32445);
nand U33873 (N_33873,N_30377,N_31944);
nand U33874 (N_33874,N_31918,N_31394);
nor U33875 (N_33875,N_32186,N_31562);
nor U33876 (N_33876,N_30982,N_31148);
and U33877 (N_33877,N_31139,N_31828);
xnor U33878 (N_33878,N_30862,N_31857);
or U33879 (N_33879,N_30126,N_32070);
or U33880 (N_33880,N_30748,N_32456);
nand U33881 (N_33881,N_30128,N_30290);
or U33882 (N_33882,N_31094,N_32480);
xor U33883 (N_33883,N_31276,N_32308);
nand U33884 (N_33884,N_30854,N_31948);
xor U33885 (N_33885,N_32035,N_31868);
and U33886 (N_33886,N_30118,N_30741);
nor U33887 (N_33887,N_30256,N_31925);
or U33888 (N_33888,N_31541,N_31544);
or U33889 (N_33889,N_31483,N_31280);
and U33890 (N_33890,N_32353,N_30895);
nand U33891 (N_33891,N_31727,N_31386);
or U33892 (N_33892,N_30911,N_30442);
nand U33893 (N_33893,N_32389,N_30518);
and U33894 (N_33894,N_30516,N_31891);
and U33895 (N_33895,N_31718,N_31842);
or U33896 (N_33896,N_30842,N_30370);
nor U33897 (N_33897,N_32313,N_31999);
and U33898 (N_33898,N_32205,N_31466);
nor U33899 (N_33899,N_30176,N_31889);
and U33900 (N_33900,N_31144,N_32149);
or U33901 (N_33901,N_30972,N_31194);
xnor U33902 (N_33902,N_30697,N_31518);
and U33903 (N_33903,N_31856,N_31097);
or U33904 (N_33904,N_31548,N_30202);
nor U33905 (N_33905,N_30165,N_31188);
or U33906 (N_33906,N_31531,N_30443);
or U33907 (N_33907,N_30384,N_31438);
and U33908 (N_33908,N_30515,N_30165);
xor U33909 (N_33909,N_31489,N_31507);
xnor U33910 (N_33910,N_30841,N_32359);
and U33911 (N_33911,N_31501,N_30341);
and U33912 (N_33912,N_31761,N_30401);
nand U33913 (N_33913,N_30325,N_31106);
nand U33914 (N_33914,N_30707,N_32297);
or U33915 (N_33915,N_30495,N_30599);
nor U33916 (N_33916,N_30144,N_30286);
and U33917 (N_33917,N_30320,N_31565);
nor U33918 (N_33918,N_31388,N_30874);
or U33919 (N_33919,N_31163,N_31070);
and U33920 (N_33920,N_30086,N_30886);
or U33921 (N_33921,N_31913,N_30657);
xnor U33922 (N_33922,N_31878,N_30185);
or U33923 (N_33923,N_31634,N_30484);
xnor U33924 (N_33924,N_31110,N_32225);
nand U33925 (N_33925,N_30724,N_30548);
nand U33926 (N_33926,N_30428,N_31379);
and U33927 (N_33927,N_32290,N_31149);
or U33928 (N_33928,N_31469,N_31329);
nand U33929 (N_33929,N_31725,N_31878);
and U33930 (N_33930,N_31484,N_30816);
nand U33931 (N_33931,N_31441,N_30386);
nor U33932 (N_33932,N_30976,N_30708);
nor U33933 (N_33933,N_32222,N_30195);
nor U33934 (N_33934,N_30400,N_30946);
nand U33935 (N_33935,N_32402,N_32396);
nand U33936 (N_33936,N_31981,N_31224);
and U33937 (N_33937,N_30301,N_32175);
nor U33938 (N_33938,N_32137,N_32337);
and U33939 (N_33939,N_31909,N_31227);
and U33940 (N_33940,N_30533,N_31332);
and U33941 (N_33941,N_31360,N_32447);
nor U33942 (N_33942,N_31244,N_31169);
or U33943 (N_33943,N_31748,N_31650);
nand U33944 (N_33944,N_30837,N_30962);
nor U33945 (N_33945,N_31385,N_30648);
xor U33946 (N_33946,N_32431,N_30740);
xnor U33947 (N_33947,N_30098,N_31451);
nor U33948 (N_33948,N_32276,N_31598);
and U33949 (N_33949,N_30265,N_30412);
or U33950 (N_33950,N_30034,N_32028);
nor U33951 (N_33951,N_31952,N_31706);
and U33952 (N_33952,N_32358,N_31306);
xor U33953 (N_33953,N_31581,N_31704);
and U33954 (N_33954,N_32068,N_31224);
nand U33955 (N_33955,N_32371,N_31833);
or U33956 (N_33956,N_31056,N_30991);
or U33957 (N_33957,N_30668,N_31995);
or U33958 (N_33958,N_31309,N_32005);
nand U33959 (N_33959,N_31401,N_31428);
nor U33960 (N_33960,N_32495,N_30489);
or U33961 (N_33961,N_31842,N_32350);
and U33962 (N_33962,N_32429,N_31650);
nand U33963 (N_33963,N_32013,N_31146);
nor U33964 (N_33964,N_32221,N_30548);
or U33965 (N_33965,N_31382,N_30082);
or U33966 (N_33966,N_32069,N_31974);
nand U33967 (N_33967,N_30124,N_30165);
nand U33968 (N_33968,N_30444,N_30701);
and U33969 (N_33969,N_31398,N_32346);
nand U33970 (N_33970,N_31764,N_32054);
and U33971 (N_33971,N_31267,N_30183);
and U33972 (N_33972,N_32112,N_31818);
xor U33973 (N_33973,N_32307,N_31030);
and U33974 (N_33974,N_30930,N_31993);
nor U33975 (N_33975,N_30170,N_30489);
and U33976 (N_33976,N_30300,N_31622);
or U33977 (N_33977,N_30026,N_30958);
nor U33978 (N_33978,N_30733,N_31891);
nor U33979 (N_33979,N_30310,N_31876);
nand U33980 (N_33980,N_30088,N_32493);
nor U33981 (N_33981,N_31005,N_31394);
xor U33982 (N_33982,N_30549,N_31536);
xor U33983 (N_33983,N_31132,N_32085);
and U33984 (N_33984,N_32159,N_31689);
nor U33985 (N_33985,N_30938,N_32145);
and U33986 (N_33986,N_32162,N_30572);
nor U33987 (N_33987,N_30270,N_31758);
nor U33988 (N_33988,N_31452,N_31334);
xnor U33989 (N_33989,N_31044,N_32480);
nor U33990 (N_33990,N_31199,N_31637);
xor U33991 (N_33991,N_32009,N_31871);
or U33992 (N_33992,N_31470,N_30484);
or U33993 (N_33993,N_32219,N_31752);
xor U33994 (N_33994,N_31597,N_30999);
nand U33995 (N_33995,N_31889,N_30793);
and U33996 (N_33996,N_30645,N_31687);
or U33997 (N_33997,N_31541,N_32473);
and U33998 (N_33998,N_30671,N_30275);
nor U33999 (N_33999,N_31391,N_32060);
or U34000 (N_34000,N_31677,N_30079);
or U34001 (N_34001,N_31737,N_32163);
nand U34002 (N_34002,N_31535,N_31353);
or U34003 (N_34003,N_32245,N_31339);
nand U34004 (N_34004,N_31733,N_32336);
nand U34005 (N_34005,N_30941,N_30870);
nand U34006 (N_34006,N_30604,N_30534);
and U34007 (N_34007,N_32260,N_32032);
nand U34008 (N_34008,N_30880,N_30784);
or U34009 (N_34009,N_30745,N_31966);
nor U34010 (N_34010,N_31668,N_30690);
or U34011 (N_34011,N_31549,N_31001);
and U34012 (N_34012,N_30013,N_32004);
or U34013 (N_34013,N_30694,N_30408);
and U34014 (N_34014,N_30101,N_31659);
nand U34015 (N_34015,N_30926,N_31277);
and U34016 (N_34016,N_30589,N_31799);
nor U34017 (N_34017,N_30271,N_32237);
nor U34018 (N_34018,N_31251,N_30154);
and U34019 (N_34019,N_30034,N_30788);
or U34020 (N_34020,N_32036,N_32264);
or U34021 (N_34021,N_31084,N_31770);
or U34022 (N_34022,N_31818,N_31417);
and U34023 (N_34023,N_31872,N_32169);
or U34024 (N_34024,N_31449,N_31208);
nand U34025 (N_34025,N_30622,N_30557);
nor U34026 (N_34026,N_31836,N_32081);
nand U34027 (N_34027,N_30015,N_31596);
xnor U34028 (N_34028,N_31077,N_30158);
xnor U34029 (N_34029,N_32109,N_31469);
nand U34030 (N_34030,N_30105,N_31846);
and U34031 (N_34031,N_30493,N_32008);
nor U34032 (N_34032,N_31707,N_32470);
and U34033 (N_34033,N_30119,N_30669);
or U34034 (N_34034,N_31458,N_31059);
or U34035 (N_34035,N_31935,N_31464);
nand U34036 (N_34036,N_32322,N_31801);
nor U34037 (N_34037,N_31228,N_32499);
and U34038 (N_34038,N_30781,N_30633);
xor U34039 (N_34039,N_30765,N_32480);
and U34040 (N_34040,N_31192,N_30383);
nand U34041 (N_34041,N_31646,N_30952);
nor U34042 (N_34042,N_30046,N_31028);
or U34043 (N_34043,N_31862,N_31202);
xor U34044 (N_34044,N_30371,N_32378);
and U34045 (N_34045,N_32419,N_31261);
and U34046 (N_34046,N_30208,N_30847);
and U34047 (N_34047,N_31302,N_30367);
nor U34048 (N_34048,N_32231,N_31058);
nor U34049 (N_34049,N_31096,N_30616);
nor U34050 (N_34050,N_30582,N_31001);
and U34051 (N_34051,N_30416,N_32357);
nand U34052 (N_34052,N_32218,N_30530);
nand U34053 (N_34053,N_31736,N_32371);
nand U34054 (N_34054,N_30945,N_31411);
nand U34055 (N_34055,N_31835,N_30534);
and U34056 (N_34056,N_30261,N_30439);
or U34057 (N_34057,N_30786,N_32361);
or U34058 (N_34058,N_30249,N_31042);
nor U34059 (N_34059,N_31251,N_32380);
or U34060 (N_34060,N_31800,N_30145);
nand U34061 (N_34061,N_30496,N_31038);
and U34062 (N_34062,N_31246,N_32061);
nand U34063 (N_34063,N_31667,N_32485);
nor U34064 (N_34064,N_31973,N_30243);
nand U34065 (N_34065,N_32000,N_30483);
or U34066 (N_34066,N_31092,N_30646);
and U34067 (N_34067,N_31426,N_30162);
or U34068 (N_34068,N_31374,N_30198);
or U34069 (N_34069,N_30020,N_31485);
nand U34070 (N_34070,N_31463,N_31670);
nor U34071 (N_34071,N_30673,N_30363);
nor U34072 (N_34072,N_30029,N_31675);
or U34073 (N_34073,N_31546,N_30655);
nand U34074 (N_34074,N_30299,N_30507);
nand U34075 (N_34075,N_30900,N_32188);
nor U34076 (N_34076,N_30882,N_32120);
nor U34077 (N_34077,N_31076,N_31334);
or U34078 (N_34078,N_31732,N_30606);
nor U34079 (N_34079,N_30197,N_31366);
xor U34080 (N_34080,N_31344,N_31150);
nor U34081 (N_34081,N_32453,N_30748);
and U34082 (N_34082,N_30610,N_32309);
nand U34083 (N_34083,N_31209,N_30190);
or U34084 (N_34084,N_32211,N_30650);
nand U34085 (N_34085,N_32321,N_30209);
nand U34086 (N_34086,N_30031,N_30319);
nand U34087 (N_34087,N_30850,N_30889);
or U34088 (N_34088,N_30942,N_30354);
nand U34089 (N_34089,N_30369,N_30119);
xor U34090 (N_34090,N_31835,N_32190);
and U34091 (N_34091,N_32211,N_31167);
nand U34092 (N_34092,N_31202,N_31025);
and U34093 (N_34093,N_32264,N_30230);
and U34094 (N_34094,N_32132,N_32498);
and U34095 (N_34095,N_30137,N_31586);
and U34096 (N_34096,N_30171,N_31085);
or U34097 (N_34097,N_31176,N_31462);
nand U34098 (N_34098,N_31963,N_30428);
nor U34099 (N_34099,N_31424,N_30706);
nand U34100 (N_34100,N_30285,N_31012);
xnor U34101 (N_34101,N_30203,N_30631);
or U34102 (N_34102,N_31910,N_31048);
nor U34103 (N_34103,N_31729,N_32232);
nor U34104 (N_34104,N_30276,N_31620);
nor U34105 (N_34105,N_31594,N_30563);
nor U34106 (N_34106,N_30121,N_30596);
xor U34107 (N_34107,N_31413,N_31092);
and U34108 (N_34108,N_30341,N_31819);
and U34109 (N_34109,N_31482,N_30530);
nor U34110 (N_34110,N_30207,N_30578);
nor U34111 (N_34111,N_30625,N_30238);
nand U34112 (N_34112,N_30458,N_31375);
or U34113 (N_34113,N_31378,N_31458);
or U34114 (N_34114,N_32371,N_32420);
or U34115 (N_34115,N_31197,N_31988);
or U34116 (N_34116,N_30857,N_32119);
nand U34117 (N_34117,N_32280,N_30588);
nor U34118 (N_34118,N_31706,N_31488);
and U34119 (N_34119,N_30973,N_31127);
nor U34120 (N_34120,N_31373,N_31604);
and U34121 (N_34121,N_30795,N_32495);
nor U34122 (N_34122,N_31981,N_30885);
and U34123 (N_34123,N_32211,N_30888);
nand U34124 (N_34124,N_31095,N_32047);
or U34125 (N_34125,N_32187,N_30604);
nand U34126 (N_34126,N_31110,N_31196);
nand U34127 (N_34127,N_31890,N_31567);
and U34128 (N_34128,N_31851,N_31160);
and U34129 (N_34129,N_32432,N_31722);
and U34130 (N_34130,N_31135,N_32143);
and U34131 (N_34131,N_31858,N_32366);
or U34132 (N_34132,N_30069,N_32036);
nand U34133 (N_34133,N_31824,N_31163);
nand U34134 (N_34134,N_31075,N_32213);
nor U34135 (N_34135,N_31985,N_30788);
and U34136 (N_34136,N_32182,N_30325);
nand U34137 (N_34137,N_32180,N_30951);
and U34138 (N_34138,N_30750,N_30628);
nor U34139 (N_34139,N_30129,N_32085);
xor U34140 (N_34140,N_31348,N_31759);
nand U34141 (N_34141,N_31904,N_30467);
and U34142 (N_34142,N_31746,N_30415);
nand U34143 (N_34143,N_32195,N_31959);
nand U34144 (N_34144,N_32086,N_30438);
or U34145 (N_34145,N_30989,N_30959);
nand U34146 (N_34146,N_30142,N_31506);
xor U34147 (N_34147,N_32109,N_30306);
nor U34148 (N_34148,N_30792,N_30530);
and U34149 (N_34149,N_31785,N_31126);
or U34150 (N_34150,N_31452,N_32252);
nand U34151 (N_34151,N_31016,N_32189);
or U34152 (N_34152,N_32249,N_31984);
xnor U34153 (N_34153,N_31985,N_31359);
or U34154 (N_34154,N_31872,N_30437);
nor U34155 (N_34155,N_30632,N_30242);
and U34156 (N_34156,N_32139,N_31272);
nor U34157 (N_34157,N_30936,N_30968);
and U34158 (N_34158,N_32386,N_31875);
or U34159 (N_34159,N_30391,N_31418);
nor U34160 (N_34160,N_32011,N_30577);
nor U34161 (N_34161,N_30485,N_32086);
and U34162 (N_34162,N_31942,N_31328);
nor U34163 (N_34163,N_30769,N_31028);
and U34164 (N_34164,N_32044,N_31521);
or U34165 (N_34165,N_31901,N_30843);
or U34166 (N_34166,N_30470,N_32070);
nor U34167 (N_34167,N_30799,N_31062);
nor U34168 (N_34168,N_30894,N_32281);
xnor U34169 (N_34169,N_32492,N_31705);
nand U34170 (N_34170,N_31442,N_31493);
nor U34171 (N_34171,N_30612,N_31089);
or U34172 (N_34172,N_30168,N_31424);
and U34173 (N_34173,N_31418,N_30051);
and U34174 (N_34174,N_32103,N_32068);
nor U34175 (N_34175,N_32435,N_30057);
xor U34176 (N_34176,N_31820,N_30689);
and U34177 (N_34177,N_31201,N_32425);
and U34178 (N_34178,N_30652,N_31372);
nor U34179 (N_34179,N_30067,N_31430);
nand U34180 (N_34180,N_32260,N_31683);
nand U34181 (N_34181,N_31378,N_31107);
xor U34182 (N_34182,N_30556,N_32184);
xnor U34183 (N_34183,N_32383,N_32143);
or U34184 (N_34184,N_32416,N_30118);
and U34185 (N_34185,N_31024,N_31923);
nor U34186 (N_34186,N_31352,N_31344);
xnor U34187 (N_34187,N_31588,N_31757);
nand U34188 (N_34188,N_32457,N_31531);
nand U34189 (N_34189,N_30493,N_30735);
nand U34190 (N_34190,N_31287,N_32172);
nand U34191 (N_34191,N_30476,N_31310);
nor U34192 (N_34192,N_30535,N_31399);
nand U34193 (N_34193,N_32404,N_30255);
nand U34194 (N_34194,N_31048,N_31152);
nor U34195 (N_34195,N_31002,N_30301);
xor U34196 (N_34196,N_30168,N_31944);
nand U34197 (N_34197,N_30489,N_31472);
nand U34198 (N_34198,N_30972,N_32452);
nand U34199 (N_34199,N_30761,N_31630);
nor U34200 (N_34200,N_32241,N_31883);
xnor U34201 (N_34201,N_32397,N_30914);
nand U34202 (N_34202,N_30716,N_32248);
and U34203 (N_34203,N_30332,N_30331);
nor U34204 (N_34204,N_30507,N_32181);
nand U34205 (N_34205,N_31399,N_30383);
and U34206 (N_34206,N_31187,N_30316);
nor U34207 (N_34207,N_30628,N_31306);
and U34208 (N_34208,N_32232,N_31999);
nand U34209 (N_34209,N_30331,N_32172);
nand U34210 (N_34210,N_30545,N_31794);
nor U34211 (N_34211,N_30858,N_32128);
or U34212 (N_34212,N_31681,N_31279);
nand U34213 (N_34213,N_30271,N_31325);
nand U34214 (N_34214,N_32242,N_31103);
nor U34215 (N_34215,N_32076,N_31997);
nand U34216 (N_34216,N_32448,N_31629);
nor U34217 (N_34217,N_31289,N_30143);
or U34218 (N_34218,N_31196,N_30016);
and U34219 (N_34219,N_31538,N_30191);
nor U34220 (N_34220,N_30521,N_31006);
nor U34221 (N_34221,N_31853,N_32029);
and U34222 (N_34222,N_31821,N_31956);
xor U34223 (N_34223,N_32453,N_31602);
and U34224 (N_34224,N_30206,N_31562);
nor U34225 (N_34225,N_31522,N_32121);
nor U34226 (N_34226,N_30312,N_30776);
and U34227 (N_34227,N_30467,N_30647);
xnor U34228 (N_34228,N_32363,N_30794);
and U34229 (N_34229,N_31040,N_31511);
or U34230 (N_34230,N_30730,N_32231);
and U34231 (N_34231,N_30633,N_31699);
nand U34232 (N_34232,N_30189,N_31623);
or U34233 (N_34233,N_32384,N_31599);
xnor U34234 (N_34234,N_30757,N_31955);
nand U34235 (N_34235,N_32259,N_31490);
or U34236 (N_34236,N_31401,N_30007);
xor U34237 (N_34237,N_30189,N_32143);
xor U34238 (N_34238,N_30845,N_31400);
and U34239 (N_34239,N_30012,N_31791);
xnor U34240 (N_34240,N_32443,N_30388);
and U34241 (N_34241,N_30295,N_30263);
or U34242 (N_34242,N_31568,N_31001);
xnor U34243 (N_34243,N_32053,N_30920);
and U34244 (N_34244,N_31262,N_30575);
and U34245 (N_34245,N_30424,N_30292);
xnor U34246 (N_34246,N_32184,N_30872);
and U34247 (N_34247,N_31502,N_31978);
xor U34248 (N_34248,N_30493,N_31408);
nor U34249 (N_34249,N_31371,N_30809);
or U34250 (N_34250,N_30022,N_31142);
or U34251 (N_34251,N_31642,N_31401);
nor U34252 (N_34252,N_31596,N_30056);
xnor U34253 (N_34253,N_30421,N_30859);
nand U34254 (N_34254,N_30236,N_30699);
or U34255 (N_34255,N_32479,N_32237);
and U34256 (N_34256,N_30938,N_31730);
nor U34257 (N_34257,N_32121,N_30302);
nor U34258 (N_34258,N_31673,N_31809);
nor U34259 (N_34259,N_30744,N_30347);
nor U34260 (N_34260,N_30455,N_31689);
xnor U34261 (N_34261,N_31515,N_30384);
and U34262 (N_34262,N_31403,N_30772);
or U34263 (N_34263,N_30691,N_31780);
and U34264 (N_34264,N_32474,N_31791);
or U34265 (N_34265,N_32059,N_31217);
and U34266 (N_34266,N_32009,N_31777);
xnor U34267 (N_34267,N_32351,N_30658);
nor U34268 (N_34268,N_31243,N_30353);
nor U34269 (N_34269,N_30576,N_31576);
nor U34270 (N_34270,N_31402,N_31353);
and U34271 (N_34271,N_32202,N_32027);
nor U34272 (N_34272,N_31500,N_30558);
or U34273 (N_34273,N_30672,N_30573);
nor U34274 (N_34274,N_31646,N_31142);
nand U34275 (N_34275,N_32116,N_30689);
or U34276 (N_34276,N_31454,N_30511);
nor U34277 (N_34277,N_30325,N_30172);
or U34278 (N_34278,N_31648,N_31108);
and U34279 (N_34279,N_30285,N_31332);
or U34280 (N_34280,N_31475,N_30751);
and U34281 (N_34281,N_31394,N_31127);
nand U34282 (N_34282,N_32295,N_32213);
nand U34283 (N_34283,N_30092,N_30216);
nand U34284 (N_34284,N_31399,N_30103);
or U34285 (N_34285,N_31492,N_32158);
nand U34286 (N_34286,N_31141,N_31955);
and U34287 (N_34287,N_32041,N_31696);
nor U34288 (N_34288,N_32356,N_32148);
or U34289 (N_34289,N_30658,N_32098);
or U34290 (N_34290,N_30308,N_30230);
nor U34291 (N_34291,N_30826,N_32104);
and U34292 (N_34292,N_31613,N_30383);
nor U34293 (N_34293,N_30093,N_32185);
or U34294 (N_34294,N_32218,N_30498);
nor U34295 (N_34295,N_30654,N_32161);
nor U34296 (N_34296,N_30181,N_30561);
nor U34297 (N_34297,N_32395,N_31698);
or U34298 (N_34298,N_30163,N_31352);
or U34299 (N_34299,N_31924,N_30083);
and U34300 (N_34300,N_31407,N_30201);
and U34301 (N_34301,N_31011,N_32469);
or U34302 (N_34302,N_31181,N_31218);
nor U34303 (N_34303,N_32260,N_32349);
and U34304 (N_34304,N_30421,N_32144);
nor U34305 (N_34305,N_30266,N_30433);
or U34306 (N_34306,N_32441,N_31201);
nand U34307 (N_34307,N_31181,N_30086);
nand U34308 (N_34308,N_30177,N_32080);
nor U34309 (N_34309,N_31917,N_32183);
and U34310 (N_34310,N_30935,N_31835);
nand U34311 (N_34311,N_31397,N_31587);
or U34312 (N_34312,N_31489,N_31143);
or U34313 (N_34313,N_31488,N_31747);
nand U34314 (N_34314,N_31391,N_30799);
or U34315 (N_34315,N_30038,N_31560);
or U34316 (N_34316,N_31422,N_32278);
xnor U34317 (N_34317,N_31211,N_31960);
nor U34318 (N_34318,N_31820,N_31232);
and U34319 (N_34319,N_30746,N_31622);
or U34320 (N_34320,N_30081,N_30850);
or U34321 (N_34321,N_32433,N_30988);
nor U34322 (N_34322,N_31640,N_31986);
xnor U34323 (N_34323,N_31194,N_31470);
xnor U34324 (N_34324,N_31098,N_31629);
nand U34325 (N_34325,N_32235,N_30912);
xor U34326 (N_34326,N_32094,N_32481);
or U34327 (N_34327,N_31064,N_30737);
or U34328 (N_34328,N_32279,N_31145);
and U34329 (N_34329,N_32224,N_31710);
or U34330 (N_34330,N_32471,N_30841);
nor U34331 (N_34331,N_30127,N_31376);
or U34332 (N_34332,N_32071,N_30394);
nor U34333 (N_34333,N_31195,N_32120);
or U34334 (N_34334,N_30468,N_31587);
or U34335 (N_34335,N_31843,N_31085);
nand U34336 (N_34336,N_31054,N_30366);
or U34337 (N_34337,N_30826,N_30639);
or U34338 (N_34338,N_30466,N_32180);
or U34339 (N_34339,N_30892,N_32284);
xor U34340 (N_34340,N_30417,N_30442);
nor U34341 (N_34341,N_31340,N_31433);
and U34342 (N_34342,N_31814,N_31193);
or U34343 (N_34343,N_32218,N_31877);
and U34344 (N_34344,N_31487,N_32436);
or U34345 (N_34345,N_32043,N_31604);
nor U34346 (N_34346,N_31738,N_30575);
and U34347 (N_34347,N_30454,N_30371);
nand U34348 (N_34348,N_31304,N_30286);
xor U34349 (N_34349,N_31812,N_30668);
and U34350 (N_34350,N_31284,N_30528);
nand U34351 (N_34351,N_30303,N_30107);
nor U34352 (N_34352,N_31696,N_30808);
nand U34353 (N_34353,N_32338,N_32416);
and U34354 (N_34354,N_32236,N_30642);
nor U34355 (N_34355,N_31023,N_30670);
nor U34356 (N_34356,N_30328,N_30245);
or U34357 (N_34357,N_30406,N_31536);
nand U34358 (N_34358,N_31662,N_31128);
and U34359 (N_34359,N_32431,N_31093);
or U34360 (N_34360,N_31939,N_31762);
xor U34361 (N_34361,N_32461,N_30205);
nor U34362 (N_34362,N_30596,N_30508);
xnor U34363 (N_34363,N_32232,N_30684);
xnor U34364 (N_34364,N_31857,N_30775);
nand U34365 (N_34365,N_31961,N_32256);
nor U34366 (N_34366,N_31376,N_31131);
and U34367 (N_34367,N_31879,N_31070);
nand U34368 (N_34368,N_30929,N_32491);
and U34369 (N_34369,N_32276,N_30157);
nand U34370 (N_34370,N_30395,N_30359);
nand U34371 (N_34371,N_30929,N_30637);
nor U34372 (N_34372,N_31365,N_31180);
nand U34373 (N_34373,N_32491,N_30354);
nand U34374 (N_34374,N_30609,N_30542);
nor U34375 (N_34375,N_31951,N_30277);
or U34376 (N_34376,N_30475,N_30667);
and U34377 (N_34377,N_31887,N_32296);
or U34378 (N_34378,N_30859,N_32350);
or U34379 (N_34379,N_31971,N_30290);
nor U34380 (N_34380,N_31519,N_31000);
nand U34381 (N_34381,N_30171,N_31986);
nand U34382 (N_34382,N_31567,N_31371);
nor U34383 (N_34383,N_31479,N_30622);
and U34384 (N_34384,N_31007,N_30875);
nor U34385 (N_34385,N_31478,N_30065);
and U34386 (N_34386,N_30273,N_31880);
xor U34387 (N_34387,N_31150,N_30514);
and U34388 (N_34388,N_32087,N_30263);
nor U34389 (N_34389,N_30366,N_30374);
and U34390 (N_34390,N_31656,N_32213);
or U34391 (N_34391,N_32474,N_30692);
xnor U34392 (N_34392,N_30093,N_32466);
nand U34393 (N_34393,N_31335,N_31296);
nor U34394 (N_34394,N_32217,N_32314);
and U34395 (N_34395,N_31159,N_32359);
or U34396 (N_34396,N_30611,N_30353);
nor U34397 (N_34397,N_31228,N_31302);
and U34398 (N_34398,N_30524,N_30789);
xor U34399 (N_34399,N_30972,N_30414);
nand U34400 (N_34400,N_31728,N_32293);
nor U34401 (N_34401,N_31185,N_30843);
nand U34402 (N_34402,N_31971,N_30378);
or U34403 (N_34403,N_30167,N_30305);
nand U34404 (N_34404,N_32487,N_32259);
and U34405 (N_34405,N_32106,N_30275);
nand U34406 (N_34406,N_30232,N_30667);
and U34407 (N_34407,N_32347,N_30724);
and U34408 (N_34408,N_31551,N_31717);
nor U34409 (N_34409,N_32329,N_31542);
or U34410 (N_34410,N_30959,N_30813);
nand U34411 (N_34411,N_32391,N_30942);
or U34412 (N_34412,N_31425,N_30740);
and U34413 (N_34413,N_30291,N_30532);
xor U34414 (N_34414,N_31033,N_32116);
nor U34415 (N_34415,N_31421,N_30921);
nor U34416 (N_34416,N_31468,N_32476);
and U34417 (N_34417,N_31169,N_31306);
nand U34418 (N_34418,N_30587,N_30968);
and U34419 (N_34419,N_32364,N_30710);
and U34420 (N_34420,N_31614,N_31466);
nor U34421 (N_34421,N_32331,N_31232);
nor U34422 (N_34422,N_31805,N_32171);
nand U34423 (N_34423,N_32249,N_30507);
and U34424 (N_34424,N_32053,N_31716);
or U34425 (N_34425,N_32290,N_31768);
and U34426 (N_34426,N_31677,N_30105);
xnor U34427 (N_34427,N_30918,N_31356);
or U34428 (N_34428,N_31142,N_31954);
nand U34429 (N_34429,N_30775,N_31958);
and U34430 (N_34430,N_32041,N_32409);
or U34431 (N_34431,N_30731,N_30353);
xnor U34432 (N_34432,N_30215,N_31374);
nor U34433 (N_34433,N_30975,N_30374);
nand U34434 (N_34434,N_30131,N_31429);
nand U34435 (N_34435,N_30611,N_30686);
nor U34436 (N_34436,N_30784,N_30821);
nor U34437 (N_34437,N_30687,N_30900);
nor U34438 (N_34438,N_30970,N_30140);
and U34439 (N_34439,N_32434,N_31984);
or U34440 (N_34440,N_31181,N_30663);
nand U34441 (N_34441,N_30014,N_31111);
and U34442 (N_34442,N_30460,N_30729);
nand U34443 (N_34443,N_30814,N_32147);
and U34444 (N_34444,N_31529,N_31079);
xnor U34445 (N_34445,N_30416,N_30261);
or U34446 (N_34446,N_31816,N_30231);
or U34447 (N_34447,N_31021,N_31625);
and U34448 (N_34448,N_32149,N_31547);
nand U34449 (N_34449,N_30948,N_30105);
nand U34450 (N_34450,N_32420,N_30053);
nand U34451 (N_34451,N_31266,N_31299);
nor U34452 (N_34452,N_32312,N_31134);
nor U34453 (N_34453,N_31629,N_30987);
and U34454 (N_34454,N_31968,N_32094);
or U34455 (N_34455,N_30510,N_31042);
and U34456 (N_34456,N_31009,N_32491);
nor U34457 (N_34457,N_31080,N_31285);
nor U34458 (N_34458,N_32195,N_30050);
nand U34459 (N_34459,N_31550,N_32347);
nand U34460 (N_34460,N_30884,N_30822);
or U34461 (N_34461,N_30329,N_32346);
and U34462 (N_34462,N_31969,N_32478);
or U34463 (N_34463,N_32494,N_31761);
or U34464 (N_34464,N_31607,N_30592);
nand U34465 (N_34465,N_32019,N_31617);
and U34466 (N_34466,N_31628,N_31011);
or U34467 (N_34467,N_30853,N_30611);
nor U34468 (N_34468,N_32344,N_30370);
and U34469 (N_34469,N_30557,N_30458);
nand U34470 (N_34470,N_30466,N_30960);
and U34471 (N_34471,N_30307,N_31468);
and U34472 (N_34472,N_30588,N_30898);
nand U34473 (N_34473,N_31060,N_31118);
nor U34474 (N_34474,N_32045,N_30374);
nor U34475 (N_34475,N_32271,N_31720);
nand U34476 (N_34476,N_30261,N_30386);
nor U34477 (N_34477,N_31963,N_31020);
nor U34478 (N_34478,N_32055,N_30922);
xor U34479 (N_34479,N_30775,N_32209);
nor U34480 (N_34480,N_30404,N_32139);
nand U34481 (N_34481,N_30387,N_31062);
or U34482 (N_34482,N_31684,N_30089);
nor U34483 (N_34483,N_30473,N_31418);
or U34484 (N_34484,N_31010,N_30464);
xnor U34485 (N_34485,N_30828,N_31276);
or U34486 (N_34486,N_32243,N_31535);
or U34487 (N_34487,N_31235,N_31234);
nor U34488 (N_34488,N_31004,N_30107);
or U34489 (N_34489,N_30176,N_30504);
and U34490 (N_34490,N_31997,N_32100);
or U34491 (N_34491,N_32205,N_30743);
and U34492 (N_34492,N_31118,N_32130);
xor U34493 (N_34493,N_30007,N_32455);
and U34494 (N_34494,N_31062,N_31315);
or U34495 (N_34495,N_32452,N_30820);
nor U34496 (N_34496,N_30978,N_30057);
xor U34497 (N_34497,N_31646,N_31362);
or U34498 (N_34498,N_30169,N_31255);
nor U34499 (N_34499,N_31635,N_30565);
nand U34500 (N_34500,N_31499,N_32082);
or U34501 (N_34501,N_32202,N_31107);
and U34502 (N_34502,N_31141,N_31574);
and U34503 (N_34503,N_30254,N_31510);
xor U34504 (N_34504,N_30665,N_31788);
nand U34505 (N_34505,N_30559,N_32127);
nand U34506 (N_34506,N_31710,N_31438);
and U34507 (N_34507,N_30300,N_32474);
and U34508 (N_34508,N_31142,N_30064);
or U34509 (N_34509,N_30767,N_31934);
or U34510 (N_34510,N_30885,N_31559);
or U34511 (N_34511,N_31621,N_32326);
xnor U34512 (N_34512,N_31630,N_31204);
nor U34513 (N_34513,N_31006,N_30887);
or U34514 (N_34514,N_32061,N_32195);
and U34515 (N_34515,N_30234,N_31996);
nand U34516 (N_34516,N_30438,N_31601);
nor U34517 (N_34517,N_32230,N_30025);
and U34518 (N_34518,N_30731,N_30053);
xnor U34519 (N_34519,N_30568,N_32071);
and U34520 (N_34520,N_32368,N_30195);
and U34521 (N_34521,N_32089,N_30500);
or U34522 (N_34522,N_32336,N_30183);
and U34523 (N_34523,N_30142,N_31264);
nor U34524 (N_34524,N_30888,N_31109);
or U34525 (N_34525,N_30510,N_30688);
and U34526 (N_34526,N_30952,N_30909);
or U34527 (N_34527,N_30182,N_32269);
nor U34528 (N_34528,N_30128,N_31547);
nand U34529 (N_34529,N_32495,N_30474);
nand U34530 (N_34530,N_31713,N_30312);
xnor U34531 (N_34531,N_31475,N_31066);
or U34532 (N_34532,N_30088,N_32397);
or U34533 (N_34533,N_30892,N_30543);
nand U34534 (N_34534,N_31517,N_31542);
xnor U34535 (N_34535,N_31059,N_32122);
nor U34536 (N_34536,N_30723,N_30489);
nand U34537 (N_34537,N_30514,N_31001);
nand U34538 (N_34538,N_31007,N_30068);
nand U34539 (N_34539,N_31559,N_31789);
nor U34540 (N_34540,N_32292,N_30722);
and U34541 (N_34541,N_31423,N_32173);
nor U34542 (N_34542,N_32493,N_31160);
nor U34543 (N_34543,N_31206,N_32278);
or U34544 (N_34544,N_32097,N_30092);
xnor U34545 (N_34545,N_32048,N_30174);
or U34546 (N_34546,N_31257,N_32129);
and U34547 (N_34547,N_31577,N_31111);
or U34548 (N_34548,N_32405,N_32410);
or U34549 (N_34549,N_32382,N_32301);
and U34550 (N_34550,N_31476,N_31045);
nand U34551 (N_34551,N_30088,N_30590);
and U34552 (N_34552,N_32499,N_30134);
nor U34553 (N_34553,N_31464,N_32317);
and U34554 (N_34554,N_30440,N_30379);
and U34555 (N_34555,N_32442,N_30392);
xnor U34556 (N_34556,N_30807,N_31259);
xnor U34557 (N_34557,N_32059,N_31603);
or U34558 (N_34558,N_31789,N_31288);
nand U34559 (N_34559,N_30393,N_30237);
nand U34560 (N_34560,N_31008,N_31809);
nand U34561 (N_34561,N_30531,N_30057);
or U34562 (N_34562,N_31984,N_30783);
nor U34563 (N_34563,N_32038,N_30036);
and U34564 (N_34564,N_30710,N_30765);
or U34565 (N_34565,N_30311,N_31395);
nand U34566 (N_34566,N_32173,N_30017);
nand U34567 (N_34567,N_30391,N_32193);
nor U34568 (N_34568,N_31353,N_31272);
nor U34569 (N_34569,N_31405,N_30438);
nor U34570 (N_34570,N_30696,N_30015);
nand U34571 (N_34571,N_31956,N_31966);
and U34572 (N_34572,N_30411,N_31274);
xor U34573 (N_34573,N_30651,N_30829);
or U34574 (N_34574,N_32188,N_31661);
and U34575 (N_34575,N_30403,N_30143);
and U34576 (N_34576,N_31644,N_32253);
xor U34577 (N_34577,N_31493,N_31193);
nand U34578 (N_34578,N_30775,N_31757);
nor U34579 (N_34579,N_31354,N_30568);
or U34580 (N_34580,N_31418,N_31181);
nor U34581 (N_34581,N_31737,N_31930);
nand U34582 (N_34582,N_31266,N_31051);
nand U34583 (N_34583,N_32316,N_31043);
and U34584 (N_34584,N_31444,N_30251);
nand U34585 (N_34585,N_30715,N_31829);
or U34586 (N_34586,N_32035,N_31666);
or U34587 (N_34587,N_32397,N_31036);
xnor U34588 (N_34588,N_32075,N_30189);
nand U34589 (N_34589,N_31497,N_32225);
nor U34590 (N_34590,N_31834,N_31981);
or U34591 (N_34591,N_31030,N_32014);
or U34592 (N_34592,N_31389,N_31328);
and U34593 (N_34593,N_31209,N_30280);
or U34594 (N_34594,N_30948,N_32340);
and U34595 (N_34595,N_31247,N_32333);
nor U34596 (N_34596,N_31649,N_30115);
nor U34597 (N_34597,N_32415,N_32281);
and U34598 (N_34598,N_30349,N_31887);
or U34599 (N_34599,N_31643,N_30298);
and U34600 (N_34600,N_30233,N_32367);
or U34601 (N_34601,N_31154,N_32342);
xor U34602 (N_34602,N_31910,N_31205);
nand U34603 (N_34603,N_31011,N_30542);
nor U34604 (N_34604,N_30576,N_31737);
or U34605 (N_34605,N_30489,N_31831);
nor U34606 (N_34606,N_31711,N_32417);
nor U34607 (N_34607,N_32164,N_32484);
xor U34608 (N_34608,N_32145,N_31337);
or U34609 (N_34609,N_30495,N_32151);
and U34610 (N_34610,N_31223,N_32152);
nor U34611 (N_34611,N_31814,N_30830);
nor U34612 (N_34612,N_32240,N_31519);
nand U34613 (N_34613,N_32042,N_30389);
or U34614 (N_34614,N_31545,N_32163);
nand U34615 (N_34615,N_32393,N_32247);
and U34616 (N_34616,N_30516,N_32381);
and U34617 (N_34617,N_31478,N_32434);
nor U34618 (N_34618,N_32434,N_31129);
xnor U34619 (N_34619,N_32031,N_30112);
nand U34620 (N_34620,N_31965,N_31879);
or U34621 (N_34621,N_31082,N_30533);
or U34622 (N_34622,N_31235,N_31400);
xnor U34623 (N_34623,N_30068,N_30518);
and U34624 (N_34624,N_30048,N_30670);
nor U34625 (N_34625,N_30154,N_30323);
xor U34626 (N_34626,N_31946,N_32041);
nor U34627 (N_34627,N_32438,N_31425);
nand U34628 (N_34628,N_32152,N_31673);
nand U34629 (N_34629,N_30749,N_30823);
nor U34630 (N_34630,N_31898,N_30668);
nand U34631 (N_34631,N_30680,N_30133);
nand U34632 (N_34632,N_31363,N_31404);
nand U34633 (N_34633,N_32292,N_32390);
or U34634 (N_34634,N_31932,N_31968);
nand U34635 (N_34635,N_31251,N_32429);
nor U34636 (N_34636,N_31790,N_31075);
nor U34637 (N_34637,N_31223,N_32156);
or U34638 (N_34638,N_32431,N_31913);
xnor U34639 (N_34639,N_30966,N_30007);
nor U34640 (N_34640,N_31947,N_31754);
or U34641 (N_34641,N_31803,N_30791);
and U34642 (N_34642,N_31302,N_30454);
xnor U34643 (N_34643,N_30166,N_30215);
and U34644 (N_34644,N_30363,N_31474);
or U34645 (N_34645,N_31897,N_31711);
or U34646 (N_34646,N_30787,N_31156);
nor U34647 (N_34647,N_31281,N_30701);
nor U34648 (N_34648,N_31447,N_31823);
nand U34649 (N_34649,N_31792,N_31463);
and U34650 (N_34650,N_30228,N_31945);
and U34651 (N_34651,N_31827,N_32257);
or U34652 (N_34652,N_30904,N_31636);
or U34653 (N_34653,N_31496,N_31787);
or U34654 (N_34654,N_31605,N_30139);
nor U34655 (N_34655,N_30130,N_30648);
or U34656 (N_34656,N_31578,N_32269);
nor U34657 (N_34657,N_31804,N_30379);
or U34658 (N_34658,N_31740,N_31162);
nor U34659 (N_34659,N_30469,N_32177);
nor U34660 (N_34660,N_32437,N_31687);
nor U34661 (N_34661,N_32112,N_30660);
and U34662 (N_34662,N_31665,N_30487);
and U34663 (N_34663,N_31351,N_30231);
or U34664 (N_34664,N_30865,N_30719);
xnor U34665 (N_34665,N_31699,N_30167);
and U34666 (N_34666,N_31783,N_31232);
nand U34667 (N_34667,N_30768,N_31157);
and U34668 (N_34668,N_31982,N_31452);
xor U34669 (N_34669,N_30196,N_30755);
or U34670 (N_34670,N_30877,N_31382);
and U34671 (N_34671,N_30487,N_31198);
and U34672 (N_34672,N_31141,N_31525);
or U34673 (N_34673,N_32428,N_30594);
nor U34674 (N_34674,N_30768,N_31643);
and U34675 (N_34675,N_32362,N_32376);
and U34676 (N_34676,N_30183,N_30335);
or U34677 (N_34677,N_32349,N_32441);
or U34678 (N_34678,N_31098,N_31263);
and U34679 (N_34679,N_30779,N_30274);
and U34680 (N_34680,N_30363,N_32178);
and U34681 (N_34681,N_31199,N_31593);
or U34682 (N_34682,N_30796,N_30876);
or U34683 (N_34683,N_32458,N_30632);
nand U34684 (N_34684,N_31801,N_31538);
or U34685 (N_34685,N_30106,N_31831);
nand U34686 (N_34686,N_32419,N_32405);
and U34687 (N_34687,N_32375,N_32392);
or U34688 (N_34688,N_31549,N_31772);
nand U34689 (N_34689,N_32421,N_32363);
nor U34690 (N_34690,N_30514,N_31545);
nor U34691 (N_34691,N_30778,N_32390);
nor U34692 (N_34692,N_30108,N_30935);
nor U34693 (N_34693,N_31945,N_32245);
or U34694 (N_34694,N_30877,N_30380);
nand U34695 (N_34695,N_30733,N_30459);
nand U34696 (N_34696,N_31829,N_30551);
and U34697 (N_34697,N_31021,N_32470);
or U34698 (N_34698,N_32265,N_31063);
or U34699 (N_34699,N_30508,N_30128);
or U34700 (N_34700,N_30246,N_31398);
or U34701 (N_34701,N_30806,N_31726);
and U34702 (N_34702,N_30739,N_32010);
nand U34703 (N_34703,N_30053,N_30319);
xor U34704 (N_34704,N_30495,N_31915);
nor U34705 (N_34705,N_32421,N_31272);
nand U34706 (N_34706,N_31744,N_31458);
or U34707 (N_34707,N_32064,N_31100);
or U34708 (N_34708,N_30063,N_32291);
and U34709 (N_34709,N_31467,N_30530);
and U34710 (N_34710,N_32295,N_30223);
and U34711 (N_34711,N_31554,N_31705);
nor U34712 (N_34712,N_32320,N_31992);
and U34713 (N_34713,N_31076,N_31813);
or U34714 (N_34714,N_30552,N_31797);
nor U34715 (N_34715,N_32374,N_30897);
nand U34716 (N_34716,N_31600,N_30141);
nand U34717 (N_34717,N_31234,N_30267);
xor U34718 (N_34718,N_31396,N_31360);
or U34719 (N_34719,N_31094,N_30546);
nand U34720 (N_34720,N_30982,N_31904);
and U34721 (N_34721,N_32017,N_30132);
and U34722 (N_34722,N_30235,N_30135);
nor U34723 (N_34723,N_32037,N_32313);
xnor U34724 (N_34724,N_32416,N_30484);
and U34725 (N_34725,N_32161,N_30816);
nor U34726 (N_34726,N_32185,N_31081);
and U34727 (N_34727,N_30036,N_30492);
or U34728 (N_34728,N_30607,N_30023);
and U34729 (N_34729,N_31192,N_31058);
nand U34730 (N_34730,N_31585,N_32248);
and U34731 (N_34731,N_30479,N_30220);
xor U34732 (N_34732,N_30761,N_31694);
xor U34733 (N_34733,N_32077,N_32442);
nand U34734 (N_34734,N_30627,N_30172);
nor U34735 (N_34735,N_30941,N_30897);
or U34736 (N_34736,N_32286,N_30162);
or U34737 (N_34737,N_31483,N_30196);
or U34738 (N_34738,N_31655,N_31716);
and U34739 (N_34739,N_30040,N_31415);
nand U34740 (N_34740,N_30912,N_31370);
nand U34741 (N_34741,N_30742,N_30540);
nor U34742 (N_34742,N_31004,N_30237);
or U34743 (N_34743,N_32049,N_31668);
nand U34744 (N_34744,N_31462,N_31184);
nand U34745 (N_34745,N_30873,N_30044);
nor U34746 (N_34746,N_30697,N_31771);
and U34747 (N_34747,N_30468,N_30198);
or U34748 (N_34748,N_30051,N_31729);
nand U34749 (N_34749,N_30993,N_32036);
nor U34750 (N_34750,N_30383,N_30147);
and U34751 (N_34751,N_31765,N_31306);
nand U34752 (N_34752,N_31912,N_31251);
and U34753 (N_34753,N_30364,N_30570);
and U34754 (N_34754,N_30209,N_30796);
and U34755 (N_34755,N_30054,N_30298);
nand U34756 (N_34756,N_31804,N_32233);
or U34757 (N_34757,N_31620,N_31129);
and U34758 (N_34758,N_31954,N_32355);
or U34759 (N_34759,N_31492,N_32177);
and U34760 (N_34760,N_31801,N_31593);
nand U34761 (N_34761,N_31072,N_31650);
and U34762 (N_34762,N_31432,N_31007);
nor U34763 (N_34763,N_32436,N_30996);
and U34764 (N_34764,N_32484,N_31981);
or U34765 (N_34765,N_30043,N_30905);
xor U34766 (N_34766,N_30279,N_30549);
and U34767 (N_34767,N_31952,N_30125);
or U34768 (N_34768,N_32325,N_30953);
or U34769 (N_34769,N_30892,N_31251);
nand U34770 (N_34770,N_30922,N_30677);
nand U34771 (N_34771,N_31890,N_31645);
or U34772 (N_34772,N_31656,N_30943);
nand U34773 (N_34773,N_31747,N_30563);
nor U34774 (N_34774,N_31551,N_31252);
nor U34775 (N_34775,N_30127,N_30653);
nand U34776 (N_34776,N_30430,N_32227);
or U34777 (N_34777,N_31671,N_31890);
xnor U34778 (N_34778,N_30200,N_31183);
nor U34779 (N_34779,N_31363,N_32097);
xor U34780 (N_34780,N_30674,N_32340);
nand U34781 (N_34781,N_31918,N_30999);
or U34782 (N_34782,N_32424,N_32370);
nor U34783 (N_34783,N_30118,N_31150);
nor U34784 (N_34784,N_31432,N_31269);
nor U34785 (N_34785,N_31788,N_30012);
and U34786 (N_34786,N_30083,N_32186);
or U34787 (N_34787,N_30774,N_30703);
and U34788 (N_34788,N_32004,N_30829);
and U34789 (N_34789,N_30759,N_32159);
and U34790 (N_34790,N_31477,N_31699);
and U34791 (N_34791,N_30481,N_30730);
nor U34792 (N_34792,N_30689,N_30320);
and U34793 (N_34793,N_30841,N_30471);
nand U34794 (N_34794,N_30883,N_30393);
or U34795 (N_34795,N_31206,N_32007);
nor U34796 (N_34796,N_32135,N_30796);
nor U34797 (N_34797,N_31054,N_31618);
or U34798 (N_34798,N_30325,N_31389);
xnor U34799 (N_34799,N_32097,N_32460);
nand U34800 (N_34800,N_30811,N_30055);
xnor U34801 (N_34801,N_31532,N_30223);
nor U34802 (N_34802,N_30914,N_31355);
xnor U34803 (N_34803,N_30948,N_30055);
and U34804 (N_34804,N_30530,N_30870);
xnor U34805 (N_34805,N_30204,N_30192);
nor U34806 (N_34806,N_31219,N_31307);
nand U34807 (N_34807,N_30529,N_30143);
or U34808 (N_34808,N_30066,N_32286);
or U34809 (N_34809,N_30411,N_30339);
or U34810 (N_34810,N_30383,N_31231);
or U34811 (N_34811,N_30413,N_30495);
or U34812 (N_34812,N_30310,N_32335);
nor U34813 (N_34813,N_30927,N_30438);
xnor U34814 (N_34814,N_32053,N_32416);
nand U34815 (N_34815,N_30826,N_32019);
and U34816 (N_34816,N_31807,N_30586);
or U34817 (N_34817,N_30139,N_31263);
and U34818 (N_34818,N_30281,N_30125);
nand U34819 (N_34819,N_31013,N_31282);
nor U34820 (N_34820,N_32356,N_32104);
and U34821 (N_34821,N_30603,N_32116);
and U34822 (N_34822,N_32305,N_31188);
nand U34823 (N_34823,N_30971,N_30411);
or U34824 (N_34824,N_31749,N_32010);
nor U34825 (N_34825,N_31453,N_31021);
and U34826 (N_34826,N_30765,N_31027);
and U34827 (N_34827,N_31062,N_30095);
nand U34828 (N_34828,N_30089,N_30229);
or U34829 (N_34829,N_32049,N_30345);
nor U34830 (N_34830,N_30891,N_31787);
and U34831 (N_34831,N_30188,N_31846);
or U34832 (N_34832,N_30501,N_31423);
nand U34833 (N_34833,N_30691,N_30446);
and U34834 (N_34834,N_30545,N_30186);
or U34835 (N_34835,N_31177,N_32268);
or U34836 (N_34836,N_31058,N_31794);
or U34837 (N_34837,N_30835,N_30187);
or U34838 (N_34838,N_30667,N_32114);
or U34839 (N_34839,N_32329,N_32027);
nor U34840 (N_34840,N_32055,N_31708);
or U34841 (N_34841,N_30939,N_31733);
and U34842 (N_34842,N_30935,N_30148);
nand U34843 (N_34843,N_30842,N_30464);
and U34844 (N_34844,N_30700,N_31942);
nor U34845 (N_34845,N_30504,N_30027);
and U34846 (N_34846,N_31528,N_30101);
or U34847 (N_34847,N_30329,N_30900);
xnor U34848 (N_34848,N_30645,N_30865);
nor U34849 (N_34849,N_32460,N_30279);
and U34850 (N_34850,N_31264,N_30148);
or U34851 (N_34851,N_31935,N_30382);
and U34852 (N_34852,N_31390,N_31807);
and U34853 (N_34853,N_30342,N_30950);
nand U34854 (N_34854,N_31083,N_31132);
or U34855 (N_34855,N_30042,N_31147);
nand U34856 (N_34856,N_30750,N_32451);
or U34857 (N_34857,N_30131,N_30963);
nor U34858 (N_34858,N_31439,N_30921);
nor U34859 (N_34859,N_32031,N_32087);
nor U34860 (N_34860,N_31449,N_30382);
and U34861 (N_34861,N_30366,N_31344);
nand U34862 (N_34862,N_30731,N_30821);
nor U34863 (N_34863,N_32485,N_30826);
and U34864 (N_34864,N_32170,N_32034);
nand U34865 (N_34865,N_31940,N_32142);
or U34866 (N_34866,N_31335,N_30595);
nand U34867 (N_34867,N_30038,N_31305);
and U34868 (N_34868,N_30520,N_31252);
nand U34869 (N_34869,N_30421,N_30635);
nand U34870 (N_34870,N_31653,N_32139);
or U34871 (N_34871,N_31457,N_32036);
nand U34872 (N_34872,N_30360,N_31175);
nand U34873 (N_34873,N_31280,N_31304);
and U34874 (N_34874,N_31381,N_30197);
or U34875 (N_34875,N_30792,N_32043);
and U34876 (N_34876,N_31131,N_30798);
nor U34877 (N_34877,N_31544,N_31651);
nand U34878 (N_34878,N_32485,N_30189);
nor U34879 (N_34879,N_31932,N_31139);
and U34880 (N_34880,N_30903,N_31956);
nand U34881 (N_34881,N_32447,N_31621);
and U34882 (N_34882,N_30400,N_30670);
and U34883 (N_34883,N_30134,N_31571);
nand U34884 (N_34884,N_31346,N_31564);
nor U34885 (N_34885,N_31321,N_30908);
nand U34886 (N_34886,N_31467,N_31678);
and U34887 (N_34887,N_31991,N_31670);
nor U34888 (N_34888,N_30265,N_30628);
nor U34889 (N_34889,N_31859,N_31491);
or U34890 (N_34890,N_31990,N_31314);
and U34891 (N_34891,N_30515,N_30754);
or U34892 (N_34892,N_31355,N_31590);
or U34893 (N_34893,N_32259,N_31856);
or U34894 (N_34894,N_30911,N_30779);
and U34895 (N_34895,N_31275,N_32294);
or U34896 (N_34896,N_31413,N_31948);
nand U34897 (N_34897,N_31596,N_32328);
nand U34898 (N_34898,N_31775,N_31506);
nand U34899 (N_34899,N_31523,N_31213);
nor U34900 (N_34900,N_32061,N_31805);
and U34901 (N_34901,N_32262,N_30097);
nand U34902 (N_34902,N_32333,N_31455);
nor U34903 (N_34903,N_32482,N_31559);
nor U34904 (N_34904,N_31534,N_31224);
nand U34905 (N_34905,N_30280,N_31416);
nor U34906 (N_34906,N_30860,N_30620);
nand U34907 (N_34907,N_31754,N_30457);
and U34908 (N_34908,N_30294,N_31982);
or U34909 (N_34909,N_30039,N_30382);
nand U34910 (N_34910,N_31878,N_30932);
nor U34911 (N_34911,N_31956,N_30731);
nand U34912 (N_34912,N_30673,N_30006);
nand U34913 (N_34913,N_31128,N_31544);
nor U34914 (N_34914,N_31160,N_32324);
nand U34915 (N_34915,N_30265,N_30991);
nand U34916 (N_34916,N_30616,N_31585);
or U34917 (N_34917,N_31359,N_32210);
and U34918 (N_34918,N_31285,N_31848);
nor U34919 (N_34919,N_30846,N_30978);
nor U34920 (N_34920,N_32447,N_30472);
xnor U34921 (N_34921,N_30252,N_31024);
or U34922 (N_34922,N_32091,N_31926);
nand U34923 (N_34923,N_30753,N_32422);
or U34924 (N_34924,N_32418,N_31942);
or U34925 (N_34925,N_32416,N_32268);
nor U34926 (N_34926,N_31405,N_30851);
xor U34927 (N_34927,N_30478,N_31543);
or U34928 (N_34928,N_30935,N_32266);
or U34929 (N_34929,N_32094,N_31302);
or U34930 (N_34930,N_31080,N_31296);
and U34931 (N_34931,N_30634,N_31071);
or U34932 (N_34932,N_30568,N_32266);
xnor U34933 (N_34933,N_30036,N_32009);
nand U34934 (N_34934,N_30315,N_31417);
and U34935 (N_34935,N_31101,N_31142);
nor U34936 (N_34936,N_30557,N_32016);
nand U34937 (N_34937,N_30474,N_31373);
and U34938 (N_34938,N_32224,N_31340);
nor U34939 (N_34939,N_31493,N_31289);
and U34940 (N_34940,N_30795,N_30668);
nor U34941 (N_34941,N_31358,N_31378);
nor U34942 (N_34942,N_31642,N_30972);
xnor U34943 (N_34943,N_31160,N_32490);
or U34944 (N_34944,N_31600,N_31895);
nor U34945 (N_34945,N_32266,N_31154);
nand U34946 (N_34946,N_31900,N_31578);
or U34947 (N_34947,N_30320,N_30657);
nor U34948 (N_34948,N_31522,N_30181);
nand U34949 (N_34949,N_31410,N_30256);
or U34950 (N_34950,N_30653,N_31965);
nand U34951 (N_34951,N_30539,N_30668);
or U34952 (N_34952,N_30126,N_30180);
nor U34953 (N_34953,N_30517,N_31150);
or U34954 (N_34954,N_30279,N_31395);
or U34955 (N_34955,N_32013,N_30053);
or U34956 (N_34956,N_32065,N_31287);
and U34957 (N_34957,N_30370,N_30231);
nor U34958 (N_34958,N_31455,N_30797);
or U34959 (N_34959,N_30980,N_32324);
nand U34960 (N_34960,N_31502,N_31012);
nand U34961 (N_34961,N_32248,N_30553);
nor U34962 (N_34962,N_30563,N_30303);
xnor U34963 (N_34963,N_30345,N_30247);
nor U34964 (N_34964,N_30556,N_31220);
and U34965 (N_34965,N_31888,N_30942);
nor U34966 (N_34966,N_30213,N_31636);
nand U34967 (N_34967,N_31908,N_31048);
nand U34968 (N_34968,N_30643,N_30467);
or U34969 (N_34969,N_32356,N_32300);
nor U34970 (N_34970,N_32304,N_31460);
and U34971 (N_34971,N_30429,N_30682);
or U34972 (N_34972,N_30180,N_30790);
and U34973 (N_34973,N_32033,N_30299);
and U34974 (N_34974,N_32092,N_30874);
or U34975 (N_34975,N_31921,N_30432);
and U34976 (N_34976,N_32284,N_31948);
nor U34977 (N_34977,N_32361,N_31785);
or U34978 (N_34978,N_30998,N_30180);
nor U34979 (N_34979,N_31845,N_30149);
and U34980 (N_34980,N_31669,N_31628);
or U34981 (N_34981,N_32451,N_30866);
and U34982 (N_34982,N_30924,N_31718);
xnor U34983 (N_34983,N_31788,N_30049);
or U34984 (N_34984,N_32212,N_30064);
and U34985 (N_34985,N_31452,N_30596);
or U34986 (N_34986,N_31688,N_31734);
nor U34987 (N_34987,N_31232,N_30129);
nor U34988 (N_34988,N_30321,N_30229);
nand U34989 (N_34989,N_32072,N_31499);
nand U34990 (N_34990,N_30984,N_30821);
nor U34991 (N_34991,N_30072,N_31160);
xnor U34992 (N_34992,N_31369,N_32163);
and U34993 (N_34993,N_31762,N_30902);
or U34994 (N_34994,N_31288,N_30839);
nand U34995 (N_34995,N_30624,N_30460);
and U34996 (N_34996,N_30401,N_32095);
nor U34997 (N_34997,N_30172,N_31639);
nor U34998 (N_34998,N_30208,N_32024);
nand U34999 (N_34999,N_31843,N_30226);
nor U35000 (N_35000,N_34388,N_34889);
xor U35001 (N_35001,N_33845,N_34096);
or U35002 (N_35002,N_34758,N_32666);
nand U35003 (N_35003,N_32864,N_32827);
nand U35004 (N_35004,N_33344,N_32620);
nor U35005 (N_35005,N_33319,N_32786);
nand U35006 (N_35006,N_33494,N_34979);
nand U35007 (N_35007,N_34586,N_34142);
nor U35008 (N_35008,N_34613,N_33604);
nor U35009 (N_35009,N_33807,N_34249);
xor U35010 (N_35010,N_34293,N_33918);
or U35011 (N_35011,N_34395,N_33191);
nand U35012 (N_35012,N_32761,N_33956);
and U35013 (N_35013,N_34159,N_34163);
nand U35014 (N_35014,N_34632,N_34377);
nor U35015 (N_35015,N_34458,N_33819);
and U35016 (N_35016,N_34993,N_34480);
and U35017 (N_35017,N_33505,N_33618);
nand U35018 (N_35018,N_33353,N_32590);
nand U35019 (N_35019,N_34174,N_33431);
nand U35020 (N_35020,N_34024,N_32759);
or U35021 (N_35021,N_33787,N_33904);
and U35022 (N_35022,N_34963,N_34074);
or U35023 (N_35023,N_34802,N_34896);
nor U35024 (N_35024,N_32867,N_33728);
nor U35025 (N_35025,N_34140,N_33302);
and U35026 (N_35026,N_33199,N_34751);
and U35027 (N_35027,N_33278,N_34723);
and U35028 (N_35028,N_34981,N_33452);
nand U35029 (N_35029,N_34176,N_34004);
nand U35030 (N_35030,N_34481,N_34513);
nor U35031 (N_35031,N_33055,N_33210);
nand U35032 (N_35032,N_32605,N_32778);
or U35033 (N_35033,N_33391,N_34591);
and U35034 (N_35034,N_32598,N_32911);
nor U35035 (N_35035,N_34523,N_34726);
or U35036 (N_35036,N_34210,N_33409);
nand U35037 (N_35037,N_32965,N_32527);
or U35038 (N_35038,N_33639,N_34029);
nor U35039 (N_35039,N_34309,N_34128);
nor U35040 (N_35040,N_32797,N_32767);
and U35041 (N_35041,N_33980,N_34023);
nor U35042 (N_35042,N_33388,N_33635);
and U35043 (N_35043,N_33272,N_34903);
or U35044 (N_35044,N_32947,N_34961);
nor U35045 (N_35045,N_32564,N_33362);
nor U35046 (N_35046,N_34930,N_32983);
nand U35047 (N_35047,N_32512,N_32636);
or U35048 (N_35048,N_34100,N_32972);
nor U35049 (N_35049,N_32630,N_32897);
nor U35050 (N_35050,N_33258,N_32889);
xnor U35051 (N_35051,N_33966,N_33839);
nor U35052 (N_35052,N_33153,N_33252);
nor U35053 (N_35053,N_33954,N_33912);
nand U35054 (N_35054,N_34273,N_34967);
nand U35055 (N_35055,N_33856,N_33069);
and U35056 (N_35056,N_33203,N_34925);
nor U35057 (N_35057,N_33529,N_33212);
and U35058 (N_35058,N_33481,N_33827);
and U35059 (N_35059,N_32702,N_33123);
nor U35060 (N_35060,N_34404,N_34693);
and U35061 (N_35061,N_33475,N_32891);
nand U35062 (N_35062,N_34265,N_32751);
or U35063 (N_35063,N_34561,N_33242);
nand U35064 (N_35064,N_32909,N_34356);
nand U35065 (N_35065,N_34972,N_34824);
nor U35066 (N_35066,N_34821,N_33401);
nor U35067 (N_35067,N_34784,N_34566);
nor U35068 (N_35068,N_33235,N_34699);
or U35069 (N_35069,N_33638,N_32775);
and U35070 (N_35070,N_34076,N_33988);
nand U35071 (N_35071,N_33854,N_33369);
or U35072 (N_35072,N_33150,N_34679);
nor U35073 (N_35073,N_33117,N_33585);
and U35074 (N_35074,N_33818,N_34898);
nor U35075 (N_35075,N_34522,N_34563);
or U35076 (N_35076,N_33310,N_33681);
and U35077 (N_35077,N_32752,N_32510);
and U35078 (N_35078,N_33370,N_32612);
or U35079 (N_35079,N_33642,N_34757);
or U35080 (N_35080,N_33326,N_34197);
and U35081 (N_35081,N_32791,N_34292);
and U35082 (N_35082,N_32503,N_33159);
or U35083 (N_35083,N_33755,N_34126);
nor U35084 (N_35084,N_33135,N_33865);
nand U35085 (N_35085,N_34676,N_32648);
nor U35086 (N_35086,N_32741,N_34349);
nand U35087 (N_35087,N_34158,N_34841);
and U35088 (N_35088,N_34028,N_34101);
nor U35089 (N_35089,N_34230,N_34031);
nand U35090 (N_35090,N_33567,N_32705);
and U35091 (N_35091,N_33853,N_34242);
nor U35092 (N_35092,N_33944,N_34663);
and U35093 (N_35093,N_32899,N_34316);
nor U35094 (N_35094,N_34867,N_32833);
and U35095 (N_35095,N_32764,N_34907);
or U35096 (N_35096,N_34648,N_32959);
or U35097 (N_35097,N_32933,N_34295);
nand U35098 (N_35098,N_34402,N_32878);
or U35099 (N_35099,N_32927,N_33561);
nand U35100 (N_35100,N_34696,N_33596);
xnor U35101 (N_35101,N_33793,N_34593);
xor U35102 (N_35102,N_34562,N_33520);
or U35103 (N_35103,N_32599,N_34542);
or U35104 (N_35104,N_34799,N_32543);
or U35105 (N_35105,N_34618,N_33393);
nand U35106 (N_35106,N_34569,N_32828);
nor U35107 (N_35107,N_34653,N_34521);
xnor U35108 (N_35108,N_33611,N_34836);
or U35109 (N_35109,N_34118,N_34897);
and U35110 (N_35110,N_32603,N_34116);
and U35111 (N_35111,N_32766,N_34795);
or U35112 (N_35112,N_32614,N_34037);
nand U35113 (N_35113,N_34073,N_34672);
nor U35114 (N_35114,N_33586,N_34279);
nor U35115 (N_35115,N_32868,N_34235);
and U35116 (N_35116,N_34188,N_33994);
and U35117 (N_35117,N_33027,N_33072);
and U35118 (N_35118,N_33770,N_33679);
and U35119 (N_35119,N_33260,N_34716);
nor U35120 (N_35120,N_34734,N_34831);
and U35121 (N_35121,N_34424,N_33958);
nand U35122 (N_35122,N_34280,N_34690);
and U35123 (N_35123,N_32780,N_34386);
nand U35124 (N_35124,N_32526,N_32934);
nor U35125 (N_35125,N_33795,N_34717);
xor U35126 (N_35126,N_32967,N_34435);
nand U35127 (N_35127,N_33894,N_34953);
nand U35128 (N_35128,N_33646,N_32872);
nand U35129 (N_35129,N_34772,N_33716);
nor U35130 (N_35130,N_33910,N_34305);
or U35131 (N_35131,N_34426,N_33552);
nor U35132 (N_35132,N_34874,N_33985);
and U35133 (N_35133,N_33050,N_32976);
or U35134 (N_35134,N_33659,N_34661);
or U35135 (N_35135,N_32701,N_33566);
nand U35136 (N_35136,N_34484,N_33935);
nand U35137 (N_35137,N_33809,N_34588);
or U35138 (N_35138,N_34208,N_32755);
and U35139 (N_35139,N_32670,N_34880);
nand U35140 (N_35140,N_33024,N_33390);
and U35141 (N_35141,N_33884,N_34928);
nor U35142 (N_35142,N_33136,N_32771);
nand U35143 (N_35143,N_33211,N_34936);
nand U35144 (N_35144,N_34674,N_32726);
nand U35145 (N_35145,N_34636,N_32516);
and U35146 (N_35146,N_33957,N_32578);
or U35147 (N_35147,N_34289,N_33231);
nor U35148 (N_35148,N_34317,N_34406);
or U35149 (N_35149,N_33164,N_34145);
nor U35150 (N_35150,N_33998,N_34493);
nor U35151 (N_35151,N_34638,N_34336);
nor U35152 (N_35152,N_34442,N_33553);
or U35153 (N_35153,N_32749,N_33620);
nor U35154 (N_35154,N_34006,N_32896);
and U35155 (N_35155,N_33876,N_34518);
or U35156 (N_35156,N_33906,N_34822);
nor U35157 (N_35157,N_34740,N_33513);
xor U35158 (N_35158,N_34320,N_34590);
nor U35159 (N_35159,N_33925,N_33348);
or U35160 (N_35160,N_34269,N_34177);
nor U35161 (N_35161,N_33852,N_33148);
or U35162 (N_35162,N_34474,N_32687);
or U35163 (N_35163,N_32577,N_34560);
and U35164 (N_35164,N_34344,N_34200);
nor U35165 (N_35165,N_34985,N_34014);
or U35166 (N_35166,N_34189,N_33116);
nor U35167 (N_35167,N_34156,N_34725);
nor U35168 (N_35168,N_34505,N_34570);
nand U35169 (N_35169,N_34828,N_34598);
nor U35170 (N_35170,N_34497,N_34463);
and U35171 (N_35171,N_33568,N_33127);
nor U35172 (N_35172,N_33195,N_32692);
or U35173 (N_35173,N_33527,N_34504);
and U35174 (N_35174,N_33170,N_33228);
nor U35175 (N_35175,N_33207,N_33803);
nor U35176 (N_35176,N_32672,N_34703);
and U35177 (N_35177,N_34328,N_32796);
or U35178 (N_35178,N_33506,N_34358);
nor U35179 (N_35179,N_32831,N_33546);
and U35180 (N_35180,N_33885,N_34579);
nor U35181 (N_35181,N_33842,N_33942);
and U35182 (N_35182,N_32641,N_32628);
nor U35183 (N_35183,N_33768,N_34043);
and U35184 (N_35184,N_33355,N_34138);
nand U35185 (N_35185,N_34027,N_34960);
nand U35186 (N_35186,N_33090,N_34133);
nand U35187 (N_35187,N_34478,N_33653);
xor U35188 (N_35188,N_33379,N_33104);
xnor U35189 (N_35189,N_34275,N_33114);
or U35190 (N_35190,N_33759,N_32869);
nand U35191 (N_35191,N_34257,N_33821);
nor U35192 (N_35192,N_33323,N_34072);
nand U35193 (N_35193,N_32645,N_34173);
or U35194 (N_35194,N_32974,N_34729);
xnor U35195 (N_35195,N_33383,N_33514);
and U35196 (N_35196,N_34583,N_32584);
or U35197 (N_35197,N_34206,N_34340);
nand U35198 (N_35198,N_34185,N_33970);
nor U35199 (N_35199,N_33573,N_33824);
and U35200 (N_35200,N_34952,N_33306);
nand U35201 (N_35201,N_32519,N_34094);
nand U35202 (N_35202,N_33049,N_33697);
or U35203 (N_35203,N_32875,N_34170);
nor U35204 (N_35204,N_34851,N_34240);
and U35205 (N_35205,N_34355,N_32905);
or U35206 (N_35206,N_33928,N_33301);
or U35207 (N_35207,N_33205,N_32714);
and U35208 (N_35208,N_33143,N_33631);
xnor U35209 (N_35209,N_32781,N_32654);
xor U35210 (N_35210,N_34905,N_34372);
or U35211 (N_35211,N_34529,N_33564);
nor U35212 (N_35212,N_34466,N_32830);
nand U35213 (N_35213,N_34741,N_33182);
nor U35214 (N_35214,N_32684,N_33089);
nor U35215 (N_35215,N_32818,N_32801);
nand U35216 (N_35216,N_32921,N_34973);
and U35217 (N_35217,N_32842,N_33720);
nor U35218 (N_35218,N_33414,N_32721);
nand U35219 (N_35219,N_33196,N_34511);
nand U35220 (N_35220,N_33423,N_34535);
nand U35221 (N_35221,N_33023,N_34362);
and U35222 (N_35222,N_33979,N_33895);
nand U35223 (N_35223,N_33396,N_33464);
nand U35224 (N_35224,N_34589,N_33351);
nand U35225 (N_35225,N_33308,N_34689);
or U35226 (N_35226,N_34630,N_33218);
or U35227 (N_35227,N_33330,N_33889);
nor U35228 (N_35228,N_33751,N_34846);
and U35229 (N_35229,N_33727,N_32784);
nor U35230 (N_35230,N_34614,N_34139);
or U35231 (N_35231,N_33840,N_32623);
nor U35232 (N_35232,N_34272,N_33099);
nor U35233 (N_35233,N_33487,N_33336);
nand U35234 (N_35234,N_34752,N_33669);
nor U35235 (N_35235,N_33965,N_32566);
and U35236 (N_35236,N_32880,N_33359);
and U35237 (N_35237,N_32887,N_33990);
and U35238 (N_35238,N_34833,N_33562);
nor U35239 (N_35239,N_33031,N_32817);
xor U35240 (N_35240,N_34516,N_33643);
nand U35241 (N_35241,N_34942,N_34067);
and U35242 (N_35242,N_33934,N_34983);
or U35243 (N_35243,N_33713,N_33919);
xor U35244 (N_35244,N_33792,N_33482);
nand U35245 (N_35245,N_34684,N_34053);
nand U35246 (N_35246,N_34055,N_34410);
nand U35247 (N_35247,N_33696,N_32754);
nand U35248 (N_35248,N_34901,N_34397);
nor U35249 (N_35249,N_33134,N_33775);
or U35250 (N_35250,N_33316,N_33189);
and U35251 (N_35251,N_34544,N_34909);
nor U35252 (N_35252,N_33453,N_34595);
and U35253 (N_35253,N_33357,N_33743);
and U35254 (N_35254,N_32571,N_33053);
or U35255 (N_35255,N_34254,N_34754);
nor U35256 (N_35256,N_32546,N_34123);
nor U35257 (N_35257,N_33402,N_33377);
nand U35258 (N_35258,N_34515,N_32552);
or U35259 (N_35259,N_33113,N_33285);
or U35260 (N_35260,N_34884,N_34443);
nand U35261 (N_35261,N_33943,N_33929);
nor U35262 (N_35262,N_34022,N_33038);
xnor U35263 (N_35263,N_34719,N_34675);
and U35264 (N_35264,N_32624,N_33341);
nand U35265 (N_35265,N_33786,N_34314);
nor U35266 (N_35266,N_33866,N_32882);
and U35267 (N_35267,N_32849,N_34642);
and U35268 (N_35268,N_34639,N_34848);
nand U35269 (N_35269,N_33614,N_34187);
nand U35270 (N_35270,N_34708,N_33896);
xnor U35271 (N_35271,N_32522,N_33634);
xnor U35272 (N_35272,N_34099,N_33157);
and U35273 (N_35273,N_33244,N_33756);
or U35274 (N_35274,N_33796,N_34207);
nand U35275 (N_35275,N_33913,N_34870);
nand U35276 (N_35276,N_32524,N_34556);
xnor U35277 (N_35277,N_32728,N_34711);
nor U35278 (N_35278,N_34036,N_32550);
and U35279 (N_35279,N_34268,N_33365);
nand U35280 (N_35280,N_34062,N_32844);
nor U35281 (N_35281,N_34436,N_32924);
and U35282 (N_35282,N_34135,N_34769);
nor U35283 (N_35283,N_34955,N_32829);
or U35284 (N_35284,N_33045,N_33217);
and U35285 (N_35285,N_33447,N_34996);
xor U35286 (N_35286,N_33420,N_34750);
and U35287 (N_35287,N_33719,N_34374);
nor U35288 (N_35288,N_33654,N_34255);
or U35289 (N_35289,N_34256,N_32795);
nand U35290 (N_35290,N_33129,N_33125);
nor U35291 (N_35291,N_34124,N_34987);
nor U35292 (N_35292,N_34771,N_34959);
or U35293 (N_35293,N_34997,N_32711);
or U35294 (N_35294,N_32696,N_33015);
nor U35295 (N_35295,N_33467,N_34282);
or U35296 (N_35296,N_33788,N_34510);
or U35297 (N_35297,N_33040,N_33848);
nand U35298 (N_35298,N_32873,N_33804);
xor U35299 (N_35299,N_34449,N_34168);
and U35300 (N_35300,N_34659,N_32988);
nand U35301 (N_35301,N_32855,N_33960);
nand U35302 (N_35302,N_33378,N_33544);
nand U35303 (N_35303,N_33386,N_34112);
nor U35304 (N_35304,N_33732,N_32936);
and U35305 (N_35305,N_34707,N_32760);
nand U35306 (N_35306,N_34121,N_33297);
or U35307 (N_35307,N_33264,N_33112);
nand U35308 (N_35308,N_33173,N_32635);
nand U35309 (N_35309,N_34003,N_34477);
and U35310 (N_35310,N_34283,N_33644);
nor U35311 (N_35311,N_33374,N_32660);
or U35312 (N_35312,N_34047,N_34298);
nand U35313 (N_35313,N_34567,N_34161);
nand U35314 (N_35314,N_33474,N_33504);
xor U35315 (N_35315,N_32876,N_32860);
xor U35316 (N_35316,N_34486,N_34199);
or U35317 (N_35317,N_33128,N_34019);
or U35318 (N_35318,N_32607,N_34850);
or U35319 (N_35319,N_33662,N_34227);
or U35320 (N_35320,N_33448,N_34370);
nand U35321 (N_35321,N_34038,N_33789);
or U35322 (N_35322,N_33937,N_34231);
nor U35323 (N_35323,N_32528,N_32673);
nor U35324 (N_35324,N_34218,N_32720);
nor U35325 (N_35325,N_33594,N_32662);
nand U35326 (N_35326,N_32832,N_33836);
and U35327 (N_35327,N_34492,N_32854);
and U35328 (N_35328,N_32639,N_34437);
nand U35329 (N_35329,N_34748,N_32734);
and U35330 (N_35330,N_33741,N_34788);
or U35331 (N_35331,N_32906,N_34612);
or U35332 (N_35332,N_34333,N_33209);
nand U35333 (N_35333,N_34815,N_33718);
nand U35334 (N_35334,N_33176,N_32677);
nor U35335 (N_35335,N_32834,N_34976);
nor U35336 (N_35336,N_32920,N_32835);
nand U35337 (N_35337,N_34594,N_33999);
and U35338 (N_35338,N_34818,N_34318);
nor U35339 (N_35339,N_33253,N_34929);
nand U35340 (N_35340,N_33108,N_34366);
nor U35341 (N_35341,N_34115,N_33346);
and U35342 (N_35342,N_34380,N_33304);
and U35343 (N_35343,N_33621,N_34829);
nor U35344 (N_35344,N_34239,N_34383);
xnor U35345 (N_35345,N_32713,N_33291);
nor U35346 (N_35346,N_32858,N_33676);
or U35347 (N_35347,N_33597,N_32857);
nand U35348 (N_35348,N_34680,N_33476);
or U35349 (N_35349,N_32953,N_33438);
and U35350 (N_35350,N_34800,N_34445);
or U35351 (N_35351,N_32790,N_33811);
and U35352 (N_35352,N_32514,N_33488);
and U35353 (N_35353,N_33758,N_33622);
nor U35354 (N_35354,N_34702,N_34129);
or U35355 (N_35355,N_33295,N_32912);
nor U35356 (N_35356,N_33457,N_32787);
nand U35357 (N_35357,N_34651,N_32802);
or U35358 (N_35358,N_34302,N_32865);
and U35359 (N_35359,N_32966,N_34194);
nor U35360 (N_35360,N_33097,N_33313);
and U35361 (N_35361,N_33299,N_33080);
or U35362 (N_35362,N_34810,N_34709);
xnor U35363 (N_35363,N_33801,N_34456);
nand U35364 (N_35364,N_33695,N_33592);
or U35365 (N_35365,N_34202,N_34695);
and U35366 (N_35366,N_33007,N_34777);
and U35367 (N_35367,N_32710,N_32649);
and U35368 (N_35368,N_33335,N_32937);
nor U35369 (N_35369,N_32861,N_34487);
and U35370 (N_35370,N_33602,N_34414);
nand U35371 (N_35371,N_34245,N_34749);
nand U35372 (N_35372,N_34311,N_34611);
and U35373 (N_35373,N_33745,N_33156);
nor U35374 (N_35374,N_34162,N_33826);
or U35375 (N_35375,N_34285,N_32644);
nor U35376 (N_35376,N_33891,N_33034);
nand U35377 (N_35377,N_34806,N_33293);
xnor U35378 (N_35378,N_33973,N_34649);
or U35379 (N_35379,N_34877,N_34219);
and U35380 (N_35380,N_34667,N_33082);
nor U35381 (N_35381,N_33986,N_33589);
nand U35382 (N_35382,N_33110,N_33522);
nand U35383 (N_35383,N_33047,N_32658);
xnor U35384 (N_35384,N_33774,N_34444);
or U35385 (N_35385,N_33802,N_34731);
nor U35386 (N_35386,N_34369,N_33282);
and U35387 (N_35387,N_32957,N_32632);
nor U35388 (N_35388,N_33830,N_34382);
xnor U35389 (N_35389,N_33822,N_34032);
nand U35390 (N_35390,N_33779,N_34943);
or U35391 (N_35391,N_33729,N_32807);
nor U35392 (N_35392,N_32826,N_34982);
nor U35393 (N_35393,N_33035,N_34009);
nand U35394 (N_35394,N_33276,N_34224);
nor U35395 (N_35395,N_33724,N_34450);
and U35396 (N_35396,N_33003,N_34214);
and U35397 (N_35397,N_33581,N_34205);
and U35398 (N_35398,N_34034,N_34000);
nor U35399 (N_35399,N_33172,N_34106);
or U35400 (N_35400,N_32511,N_32812);
and U35401 (N_35401,N_33813,N_34839);
nor U35402 (N_35402,N_32777,N_34575);
or U35403 (N_35403,N_34826,N_32539);
and U35404 (N_35404,N_32567,N_33938);
and U35405 (N_35405,N_34937,N_32515);
and U35406 (N_35406,N_34817,N_32657);
or U35407 (N_35407,N_33871,N_33577);
or U35408 (N_35408,N_34704,N_34507);
nand U35409 (N_35409,N_34005,N_33685);
or U35410 (N_35410,N_34296,N_33927);
or U35411 (N_35411,N_32587,N_32706);
and U35412 (N_35412,N_32529,N_33410);
nand U35413 (N_35413,N_34706,N_34580);
nor U35414 (N_35414,N_33740,N_34863);
and U35415 (N_35415,N_34013,N_32910);
nor U35416 (N_35416,N_34367,N_33584);
xor U35417 (N_35417,N_34732,N_33735);
nor U35418 (N_35418,N_33851,N_33177);
or U35419 (N_35419,N_34520,N_33610);
xor U35420 (N_35420,N_34917,N_34419);
nand U35421 (N_35421,N_33909,N_34974);
nand U35422 (N_35422,N_33236,N_32883);
or U35423 (N_35423,N_33287,N_34151);
and U35424 (N_35424,N_34615,N_34095);
and U35425 (N_35425,N_34204,N_32568);
or U35426 (N_35426,N_34276,N_34136);
and U35427 (N_35427,N_34330,N_34048);
nand U35428 (N_35428,N_34315,N_34512);
and U35429 (N_35429,N_34883,N_32870);
nor U35430 (N_35430,N_33430,N_33325);
or U35431 (N_35431,N_33144,N_33778);
nand U35432 (N_35432,N_34564,N_34071);
and U35433 (N_35433,N_33632,N_32504);
nor U35434 (N_35434,N_34629,N_32680);
nor U35435 (N_35435,N_33615,N_32731);
and U35436 (N_35436,N_34002,N_34070);
or U35437 (N_35437,N_33419,N_34820);
or U35438 (N_35438,N_33923,N_34845);
nand U35439 (N_35439,N_33900,N_34572);
nor U35440 (N_35440,N_34687,N_33701);
nor U35441 (N_35441,N_32592,N_34113);
xor U35442 (N_35442,N_33946,N_33645);
nand U35443 (N_35443,N_33139,N_33363);
and U35444 (N_35444,N_32533,N_34809);
and U35445 (N_35445,N_34464,N_33808);
and U35446 (N_35446,N_33883,N_34323);
or U35447 (N_35447,N_33171,N_34710);
and U35448 (N_35448,N_34376,N_33041);
or U35449 (N_35449,N_33399,N_32888);
or U35450 (N_35450,N_34652,N_34503);
nor U35451 (N_35451,N_34496,N_34608);
nand U35452 (N_35452,N_32517,N_34554);
and U35453 (N_35453,N_34975,N_33070);
or U35454 (N_35454,N_34303,N_32960);
nand U35455 (N_35455,N_33650,N_34428);
nand U35456 (N_35456,N_34519,N_34781);
or U35457 (N_35457,N_33550,N_33843);
nor U35458 (N_35458,N_32556,N_34691);
nor U35459 (N_35459,N_32762,N_32554);
nor U35460 (N_35460,N_33454,N_33587);
or U35461 (N_35461,N_34084,N_33785);
or U35462 (N_35462,N_34600,N_34104);
xor U35463 (N_35463,N_33436,N_33232);
nor U35464 (N_35464,N_34670,N_34573);
or U35465 (N_35465,N_33307,N_33503);
and U35466 (N_35466,N_33899,N_34525);
nand U35467 (N_35467,N_34134,N_33265);
nand U35468 (N_35468,N_34881,N_32656);
and U35469 (N_35469,N_33771,N_32982);
or U35470 (N_35470,N_33255,N_33941);
nor U35471 (N_35471,N_32569,N_34647);
nand U35472 (N_35472,N_33569,N_32923);
and U35473 (N_35473,N_32836,N_34657);
nor U35474 (N_35474,N_34117,N_33032);
and U35475 (N_35475,N_34683,N_33625);
nor U35476 (N_35476,N_33936,N_34146);
nor U35477 (N_35477,N_34728,N_33582);
or U35478 (N_35478,N_34291,N_33305);
nand U35479 (N_35479,N_33096,N_34381);
or U35480 (N_35480,N_34216,N_34773);
and U35481 (N_35481,N_32997,N_32678);
and U35482 (N_35482,N_33426,N_33271);
or U35483 (N_35483,N_33017,N_34310);
or U35484 (N_35484,N_32708,N_34109);
and U35485 (N_35485,N_33598,N_34041);
or U35486 (N_35486,N_34483,N_33303);
nand U35487 (N_35487,N_32742,N_32823);
nor U35488 (N_35488,N_33094,N_32574);
and U35489 (N_35489,N_34501,N_34488);
nand U35490 (N_35490,N_33630,N_33208);
or U35491 (N_35491,N_33149,N_32686);
and U35492 (N_35492,N_32585,N_34932);
and U35493 (N_35493,N_33769,N_33640);
or U35494 (N_35494,N_34234,N_33048);
or U35495 (N_35495,N_32596,N_33543);
nand U35496 (N_35496,N_33284,N_34423);
nor U35497 (N_35497,N_32984,N_34727);
or U35498 (N_35498,N_32621,N_33797);
and U35499 (N_35499,N_33607,N_34927);
and U35500 (N_35500,N_33400,N_33969);
or U35501 (N_35501,N_33628,N_34637);
nand U35502 (N_35502,N_34609,N_32681);
nor U35503 (N_35503,N_34837,N_33715);
or U35504 (N_35504,N_34966,N_32916);
nor U35505 (N_35505,N_34541,N_32946);
and U35506 (N_35506,N_32676,N_33794);
or U35507 (N_35507,N_33138,N_32989);
nand U35508 (N_35508,N_32848,N_34857);
or U35509 (N_35509,N_32540,N_34455);
nor U35510 (N_35510,N_33352,N_32768);
xor U35511 (N_35511,N_32977,N_34838);
nor U35512 (N_35512,N_32951,N_33187);
xnor U35513 (N_35513,N_34890,N_32846);
nand U35514 (N_35514,N_34287,N_33130);
nand U35515 (N_35515,N_33269,N_32616);
nand U35516 (N_35516,N_32845,N_33052);
and U35517 (N_35517,N_33491,N_32881);
nor U35518 (N_35518,N_34791,N_32682);
nor U35519 (N_35519,N_33121,N_33525);
nand U35520 (N_35520,N_34694,N_34401);
or U35521 (N_35521,N_33256,N_34054);
or U35522 (N_35522,N_33100,N_33407);
xor U35523 (N_35523,N_33626,N_32987);
and U35524 (N_35524,N_32992,N_33555);
xor U35525 (N_35525,N_33219,N_34764);
nor U35526 (N_35526,N_34582,N_34348);
nor U35527 (N_35527,N_33202,N_34228);
xor U35528 (N_35528,N_33518,N_34517);
or U35529 (N_35529,N_33688,N_32985);
nand U35530 (N_35530,N_33993,N_34237);
nor U35531 (N_35531,N_33499,N_34776);
nand U35532 (N_35532,N_33155,N_33828);
xor U35533 (N_35533,N_34778,N_32611);
or U35534 (N_35534,N_33914,N_32652);
or U35535 (N_35535,N_33780,N_33234);
nor U35536 (N_35536,N_33066,N_32890);
and U35537 (N_35537,N_34337,N_32904);
nor U35538 (N_35538,N_32549,N_32914);
and U35539 (N_35539,N_33437,N_33194);
and U35540 (N_35540,N_33019,N_33327);
xnor U35541 (N_35541,N_33726,N_33263);
nor U35542 (N_35542,N_33318,N_34092);
xor U35543 (N_35543,N_33548,N_34499);
nor U35544 (N_35544,N_34063,N_34832);
nand U35545 (N_35545,N_32573,N_33215);
nor U35546 (N_35546,N_32748,N_34441);
nor U35547 (N_35547,N_33705,N_34169);
or U35548 (N_35548,N_34882,N_32646);
nand U35549 (N_35549,N_34968,N_34465);
or U35550 (N_35550,N_33672,N_33167);
and U35551 (N_35551,N_33526,N_34253);
nand U35552 (N_35552,N_33286,N_32638);
nand U35553 (N_35553,N_33747,N_34656);
or U35554 (N_35554,N_34258,N_33440);
or U35555 (N_35555,N_32627,N_33572);
or U35556 (N_35556,N_32694,N_33043);
nor U35557 (N_35557,N_34945,N_34980);
nand U35558 (N_35558,N_34087,N_34797);
nor U35559 (N_35559,N_33412,N_33190);
and U35560 (N_35560,N_34713,N_32782);
and U35561 (N_35561,N_34290,N_33507);
nor U35562 (N_35562,N_33545,N_34485);
nor U35563 (N_35563,N_34078,N_33971);
nor U35564 (N_35564,N_33289,N_34673);
xnor U35565 (N_35565,N_33509,N_34946);
and U35566 (N_35566,N_32944,N_34892);
nor U35567 (N_35567,N_32939,N_33905);
nor U35568 (N_35568,N_32756,N_32633);
xor U35569 (N_35569,N_33721,N_33575);
nand U35570 (N_35570,N_33441,N_34762);
nand U35571 (N_35571,N_34415,N_33337);
nor U35572 (N_35572,N_32968,N_32723);
nor U35573 (N_35573,N_34559,N_33549);
or U35574 (N_35574,N_33434,N_32779);
xor U35575 (N_35575,N_34182,N_33033);
nor U35576 (N_35576,N_33483,N_34605);
xor U35577 (N_35577,N_34876,N_34172);
nor U35578 (N_35578,N_33339,N_34077);
nand U35579 (N_35579,N_34011,N_34830);
nand U35580 (N_35580,N_34803,N_33838);
or U35581 (N_35581,N_34165,N_34213);
and U35582 (N_35582,N_34549,N_34603);
or U35583 (N_35583,N_33508,N_32561);
or U35584 (N_35584,N_32931,N_33921);
or U35585 (N_35585,N_34500,N_34664);
and U35586 (N_35586,N_34387,N_34180);
or U35587 (N_35587,N_34743,N_34016);
or U35588 (N_35588,N_33331,N_33312);
or U35589 (N_35589,N_34304,N_32954);
nor U35590 (N_35590,N_33036,N_33012);
and U35591 (N_35591,N_34020,N_33930);
or U35592 (N_35592,N_34714,N_33652);
or U35593 (N_35593,N_33324,N_32520);
or U35594 (N_35594,N_34530,N_34783);
nand U35595 (N_35595,N_33061,N_34451);
nor U35596 (N_35596,N_34532,N_33558);
nand U35597 (N_35597,N_33570,N_33523);
nand U35598 (N_35598,N_33897,N_33893);
nand U35599 (N_35599,N_34753,N_33933);
nor U35600 (N_35600,N_32770,N_33465);
or U35601 (N_35601,N_32964,N_34962);
or U35602 (N_35602,N_34430,N_32816);
nand U35603 (N_35603,N_34508,N_33733);
and U35604 (N_35604,N_33485,N_34385);
or U35605 (N_35605,N_34015,N_32772);
nor U35606 (N_35606,N_34969,N_33815);
nand U35607 (N_35607,N_32773,N_32575);
or U35608 (N_35608,N_33704,N_32794);
nand U35609 (N_35609,N_34150,N_34823);
or U35610 (N_35610,N_32879,N_34804);
nand U35611 (N_35611,N_34425,N_33898);
nand U35612 (N_35612,N_33425,N_34457);
and U35613 (N_35613,N_33008,N_33903);
and U35614 (N_35614,N_33473,N_34396);
nand U35615 (N_35615,N_33799,N_33908);
nand U35616 (N_35616,N_32808,N_34954);
xor U35617 (N_35617,N_34599,N_34127);
or U35618 (N_35618,N_32971,N_34058);
xor U35619 (N_35619,N_34666,N_34574);
or U35620 (N_35620,N_33422,N_32928);
xor U35621 (N_35621,N_34389,N_33831);
and U35622 (N_35622,N_34644,N_34331);
nand U35623 (N_35623,N_32769,N_34842);
or U35624 (N_35624,N_34264,N_34744);
nand U35625 (N_35625,N_34558,N_32862);
or U35626 (N_35626,N_33590,N_32562);
or U35627 (N_35627,N_33554,N_33798);
or U35628 (N_35628,N_33725,N_33517);
nor U35629 (N_35629,N_32588,N_32800);
nor U35630 (N_35630,N_33342,N_34225);
and U35631 (N_35631,N_34875,N_33078);
nor U35632 (N_35632,N_32851,N_32541);
and U35633 (N_35633,N_33180,N_34440);
and U35634 (N_35634,N_33216,N_33761);
nor U35635 (N_35635,N_33120,N_32739);
xnor U35636 (N_35636,N_34346,N_33950);
nor U35637 (N_35637,N_32600,N_34352);
and U35638 (N_35638,N_33677,N_33141);
or U35639 (N_35639,N_34160,N_33757);
and U35640 (N_35640,N_34509,N_33384);
or U35641 (N_35641,N_33781,N_34393);
or U35642 (N_35642,N_32542,N_34825);
and U35643 (N_35643,N_32792,N_33262);
nand U35644 (N_35644,N_33459,N_34193);
nand U35645 (N_35645,N_34855,N_33578);
xnor U35646 (N_35646,N_34633,N_34196);
nor U35647 (N_35647,N_34548,N_33206);
and U35648 (N_35648,N_34970,N_32747);
or U35649 (N_35649,N_33460,N_32634);
nor U35650 (N_35650,N_33372,N_34634);
nand U35651 (N_35651,N_32942,N_33707);
nor U35652 (N_35652,N_32523,N_32819);
xor U35653 (N_35653,N_34050,N_33730);
nand U35654 (N_35654,N_33261,N_33484);
or U35655 (N_35655,N_32558,N_33131);
nor U35656 (N_35656,N_33468,N_34956);
nand U35657 (N_35657,N_33663,N_33408);
nor U35658 (N_35658,N_34433,N_34226);
nor U35659 (N_35659,N_33535,N_33178);
or U35660 (N_35660,N_34601,N_32689);
nor U35661 (N_35661,N_33201,N_34171);
or U35662 (N_35662,N_32941,N_34722);
nor U35663 (N_35663,N_32841,N_33223);
nand U35664 (N_35664,N_34834,N_32507);
nor U35665 (N_35665,N_33841,N_34992);
or U35666 (N_35666,N_33037,N_33181);
and U35667 (N_35667,N_33832,N_32935);
nand U35668 (N_35668,N_32994,N_33661);
nor U35669 (N_35669,N_32553,N_34375);
xor U35670 (N_35670,N_34587,N_34964);
nand U35671 (N_35671,N_33381,N_33500);
and U35672 (N_35672,N_34083,N_33559);
nor U35673 (N_35673,N_33079,N_34064);
nand U35674 (N_35674,N_32810,N_34920);
xnor U35675 (N_35675,N_34244,N_34958);
nand U35676 (N_35676,N_34782,N_33480);
nor U35677 (N_35677,N_32981,N_32895);
nand U35678 (N_35678,N_34057,N_33557);
or U35679 (N_35679,N_33119,N_33619);
nand U35680 (N_35680,N_34990,N_34765);
nor U35681 (N_35681,N_33446,N_34175);
nand U35682 (N_35682,N_34911,N_33823);
nor U35683 (N_35683,N_33226,N_32629);
nand U35684 (N_35684,N_34787,N_34363);
nor U35685 (N_35685,N_34447,N_33783);
and U35686 (N_35686,N_34413,N_33000);
nor U35687 (N_35687,N_33878,N_32962);
nand U35688 (N_35688,N_34052,N_34212);
and U35689 (N_35689,N_34852,N_34999);
nor U35690 (N_35690,N_32753,N_32525);
nand U35691 (N_35691,N_32986,N_33537);
or U35692 (N_35692,N_33975,N_33877);
and U35693 (N_35693,N_33056,N_33338);
nor U35694 (N_35694,N_34844,N_34720);
or U35695 (N_35695,N_34931,N_33489);
and U35696 (N_35696,N_33225,N_33411);
and U35697 (N_35697,N_33162,N_34467);
and U35698 (N_35698,N_33071,N_33524);
nor U35699 (N_35699,N_33067,N_33101);
nor U35700 (N_35700,N_32863,N_34768);
or U35701 (N_35701,N_34533,N_33493);
nor U35702 (N_35702,N_32602,N_32530);
and U35703 (N_35703,N_34181,N_33463);
nor U35704 (N_35704,N_33039,N_32669);
or U35705 (N_35705,N_33606,N_33911);
and U35706 (N_35706,N_33321,N_34007);
nand U35707 (N_35707,N_34220,N_34326);
or U35708 (N_35708,N_32809,N_33340);
nor U35709 (N_35709,N_33309,N_34551);
or U35710 (N_35710,N_33490,N_34550);
or U35711 (N_35711,N_33268,N_32940);
or U35712 (N_35712,N_32647,N_34325);
nand U35713 (N_35713,N_34035,N_34324);
and U35714 (N_35714,N_32651,N_33717);
nand U35715 (N_35715,N_32663,N_33648);
or U35716 (N_35716,N_32852,N_33275);
xor U35717 (N_35717,N_33020,N_32730);
nor U35718 (N_35718,N_32788,N_34452);
nor U35719 (N_35719,N_32838,N_33817);
nor U35720 (N_35720,N_34918,N_33637);
or U35721 (N_35721,N_34868,N_32709);
and U35722 (N_35722,N_32679,N_34357);
nand U35723 (N_35723,N_33166,N_34902);
nor U35724 (N_35724,N_34658,N_33140);
nor U35725 (N_35725,N_33394,N_32544);
nand U35726 (N_35726,N_32837,N_33088);
nor U35727 (N_35727,N_33687,N_34494);
nor U35728 (N_35728,N_33748,N_34737);
nand U35729 (N_35729,N_33389,N_34665);
or U35730 (N_35730,N_34701,N_33270);
or U35731 (N_35731,N_32591,N_33764);
nor U35732 (N_35732,N_34977,N_34307);
and U35733 (N_35733,N_32671,N_33095);
nor U35734 (N_35734,N_32589,N_34319);
or U35735 (N_35735,N_33179,N_34641);
nand U35736 (N_35736,N_34915,N_33492);
xor U35737 (N_35737,N_33784,N_32615);
nor U35738 (N_35738,N_33298,N_32963);
and U35739 (N_35739,N_33371,N_34733);
and U35740 (N_35740,N_32776,N_32697);
xor U35741 (N_35741,N_32811,N_33686);
and U35742 (N_35742,N_33556,N_33317);
nor U35743 (N_35743,N_33174,N_32700);
or U35744 (N_35744,N_32900,N_33888);
nand U35745 (N_35745,N_34526,N_33887);
nor U35746 (N_35746,N_33773,N_33433);
and U35747 (N_35747,N_33700,N_34394);
nor U35748 (N_35748,N_34184,N_34557);
nor U35749 (N_35749,N_34965,N_33087);
and U35750 (N_35750,N_32969,N_33380);
nor U35751 (N_35751,N_32793,N_34312);
nor U35752 (N_35752,N_33002,N_33940);
and U35753 (N_35753,N_34607,N_33563);
and U35754 (N_35754,N_32565,N_34668);
xnor U35755 (N_35755,N_33693,N_33240);
or U35756 (N_35756,N_34894,N_32537);
nor U35757 (N_35757,N_32978,N_34025);
or U35758 (N_35758,N_33579,N_32501);
nand U35759 (N_35759,N_32665,N_34984);
and U35760 (N_35760,N_33599,N_33501);
and U35761 (N_35761,N_33833,N_34893);
and U35762 (N_35762,N_32740,N_33989);
or U35763 (N_35763,N_34552,N_33314);
xor U35764 (N_35764,N_32659,N_32625);
nor U35765 (N_35765,N_34001,N_33984);
nor U35766 (N_35766,N_33220,N_32824);
or U35767 (N_35767,N_32593,N_33461);
and U35768 (N_35768,N_34577,N_34042);
and U35769 (N_35769,N_33392,N_34847);
nand U35770 (N_35770,N_34610,N_34010);
nand U35771 (N_35771,N_34628,N_34735);
nor U35772 (N_35772,N_33188,N_34033);
nor U35773 (N_35773,N_34335,N_33185);
nor U35774 (N_35774,N_33026,N_34926);
nand U35775 (N_35775,N_33118,N_33846);
or U35776 (N_35776,N_33541,N_34399);
nor U35777 (N_35777,N_33706,N_34154);
or U35778 (N_35778,N_33870,N_34576);
nor U35779 (N_35779,N_33825,N_33671);
or U35780 (N_35780,N_33699,N_33519);
or U35781 (N_35781,N_33875,N_34137);
nor U35782 (N_35782,N_33200,N_33063);
or U35783 (N_35783,N_32560,N_33560);
nand U35784 (N_35784,N_34297,N_33710);
or U35785 (N_35785,N_34232,N_32722);
and U35786 (N_35786,N_33961,N_34097);
and U35787 (N_35787,N_32535,N_34306);
and U35788 (N_35788,N_34531,N_34715);
or U35789 (N_35789,N_34403,N_34091);
nor U35790 (N_35790,N_32674,N_33249);
xor U35791 (N_35791,N_33987,N_33947);
or U35792 (N_35792,N_32518,N_33266);
and U35793 (N_35793,N_34645,N_32610);
or U35794 (N_35794,N_34469,N_33805);
and U35795 (N_35795,N_34329,N_33497);
xor U35796 (N_35796,N_33902,N_33029);
nand U35797 (N_35797,N_34471,N_34616);
nor U35798 (N_35798,N_32820,N_34947);
nand U35799 (N_35799,N_33245,N_34669);
nand U35800 (N_35800,N_34697,N_33651);
and U35801 (N_35801,N_34473,N_34412);
or U35802 (N_35802,N_33692,N_32712);
nand U35803 (N_35803,N_33081,N_32707);
xor U35804 (N_35804,N_33666,N_33334);
or U35805 (N_35805,N_34502,N_32943);
nor U35806 (N_35806,N_33588,N_33005);
and U35807 (N_35807,N_32871,N_34730);
and U35808 (N_35808,N_32785,N_34086);
and U35809 (N_35809,N_32743,N_34248);
or U35810 (N_35810,N_33449,N_33111);
and U35811 (N_35811,N_33322,N_33175);
nand U35812 (N_35812,N_33001,N_32949);
nor U35813 (N_35813,N_34049,N_33239);
nor U35814 (N_35814,N_33673,N_33442);
nand U35815 (N_35815,N_33624,N_34338);
nand U35816 (N_35816,N_32894,N_34046);
nor U35817 (N_35817,N_34472,N_33233);
or U35818 (N_35818,N_32840,N_33385);
nor U35819 (N_35819,N_33277,N_32856);
or U35820 (N_35820,N_34183,N_32548);
nor U35821 (N_35821,N_34546,N_33288);
nand U35822 (N_35822,N_32703,N_32693);
or U35823 (N_35823,N_33479,N_34069);
nor U35824 (N_35824,N_33098,N_33861);
and U35825 (N_35825,N_34354,N_34700);
nor U35826 (N_35826,N_34270,N_34807);
xor U35827 (N_35827,N_33812,N_34514);
and U35828 (N_35828,N_33243,N_34816);
or U35829 (N_35829,N_32893,N_32668);
or U35830 (N_35830,N_34862,N_33084);
nor U35831 (N_35831,N_33963,N_34592);
nand U35832 (N_35832,N_34479,N_33924);
and U35833 (N_35833,N_33613,N_34439);
nand U35834 (N_35834,N_33532,N_34018);
nand U35835 (N_35835,N_32877,N_33512);
xnor U35836 (N_35836,N_34085,N_32500);
or U35837 (N_35837,N_33418,N_33350);
or U35838 (N_35838,N_33976,N_33542);
nor U35839 (N_35839,N_33042,N_33347);
and U35840 (N_35840,N_33398,N_33886);
or U35841 (N_35841,N_34861,N_32661);
nor U35842 (N_35842,N_33450,N_33521);
or U35843 (N_35843,N_34361,N_33329);
and U35844 (N_35844,N_34662,N_33142);
nand U35845 (N_35845,N_33469,N_34278);
xnor U35846 (N_35846,N_34026,N_34261);
nor U35847 (N_35847,N_34763,N_33879);
nand U35848 (N_35848,N_33466,N_33683);
and U35849 (N_35849,N_33105,N_32886);
nor U35850 (N_35850,N_34195,N_32898);
xnor U35851 (N_35851,N_34949,N_34796);
nand U35852 (N_35852,N_33674,N_33534);
and U35853 (N_35853,N_34957,N_33868);
or U35854 (N_35854,N_34039,N_33332);
or U35855 (N_35855,N_33146,N_33547);
nor U35856 (N_35856,N_34045,N_34814);
nand U35857 (N_35857,N_32698,N_33657);
or U35858 (N_35858,N_33058,N_33230);
nand U35859 (N_35859,N_34470,N_34427);
or U35860 (N_35860,N_34650,N_33890);
nor U35861 (N_35861,N_33763,N_34646);
nor U35862 (N_35862,N_32922,N_33580);
nand U35863 (N_35863,N_33073,N_33591);
or U35864 (N_35864,N_34950,N_33193);
and U35865 (N_35865,N_33443,N_34409);
nor U35866 (N_35866,N_34860,N_34243);
nand U35867 (N_35867,N_32716,N_32685);
nand U35868 (N_35868,N_32631,N_33742);
nand U35869 (N_35869,N_32545,N_34998);
xnor U35870 (N_35870,N_33022,N_34886);
nand U35871 (N_35871,N_34102,N_32961);
nor U35872 (N_35872,N_34012,N_34819);
nor U35873 (N_35873,N_34534,N_32945);
xor U35874 (N_35874,N_34627,N_34840);
nand U35875 (N_35875,N_33062,N_32806);
or U35876 (N_35876,N_34373,N_34178);
xor U35877 (N_35877,N_32640,N_33791);
or U35878 (N_35878,N_32738,N_33880);
xnor U35879 (N_35879,N_34313,N_32637);
nand U35880 (N_35880,N_34766,N_33738);
nand U35881 (N_35881,N_34565,N_34429);
and U35882 (N_35882,N_32932,N_34420);
xor U35883 (N_35883,N_34671,N_33059);
xnor U35884 (N_35884,N_34878,N_34274);
nor U35885 (N_35885,N_32643,N_34068);
or U35886 (N_35886,N_34895,N_33922);
nor U35887 (N_35887,N_34760,N_32737);
nand U35888 (N_35888,N_32655,N_34524);
and U35889 (N_35889,N_34164,N_34739);
nor U35890 (N_35890,N_32586,N_33472);
nor U35891 (N_35891,N_33361,N_33122);
nor U35892 (N_35892,N_33290,N_34359);
nor U35893 (N_35893,N_33617,N_33511);
or U35894 (N_35894,N_32736,N_33762);
nor U35895 (N_35895,N_33168,N_33292);
xor U35896 (N_35896,N_33083,N_33714);
nand U35897 (N_35897,N_32521,N_34738);
or U35898 (N_35898,N_34149,N_34334);
nor U35899 (N_35899,N_32746,N_33151);
xor U35900 (N_35900,N_34780,N_33668);
xor U35901 (N_35901,N_34153,N_33945);
and U35902 (N_35902,N_34157,N_32908);
or U35903 (N_35903,N_32536,N_32815);
xnor U35904 (N_35904,N_34201,N_34215);
nand U35905 (N_35905,N_32917,N_33435);
nor U35906 (N_35906,N_34745,N_33405);
nor U35907 (N_35907,N_32699,N_33247);
nand U35908 (N_35908,N_33267,N_33367);
nor U35909 (N_35909,N_33882,N_33315);
nand U35910 (N_35910,N_33670,N_33702);
and U35911 (N_35911,N_32609,N_34368);
or U35912 (N_35912,N_34631,N_33126);
nand U35913 (N_35913,N_33595,N_34343);
xnor U35914 (N_35914,N_32557,N_33011);
xor U35915 (N_35915,N_33665,N_33533);
and U35916 (N_35916,N_33623,N_32874);
and U35917 (N_35917,N_33091,N_34263);
nand U35918 (N_35918,N_34571,N_33427);
nand U35919 (N_35919,N_33767,N_33075);
nand U35920 (N_35920,N_32688,N_34718);
or U35921 (N_35921,N_33360,N_32667);
nand U35922 (N_35922,N_34635,N_34827);
nor U35923 (N_35923,N_34989,N_34490);
and U35924 (N_35924,N_33241,N_33382);
nor U35925 (N_35925,N_33404,N_32744);
nor U35926 (N_35926,N_34093,N_34284);
or U35927 (N_35927,N_34148,N_34948);
and U35928 (N_35928,N_34621,N_32973);
nand U35929 (N_35929,N_33816,N_34247);
nand U35930 (N_35930,N_34390,N_34798);
or U35931 (N_35931,N_34756,N_34871);
nand U35932 (N_35932,N_32502,N_32799);
nor U35933 (N_35933,N_34251,N_34789);
nor U35934 (N_35934,N_32926,N_33857);
nand U35935 (N_35935,N_34342,N_33601);
nand U35936 (N_35936,N_32580,N_32763);
and U35937 (N_35937,N_33366,N_34995);
nand U35938 (N_35938,N_33656,N_34678);
and U35939 (N_35939,N_34935,N_32813);
nor U35940 (N_35940,N_34371,N_33133);
or U35941 (N_35941,N_33974,N_34940);
or U35942 (N_35942,N_33863,N_34082);
nor U35943 (N_35943,N_32718,N_34107);
nand U35944 (N_35944,N_34110,N_32683);
nand U35945 (N_35945,N_33538,N_32619);
nand U35946 (N_35946,N_33044,N_33213);
nor U35947 (N_35947,N_33603,N_32555);
or U35948 (N_35948,N_33057,N_34939);
and U35949 (N_35949,N_32998,N_33496);
nand U35950 (N_35950,N_34065,N_34103);
and U35951 (N_35951,N_34888,N_33873);
nor U35952 (N_35952,N_34543,N_32929);
and U35953 (N_35953,N_34453,N_33782);
xor U35954 (N_35954,N_33977,N_33703);
or U35955 (N_35955,N_34417,N_32531);
or U35956 (N_35956,N_33137,N_33354);
nor U35957 (N_35957,N_34794,N_33565);
xnor U35958 (N_35958,N_33722,N_33892);
and U35959 (N_35959,N_34286,N_33163);
and U35960 (N_35960,N_33867,N_32843);
nor U35961 (N_35961,N_33106,N_34098);
or U35962 (N_35962,N_32650,N_33154);
or U35963 (N_35963,N_33995,N_33085);
and U35964 (N_35964,N_34347,N_33736);
and U35965 (N_35965,N_33608,N_34604);
or U35966 (N_35966,N_34217,N_33345);
and U35967 (N_35967,N_33051,N_34392);
or U35968 (N_35968,N_34044,N_33030);
nand U35969 (N_35969,N_33158,N_34712);
nand U35970 (N_35970,N_33616,N_33531);
nand U35971 (N_35971,N_32579,N_34259);
nand U35972 (N_35972,N_32617,N_33406);
xor U35973 (N_35973,N_32653,N_33574);
xnor U35974 (N_35974,N_33165,N_33403);
nand U35975 (N_35975,N_33997,N_34682);
or U35976 (N_35976,N_34681,N_34209);
nor U35977 (N_35977,N_32725,N_33855);
nand U35978 (N_35978,N_32915,N_33874);
nand U35979 (N_35979,N_34030,N_33917);
nand U35980 (N_35980,N_33439,N_32532);
xor U35981 (N_35981,N_33869,N_32938);
xnor U35982 (N_35982,N_32789,N_34620);
nand U35983 (N_35983,N_34655,N_32729);
and U35984 (N_35984,N_34434,N_34853);
and U35985 (N_35985,N_33432,N_34482);
and U35986 (N_35986,N_34407,N_33800);
nor U35987 (N_35987,N_33920,N_33739);
and U35988 (N_35988,N_34322,N_34916);
and U35989 (N_35989,N_34405,N_34203);
nor U35990 (N_35990,N_32750,N_34924);
or U35991 (N_35991,N_33009,N_33021);
or U35992 (N_35992,N_34978,N_33991);
or U35993 (N_35993,N_34879,N_32948);
nor U35994 (N_35994,N_34061,N_33102);
nand U35995 (N_35995,N_33684,N_33765);
nand U35996 (N_35996,N_34365,N_33281);
or U35997 (N_35997,N_33907,N_32884);
xnor U35998 (N_35998,N_33018,N_33115);
and U35999 (N_35999,N_34578,N_33996);
nor U36000 (N_36000,N_33221,N_33214);
or U36001 (N_36001,N_33658,N_34364);
xnor U36002 (N_36002,N_34398,N_33429);
nand U36003 (N_36003,N_33820,N_32783);
nand U36004 (N_36004,N_33376,N_33939);
nor U36005 (N_36005,N_33709,N_33636);
nor U36006 (N_36006,N_34416,N_32597);
nand U36007 (N_36007,N_34400,N_33197);
or U36008 (N_36008,N_34770,N_34294);
or U36009 (N_36009,N_34190,N_33495);
and U36010 (N_36010,N_32551,N_34152);
nor U36011 (N_36011,N_34619,N_34271);
and U36012 (N_36012,N_34353,N_32901);
nor U36013 (N_36013,N_32798,N_32538);
nand U36014 (N_36014,N_34379,N_32581);
xnor U36015 (N_36015,N_33723,N_34114);
nand U36016 (N_36016,N_34912,N_33810);
or U36017 (N_36017,N_32913,N_34066);
or U36018 (N_36018,N_34468,N_33711);
and U36019 (N_36019,N_34891,N_33760);
nor U36020 (N_36020,N_33664,N_34568);
or U36021 (N_36021,N_34606,N_32774);
nand U36022 (N_36022,N_33424,N_32534);
nor U36023 (N_36023,N_33477,N_34236);
or U36024 (N_36024,N_33025,N_33528);
nand U36025 (N_36025,N_34747,N_32508);
xnor U36026 (N_36026,N_34677,N_33829);
xor U36027 (N_36027,N_34246,N_33901);
xor U36028 (N_36028,N_33198,N_34351);
nand U36029 (N_36029,N_33458,N_33835);
and U36030 (N_36030,N_34721,N_33283);
and U36031 (N_36031,N_32814,N_33147);
xor U36032 (N_36032,N_33444,N_34233);
xor U36033 (N_36033,N_34079,N_33837);
nor U36034 (N_36034,N_34793,N_33356);
nand U36035 (N_36035,N_32952,N_33224);
nand U36036 (N_36036,N_32903,N_34904);
or U36037 (N_36037,N_33152,N_33373);
or U36038 (N_36038,N_33959,N_34705);
nand U36039 (N_36039,N_34872,N_33766);
or U36040 (N_36040,N_33238,N_34422);
nand U36041 (N_36041,N_33478,N_33680);
and U36042 (N_36042,N_34462,N_32604);
nand U36043 (N_36043,N_32735,N_33010);
nand U36044 (N_36044,N_33916,N_34301);
or U36045 (N_36045,N_33931,N_34384);
nand U36046 (N_36046,N_34547,N_33065);
nor U36047 (N_36047,N_33103,N_33967);
nor U36048 (N_36048,N_34685,N_33428);
nor U36049 (N_36049,N_34125,N_34120);
nand U36050 (N_36050,N_34418,N_32724);
and U36051 (N_36051,N_33847,N_32970);
nand U36052 (N_36052,N_34391,N_34059);
or U36053 (N_36053,N_33183,N_33862);
xnor U36054 (N_36054,N_33387,N_33536);
or U36055 (N_36055,N_33731,N_32975);
xnor U36056 (N_36056,N_34446,N_32918);
or U36057 (N_36057,N_33675,N_33222);
xor U36058 (N_36058,N_34080,N_32576);
nor U36059 (N_36059,N_34538,N_33375);
xnor U36060 (N_36060,N_34299,N_34438);
nand U36061 (N_36061,N_34223,N_34971);
nor U36062 (N_36062,N_34260,N_33834);
xor U36063 (N_36063,N_32618,N_33074);
or U36064 (N_36064,N_34991,N_34105);
nor U36065 (N_36065,N_33451,N_33953);
or U36066 (N_36066,N_34923,N_34921);
and U36067 (N_36067,N_33413,N_34843);
nor U36068 (N_36068,N_33849,N_34596);
xnor U36069 (N_36069,N_33844,N_32717);
and U36070 (N_36070,N_33754,N_34432);
nand U36071 (N_36071,N_34540,N_34167);
xor U36072 (N_36072,N_34088,N_32719);
or U36073 (N_36073,N_33600,N_34617);
nor U36074 (N_36074,N_33161,N_33054);
nand U36075 (N_36075,N_34179,N_33689);
xor U36076 (N_36076,N_32892,N_34919);
and U36077 (N_36077,N_33169,N_34308);
and U36078 (N_36078,N_32715,N_33250);
and U36079 (N_36079,N_32956,N_33028);
nor U36080 (N_36080,N_33814,N_32570);
and U36081 (N_36081,N_34686,N_33364);
nor U36082 (N_36082,N_34475,N_33647);
nand U36083 (N_36083,N_34698,N_33633);
nand U36084 (N_36084,N_33358,N_33192);
nand U36085 (N_36085,N_33609,N_34640);
and U36086 (N_36086,N_32559,N_34489);
and U36087 (N_36087,N_34528,N_34938);
and U36088 (N_36088,N_34654,N_34021);
nor U36089 (N_36089,N_33915,N_33964);
nand U36090 (N_36090,N_34459,N_33744);
nand U36091 (N_36091,N_34835,N_34986);
xnor U36092 (N_36092,N_34914,N_34192);
nand U36093 (N_36093,N_32958,N_34075);
nand U36094 (N_36094,N_33445,N_33708);
and U36095 (N_36095,N_34746,N_34506);
nand U36096 (N_36096,N_32850,N_33948);
and U36097 (N_36097,N_33300,N_34887);
or U36098 (N_36098,N_33858,N_34090);
nor U36099 (N_36099,N_34792,N_34111);
nand U36100 (N_36100,N_33850,N_33455);
nor U36101 (N_36101,N_34581,N_32991);
and U36102 (N_36102,N_33237,N_34252);
nor U36103 (N_36103,N_34460,N_32583);
and U36104 (N_36104,N_33320,N_33962);
nor U36105 (N_36105,N_33124,N_33184);
nand U36106 (N_36106,N_33678,N_33629);
xnor U36107 (N_36107,N_33982,N_33859);
and U36108 (N_36108,N_34779,N_34584);
and U36109 (N_36109,N_33571,N_32919);
or U36110 (N_36110,N_33772,N_33160);
nand U36111 (N_36111,N_34360,N_33691);
nor U36112 (N_36112,N_34775,N_32695);
nor U36113 (N_36113,N_34910,N_34813);
nor U36114 (N_36114,N_34913,N_34332);
and U36115 (N_36115,N_34144,N_33248);
nand U36116 (N_36116,N_33978,N_33415);
or U36117 (N_36117,N_33132,N_34933);
or U36118 (N_36118,N_34994,N_33881);
nor U36119 (N_36119,N_34626,N_33593);
and U36120 (N_36120,N_33145,N_33649);
nand U36121 (N_36121,N_32690,N_33516);
or U36122 (N_36122,N_33328,N_33949);
nand U36123 (N_36123,N_34908,N_33605);
and U36124 (N_36124,N_34790,N_33682);
and U36125 (N_36125,N_34759,N_34454);
nand U36126 (N_36126,N_32594,N_33712);
xnor U36127 (N_36127,N_32595,N_33368);
and U36128 (N_36128,N_33274,N_34537);
and U36129 (N_36129,N_34785,N_33092);
or U36130 (N_36130,N_33107,N_34461);
nand U36131 (N_36131,N_34495,N_34040);
xor U36132 (N_36132,N_33968,N_34262);
and U36133 (N_36133,N_34724,N_34858);
nor U36134 (N_36134,N_33470,N_33077);
and U36135 (N_36135,N_33109,N_33627);
or U36136 (N_36136,N_34250,N_33349);
nand U36137 (N_36137,N_34869,N_34132);
or U36138 (N_36138,N_33698,N_33776);
nand U36139 (N_36139,N_32626,N_34222);
xor U36140 (N_36140,N_33046,N_34131);
or U36141 (N_36141,N_33076,N_33734);
nor U36142 (N_36142,N_34281,N_32805);
and U36143 (N_36143,N_32506,N_32606);
nand U36144 (N_36144,N_34238,N_34597);
and U36145 (N_36145,N_33004,N_34056);
or U36146 (N_36146,N_34350,N_34017);
nor U36147 (N_36147,N_34660,N_32839);
and U36148 (N_36148,N_33952,N_34191);
xnor U36149 (N_36149,N_34951,N_33257);
nor U36150 (N_36150,N_32803,N_34864);
nor U36151 (N_36151,N_33273,N_34555);
nor U36152 (N_36152,N_33498,N_34624);
nand U36153 (N_36153,N_32622,N_34411);
nand U36154 (N_36154,N_33752,N_34801);
nand U36155 (N_36155,N_33932,N_34941);
and U36156 (N_36156,N_33694,N_33333);
and U36157 (N_36157,N_32885,N_32930);
nand U36158 (N_36158,N_34147,N_32547);
xnor U36159 (N_36159,N_34906,N_34859);
nor U36160 (N_36160,N_32732,N_34341);
and U36161 (N_36161,N_32642,N_33294);
or U36162 (N_36162,N_33583,N_34553);
or U36163 (N_36163,N_34186,N_33204);
or U36164 (N_36164,N_32765,N_34491);
or U36165 (N_36165,N_32996,N_34408);
nand U36166 (N_36166,N_33981,N_32825);
or U36167 (N_36167,N_34811,N_33016);
and U36168 (N_36168,N_33983,N_33014);
or U36169 (N_36169,N_32745,N_34119);
or U36170 (N_36170,N_33254,N_32866);
xnor U36171 (N_36171,N_33229,N_34742);
nor U36172 (N_36172,N_32675,N_34688);
nand U36173 (N_36173,N_33576,N_33667);
nand U36174 (N_36174,N_34922,N_34155);
nor U36175 (N_36175,N_32804,N_32980);
xor U36176 (N_36176,N_34051,N_32821);
xnor U36177 (N_36177,N_33864,N_32513);
nor U36178 (N_36178,N_34339,N_34944);
or U36179 (N_36179,N_33471,N_32990);
or U36180 (N_36180,N_34008,N_33395);
nand U36181 (N_36181,N_33486,N_34267);
nand U36182 (N_36182,N_33251,N_32993);
or U36183 (N_36183,N_34288,N_34081);
and U36184 (N_36184,N_34421,N_34378);
or U36185 (N_36185,N_34321,N_34643);
nand U36186 (N_36186,N_32582,N_34143);
or U36187 (N_36187,N_32853,N_33530);
xor U36188 (N_36188,N_33955,N_34141);
or U36189 (N_36189,N_32757,N_32613);
nor U36190 (N_36190,N_33806,N_34899);
or U36191 (N_36191,N_32979,N_33013);
and U36192 (N_36192,N_34448,N_34327);
nand U36193 (N_36193,N_32955,N_32902);
nand U36194 (N_36194,N_34866,N_34300);
nand U36195 (N_36195,N_33259,N_33641);
nand U36196 (N_36196,N_32822,N_33750);
nor U36197 (N_36197,N_33992,N_33655);
nor U36198 (N_36198,N_32704,N_32847);
nor U36199 (N_36199,N_33551,N_33540);
and U36200 (N_36200,N_33006,N_34130);
nand U36201 (N_36201,N_32601,N_32733);
nand U36202 (N_36202,N_33510,N_32727);
nand U36203 (N_36203,N_34108,N_33749);
nor U36204 (N_36204,N_34527,N_33416);
and U36205 (N_36205,N_33186,N_33296);
nand U36206 (N_36206,N_32995,N_33068);
and U36207 (N_36207,N_33456,N_32505);
nor U36208 (N_36208,N_34539,N_34885);
xor U36209 (N_36209,N_33951,N_34585);
and U36210 (N_36210,N_34767,N_34808);
or U36211 (N_36211,N_34266,N_34865);
nor U36212 (N_36212,N_34786,N_34277);
and U36213 (N_36213,N_34345,N_33790);
or U36214 (N_36214,N_34873,N_33737);
nor U36215 (N_36215,N_32572,N_32925);
or U36216 (N_36216,N_33343,N_33311);
and U36217 (N_36217,N_34736,N_33462);
nand U36218 (N_36218,N_33397,N_34211);
and U36219 (N_36219,N_34622,N_34854);
and U36220 (N_36220,N_32907,N_33539);
xnor U36221 (N_36221,N_34545,N_33086);
nor U36222 (N_36222,N_33279,N_34060);
xnor U36223 (N_36223,N_34166,N_34849);
or U36224 (N_36224,N_34761,N_33690);
nand U36225 (N_36225,N_33746,N_32758);
and U36226 (N_36226,N_33660,N_32563);
and U36227 (N_36227,N_32950,N_34122);
xor U36228 (N_36228,N_32608,N_32509);
nor U36229 (N_36229,N_33972,N_33926);
nor U36230 (N_36230,N_32999,N_34755);
nor U36231 (N_36231,N_34623,N_34089);
and U36232 (N_36232,N_34774,N_32691);
or U36233 (N_36233,N_34692,N_33280);
nand U36234 (N_36234,N_32664,N_34856);
nor U36235 (N_36235,N_34536,N_34198);
or U36236 (N_36236,N_34625,N_33417);
and U36237 (N_36237,N_34241,N_34498);
nor U36238 (N_36238,N_34221,N_34229);
nand U36239 (N_36239,N_33227,N_34476);
nor U36240 (N_36240,N_34602,N_33612);
nand U36241 (N_36241,N_34431,N_32859);
nand U36242 (N_36242,N_33093,N_33064);
and U36243 (N_36243,N_33502,N_33246);
and U36244 (N_36244,N_33060,N_33421);
and U36245 (N_36245,N_34805,N_33753);
xor U36246 (N_36246,N_34812,N_34934);
nor U36247 (N_36247,N_33777,N_34900);
or U36248 (N_36248,N_34988,N_33515);
nand U36249 (N_36249,N_33872,N_33860);
and U36250 (N_36250,N_34958,N_33466);
nor U36251 (N_36251,N_32905,N_34690);
nor U36252 (N_36252,N_33673,N_34416);
or U36253 (N_36253,N_33411,N_33651);
xnor U36254 (N_36254,N_32779,N_33861);
or U36255 (N_36255,N_33589,N_33577);
nor U36256 (N_36256,N_33309,N_34327);
nor U36257 (N_36257,N_32831,N_32837);
xor U36258 (N_36258,N_32802,N_32537);
or U36259 (N_36259,N_32664,N_33989);
or U36260 (N_36260,N_34697,N_34064);
nor U36261 (N_36261,N_34673,N_33529);
and U36262 (N_36262,N_33799,N_34112);
or U36263 (N_36263,N_32909,N_32807);
nor U36264 (N_36264,N_33069,N_32987);
and U36265 (N_36265,N_33982,N_32792);
or U36266 (N_36266,N_33293,N_34190);
and U36267 (N_36267,N_34059,N_34578);
xor U36268 (N_36268,N_33552,N_34771);
nand U36269 (N_36269,N_34698,N_33014);
nand U36270 (N_36270,N_33469,N_34945);
nand U36271 (N_36271,N_34354,N_34636);
nor U36272 (N_36272,N_34834,N_33321);
or U36273 (N_36273,N_34389,N_34760);
and U36274 (N_36274,N_33684,N_33319);
nor U36275 (N_36275,N_32812,N_33886);
or U36276 (N_36276,N_33636,N_32850);
and U36277 (N_36277,N_34816,N_32810);
nor U36278 (N_36278,N_34968,N_34503);
or U36279 (N_36279,N_34500,N_32676);
nor U36280 (N_36280,N_33698,N_33952);
and U36281 (N_36281,N_34419,N_34219);
nor U36282 (N_36282,N_33796,N_33411);
or U36283 (N_36283,N_32821,N_33189);
nor U36284 (N_36284,N_34934,N_33211);
and U36285 (N_36285,N_33881,N_34997);
or U36286 (N_36286,N_34582,N_33773);
nand U36287 (N_36287,N_33243,N_34890);
and U36288 (N_36288,N_34833,N_34296);
and U36289 (N_36289,N_32782,N_34914);
nor U36290 (N_36290,N_32953,N_32515);
and U36291 (N_36291,N_32556,N_33987);
nor U36292 (N_36292,N_32504,N_33478);
and U36293 (N_36293,N_34062,N_34033);
or U36294 (N_36294,N_34276,N_34751);
or U36295 (N_36295,N_32627,N_32592);
nand U36296 (N_36296,N_34116,N_33773);
nor U36297 (N_36297,N_33256,N_33049);
or U36298 (N_36298,N_33078,N_33945);
nor U36299 (N_36299,N_34354,N_33411);
or U36300 (N_36300,N_33173,N_33693);
xor U36301 (N_36301,N_33814,N_33294);
nand U36302 (N_36302,N_32953,N_34424);
nor U36303 (N_36303,N_33992,N_34752);
nor U36304 (N_36304,N_34724,N_32718);
nor U36305 (N_36305,N_33910,N_32772);
xnor U36306 (N_36306,N_34700,N_34912);
and U36307 (N_36307,N_33271,N_34784);
nor U36308 (N_36308,N_33746,N_33717);
nor U36309 (N_36309,N_34256,N_32587);
or U36310 (N_36310,N_32979,N_33997);
nor U36311 (N_36311,N_33386,N_33758);
or U36312 (N_36312,N_34854,N_32934);
nand U36313 (N_36313,N_33456,N_34316);
nand U36314 (N_36314,N_34322,N_34791);
nor U36315 (N_36315,N_34448,N_34467);
or U36316 (N_36316,N_32544,N_33294);
or U36317 (N_36317,N_32526,N_34078);
or U36318 (N_36318,N_34809,N_33070);
xor U36319 (N_36319,N_34131,N_34192);
and U36320 (N_36320,N_33128,N_34033);
nand U36321 (N_36321,N_34217,N_34970);
xnor U36322 (N_36322,N_34862,N_34199);
or U36323 (N_36323,N_34848,N_33070);
and U36324 (N_36324,N_33799,N_33766);
nor U36325 (N_36325,N_34737,N_32762);
or U36326 (N_36326,N_34794,N_32644);
and U36327 (N_36327,N_32682,N_33968);
and U36328 (N_36328,N_33683,N_33110);
and U36329 (N_36329,N_32955,N_34120);
nor U36330 (N_36330,N_32925,N_33874);
nor U36331 (N_36331,N_32728,N_34739);
nand U36332 (N_36332,N_34538,N_32538);
and U36333 (N_36333,N_32740,N_34803);
nor U36334 (N_36334,N_32564,N_34957);
nor U36335 (N_36335,N_33922,N_34394);
and U36336 (N_36336,N_33274,N_34829);
nand U36337 (N_36337,N_34955,N_33488);
and U36338 (N_36338,N_33916,N_34521);
or U36339 (N_36339,N_34470,N_33818);
and U36340 (N_36340,N_34508,N_33399);
and U36341 (N_36341,N_33043,N_33798);
nor U36342 (N_36342,N_34727,N_32693);
and U36343 (N_36343,N_33211,N_34542);
nand U36344 (N_36344,N_34078,N_33624);
nor U36345 (N_36345,N_32740,N_34505);
nand U36346 (N_36346,N_34875,N_32657);
or U36347 (N_36347,N_34557,N_34547);
nand U36348 (N_36348,N_34269,N_34368);
and U36349 (N_36349,N_34269,N_34427);
nand U36350 (N_36350,N_33309,N_32554);
xor U36351 (N_36351,N_34455,N_33565);
and U36352 (N_36352,N_33966,N_34899);
and U36353 (N_36353,N_34385,N_33665);
nor U36354 (N_36354,N_33640,N_33251);
or U36355 (N_36355,N_34782,N_32564);
nand U36356 (N_36356,N_34086,N_33149);
nor U36357 (N_36357,N_33486,N_34170);
and U36358 (N_36358,N_32895,N_32511);
and U36359 (N_36359,N_34266,N_34836);
nor U36360 (N_36360,N_34876,N_34862);
nand U36361 (N_36361,N_33420,N_34596);
nand U36362 (N_36362,N_34008,N_33975);
nor U36363 (N_36363,N_33535,N_34673);
nand U36364 (N_36364,N_34324,N_33684);
nand U36365 (N_36365,N_33532,N_34280);
nor U36366 (N_36366,N_34984,N_32956);
nor U36367 (N_36367,N_34462,N_32944);
nand U36368 (N_36368,N_33916,N_33011);
nor U36369 (N_36369,N_34023,N_34510);
nand U36370 (N_36370,N_33365,N_33829);
and U36371 (N_36371,N_32525,N_33614);
nand U36372 (N_36372,N_34958,N_33848);
xnor U36373 (N_36373,N_34588,N_33972);
nor U36374 (N_36374,N_33800,N_34874);
and U36375 (N_36375,N_33355,N_33672);
and U36376 (N_36376,N_32847,N_33434);
and U36377 (N_36377,N_34372,N_33712);
nand U36378 (N_36378,N_32533,N_34384);
nor U36379 (N_36379,N_33162,N_33426);
or U36380 (N_36380,N_32584,N_34685);
nor U36381 (N_36381,N_34867,N_33810);
and U36382 (N_36382,N_34493,N_34668);
nor U36383 (N_36383,N_34657,N_33509);
nand U36384 (N_36384,N_32598,N_34896);
nand U36385 (N_36385,N_33742,N_33026);
or U36386 (N_36386,N_32999,N_34600);
nor U36387 (N_36387,N_34635,N_34433);
and U36388 (N_36388,N_34457,N_32957);
and U36389 (N_36389,N_32836,N_33907);
nand U36390 (N_36390,N_33961,N_34470);
xnor U36391 (N_36391,N_34196,N_34433);
nand U36392 (N_36392,N_33130,N_33934);
and U36393 (N_36393,N_34403,N_34991);
or U36394 (N_36394,N_33722,N_34325);
and U36395 (N_36395,N_33451,N_32956);
and U36396 (N_36396,N_34860,N_34531);
or U36397 (N_36397,N_32985,N_32786);
nand U36398 (N_36398,N_33432,N_33107);
or U36399 (N_36399,N_33091,N_32980);
and U36400 (N_36400,N_34822,N_34494);
xnor U36401 (N_36401,N_33622,N_33824);
nand U36402 (N_36402,N_33751,N_34923);
nor U36403 (N_36403,N_34300,N_33252);
nor U36404 (N_36404,N_34734,N_33393);
nand U36405 (N_36405,N_32524,N_34664);
and U36406 (N_36406,N_33489,N_33754);
and U36407 (N_36407,N_33600,N_34386);
nor U36408 (N_36408,N_32519,N_32607);
nand U36409 (N_36409,N_32589,N_33073);
nand U36410 (N_36410,N_34920,N_32575);
or U36411 (N_36411,N_34220,N_32693);
or U36412 (N_36412,N_34375,N_32601);
nor U36413 (N_36413,N_34328,N_33528);
nand U36414 (N_36414,N_34441,N_33514);
nand U36415 (N_36415,N_33045,N_32841);
or U36416 (N_36416,N_33418,N_32681);
xnor U36417 (N_36417,N_34850,N_34542);
xnor U36418 (N_36418,N_33441,N_34026);
nand U36419 (N_36419,N_33080,N_33848);
nand U36420 (N_36420,N_34434,N_32943);
nand U36421 (N_36421,N_34531,N_33792);
nor U36422 (N_36422,N_34076,N_34732);
nor U36423 (N_36423,N_32645,N_33156);
xnor U36424 (N_36424,N_33123,N_33365);
nor U36425 (N_36425,N_34786,N_34177);
nor U36426 (N_36426,N_33062,N_34690);
xor U36427 (N_36427,N_32625,N_33406);
nand U36428 (N_36428,N_34104,N_33886);
nor U36429 (N_36429,N_33571,N_34218);
or U36430 (N_36430,N_32958,N_34990);
nor U36431 (N_36431,N_33909,N_32546);
nor U36432 (N_36432,N_34341,N_33921);
nand U36433 (N_36433,N_34215,N_33704);
or U36434 (N_36434,N_34710,N_33309);
nand U36435 (N_36435,N_32942,N_33873);
xor U36436 (N_36436,N_33874,N_34170);
nand U36437 (N_36437,N_32748,N_33196);
nor U36438 (N_36438,N_32639,N_32699);
nand U36439 (N_36439,N_32627,N_33661);
nor U36440 (N_36440,N_33195,N_33786);
xor U36441 (N_36441,N_32926,N_32780);
nand U36442 (N_36442,N_34834,N_34614);
nor U36443 (N_36443,N_33057,N_33302);
nor U36444 (N_36444,N_33554,N_32963);
nor U36445 (N_36445,N_32779,N_34064);
xnor U36446 (N_36446,N_33898,N_33859);
nor U36447 (N_36447,N_33501,N_34693);
and U36448 (N_36448,N_34984,N_33950);
nand U36449 (N_36449,N_32703,N_34307);
nand U36450 (N_36450,N_34176,N_33644);
and U36451 (N_36451,N_34454,N_34896);
and U36452 (N_36452,N_33025,N_34792);
nor U36453 (N_36453,N_32955,N_33353);
xor U36454 (N_36454,N_34187,N_32801);
or U36455 (N_36455,N_33870,N_34658);
or U36456 (N_36456,N_33654,N_33453);
or U36457 (N_36457,N_33873,N_32834);
and U36458 (N_36458,N_33829,N_34100);
and U36459 (N_36459,N_34112,N_32709);
nor U36460 (N_36460,N_34625,N_33887);
or U36461 (N_36461,N_34147,N_34157);
nor U36462 (N_36462,N_32722,N_32992);
xnor U36463 (N_36463,N_33412,N_33445);
and U36464 (N_36464,N_34356,N_34040);
or U36465 (N_36465,N_34913,N_33847);
and U36466 (N_36466,N_33447,N_33287);
and U36467 (N_36467,N_32837,N_33813);
xor U36468 (N_36468,N_33679,N_34704);
or U36469 (N_36469,N_34296,N_33447);
nand U36470 (N_36470,N_33036,N_32587);
nor U36471 (N_36471,N_32653,N_34758);
or U36472 (N_36472,N_33252,N_34839);
nand U36473 (N_36473,N_33688,N_32969);
nor U36474 (N_36474,N_33392,N_34872);
or U36475 (N_36475,N_33958,N_32620);
or U36476 (N_36476,N_34831,N_34889);
nor U36477 (N_36477,N_33163,N_33096);
or U36478 (N_36478,N_34896,N_33330);
nand U36479 (N_36479,N_32801,N_32849);
or U36480 (N_36480,N_34157,N_33334);
nor U36481 (N_36481,N_33453,N_32614);
nand U36482 (N_36482,N_33791,N_32706);
and U36483 (N_36483,N_34536,N_33188);
and U36484 (N_36484,N_33769,N_32973);
nor U36485 (N_36485,N_33026,N_33544);
nor U36486 (N_36486,N_34415,N_34075);
and U36487 (N_36487,N_33251,N_33322);
and U36488 (N_36488,N_34513,N_33176);
nand U36489 (N_36489,N_34393,N_34885);
xnor U36490 (N_36490,N_33881,N_32560);
nor U36491 (N_36491,N_33113,N_33370);
nand U36492 (N_36492,N_33849,N_33086);
nand U36493 (N_36493,N_34550,N_34090);
and U36494 (N_36494,N_33143,N_34528);
nor U36495 (N_36495,N_32756,N_32971);
nor U36496 (N_36496,N_34353,N_32739);
nor U36497 (N_36497,N_32952,N_34037);
and U36498 (N_36498,N_33953,N_34260);
nor U36499 (N_36499,N_33459,N_34849);
or U36500 (N_36500,N_32854,N_34853);
or U36501 (N_36501,N_34537,N_34684);
or U36502 (N_36502,N_32708,N_33183);
or U36503 (N_36503,N_34691,N_32504);
nand U36504 (N_36504,N_33629,N_33431);
or U36505 (N_36505,N_32679,N_34594);
or U36506 (N_36506,N_33761,N_32523);
nor U36507 (N_36507,N_32628,N_32992);
nand U36508 (N_36508,N_32987,N_33502);
and U36509 (N_36509,N_33690,N_34303);
nor U36510 (N_36510,N_32595,N_33900);
and U36511 (N_36511,N_34402,N_33692);
and U36512 (N_36512,N_34871,N_34570);
nor U36513 (N_36513,N_33444,N_34988);
nand U36514 (N_36514,N_34530,N_34819);
or U36515 (N_36515,N_33141,N_32923);
nand U36516 (N_36516,N_33759,N_32767);
nor U36517 (N_36517,N_33420,N_33524);
and U36518 (N_36518,N_34967,N_33407);
xor U36519 (N_36519,N_33160,N_34344);
or U36520 (N_36520,N_33114,N_33637);
nor U36521 (N_36521,N_34849,N_34566);
nor U36522 (N_36522,N_34477,N_33185);
nor U36523 (N_36523,N_34258,N_34395);
nor U36524 (N_36524,N_34833,N_34506);
nor U36525 (N_36525,N_33580,N_34054);
or U36526 (N_36526,N_34291,N_34451);
nor U36527 (N_36527,N_32657,N_33431);
and U36528 (N_36528,N_33971,N_34258);
or U36529 (N_36529,N_34028,N_33254);
or U36530 (N_36530,N_33210,N_33441);
nor U36531 (N_36531,N_33280,N_34346);
nor U36532 (N_36532,N_33696,N_34990);
or U36533 (N_36533,N_32776,N_33483);
nor U36534 (N_36534,N_33151,N_34245);
nand U36535 (N_36535,N_32913,N_34238);
nand U36536 (N_36536,N_32635,N_34911);
xor U36537 (N_36537,N_33600,N_34425);
nand U36538 (N_36538,N_33589,N_33816);
xnor U36539 (N_36539,N_33438,N_34407);
nor U36540 (N_36540,N_33564,N_34746);
xnor U36541 (N_36541,N_33755,N_34555);
or U36542 (N_36542,N_34029,N_33826);
nand U36543 (N_36543,N_33721,N_34666);
nor U36544 (N_36544,N_32941,N_34823);
or U36545 (N_36545,N_34096,N_34950);
or U36546 (N_36546,N_33221,N_34561);
nand U36547 (N_36547,N_32808,N_34998);
or U36548 (N_36548,N_34439,N_33689);
xnor U36549 (N_36549,N_32512,N_32978);
nor U36550 (N_36550,N_32680,N_34738);
and U36551 (N_36551,N_34479,N_32887);
nand U36552 (N_36552,N_34853,N_34134);
and U36553 (N_36553,N_34090,N_34909);
nor U36554 (N_36554,N_33372,N_34438);
nand U36555 (N_36555,N_32670,N_34550);
nor U36556 (N_36556,N_33533,N_33130);
and U36557 (N_36557,N_34137,N_33730);
or U36558 (N_36558,N_34021,N_34066);
and U36559 (N_36559,N_33436,N_33314);
or U36560 (N_36560,N_34868,N_34733);
and U36561 (N_36561,N_32644,N_33550);
nand U36562 (N_36562,N_32881,N_33812);
nor U36563 (N_36563,N_33773,N_34757);
nand U36564 (N_36564,N_34697,N_34380);
nor U36565 (N_36565,N_32518,N_32867);
nor U36566 (N_36566,N_34367,N_34110);
nor U36567 (N_36567,N_33703,N_33313);
xnor U36568 (N_36568,N_34961,N_33516);
and U36569 (N_36569,N_34736,N_33794);
or U36570 (N_36570,N_34628,N_33283);
or U36571 (N_36571,N_34937,N_34361);
xor U36572 (N_36572,N_34631,N_34480);
nand U36573 (N_36573,N_33879,N_32594);
or U36574 (N_36574,N_34498,N_33026);
nand U36575 (N_36575,N_34435,N_34081);
nor U36576 (N_36576,N_33671,N_33599);
or U36577 (N_36577,N_33532,N_32825);
nor U36578 (N_36578,N_33488,N_32757);
or U36579 (N_36579,N_34790,N_34602);
or U36580 (N_36580,N_32882,N_32979);
nand U36581 (N_36581,N_33356,N_32636);
and U36582 (N_36582,N_33555,N_32658);
or U36583 (N_36583,N_33008,N_33478);
or U36584 (N_36584,N_33975,N_33426);
or U36585 (N_36585,N_34188,N_34047);
nand U36586 (N_36586,N_34358,N_33354);
or U36587 (N_36587,N_33167,N_33466);
nor U36588 (N_36588,N_34989,N_34049);
nand U36589 (N_36589,N_33447,N_33532);
nand U36590 (N_36590,N_34562,N_34613);
and U36591 (N_36591,N_32805,N_33150);
nand U36592 (N_36592,N_33733,N_33904);
nand U36593 (N_36593,N_32726,N_32609);
nor U36594 (N_36594,N_34127,N_32663);
or U36595 (N_36595,N_34996,N_33261);
nand U36596 (N_36596,N_32757,N_34183);
nand U36597 (N_36597,N_33688,N_34188);
nor U36598 (N_36598,N_34832,N_33911);
and U36599 (N_36599,N_33447,N_33716);
nor U36600 (N_36600,N_32942,N_33811);
and U36601 (N_36601,N_32775,N_34480);
or U36602 (N_36602,N_32565,N_34940);
and U36603 (N_36603,N_33870,N_34207);
and U36604 (N_36604,N_32873,N_33771);
nand U36605 (N_36605,N_34428,N_34656);
nand U36606 (N_36606,N_34610,N_34885);
nand U36607 (N_36607,N_34956,N_33637);
and U36608 (N_36608,N_34250,N_34292);
or U36609 (N_36609,N_32610,N_33457);
nor U36610 (N_36610,N_34270,N_32794);
and U36611 (N_36611,N_33035,N_34367);
nand U36612 (N_36612,N_32588,N_34372);
or U36613 (N_36613,N_34635,N_32930);
nand U36614 (N_36614,N_33688,N_33784);
and U36615 (N_36615,N_33555,N_34933);
and U36616 (N_36616,N_34618,N_32885);
nor U36617 (N_36617,N_34314,N_34550);
xnor U36618 (N_36618,N_33962,N_32532);
nor U36619 (N_36619,N_33105,N_33987);
nor U36620 (N_36620,N_34592,N_32685);
nor U36621 (N_36621,N_33227,N_34198);
or U36622 (N_36622,N_34724,N_34619);
nand U36623 (N_36623,N_33483,N_33438);
nor U36624 (N_36624,N_34303,N_34891);
and U36625 (N_36625,N_34980,N_33016);
nor U36626 (N_36626,N_34386,N_32521);
nand U36627 (N_36627,N_33240,N_32882);
and U36628 (N_36628,N_33377,N_32835);
xor U36629 (N_36629,N_33790,N_34867);
nor U36630 (N_36630,N_33714,N_33549);
and U36631 (N_36631,N_34822,N_32515);
nor U36632 (N_36632,N_33737,N_34858);
nor U36633 (N_36633,N_33674,N_34324);
and U36634 (N_36634,N_33601,N_33250);
or U36635 (N_36635,N_33487,N_34995);
or U36636 (N_36636,N_33804,N_34620);
nand U36637 (N_36637,N_32927,N_32665);
xor U36638 (N_36638,N_34684,N_34954);
nor U36639 (N_36639,N_33994,N_33806);
nand U36640 (N_36640,N_33869,N_34754);
nor U36641 (N_36641,N_34253,N_32862);
or U36642 (N_36642,N_32633,N_32737);
nor U36643 (N_36643,N_33359,N_32784);
nand U36644 (N_36644,N_34011,N_33381);
nor U36645 (N_36645,N_33426,N_32752);
and U36646 (N_36646,N_34772,N_34510);
nor U36647 (N_36647,N_34650,N_34270);
nor U36648 (N_36648,N_32865,N_32859);
or U36649 (N_36649,N_34764,N_32557);
nand U36650 (N_36650,N_32832,N_33690);
or U36651 (N_36651,N_34242,N_34049);
and U36652 (N_36652,N_34883,N_32827);
nand U36653 (N_36653,N_33927,N_32874);
or U36654 (N_36654,N_33942,N_32560);
xor U36655 (N_36655,N_34105,N_34578);
or U36656 (N_36656,N_33909,N_32645);
and U36657 (N_36657,N_34144,N_34408);
and U36658 (N_36658,N_34301,N_33478);
xor U36659 (N_36659,N_33450,N_33473);
nor U36660 (N_36660,N_34475,N_34988);
or U36661 (N_36661,N_33230,N_33337);
and U36662 (N_36662,N_33841,N_33862);
nand U36663 (N_36663,N_33877,N_33740);
nor U36664 (N_36664,N_33906,N_32815);
xor U36665 (N_36665,N_34979,N_34152);
nand U36666 (N_36666,N_32841,N_34757);
nand U36667 (N_36667,N_34123,N_32854);
or U36668 (N_36668,N_34102,N_34148);
and U36669 (N_36669,N_34292,N_34455);
or U36670 (N_36670,N_32517,N_34252);
and U36671 (N_36671,N_34365,N_32796);
nor U36672 (N_36672,N_32731,N_33687);
and U36673 (N_36673,N_33253,N_34029);
nand U36674 (N_36674,N_33793,N_33768);
and U36675 (N_36675,N_34160,N_32980);
or U36676 (N_36676,N_34136,N_33458);
and U36677 (N_36677,N_32962,N_33053);
and U36678 (N_36678,N_34669,N_34074);
and U36679 (N_36679,N_33875,N_34743);
nand U36680 (N_36680,N_34514,N_33666);
and U36681 (N_36681,N_33448,N_34276);
nor U36682 (N_36682,N_32596,N_32877);
nor U36683 (N_36683,N_34107,N_32602);
and U36684 (N_36684,N_34514,N_32603);
and U36685 (N_36685,N_33786,N_32528);
xor U36686 (N_36686,N_34549,N_33247);
and U36687 (N_36687,N_34159,N_32503);
xnor U36688 (N_36688,N_34614,N_32804);
nand U36689 (N_36689,N_34051,N_33413);
and U36690 (N_36690,N_32581,N_34690);
or U36691 (N_36691,N_33354,N_32808);
nor U36692 (N_36692,N_34370,N_34163);
nor U36693 (N_36693,N_33744,N_33493);
nand U36694 (N_36694,N_32652,N_33320);
and U36695 (N_36695,N_34018,N_32870);
nand U36696 (N_36696,N_33618,N_33183);
or U36697 (N_36697,N_33311,N_34617);
and U36698 (N_36698,N_34041,N_34349);
nand U36699 (N_36699,N_34714,N_33437);
or U36700 (N_36700,N_33318,N_34609);
and U36701 (N_36701,N_32522,N_34546);
and U36702 (N_36702,N_33525,N_33606);
nand U36703 (N_36703,N_34536,N_33466);
or U36704 (N_36704,N_33782,N_34306);
xnor U36705 (N_36705,N_32781,N_34628);
nor U36706 (N_36706,N_32541,N_34357);
or U36707 (N_36707,N_34796,N_33127);
or U36708 (N_36708,N_34464,N_33668);
xnor U36709 (N_36709,N_32813,N_33977);
and U36710 (N_36710,N_34108,N_33636);
xor U36711 (N_36711,N_34977,N_32555);
or U36712 (N_36712,N_34743,N_33337);
nor U36713 (N_36713,N_34107,N_34048);
xor U36714 (N_36714,N_33132,N_33138);
nor U36715 (N_36715,N_33837,N_32764);
and U36716 (N_36716,N_33923,N_34885);
or U36717 (N_36717,N_33319,N_32956);
nand U36718 (N_36718,N_34884,N_34200);
or U36719 (N_36719,N_33393,N_32501);
nor U36720 (N_36720,N_33376,N_32725);
nand U36721 (N_36721,N_32884,N_32965);
nor U36722 (N_36722,N_33312,N_34341);
nand U36723 (N_36723,N_32791,N_32634);
and U36724 (N_36724,N_33029,N_33699);
or U36725 (N_36725,N_33188,N_34539);
or U36726 (N_36726,N_33808,N_34805);
nor U36727 (N_36727,N_34955,N_32835);
and U36728 (N_36728,N_32930,N_33184);
nor U36729 (N_36729,N_34853,N_33972);
or U36730 (N_36730,N_33028,N_34728);
and U36731 (N_36731,N_33956,N_34819);
nand U36732 (N_36732,N_34952,N_34054);
xor U36733 (N_36733,N_32961,N_33791);
nand U36734 (N_36734,N_33721,N_34613);
and U36735 (N_36735,N_34246,N_34485);
nand U36736 (N_36736,N_34968,N_32670);
or U36737 (N_36737,N_32666,N_34058);
nand U36738 (N_36738,N_32571,N_34179);
or U36739 (N_36739,N_34165,N_34163);
nor U36740 (N_36740,N_34301,N_34546);
nor U36741 (N_36741,N_32758,N_34555);
nor U36742 (N_36742,N_33350,N_33234);
or U36743 (N_36743,N_33523,N_34017);
and U36744 (N_36744,N_32912,N_32525);
nor U36745 (N_36745,N_33065,N_32578);
nor U36746 (N_36746,N_32813,N_32698);
and U36747 (N_36747,N_32969,N_33565);
and U36748 (N_36748,N_34620,N_32674);
or U36749 (N_36749,N_32800,N_32766);
nor U36750 (N_36750,N_34169,N_33677);
nand U36751 (N_36751,N_34706,N_34105);
nand U36752 (N_36752,N_33638,N_33373);
and U36753 (N_36753,N_34451,N_34917);
nor U36754 (N_36754,N_33679,N_33126);
or U36755 (N_36755,N_34471,N_33975);
nor U36756 (N_36756,N_34622,N_32973);
or U36757 (N_36757,N_34298,N_33914);
or U36758 (N_36758,N_34755,N_34148);
nor U36759 (N_36759,N_34085,N_32610);
nand U36760 (N_36760,N_34361,N_34801);
xor U36761 (N_36761,N_33131,N_33509);
and U36762 (N_36762,N_34422,N_34854);
nand U36763 (N_36763,N_33512,N_33832);
and U36764 (N_36764,N_33961,N_33036);
nor U36765 (N_36765,N_32698,N_34161);
nor U36766 (N_36766,N_34135,N_32838);
nor U36767 (N_36767,N_33678,N_33617);
nand U36768 (N_36768,N_33398,N_32574);
nand U36769 (N_36769,N_34719,N_33627);
and U36770 (N_36770,N_34027,N_34422);
xor U36771 (N_36771,N_33214,N_34068);
and U36772 (N_36772,N_33254,N_32507);
nor U36773 (N_36773,N_34330,N_32923);
nand U36774 (N_36774,N_32638,N_32689);
nor U36775 (N_36775,N_33752,N_33288);
or U36776 (N_36776,N_34345,N_34604);
nand U36777 (N_36777,N_33710,N_33800);
nand U36778 (N_36778,N_32505,N_33246);
and U36779 (N_36779,N_33080,N_34364);
nand U36780 (N_36780,N_33077,N_34097);
and U36781 (N_36781,N_32804,N_32992);
nor U36782 (N_36782,N_34701,N_33003);
xor U36783 (N_36783,N_33254,N_34532);
nor U36784 (N_36784,N_34972,N_34577);
nand U36785 (N_36785,N_33476,N_33596);
or U36786 (N_36786,N_34338,N_32874);
nand U36787 (N_36787,N_34860,N_32669);
nor U36788 (N_36788,N_33916,N_33002);
or U36789 (N_36789,N_33337,N_32701);
and U36790 (N_36790,N_33688,N_32609);
or U36791 (N_36791,N_34872,N_34813);
nand U36792 (N_36792,N_34067,N_32860);
nand U36793 (N_36793,N_34296,N_32968);
or U36794 (N_36794,N_32641,N_34404);
nor U36795 (N_36795,N_33484,N_33757);
nand U36796 (N_36796,N_34690,N_33190);
nor U36797 (N_36797,N_33579,N_32641);
nor U36798 (N_36798,N_34326,N_33622);
xnor U36799 (N_36799,N_34372,N_33793);
or U36800 (N_36800,N_34560,N_33681);
and U36801 (N_36801,N_34500,N_33655);
nand U36802 (N_36802,N_34070,N_34456);
nor U36803 (N_36803,N_33034,N_33841);
or U36804 (N_36804,N_33144,N_33419);
and U36805 (N_36805,N_33619,N_33803);
and U36806 (N_36806,N_33706,N_33141);
xnor U36807 (N_36807,N_33638,N_34858);
or U36808 (N_36808,N_33362,N_33332);
nand U36809 (N_36809,N_34690,N_33400);
xor U36810 (N_36810,N_34074,N_32840);
nand U36811 (N_36811,N_33651,N_34119);
and U36812 (N_36812,N_33256,N_34924);
or U36813 (N_36813,N_33407,N_33903);
nand U36814 (N_36814,N_34129,N_34220);
nand U36815 (N_36815,N_32868,N_33425);
nand U36816 (N_36816,N_34778,N_33295);
and U36817 (N_36817,N_33342,N_33598);
and U36818 (N_36818,N_33706,N_33196);
nand U36819 (N_36819,N_32921,N_34790);
or U36820 (N_36820,N_33227,N_34702);
nor U36821 (N_36821,N_33945,N_33465);
nor U36822 (N_36822,N_33346,N_33348);
nand U36823 (N_36823,N_32852,N_34901);
nor U36824 (N_36824,N_33558,N_34438);
xnor U36825 (N_36825,N_33284,N_33964);
nand U36826 (N_36826,N_34008,N_34198);
or U36827 (N_36827,N_32919,N_33681);
and U36828 (N_36828,N_33496,N_32507);
nand U36829 (N_36829,N_33911,N_33598);
or U36830 (N_36830,N_34605,N_34255);
and U36831 (N_36831,N_33771,N_32573);
nor U36832 (N_36832,N_34555,N_34438);
or U36833 (N_36833,N_32666,N_32993);
or U36834 (N_36834,N_34727,N_33807);
nor U36835 (N_36835,N_33666,N_33633);
nand U36836 (N_36836,N_33704,N_32762);
nand U36837 (N_36837,N_34940,N_33122);
and U36838 (N_36838,N_32699,N_34884);
and U36839 (N_36839,N_34915,N_33417);
xnor U36840 (N_36840,N_34359,N_34228);
nor U36841 (N_36841,N_34608,N_33282);
nand U36842 (N_36842,N_33781,N_32682);
xnor U36843 (N_36843,N_34368,N_34620);
nand U36844 (N_36844,N_34209,N_33818);
xnor U36845 (N_36845,N_32700,N_33158);
nand U36846 (N_36846,N_32583,N_34764);
or U36847 (N_36847,N_33680,N_34517);
or U36848 (N_36848,N_34732,N_34928);
and U36849 (N_36849,N_34986,N_33443);
nand U36850 (N_36850,N_34180,N_34267);
xnor U36851 (N_36851,N_33823,N_33352);
nor U36852 (N_36852,N_33030,N_32628);
or U36853 (N_36853,N_33135,N_34973);
nor U36854 (N_36854,N_34043,N_34550);
nand U36855 (N_36855,N_33647,N_33293);
xor U36856 (N_36856,N_34287,N_34522);
nand U36857 (N_36857,N_32764,N_34358);
nand U36858 (N_36858,N_32939,N_34064);
or U36859 (N_36859,N_33129,N_33244);
nor U36860 (N_36860,N_33240,N_32864);
nand U36861 (N_36861,N_34154,N_34148);
or U36862 (N_36862,N_34151,N_32562);
and U36863 (N_36863,N_33236,N_33186);
or U36864 (N_36864,N_32618,N_33371);
nor U36865 (N_36865,N_34926,N_32604);
nor U36866 (N_36866,N_33123,N_34609);
or U36867 (N_36867,N_32887,N_34713);
and U36868 (N_36868,N_34000,N_33065);
and U36869 (N_36869,N_33619,N_34588);
or U36870 (N_36870,N_34234,N_34459);
nand U36871 (N_36871,N_33638,N_34861);
nand U36872 (N_36872,N_33692,N_32951);
or U36873 (N_36873,N_34500,N_33056);
or U36874 (N_36874,N_34252,N_33384);
and U36875 (N_36875,N_33971,N_32906);
nor U36876 (N_36876,N_34696,N_34429);
and U36877 (N_36877,N_34858,N_33867);
and U36878 (N_36878,N_33138,N_33532);
and U36879 (N_36879,N_32994,N_34895);
or U36880 (N_36880,N_33828,N_32874);
xnor U36881 (N_36881,N_34745,N_34145);
or U36882 (N_36882,N_33711,N_34799);
or U36883 (N_36883,N_32978,N_34069);
nor U36884 (N_36884,N_33767,N_34774);
nand U36885 (N_36885,N_32788,N_34287);
nand U36886 (N_36886,N_33828,N_33567);
nor U36887 (N_36887,N_34870,N_33248);
or U36888 (N_36888,N_32509,N_33942);
nand U36889 (N_36889,N_34356,N_33036);
or U36890 (N_36890,N_34126,N_34046);
xor U36891 (N_36891,N_34093,N_33377);
and U36892 (N_36892,N_33130,N_34417);
nor U36893 (N_36893,N_33708,N_34184);
nor U36894 (N_36894,N_34849,N_34663);
nand U36895 (N_36895,N_33816,N_34455);
nand U36896 (N_36896,N_34119,N_32824);
nor U36897 (N_36897,N_33182,N_34209);
xnor U36898 (N_36898,N_33038,N_34620);
and U36899 (N_36899,N_33526,N_32672);
nor U36900 (N_36900,N_34857,N_33134);
or U36901 (N_36901,N_33034,N_32868);
and U36902 (N_36902,N_34521,N_32990);
xor U36903 (N_36903,N_33824,N_33635);
nor U36904 (N_36904,N_34473,N_33299);
nand U36905 (N_36905,N_34945,N_34413);
and U36906 (N_36906,N_33094,N_34060);
or U36907 (N_36907,N_33450,N_33634);
and U36908 (N_36908,N_32501,N_33818);
nor U36909 (N_36909,N_34542,N_34237);
nand U36910 (N_36910,N_33696,N_33850);
nor U36911 (N_36911,N_33834,N_34402);
xnor U36912 (N_36912,N_33823,N_33591);
nand U36913 (N_36913,N_34887,N_33123);
nor U36914 (N_36914,N_32779,N_34442);
and U36915 (N_36915,N_34025,N_33049);
nand U36916 (N_36916,N_32901,N_34098);
and U36917 (N_36917,N_34991,N_32537);
and U36918 (N_36918,N_34891,N_34892);
and U36919 (N_36919,N_34653,N_32951);
and U36920 (N_36920,N_33039,N_34647);
nand U36921 (N_36921,N_32606,N_33501);
nand U36922 (N_36922,N_32572,N_32905);
and U36923 (N_36923,N_34975,N_32922);
or U36924 (N_36924,N_32986,N_34032);
and U36925 (N_36925,N_33649,N_32928);
xor U36926 (N_36926,N_33943,N_33620);
nor U36927 (N_36927,N_32680,N_32596);
and U36928 (N_36928,N_33591,N_34935);
xnor U36929 (N_36929,N_33858,N_34714);
or U36930 (N_36930,N_32786,N_34610);
nor U36931 (N_36931,N_34384,N_32978);
nor U36932 (N_36932,N_34048,N_33673);
nand U36933 (N_36933,N_33770,N_33489);
and U36934 (N_36934,N_32996,N_34690);
xor U36935 (N_36935,N_34838,N_32511);
or U36936 (N_36936,N_33402,N_34148);
and U36937 (N_36937,N_33227,N_34061);
nor U36938 (N_36938,N_34954,N_33025);
nor U36939 (N_36939,N_33901,N_32743);
or U36940 (N_36940,N_33123,N_34188);
and U36941 (N_36941,N_33169,N_32998);
nand U36942 (N_36942,N_32693,N_34850);
nor U36943 (N_36943,N_33918,N_33175);
and U36944 (N_36944,N_34139,N_34151);
and U36945 (N_36945,N_34097,N_33185);
nand U36946 (N_36946,N_32533,N_33981);
nand U36947 (N_36947,N_34929,N_33948);
nor U36948 (N_36948,N_33222,N_32711);
nand U36949 (N_36949,N_32698,N_32856);
or U36950 (N_36950,N_32781,N_34383);
nor U36951 (N_36951,N_34051,N_33254);
nor U36952 (N_36952,N_33333,N_34083);
nor U36953 (N_36953,N_34385,N_33306);
nor U36954 (N_36954,N_34936,N_33733);
nor U36955 (N_36955,N_34427,N_33394);
or U36956 (N_36956,N_34550,N_34615);
or U36957 (N_36957,N_33016,N_33154);
nor U36958 (N_36958,N_34917,N_34340);
nor U36959 (N_36959,N_32784,N_32872);
or U36960 (N_36960,N_33281,N_34031);
xor U36961 (N_36961,N_32697,N_34064);
and U36962 (N_36962,N_34358,N_33395);
nor U36963 (N_36963,N_34934,N_33638);
nand U36964 (N_36964,N_33809,N_34977);
xnor U36965 (N_36965,N_33855,N_34537);
and U36966 (N_36966,N_32584,N_32556);
nor U36967 (N_36967,N_33631,N_34283);
nand U36968 (N_36968,N_34744,N_32507);
and U36969 (N_36969,N_32523,N_34753);
nor U36970 (N_36970,N_33079,N_34280);
xor U36971 (N_36971,N_33941,N_32847);
and U36972 (N_36972,N_33198,N_33796);
and U36973 (N_36973,N_33841,N_33967);
or U36974 (N_36974,N_32879,N_33093);
or U36975 (N_36975,N_32801,N_33963);
nand U36976 (N_36976,N_32571,N_33915);
nor U36977 (N_36977,N_33234,N_32683);
and U36978 (N_36978,N_34673,N_34300);
and U36979 (N_36979,N_33574,N_32690);
and U36980 (N_36980,N_32949,N_34576);
nand U36981 (N_36981,N_33696,N_33076);
nor U36982 (N_36982,N_33177,N_34824);
nand U36983 (N_36983,N_34664,N_33948);
nor U36984 (N_36984,N_34376,N_32965);
and U36985 (N_36985,N_34497,N_33909);
nand U36986 (N_36986,N_32845,N_32698);
or U36987 (N_36987,N_33809,N_34812);
nand U36988 (N_36988,N_34784,N_33636);
xnor U36989 (N_36989,N_32712,N_32835);
nand U36990 (N_36990,N_33914,N_33329);
nand U36991 (N_36991,N_34148,N_33565);
nor U36992 (N_36992,N_32572,N_32829);
nor U36993 (N_36993,N_34598,N_33433);
xor U36994 (N_36994,N_32686,N_32523);
nand U36995 (N_36995,N_34461,N_32795);
and U36996 (N_36996,N_33609,N_34939);
nand U36997 (N_36997,N_34773,N_32839);
nor U36998 (N_36998,N_33843,N_34380);
and U36999 (N_36999,N_34101,N_33237);
nand U37000 (N_37000,N_32584,N_33930);
and U37001 (N_37001,N_33063,N_33959);
and U37002 (N_37002,N_33725,N_34249);
nor U37003 (N_37003,N_33942,N_33587);
or U37004 (N_37004,N_32984,N_34978);
and U37005 (N_37005,N_34246,N_34783);
or U37006 (N_37006,N_34787,N_32976);
nor U37007 (N_37007,N_33149,N_32562);
nand U37008 (N_37008,N_32616,N_32826);
and U37009 (N_37009,N_32925,N_33879);
and U37010 (N_37010,N_34534,N_34895);
and U37011 (N_37011,N_32836,N_33848);
or U37012 (N_37012,N_34568,N_34401);
or U37013 (N_37013,N_32571,N_33098);
or U37014 (N_37014,N_33841,N_34860);
or U37015 (N_37015,N_33513,N_34494);
and U37016 (N_37016,N_34594,N_33205);
nor U37017 (N_37017,N_34868,N_34612);
nor U37018 (N_37018,N_34902,N_34117);
nor U37019 (N_37019,N_33214,N_34184);
or U37020 (N_37020,N_34849,N_34003);
and U37021 (N_37021,N_32508,N_32641);
or U37022 (N_37022,N_34817,N_33838);
xor U37023 (N_37023,N_32656,N_33862);
or U37024 (N_37024,N_34551,N_33760);
nor U37025 (N_37025,N_33516,N_33197);
and U37026 (N_37026,N_34551,N_33334);
or U37027 (N_37027,N_32768,N_33655);
or U37028 (N_37028,N_32610,N_32948);
or U37029 (N_37029,N_34334,N_33027);
or U37030 (N_37030,N_33166,N_33616);
or U37031 (N_37031,N_34543,N_33162);
and U37032 (N_37032,N_33505,N_34104);
or U37033 (N_37033,N_33922,N_33556);
and U37034 (N_37034,N_34462,N_34082);
nand U37035 (N_37035,N_33950,N_33845);
or U37036 (N_37036,N_33071,N_34438);
or U37037 (N_37037,N_34506,N_33344);
nand U37038 (N_37038,N_33980,N_32773);
and U37039 (N_37039,N_33862,N_32679);
and U37040 (N_37040,N_34193,N_33940);
nor U37041 (N_37041,N_32884,N_33412);
and U37042 (N_37042,N_32987,N_32663);
and U37043 (N_37043,N_33184,N_32953);
or U37044 (N_37044,N_32825,N_33040);
and U37045 (N_37045,N_34490,N_32507);
nor U37046 (N_37046,N_32625,N_34842);
and U37047 (N_37047,N_33935,N_34011);
nand U37048 (N_37048,N_34748,N_33234);
and U37049 (N_37049,N_33982,N_34371);
nor U37050 (N_37050,N_33835,N_32620);
nor U37051 (N_37051,N_34651,N_32644);
nand U37052 (N_37052,N_34738,N_33817);
xnor U37053 (N_37053,N_34820,N_33118);
and U37054 (N_37054,N_32959,N_34478);
nand U37055 (N_37055,N_34774,N_33795);
nor U37056 (N_37056,N_33283,N_34574);
and U37057 (N_37057,N_34583,N_33176);
nor U37058 (N_37058,N_34953,N_33935);
nor U37059 (N_37059,N_33751,N_32795);
nand U37060 (N_37060,N_32532,N_33166);
nor U37061 (N_37061,N_33310,N_33041);
nor U37062 (N_37062,N_33329,N_33108);
or U37063 (N_37063,N_34472,N_33938);
and U37064 (N_37064,N_32698,N_33662);
or U37065 (N_37065,N_33985,N_32979);
and U37066 (N_37066,N_33215,N_33418);
xnor U37067 (N_37067,N_32537,N_34081);
nand U37068 (N_37068,N_34341,N_33321);
nand U37069 (N_37069,N_34762,N_33638);
and U37070 (N_37070,N_32876,N_33437);
or U37071 (N_37071,N_33151,N_33136);
and U37072 (N_37072,N_32891,N_33554);
and U37073 (N_37073,N_33910,N_34347);
xor U37074 (N_37074,N_32672,N_33018);
or U37075 (N_37075,N_34862,N_34157);
xor U37076 (N_37076,N_33414,N_34143);
or U37077 (N_37077,N_34873,N_33723);
and U37078 (N_37078,N_34422,N_32665);
and U37079 (N_37079,N_33338,N_33933);
nor U37080 (N_37080,N_33291,N_33592);
or U37081 (N_37081,N_34037,N_34226);
nor U37082 (N_37082,N_34058,N_33215);
and U37083 (N_37083,N_33063,N_34909);
and U37084 (N_37084,N_33643,N_32504);
nor U37085 (N_37085,N_34623,N_32656);
or U37086 (N_37086,N_34327,N_34105);
and U37087 (N_37087,N_34737,N_33112);
and U37088 (N_37088,N_34390,N_33186);
or U37089 (N_37089,N_33390,N_34393);
nor U37090 (N_37090,N_34327,N_34489);
or U37091 (N_37091,N_32593,N_34531);
nor U37092 (N_37092,N_34731,N_34524);
nand U37093 (N_37093,N_32587,N_34705);
and U37094 (N_37094,N_34319,N_34781);
xnor U37095 (N_37095,N_32509,N_32804);
and U37096 (N_37096,N_34490,N_32633);
nand U37097 (N_37097,N_34798,N_34972);
nor U37098 (N_37098,N_33512,N_34455);
nor U37099 (N_37099,N_32622,N_34831);
or U37100 (N_37100,N_33054,N_33268);
or U37101 (N_37101,N_34589,N_33281);
nor U37102 (N_37102,N_32745,N_33206);
and U37103 (N_37103,N_33024,N_32973);
or U37104 (N_37104,N_33763,N_34256);
nor U37105 (N_37105,N_34626,N_32680);
or U37106 (N_37106,N_34546,N_34135);
nor U37107 (N_37107,N_32750,N_33074);
nor U37108 (N_37108,N_33085,N_32907);
or U37109 (N_37109,N_33771,N_34074);
or U37110 (N_37110,N_34474,N_34071);
nand U37111 (N_37111,N_34601,N_33458);
xnor U37112 (N_37112,N_33816,N_33392);
xnor U37113 (N_37113,N_33977,N_33571);
or U37114 (N_37114,N_34894,N_34096);
nand U37115 (N_37115,N_33164,N_33630);
nand U37116 (N_37116,N_33640,N_34709);
and U37117 (N_37117,N_34681,N_33471);
and U37118 (N_37118,N_34993,N_33811);
and U37119 (N_37119,N_34506,N_33619);
nand U37120 (N_37120,N_33613,N_34324);
or U37121 (N_37121,N_34032,N_33646);
and U37122 (N_37122,N_33881,N_34668);
nand U37123 (N_37123,N_33881,N_34794);
and U37124 (N_37124,N_34528,N_33142);
nand U37125 (N_37125,N_34644,N_34461);
and U37126 (N_37126,N_33337,N_33172);
nor U37127 (N_37127,N_34074,N_34950);
or U37128 (N_37128,N_34018,N_34363);
xor U37129 (N_37129,N_34638,N_34749);
nor U37130 (N_37130,N_32792,N_33151);
nor U37131 (N_37131,N_32986,N_33512);
nor U37132 (N_37132,N_33405,N_32675);
and U37133 (N_37133,N_34604,N_33510);
nand U37134 (N_37134,N_33052,N_32707);
or U37135 (N_37135,N_33479,N_34272);
nand U37136 (N_37136,N_32825,N_34960);
and U37137 (N_37137,N_34265,N_34610);
nor U37138 (N_37138,N_33108,N_33575);
or U37139 (N_37139,N_33049,N_32857);
and U37140 (N_37140,N_32559,N_33869);
and U37141 (N_37141,N_33820,N_32966);
or U37142 (N_37142,N_32779,N_34521);
nand U37143 (N_37143,N_33221,N_33039);
or U37144 (N_37144,N_34399,N_34183);
nand U37145 (N_37145,N_34857,N_33979);
xor U37146 (N_37146,N_33732,N_33247);
nand U37147 (N_37147,N_34036,N_34557);
and U37148 (N_37148,N_33443,N_34678);
and U37149 (N_37149,N_34295,N_33597);
or U37150 (N_37150,N_34829,N_33753);
or U37151 (N_37151,N_32571,N_32643);
or U37152 (N_37152,N_32725,N_34409);
or U37153 (N_37153,N_34410,N_33437);
nor U37154 (N_37154,N_32949,N_34413);
nand U37155 (N_37155,N_33975,N_32588);
and U37156 (N_37156,N_34547,N_33400);
nand U37157 (N_37157,N_33933,N_32595);
and U37158 (N_37158,N_33201,N_33405);
or U37159 (N_37159,N_34397,N_33966);
xnor U37160 (N_37160,N_34790,N_34355);
nor U37161 (N_37161,N_32824,N_33299);
nand U37162 (N_37162,N_33088,N_33187);
nand U37163 (N_37163,N_34315,N_33160);
and U37164 (N_37164,N_33805,N_33878);
or U37165 (N_37165,N_34718,N_33986);
and U37166 (N_37166,N_34002,N_34176);
or U37167 (N_37167,N_33089,N_32546);
nand U37168 (N_37168,N_32537,N_32605);
nand U37169 (N_37169,N_33608,N_32627);
xor U37170 (N_37170,N_33075,N_33932);
or U37171 (N_37171,N_33552,N_33853);
or U37172 (N_37172,N_34273,N_32656);
or U37173 (N_37173,N_32660,N_32620);
or U37174 (N_37174,N_33545,N_33488);
and U37175 (N_37175,N_34872,N_34046);
nand U37176 (N_37176,N_32599,N_34305);
and U37177 (N_37177,N_34220,N_32520);
or U37178 (N_37178,N_33233,N_32876);
and U37179 (N_37179,N_34196,N_34885);
and U37180 (N_37180,N_32697,N_34969);
nor U37181 (N_37181,N_34862,N_34819);
and U37182 (N_37182,N_33591,N_33256);
or U37183 (N_37183,N_32998,N_32629);
nor U37184 (N_37184,N_33750,N_34777);
nand U37185 (N_37185,N_34526,N_33634);
and U37186 (N_37186,N_34848,N_34334);
nor U37187 (N_37187,N_33526,N_33995);
or U37188 (N_37188,N_34969,N_33224);
nor U37189 (N_37189,N_34263,N_32881);
nor U37190 (N_37190,N_32839,N_34421);
nand U37191 (N_37191,N_33029,N_34541);
xnor U37192 (N_37192,N_32960,N_33374);
and U37193 (N_37193,N_34513,N_33522);
or U37194 (N_37194,N_34031,N_33188);
nand U37195 (N_37195,N_33800,N_34048);
and U37196 (N_37196,N_32556,N_32546);
or U37197 (N_37197,N_34861,N_34399);
or U37198 (N_37198,N_34914,N_32934);
and U37199 (N_37199,N_33264,N_34641);
nor U37200 (N_37200,N_33618,N_32618);
or U37201 (N_37201,N_32580,N_33844);
or U37202 (N_37202,N_34956,N_33301);
and U37203 (N_37203,N_32549,N_32510);
or U37204 (N_37204,N_33621,N_34054);
or U37205 (N_37205,N_34168,N_33567);
nor U37206 (N_37206,N_33116,N_32538);
or U37207 (N_37207,N_32882,N_32612);
or U37208 (N_37208,N_33503,N_32891);
xor U37209 (N_37209,N_34249,N_33758);
nor U37210 (N_37210,N_34838,N_32795);
nor U37211 (N_37211,N_34878,N_34787);
xnor U37212 (N_37212,N_34897,N_34807);
and U37213 (N_37213,N_33026,N_34672);
nor U37214 (N_37214,N_34993,N_33539);
nor U37215 (N_37215,N_33711,N_33789);
or U37216 (N_37216,N_32751,N_33462);
nor U37217 (N_37217,N_32505,N_33039);
nand U37218 (N_37218,N_32910,N_33973);
or U37219 (N_37219,N_33519,N_33479);
or U37220 (N_37220,N_34242,N_33211);
and U37221 (N_37221,N_32538,N_34494);
or U37222 (N_37222,N_33191,N_32712);
nor U37223 (N_37223,N_33001,N_32952);
and U37224 (N_37224,N_33256,N_34607);
nor U37225 (N_37225,N_34506,N_34976);
nor U37226 (N_37226,N_33629,N_32982);
or U37227 (N_37227,N_33208,N_33780);
nand U37228 (N_37228,N_33310,N_34508);
and U37229 (N_37229,N_34922,N_33751);
and U37230 (N_37230,N_34666,N_33541);
and U37231 (N_37231,N_34869,N_34912);
nand U37232 (N_37232,N_34060,N_34456);
nand U37233 (N_37233,N_33114,N_34914);
xnor U37234 (N_37234,N_33132,N_33083);
nand U37235 (N_37235,N_34442,N_33919);
and U37236 (N_37236,N_34899,N_34530);
xnor U37237 (N_37237,N_34403,N_33160);
and U37238 (N_37238,N_32886,N_33703);
and U37239 (N_37239,N_33111,N_33101);
and U37240 (N_37240,N_33451,N_33078);
xor U37241 (N_37241,N_34481,N_34893);
nor U37242 (N_37242,N_33568,N_33081);
and U37243 (N_37243,N_34324,N_32878);
and U37244 (N_37244,N_34500,N_34632);
nand U37245 (N_37245,N_34828,N_33360);
xnor U37246 (N_37246,N_33973,N_33215);
nand U37247 (N_37247,N_33433,N_32733);
nor U37248 (N_37248,N_34784,N_34054);
nor U37249 (N_37249,N_33399,N_32608);
nand U37250 (N_37250,N_33207,N_33942);
and U37251 (N_37251,N_33310,N_33668);
or U37252 (N_37252,N_33409,N_34527);
or U37253 (N_37253,N_33569,N_34065);
nand U37254 (N_37254,N_33501,N_32644);
xor U37255 (N_37255,N_33228,N_33955);
and U37256 (N_37256,N_32865,N_33308);
nor U37257 (N_37257,N_34704,N_33735);
nand U37258 (N_37258,N_32659,N_32901);
or U37259 (N_37259,N_34643,N_32649);
and U37260 (N_37260,N_34632,N_32634);
xor U37261 (N_37261,N_34177,N_33627);
or U37262 (N_37262,N_34609,N_33732);
nand U37263 (N_37263,N_32804,N_33607);
nor U37264 (N_37264,N_33646,N_33802);
nor U37265 (N_37265,N_32575,N_33528);
and U37266 (N_37266,N_32885,N_32888);
or U37267 (N_37267,N_34852,N_32912);
nand U37268 (N_37268,N_34799,N_32710);
or U37269 (N_37269,N_33693,N_33504);
nor U37270 (N_37270,N_33165,N_34705);
or U37271 (N_37271,N_34752,N_34842);
xnor U37272 (N_37272,N_32650,N_32928);
or U37273 (N_37273,N_34335,N_34043);
or U37274 (N_37274,N_33657,N_32896);
and U37275 (N_37275,N_33280,N_33938);
and U37276 (N_37276,N_33540,N_34262);
or U37277 (N_37277,N_34089,N_33447);
or U37278 (N_37278,N_33213,N_33205);
and U37279 (N_37279,N_33063,N_34827);
or U37280 (N_37280,N_33337,N_34944);
nand U37281 (N_37281,N_33390,N_34968);
xnor U37282 (N_37282,N_33492,N_33470);
or U37283 (N_37283,N_33402,N_33739);
xor U37284 (N_37284,N_33343,N_33040);
nor U37285 (N_37285,N_33336,N_32541);
and U37286 (N_37286,N_34169,N_34097);
nand U37287 (N_37287,N_32519,N_33208);
and U37288 (N_37288,N_34867,N_33447);
or U37289 (N_37289,N_33258,N_33091);
xor U37290 (N_37290,N_32987,N_34899);
nor U37291 (N_37291,N_32597,N_32827);
nor U37292 (N_37292,N_34456,N_34946);
nor U37293 (N_37293,N_32608,N_32897);
nor U37294 (N_37294,N_33698,N_34169);
and U37295 (N_37295,N_32678,N_33434);
nor U37296 (N_37296,N_33924,N_34215);
nor U37297 (N_37297,N_33180,N_33642);
xor U37298 (N_37298,N_33561,N_33993);
and U37299 (N_37299,N_33287,N_34822);
nand U37300 (N_37300,N_34798,N_32958);
or U37301 (N_37301,N_34211,N_34279);
nand U37302 (N_37302,N_32795,N_32532);
and U37303 (N_37303,N_34437,N_32868);
nor U37304 (N_37304,N_33863,N_33667);
and U37305 (N_37305,N_33729,N_34756);
nand U37306 (N_37306,N_32636,N_33891);
nor U37307 (N_37307,N_33430,N_34925);
and U37308 (N_37308,N_34859,N_34846);
nor U37309 (N_37309,N_34629,N_34494);
or U37310 (N_37310,N_34591,N_32603);
nor U37311 (N_37311,N_33086,N_32902);
and U37312 (N_37312,N_32624,N_34920);
and U37313 (N_37313,N_32588,N_32560);
nor U37314 (N_37314,N_33469,N_34217);
nor U37315 (N_37315,N_33706,N_32548);
and U37316 (N_37316,N_34415,N_33277);
xor U37317 (N_37317,N_32873,N_34008);
nor U37318 (N_37318,N_33021,N_33986);
nand U37319 (N_37319,N_34021,N_33125);
and U37320 (N_37320,N_34155,N_33272);
or U37321 (N_37321,N_33271,N_33419);
and U37322 (N_37322,N_32631,N_34326);
or U37323 (N_37323,N_32591,N_34852);
nor U37324 (N_37324,N_33349,N_34081);
nand U37325 (N_37325,N_32568,N_33163);
and U37326 (N_37326,N_32919,N_32981);
nor U37327 (N_37327,N_33862,N_34884);
and U37328 (N_37328,N_32711,N_34789);
or U37329 (N_37329,N_32904,N_33466);
nor U37330 (N_37330,N_34363,N_34509);
nand U37331 (N_37331,N_33959,N_33284);
xor U37332 (N_37332,N_34972,N_32973);
and U37333 (N_37333,N_33353,N_32617);
xor U37334 (N_37334,N_34618,N_33778);
and U37335 (N_37335,N_32858,N_34666);
xnor U37336 (N_37336,N_34971,N_33984);
nor U37337 (N_37337,N_34094,N_33177);
and U37338 (N_37338,N_33246,N_34217);
or U37339 (N_37339,N_34296,N_33389);
nand U37340 (N_37340,N_34689,N_34099);
and U37341 (N_37341,N_33945,N_33457);
and U37342 (N_37342,N_33526,N_34220);
or U37343 (N_37343,N_32733,N_33721);
or U37344 (N_37344,N_32920,N_32647);
nand U37345 (N_37345,N_33626,N_34725);
nor U37346 (N_37346,N_32919,N_34803);
nand U37347 (N_37347,N_34010,N_32777);
or U37348 (N_37348,N_33954,N_34666);
or U37349 (N_37349,N_34280,N_33477);
and U37350 (N_37350,N_33710,N_32583);
xor U37351 (N_37351,N_34080,N_33048);
and U37352 (N_37352,N_33552,N_32835);
or U37353 (N_37353,N_34593,N_33079);
or U37354 (N_37354,N_33017,N_33746);
nand U37355 (N_37355,N_33461,N_33250);
or U37356 (N_37356,N_33239,N_33306);
or U37357 (N_37357,N_33112,N_33714);
or U37358 (N_37358,N_34160,N_33105);
xnor U37359 (N_37359,N_33261,N_33836);
or U37360 (N_37360,N_34392,N_34876);
nor U37361 (N_37361,N_33129,N_33364);
or U37362 (N_37362,N_34563,N_32695);
nor U37363 (N_37363,N_34575,N_34439);
nand U37364 (N_37364,N_33745,N_34645);
and U37365 (N_37365,N_32877,N_34623);
and U37366 (N_37366,N_34128,N_34291);
nor U37367 (N_37367,N_33515,N_32860);
nand U37368 (N_37368,N_34124,N_32716);
nand U37369 (N_37369,N_32626,N_33351);
or U37370 (N_37370,N_34142,N_33893);
nand U37371 (N_37371,N_33412,N_33446);
nand U37372 (N_37372,N_34968,N_32532);
nor U37373 (N_37373,N_33612,N_34971);
or U37374 (N_37374,N_33726,N_33773);
or U37375 (N_37375,N_34691,N_33118);
or U37376 (N_37376,N_34403,N_32917);
and U37377 (N_37377,N_32569,N_34495);
nor U37378 (N_37378,N_33505,N_32575);
nand U37379 (N_37379,N_32902,N_34607);
nand U37380 (N_37380,N_33189,N_33650);
or U37381 (N_37381,N_33882,N_34080);
and U37382 (N_37382,N_33261,N_32775);
or U37383 (N_37383,N_32905,N_34652);
or U37384 (N_37384,N_33745,N_32954);
or U37385 (N_37385,N_33581,N_33875);
nand U37386 (N_37386,N_33946,N_34048);
or U37387 (N_37387,N_33689,N_34170);
or U37388 (N_37388,N_34796,N_34369);
and U37389 (N_37389,N_33068,N_32889);
or U37390 (N_37390,N_33775,N_33661);
nor U37391 (N_37391,N_32612,N_33539);
nor U37392 (N_37392,N_34932,N_33430);
and U37393 (N_37393,N_32516,N_32649);
nand U37394 (N_37394,N_33851,N_32977);
and U37395 (N_37395,N_34180,N_33244);
nor U37396 (N_37396,N_34931,N_34113);
or U37397 (N_37397,N_34367,N_33164);
nor U37398 (N_37398,N_32948,N_34914);
or U37399 (N_37399,N_32698,N_33688);
nor U37400 (N_37400,N_33754,N_33706);
or U37401 (N_37401,N_33925,N_33724);
or U37402 (N_37402,N_34638,N_34270);
or U37403 (N_37403,N_33247,N_34483);
nor U37404 (N_37404,N_34887,N_33530);
and U37405 (N_37405,N_32809,N_34450);
or U37406 (N_37406,N_33184,N_34141);
or U37407 (N_37407,N_34038,N_33653);
xnor U37408 (N_37408,N_32583,N_34859);
nor U37409 (N_37409,N_34892,N_33965);
or U37410 (N_37410,N_33311,N_32696);
nand U37411 (N_37411,N_33781,N_33370);
and U37412 (N_37412,N_33012,N_32958);
nor U37413 (N_37413,N_33530,N_34723);
nor U37414 (N_37414,N_33610,N_33215);
nor U37415 (N_37415,N_33748,N_32766);
or U37416 (N_37416,N_34007,N_33079);
xor U37417 (N_37417,N_34675,N_33855);
nand U37418 (N_37418,N_33669,N_34112);
or U37419 (N_37419,N_32526,N_32644);
xor U37420 (N_37420,N_33018,N_32548);
nand U37421 (N_37421,N_33592,N_34522);
or U37422 (N_37422,N_33917,N_33968);
and U37423 (N_37423,N_33103,N_32500);
or U37424 (N_37424,N_34336,N_33381);
xor U37425 (N_37425,N_34911,N_32982);
or U37426 (N_37426,N_32916,N_33461);
nor U37427 (N_37427,N_32978,N_33631);
nand U37428 (N_37428,N_34653,N_32758);
xor U37429 (N_37429,N_33822,N_34373);
and U37430 (N_37430,N_34564,N_33965);
nor U37431 (N_37431,N_33036,N_34752);
and U37432 (N_37432,N_34814,N_33865);
nor U37433 (N_37433,N_33742,N_33056);
nand U37434 (N_37434,N_34585,N_32525);
xor U37435 (N_37435,N_33213,N_33176);
or U37436 (N_37436,N_33696,N_34069);
or U37437 (N_37437,N_33936,N_34113);
nand U37438 (N_37438,N_33701,N_34976);
xor U37439 (N_37439,N_32699,N_33143);
nand U37440 (N_37440,N_34502,N_34866);
nand U37441 (N_37441,N_34315,N_32748);
nor U37442 (N_37442,N_33768,N_33759);
and U37443 (N_37443,N_33246,N_34123);
and U37444 (N_37444,N_34827,N_33010);
nor U37445 (N_37445,N_33842,N_33228);
and U37446 (N_37446,N_32609,N_32985);
or U37447 (N_37447,N_33581,N_33880);
and U37448 (N_37448,N_34413,N_34112);
nor U37449 (N_37449,N_32846,N_34222);
xor U37450 (N_37450,N_33875,N_33158);
nand U37451 (N_37451,N_33294,N_33915);
and U37452 (N_37452,N_32766,N_33247);
and U37453 (N_37453,N_34834,N_33528);
and U37454 (N_37454,N_32644,N_34335);
nor U37455 (N_37455,N_33483,N_32581);
and U37456 (N_37456,N_33656,N_34487);
or U37457 (N_37457,N_34669,N_33196);
xor U37458 (N_37458,N_32836,N_34304);
and U37459 (N_37459,N_33724,N_33900);
or U37460 (N_37460,N_34720,N_33739);
nor U37461 (N_37461,N_33143,N_33713);
xor U37462 (N_37462,N_33599,N_32907);
nand U37463 (N_37463,N_34480,N_34660);
and U37464 (N_37464,N_34940,N_33436);
nand U37465 (N_37465,N_34492,N_33486);
nor U37466 (N_37466,N_34137,N_33040);
nand U37467 (N_37467,N_34153,N_33475);
and U37468 (N_37468,N_34341,N_33208);
nor U37469 (N_37469,N_34018,N_34664);
or U37470 (N_37470,N_32523,N_32592);
or U37471 (N_37471,N_34913,N_32518);
nand U37472 (N_37472,N_34090,N_33797);
and U37473 (N_37473,N_33297,N_33161);
nor U37474 (N_37474,N_34146,N_34466);
nand U37475 (N_37475,N_33629,N_34518);
and U37476 (N_37476,N_34150,N_34226);
or U37477 (N_37477,N_32584,N_33632);
nand U37478 (N_37478,N_33780,N_32998);
nor U37479 (N_37479,N_34406,N_33233);
xor U37480 (N_37480,N_34007,N_33837);
or U37481 (N_37481,N_33627,N_32613);
nand U37482 (N_37482,N_34547,N_33752);
nor U37483 (N_37483,N_32894,N_34652);
nand U37484 (N_37484,N_32988,N_33554);
and U37485 (N_37485,N_33445,N_34522);
or U37486 (N_37486,N_32961,N_32599);
or U37487 (N_37487,N_32630,N_34313);
or U37488 (N_37488,N_32735,N_32500);
or U37489 (N_37489,N_33624,N_34717);
or U37490 (N_37490,N_34030,N_32840);
nand U37491 (N_37491,N_32947,N_32618);
nor U37492 (N_37492,N_33844,N_33617);
or U37493 (N_37493,N_34257,N_33367);
or U37494 (N_37494,N_33149,N_34525);
nand U37495 (N_37495,N_34139,N_33541);
and U37496 (N_37496,N_32946,N_33517);
nand U37497 (N_37497,N_32689,N_33027);
xnor U37498 (N_37498,N_34477,N_34993);
nand U37499 (N_37499,N_32923,N_33428);
or U37500 (N_37500,N_36529,N_35470);
and U37501 (N_37501,N_35825,N_35147);
xor U37502 (N_37502,N_36294,N_36199);
nor U37503 (N_37503,N_35542,N_37166);
nand U37504 (N_37504,N_35175,N_35808);
and U37505 (N_37505,N_37318,N_36342);
and U37506 (N_37506,N_36335,N_36413);
and U37507 (N_37507,N_35894,N_36740);
nand U37508 (N_37508,N_35251,N_37143);
xor U37509 (N_37509,N_37478,N_37025);
nand U37510 (N_37510,N_36822,N_37177);
xor U37511 (N_37511,N_35543,N_36912);
and U37512 (N_37512,N_35621,N_36557);
nand U37513 (N_37513,N_37098,N_37003);
nor U37514 (N_37514,N_37195,N_35582);
nor U37515 (N_37515,N_36119,N_35828);
nor U37516 (N_37516,N_37454,N_37404);
nand U37517 (N_37517,N_35047,N_36428);
xnor U37518 (N_37518,N_37191,N_37043);
or U37519 (N_37519,N_36861,N_35136);
nand U37520 (N_37520,N_36215,N_35066);
and U37521 (N_37521,N_35286,N_37137);
nor U37522 (N_37522,N_35193,N_37226);
nor U37523 (N_37523,N_35109,N_36799);
nor U37524 (N_37524,N_35763,N_36584);
nor U37525 (N_37525,N_36130,N_35531);
and U37526 (N_37526,N_35197,N_35395);
and U37527 (N_37527,N_35586,N_36600);
nand U37528 (N_37528,N_35304,N_35740);
nand U37529 (N_37529,N_37299,N_36292);
or U37530 (N_37530,N_35669,N_36061);
nor U37531 (N_37531,N_35213,N_35300);
xnor U37532 (N_37532,N_37080,N_37475);
nand U37533 (N_37533,N_35830,N_37261);
and U37534 (N_37534,N_36873,N_35823);
and U37535 (N_37535,N_36709,N_35118);
nor U37536 (N_37536,N_35003,N_35559);
or U37537 (N_37537,N_35617,N_35581);
xnor U37538 (N_37538,N_36945,N_36323);
nand U37539 (N_37539,N_36089,N_37497);
nor U37540 (N_37540,N_37019,N_36427);
or U37541 (N_37541,N_36242,N_36574);
nor U37542 (N_37542,N_35496,N_35489);
nand U37543 (N_37543,N_35218,N_36743);
or U37544 (N_37544,N_36484,N_36804);
nand U37545 (N_37545,N_36990,N_36620);
and U37546 (N_37546,N_35195,N_37124);
and U37547 (N_37547,N_37060,N_35523);
nor U37548 (N_37548,N_35231,N_36312);
nand U37549 (N_37549,N_35524,N_35296);
nand U37550 (N_37550,N_35682,N_37348);
or U37551 (N_37551,N_36689,N_37131);
nor U37552 (N_37552,N_36617,N_35051);
and U37553 (N_37553,N_36223,N_36702);
nor U37554 (N_37554,N_37198,N_35796);
nand U37555 (N_37555,N_35623,N_35842);
nand U37556 (N_37556,N_35292,N_36004);
nor U37557 (N_37557,N_37008,N_35095);
xnor U37558 (N_37558,N_36103,N_36008);
nor U37559 (N_37559,N_35941,N_37259);
nor U37560 (N_37560,N_35172,N_36001);
or U37561 (N_37561,N_36489,N_37160);
or U37562 (N_37562,N_36553,N_35098);
nor U37563 (N_37563,N_36576,N_36791);
and U37564 (N_37564,N_36346,N_35085);
xor U37565 (N_37565,N_37347,N_37040);
xnor U37566 (N_37566,N_36712,N_35865);
or U37567 (N_37567,N_37213,N_35848);
xor U37568 (N_37568,N_36780,N_35918);
and U37569 (N_37569,N_35824,N_35752);
or U37570 (N_37570,N_35431,N_36338);
nand U37571 (N_37571,N_35082,N_35616);
and U37572 (N_37572,N_35539,N_35155);
xor U37573 (N_37573,N_37157,N_36601);
and U37574 (N_37574,N_36925,N_35746);
nand U37575 (N_37575,N_35603,N_35441);
nand U37576 (N_37576,N_36858,N_36905);
xor U37577 (N_37577,N_37422,N_37158);
or U37578 (N_37578,N_35913,N_36979);
nor U37579 (N_37579,N_35281,N_35955);
nor U37580 (N_37580,N_35620,N_35505);
nand U37581 (N_37581,N_35233,N_35159);
and U37582 (N_37582,N_36101,N_35593);
or U37583 (N_37583,N_35550,N_37076);
nor U37584 (N_37584,N_35897,N_36632);
nand U37585 (N_37585,N_37114,N_35312);
nand U37586 (N_37586,N_36118,N_35378);
nor U37587 (N_37587,N_35856,N_36759);
and U37588 (N_37588,N_35417,N_35203);
and U37589 (N_37589,N_37267,N_36677);
nor U37590 (N_37590,N_36835,N_35374);
or U37591 (N_37591,N_36781,N_35475);
nor U37592 (N_37592,N_35349,N_35498);
nor U37593 (N_37593,N_37310,N_36081);
and U37594 (N_37594,N_37154,N_36286);
xor U37595 (N_37595,N_37009,N_37304);
and U37596 (N_37596,N_37345,N_36234);
nor U37597 (N_37597,N_37439,N_35259);
nand U37598 (N_37598,N_36871,N_36830);
or U37599 (N_37599,N_36594,N_36832);
nand U37600 (N_37600,N_35812,N_35833);
and U37601 (N_37601,N_36167,N_35392);
or U37602 (N_37602,N_36104,N_36284);
nand U37603 (N_37603,N_36967,N_35210);
nand U37604 (N_37604,N_35912,N_37051);
nand U37605 (N_37605,N_36051,N_37321);
and U37606 (N_37606,N_36706,N_35841);
and U37607 (N_37607,N_35090,N_35948);
xnor U37608 (N_37608,N_35450,N_35403);
nor U37609 (N_37609,N_35507,N_35872);
nor U37610 (N_37610,N_36634,N_37207);
nor U37611 (N_37611,N_35692,N_35696);
and U37612 (N_37612,N_36604,N_36980);
nor U37613 (N_37613,N_36813,N_35226);
and U37614 (N_37614,N_36650,N_35027);
or U37615 (N_37615,N_37190,N_36828);
xnor U37616 (N_37616,N_35555,N_35990);
nand U37617 (N_37617,N_36193,N_36341);
and U37618 (N_37618,N_36825,N_36394);
or U37619 (N_37619,N_35837,N_36356);
and U37620 (N_37620,N_36085,N_35774);
or U37621 (N_37621,N_35334,N_36416);
nor U37622 (N_37622,N_35921,N_35803);
and U37623 (N_37623,N_37353,N_36672);
or U37624 (N_37624,N_35444,N_35923);
nor U37625 (N_37625,N_35693,N_36908);
or U37626 (N_37626,N_37017,N_37322);
or U37627 (N_37627,N_36451,N_35704);
or U37628 (N_37628,N_36571,N_35722);
nand U37629 (N_37629,N_36724,N_36329);
or U37630 (N_37630,N_35922,N_35119);
nor U37631 (N_37631,N_36330,N_37020);
nor U37632 (N_37632,N_36836,N_35942);
nand U37633 (N_37633,N_35255,N_36433);
nand U37634 (N_37634,N_35084,N_36239);
and U37635 (N_37635,N_37397,N_36315);
nor U37636 (N_37636,N_36477,N_37185);
and U37637 (N_37637,N_36090,N_35002);
xor U37638 (N_37638,N_35769,N_36555);
and U37639 (N_37639,N_36847,N_37334);
and U37640 (N_37640,N_37270,N_36889);
nand U37641 (N_37641,N_35293,N_35951);
nor U37642 (N_37642,N_37385,N_35855);
and U37643 (N_37643,N_35646,N_36705);
and U37644 (N_37644,N_36269,N_35310);
xor U37645 (N_37645,N_37390,N_36808);
xnor U37646 (N_37646,N_35198,N_35663);
or U37647 (N_37647,N_36088,N_37180);
nor U37648 (N_37648,N_35199,N_37168);
nor U37649 (N_37649,N_35329,N_36038);
nor U37650 (N_37650,N_36996,N_37193);
nand U37651 (N_37651,N_35919,N_35584);
and U37652 (N_37652,N_36638,N_35468);
nor U37653 (N_37653,N_36408,N_36875);
and U37654 (N_37654,N_37273,N_36328);
nor U37655 (N_37655,N_36640,N_35326);
nor U37656 (N_37656,N_35303,N_35479);
nor U37657 (N_37657,N_36974,N_37256);
xnor U37658 (N_37658,N_37028,N_35430);
or U37659 (N_37659,N_35510,N_37292);
or U37660 (N_37660,N_36448,N_36998);
or U37661 (N_37661,N_37389,N_36078);
xnor U37662 (N_37662,N_36044,N_36045);
and U37663 (N_37663,N_36100,N_35548);
nand U37664 (N_37664,N_37225,N_36073);
or U37665 (N_37665,N_37332,N_35654);
or U37666 (N_37666,N_36107,N_36157);
or U37667 (N_37667,N_37377,N_35228);
nor U37668 (N_37668,N_37372,N_35173);
nand U37669 (N_37669,N_37361,N_35766);
or U37670 (N_37670,N_36497,N_37352);
and U37671 (N_37671,N_36578,N_35596);
nand U37672 (N_37672,N_36610,N_35836);
nand U37673 (N_37673,N_35698,N_36521);
or U37674 (N_37674,N_36469,N_36375);
or U37675 (N_37675,N_36019,N_36520);
nand U37676 (N_37676,N_36492,N_35151);
xnor U37677 (N_37677,N_35628,N_37314);
and U37678 (N_37678,N_35989,N_36391);
and U37679 (N_37679,N_36915,N_36172);
nor U37680 (N_37680,N_35052,N_37083);
or U37681 (N_37681,N_35362,N_36953);
nor U37682 (N_37682,N_35831,N_36210);
and U37683 (N_37683,N_35045,N_35860);
and U37684 (N_37684,N_35854,N_35284);
nor U37685 (N_37685,N_36499,N_35914);
and U37686 (N_37686,N_36788,N_36271);
or U37687 (N_37687,N_35979,N_36570);
and U37688 (N_37688,N_36994,N_36374);
or U37689 (N_37689,N_37159,N_37142);
nor U37690 (N_37690,N_36093,N_37209);
or U37691 (N_37691,N_35443,N_35471);
or U37692 (N_37692,N_37243,N_36802);
nand U37693 (N_37693,N_36968,N_36538);
or U37694 (N_37694,N_37224,N_37184);
or U37695 (N_37695,N_36961,N_35017);
nand U37696 (N_37696,N_36854,N_36755);
nor U37697 (N_37697,N_37179,N_35217);
and U37698 (N_37698,N_36083,N_37471);
or U37699 (N_37699,N_35071,N_36603);
or U37700 (N_37700,N_35375,N_36295);
nor U37701 (N_37701,N_36868,N_35762);
and U37702 (N_37702,N_36462,N_35414);
nor U37703 (N_37703,N_35360,N_35689);
nor U37704 (N_37704,N_35216,N_35194);
or U37705 (N_37705,N_35956,N_36774);
nor U37706 (N_37706,N_36411,N_36176);
nor U37707 (N_37707,N_37097,N_36704);
nand U37708 (N_37708,N_37441,N_36815);
or U37709 (N_37709,N_35074,N_36692);
nand U37710 (N_37710,N_35120,N_37230);
nand U37711 (N_37711,N_35633,N_36343);
nand U37712 (N_37712,N_35130,N_37127);
xor U37713 (N_37713,N_36886,N_36568);
nor U37714 (N_37714,N_37424,N_35925);
and U37715 (N_37715,N_35315,N_36674);
or U37716 (N_37716,N_35985,N_37487);
or U37717 (N_37717,N_35469,N_35037);
nand U37718 (N_37718,N_36153,N_36695);
nor U37719 (N_37719,N_35248,N_37489);
nand U37720 (N_37720,N_36931,N_36919);
or U37721 (N_37721,N_37410,N_35567);
nand U37722 (N_37722,N_37455,N_36734);
nand U37723 (N_37723,N_35062,N_36410);
or U37724 (N_37724,N_35018,N_36765);
or U37725 (N_37725,N_37032,N_36987);
and U37726 (N_37726,N_36645,N_36397);
and U37727 (N_37727,N_35322,N_37447);
nor U37728 (N_37728,N_37434,N_35573);
or U37729 (N_37729,N_37182,N_35535);
nor U37730 (N_37730,N_35685,N_36591);
or U37731 (N_37731,N_36426,N_36707);
or U37732 (N_37732,N_35088,N_36097);
and U37733 (N_37733,N_35010,N_35289);
nand U37734 (N_37734,N_37286,N_37470);
nand U37735 (N_37735,N_36062,N_36137);
xor U37736 (N_37736,N_35318,N_37363);
nor U37737 (N_37737,N_35647,N_36794);
nor U37738 (N_37738,N_36778,N_35008);
or U37739 (N_37739,N_36259,N_37388);
and U37740 (N_37740,N_35641,N_35827);
or U37741 (N_37741,N_35602,N_35517);
or U37742 (N_37742,N_35401,N_35004);
nand U37743 (N_37743,N_35892,N_37045);
nor U37744 (N_37744,N_37350,N_37088);
and U37745 (N_37745,N_37050,N_36279);
or U37746 (N_37746,N_35046,N_37281);
nand U37747 (N_37747,N_36454,N_36091);
nor U37748 (N_37748,N_36291,N_35342);
or U37749 (N_37749,N_36727,N_37414);
and U37750 (N_37750,N_37403,N_36726);
or U37751 (N_37751,N_36586,N_35648);
and U37752 (N_37752,N_37162,N_37092);
or U37753 (N_37753,N_36249,N_35274);
nand U37754 (N_37754,N_36068,N_36527);
nor U37755 (N_37755,N_36962,N_37467);
nand U37756 (N_37756,N_35664,N_35954);
nor U37757 (N_37757,N_36055,N_36934);
nand U37758 (N_37758,N_36457,N_37284);
nor U37759 (N_37759,N_35768,N_36444);
and U37760 (N_37760,N_36404,N_36685);
or U37761 (N_37761,N_37202,N_36798);
nor U37762 (N_37762,N_36892,N_35133);
or U37763 (N_37763,N_37399,N_36652);
and U37764 (N_37764,N_36053,N_36764);
or U37765 (N_37765,N_36123,N_35670);
or U37766 (N_37766,N_35592,N_35600);
and U37767 (N_37767,N_36885,N_36367);
and U37768 (N_37768,N_37250,N_36377);
or U37769 (N_37769,N_35439,N_35929);
or U37770 (N_37770,N_36503,N_36487);
or U37771 (N_37771,N_36385,N_35684);
nor U37772 (N_37772,N_37375,N_35667);
and U37773 (N_37773,N_35960,N_35207);
nor U37774 (N_37774,N_35554,N_37477);
nand U37775 (N_37775,N_36441,N_35562);
nor U37776 (N_37776,N_35566,N_35934);
or U37777 (N_37777,N_35308,N_36547);
nand U37778 (N_37778,N_37498,N_36869);
and U37779 (N_37779,N_37445,N_36616);
and U37780 (N_37780,N_35904,N_37016);
xnor U37781 (N_37781,N_36579,N_37435);
xor U37782 (N_37782,N_36029,N_36633);
nand U37783 (N_37783,N_35819,N_36627);
and U37784 (N_37784,N_36659,N_36370);
and U37785 (N_37785,N_35427,N_35797);
or U37786 (N_37786,N_35552,N_35787);
nor U37787 (N_37787,N_36033,N_35939);
xor U37788 (N_37788,N_36753,N_35643);
nor U37789 (N_37789,N_37462,N_35858);
or U37790 (N_37790,N_37205,N_36461);
and U37791 (N_37791,N_37287,N_37176);
nor U37792 (N_37792,N_36420,N_37457);
and U37793 (N_37793,N_35116,N_37163);
nand U37794 (N_37794,N_36725,N_36296);
nand U37795 (N_37795,N_35246,N_36253);
or U37796 (N_37796,N_35634,N_37094);
or U37797 (N_37797,N_37105,N_35278);
or U37798 (N_37798,N_36219,N_36324);
and U37799 (N_37799,N_36893,N_36003);
and U37800 (N_37800,N_35391,N_37164);
or U37801 (N_37801,N_37242,N_37188);
or U37802 (N_37802,N_35258,N_36658);
nor U37803 (N_37803,N_35314,N_35813);
nor U37804 (N_37804,N_37161,N_35723);
and U37805 (N_37805,N_37129,N_36422);
nand U37806 (N_37806,N_36120,N_37476);
or U37807 (N_37807,N_36163,N_35619);
xor U37808 (N_37808,N_36720,N_36195);
nor U37809 (N_37809,N_36630,N_35908);
and U37810 (N_37810,N_37279,N_35782);
nor U37811 (N_37811,N_36010,N_35578);
xnor U37812 (N_37812,N_35741,N_35168);
xnor U37813 (N_37813,N_37373,N_35866);
xnor U37814 (N_37814,N_35614,N_37264);
and U37815 (N_37815,N_37355,N_36299);
or U37816 (N_37816,N_36285,N_35393);
or U37817 (N_37817,N_36403,N_36949);
nand U37818 (N_37818,N_35984,N_36673);
nor U37819 (N_37819,N_35672,N_37071);
and U37820 (N_37820,N_36087,N_37326);
or U37821 (N_37821,N_36216,N_36818);
xnor U37822 (N_37822,N_35958,N_37418);
or U37823 (N_37823,N_37208,N_37252);
xor U37824 (N_37824,N_37062,N_35805);
nor U37825 (N_37825,N_35232,N_35745);
and U37826 (N_37826,N_35126,N_37432);
nor U37827 (N_37827,N_35013,N_36595);
or U37828 (N_37828,N_36544,N_37089);
nor U37829 (N_37829,N_35515,N_36429);
nor U37830 (N_37830,N_36878,N_37150);
nor U37831 (N_37831,N_36840,N_36151);
or U37832 (N_37832,N_36509,N_35466);
nor U37833 (N_37833,N_35264,N_36516);
or U37834 (N_37834,N_35324,N_36070);
or U37835 (N_37835,N_35732,N_37419);
and U37836 (N_37836,N_36981,N_37054);
or U37837 (N_37837,N_37362,N_35844);
and U37838 (N_37838,N_35590,N_36959);
or U37839 (N_37839,N_35164,N_36845);
nand U37840 (N_37840,N_35760,N_36988);
nand U37841 (N_37841,N_37496,N_35177);
nor U37842 (N_37842,N_36504,N_36843);
nand U37843 (N_37843,N_36749,N_35834);
and U37844 (N_37844,N_35112,N_36665);
or U37845 (N_37845,N_35055,N_35270);
nor U37846 (N_37846,N_36510,N_37049);
nor U37847 (N_37847,N_36738,N_35716);
nor U37848 (N_37848,N_36471,N_36214);
or U37849 (N_37849,N_36711,N_35765);
or U37850 (N_37850,N_37244,N_37211);
nor U37851 (N_37851,N_36201,N_35871);
nand U37852 (N_37852,N_36230,N_37147);
nand U37853 (N_37853,N_36537,N_35815);
nor U37854 (N_37854,N_36648,N_36144);
or U37855 (N_37855,N_36663,N_37479);
and U37856 (N_37856,N_36635,N_36190);
xnor U37857 (N_37857,N_37030,N_35452);
and U37858 (N_37858,N_35537,N_36275);
nor U37859 (N_37859,N_36754,N_35793);
or U37860 (N_37860,N_35068,N_36517);
nand U37861 (N_37861,N_36014,N_35712);
and U37862 (N_37862,N_36577,N_36252);
nand U37863 (N_37863,N_35840,N_35072);
and U37864 (N_37864,N_36552,N_36336);
and U37865 (N_37865,N_36588,N_35309);
nand U37866 (N_37866,N_35553,N_36564);
xnor U37867 (N_37867,N_36697,N_36389);
or U37868 (N_37868,N_36647,N_36768);
nand U37869 (N_37869,N_35843,N_36913);
xor U37870 (N_37870,N_35208,N_37012);
and U37871 (N_37871,N_35212,N_35783);
and U37872 (N_37872,N_36866,N_35327);
nor U37873 (N_37873,N_35546,N_35316);
nor U37874 (N_37874,N_36842,N_35178);
nor U37875 (N_37875,N_36418,N_35019);
nor U37876 (N_37876,N_37265,N_36926);
nor U37877 (N_37877,N_36020,N_35005);
and U37878 (N_37878,N_37282,N_35012);
and U37879 (N_37879,N_35601,N_35371);
or U37880 (N_37880,N_35477,N_35968);
nand U37881 (N_37881,N_36146,N_35191);
nor U37882 (N_37882,N_36668,N_35273);
nand U37883 (N_37883,N_37319,N_36823);
nand U37884 (N_37884,N_37301,N_35711);
nand U37885 (N_37885,N_36479,N_36614);
or U37886 (N_37886,N_37113,N_36948);
or U37887 (N_37887,N_35887,N_37215);
or U37888 (N_37888,N_36009,N_36475);
nand U37889 (N_37889,N_35369,N_35454);
or U37890 (N_37890,N_35429,N_36362);
nor U37891 (N_37891,N_35511,N_35291);
or U37892 (N_37892,N_36969,N_35145);
nor U37893 (N_37893,N_35041,N_35649);
nor U37894 (N_37894,N_36699,N_35026);
and U37895 (N_37895,N_36265,N_36183);
or U37896 (N_37896,N_35049,N_36606);
nand U37897 (N_37897,N_35952,N_35000);
and U37898 (N_37898,N_35087,N_36972);
or U37899 (N_37899,N_35038,N_36501);
and U37900 (N_37900,N_36072,N_36863);
nor U37901 (N_37901,N_36716,N_37070);
or U37902 (N_37902,N_36174,N_36752);
nor U37903 (N_37903,N_36540,N_36899);
nor U37904 (N_37904,N_35632,N_35933);
xor U37905 (N_37905,N_36125,N_37075);
or U37906 (N_37906,N_36181,N_36751);
nand U37907 (N_37907,N_36358,N_35972);
and U37908 (N_37908,N_36874,N_36746);
nand U37909 (N_37909,N_35238,N_36227);
or U37910 (N_37910,N_36450,N_36278);
or U37911 (N_37911,N_37135,N_36793);
or U37912 (N_37912,N_37383,N_36327);
nor U37913 (N_37913,N_35551,N_36762);
nor U37914 (N_37914,N_36316,N_35743);
or U37915 (N_37915,N_36850,N_37084);
and U37916 (N_37916,N_36491,N_37459);
xnor U37917 (N_37917,N_36563,N_35405);
and U37918 (N_37918,N_35434,N_37364);
xnor U37919 (N_37919,N_37172,N_35736);
or U37920 (N_37920,N_36322,N_35335);
or U37921 (N_37921,N_36363,N_36565);
nor U37922 (N_37922,N_36841,N_35142);
nand U37923 (N_37923,N_37116,N_36985);
and U37924 (N_37924,N_36519,N_36071);
nor U37925 (N_37925,N_36430,N_35379);
nor U37926 (N_37926,N_35859,N_36026);
nand U37927 (N_37927,N_36852,N_36117);
or U37928 (N_37928,N_35404,N_35626);
or U37929 (N_37929,N_35307,N_36349);
and U37930 (N_37930,N_35675,N_35236);
or U37931 (N_37931,N_36918,N_37450);
and U37932 (N_37932,N_36896,N_35157);
or U37933 (N_37933,N_36927,N_35635);
or U37934 (N_37934,N_36340,N_36870);
and U37935 (N_37935,N_35104,N_37338);
and U37936 (N_37936,N_35656,N_35905);
nor U37937 (N_37937,N_36007,N_35458);
or U37938 (N_37938,N_37240,N_37181);
nand U37939 (N_37939,N_36069,N_35478);
nor U37940 (N_37940,N_35180,N_37472);
nor U37941 (N_37941,N_36277,N_37067);
and U37942 (N_37942,N_36392,N_36760);
nor U37943 (N_37943,N_35416,N_36680);
nand U37944 (N_37944,N_37153,N_36867);
and U37945 (N_37945,N_36459,N_37354);
or U37946 (N_37946,N_36795,N_36453);
nand U37947 (N_37947,N_35575,N_37351);
nor U37948 (N_37948,N_36446,N_36928);
nor U37949 (N_37949,N_35791,N_35986);
nand U37950 (N_37950,N_35677,N_37149);
xnor U37951 (N_37951,N_35227,N_35402);
nor U37952 (N_37952,N_35868,N_37433);
nor U37953 (N_37953,N_35863,N_36732);
and U37954 (N_37954,N_37342,N_35651);
nor U37955 (N_37955,N_37401,N_36801);
or U37956 (N_37956,N_36447,N_35758);
nor U37957 (N_37957,N_36582,N_36102);
nor U37958 (N_37958,N_36386,N_37241);
nor U37959 (N_37959,N_35294,N_36952);
nor U37960 (N_37960,N_36364,N_36733);
or U37961 (N_37961,N_36115,N_37484);
nor U37962 (N_37962,N_36351,N_35418);
nand U37963 (N_37963,N_35792,N_37438);
nor U37964 (N_37964,N_36139,N_37307);
xnor U37965 (N_37965,N_35560,N_37288);
or U37966 (N_37966,N_37011,N_37278);
nand U37967 (N_37967,N_35209,N_36785);
and U37968 (N_37968,N_36621,N_35604);
nor U37969 (N_37969,N_36406,N_36378);
or U37970 (N_37970,N_37041,N_37442);
nand U37971 (N_37971,N_35338,N_35987);
and U37972 (N_37972,N_36182,N_36145);
nand U37973 (N_37973,N_36637,N_35637);
nand U37974 (N_37974,N_35901,N_35247);
xor U37975 (N_37975,N_36047,N_35476);
nor U37976 (N_37976,N_36623,N_35200);
nor U37977 (N_37977,N_35211,N_36525);
xor U37978 (N_37978,N_35297,N_36046);
or U37979 (N_37979,N_36016,N_35370);
xnor U37980 (N_37980,N_35124,N_36483);
or U37981 (N_37981,N_37134,N_36463);
or U37982 (N_37982,N_35170,N_37469);
nor U37983 (N_37983,N_36439,N_35927);
nor U37984 (N_37984,N_36826,N_35719);
nand U37985 (N_37985,N_35150,N_37376);
nand U37986 (N_37986,N_37056,N_35482);
nor U37987 (N_37987,N_35742,N_37223);
and U37988 (N_37988,N_36466,N_36941);
or U37989 (N_37989,N_36436,N_35015);
or U37990 (N_37990,N_35364,N_35202);
nor U37991 (N_37991,N_37405,N_35845);
and U37992 (N_37992,N_36993,N_35563);
or U37993 (N_37993,N_36465,N_36023);
nand U37994 (N_37994,N_36728,N_36131);
and U37995 (N_37995,N_36098,N_35165);
nor U37996 (N_37996,N_35382,N_37408);
and U37997 (N_37997,N_36831,N_35048);
and U37998 (N_37998,N_36856,N_37238);
nand U37999 (N_37999,N_35810,N_35389);
and U38000 (N_38000,N_37323,N_37371);
nor U38001 (N_38001,N_35816,N_35261);
and U38002 (N_38002,N_35260,N_36587);
nand U38003 (N_38003,N_35028,N_35893);
and U38004 (N_38004,N_36084,N_36901);
nand U38005 (N_38005,N_37210,N_35492);
nand U38006 (N_38006,N_35295,N_37144);
nand U38007 (N_38007,N_36718,N_36359);
or U38008 (N_38008,N_35789,N_35093);
nor U38009 (N_38009,N_36846,N_37429);
nor U38010 (N_38010,N_36231,N_35588);
nand U38011 (N_38011,N_36964,N_35911);
nand U38012 (N_38012,N_36951,N_37115);
or U38013 (N_38013,N_36498,N_35847);
or U38014 (N_38014,N_36470,N_37233);
or U38015 (N_38015,N_35453,N_36670);
nor U38016 (N_38016,N_36177,N_36025);
nor U38017 (N_38017,N_35493,N_35396);
nor U38018 (N_38018,N_36589,N_36569);
nand U38019 (N_38019,N_36095,N_37068);
nor U38020 (N_38020,N_36387,N_35472);
and U38021 (N_38021,N_37170,N_35606);
or U38022 (N_38022,N_35386,N_35257);
and U38023 (N_38023,N_35680,N_37053);
xnor U38024 (N_38024,N_35595,N_37253);
xnor U38025 (N_38025,N_36302,N_36467);
or U38026 (N_38026,N_36664,N_37010);
nor U38027 (N_38027,N_36353,N_37298);
nor U38028 (N_38028,N_36715,N_35446);
and U38029 (N_38029,N_36803,N_35328);
or U38030 (N_38030,N_36661,N_36297);
nand U38031 (N_38031,N_36615,N_36383);
nand U38032 (N_38032,N_36766,N_36188);
nor U38033 (N_38033,N_37346,N_36405);
nand U38034 (N_38034,N_36175,N_37033);
and U38035 (N_38035,N_35121,N_36272);
nand U38036 (N_38036,N_36369,N_35179);
or U38037 (N_38037,N_35678,N_36897);
and U38038 (N_38038,N_37123,N_36522);
or U38039 (N_38039,N_37263,N_36320);
or U38040 (N_38040,N_35313,N_35244);
nand U38041 (N_38041,N_35081,N_35140);
or U38042 (N_38042,N_35501,N_35245);
or U38043 (N_38043,N_37411,N_35290);
or U38044 (N_38044,N_37473,N_36222);
nand U38045 (N_38045,N_35755,N_36776);
nand U38046 (N_38046,N_36065,N_35661);
nor U38047 (N_38047,N_37141,N_36162);
xnor U38048 (N_38048,N_37126,N_37339);
and U38049 (N_38049,N_36233,N_35407);
nand U38050 (N_38050,N_35024,N_36414);
and U38051 (N_38051,N_37189,N_37206);
or U38052 (N_38052,N_35388,N_35445);
nor U38053 (N_38053,N_36771,N_36700);
nand U38054 (N_38054,N_35148,N_36236);
nor U38055 (N_38055,N_36360,N_36124);
nor U38056 (N_38056,N_37294,N_35306);
and U38057 (N_38057,N_35101,N_37290);
xor U38058 (N_38058,N_36947,N_35001);
xnor U38059 (N_38059,N_35920,N_35618);
or U38060 (N_38060,N_36380,N_35738);
or U38061 (N_38061,N_36942,N_36099);
nor U38062 (N_38062,N_36197,N_36769);
or U38063 (N_38063,N_35756,N_37400);
or U38064 (N_38064,N_35609,N_36485);
xnor U38065 (N_38065,N_35448,N_37395);
nand U38066 (N_38066,N_36154,N_35353);
or U38067 (N_38067,N_37231,N_36950);
nand U38068 (N_38068,N_36274,N_36696);
nand U38069 (N_38069,N_35973,N_36810);
and U38070 (N_38070,N_37194,N_35924);
and U38071 (N_38071,N_35525,N_35549);
and U38072 (N_38072,N_35638,N_35384);
or U38073 (N_38073,N_36423,N_36879);
nand U38074 (N_38074,N_37249,N_35190);
nand U38075 (N_38075,N_37167,N_37111);
or U38076 (N_38076,N_35850,N_35262);
nand U38077 (N_38077,N_35671,N_35583);
nand U38078 (N_38078,N_36220,N_36622);
nand U38079 (N_38079,N_36936,N_37456);
xor U38080 (N_38080,N_35978,N_35381);
nor U38081 (N_38081,N_35139,N_35330);
nor U38082 (N_38082,N_36671,N_37421);
nor U38083 (N_38083,N_35484,N_37343);
nand U38084 (N_38084,N_35486,N_36114);
nor U38085 (N_38085,N_37024,N_36357);
nor U38086 (N_38086,N_35702,N_36347);
nand U38087 (N_38087,N_35718,N_37148);
or U38088 (N_38088,N_36057,N_37327);
and U38089 (N_38089,N_36445,N_35709);
and U38090 (N_38090,N_35214,N_36957);
or U38091 (N_38091,N_37118,N_37413);
and U38092 (N_38092,N_35645,N_36864);
nor U38093 (N_38093,N_35864,N_36602);
nand U38094 (N_38094,N_35891,N_36562);
and U38095 (N_38095,N_37274,N_37090);
or U38096 (N_38096,N_35714,N_35154);
nor U38097 (N_38097,N_35852,N_36687);
xor U38098 (N_38098,N_36108,N_37464);
nand U38099 (N_38099,N_35778,N_35967);
and U38100 (N_38100,N_35215,N_35132);
or U38101 (N_38101,N_35237,N_36412);
and U38102 (N_38102,N_36597,N_35976);
and U38103 (N_38103,N_37335,N_36005);
and U38104 (N_38104,N_36140,N_37027);
or U38105 (N_38105,N_36824,N_36368);
nand U38106 (N_38106,N_37276,N_37186);
and U38107 (N_38107,N_36141,N_36399);
nor U38108 (N_38108,N_37101,N_37295);
or U38109 (N_38109,N_35737,N_37133);
nor U38110 (N_38110,N_37396,N_37380);
or U38111 (N_38111,N_35729,N_36682);
nand U38112 (N_38112,N_36737,N_37481);
xnor U38113 (N_38113,N_35749,N_35589);
and U38114 (N_38114,N_36703,N_36390);
nor U38115 (N_38115,N_37140,N_37023);
or U38116 (N_38116,N_35376,N_35415);
nor U38117 (N_38117,N_35639,N_37069);
and U38118 (N_38118,N_35561,N_35467);
and U38119 (N_38119,N_36877,N_36937);
and U38120 (N_38120,N_35903,N_37406);
and U38121 (N_38121,N_37437,N_37258);
or U38122 (N_38122,N_36432,N_35413);
and U38123 (N_38123,N_35694,N_36898);
and U38124 (N_38124,N_36807,N_36678);
nand U38125 (N_38125,N_35761,N_35720);
nand U38126 (N_38126,N_35556,N_37128);
nand U38127 (N_38127,N_35818,N_37047);
nor U38128 (N_38128,N_36207,N_35683);
and U38129 (N_38129,N_36880,N_36618);
nor U38130 (N_38130,N_37156,N_35063);
and U38131 (N_38131,N_37064,N_36922);
nand U38132 (N_38132,N_36407,N_37104);
or U38133 (N_38133,N_36455,N_36419);
and U38134 (N_38134,N_35039,N_35896);
xnor U38135 (N_38135,N_36513,N_36229);
xnor U38136 (N_38136,N_36398,N_35801);
or U38137 (N_38137,N_36742,N_35530);
nand U38138 (N_38138,N_37038,N_35994);
nand U38139 (N_38139,N_35096,N_35461);
nand U38140 (N_38140,N_35506,N_36192);
and U38141 (N_38141,N_36923,N_36844);
or U38142 (N_38142,N_36160,N_36739);
and U38143 (N_38143,N_35715,N_36321);
nand U38144 (N_38144,N_36554,N_35428);
nor U38145 (N_38145,N_37037,N_35807);
nor U38146 (N_38146,N_36646,N_36168);
nand U38147 (N_38147,N_36611,N_36816);
nor U38148 (N_38148,N_35974,N_35577);
nor U38149 (N_38149,N_36307,N_37187);
nand U38150 (N_38150,N_36556,N_36464);
and U38151 (N_38151,N_37333,N_36723);
nor U38152 (N_38152,N_36502,N_36829);
nand U38153 (N_38153,N_35876,N_36147);
nand U38154 (N_38154,N_35464,N_35953);
nand U38155 (N_38155,N_35161,N_35103);
and U38156 (N_38156,N_36790,N_35707);
and U38157 (N_38157,N_36992,N_36655);
xnor U38158 (N_38158,N_37452,N_37296);
nand U38159 (N_38159,N_36437,N_37200);
nand U38160 (N_38160,N_35611,N_35457);
or U38161 (N_38161,N_35977,N_35011);
nand U38162 (N_38162,N_35187,N_35570);
and U38163 (N_38163,N_36911,N_35534);
nand U38164 (N_38164,N_36654,N_35499);
and U38165 (N_38165,N_35412,N_35359);
or U38166 (N_38166,N_35795,N_37280);
or U38167 (N_38167,N_36545,N_35323);
or U38168 (N_38168,N_35239,N_35372);
and U38169 (N_38169,N_35282,N_37340);
or U38170 (N_38170,N_36958,N_35655);
nor U38171 (N_38171,N_36178,N_35660);
or U38172 (N_38172,N_36558,N_36651);
nand U38173 (N_38173,N_36644,N_35169);
nand U38174 (N_38174,N_36076,N_35069);
nand U38175 (N_38175,N_36493,N_35421);
and U38176 (N_38176,N_36683,N_36944);
and U38177 (N_38177,N_37458,N_36982);
nand U38178 (N_38178,N_36226,N_37359);
nor U38179 (N_38179,N_36121,N_36773);
and U38180 (N_38180,N_36543,N_35144);
nand U38181 (N_38181,N_35057,N_36792);
nand U38182 (N_38182,N_35679,N_36585);
nand U38183 (N_38183,N_37183,N_35995);
nor U38184 (N_38184,N_35181,N_35727);
and U38185 (N_38185,N_35811,N_37146);
or U38186 (N_38186,N_37048,N_35158);
nor U38187 (N_38187,N_35035,N_37145);
and U38188 (N_38188,N_36698,N_35532);
nor U38189 (N_38189,N_35775,N_35332);
and U38190 (N_38190,N_36354,N_35615);
and U38191 (N_38191,N_35757,N_36080);
or U38192 (N_38192,N_36159,N_36657);
or U38193 (N_38193,N_35350,N_36250);
xnor U38194 (N_38194,N_36821,N_37039);
nor U38195 (N_38195,N_35610,N_35363);
or U38196 (N_38196,N_37031,N_36884);
or U38197 (N_38197,N_36806,N_36533);
nand U38198 (N_38198,N_37336,N_36921);
nand U38199 (N_38199,N_35077,N_36667);
xor U38200 (N_38200,N_37416,N_35117);
nor U38201 (N_38201,N_35784,N_37035);
or U38202 (N_38202,N_36138,N_36331);
xnor U38203 (N_38203,N_36196,N_37106);
nand U38204 (N_38204,N_35947,N_35790);
and U38205 (N_38205,N_36750,N_36581);
nand U38206 (N_38206,N_35241,N_37269);
nor U38207 (N_38207,N_35111,N_35050);
and U38208 (N_38208,N_37108,N_35817);
nand U38209 (N_38209,N_35992,N_37349);
nor U38210 (N_38210,N_36817,N_36251);
nand U38211 (N_38211,N_35256,N_35520);
nand U38212 (N_38212,N_35910,N_36745);
nor U38213 (N_38213,N_35138,N_36719);
and U38214 (N_38214,N_35192,N_35673);
nor U38215 (N_38215,N_36666,N_36381);
nor U38216 (N_38216,N_35185,N_36512);
and U38217 (N_38217,N_37197,N_35107);
nand U38218 (N_38218,N_35945,N_37122);
nand U38219 (N_38219,N_35906,N_36995);
or U38220 (N_38220,N_35115,N_37155);
nor U38221 (N_38221,N_37237,N_37444);
xor U38222 (N_38222,N_35770,N_36736);
or U38223 (N_38223,N_37222,N_36317);
nor U38224 (N_38224,N_35337,N_37026);
nor U38225 (N_38225,N_35383,N_36241);
or U38226 (N_38226,N_37365,N_36049);
and U38227 (N_38227,N_35275,N_35234);
nor U38228 (N_38228,N_35870,N_35016);
xnor U38229 (N_38229,N_36656,N_35495);
xnor U38230 (N_38230,N_36914,N_35276);
nand U38231 (N_38231,N_35579,N_37034);
and U38232 (N_38232,N_35750,N_35320);
nor U38233 (N_38233,N_36721,N_35771);
xor U38234 (N_38234,N_36031,N_35073);
or U38235 (N_38235,N_35419,N_35629);
nand U38236 (N_38236,N_36258,N_36938);
or U38237 (N_38237,N_36170,N_37074);
xor U38238 (N_38238,N_35930,N_37398);
nor U38239 (N_38239,N_36415,N_37007);
nand U38240 (N_38240,N_36599,N_37443);
or U38241 (N_38241,N_36876,N_37220);
or U38242 (N_38242,N_35949,N_36366);
nand U38243 (N_38243,N_37004,N_35591);
nand U38244 (N_38244,N_36474,N_35959);
nor U38245 (N_38245,N_35527,N_37109);
and U38246 (N_38246,N_36596,N_37130);
and U38247 (N_38247,N_35385,N_36904);
and U38248 (N_38248,N_36946,N_35127);
or U38249 (N_38249,N_36202,N_37329);
nor U38250 (N_38250,N_35188,N_37218);
xor U38251 (N_38251,N_35565,N_37431);
nor U38252 (N_38252,N_35653,N_35730);
nand U38253 (N_38253,N_37311,N_37331);
and U38254 (N_38254,N_36187,N_36984);
nand U38255 (N_38255,N_36434,N_35409);
nor U38256 (N_38256,N_36975,N_36268);
and U38257 (N_38257,N_37305,N_37103);
nand U38258 (N_38258,N_37214,N_36991);
nand U38259 (N_38259,N_37139,N_36833);
nand U38260 (N_38260,N_36862,N_35345);
nand U38261 (N_38261,N_35250,N_36246);
or U38262 (N_38262,N_37446,N_35059);
nand U38263 (N_38263,N_35176,N_37494);
xnor U38264 (N_38264,N_35174,N_36940);
xor U38265 (N_38265,N_37000,N_35221);
nand U38266 (N_38266,N_36189,N_35344);
nor U38267 (N_38267,N_35442,N_37212);
xor U38268 (N_38268,N_36730,N_36240);
nor U38269 (N_38269,N_35717,N_36401);
nand U38270 (N_38270,N_35252,N_35220);
or U38271 (N_38271,N_37006,N_35435);
or U38272 (N_38272,N_36694,N_37262);
and U38273 (N_38273,N_35886,N_35020);
or U38274 (N_38274,N_36311,N_35594);
nand U38275 (N_38275,N_35564,N_35613);
or U38276 (N_38276,N_35253,N_35043);
xnor U38277 (N_38277,N_36156,N_35713);
nand U38278 (N_38278,N_36289,N_35734);
and U38279 (N_38279,N_37095,N_36508);
nor U38280 (N_38280,N_35229,N_35317);
or U38281 (N_38281,N_35243,N_36326);
and U38282 (N_38282,N_36693,N_35030);
nand U38283 (N_38283,N_36079,N_36135);
nor U38284 (N_38284,N_35806,N_35368);
and U38285 (N_38285,N_37171,N_35285);
or U38286 (N_38286,N_35356,N_36060);
nand U38287 (N_38287,N_35025,N_36690);
and U38288 (N_38288,N_36106,N_36838);
or U38289 (N_38289,N_35503,N_36748);
or U38290 (N_38290,N_37268,N_35219);
or U38291 (N_38291,N_35424,N_37239);
nand U38292 (N_38292,N_35459,N_36303);
or U38293 (N_38293,N_35697,N_36935);
nand U38294 (N_38294,N_36691,N_35036);
and U38295 (N_38295,N_35659,N_35449);
or U38296 (N_38296,N_35465,N_37368);
nor U38297 (N_38297,N_37175,N_35420);
or U38298 (N_38298,N_36973,N_35137);
or U38299 (N_38299,N_36313,N_35267);
xor U38300 (N_38300,N_35277,N_35981);
or U38301 (N_38301,N_37221,N_36613);
nand U38302 (N_38302,N_37366,N_35991);
nor U38303 (N_38303,N_37072,N_35007);
nor U38304 (N_38304,N_37100,N_35205);
or U38305 (N_38305,N_37059,N_36480);
nor U38306 (N_38306,N_37248,N_36989);
xor U38307 (N_38307,N_35451,N_37466);
or U38308 (N_38308,N_35881,N_36848);
nor U38309 (N_38309,N_36203,N_35067);
nand U38310 (N_38310,N_36767,N_36684);
or U38311 (N_38311,N_36701,N_35612);
xnor U38312 (N_38312,N_35666,N_36094);
and U38313 (N_38313,N_35113,N_36247);
nor U38314 (N_38314,N_37436,N_35705);
xor U38315 (N_38315,N_36643,N_36421);
nand U38316 (N_38316,N_35839,N_37219);
or U38317 (N_38317,N_36903,N_36482);
and U38318 (N_38318,N_36626,N_36225);
nand U38319 (N_38319,N_36221,N_36572);
nand U38320 (N_38320,N_36811,N_35283);
nand U38321 (N_38321,N_35587,N_35544);
nor U38322 (N_38322,N_35788,N_36344);
nor U38323 (N_38323,N_36789,N_35080);
and U38324 (N_38324,N_36714,N_37246);
or U38325 (N_38325,N_36264,N_36395);
or U38326 (N_38326,N_36933,N_36166);
xnor U38327 (N_38327,N_36530,N_36561);
or U38328 (N_38328,N_35869,N_35040);
nand U38329 (N_38329,N_36355,N_37138);
or U38330 (N_38330,N_36756,N_35607);
nand U38331 (N_38331,N_37227,N_35777);
and U38332 (N_38332,N_35625,N_35106);
and U38333 (N_38333,N_37096,N_35877);
xnor U38334 (N_38334,N_35331,N_36717);
or U38335 (N_38335,N_35781,N_35436);
or U38336 (N_38336,N_36133,N_35058);
nand U38337 (N_38337,N_37102,N_36495);
nand U38338 (N_38338,N_36293,N_36534);
or U38339 (N_38339,N_36546,N_37493);
and U38340 (N_38340,N_36853,N_36514);
and U38341 (N_38341,N_35473,N_35189);
or U38342 (N_38342,N_36013,N_36002);
xor U38343 (N_38343,N_37379,N_35065);
or U38344 (N_38344,N_35576,N_35006);
and U38345 (N_38345,N_36345,N_37302);
xor U38346 (N_38346,N_36955,N_36384);
and U38347 (N_38347,N_35572,N_35230);
nand U38348 (N_38348,N_37428,N_36779);
xnor U38349 (N_38349,N_36198,N_36649);
or U38350 (N_38350,N_35747,N_35970);
nor U38351 (N_38351,N_35971,N_36171);
and U38352 (N_38352,N_35998,N_37465);
or U38353 (N_38353,N_36043,N_35846);
or U38354 (N_38354,N_35794,N_35512);
nor U38355 (N_38355,N_37392,N_37468);
nor U38356 (N_38356,N_36747,N_37093);
xnor U38357 (N_38357,N_37423,N_35681);
or U38358 (N_38358,N_35853,N_36783);
nor U38359 (N_38359,N_37451,N_37289);
nand U38360 (N_38360,N_35516,N_35029);
nand U38361 (N_38361,N_36169,N_36710);
or U38362 (N_38362,N_35097,N_35336);
xnor U38363 (N_38363,N_36037,N_35422);
and U38364 (N_38364,N_35146,N_37099);
and U38365 (N_38365,N_35862,N_36676);
or U38366 (N_38366,N_36965,N_36488);
or U38367 (N_38367,N_35271,N_35772);
nor U38368 (N_38368,N_36551,N_35875);
or U38369 (N_38369,N_36113,N_37387);
xor U38370 (N_38370,N_35975,N_36213);
and U38371 (N_38371,N_35398,N_35786);
nand U38372 (N_38372,N_36024,N_36909);
nor U38373 (N_38373,N_36629,N_35802);
nand U38374 (N_38374,N_37078,N_35928);
and U38375 (N_38375,N_36518,N_36211);
xor U38376 (N_38376,N_35993,N_37369);
xor U38377 (N_38377,N_37234,N_37013);
nand U38378 (N_38378,N_36400,N_37485);
nor U38379 (N_38379,N_37341,N_35931);
xnor U38380 (N_38380,N_37407,N_35879);
nand U38381 (N_38381,N_36970,N_37018);
nand U38382 (N_38382,N_35691,N_37480);
and U38383 (N_38383,N_37228,N_35814);
and U38384 (N_38384,N_36438,N_35094);
nor U38385 (N_38385,N_37061,N_35538);
nand U38386 (N_38386,N_36402,N_35821);
and U38387 (N_38387,N_35988,N_36263);
nor U38388 (N_38388,N_37461,N_36624);
nand U38389 (N_38389,N_35631,N_35700);
and U38390 (N_38390,N_35540,N_37029);
or U38391 (N_38391,N_35776,N_35367);
and U38392 (N_38392,N_35686,N_35688);
or U38393 (N_38393,N_35225,N_35726);
and U38394 (N_38394,N_36609,N_36281);
nand U38395 (N_38395,N_36164,N_37174);
and U38396 (N_38396,N_35739,N_36122);
and U38397 (N_38397,N_35878,N_35857);
nand U38398 (N_38398,N_35725,N_36625);
and U38399 (N_38399,N_35969,N_35042);
xnor U38400 (N_38400,N_36238,N_37463);
nand U38401 (N_38401,N_35021,N_37112);
and U38402 (N_38402,N_35110,N_35485);
or U38403 (N_38403,N_36388,N_37235);
xor U38404 (N_38404,N_35630,N_35703);
or U38405 (N_38405,N_35497,N_35547);
nor U38406 (N_38406,N_35408,N_35748);
and U38407 (N_38407,N_37312,N_36920);
xnor U38408 (N_38408,N_35889,N_35196);
nand U38409 (N_38409,N_36155,N_35108);
and U38410 (N_38410,N_36012,N_37036);
nor U38411 (N_38411,N_37449,N_35319);
nor U38412 (N_38412,N_35509,N_36161);
xor U38413 (N_38413,N_36929,N_35500);
nand U38414 (N_38414,N_37266,N_37453);
and U38415 (N_38415,N_36907,N_37358);
nand U38416 (N_38416,N_35961,N_35460);
nor U38417 (N_38417,N_36851,N_37330);
and U38418 (N_38418,N_35204,N_36560);
and U38419 (N_38419,N_35488,N_36924);
and U38420 (N_38420,N_37257,N_37079);
nor U38421 (N_38421,N_35483,N_36524);
nor U38422 (N_38422,N_36128,N_36713);
nand U38423 (N_38423,N_36435,N_36796);
and U38424 (N_38424,N_36532,N_36978);
nor U38425 (N_38425,N_36476,N_35902);
or U38426 (N_38426,N_35152,N_35182);
or U38427 (N_38427,N_36515,N_35487);
nand U38428 (N_38428,N_36782,N_36126);
nor U38429 (N_38429,N_35999,N_35701);
xnor U38430 (N_38430,N_35529,N_36074);
xnor U38431 (N_38431,N_35423,N_36456);
nor U38432 (N_38432,N_36243,N_35804);
and U38433 (N_38433,N_36681,N_35508);
and U38434 (N_38434,N_35135,N_35075);
nand U38435 (N_38435,N_37216,N_36507);
or U38436 (N_38436,N_35785,N_36149);
nor U38437 (N_38437,N_37303,N_35608);
and U38438 (N_38438,N_37251,N_37306);
nand U38439 (N_38439,N_37173,N_35938);
and U38440 (N_38440,N_36050,N_36365);
nor U38441 (N_38441,N_35287,N_37217);
or U38442 (N_38442,N_37005,N_35822);
nor U38443 (N_38443,N_35657,N_35125);
or U38444 (N_38444,N_36590,N_35092);
nor U38445 (N_38445,N_35571,N_37382);
and U38446 (N_38446,N_36496,N_36425);
and U38447 (N_38447,N_35940,N_36583);
and U38448 (N_38448,N_37427,N_37117);
nor U38449 (N_38449,N_35440,N_36608);
nand U38450 (N_38450,N_35733,N_36132);
or U38451 (N_38451,N_35397,N_35054);
nand U38452 (N_38452,N_37490,N_36784);
xnor U38453 (N_38453,N_36194,N_36639);
and U38454 (N_38454,N_35907,N_37386);
xnor U38455 (N_38455,N_35983,N_35627);
nand U38456 (N_38456,N_37152,N_36449);
nor U38457 (N_38457,N_35568,N_36686);
or U38458 (N_38458,N_35557,N_36254);
or U38459 (N_38459,N_36267,N_37495);
and U38460 (N_38460,N_35521,N_35735);
or U38461 (N_38461,N_37201,N_35585);
and U38462 (N_38462,N_37297,N_36452);
and U38463 (N_38463,N_36000,N_37426);
and U38464 (N_38464,N_36567,N_36337);
or U38465 (N_38465,N_36528,N_37391);
and U38466 (N_38466,N_36309,N_36539);
or U38467 (N_38467,N_35574,N_37204);
nand U38468 (N_38468,N_36834,N_35880);
nor U38469 (N_38469,N_35751,N_35605);
nor U38470 (N_38470,N_35829,N_36971);
nor U38471 (N_38471,N_36217,N_36109);
nand U38472 (N_38472,N_36300,N_35502);
and U38473 (N_38473,N_36523,N_35355);
nand U38474 (N_38474,N_35456,N_35380);
xnor U38475 (N_38475,N_36642,N_35298);
and U38476 (N_38476,N_35622,N_35078);
and U38477 (N_38477,N_35102,N_36775);
nor U38478 (N_38478,N_36809,N_36910);
or U38479 (N_38479,N_36310,N_36494);
nor U38480 (N_38480,N_36255,N_37402);
and U38481 (N_38481,N_35687,N_36478);
and U38482 (N_38482,N_36882,N_35166);
and U38483 (N_38483,N_37315,N_36860);
xnor U38484 (N_38484,N_35533,N_36301);
or U38485 (N_38485,N_35935,N_35280);
or U38486 (N_38486,N_36443,N_36305);
nand U38487 (N_38487,N_36371,N_35056);
and U38488 (N_38488,N_37232,N_36636);
and U38489 (N_38489,N_37136,N_35963);
and U38490 (N_38490,N_36200,N_35333);
nand U38491 (N_38491,N_36486,N_36054);
xnor U38492 (N_38492,N_35874,N_36688);
nor U38493 (N_38493,N_36506,N_35268);
and U38494 (N_38494,N_35528,N_35162);
nand U38495 (N_38495,N_37393,N_36573);
nand U38496 (N_38496,N_37196,N_36039);
and U38497 (N_38497,N_36290,N_36056);
or U38498 (N_38498,N_36966,N_36244);
nor U38499 (N_38499,N_36857,N_36308);
nor U38500 (N_38500,N_36827,N_36763);
and U38501 (N_38501,N_35361,N_35143);
xnor U38502 (N_38502,N_35826,N_37073);
nor U38503 (N_38503,N_35569,N_35513);
nand U38504 (N_38504,N_37448,N_37344);
xnor U38505 (N_38505,N_37482,N_35504);
and U38506 (N_38506,N_35348,N_35053);
and U38507 (N_38507,N_36839,N_35599);
nand U38508 (N_38508,N_36066,N_35183);
nor U38509 (N_38509,N_36800,N_36986);
nor U38510 (N_38510,N_35438,N_35463);
xor U38511 (N_38511,N_35201,N_35086);
and U38512 (N_38512,N_36116,N_36735);
or U38513 (N_38513,N_35076,N_36040);
and U38514 (N_38514,N_35779,N_35536);
and U38515 (N_38515,N_36086,N_35946);
or U38516 (N_38516,N_35883,N_35410);
or U38517 (N_38517,N_36431,N_35668);
or U38518 (N_38518,N_36559,N_36888);
nand U38519 (N_38519,N_37308,N_36468);
and U38520 (N_38520,N_36976,N_35437);
or U38521 (N_38521,N_37058,N_36143);
and U38522 (N_38522,N_35888,N_35773);
nor U38523 (N_38523,N_36333,N_35105);
and U38524 (N_38524,N_36261,N_37415);
nand U38525 (N_38525,N_37255,N_35083);
or U38526 (N_38526,N_35966,N_35279);
nand U38527 (N_38527,N_37271,N_36185);
nand U38528 (N_38528,N_37474,N_37066);
nand U38529 (N_38529,N_35426,N_36956);
nor U38530 (N_38530,N_37374,N_36511);
nand U38531 (N_38531,N_35167,N_35023);
and U38532 (N_38532,N_35141,N_36548);
nand U38533 (N_38533,N_35357,N_37313);
nand U38534 (N_38534,N_35134,N_35662);
nand U38535 (N_38535,N_36042,N_36442);
nand U38536 (N_38536,N_36052,N_37430);
nor U38537 (N_38537,N_37021,N_36612);
or U38538 (N_38538,N_36679,N_35091);
xor U38539 (N_38539,N_35915,N_37247);
nor U38540 (N_38540,N_36022,N_37440);
or U38541 (N_38541,N_35022,N_35980);
and U38542 (N_38542,N_35699,N_35964);
and U38543 (N_38543,N_36191,N_35957);
nor U38544 (N_38544,N_36212,N_35731);
and U38545 (N_38545,N_35835,N_35997);
xnor U38546 (N_38546,N_36288,N_37107);
nand U38547 (N_38547,N_35373,N_35598);
nor U38548 (N_38548,N_35122,N_37293);
and U38549 (N_38549,N_37192,N_35753);
or U38550 (N_38550,N_35640,N_35898);
nand U38551 (N_38551,N_35366,N_37483);
nand U38552 (N_38552,N_37015,N_36262);
nand U38553 (N_38553,N_36218,N_36906);
nor U38554 (N_38554,N_35400,N_37394);
xor U38555 (N_38555,N_35832,N_37283);
nor U38556 (N_38556,N_35799,N_35341);
and U38557 (N_38557,N_36011,N_35406);
nor U38558 (N_38558,N_37169,N_37119);
xor U38559 (N_38559,N_36758,N_36490);
nand U38560 (N_38560,N_37151,N_36542);
and U38561 (N_38561,N_36319,N_36173);
nand U38562 (N_38562,N_36472,N_37057);
or U38563 (N_38563,N_36209,N_35895);
and U38564 (N_38564,N_37337,N_35580);
nor U38565 (N_38565,N_35526,N_35070);
and U38566 (N_38566,N_35491,N_35624);
or U38567 (N_38567,N_36814,N_35149);
nand U38568 (N_38568,N_36206,N_35206);
nand U38569 (N_38569,N_37420,N_36136);
nand U38570 (N_38570,N_35644,N_35346);
nand U38571 (N_38571,N_35343,N_35153);
or U38572 (N_38572,N_35223,N_36481);
nor U38573 (N_38573,N_36058,N_36458);
nand U38574 (N_38574,N_35064,N_35044);
nor U38575 (N_38575,N_37110,N_35728);
nand U38576 (N_38576,N_37357,N_36939);
or U38577 (N_38577,N_37052,N_36741);
or U38578 (N_38578,N_35347,N_36930);
and U38579 (N_38579,N_35642,N_36598);
nand U38580 (N_38580,N_35325,N_36298);
nand U38581 (N_38581,N_36999,N_37077);
nor U38582 (N_38582,N_36075,N_36550);
nor U38583 (N_38583,N_36036,N_36248);
or U38584 (N_38584,N_36134,N_36820);
and U38585 (N_38585,N_35759,N_36245);
nand U38586 (N_38586,N_36777,N_35411);
and U38587 (N_38587,N_36536,N_36669);
nand U38588 (N_38588,N_35358,N_35299);
xnor U38589 (N_38589,N_35263,N_35519);
nor U38590 (N_38590,N_36232,N_37002);
nand U38591 (N_38591,N_37378,N_35339);
or U38592 (N_38592,N_36902,N_35184);
nor U38593 (N_38593,N_36865,N_35721);
and U38594 (N_38594,N_36287,N_36082);
nand U38595 (N_38595,N_36440,N_36894);
nand U38596 (N_38596,N_36063,N_35009);
nor U38597 (N_38597,N_37384,N_36891);
and U38598 (N_38598,N_35447,N_35160);
or U38599 (N_38599,N_36152,N_35302);
nand U38600 (N_38600,N_35034,N_35455);
or U38601 (N_38601,N_37254,N_35390);
nor U38602 (N_38602,N_35481,N_35943);
and U38603 (N_38603,N_36653,N_36372);
nand U38604 (N_38604,N_36849,N_35474);
nand U38605 (N_38605,N_36722,N_36424);
and U38606 (N_38606,N_35265,N_35352);
nor U38607 (N_38607,N_36960,N_37260);
nor U38608 (N_38608,N_36549,N_37488);
nand U38609 (N_38609,N_36256,N_36917);
and U38610 (N_38610,N_37055,N_35724);
or U38611 (N_38611,N_36619,N_36105);
nand U38612 (N_38612,N_35965,N_35365);
and U38613 (N_38613,N_37125,N_36204);
or U38614 (N_38614,N_35676,N_35131);
and U38615 (N_38615,N_37275,N_36028);
and U38616 (N_38616,N_35518,N_36276);
nand U38617 (N_38617,N_37370,N_35014);
nor U38618 (N_38618,N_36797,N_37491);
or U38619 (N_38619,N_35899,N_36887);
nand U38620 (N_38620,N_35944,N_35462);
nand U38621 (N_38621,N_35780,N_35377);
xnor U38622 (N_38622,N_35514,N_37486);
xor U38623 (N_38623,N_36772,N_36127);
and U38624 (N_38624,N_36280,N_37132);
or U38625 (N_38625,N_36473,N_37309);
nor U38626 (N_38626,N_35932,N_36092);
and U38627 (N_38627,N_35128,N_37199);
nor U38628 (N_38628,N_35674,N_35882);
or U38629 (N_38629,N_37460,N_35433);
nand U38630 (N_38630,N_35800,N_36142);
xor U38631 (N_38631,N_37285,N_36283);
and U38632 (N_38632,N_35340,N_36631);
xnor U38633 (N_38633,N_36270,N_35658);
or U38634 (N_38634,N_36224,N_36744);
xnor U38635 (N_38635,N_35936,N_35744);
nand U38636 (N_38636,N_35926,N_35224);
nor U38637 (N_38637,N_36593,N_37300);
nor U38638 (N_38638,N_37082,N_36041);
and U38639 (N_38639,N_36318,N_36304);
and U38640 (N_38640,N_35809,N_36382);
or U38641 (N_38641,N_35851,N_35652);
nor U38642 (N_38642,N_35061,N_36018);
nor U38643 (N_38643,N_36541,N_36977);
nand U38644 (N_38644,N_37236,N_35494);
and U38645 (N_38645,N_36872,N_36067);
and U38646 (N_38646,N_35885,N_35541);
nand U38647 (N_38647,N_35665,N_36273);
nand U38648 (N_38648,N_36805,N_36628);
nand U38649 (N_38649,N_37328,N_37229);
nor U38650 (N_38650,N_35186,N_35163);
nor U38651 (N_38651,N_35079,N_36035);
or U38652 (N_38652,N_36660,N_36396);
nand U38653 (N_38653,N_36059,N_36409);
and U38654 (N_38654,N_37425,N_35767);
nand U38655 (N_38655,N_36376,N_35861);
xor U38656 (N_38656,N_36096,N_36179);
nand U38657 (N_38657,N_36675,N_36373);
or U38658 (N_38658,N_36077,N_36334);
nand U38659 (N_38659,N_36237,N_36729);
xnor U38660 (N_38660,N_35305,N_35636);
nand U38661 (N_38661,N_35301,N_35996);
nand U38662 (N_38662,N_36021,N_35387);
or U38663 (N_38663,N_37409,N_36027);
nor U38664 (N_38664,N_36348,N_36535);
and U38665 (N_38665,N_35249,N_35114);
nor U38666 (N_38666,N_36361,N_35321);
and U38667 (N_38667,N_37317,N_36531);
or U38668 (N_38668,N_36332,N_36112);
nand U38669 (N_38669,N_36526,N_35425);
xnor U38670 (N_38670,N_37085,N_35129);
nand U38671 (N_38671,N_35867,N_36812);
xnor U38672 (N_38672,N_35480,N_36393);
nor U38673 (N_38673,N_36030,N_37245);
nand U38674 (N_38674,N_35156,N_37046);
or U38675 (N_38675,N_37277,N_36757);
or U38676 (N_38676,N_35754,N_35650);
and U38677 (N_38677,N_35235,N_35222);
nand U38678 (N_38678,N_35432,N_35033);
or U38679 (N_38679,N_36417,N_35950);
and U38680 (N_38680,N_35849,N_35032);
and U38681 (N_38681,N_35695,N_36916);
nor U38682 (N_38682,N_36257,N_36460);
nor U38683 (N_38683,N_35490,N_37081);
and U38684 (N_38684,N_37412,N_36339);
and U38685 (N_38685,N_36350,N_35982);
or U38686 (N_38686,N_35269,N_37087);
nor U38687 (N_38687,N_35171,N_36048);
nand U38688 (N_38688,N_36500,N_35838);
xnor U38689 (N_38689,N_37324,N_35916);
and U38690 (N_38690,N_35272,N_35240);
or U38691 (N_38691,N_37325,N_35558);
nor U38692 (N_38692,N_37360,N_35288);
nor U38693 (N_38693,N_37042,N_37014);
and U38694 (N_38694,N_36325,N_36943);
nor U38695 (N_38695,N_35937,N_35900);
nand U38696 (N_38696,N_36607,N_35597);
nor U38697 (N_38697,N_36111,N_36605);
and U38698 (N_38698,N_37178,N_36566);
and U38699 (N_38699,N_35399,N_35798);
or U38700 (N_38700,N_36017,N_35706);
nor U38701 (N_38701,N_37086,N_35909);
xnor U38702 (N_38702,N_35266,N_37356);
nor U38703 (N_38703,N_36641,N_35254);
or U38704 (N_38704,N_36819,N_36184);
or U38705 (N_38705,N_35354,N_36306);
nor U38706 (N_38706,N_36006,N_37272);
or U38707 (N_38707,N_36786,N_36505);
nand U38708 (N_38708,N_36731,N_37320);
or U38709 (N_38709,N_37367,N_37121);
and U38710 (N_38710,N_35100,N_35917);
nor U38711 (N_38711,N_35873,N_36761);
or U38712 (N_38712,N_36708,N_37022);
or U38713 (N_38713,N_36881,N_36662);
or U38714 (N_38714,N_36932,N_36787);
nand U38715 (N_38715,N_36580,N_35089);
xnor U38716 (N_38716,N_35242,N_36180);
nand U38717 (N_38717,N_35123,N_36859);
xor U38718 (N_38718,N_35890,N_35962);
nor U38719 (N_38719,N_36148,N_37316);
and U38720 (N_38720,N_35710,N_36895);
and U38721 (N_38721,N_35060,N_36352);
nand U38722 (N_38722,N_35099,N_36314);
nor U38723 (N_38723,N_36260,N_37499);
or U38724 (N_38724,N_37381,N_35311);
or U38725 (N_38725,N_36034,N_36165);
nand U38726 (N_38726,N_36983,N_36883);
nand U38727 (N_38727,N_36235,N_35764);
nand U38728 (N_38728,N_36890,N_37065);
and U38729 (N_38729,N_37165,N_36150);
nand U38730 (N_38730,N_36575,N_35351);
or U38731 (N_38731,N_37001,N_37063);
xnor U38732 (N_38732,N_37203,N_36997);
xor U38733 (N_38733,N_37492,N_36015);
or U38734 (N_38734,N_35394,N_36900);
and U38735 (N_38735,N_36032,N_36266);
or U38736 (N_38736,N_36158,N_35545);
xor U38737 (N_38737,N_35884,N_36208);
xor U38738 (N_38738,N_36592,N_37120);
nor U38739 (N_38739,N_36963,N_35031);
and U38740 (N_38740,N_36228,N_36837);
nand U38741 (N_38741,N_37091,N_35820);
and U38742 (N_38742,N_35690,N_36954);
or U38743 (N_38743,N_36770,N_36282);
or U38744 (N_38744,N_36186,N_36110);
and U38745 (N_38745,N_37417,N_36129);
xnor U38746 (N_38746,N_36205,N_36064);
or U38747 (N_38747,N_36379,N_35522);
nor U38748 (N_38748,N_37044,N_36855);
or U38749 (N_38749,N_35708,N_37291);
and U38750 (N_38750,N_37331,N_37490);
nor U38751 (N_38751,N_36677,N_35391);
or U38752 (N_38752,N_36008,N_37470);
nor U38753 (N_38753,N_35539,N_37181);
and U38754 (N_38754,N_36856,N_36592);
and U38755 (N_38755,N_37270,N_36707);
nor U38756 (N_38756,N_36317,N_35951);
and U38757 (N_38757,N_35421,N_36558);
nand U38758 (N_38758,N_37056,N_36571);
nand U38759 (N_38759,N_35510,N_36618);
nor U38760 (N_38760,N_37013,N_35153);
nand U38761 (N_38761,N_35673,N_37303);
xnor U38762 (N_38762,N_37211,N_35507);
nor U38763 (N_38763,N_36969,N_36121);
nand U38764 (N_38764,N_35527,N_35426);
nor U38765 (N_38765,N_37157,N_35874);
nand U38766 (N_38766,N_36842,N_36919);
nor U38767 (N_38767,N_35030,N_35255);
xnor U38768 (N_38768,N_36177,N_36139);
nor U38769 (N_38769,N_35827,N_37082);
nand U38770 (N_38770,N_36958,N_35079);
nand U38771 (N_38771,N_35878,N_37004);
or U38772 (N_38772,N_37075,N_36092);
xnor U38773 (N_38773,N_36217,N_35706);
nor U38774 (N_38774,N_37365,N_36571);
and U38775 (N_38775,N_35225,N_37472);
nor U38776 (N_38776,N_35108,N_36975);
and U38777 (N_38777,N_36167,N_37305);
and U38778 (N_38778,N_36832,N_35738);
nand U38779 (N_38779,N_36185,N_36816);
nand U38780 (N_38780,N_36007,N_36263);
or U38781 (N_38781,N_36804,N_35262);
and U38782 (N_38782,N_35827,N_35244);
nor U38783 (N_38783,N_35708,N_36645);
nor U38784 (N_38784,N_36889,N_35219);
nor U38785 (N_38785,N_36265,N_35286);
nor U38786 (N_38786,N_35332,N_36131);
nand U38787 (N_38787,N_37304,N_35365);
nand U38788 (N_38788,N_35724,N_36924);
and U38789 (N_38789,N_35222,N_35588);
nand U38790 (N_38790,N_36503,N_36293);
nand U38791 (N_38791,N_36181,N_37441);
or U38792 (N_38792,N_35467,N_36831);
or U38793 (N_38793,N_36333,N_36942);
or U38794 (N_38794,N_37061,N_37348);
nor U38795 (N_38795,N_36234,N_36161);
xnor U38796 (N_38796,N_35650,N_35549);
xor U38797 (N_38797,N_36320,N_36398);
and U38798 (N_38798,N_36473,N_36751);
and U38799 (N_38799,N_36718,N_35389);
nand U38800 (N_38800,N_35597,N_36235);
nand U38801 (N_38801,N_36052,N_36543);
xor U38802 (N_38802,N_35259,N_36648);
nor U38803 (N_38803,N_35070,N_35187);
nand U38804 (N_38804,N_36646,N_35166);
nand U38805 (N_38805,N_36287,N_35014);
and U38806 (N_38806,N_36692,N_35446);
xor U38807 (N_38807,N_35598,N_35397);
and U38808 (N_38808,N_37264,N_36911);
xnor U38809 (N_38809,N_35320,N_37176);
nor U38810 (N_38810,N_37364,N_35977);
nand U38811 (N_38811,N_37242,N_36309);
or U38812 (N_38812,N_37136,N_36180);
and U38813 (N_38813,N_37444,N_36969);
nor U38814 (N_38814,N_36669,N_36803);
and U38815 (N_38815,N_36834,N_37444);
or U38816 (N_38816,N_35519,N_35000);
or U38817 (N_38817,N_36248,N_35299);
or U38818 (N_38818,N_36285,N_35941);
nand U38819 (N_38819,N_35547,N_35802);
nor U38820 (N_38820,N_36952,N_35711);
nor U38821 (N_38821,N_36865,N_36221);
and U38822 (N_38822,N_36691,N_35433);
and U38823 (N_38823,N_36776,N_35310);
xor U38824 (N_38824,N_35485,N_37462);
or U38825 (N_38825,N_35515,N_35840);
and U38826 (N_38826,N_35543,N_35116);
nor U38827 (N_38827,N_36420,N_35024);
and U38828 (N_38828,N_37049,N_37308);
nor U38829 (N_38829,N_35520,N_35805);
nand U38830 (N_38830,N_36559,N_36015);
nand U38831 (N_38831,N_36658,N_36066);
nand U38832 (N_38832,N_37142,N_36813);
and U38833 (N_38833,N_35886,N_36442);
or U38834 (N_38834,N_37173,N_35178);
or U38835 (N_38835,N_36128,N_35906);
nor U38836 (N_38836,N_36120,N_35747);
or U38837 (N_38837,N_36565,N_37368);
nand U38838 (N_38838,N_37141,N_36833);
nand U38839 (N_38839,N_37437,N_36884);
and U38840 (N_38840,N_36296,N_36942);
and U38841 (N_38841,N_35991,N_35095);
nor U38842 (N_38842,N_36801,N_37409);
nand U38843 (N_38843,N_35822,N_35168);
nand U38844 (N_38844,N_36837,N_36634);
or U38845 (N_38845,N_37193,N_35076);
and U38846 (N_38846,N_36107,N_36791);
and U38847 (N_38847,N_36821,N_35299);
or U38848 (N_38848,N_37058,N_35180);
and U38849 (N_38849,N_36800,N_35829);
nor U38850 (N_38850,N_36170,N_35912);
nor U38851 (N_38851,N_35638,N_35263);
or U38852 (N_38852,N_37123,N_35603);
and U38853 (N_38853,N_36051,N_36577);
nor U38854 (N_38854,N_36535,N_35381);
nand U38855 (N_38855,N_36625,N_35695);
nand U38856 (N_38856,N_36579,N_36232);
or U38857 (N_38857,N_35562,N_36545);
xor U38858 (N_38858,N_37491,N_36701);
or U38859 (N_38859,N_37099,N_35984);
xnor U38860 (N_38860,N_35457,N_36345);
and U38861 (N_38861,N_36502,N_35804);
or U38862 (N_38862,N_35112,N_37310);
xor U38863 (N_38863,N_37465,N_37262);
nand U38864 (N_38864,N_36806,N_35362);
or U38865 (N_38865,N_36241,N_35553);
or U38866 (N_38866,N_37184,N_36497);
or U38867 (N_38867,N_35588,N_35420);
nor U38868 (N_38868,N_35582,N_35221);
or U38869 (N_38869,N_35137,N_35335);
and U38870 (N_38870,N_35669,N_35115);
and U38871 (N_38871,N_35690,N_36442);
or U38872 (N_38872,N_36837,N_35349);
nor U38873 (N_38873,N_36535,N_37338);
xor U38874 (N_38874,N_35225,N_36675);
or U38875 (N_38875,N_35499,N_35470);
and U38876 (N_38876,N_37414,N_36942);
nor U38877 (N_38877,N_35925,N_37204);
nand U38878 (N_38878,N_36433,N_35256);
and U38879 (N_38879,N_35959,N_35789);
nand U38880 (N_38880,N_37222,N_36008);
nand U38881 (N_38881,N_37344,N_37106);
nor U38882 (N_38882,N_35502,N_36175);
nand U38883 (N_38883,N_35227,N_36143);
nand U38884 (N_38884,N_35718,N_35528);
nor U38885 (N_38885,N_35813,N_36366);
nand U38886 (N_38886,N_36461,N_36852);
and U38887 (N_38887,N_35198,N_36714);
or U38888 (N_38888,N_35342,N_37272);
xor U38889 (N_38889,N_35027,N_36084);
nor U38890 (N_38890,N_35954,N_35805);
and U38891 (N_38891,N_36157,N_37351);
nand U38892 (N_38892,N_35826,N_36898);
nor U38893 (N_38893,N_36833,N_35531);
and U38894 (N_38894,N_35676,N_35357);
and U38895 (N_38895,N_35762,N_37079);
and U38896 (N_38896,N_36446,N_35712);
or U38897 (N_38897,N_35649,N_36350);
nand U38898 (N_38898,N_36587,N_37139);
and U38899 (N_38899,N_37034,N_36151);
nand U38900 (N_38900,N_37196,N_36571);
nor U38901 (N_38901,N_36842,N_35228);
nand U38902 (N_38902,N_37170,N_36614);
or U38903 (N_38903,N_35834,N_36489);
nor U38904 (N_38904,N_35189,N_35011);
or U38905 (N_38905,N_36191,N_35047);
or U38906 (N_38906,N_36261,N_35567);
or U38907 (N_38907,N_36085,N_36745);
nor U38908 (N_38908,N_36250,N_37219);
nand U38909 (N_38909,N_37368,N_35396);
nor U38910 (N_38910,N_36601,N_35230);
or U38911 (N_38911,N_36753,N_35369);
nor U38912 (N_38912,N_35360,N_37434);
or U38913 (N_38913,N_37083,N_35478);
and U38914 (N_38914,N_35923,N_37053);
nor U38915 (N_38915,N_36053,N_36769);
and U38916 (N_38916,N_37016,N_35222);
and U38917 (N_38917,N_35023,N_36006);
nand U38918 (N_38918,N_35934,N_37363);
and U38919 (N_38919,N_35363,N_37436);
or U38920 (N_38920,N_37220,N_37063);
nor U38921 (N_38921,N_35135,N_36167);
and U38922 (N_38922,N_35865,N_35984);
and U38923 (N_38923,N_36046,N_36076);
xnor U38924 (N_38924,N_35364,N_37431);
nor U38925 (N_38925,N_35554,N_36250);
nor U38926 (N_38926,N_37059,N_36858);
or U38927 (N_38927,N_36579,N_36623);
and U38928 (N_38928,N_37239,N_36541);
xnor U38929 (N_38929,N_35079,N_35868);
nand U38930 (N_38930,N_35999,N_36393);
or U38931 (N_38931,N_35405,N_35827);
nor U38932 (N_38932,N_36706,N_35157);
nor U38933 (N_38933,N_35333,N_36457);
xnor U38934 (N_38934,N_36828,N_35153);
or U38935 (N_38935,N_35094,N_36341);
nor U38936 (N_38936,N_36627,N_35123);
nand U38937 (N_38937,N_36724,N_37423);
or U38938 (N_38938,N_37360,N_36871);
nand U38939 (N_38939,N_35009,N_35731);
or U38940 (N_38940,N_35898,N_37355);
xnor U38941 (N_38941,N_36468,N_36941);
nand U38942 (N_38942,N_35837,N_36419);
xnor U38943 (N_38943,N_37182,N_37054);
and U38944 (N_38944,N_37175,N_36494);
nor U38945 (N_38945,N_36642,N_36897);
nand U38946 (N_38946,N_36427,N_36703);
or U38947 (N_38947,N_36607,N_36037);
and U38948 (N_38948,N_36929,N_35270);
nand U38949 (N_38949,N_36831,N_36623);
xnor U38950 (N_38950,N_37385,N_35436);
and U38951 (N_38951,N_36701,N_36003);
and U38952 (N_38952,N_37407,N_36608);
and U38953 (N_38953,N_35484,N_36907);
and U38954 (N_38954,N_36875,N_35770);
xor U38955 (N_38955,N_37474,N_36935);
or U38956 (N_38956,N_35169,N_36454);
and U38957 (N_38957,N_36849,N_37464);
xnor U38958 (N_38958,N_36894,N_35076);
nor U38959 (N_38959,N_36669,N_36998);
or U38960 (N_38960,N_35166,N_35471);
xor U38961 (N_38961,N_37447,N_37135);
or U38962 (N_38962,N_35013,N_37375);
nand U38963 (N_38963,N_36023,N_36770);
or U38964 (N_38964,N_35292,N_36738);
and U38965 (N_38965,N_36058,N_35355);
or U38966 (N_38966,N_35961,N_36780);
nand U38967 (N_38967,N_35181,N_37205);
or U38968 (N_38968,N_36682,N_36984);
or U38969 (N_38969,N_37295,N_36909);
and U38970 (N_38970,N_36648,N_35174);
or U38971 (N_38971,N_35128,N_35822);
nor U38972 (N_38972,N_35560,N_35955);
or U38973 (N_38973,N_36295,N_36531);
nor U38974 (N_38974,N_35921,N_35701);
nor U38975 (N_38975,N_37162,N_35858);
or U38976 (N_38976,N_36912,N_35646);
nor U38977 (N_38977,N_35148,N_35330);
nand U38978 (N_38978,N_36064,N_35212);
and U38979 (N_38979,N_35080,N_37046);
nand U38980 (N_38980,N_35767,N_36450);
nand U38981 (N_38981,N_36764,N_36501);
or U38982 (N_38982,N_36834,N_35562);
xor U38983 (N_38983,N_36729,N_35594);
or U38984 (N_38984,N_36186,N_35680);
or U38985 (N_38985,N_37057,N_35544);
and U38986 (N_38986,N_36661,N_36726);
or U38987 (N_38987,N_35733,N_35911);
and U38988 (N_38988,N_35592,N_36563);
or U38989 (N_38989,N_36635,N_36163);
or U38990 (N_38990,N_35742,N_36207);
or U38991 (N_38991,N_36295,N_37133);
or U38992 (N_38992,N_36508,N_35865);
or U38993 (N_38993,N_35962,N_35518);
and U38994 (N_38994,N_37037,N_37301);
and U38995 (N_38995,N_35060,N_37344);
or U38996 (N_38996,N_36418,N_35759);
nand U38997 (N_38997,N_36188,N_35592);
nor U38998 (N_38998,N_36111,N_35331);
nand U38999 (N_38999,N_36465,N_36078);
nor U39000 (N_39000,N_35121,N_36287);
nand U39001 (N_39001,N_36786,N_36001);
nand U39002 (N_39002,N_36186,N_36596);
xor U39003 (N_39003,N_35226,N_35143);
and U39004 (N_39004,N_35962,N_36982);
nand U39005 (N_39005,N_36145,N_35379);
nand U39006 (N_39006,N_37107,N_36198);
and U39007 (N_39007,N_37272,N_36698);
or U39008 (N_39008,N_36735,N_36995);
or U39009 (N_39009,N_36859,N_35517);
nand U39010 (N_39010,N_35920,N_35014);
and U39011 (N_39011,N_35805,N_37319);
xor U39012 (N_39012,N_35795,N_35327);
xor U39013 (N_39013,N_37366,N_36026);
and U39014 (N_39014,N_36398,N_37179);
and U39015 (N_39015,N_37184,N_36360);
or U39016 (N_39016,N_35109,N_35723);
nand U39017 (N_39017,N_35423,N_37466);
nor U39018 (N_39018,N_37229,N_37147);
and U39019 (N_39019,N_36143,N_35725);
and U39020 (N_39020,N_35864,N_36662);
nand U39021 (N_39021,N_35055,N_36314);
xnor U39022 (N_39022,N_35166,N_36085);
and U39023 (N_39023,N_35338,N_36930);
nand U39024 (N_39024,N_35255,N_35822);
and U39025 (N_39025,N_37493,N_36481);
nand U39026 (N_39026,N_37438,N_36980);
nor U39027 (N_39027,N_36550,N_36296);
nand U39028 (N_39028,N_37084,N_36317);
nand U39029 (N_39029,N_35213,N_36498);
and U39030 (N_39030,N_35908,N_35914);
xnor U39031 (N_39031,N_36232,N_36781);
and U39032 (N_39032,N_35783,N_37448);
nand U39033 (N_39033,N_35372,N_36521);
xor U39034 (N_39034,N_36437,N_36654);
xnor U39035 (N_39035,N_37411,N_37259);
or U39036 (N_39036,N_35727,N_36005);
or U39037 (N_39037,N_35072,N_37309);
nand U39038 (N_39038,N_37018,N_35758);
nand U39039 (N_39039,N_35801,N_36355);
or U39040 (N_39040,N_35681,N_35318);
xnor U39041 (N_39041,N_35953,N_36026);
nand U39042 (N_39042,N_36698,N_36404);
or U39043 (N_39043,N_36788,N_37467);
nor U39044 (N_39044,N_35115,N_36795);
or U39045 (N_39045,N_36180,N_35388);
and U39046 (N_39046,N_36394,N_35552);
and U39047 (N_39047,N_37495,N_36684);
nand U39048 (N_39048,N_37225,N_36578);
nor U39049 (N_39049,N_35668,N_36504);
and U39050 (N_39050,N_35276,N_35310);
nand U39051 (N_39051,N_35148,N_37495);
nand U39052 (N_39052,N_36570,N_35943);
nand U39053 (N_39053,N_36512,N_35816);
nor U39054 (N_39054,N_36877,N_35255);
and U39055 (N_39055,N_35790,N_37217);
nor U39056 (N_39056,N_37319,N_37282);
and U39057 (N_39057,N_36527,N_35905);
or U39058 (N_39058,N_35505,N_37171);
nor U39059 (N_39059,N_35439,N_35993);
nor U39060 (N_39060,N_36938,N_36682);
or U39061 (N_39061,N_36227,N_35742);
and U39062 (N_39062,N_35688,N_35871);
nand U39063 (N_39063,N_35462,N_37048);
nor U39064 (N_39064,N_36521,N_35064);
xor U39065 (N_39065,N_35169,N_35136);
nand U39066 (N_39066,N_36723,N_36323);
and U39067 (N_39067,N_36083,N_37063);
and U39068 (N_39068,N_35403,N_35637);
nor U39069 (N_39069,N_35411,N_35423);
and U39070 (N_39070,N_36570,N_36638);
and U39071 (N_39071,N_35348,N_36845);
or U39072 (N_39072,N_35837,N_36721);
nor U39073 (N_39073,N_37168,N_36828);
and U39074 (N_39074,N_37417,N_37087);
xor U39075 (N_39075,N_35409,N_37347);
and U39076 (N_39076,N_36467,N_37390);
nor U39077 (N_39077,N_35977,N_37380);
nand U39078 (N_39078,N_36552,N_35155);
xor U39079 (N_39079,N_36376,N_36380);
nand U39080 (N_39080,N_35298,N_36738);
nand U39081 (N_39081,N_35225,N_37491);
and U39082 (N_39082,N_35024,N_37444);
or U39083 (N_39083,N_35314,N_35333);
or U39084 (N_39084,N_37400,N_37451);
xnor U39085 (N_39085,N_36811,N_36895);
or U39086 (N_39086,N_35107,N_35031);
nand U39087 (N_39087,N_35859,N_35225);
nor U39088 (N_39088,N_36406,N_35881);
or U39089 (N_39089,N_35917,N_36660);
xnor U39090 (N_39090,N_37205,N_36758);
nor U39091 (N_39091,N_35417,N_37123);
and U39092 (N_39092,N_35081,N_35379);
nand U39093 (N_39093,N_37034,N_36755);
nor U39094 (N_39094,N_35718,N_36338);
and U39095 (N_39095,N_36130,N_35834);
or U39096 (N_39096,N_36240,N_35208);
nand U39097 (N_39097,N_36732,N_35677);
nor U39098 (N_39098,N_36028,N_35408);
nor U39099 (N_39099,N_35283,N_35137);
and U39100 (N_39100,N_35532,N_36528);
and U39101 (N_39101,N_35554,N_37334);
or U39102 (N_39102,N_36528,N_37428);
nand U39103 (N_39103,N_37307,N_36852);
xor U39104 (N_39104,N_35441,N_36563);
and U39105 (N_39105,N_36052,N_35069);
nor U39106 (N_39106,N_35804,N_37223);
nand U39107 (N_39107,N_35214,N_37383);
and U39108 (N_39108,N_37379,N_37016);
nor U39109 (N_39109,N_35107,N_35825);
nand U39110 (N_39110,N_37270,N_35405);
nor U39111 (N_39111,N_36922,N_37270);
or U39112 (N_39112,N_36271,N_35545);
nand U39113 (N_39113,N_36975,N_36166);
nand U39114 (N_39114,N_36717,N_35901);
or U39115 (N_39115,N_35560,N_35044);
or U39116 (N_39116,N_37362,N_35289);
and U39117 (N_39117,N_35774,N_36422);
or U39118 (N_39118,N_36313,N_35294);
xnor U39119 (N_39119,N_36247,N_36327);
nor U39120 (N_39120,N_37215,N_35254);
and U39121 (N_39121,N_36447,N_35495);
and U39122 (N_39122,N_37201,N_37021);
and U39123 (N_39123,N_36912,N_35771);
and U39124 (N_39124,N_36422,N_36736);
and U39125 (N_39125,N_37328,N_37330);
or U39126 (N_39126,N_35856,N_35157);
or U39127 (N_39127,N_36907,N_35807);
nor U39128 (N_39128,N_35323,N_35186);
nand U39129 (N_39129,N_36637,N_35370);
nor U39130 (N_39130,N_35444,N_36078);
nand U39131 (N_39131,N_35345,N_36605);
or U39132 (N_39132,N_35788,N_37395);
and U39133 (N_39133,N_36585,N_35380);
nor U39134 (N_39134,N_35010,N_37114);
or U39135 (N_39135,N_35430,N_37014);
and U39136 (N_39136,N_35143,N_36698);
nand U39137 (N_39137,N_36463,N_37249);
nor U39138 (N_39138,N_36208,N_37413);
or U39139 (N_39139,N_35234,N_36352);
nand U39140 (N_39140,N_35680,N_37189);
xor U39141 (N_39141,N_36288,N_35282);
nor U39142 (N_39142,N_36023,N_36835);
nand U39143 (N_39143,N_37429,N_36856);
nor U39144 (N_39144,N_35030,N_36297);
and U39145 (N_39145,N_36784,N_36714);
nand U39146 (N_39146,N_35779,N_35226);
nor U39147 (N_39147,N_35262,N_35569);
nand U39148 (N_39148,N_37143,N_35116);
xnor U39149 (N_39149,N_37152,N_36859);
or U39150 (N_39150,N_35108,N_36912);
nand U39151 (N_39151,N_35738,N_37161);
nand U39152 (N_39152,N_37303,N_35128);
nor U39153 (N_39153,N_35821,N_35968);
xnor U39154 (N_39154,N_37229,N_37454);
and U39155 (N_39155,N_37448,N_36131);
or U39156 (N_39156,N_36921,N_36739);
nand U39157 (N_39157,N_37452,N_37381);
or U39158 (N_39158,N_35086,N_37138);
or U39159 (N_39159,N_36786,N_35291);
nor U39160 (N_39160,N_36328,N_36173);
nor U39161 (N_39161,N_35276,N_36165);
nor U39162 (N_39162,N_35961,N_36470);
nand U39163 (N_39163,N_37348,N_35919);
nand U39164 (N_39164,N_35923,N_36765);
nor U39165 (N_39165,N_36159,N_36648);
nand U39166 (N_39166,N_35872,N_35431);
nand U39167 (N_39167,N_35601,N_35854);
nand U39168 (N_39168,N_36297,N_35354);
or U39169 (N_39169,N_35560,N_36738);
nand U39170 (N_39170,N_36887,N_36855);
xor U39171 (N_39171,N_35122,N_37408);
or U39172 (N_39172,N_36846,N_36842);
nor U39173 (N_39173,N_36134,N_36374);
nand U39174 (N_39174,N_35818,N_37265);
and U39175 (N_39175,N_35772,N_36446);
nand U39176 (N_39176,N_37242,N_35712);
and U39177 (N_39177,N_36753,N_35506);
or U39178 (N_39178,N_35215,N_35776);
nand U39179 (N_39179,N_35371,N_36122);
and U39180 (N_39180,N_37257,N_35309);
xor U39181 (N_39181,N_35921,N_37096);
or U39182 (N_39182,N_35841,N_35033);
nand U39183 (N_39183,N_37016,N_36588);
nand U39184 (N_39184,N_35768,N_36587);
nand U39185 (N_39185,N_35011,N_35689);
nor U39186 (N_39186,N_35885,N_35263);
nor U39187 (N_39187,N_36678,N_36813);
nor U39188 (N_39188,N_36453,N_36132);
nand U39189 (N_39189,N_35689,N_36275);
nand U39190 (N_39190,N_35758,N_35714);
or U39191 (N_39191,N_35386,N_35625);
or U39192 (N_39192,N_35527,N_35574);
or U39193 (N_39193,N_35300,N_36748);
and U39194 (N_39194,N_37396,N_37005);
and U39195 (N_39195,N_35222,N_37329);
nor U39196 (N_39196,N_35269,N_37133);
nor U39197 (N_39197,N_37178,N_35060);
and U39198 (N_39198,N_35355,N_36262);
nor U39199 (N_39199,N_36947,N_36563);
nor U39200 (N_39200,N_36470,N_35219);
nand U39201 (N_39201,N_35258,N_35439);
nor U39202 (N_39202,N_35935,N_36652);
nand U39203 (N_39203,N_35462,N_36483);
nor U39204 (N_39204,N_36782,N_37368);
nand U39205 (N_39205,N_35040,N_35448);
and U39206 (N_39206,N_35312,N_35375);
xor U39207 (N_39207,N_36943,N_36142);
and U39208 (N_39208,N_35024,N_35126);
and U39209 (N_39209,N_37127,N_35189);
nand U39210 (N_39210,N_36072,N_35299);
nor U39211 (N_39211,N_36190,N_35622);
and U39212 (N_39212,N_36548,N_35757);
xnor U39213 (N_39213,N_36859,N_36832);
or U39214 (N_39214,N_35309,N_36106);
and U39215 (N_39215,N_35017,N_35537);
nand U39216 (N_39216,N_36986,N_37143);
or U39217 (N_39217,N_37027,N_36490);
nor U39218 (N_39218,N_37242,N_36129);
xor U39219 (N_39219,N_36423,N_36425);
nor U39220 (N_39220,N_35342,N_35076);
nand U39221 (N_39221,N_37096,N_35565);
and U39222 (N_39222,N_37111,N_36330);
xor U39223 (N_39223,N_35615,N_36777);
nand U39224 (N_39224,N_36973,N_36270);
nand U39225 (N_39225,N_36849,N_36797);
nand U39226 (N_39226,N_36403,N_36296);
nand U39227 (N_39227,N_36211,N_36392);
and U39228 (N_39228,N_36298,N_35131);
or U39229 (N_39229,N_36870,N_37154);
or U39230 (N_39230,N_36674,N_36788);
nand U39231 (N_39231,N_36374,N_35175);
nand U39232 (N_39232,N_36830,N_37359);
or U39233 (N_39233,N_36537,N_35593);
or U39234 (N_39234,N_35276,N_37479);
and U39235 (N_39235,N_36222,N_35258);
or U39236 (N_39236,N_36790,N_36670);
and U39237 (N_39237,N_36462,N_36217);
or U39238 (N_39238,N_37086,N_36830);
and U39239 (N_39239,N_36042,N_35669);
nand U39240 (N_39240,N_37330,N_36287);
nor U39241 (N_39241,N_35801,N_36105);
nand U39242 (N_39242,N_36483,N_35515);
nor U39243 (N_39243,N_37208,N_36004);
nand U39244 (N_39244,N_35553,N_36960);
and U39245 (N_39245,N_36791,N_35867);
nand U39246 (N_39246,N_36790,N_35785);
and U39247 (N_39247,N_36710,N_36035);
nand U39248 (N_39248,N_35674,N_36623);
nand U39249 (N_39249,N_35124,N_37329);
and U39250 (N_39250,N_35905,N_37355);
xnor U39251 (N_39251,N_36762,N_36987);
and U39252 (N_39252,N_36953,N_35509);
nor U39253 (N_39253,N_37289,N_35782);
or U39254 (N_39254,N_36206,N_36600);
and U39255 (N_39255,N_35675,N_35185);
nand U39256 (N_39256,N_36534,N_36098);
nand U39257 (N_39257,N_37259,N_35639);
xnor U39258 (N_39258,N_36439,N_36496);
and U39259 (N_39259,N_36803,N_35531);
and U39260 (N_39260,N_36458,N_36898);
or U39261 (N_39261,N_37280,N_37308);
and U39262 (N_39262,N_35862,N_35627);
and U39263 (N_39263,N_36653,N_35133);
and U39264 (N_39264,N_35370,N_36459);
and U39265 (N_39265,N_36276,N_35327);
xor U39266 (N_39266,N_36614,N_35609);
xnor U39267 (N_39267,N_36421,N_36145);
or U39268 (N_39268,N_36025,N_36336);
nand U39269 (N_39269,N_37099,N_35354);
xnor U39270 (N_39270,N_35363,N_36783);
nand U39271 (N_39271,N_35091,N_36757);
or U39272 (N_39272,N_35995,N_36003);
nor U39273 (N_39273,N_36599,N_37285);
nor U39274 (N_39274,N_36369,N_35552);
nand U39275 (N_39275,N_36438,N_36891);
nor U39276 (N_39276,N_36536,N_35425);
nor U39277 (N_39277,N_35771,N_35305);
or U39278 (N_39278,N_35843,N_36479);
or U39279 (N_39279,N_35249,N_36855);
and U39280 (N_39280,N_36089,N_36116);
nor U39281 (N_39281,N_35820,N_36871);
nand U39282 (N_39282,N_35355,N_36937);
xor U39283 (N_39283,N_36804,N_37115);
or U39284 (N_39284,N_36411,N_37046);
nand U39285 (N_39285,N_37264,N_35392);
and U39286 (N_39286,N_35660,N_37488);
nand U39287 (N_39287,N_36679,N_36216);
nor U39288 (N_39288,N_35874,N_35185);
nor U39289 (N_39289,N_37176,N_37485);
nor U39290 (N_39290,N_35013,N_37474);
and U39291 (N_39291,N_37269,N_36191);
and U39292 (N_39292,N_37321,N_35598);
or U39293 (N_39293,N_36796,N_36596);
nand U39294 (N_39294,N_35400,N_35249);
and U39295 (N_39295,N_36098,N_35096);
nor U39296 (N_39296,N_36511,N_35048);
nand U39297 (N_39297,N_36084,N_35896);
xnor U39298 (N_39298,N_35618,N_35812);
nand U39299 (N_39299,N_35003,N_36893);
nor U39300 (N_39300,N_36934,N_35482);
or U39301 (N_39301,N_35857,N_37185);
or U39302 (N_39302,N_37119,N_37013);
nand U39303 (N_39303,N_37421,N_36133);
nor U39304 (N_39304,N_35272,N_35017);
xor U39305 (N_39305,N_35717,N_35168);
nor U39306 (N_39306,N_37268,N_35195);
nor U39307 (N_39307,N_35379,N_35031);
or U39308 (N_39308,N_36977,N_35927);
and U39309 (N_39309,N_36298,N_36818);
nor U39310 (N_39310,N_35589,N_36105);
nor U39311 (N_39311,N_36141,N_36095);
nand U39312 (N_39312,N_35359,N_36193);
nor U39313 (N_39313,N_36726,N_36470);
nand U39314 (N_39314,N_36566,N_35451);
or U39315 (N_39315,N_36552,N_37171);
xor U39316 (N_39316,N_37305,N_36282);
nand U39317 (N_39317,N_35082,N_36418);
nand U39318 (N_39318,N_35176,N_36909);
nor U39319 (N_39319,N_37038,N_36192);
nor U39320 (N_39320,N_35511,N_36576);
and U39321 (N_39321,N_35795,N_37369);
and U39322 (N_39322,N_35831,N_36247);
nand U39323 (N_39323,N_37194,N_37121);
and U39324 (N_39324,N_35272,N_35101);
nand U39325 (N_39325,N_36358,N_37392);
or U39326 (N_39326,N_37384,N_36091);
and U39327 (N_39327,N_36075,N_36732);
and U39328 (N_39328,N_36670,N_36813);
or U39329 (N_39329,N_36027,N_36015);
nor U39330 (N_39330,N_35852,N_35574);
or U39331 (N_39331,N_36898,N_35715);
xor U39332 (N_39332,N_36875,N_35766);
or U39333 (N_39333,N_36806,N_36942);
xor U39334 (N_39334,N_37334,N_36212);
and U39335 (N_39335,N_36578,N_35933);
or U39336 (N_39336,N_35594,N_35633);
nor U39337 (N_39337,N_37330,N_36133);
or U39338 (N_39338,N_36163,N_35188);
and U39339 (N_39339,N_36474,N_35505);
and U39340 (N_39340,N_36662,N_35451);
and U39341 (N_39341,N_37019,N_36739);
nor U39342 (N_39342,N_35587,N_37065);
and U39343 (N_39343,N_35875,N_35543);
xnor U39344 (N_39344,N_35102,N_36002);
or U39345 (N_39345,N_35379,N_36190);
xnor U39346 (N_39346,N_35251,N_36357);
nor U39347 (N_39347,N_37047,N_36565);
and U39348 (N_39348,N_36574,N_36244);
and U39349 (N_39349,N_36989,N_35651);
nor U39350 (N_39350,N_36189,N_35639);
nor U39351 (N_39351,N_35663,N_37136);
nor U39352 (N_39352,N_35298,N_35519);
or U39353 (N_39353,N_35684,N_36375);
nand U39354 (N_39354,N_37484,N_36002);
and U39355 (N_39355,N_36834,N_35144);
nand U39356 (N_39356,N_37251,N_35562);
nor U39357 (N_39357,N_37086,N_35979);
nand U39358 (N_39358,N_35863,N_35038);
or U39359 (N_39359,N_37044,N_36017);
nor U39360 (N_39360,N_37278,N_35089);
nor U39361 (N_39361,N_36250,N_37174);
or U39362 (N_39362,N_36029,N_36200);
nor U39363 (N_39363,N_36404,N_35516);
nor U39364 (N_39364,N_35755,N_35966);
or U39365 (N_39365,N_36199,N_36740);
or U39366 (N_39366,N_36605,N_35253);
xnor U39367 (N_39367,N_36394,N_36673);
xnor U39368 (N_39368,N_35500,N_36806);
and U39369 (N_39369,N_36664,N_35192);
nor U39370 (N_39370,N_36738,N_35027);
and U39371 (N_39371,N_35938,N_35041);
nor U39372 (N_39372,N_35293,N_35411);
and U39373 (N_39373,N_36342,N_35613);
nand U39374 (N_39374,N_35862,N_36483);
nor U39375 (N_39375,N_36711,N_35822);
and U39376 (N_39376,N_36321,N_36638);
or U39377 (N_39377,N_36190,N_36260);
nand U39378 (N_39378,N_36589,N_35004);
and U39379 (N_39379,N_36305,N_37398);
nand U39380 (N_39380,N_37242,N_37341);
and U39381 (N_39381,N_37148,N_36128);
or U39382 (N_39382,N_35920,N_36406);
nand U39383 (N_39383,N_36860,N_36385);
nor U39384 (N_39384,N_36048,N_37097);
nor U39385 (N_39385,N_35012,N_35352);
or U39386 (N_39386,N_35277,N_35843);
and U39387 (N_39387,N_36758,N_35853);
and U39388 (N_39388,N_36985,N_37412);
nor U39389 (N_39389,N_36810,N_36784);
and U39390 (N_39390,N_36430,N_37437);
nor U39391 (N_39391,N_35859,N_35428);
nand U39392 (N_39392,N_35762,N_36362);
and U39393 (N_39393,N_37158,N_35719);
and U39394 (N_39394,N_36386,N_36278);
nand U39395 (N_39395,N_36553,N_36208);
and U39396 (N_39396,N_36633,N_36634);
and U39397 (N_39397,N_36381,N_36472);
and U39398 (N_39398,N_36542,N_36075);
xnor U39399 (N_39399,N_36097,N_35657);
xor U39400 (N_39400,N_37071,N_35745);
nor U39401 (N_39401,N_36519,N_36884);
xor U39402 (N_39402,N_35149,N_36962);
xor U39403 (N_39403,N_36892,N_36135);
or U39404 (N_39404,N_35602,N_35078);
or U39405 (N_39405,N_36472,N_36444);
or U39406 (N_39406,N_37146,N_36954);
nand U39407 (N_39407,N_37056,N_35951);
nor U39408 (N_39408,N_36208,N_35318);
nor U39409 (N_39409,N_35035,N_36499);
and U39410 (N_39410,N_35737,N_36683);
or U39411 (N_39411,N_37135,N_36310);
nor U39412 (N_39412,N_36471,N_35511);
and U39413 (N_39413,N_36575,N_37162);
or U39414 (N_39414,N_35900,N_36060);
nor U39415 (N_39415,N_37020,N_35398);
and U39416 (N_39416,N_35142,N_35205);
xnor U39417 (N_39417,N_37334,N_36449);
or U39418 (N_39418,N_37227,N_35534);
nand U39419 (N_39419,N_35275,N_35470);
and U39420 (N_39420,N_37421,N_36391);
or U39421 (N_39421,N_36058,N_37431);
or U39422 (N_39422,N_37301,N_35011);
nand U39423 (N_39423,N_35589,N_36259);
and U39424 (N_39424,N_37274,N_35028);
and U39425 (N_39425,N_35404,N_35216);
nor U39426 (N_39426,N_36449,N_35712);
nor U39427 (N_39427,N_36286,N_35555);
nor U39428 (N_39428,N_37238,N_36747);
and U39429 (N_39429,N_35655,N_37439);
or U39430 (N_39430,N_37364,N_35104);
nand U39431 (N_39431,N_37271,N_35415);
and U39432 (N_39432,N_37112,N_36315);
and U39433 (N_39433,N_35113,N_35383);
nor U39434 (N_39434,N_35208,N_36245);
nand U39435 (N_39435,N_35346,N_35332);
nor U39436 (N_39436,N_37429,N_36005);
or U39437 (N_39437,N_35700,N_35213);
nand U39438 (N_39438,N_35416,N_35095);
or U39439 (N_39439,N_37382,N_36784);
xor U39440 (N_39440,N_36810,N_35195);
xor U39441 (N_39441,N_36294,N_35196);
nor U39442 (N_39442,N_36034,N_37181);
nand U39443 (N_39443,N_35353,N_36741);
nor U39444 (N_39444,N_35260,N_36423);
and U39445 (N_39445,N_36823,N_37041);
nor U39446 (N_39446,N_36693,N_36833);
nor U39447 (N_39447,N_35322,N_36951);
or U39448 (N_39448,N_36958,N_35952);
or U39449 (N_39449,N_36354,N_35293);
nand U39450 (N_39450,N_36702,N_35654);
xor U39451 (N_39451,N_35016,N_36892);
nand U39452 (N_39452,N_36176,N_37249);
and U39453 (N_39453,N_36038,N_35543);
nand U39454 (N_39454,N_36661,N_36305);
nand U39455 (N_39455,N_35282,N_37232);
and U39456 (N_39456,N_37314,N_37109);
or U39457 (N_39457,N_35800,N_35104);
or U39458 (N_39458,N_36594,N_36680);
xnor U39459 (N_39459,N_35443,N_37479);
nor U39460 (N_39460,N_35121,N_37356);
nor U39461 (N_39461,N_35722,N_36298);
nand U39462 (N_39462,N_36443,N_35869);
and U39463 (N_39463,N_36986,N_37461);
nand U39464 (N_39464,N_35776,N_36329);
or U39465 (N_39465,N_36656,N_37133);
nand U39466 (N_39466,N_37299,N_36225);
nor U39467 (N_39467,N_36575,N_36084);
and U39468 (N_39468,N_35801,N_37026);
nor U39469 (N_39469,N_36666,N_35508);
and U39470 (N_39470,N_35154,N_35620);
nor U39471 (N_39471,N_35536,N_36654);
or U39472 (N_39472,N_36481,N_37436);
and U39473 (N_39473,N_35544,N_35843);
or U39474 (N_39474,N_36415,N_35311);
nand U39475 (N_39475,N_36598,N_35856);
nand U39476 (N_39476,N_35140,N_37212);
and U39477 (N_39477,N_37054,N_36074);
nor U39478 (N_39478,N_35707,N_36975);
xnor U39479 (N_39479,N_37167,N_36659);
or U39480 (N_39480,N_35247,N_35240);
nor U39481 (N_39481,N_36958,N_35815);
or U39482 (N_39482,N_35571,N_37366);
nand U39483 (N_39483,N_36249,N_36268);
nor U39484 (N_39484,N_36617,N_35586);
nand U39485 (N_39485,N_36500,N_36616);
nand U39486 (N_39486,N_35934,N_35445);
and U39487 (N_39487,N_36601,N_37059);
xnor U39488 (N_39488,N_36068,N_37408);
nor U39489 (N_39489,N_35831,N_37440);
and U39490 (N_39490,N_36949,N_35669);
nand U39491 (N_39491,N_37182,N_36735);
nor U39492 (N_39492,N_36792,N_36418);
xor U39493 (N_39493,N_37424,N_36526);
or U39494 (N_39494,N_35070,N_36764);
or U39495 (N_39495,N_36259,N_35207);
or U39496 (N_39496,N_35363,N_37308);
xor U39497 (N_39497,N_36139,N_36039);
nor U39498 (N_39498,N_35402,N_37193);
nor U39499 (N_39499,N_36046,N_37254);
and U39500 (N_39500,N_36788,N_36257);
or U39501 (N_39501,N_35483,N_35346);
nor U39502 (N_39502,N_36876,N_35092);
and U39503 (N_39503,N_36337,N_36941);
and U39504 (N_39504,N_36536,N_35507);
and U39505 (N_39505,N_36596,N_35480);
nor U39506 (N_39506,N_35131,N_37407);
nor U39507 (N_39507,N_35094,N_35585);
nand U39508 (N_39508,N_35591,N_37030);
nand U39509 (N_39509,N_35097,N_36135);
nor U39510 (N_39510,N_37388,N_36409);
nor U39511 (N_39511,N_35497,N_36430);
and U39512 (N_39512,N_36719,N_35854);
nand U39513 (N_39513,N_36036,N_35176);
and U39514 (N_39514,N_36549,N_37409);
nand U39515 (N_39515,N_36504,N_36749);
nor U39516 (N_39516,N_35575,N_36101);
nor U39517 (N_39517,N_36241,N_35869);
nor U39518 (N_39518,N_36709,N_35730);
nor U39519 (N_39519,N_35839,N_37006);
or U39520 (N_39520,N_35414,N_37326);
nor U39521 (N_39521,N_37289,N_35948);
xor U39522 (N_39522,N_37047,N_37262);
and U39523 (N_39523,N_36909,N_36982);
nand U39524 (N_39524,N_37111,N_37156);
or U39525 (N_39525,N_36236,N_37403);
nor U39526 (N_39526,N_36059,N_35027);
or U39527 (N_39527,N_35848,N_35933);
xnor U39528 (N_39528,N_35387,N_37399);
or U39529 (N_39529,N_35207,N_37317);
nand U39530 (N_39530,N_37219,N_36610);
nand U39531 (N_39531,N_35944,N_35861);
nand U39532 (N_39532,N_37232,N_37202);
and U39533 (N_39533,N_36695,N_35806);
and U39534 (N_39534,N_36438,N_35043);
or U39535 (N_39535,N_36566,N_36338);
xor U39536 (N_39536,N_37254,N_37111);
nor U39537 (N_39537,N_35648,N_35973);
nor U39538 (N_39538,N_36379,N_37048);
or U39539 (N_39539,N_35036,N_35451);
nand U39540 (N_39540,N_36119,N_36171);
and U39541 (N_39541,N_37210,N_35079);
nand U39542 (N_39542,N_36651,N_36711);
nor U39543 (N_39543,N_36274,N_35516);
nand U39544 (N_39544,N_37137,N_37052);
and U39545 (N_39545,N_36167,N_36721);
nor U39546 (N_39546,N_37235,N_35505);
or U39547 (N_39547,N_37267,N_36030);
and U39548 (N_39548,N_36412,N_37406);
and U39549 (N_39549,N_36308,N_37249);
nand U39550 (N_39550,N_36765,N_35900);
nand U39551 (N_39551,N_37109,N_36603);
and U39552 (N_39552,N_35799,N_36563);
and U39553 (N_39553,N_36708,N_37231);
and U39554 (N_39554,N_37140,N_35522);
xor U39555 (N_39555,N_36807,N_35490);
nand U39556 (N_39556,N_37414,N_36244);
nor U39557 (N_39557,N_35263,N_36286);
and U39558 (N_39558,N_37180,N_35422);
nand U39559 (N_39559,N_36507,N_36776);
xnor U39560 (N_39560,N_36342,N_36470);
and U39561 (N_39561,N_35592,N_35461);
and U39562 (N_39562,N_36140,N_35067);
and U39563 (N_39563,N_35499,N_35783);
nand U39564 (N_39564,N_37321,N_35048);
or U39565 (N_39565,N_36720,N_37317);
nand U39566 (N_39566,N_36215,N_37121);
xnor U39567 (N_39567,N_37344,N_35787);
and U39568 (N_39568,N_35901,N_36873);
or U39569 (N_39569,N_35626,N_36363);
nand U39570 (N_39570,N_36442,N_35031);
nor U39571 (N_39571,N_36809,N_37403);
nor U39572 (N_39572,N_35575,N_37485);
nor U39573 (N_39573,N_36779,N_35969);
or U39574 (N_39574,N_37092,N_36493);
and U39575 (N_39575,N_35236,N_36782);
nor U39576 (N_39576,N_36509,N_35530);
nand U39577 (N_39577,N_36109,N_36161);
nor U39578 (N_39578,N_35664,N_37491);
and U39579 (N_39579,N_36620,N_35892);
nor U39580 (N_39580,N_35176,N_36166);
nor U39581 (N_39581,N_35576,N_36046);
nor U39582 (N_39582,N_36476,N_36460);
or U39583 (N_39583,N_37361,N_36121);
nand U39584 (N_39584,N_35566,N_37401);
nor U39585 (N_39585,N_36157,N_37395);
or U39586 (N_39586,N_36657,N_37465);
and U39587 (N_39587,N_36627,N_35257);
or U39588 (N_39588,N_35233,N_36006);
xor U39589 (N_39589,N_36196,N_36379);
and U39590 (N_39590,N_35319,N_35929);
or U39591 (N_39591,N_36454,N_36855);
and U39592 (N_39592,N_36347,N_37080);
or U39593 (N_39593,N_35449,N_35215);
nand U39594 (N_39594,N_36201,N_37149);
and U39595 (N_39595,N_37426,N_35687);
nand U39596 (N_39596,N_35500,N_35452);
nor U39597 (N_39597,N_36332,N_35853);
nor U39598 (N_39598,N_37000,N_35434);
nand U39599 (N_39599,N_37419,N_35575);
or U39600 (N_39600,N_37480,N_35205);
nor U39601 (N_39601,N_35437,N_35089);
xor U39602 (N_39602,N_35647,N_35298);
nand U39603 (N_39603,N_35984,N_37155);
nor U39604 (N_39604,N_36279,N_36231);
or U39605 (N_39605,N_35602,N_36882);
and U39606 (N_39606,N_36413,N_36961);
and U39607 (N_39607,N_36428,N_35801);
xor U39608 (N_39608,N_36154,N_36896);
xnor U39609 (N_39609,N_36075,N_37385);
nor U39610 (N_39610,N_35408,N_37265);
nor U39611 (N_39611,N_36334,N_37289);
or U39612 (N_39612,N_35863,N_36574);
nor U39613 (N_39613,N_37002,N_36485);
and U39614 (N_39614,N_36322,N_37237);
or U39615 (N_39615,N_37461,N_36645);
xnor U39616 (N_39616,N_36176,N_36428);
or U39617 (N_39617,N_35900,N_35102);
nor U39618 (N_39618,N_36099,N_36261);
and U39619 (N_39619,N_36247,N_37248);
or U39620 (N_39620,N_37265,N_35543);
or U39621 (N_39621,N_36694,N_36526);
nand U39622 (N_39622,N_35844,N_37013);
nor U39623 (N_39623,N_37177,N_35115);
and U39624 (N_39624,N_35750,N_36868);
nor U39625 (N_39625,N_36259,N_37211);
nand U39626 (N_39626,N_35271,N_36599);
or U39627 (N_39627,N_35288,N_36109);
or U39628 (N_39628,N_36014,N_36128);
xor U39629 (N_39629,N_36562,N_35333);
nor U39630 (N_39630,N_36723,N_35601);
nor U39631 (N_39631,N_36234,N_36058);
nand U39632 (N_39632,N_35469,N_35948);
nor U39633 (N_39633,N_36472,N_36861);
xnor U39634 (N_39634,N_37107,N_37175);
or U39635 (N_39635,N_36920,N_36210);
nor U39636 (N_39636,N_35594,N_35813);
nand U39637 (N_39637,N_36276,N_36946);
nand U39638 (N_39638,N_36910,N_36840);
nand U39639 (N_39639,N_35287,N_36062);
nor U39640 (N_39640,N_37026,N_35070);
and U39641 (N_39641,N_37471,N_35243);
or U39642 (N_39642,N_35491,N_35560);
nor U39643 (N_39643,N_36922,N_37073);
nand U39644 (N_39644,N_35106,N_35231);
nand U39645 (N_39645,N_35758,N_35215);
nor U39646 (N_39646,N_35544,N_35946);
xnor U39647 (N_39647,N_35662,N_36600);
nand U39648 (N_39648,N_36503,N_35438);
xor U39649 (N_39649,N_37067,N_37038);
xnor U39650 (N_39650,N_36322,N_37219);
nand U39651 (N_39651,N_37480,N_36495);
nand U39652 (N_39652,N_35033,N_36695);
nor U39653 (N_39653,N_36923,N_36456);
nor U39654 (N_39654,N_35199,N_35105);
nand U39655 (N_39655,N_35154,N_36733);
nor U39656 (N_39656,N_35149,N_36679);
and U39657 (N_39657,N_36368,N_37378);
or U39658 (N_39658,N_37337,N_36249);
nor U39659 (N_39659,N_35643,N_35330);
and U39660 (N_39660,N_36207,N_35950);
nor U39661 (N_39661,N_35287,N_36800);
or U39662 (N_39662,N_35305,N_37359);
xnor U39663 (N_39663,N_36913,N_36596);
and U39664 (N_39664,N_35791,N_36743);
nor U39665 (N_39665,N_35242,N_37475);
or U39666 (N_39666,N_35051,N_36775);
xor U39667 (N_39667,N_36324,N_37384);
or U39668 (N_39668,N_36957,N_36856);
nor U39669 (N_39669,N_35880,N_36420);
nand U39670 (N_39670,N_36978,N_35745);
nand U39671 (N_39671,N_35847,N_36638);
xor U39672 (N_39672,N_36084,N_37054);
and U39673 (N_39673,N_36596,N_35098);
and U39674 (N_39674,N_35659,N_35993);
nor U39675 (N_39675,N_35440,N_37155);
or U39676 (N_39676,N_36137,N_36725);
nor U39677 (N_39677,N_36198,N_35221);
and U39678 (N_39678,N_35693,N_35062);
or U39679 (N_39679,N_35117,N_37081);
xnor U39680 (N_39680,N_36794,N_36633);
nand U39681 (N_39681,N_36568,N_36496);
and U39682 (N_39682,N_36028,N_35296);
and U39683 (N_39683,N_36082,N_36537);
or U39684 (N_39684,N_35247,N_36067);
nand U39685 (N_39685,N_35954,N_35585);
nand U39686 (N_39686,N_35956,N_35568);
xor U39687 (N_39687,N_35569,N_36356);
or U39688 (N_39688,N_35222,N_36627);
xor U39689 (N_39689,N_35342,N_37483);
nand U39690 (N_39690,N_35931,N_37198);
and U39691 (N_39691,N_36121,N_35324);
nor U39692 (N_39692,N_37462,N_36799);
or U39693 (N_39693,N_36318,N_35029);
xor U39694 (N_39694,N_35713,N_35841);
xor U39695 (N_39695,N_37493,N_37404);
and U39696 (N_39696,N_35613,N_35796);
nor U39697 (N_39697,N_35895,N_36830);
and U39698 (N_39698,N_37404,N_37110);
or U39699 (N_39699,N_37032,N_36492);
and U39700 (N_39700,N_36956,N_35402);
nand U39701 (N_39701,N_37140,N_35011);
and U39702 (N_39702,N_36599,N_35909);
or U39703 (N_39703,N_36472,N_35847);
nand U39704 (N_39704,N_35015,N_35726);
or U39705 (N_39705,N_36745,N_36919);
nor U39706 (N_39706,N_35103,N_35819);
or U39707 (N_39707,N_36294,N_35390);
or U39708 (N_39708,N_37464,N_35788);
nand U39709 (N_39709,N_35991,N_36041);
or U39710 (N_39710,N_37090,N_35655);
and U39711 (N_39711,N_36667,N_35191);
and U39712 (N_39712,N_36390,N_36314);
nand U39713 (N_39713,N_35984,N_37245);
xnor U39714 (N_39714,N_35190,N_36550);
nand U39715 (N_39715,N_37060,N_36380);
nand U39716 (N_39716,N_35921,N_36472);
nand U39717 (N_39717,N_37245,N_37110);
nor U39718 (N_39718,N_36045,N_35007);
nor U39719 (N_39719,N_36351,N_36277);
nor U39720 (N_39720,N_35023,N_37005);
xnor U39721 (N_39721,N_36727,N_35878);
nand U39722 (N_39722,N_36144,N_36655);
or U39723 (N_39723,N_36962,N_37096);
and U39724 (N_39724,N_35852,N_36729);
nand U39725 (N_39725,N_37250,N_36609);
and U39726 (N_39726,N_35513,N_37372);
or U39727 (N_39727,N_37010,N_35898);
or U39728 (N_39728,N_36037,N_36896);
nor U39729 (N_39729,N_37403,N_36009);
or U39730 (N_39730,N_36412,N_37315);
xnor U39731 (N_39731,N_35077,N_35739);
nor U39732 (N_39732,N_35463,N_35055);
nor U39733 (N_39733,N_35503,N_35539);
nand U39734 (N_39734,N_35184,N_37097);
xor U39735 (N_39735,N_36897,N_37145);
or U39736 (N_39736,N_36082,N_35544);
or U39737 (N_39737,N_35269,N_37221);
nor U39738 (N_39738,N_35035,N_35640);
nor U39739 (N_39739,N_36476,N_35063);
or U39740 (N_39740,N_36059,N_36859);
nand U39741 (N_39741,N_35772,N_35367);
and U39742 (N_39742,N_37347,N_35618);
nand U39743 (N_39743,N_35241,N_36262);
and U39744 (N_39744,N_35999,N_36418);
nand U39745 (N_39745,N_36890,N_35936);
nand U39746 (N_39746,N_36601,N_36136);
and U39747 (N_39747,N_36374,N_37422);
or U39748 (N_39748,N_36591,N_36238);
nand U39749 (N_39749,N_35959,N_35335);
and U39750 (N_39750,N_37072,N_35437);
or U39751 (N_39751,N_35576,N_35313);
nor U39752 (N_39752,N_37032,N_37479);
nor U39753 (N_39753,N_37222,N_36984);
and U39754 (N_39754,N_35703,N_35052);
nor U39755 (N_39755,N_35034,N_35579);
nand U39756 (N_39756,N_36408,N_36338);
nor U39757 (N_39757,N_36242,N_36988);
and U39758 (N_39758,N_36810,N_36841);
nor U39759 (N_39759,N_36177,N_36297);
xor U39760 (N_39760,N_37463,N_36533);
and U39761 (N_39761,N_35724,N_37290);
or U39762 (N_39762,N_37372,N_36872);
and U39763 (N_39763,N_36541,N_35964);
and U39764 (N_39764,N_37019,N_37388);
or U39765 (N_39765,N_35569,N_35321);
and U39766 (N_39766,N_35436,N_36349);
nor U39767 (N_39767,N_35370,N_35368);
nand U39768 (N_39768,N_37139,N_36539);
and U39769 (N_39769,N_35078,N_37309);
nor U39770 (N_39770,N_36597,N_36734);
and U39771 (N_39771,N_37493,N_37140);
nand U39772 (N_39772,N_35696,N_36580);
and U39773 (N_39773,N_35466,N_35270);
xor U39774 (N_39774,N_36769,N_37232);
or U39775 (N_39775,N_35745,N_35535);
and U39776 (N_39776,N_36707,N_36282);
xnor U39777 (N_39777,N_37136,N_36921);
or U39778 (N_39778,N_36837,N_36541);
or U39779 (N_39779,N_35524,N_35434);
and U39780 (N_39780,N_36244,N_35180);
or U39781 (N_39781,N_36215,N_35690);
or U39782 (N_39782,N_35741,N_35149);
nand U39783 (N_39783,N_36810,N_37019);
or U39784 (N_39784,N_36044,N_35728);
or U39785 (N_39785,N_35694,N_35987);
nor U39786 (N_39786,N_36905,N_36164);
nand U39787 (N_39787,N_35698,N_36690);
or U39788 (N_39788,N_35495,N_37210);
nor U39789 (N_39789,N_35028,N_35824);
xor U39790 (N_39790,N_37001,N_35235);
nor U39791 (N_39791,N_36968,N_35185);
and U39792 (N_39792,N_35589,N_36083);
and U39793 (N_39793,N_35549,N_35852);
xnor U39794 (N_39794,N_37217,N_36994);
or U39795 (N_39795,N_36974,N_35300);
or U39796 (N_39796,N_35237,N_35656);
nor U39797 (N_39797,N_36652,N_36029);
nand U39798 (N_39798,N_35756,N_35623);
nor U39799 (N_39799,N_37258,N_35277);
xnor U39800 (N_39800,N_37052,N_36126);
and U39801 (N_39801,N_37083,N_35884);
nor U39802 (N_39802,N_35948,N_36845);
nand U39803 (N_39803,N_35658,N_36858);
and U39804 (N_39804,N_37097,N_36066);
or U39805 (N_39805,N_37481,N_36250);
and U39806 (N_39806,N_36800,N_37450);
nor U39807 (N_39807,N_36582,N_35298);
and U39808 (N_39808,N_36461,N_36764);
nor U39809 (N_39809,N_35726,N_37202);
or U39810 (N_39810,N_35900,N_35605);
and U39811 (N_39811,N_36353,N_35681);
and U39812 (N_39812,N_36481,N_35985);
nand U39813 (N_39813,N_37345,N_35216);
nor U39814 (N_39814,N_35894,N_35826);
nor U39815 (N_39815,N_37328,N_36551);
nand U39816 (N_39816,N_35867,N_35417);
or U39817 (N_39817,N_37102,N_37192);
nand U39818 (N_39818,N_35621,N_36531);
nor U39819 (N_39819,N_37085,N_36847);
and U39820 (N_39820,N_35693,N_36290);
nor U39821 (N_39821,N_36984,N_37395);
nand U39822 (N_39822,N_36954,N_37176);
nand U39823 (N_39823,N_36836,N_35844);
xnor U39824 (N_39824,N_36043,N_36640);
or U39825 (N_39825,N_35134,N_37334);
or U39826 (N_39826,N_35966,N_35575);
nand U39827 (N_39827,N_36104,N_36409);
or U39828 (N_39828,N_35005,N_37302);
nor U39829 (N_39829,N_35049,N_35713);
nor U39830 (N_39830,N_36361,N_36727);
nor U39831 (N_39831,N_37381,N_36446);
nand U39832 (N_39832,N_35884,N_36464);
or U39833 (N_39833,N_37063,N_36247);
or U39834 (N_39834,N_35341,N_37050);
and U39835 (N_39835,N_35190,N_36873);
nand U39836 (N_39836,N_35232,N_36380);
nor U39837 (N_39837,N_37321,N_35366);
xnor U39838 (N_39838,N_36794,N_35985);
nand U39839 (N_39839,N_36990,N_37245);
or U39840 (N_39840,N_35433,N_37320);
nor U39841 (N_39841,N_35832,N_35630);
nand U39842 (N_39842,N_36967,N_35081);
nor U39843 (N_39843,N_35012,N_36065);
nand U39844 (N_39844,N_37482,N_36596);
nor U39845 (N_39845,N_36249,N_37234);
nor U39846 (N_39846,N_37495,N_36167);
nand U39847 (N_39847,N_36726,N_36655);
and U39848 (N_39848,N_36490,N_35285);
and U39849 (N_39849,N_37448,N_35185);
nand U39850 (N_39850,N_35118,N_35498);
nor U39851 (N_39851,N_36063,N_36966);
or U39852 (N_39852,N_36562,N_35707);
and U39853 (N_39853,N_37217,N_36872);
or U39854 (N_39854,N_35939,N_37004);
xor U39855 (N_39855,N_35719,N_35190);
or U39856 (N_39856,N_36311,N_35457);
nand U39857 (N_39857,N_36371,N_37302);
nor U39858 (N_39858,N_36684,N_35121);
and U39859 (N_39859,N_35455,N_36457);
or U39860 (N_39860,N_35251,N_35258);
nand U39861 (N_39861,N_35319,N_35333);
nor U39862 (N_39862,N_36035,N_36672);
or U39863 (N_39863,N_36882,N_36042);
and U39864 (N_39864,N_35364,N_37015);
nand U39865 (N_39865,N_36913,N_37368);
or U39866 (N_39866,N_35806,N_36140);
and U39867 (N_39867,N_35335,N_36630);
or U39868 (N_39868,N_36646,N_37037);
nor U39869 (N_39869,N_35771,N_37254);
xnor U39870 (N_39870,N_35757,N_35188);
xnor U39871 (N_39871,N_35993,N_36364);
nor U39872 (N_39872,N_35707,N_36130);
or U39873 (N_39873,N_36905,N_37190);
nand U39874 (N_39874,N_35821,N_35324);
or U39875 (N_39875,N_36244,N_36859);
nor U39876 (N_39876,N_35498,N_35723);
or U39877 (N_39877,N_36313,N_35611);
xor U39878 (N_39878,N_35734,N_36711);
xor U39879 (N_39879,N_36988,N_37324);
nor U39880 (N_39880,N_37022,N_36980);
and U39881 (N_39881,N_36512,N_35069);
or U39882 (N_39882,N_36889,N_37002);
nor U39883 (N_39883,N_35140,N_35084);
nand U39884 (N_39884,N_35394,N_35735);
and U39885 (N_39885,N_35627,N_36538);
nor U39886 (N_39886,N_36388,N_36363);
xor U39887 (N_39887,N_35509,N_35174);
and U39888 (N_39888,N_36294,N_36793);
and U39889 (N_39889,N_36056,N_35967);
nand U39890 (N_39890,N_37236,N_36870);
and U39891 (N_39891,N_35986,N_35412);
or U39892 (N_39892,N_36572,N_37170);
and U39893 (N_39893,N_35367,N_36532);
xor U39894 (N_39894,N_37095,N_37047);
nor U39895 (N_39895,N_35972,N_37266);
or U39896 (N_39896,N_36662,N_37169);
and U39897 (N_39897,N_36843,N_37209);
nor U39898 (N_39898,N_36627,N_37497);
or U39899 (N_39899,N_35169,N_35363);
nand U39900 (N_39900,N_35464,N_36565);
xnor U39901 (N_39901,N_35140,N_36968);
or U39902 (N_39902,N_35866,N_35438);
nor U39903 (N_39903,N_36730,N_35393);
or U39904 (N_39904,N_36488,N_36310);
nand U39905 (N_39905,N_35570,N_36426);
nand U39906 (N_39906,N_36932,N_35373);
or U39907 (N_39907,N_36492,N_35405);
or U39908 (N_39908,N_36470,N_35160);
or U39909 (N_39909,N_35302,N_35362);
nand U39910 (N_39910,N_35365,N_35061);
or U39911 (N_39911,N_36911,N_36771);
xor U39912 (N_39912,N_36061,N_37241);
or U39913 (N_39913,N_37067,N_35313);
nor U39914 (N_39914,N_37401,N_35028);
or U39915 (N_39915,N_36346,N_37268);
nand U39916 (N_39916,N_36443,N_36511);
xor U39917 (N_39917,N_36643,N_35226);
xor U39918 (N_39918,N_37035,N_36840);
nand U39919 (N_39919,N_35638,N_36369);
and U39920 (N_39920,N_37136,N_36801);
or U39921 (N_39921,N_36854,N_36296);
nor U39922 (N_39922,N_35794,N_35286);
nor U39923 (N_39923,N_36034,N_36249);
xor U39924 (N_39924,N_36165,N_36546);
nand U39925 (N_39925,N_36255,N_36303);
nand U39926 (N_39926,N_36936,N_35443);
or U39927 (N_39927,N_35693,N_35087);
and U39928 (N_39928,N_37412,N_35174);
nand U39929 (N_39929,N_35998,N_36702);
nor U39930 (N_39930,N_35727,N_35521);
nand U39931 (N_39931,N_37318,N_36969);
and U39932 (N_39932,N_36259,N_35428);
or U39933 (N_39933,N_36950,N_35684);
and U39934 (N_39934,N_36887,N_35538);
or U39935 (N_39935,N_35641,N_37016);
and U39936 (N_39936,N_35260,N_36893);
or U39937 (N_39937,N_36710,N_35888);
or U39938 (N_39938,N_36052,N_36116);
nor U39939 (N_39939,N_36809,N_37091);
or U39940 (N_39940,N_35400,N_35477);
or U39941 (N_39941,N_36336,N_36699);
nand U39942 (N_39942,N_35529,N_36814);
nand U39943 (N_39943,N_36805,N_37327);
or U39944 (N_39944,N_35938,N_36945);
nand U39945 (N_39945,N_37359,N_35195);
and U39946 (N_39946,N_37213,N_36003);
nand U39947 (N_39947,N_36848,N_35198);
or U39948 (N_39948,N_35288,N_36943);
or U39949 (N_39949,N_35374,N_36503);
nand U39950 (N_39950,N_36476,N_37160);
and U39951 (N_39951,N_35521,N_37480);
xor U39952 (N_39952,N_35645,N_36422);
nand U39953 (N_39953,N_37189,N_35311);
nor U39954 (N_39954,N_35003,N_37248);
nor U39955 (N_39955,N_35089,N_36844);
nor U39956 (N_39956,N_36451,N_36793);
nor U39957 (N_39957,N_37235,N_36549);
nor U39958 (N_39958,N_36609,N_37127);
and U39959 (N_39959,N_37081,N_37446);
nand U39960 (N_39960,N_35201,N_36055);
nand U39961 (N_39961,N_35019,N_35899);
and U39962 (N_39962,N_35925,N_35034);
nand U39963 (N_39963,N_36373,N_37130);
and U39964 (N_39964,N_36769,N_35328);
nand U39965 (N_39965,N_35749,N_37467);
nor U39966 (N_39966,N_36114,N_35990);
xor U39967 (N_39967,N_35820,N_36300);
or U39968 (N_39968,N_35008,N_36022);
and U39969 (N_39969,N_37447,N_35716);
xor U39970 (N_39970,N_35379,N_37242);
nand U39971 (N_39971,N_36995,N_35106);
or U39972 (N_39972,N_35034,N_35936);
nor U39973 (N_39973,N_36933,N_35855);
nand U39974 (N_39974,N_35540,N_36056);
xor U39975 (N_39975,N_36705,N_36850);
nand U39976 (N_39976,N_37214,N_35164);
nand U39977 (N_39977,N_35342,N_36423);
nor U39978 (N_39978,N_36094,N_37212);
or U39979 (N_39979,N_36369,N_36713);
xor U39980 (N_39980,N_36684,N_37447);
or U39981 (N_39981,N_36121,N_36323);
and U39982 (N_39982,N_36707,N_35106);
nor U39983 (N_39983,N_35007,N_36967);
xor U39984 (N_39984,N_37468,N_35579);
nand U39985 (N_39985,N_35162,N_35328);
nand U39986 (N_39986,N_35784,N_35427);
nand U39987 (N_39987,N_35118,N_35665);
and U39988 (N_39988,N_36182,N_35349);
and U39989 (N_39989,N_36817,N_35397);
nand U39990 (N_39990,N_37064,N_35060);
nor U39991 (N_39991,N_36123,N_36495);
nor U39992 (N_39992,N_35291,N_36658);
nand U39993 (N_39993,N_36973,N_37208);
or U39994 (N_39994,N_36024,N_36619);
nand U39995 (N_39995,N_35675,N_36146);
or U39996 (N_39996,N_37100,N_35031);
nand U39997 (N_39997,N_35311,N_37088);
nor U39998 (N_39998,N_36346,N_35594);
or U39999 (N_39999,N_35460,N_37062);
nor U40000 (N_40000,N_37956,N_39895);
or U40001 (N_40001,N_39301,N_38506);
nand U40002 (N_40002,N_39896,N_38002);
nor U40003 (N_40003,N_38557,N_38594);
and U40004 (N_40004,N_38826,N_39902);
nor U40005 (N_40005,N_37962,N_38700);
and U40006 (N_40006,N_38397,N_39701);
or U40007 (N_40007,N_38796,N_39345);
and U40008 (N_40008,N_37730,N_37992);
and U40009 (N_40009,N_39480,N_38113);
or U40010 (N_40010,N_37586,N_38483);
and U40011 (N_40011,N_38372,N_38346);
nand U40012 (N_40012,N_38989,N_39740);
nor U40013 (N_40013,N_37915,N_38579);
nor U40014 (N_40014,N_39202,N_39767);
nor U40015 (N_40015,N_39922,N_37789);
or U40016 (N_40016,N_37875,N_39222);
xor U40017 (N_40017,N_38086,N_38099);
nand U40018 (N_40018,N_39894,N_38772);
xnor U40019 (N_40019,N_39138,N_39231);
or U40020 (N_40020,N_38469,N_39288);
or U40021 (N_40021,N_39623,N_38495);
nand U40022 (N_40022,N_39968,N_38556);
and U40023 (N_40023,N_39314,N_39860);
or U40024 (N_40024,N_38341,N_38786);
and U40025 (N_40025,N_38932,N_38761);
nor U40026 (N_40026,N_39120,N_38953);
nand U40027 (N_40027,N_38755,N_38164);
or U40028 (N_40028,N_39006,N_38137);
or U40029 (N_40029,N_38101,N_39203);
nand U40030 (N_40030,N_39065,N_38603);
and U40031 (N_40031,N_38351,N_39640);
nand U40032 (N_40032,N_39209,N_38795);
nand U40033 (N_40033,N_39557,N_39353);
nand U40034 (N_40034,N_37859,N_38733);
nand U40035 (N_40035,N_38889,N_37712);
nor U40036 (N_40036,N_39863,N_38694);
and U40037 (N_40037,N_39490,N_38870);
nor U40038 (N_40038,N_39693,N_39530);
xnor U40039 (N_40039,N_37762,N_38460);
and U40040 (N_40040,N_38585,N_39181);
nand U40041 (N_40041,N_39672,N_38709);
and U40042 (N_40042,N_39880,N_39634);
or U40043 (N_40043,N_38388,N_38160);
nor U40044 (N_40044,N_38981,N_38587);
or U40045 (N_40045,N_38611,N_38187);
nand U40046 (N_40046,N_37944,N_39768);
or U40047 (N_40047,N_38443,N_39395);
nand U40048 (N_40048,N_38055,N_39245);
or U40049 (N_40049,N_39264,N_39846);
nand U40050 (N_40050,N_38540,N_38052);
xnor U40051 (N_40051,N_39391,N_39952);
or U40052 (N_40052,N_39124,N_39756);
or U40053 (N_40053,N_37951,N_39185);
nand U40054 (N_40054,N_38633,N_38444);
nand U40055 (N_40055,N_37668,N_38474);
and U40056 (N_40056,N_38103,N_38883);
nand U40057 (N_40057,N_39333,N_38714);
nor U40058 (N_40058,N_38596,N_38007);
nand U40059 (N_40059,N_38161,N_38138);
xnor U40060 (N_40060,N_37908,N_39268);
nand U40061 (N_40061,N_38194,N_38781);
nor U40062 (N_40062,N_37925,N_38866);
or U40063 (N_40063,N_37632,N_39698);
and U40064 (N_40064,N_38163,N_39485);
and U40065 (N_40065,N_37919,N_37893);
and U40066 (N_40066,N_37701,N_38401);
and U40067 (N_40067,N_38182,N_39388);
and U40068 (N_40068,N_38285,N_39051);
nand U40069 (N_40069,N_38745,N_37512);
and U40070 (N_40070,N_38806,N_38575);
and U40071 (N_40071,N_38931,N_39054);
and U40072 (N_40072,N_38299,N_39095);
or U40073 (N_40073,N_39063,N_38679);
nor U40074 (N_40074,N_37613,N_38669);
xnor U40075 (N_40075,N_37887,N_38956);
nand U40076 (N_40076,N_38522,N_38353);
xor U40077 (N_40077,N_37818,N_39446);
or U40078 (N_40078,N_38368,N_37928);
nor U40079 (N_40079,N_38266,N_38711);
nand U40080 (N_40080,N_38038,N_38527);
or U40081 (N_40081,N_39025,N_38671);
and U40082 (N_40082,N_38841,N_38542);
and U40083 (N_40083,N_38899,N_38442);
and U40084 (N_40084,N_39630,N_38090);
nor U40085 (N_40085,N_38972,N_39217);
or U40086 (N_40086,N_38604,N_39532);
xnor U40087 (N_40087,N_39201,N_39189);
nand U40088 (N_40088,N_38861,N_39722);
nor U40089 (N_40089,N_39242,N_39744);
and U40090 (N_40090,N_39319,N_38012);
or U40091 (N_40091,N_38272,N_39663);
or U40092 (N_40092,N_37916,N_37914);
nor U40093 (N_40093,N_39022,N_37719);
nand U40094 (N_40094,N_37782,N_39118);
or U40095 (N_40095,N_38457,N_39577);
nor U40096 (N_40096,N_37764,N_38533);
and U40097 (N_40097,N_37548,N_39590);
nor U40098 (N_40098,N_39210,N_39008);
or U40099 (N_40099,N_39145,N_38509);
nor U40100 (N_40100,N_39158,N_38015);
nor U40101 (N_40101,N_37587,N_39448);
nand U40102 (N_40102,N_37982,N_39949);
or U40103 (N_40103,N_39820,N_39782);
and U40104 (N_40104,N_37553,N_38453);
or U40105 (N_40105,N_38552,N_38029);
nor U40106 (N_40106,N_37999,N_38241);
or U40107 (N_40107,N_38063,N_38074);
nor U40108 (N_40108,N_39257,N_39838);
or U40109 (N_40109,N_39766,N_39654);
or U40110 (N_40110,N_37513,N_38140);
and U40111 (N_40111,N_39481,N_38627);
nor U40112 (N_40112,N_38348,N_38327);
nor U40113 (N_40113,N_38917,N_37829);
or U40114 (N_40114,N_38115,N_39092);
or U40115 (N_40115,N_37502,N_39169);
or U40116 (N_40116,N_38643,N_38863);
nand U40117 (N_40117,N_38938,N_39538);
nor U40118 (N_40118,N_38884,N_39897);
nor U40119 (N_40119,N_38454,N_39427);
nand U40120 (N_40120,N_37593,N_39605);
and U40121 (N_40121,N_39487,N_38895);
or U40122 (N_40122,N_38554,N_37960);
and U40123 (N_40123,N_38234,N_39582);
and U40124 (N_40124,N_39888,N_37966);
or U40125 (N_40125,N_38614,N_38652);
nand U40126 (N_40126,N_39364,N_37742);
or U40127 (N_40127,N_39821,N_37710);
or U40128 (N_40128,N_39339,N_39347);
and U40129 (N_40129,N_39650,N_38721);
or U40130 (N_40130,N_39521,N_38856);
nand U40131 (N_40131,N_39381,N_38133);
nand U40132 (N_40132,N_38854,N_39493);
nor U40133 (N_40133,N_39526,N_38110);
nor U40134 (N_40134,N_38868,N_38355);
nor U40135 (N_40135,N_39597,N_37833);
or U40136 (N_40136,N_38945,N_38468);
or U40137 (N_40137,N_39901,N_38130);
or U40138 (N_40138,N_38816,N_38690);
nor U40139 (N_40139,N_38770,N_38239);
xor U40140 (N_40140,N_37964,N_37890);
nor U40141 (N_40141,N_38172,N_38405);
nand U40142 (N_40142,N_37516,N_38612);
xor U40143 (N_40143,N_38188,N_38011);
or U40144 (N_40144,N_39932,N_37901);
xor U40145 (N_40145,N_38216,N_38717);
and U40146 (N_40146,N_39466,N_39007);
and U40147 (N_40147,N_38463,N_37766);
nand U40148 (N_40148,N_37631,N_38821);
or U40149 (N_40149,N_39473,N_37723);
nand U40150 (N_40150,N_38311,N_37942);
nand U40151 (N_40151,N_38879,N_39101);
xor U40152 (N_40152,N_39954,N_39678);
and U40153 (N_40153,N_39598,N_38148);
nand U40154 (N_40154,N_38389,N_38410);
or U40155 (N_40155,N_39046,N_39369);
and U40156 (N_40156,N_38283,N_38996);
or U40157 (N_40157,N_37564,N_39967);
nor U40158 (N_40158,N_38267,N_37791);
nor U40159 (N_40159,N_38065,N_39130);
and U40160 (N_40160,N_37788,N_39852);
nand U40161 (N_40161,N_39772,N_38901);
and U40162 (N_40162,N_38536,N_37753);
and U40163 (N_40163,N_39278,N_37538);
xor U40164 (N_40164,N_39104,N_39689);
and U40165 (N_40165,N_38087,N_39495);
nor U40166 (N_40166,N_39749,N_38304);
and U40167 (N_40167,N_38365,N_39992);
nand U40168 (N_40168,N_37577,N_38935);
or U40169 (N_40169,N_37589,N_39251);
nand U40170 (N_40170,N_39424,N_39648);
nand U40171 (N_40171,N_38277,N_39260);
nor U40172 (N_40172,N_39851,N_38149);
nor U40173 (N_40173,N_38387,N_39213);
or U40174 (N_40174,N_37612,N_39153);
nand U40175 (N_40175,N_38192,N_37660);
nor U40176 (N_40176,N_38791,N_39947);
or U40177 (N_40177,N_39474,N_39784);
or U40178 (N_40178,N_39580,N_39686);
xnor U40179 (N_40179,N_39175,N_38104);
nand U40180 (N_40180,N_38108,N_39951);
or U40181 (N_40181,N_38114,N_38619);
or U40182 (N_40182,N_38217,N_38222);
nand U40183 (N_40183,N_37824,N_39700);
xor U40184 (N_40184,N_38549,N_37812);
nor U40185 (N_40185,N_38003,N_37955);
nor U40186 (N_40186,N_39087,N_39218);
nand U40187 (N_40187,N_38497,N_39310);
or U40188 (N_40188,N_39108,N_39613);
nand U40189 (N_40189,N_39277,N_39933);
nand U40190 (N_40190,N_38815,N_39057);
nand U40191 (N_40191,N_39725,N_38697);
nand U40192 (N_40192,N_37504,N_38338);
nand U40193 (N_40193,N_37580,N_37559);
nand U40194 (N_40194,N_38837,N_39115);
and U40195 (N_40195,N_38275,N_38263);
or U40196 (N_40196,N_38922,N_37590);
nor U40197 (N_40197,N_37997,N_38936);
xnor U40198 (N_40198,N_38202,N_39511);
nand U40199 (N_40199,N_38865,N_39862);
and U40200 (N_40200,N_37821,N_38912);
nor U40201 (N_40201,N_38246,N_37633);
or U40202 (N_40202,N_37813,N_37920);
and U40203 (N_40203,N_39979,N_39870);
nand U40204 (N_40204,N_39680,N_39363);
nor U40205 (N_40205,N_38950,N_39997);
nand U40206 (N_40206,N_38551,N_39279);
nand U40207 (N_40207,N_38918,N_39872);
and U40208 (N_40208,N_38077,N_38805);
nand U40209 (N_40209,N_39077,N_37615);
nor U40210 (N_40210,N_38257,N_37662);
and U40211 (N_40211,N_39981,N_39252);
nor U40212 (N_40212,N_38985,N_39632);
nand U40213 (N_40213,N_39091,N_39034);
or U40214 (N_40214,N_39618,N_39114);
or U40215 (N_40215,N_38990,N_39327);
nor U40216 (N_40216,N_39033,N_39716);
or U40217 (N_40217,N_39738,N_38336);
or U40218 (N_40218,N_39386,N_37834);
xor U40219 (N_40219,N_38544,N_38919);
nor U40220 (N_40220,N_39940,N_39522);
nand U40221 (N_40221,N_38465,N_39558);
nand U40222 (N_40222,N_39584,N_37672);
and U40223 (N_40223,N_39696,N_38136);
nand U40224 (N_40224,N_38330,N_38846);
nor U40225 (N_40225,N_38787,N_38375);
and U40226 (N_40226,N_37971,N_39450);
nor U40227 (N_40227,N_39874,N_38672);
xor U40228 (N_40228,N_38485,N_38450);
or U40229 (N_40229,N_37679,N_39697);
nor U40230 (N_40230,N_39750,N_37871);
and U40231 (N_40231,N_39343,N_39233);
xor U40232 (N_40232,N_39800,N_37784);
nand U40233 (N_40233,N_38827,N_37697);
nor U40234 (N_40234,N_39163,N_38976);
nand U40235 (N_40235,N_39426,N_38345);
nor U40236 (N_40236,N_39876,N_38850);
xnor U40237 (N_40237,N_38606,N_39732);
xor U40238 (N_40238,N_39866,N_39362);
nand U40239 (N_40239,N_39005,N_38794);
nor U40240 (N_40240,N_37894,N_39069);
or U40241 (N_40241,N_39107,N_39170);
or U40242 (N_40242,N_39298,N_38303);
nor U40243 (N_40243,N_37692,N_38414);
and U40244 (N_40244,N_37555,N_38929);
or U40245 (N_40245,N_38916,N_39512);
and U40246 (N_40246,N_39293,N_39224);
nand U40247 (N_40247,N_38005,N_39453);
or U40248 (N_40248,N_37994,N_37560);
nor U40249 (N_40249,N_39633,N_39556);
nand U40250 (N_40250,N_38988,N_37627);
and U40251 (N_40251,N_39796,N_38296);
or U40252 (N_40252,N_38333,N_39015);
nand U40253 (N_40253,N_39075,N_39788);
nor U40254 (N_40254,N_39188,N_38008);
or U40255 (N_40255,N_39308,N_39271);
and U40256 (N_40256,N_39569,N_38888);
nor U40257 (N_40257,N_37873,N_39320);
and U40258 (N_40258,N_37600,N_38281);
nor U40259 (N_40259,N_38235,N_38419);
nand U40260 (N_40260,N_38894,N_37809);
and U40261 (N_40261,N_38847,N_38204);
nor U40262 (N_40262,N_38574,N_38572);
nand U40263 (N_40263,N_39593,N_38091);
nor U40264 (N_40264,N_39085,N_39999);
and U40265 (N_40265,N_39823,N_39978);
nand U40266 (N_40266,N_39976,N_39019);
xnor U40267 (N_40267,N_38181,N_38037);
or U40268 (N_40268,N_39083,N_38395);
and U40269 (N_40269,N_37953,N_39705);
nor U40270 (N_40270,N_39411,N_38605);
and U40271 (N_40271,N_38725,N_39884);
and U40272 (N_40272,N_37807,N_38384);
nand U40273 (N_40273,N_39950,N_37670);
nor U40274 (N_40274,N_39326,N_39229);
nand U40275 (N_40275,N_37588,N_37838);
nand U40276 (N_40276,N_38840,N_38920);
nand U40277 (N_40277,N_39877,N_39144);
or U40278 (N_40278,N_37611,N_37978);
xor U40279 (N_40279,N_37886,N_39196);
or U40280 (N_40280,N_39387,N_37514);
or U40281 (N_40281,N_39379,N_38186);
nor U40282 (N_40282,N_39977,N_38957);
nor U40283 (N_40283,N_38313,N_39548);
or U40284 (N_40284,N_37624,N_37808);
nand U40285 (N_40285,N_38155,N_39183);
nor U40286 (N_40286,N_37572,N_39709);
nor U40287 (N_40287,N_39449,N_39676);
nor U40288 (N_40288,N_39515,N_38366);
xor U40289 (N_40289,N_39325,N_38939);
nand U40290 (N_40290,N_37666,N_39093);
and U40291 (N_40291,N_38265,N_39361);
or U40292 (N_40292,N_39125,N_38417);
nor U40293 (N_40293,N_37847,N_37836);
xnor U40294 (N_40294,N_39960,N_38060);
nor U40295 (N_40295,N_37803,N_37635);
nand U40296 (N_40296,N_38952,N_39758);
nand U40297 (N_40297,N_38196,N_37987);
nand U40298 (N_40298,N_38637,N_39032);
nor U40299 (N_40299,N_39935,N_39719);
and U40300 (N_40300,N_38766,N_39924);
or U40301 (N_40301,N_37864,N_38399);
xnor U40302 (N_40302,N_38739,N_37760);
xnor U40303 (N_40303,N_38158,N_38441);
nand U40304 (N_40304,N_39399,N_39499);
nor U40305 (N_40305,N_38774,N_39404);
xor U40306 (N_40306,N_39525,N_37896);
nand U40307 (N_40307,N_37734,N_38802);
and U40308 (N_40308,N_39273,N_37831);
nand U40309 (N_40309,N_37661,N_38185);
and U40310 (N_40310,N_38666,N_37769);
nor U40311 (N_40311,N_39771,N_38479);
or U40312 (N_40312,N_39988,N_38340);
or U40313 (N_40313,N_38504,N_39024);
nor U40314 (N_40314,N_38686,N_37550);
nor U40315 (N_40315,N_38129,N_39292);
and U40316 (N_40316,N_39604,N_39524);
and U40317 (N_40317,N_39462,N_38501);
or U40318 (N_40318,N_37932,N_39142);
and U40319 (N_40319,N_38783,N_38408);
xnor U40320 (N_40320,N_38193,N_39708);
nor U40321 (N_40321,N_39778,N_38224);
xnor U40322 (N_40322,N_38043,N_39916);
nand U40323 (N_40323,N_38391,N_39047);
nor U40324 (N_40324,N_38321,N_39906);
nor U40325 (N_40325,N_39113,N_39969);
nand U40326 (N_40326,N_38219,N_38705);
or U40327 (N_40327,N_37592,N_39566);
or U40328 (N_40328,N_38083,N_38740);
or U40329 (N_40329,N_38323,N_37839);
or U40330 (N_40330,N_39467,N_37853);
xor U40331 (N_40331,N_37601,N_38560);
or U40332 (N_40332,N_39066,N_39418);
nor U40333 (N_40333,N_39122,N_39927);
or U40334 (N_40334,N_38558,N_39405);
or U40335 (N_40335,N_39998,N_37866);
nand U40336 (N_40336,N_39579,N_38287);
nor U40337 (N_40337,N_38251,N_38570);
xnor U40338 (N_40338,N_38685,N_38021);
nor U40339 (N_40339,N_38962,N_37594);
nand U40340 (N_40340,N_37968,N_39636);
and U40341 (N_40341,N_37582,N_38492);
nor U40342 (N_40342,N_39211,N_38206);
nor U40343 (N_40343,N_37775,N_37822);
and U40344 (N_40344,N_39543,N_37961);
or U40345 (N_40345,N_39148,N_39176);
and U40346 (N_40346,N_39615,N_38951);
nand U40347 (N_40347,N_37558,N_38117);
or U40348 (N_40348,N_38280,N_39811);
or U40349 (N_40349,N_39563,N_39889);
or U40350 (N_40350,N_38660,N_37904);
nor U40351 (N_40351,N_38406,N_39822);
or U40352 (N_40352,N_39416,N_39394);
and U40353 (N_40353,N_37659,N_39482);
and U40354 (N_40354,N_38902,N_37581);
nor U40355 (N_40355,N_39309,N_38017);
xor U40356 (N_40356,N_38869,N_37909);
xor U40357 (N_40357,N_37563,N_39322);
xnor U40358 (N_40358,N_38238,N_38201);
nand U40359 (N_40359,N_39174,N_38653);
or U40360 (N_40360,N_38632,N_37981);
nor U40361 (N_40361,N_37616,N_39751);
nand U40362 (N_40362,N_39535,N_39344);
nor U40363 (N_40363,N_39859,N_37561);
or U40364 (N_40364,N_38053,N_37811);
nor U40365 (N_40365,N_38526,N_38462);
or U40366 (N_40366,N_37715,N_38743);
or U40367 (N_40367,N_39845,N_38750);
or U40368 (N_40368,N_38018,N_38394);
and U40369 (N_40369,N_39652,N_38242);
or U40370 (N_40370,N_38514,N_38098);
nand U40371 (N_40371,N_38607,N_39706);
and U40372 (N_40372,N_38066,N_39139);
nand U40373 (N_40373,N_37943,N_39420);
or U40374 (N_40374,N_37696,N_39841);
xnor U40375 (N_40375,N_37658,N_38663);
nand U40376 (N_40376,N_39626,N_39374);
or U40377 (N_40377,N_37669,N_37820);
nor U40378 (N_40378,N_38374,N_39471);
and U40379 (N_40379,N_37923,N_39759);
nor U40380 (N_40380,N_37722,N_39727);
nor U40381 (N_40381,N_38314,N_39223);
or U40382 (N_40382,N_39549,N_39690);
nand U40383 (N_40383,N_38432,N_38064);
nand U40384 (N_40384,N_39945,N_38830);
nor U40385 (N_40385,N_37653,N_38857);
or U40386 (N_40386,N_38300,N_37880);
nand U40387 (N_40387,N_37801,N_37556);
and U40388 (N_40388,N_38620,N_39429);
nand U40389 (N_40389,N_38464,N_39494);
nand U40390 (N_40390,N_37619,N_39850);
and U40391 (N_40391,N_38214,N_39097);
or U40392 (N_40392,N_39507,N_39944);
nor U40393 (N_40393,N_39925,N_38523);
and U40394 (N_40394,N_38120,N_38648);
nor U40395 (N_40395,N_39397,N_39655);
nor U40396 (N_40396,N_39814,N_39358);
nor U40397 (N_40397,N_39128,N_39258);
or U40398 (N_40398,N_39567,N_37584);
or U40399 (N_40399,N_38730,N_39990);
nor U40400 (N_40400,N_39801,N_38439);
nand U40401 (N_40401,N_38531,N_39710);
xnor U40402 (N_40402,N_38264,N_38398);
and U40403 (N_40403,N_37657,N_37902);
xnor U40404 (N_40404,N_38072,N_38412);
and U40405 (N_40405,N_38131,N_39109);
nand U40406 (N_40406,N_37937,N_37900);
nor U40407 (N_40407,N_37605,N_39624);
xnor U40408 (N_40408,N_37950,N_39785);
and U40409 (N_40409,N_39383,N_38236);
nor U40410 (N_40410,N_39178,N_38487);
nand U40411 (N_40411,N_39736,N_39980);
nand U40412 (N_40412,N_39237,N_38698);
nor U40413 (N_40413,N_39100,N_38667);
or U40414 (N_40414,N_39581,N_39956);
and U40415 (N_40415,N_39376,N_38954);
and U40416 (N_40416,N_39608,N_38789);
xor U40417 (N_40417,N_38094,N_39043);
nor U40418 (N_40418,N_38416,N_38864);
nand U40419 (N_40419,N_38093,N_38143);
nor U40420 (N_40420,N_39625,N_39475);
or U40421 (N_40421,N_39910,N_39645);
and U40422 (N_40422,N_39127,N_39117);
nand U40423 (N_40423,N_39050,N_38760);
nand U40424 (N_40424,N_39657,N_38418);
or U40425 (N_40425,N_37609,N_38547);
nor U40426 (N_40426,N_38971,N_39282);
nand U40427 (N_40427,N_37816,N_39986);
and U40428 (N_40428,N_39937,N_39040);
and U40429 (N_40429,N_37979,N_39832);
xnor U40430 (N_40430,N_39726,N_38023);
nand U40431 (N_40431,N_38179,N_38727);
xnor U40432 (N_40432,N_39436,N_38986);
and U40433 (N_40433,N_39461,N_37733);
nor U40434 (N_40434,N_38765,N_38415);
and U40435 (N_40435,N_39519,N_39098);
nand U40436 (N_40436,N_38290,N_38595);
and U40437 (N_40437,N_37963,N_39221);
or U40438 (N_40438,N_39409,N_38817);
xor U40439 (N_40439,N_38413,N_38767);
and U40440 (N_40440,N_38590,N_39419);
or U40441 (N_40441,N_39915,N_39489);
nor U40442 (N_40442,N_38424,N_38360);
xnor U40443 (N_40443,N_38363,N_39247);
nor U40444 (N_40444,N_38438,N_39812);
nor U40445 (N_40445,N_38058,N_38780);
nand U40446 (N_40446,N_39509,N_38364);
nand U40447 (N_40447,N_38658,N_38451);
or U40448 (N_40448,N_39594,N_38695);
nor U40449 (N_40449,N_38613,N_39267);
nor U40450 (N_40450,N_39417,N_39235);
or U40451 (N_40451,N_38146,N_38508);
nand U40452 (N_40452,N_38703,N_37684);
nand U40453 (N_40453,N_38107,N_39350);
nor U40454 (N_40454,N_39060,N_39468);
xnor U40455 (N_40455,N_38831,N_38031);
nor U40456 (N_40456,N_37537,N_38890);
and U40457 (N_40457,N_38215,N_39226);
or U40458 (N_40458,N_38493,N_39248);
nand U40459 (N_40459,N_39488,N_39774);
nand U40460 (N_40460,N_39703,N_39317);
or U40461 (N_40461,N_37711,N_39938);
nor U40462 (N_40462,N_38842,N_39337);
nand U40463 (N_40463,N_39704,N_38271);
and U40464 (N_40464,N_38403,N_37664);
nand U40465 (N_40465,N_39370,N_39849);
nor U40466 (N_40466,N_39677,N_38472);
and U40467 (N_40467,N_38307,N_37667);
and U40468 (N_40468,N_37656,N_39441);
and U40469 (N_40469,N_38639,N_39776);
xnor U40470 (N_40470,N_38838,N_39711);
nand U40471 (N_40471,N_38390,N_39638);
or U40472 (N_40472,N_39079,N_39836);
xor U40473 (N_40473,N_39664,N_37704);
xor U40474 (N_40474,N_38045,N_39017);
nand U40475 (N_40475,N_37645,N_39962);
nand U40476 (N_40476,N_38473,N_38231);
and U40477 (N_40477,N_38250,N_37617);
or U40478 (N_40478,N_39666,N_38886);
or U40479 (N_40479,N_39354,N_37526);
xnor U40480 (N_40480,N_38975,N_38615);
nand U40481 (N_40481,N_38402,N_39452);
or U40482 (N_40482,N_39219,N_38984);
nand U40483 (N_40483,N_39428,N_37708);
and U40484 (N_40484,N_39000,N_38171);
or U40485 (N_40485,N_38726,N_39564);
nor U40486 (N_40486,N_39854,N_39537);
and U40487 (N_40487,N_37621,N_37549);
nand U40488 (N_40488,N_39742,N_38256);
nand U40489 (N_40489,N_37874,N_38423);
nand U40490 (N_40490,N_38199,N_38189);
or U40491 (N_40491,N_39160,N_38813);
or U40492 (N_40492,N_38226,N_39911);
nor U40493 (N_40493,N_38411,N_39790);
and U40494 (N_40494,N_37620,N_37910);
nor U40495 (N_40495,N_38778,N_37597);
and U40496 (N_40496,N_38371,N_38124);
nor U40497 (N_40497,N_37647,N_37576);
or U40498 (N_40498,N_38435,N_39105);
or U40499 (N_40499,N_37879,N_38383);
and U40500 (N_40500,N_39958,N_37706);
or U40501 (N_40501,N_38538,N_37828);
nor U40502 (N_40502,N_37799,N_39627);
or U40503 (N_40503,N_39439,N_37878);
or U40504 (N_40504,N_38812,N_39541);
nor U40505 (N_40505,N_39018,N_37773);
nor U40506 (N_40506,N_38208,N_38834);
nand U40507 (N_40507,N_37678,N_38753);
or U40508 (N_40508,N_39975,N_38254);
nor U40509 (N_40509,N_38561,N_39794);
or U40510 (N_40510,N_39194,N_39064);
nor U40511 (N_40511,N_39250,N_39243);
and U40512 (N_40512,N_39255,N_38312);
or U40513 (N_40513,N_37721,N_38845);
xnor U40514 (N_40514,N_39658,N_37767);
xnor U40515 (N_40515,N_39819,N_39856);
nor U40516 (N_40516,N_39674,N_39121);
and U40517 (N_40517,N_37726,N_38481);
nand U40518 (N_40518,N_37651,N_37636);
nor U40519 (N_40519,N_38820,N_37855);
nand U40520 (N_40520,N_38079,N_38262);
or U40521 (N_40521,N_39035,N_37930);
and U40522 (N_40522,N_37650,N_37736);
or U40523 (N_40523,N_38502,N_39614);
nand U40524 (N_40524,N_39571,N_39116);
and U40525 (N_40525,N_37709,N_38335);
and U40526 (N_40526,N_39484,N_39763);
xor U40527 (N_40527,N_38764,N_39656);
or U40528 (N_40528,N_37535,N_37517);
xor U40529 (N_40529,N_37644,N_37969);
nor U40530 (N_40530,N_39002,N_38218);
or U40531 (N_40531,N_37872,N_39926);
nand U40532 (N_40532,N_39197,N_37825);
or U40533 (N_40533,N_37970,N_39622);
nor U40534 (N_40534,N_38370,N_37503);
nand U40535 (N_40535,N_37935,N_38728);
and U40536 (N_40536,N_38004,N_38240);
nand U40537 (N_40537,N_38793,N_39132);
and U40538 (N_40538,N_37506,N_38881);
xor U40539 (N_40539,N_39883,N_39306);
nand U40540 (N_40540,N_39454,N_38926);
xnor U40541 (N_40541,N_39792,N_39575);
nand U40542 (N_40542,N_39225,N_39067);
nor U40543 (N_40543,N_39817,N_39510);
nand U40544 (N_40544,N_39366,N_39498);
xor U40545 (N_40545,N_38081,N_37705);
and U40546 (N_40546,N_38969,N_37856);
or U40547 (N_40547,N_37881,N_38127);
nand U40548 (N_40548,N_38059,N_39205);
and U40549 (N_40549,N_39283,N_39966);
and U40550 (N_40550,N_39336,N_38157);
or U40551 (N_40551,N_38689,N_38887);
and U40552 (N_40552,N_37727,N_38773);
and U40553 (N_40553,N_37796,N_38436);
xnor U40554 (N_40554,N_39562,N_38085);
and U40555 (N_40555,N_39761,N_39234);
or U40556 (N_40556,N_38213,N_37921);
nor U40557 (N_40557,N_38792,N_38741);
and U40558 (N_40558,N_38563,N_39440);
or U40559 (N_40559,N_37749,N_38109);
nor U40560 (N_40560,N_37747,N_39269);
nor U40561 (N_40561,N_39644,N_39029);
or U40562 (N_40562,N_38471,N_38392);
nand U40563 (N_40563,N_38162,N_39547);
or U40564 (N_40564,N_37954,N_38618);
and U40565 (N_40565,N_38332,N_37870);
nor U40566 (N_40566,N_37988,N_39013);
nor U40567 (N_40567,N_38580,N_37862);
nor U40568 (N_40568,N_38476,N_38835);
or U40569 (N_40569,N_37683,N_37579);
nand U40570 (N_40570,N_39550,N_39119);
and U40571 (N_40571,N_39016,N_38828);
nor U40572 (N_40572,N_39081,N_39500);
nand U40573 (N_40573,N_39021,N_38376);
or U40574 (N_40574,N_39639,N_37913);
or U40575 (N_40575,N_39177,N_38798);
and U40576 (N_40576,N_38165,N_38532);
nand U40577 (N_40577,N_37750,N_37628);
or U40578 (N_40578,N_37817,N_38804);
nor U40579 (N_40579,N_39036,N_39232);
or U40580 (N_40580,N_38480,N_39825);
or U40581 (N_40581,N_39685,N_39718);
or U40582 (N_40582,N_38511,N_37739);
xnor U40583 (N_40583,N_38046,N_39671);
nand U40584 (N_40584,N_38858,N_37665);
or U40585 (N_40585,N_39919,N_39037);
and U40586 (N_40586,N_39042,N_39837);
nand U40587 (N_40587,N_38974,N_39406);
nor U40588 (N_40588,N_39545,N_38422);
and U40589 (N_40589,N_38983,N_38958);
nand U40590 (N_40590,N_38317,N_39787);
or U40591 (N_40591,N_38822,N_38499);
or U40592 (N_40592,N_39433,N_39606);
and U40593 (N_40593,N_39457,N_38891);
xor U40594 (N_40594,N_39472,N_38748);
or U40595 (N_40595,N_37985,N_38684);
nor U40596 (N_40596,N_39078,N_38539);
or U40597 (N_40597,N_38885,N_39014);
and U40598 (N_40598,N_37793,N_37680);
nand U40599 (N_40599,N_39246,N_39010);
or U40600 (N_40600,N_37984,N_39723);
or U40601 (N_40601,N_38910,N_37540);
nor U40602 (N_40602,N_39199,N_39533);
nand U40603 (N_40603,N_37759,N_38132);
xnor U40604 (N_40604,N_39503,N_38738);
and U40605 (N_40605,N_37755,N_39241);
nor U40606 (N_40606,N_39403,N_39307);
nor U40607 (N_40607,N_38030,N_39076);
nand U40608 (N_40608,N_37850,N_38577);
nor U40609 (N_40609,N_38430,N_37515);
or U40610 (N_40610,N_39464,N_39961);
or U40611 (N_40611,N_38357,N_37685);
nand U40612 (N_40612,N_39848,N_39946);
xor U40613 (N_40613,N_39869,N_39920);
and U40614 (N_40614,N_39331,N_39272);
nand U40615 (N_40615,N_38420,N_39847);
or U40616 (N_40616,N_38873,N_39212);
nand U40617 (N_40617,N_39611,N_38800);
nand U40618 (N_40618,N_39721,N_37959);
nor U40619 (N_40619,N_39673,N_39463);
or U40620 (N_40620,N_38427,N_38872);
or U40621 (N_40621,N_39378,N_39330);
xor U40622 (N_40622,N_37521,N_39589);
nor U40623 (N_40623,N_39528,N_37731);
nand U40624 (N_40624,N_39367,N_39892);
nor U40625 (N_40625,N_37827,N_38067);
and U40626 (N_40626,N_38325,N_37845);
or U40627 (N_40627,N_39546,N_39755);
nor U40628 (N_40628,N_39717,N_39789);
and U40629 (N_40629,N_38924,N_38699);
and U40630 (N_40630,N_39692,N_38874);
nand U40631 (N_40631,N_39413,N_39011);
or U40632 (N_40632,N_39578,N_37851);
nor U40633 (N_40633,N_39748,N_39316);
nor U40634 (N_40634,N_39552,N_38331);
xor U40635 (N_40635,N_39099,N_38510);
nor U40636 (N_40636,N_38141,N_38853);
xor U40637 (N_40637,N_38119,N_37602);
nand U40638 (N_40638,N_39028,N_39102);
and U40639 (N_40639,N_38680,N_38810);
and U40640 (N_40640,N_39455,N_38170);
or U40641 (N_40641,N_37882,N_38452);
and U40642 (N_40642,N_39899,N_39505);
or U40643 (N_40643,N_39103,N_38803);
nor U40644 (N_40644,N_38993,N_39460);
and U40645 (N_40645,N_39745,N_38687);
and U40646 (N_40646,N_38565,N_38207);
nor U40647 (N_40647,N_38949,N_39907);
and U40648 (N_40648,N_38609,N_39694);
or U40649 (N_40649,N_38541,N_38237);
nand U40650 (N_40650,N_38723,N_38550);
and U40651 (N_40651,N_38198,N_38905);
nor U40652 (N_40652,N_39539,N_38756);
nor U40653 (N_40653,N_38070,N_37571);
nor U40654 (N_40654,N_38701,N_39074);
and U40655 (N_40655,N_39631,N_37777);
or U40656 (N_40656,N_38941,N_38807);
nor U40657 (N_40657,N_37941,N_38893);
or U40658 (N_40658,N_39536,N_39791);
and U40659 (N_40659,N_39747,N_39299);
and U40660 (N_40660,N_39263,N_39921);
nor U40661 (N_40661,N_39038,N_37877);
or U40662 (N_40662,N_39982,N_39407);
nand U40663 (N_40663,N_39291,N_38959);
and U40664 (N_40664,N_39826,N_38877);
nand U40665 (N_40665,N_38373,N_38706);
and U40666 (N_40666,N_38434,N_39172);
or U40667 (N_40667,N_38734,N_38253);
or U40668 (N_40668,N_39149,N_38319);
or U40669 (N_40669,N_39867,N_39649);
and U40670 (N_40670,N_39861,N_39094);
nand U40671 (N_40671,N_39733,N_38923);
nand U40672 (N_40672,N_38279,N_38147);
and U40673 (N_40673,N_38289,N_37934);
or U40674 (N_40674,N_39390,N_38718);
nand U40675 (N_40675,N_39502,N_39477);
xnor U40676 (N_40676,N_39560,N_39893);
nor U40677 (N_40677,N_38720,N_38844);
nor U40678 (N_40678,N_38056,N_37842);
nor U40679 (N_40679,N_38278,N_37551);
and U40680 (N_40680,N_39681,N_38100);
or U40681 (N_40681,N_39797,N_38078);
or U40682 (N_40682,N_38692,N_39086);
nand U40683 (N_40683,N_37562,N_37949);
or U40684 (N_40684,N_38284,N_37655);
nand U40685 (N_40685,N_39150,N_39583);
nand U40686 (N_40686,N_39421,N_38260);
or U40687 (N_40687,N_38505,N_39939);
or U40688 (N_40688,N_37525,N_37707);
or U40689 (N_40689,N_39970,N_38677);
nor U40690 (N_40690,N_38013,N_39904);
nor U40691 (N_40691,N_39003,N_38994);
nand U40692 (N_40692,N_38588,N_39773);
or U40693 (N_40693,N_37976,N_37618);
nor U40694 (N_40694,N_38875,N_38123);
nand U40695 (N_40695,N_39089,N_38344);
xor U40696 (N_40696,N_38904,N_38151);
or U40697 (N_40697,N_39444,N_39297);
nor U40698 (N_40698,N_38704,N_38591);
xor U40699 (N_40699,N_38092,N_38517);
nand U40700 (N_40700,N_38448,N_38139);
xnor U40701 (N_40701,N_39384,N_39828);
or U40702 (N_40702,N_38095,N_38617);
nor U40703 (N_40703,N_38788,N_38782);
nand U40704 (N_40704,N_39561,N_38674);
nor U40705 (N_40705,N_38530,N_38350);
and U40706 (N_40706,N_38210,N_38638);
nor U40707 (N_40707,N_37547,N_38174);
and U40708 (N_40708,N_38707,N_38811);
nor U40709 (N_40709,N_39635,N_38977);
nor U40710 (N_40710,N_39084,N_39059);
and U40711 (N_40711,N_39600,N_38433);
xor U40712 (N_40712,N_39542,N_38661);
and U40713 (N_40713,N_39602,N_39239);
and U40714 (N_40714,N_38553,N_39551);
xnor U40715 (N_40715,N_38573,N_39637);
nor U40716 (N_40716,N_39777,N_38166);
and U40717 (N_40717,N_37889,N_37693);
and U40718 (N_40718,N_39275,N_38440);
xnor U40719 (N_40719,N_37740,N_38691);
nor U40720 (N_40720,N_38001,N_38152);
xor U40721 (N_40721,N_39009,N_38545);
nand U40722 (N_40722,N_39827,N_38489);
xor U40723 (N_40723,N_39695,N_38946);
or U40724 (N_40724,N_39061,N_37500);
nand U40725 (N_40725,N_39422,N_37743);
or U40726 (N_40726,N_38625,N_39741);
or U40727 (N_40727,N_38144,N_37805);
and U40728 (N_40728,N_39835,N_39864);
nor U40729 (N_40729,N_38742,N_39506);
nor U40730 (N_40730,N_37614,N_39683);
and U40731 (N_40731,N_38999,N_39230);
or U40732 (N_40732,N_37929,N_39908);
or U40733 (N_40733,N_39934,N_39839);
and U40734 (N_40734,N_38955,N_38404);
nand U40735 (N_40735,N_39220,N_38156);
xor U40736 (N_40736,N_37945,N_39793);
and U40737 (N_40737,N_37840,N_38843);
nor U40738 (N_40738,N_39206,N_38566);
and U40739 (N_40739,N_39401,N_39186);
or U40740 (N_40740,N_38790,N_37897);
and U40741 (N_40741,N_39930,N_38326);
and U40742 (N_40742,N_39324,N_38683);
and U40743 (N_40743,N_39588,N_39193);
nand U40744 (N_40744,N_37792,N_38169);
nand U40745 (N_40745,N_38437,N_38369);
and U40746 (N_40746,N_39617,N_38249);
and U40747 (N_40747,N_38849,N_39171);
nor U40748 (N_40748,N_38259,N_38286);
or U40749 (N_40749,N_38963,N_38269);
and U40750 (N_40750,N_37689,N_39591);
and U40751 (N_40751,N_39200,N_38535);
xor U40752 (N_40752,N_38567,N_38032);
xnor U40753 (N_40753,N_38328,N_38042);
nor U40754 (N_40754,N_39445,N_39646);
or U40755 (N_40755,N_38537,N_39769);
nor U40756 (N_40756,N_39334,N_37639);
nand U40757 (N_40757,N_39133,N_39565);
or U40758 (N_40758,N_39599,N_39303);
nor U40759 (N_40759,N_38145,N_37732);
or U40760 (N_40760,N_38329,N_38655);
nor U40761 (N_40761,N_39244,N_37673);
nor U40762 (N_40762,N_37972,N_38731);
nand U40763 (N_40763,N_37509,N_38173);
or U40764 (N_40764,N_38656,N_39983);
xor U40765 (N_40765,N_37938,N_37823);
or U40766 (N_40766,N_39620,N_37545);
and U40767 (N_40767,N_37737,N_38759);
and U40768 (N_40768,N_38302,N_39516);
xor U40769 (N_40769,N_37952,N_38824);
nand U40770 (N_40770,N_39023,N_38543);
xnor U40771 (N_40771,N_39155,N_37931);
nand U40772 (N_40772,N_38970,N_39030);
nand U40773 (N_40773,N_39062,N_38758);
nor U40774 (N_40774,N_39216,N_39262);
xor U40775 (N_40775,N_39140,N_39451);
xnor U40776 (N_40776,N_38135,N_38668);
nand U40777 (N_40777,N_38429,N_39963);
xor U40778 (N_40778,N_38823,N_39728);
nor U40779 (N_40779,N_37531,N_38255);
nor U40780 (N_40780,N_38019,N_37637);
and U40781 (N_40781,N_38076,N_38719);
nand U40782 (N_40782,N_38722,N_37787);
xor U40783 (N_40783,N_39131,N_37883);
and U40784 (N_40784,N_38654,N_38459);
nor U40785 (N_40785,N_38771,N_38584);
xnor U40786 (N_40786,N_38754,N_37714);
and U40787 (N_40787,N_39070,N_39123);
nand U40788 (N_40788,N_37596,N_38121);
nor U40789 (N_40789,N_37677,N_37786);
and U40790 (N_40790,N_38534,N_39020);
and U40791 (N_40791,N_38168,N_38470);
or U40792 (N_40792,N_39574,N_39332);
or U40793 (N_40793,N_39110,N_39974);
and U40794 (N_40794,N_37643,N_37682);
nand U40795 (N_40795,N_39372,N_38634);
nor U40796 (N_40796,N_38597,N_37718);
nor U40797 (N_40797,N_38997,N_39443);
nand U40798 (N_40798,N_39180,N_38112);
nand U40799 (N_40799,N_38153,N_37703);
nor U40800 (N_40800,N_38608,N_38082);
nand U40801 (N_40801,N_39743,N_39295);
and U40802 (N_40802,N_37975,N_37995);
or U40803 (N_40803,N_39400,N_39004);
and U40804 (N_40804,N_38361,N_38862);
nand U40805 (N_40805,N_37663,N_38948);
and U40806 (N_40806,N_37694,N_38455);
nor U40807 (N_40807,N_39392,N_39136);
xor U40808 (N_40808,N_38292,N_39355);
or U40809 (N_40809,N_37863,N_38897);
xor U40810 (N_40810,N_38477,N_38400);
nand U40811 (N_40811,N_39688,N_39437);
xnor U40812 (N_40812,N_39568,N_37610);
nand U40813 (N_40813,N_38944,N_38628);
or U40814 (N_40814,N_37814,N_37819);
nor U40815 (N_40815,N_38961,N_38768);
or U40816 (N_40816,N_39991,N_37751);
nor U40817 (N_40817,N_37527,N_37625);
nand U40818 (N_40818,N_37757,N_37912);
nand U40819 (N_40819,N_39596,N_38518);
xnor U40820 (N_40820,N_38599,N_37848);
or U40821 (N_40821,N_39329,N_38646);
nand U40822 (N_40822,N_39668,N_38562);
and U40823 (N_40823,N_39240,N_37713);
or U40824 (N_40824,N_39520,N_39987);
nor U40825 (N_40825,N_38195,N_38947);
nand U40826 (N_40826,N_38035,N_37544);
or U40827 (N_40827,N_38930,N_38034);
nor U40828 (N_40828,N_39629,N_39643);
and U40829 (N_40829,N_38484,N_39855);
and U40830 (N_40830,N_39154,N_39830);
or U40831 (N_40831,N_38871,N_38777);
or U40832 (N_40832,N_37804,N_37505);
nand U40833 (N_40833,N_38431,N_38308);
nand U40834 (N_40834,N_38309,N_39135);
nand U40835 (N_40835,N_37738,N_39166);
nor U40836 (N_40836,N_39281,N_39164);
and U40837 (N_40837,N_38028,N_37501);
nand U40838 (N_40838,N_39729,N_38010);
or U40839 (N_40839,N_39804,N_37763);
nand U40840 (N_40840,N_38054,N_38230);
nand U40841 (N_40841,N_39973,N_38635);
nor U40842 (N_40842,N_39348,N_38651);
or U40843 (N_40843,N_38006,N_38301);
xnor U40844 (N_40844,N_39055,N_39619);
and U40845 (N_40845,N_38191,N_39529);
or U40846 (N_40846,N_37702,N_39559);
and U40847 (N_40847,N_39675,N_38040);
or U40848 (N_40848,N_37891,N_37725);
and U40849 (N_40849,N_38715,N_38244);
or U40850 (N_40850,N_37806,N_38729);
and U40851 (N_40851,N_37634,N_38449);
or U40852 (N_40852,N_37724,N_38343);
or U40853 (N_40853,N_37754,N_39799);
nand U40854 (N_40854,N_39514,N_37728);
nand U40855 (N_40855,N_39001,N_38227);
and U40856 (N_40856,N_38979,N_39423);
nor U40857 (N_40857,N_38708,N_39885);
nand U40858 (N_40858,N_38583,N_39152);
or U40859 (N_40859,N_39610,N_38428);
xor U40860 (N_40860,N_39249,N_38385);
xor U40861 (N_40861,N_38022,N_39903);
xnor U40862 (N_40862,N_38688,N_38860);
nand U40863 (N_40863,N_39368,N_38128);
xnor U40864 (N_40864,N_39868,N_39072);
xnor U40865 (N_40865,N_39518,N_38221);
and U40866 (N_40866,N_39616,N_39833);
nor U40867 (N_40867,N_38819,N_39731);
or U40868 (N_40868,N_37533,N_39184);
and U40869 (N_40869,N_38324,N_39669);
xor U40870 (N_40870,N_39586,N_38978);
and U40871 (N_40871,N_38769,N_39628);
and U40872 (N_40872,N_38111,N_37958);
or U40873 (N_40873,N_38610,N_37699);
and U40874 (N_40874,N_38673,N_38061);
nor U40875 (N_40875,N_39659,N_39816);
nor U40876 (N_40876,N_38839,N_38027);
nand U40877 (N_40877,N_39879,N_39853);
or U40878 (N_40878,N_38622,N_38273);
nor U40879 (N_40879,N_39192,N_37841);
nor U40880 (N_40880,N_39044,N_39918);
or U40881 (N_40881,N_39572,N_38713);
nand U40882 (N_40882,N_39026,N_37776);
and U40883 (N_40883,N_39276,N_37595);
and U40884 (N_40884,N_38732,N_38848);
or U40885 (N_40885,N_38797,N_39393);
nor U40886 (N_40886,N_38515,N_39434);
nand U40887 (N_40887,N_39456,N_38925);
or U40888 (N_40888,N_39715,N_38122);
or U40889 (N_40889,N_39739,N_38645);
nor U40890 (N_40890,N_38297,N_39259);
nor U40891 (N_40891,N_39813,N_38409);
nand U40892 (N_40892,N_39707,N_38937);
nand U40893 (N_40893,N_38197,N_38581);
nor U40894 (N_40894,N_37646,N_39779);
and U40895 (N_40895,N_38142,N_38928);
and U40896 (N_40896,N_39642,N_37865);
nand U40897 (N_40897,N_39346,N_39126);
xor U40898 (N_40898,N_38859,N_39878);
nand U40899 (N_40899,N_38178,N_38681);
nor U40900 (N_40900,N_38749,N_38482);
or U40901 (N_40901,N_39595,N_37604);
and U40902 (N_40902,N_38785,N_38212);
or U40903 (N_40903,N_37798,N_38657);
nor U40904 (N_40904,N_38737,N_37854);
nand U40905 (N_40905,N_38209,N_38445);
nand U40906 (N_40906,N_37688,N_39995);
nand U40907 (N_40907,N_39818,N_38068);
nand U40908 (N_40908,N_37774,N_38980);
and U40909 (N_40909,N_39576,N_39073);
or U40910 (N_40910,N_39775,N_38900);
and U40911 (N_40911,N_39730,N_39757);
nand U40912 (N_40912,N_38488,N_38576);
or U40913 (N_40913,N_38763,N_39442);
and U40914 (N_40914,N_38044,N_39215);
and U40915 (N_40915,N_37557,N_39527);
nand U40916 (N_40916,N_37846,N_39824);
xor U40917 (N_40917,N_38724,N_39491);
nand U40918 (N_40918,N_38252,N_37965);
or U40919 (N_40919,N_38282,N_39760);
nor U40920 (N_40920,N_39187,N_38682);
and U40921 (N_40921,N_39039,N_37536);
or U40922 (N_40922,N_38096,N_38228);
nand U40923 (N_40923,N_37830,N_37998);
or U40924 (N_40924,N_38229,N_38456);
and U40925 (N_40925,N_37876,N_39313);
or U40926 (N_40926,N_37837,N_38836);
or U40927 (N_40927,N_39570,N_37843);
nand U40928 (N_40928,N_38089,N_38903);
and U40929 (N_40929,N_38233,N_39517);
xor U40930 (N_40930,N_38987,N_39898);
and U40931 (N_40931,N_39815,N_38818);
nor U40932 (N_40932,N_37566,N_39195);
or U40933 (N_40933,N_37717,N_38593);
nor U40934 (N_40934,N_37917,N_38184);
and U40935 (N_40935,N_38629,N_39702);
nand U40936 (N_40936,N_37899,N_37623);
xor U40937 (N_40937,N_38568,N_38995);
or U40938 (N_40938,N_38467,N_39179);
and U40939 (N_40939,N_37543,N_39936);
nor U40940 (N_40940,N_38914,N_39753);
or U40941 (N_40941,N_38546,N_38349);
xor U40942 (N_40942,N_38559,N_38047);
and U40943 (N_40943,N_38876,N_38801);
nor U40944 (N_40944,N_37649,N_39373);
or U40945 (N_40945,N_37518,N_39173);
and U40946 (N_40946,N_39798,N_39843);
or U40947 (N_40947,N_37603,N_38106);
nor U40948 (N_40948,N_37552,N_39667);
nand U40949 (N_40949,N_38320,N_38659);
nand U40950 (N_40950,N_38513,N_37795);
or U40951 (N_40951,N_38150,N_38592);
nand U40952 (N_40952,N_39802,N_39553);
and U40953 (N_40953,N_39942,N_39377);
nor U40954 (N_40954,N_38878,N_39754);
nor U40955 (N_40955,N_38520,N_39531);
or U40956 (N_40956,N_37542,N_37642);
nor U40957 (N_40957,N_39497,N_38833);
nand U40958 (N_40958,N_38524,N_38496);
or U40959 (N_40959,N_39402,N_37940);
nor U40960 (N_40960,N_39909,N_39923);
nor U40961 (N_40961,N_39993,N_38270);
nor U40962 (N_40962,N_37752,N_37905);
or U40963 (N_40963,N_39641,N_38621);
and U40964 (N_40964,N_39890,N_39265);
nand U40965 (N_40965,N_38589,N_39691);
nor U40966 (N_40966,N_37567,N_38382);
and U40967 (N_40967,N_38102,N_38571);
and U40968 (N_40968,N_38601,N_39161);
or U40969 (N_40969,N_39555,N_37687);
nand U40970 (N_40970,N_39049,N_39972);
or U40971 (N_40971,N_39492,N_39713);
nand U40972 (N_40972,N_38943,N_39365);
nand U40973 (N_40973,N_39430,N_38203);
nand U40974 (N_40974,N_37648,N_38062);
nor U40975 (N_40975,N_38992,N_38624);
or U40976 (N_40976,N_38458,N_39943);
nor U40977 (N_40977,N_37832,N_38921);
or U40978 (N_40978,N_39398,N_39342);
xnor U40979 (N_40979,N_39661,N_39682);
nor U40980 (N_40980,N_37546,N_37583);
nor U40981 (N_40981,N_39752,N_39447);
nor U40982 (N_40982,N_39734,N_38882);
or U40983 (N_40983,N_39096,N_38982);
nand U40984 (N_40984,N_39151,N_39375);
nand U40985 (N_40985,N_39415,N_38867);
nor U40986 (N_40986,N_39665,N_39056);
nor U40987 (N_40987,N_37768,N_38446);
or U40988 (N_40988,N_39609,N_39335);
or U40989 (N_40989,N_38678,N_38116);
nor U40990 (N_40990,N_38134,N_38852);
and U40991 (N_40991,N_39746,N_39647);
nor U40992 (N_40992,N_38183,N_38245);
or U40993 (N_40993,N_37744,N_38342);
and U40994 (N_40994,N_37790,N_39380);
and U40995 (N_40995,N_38998,N_38425);
and U40996 (N_40996,N_38641,N_39053);
or U40997 (N_40997,N_39912,N_39159);
nor U40998 (N_40998,N_39735,N_39351);
or U40999 (N_40999,N_38855,N_39653);
nor U41000 (N_41000,N_38276,N_39318);
or U41001 (N_41001,N_37606,N_37511);
nor U41002 (N_41002,N_38421,N_38306);
and U41003 (N_41003,N_37520,N_39917);
nand U41004 (N_41004,N_39783,N_37911);
and U41005 (N_41005,N_37686,N_38757);
nor U41006 (N_41006,N_38675,N_38933);
or U41007 (N_41007,N_38177,N_37691);
nor U41008 (N_41008,N_39786,N_38967);
xor U41009 (N_41009,N_38243,N_37924);
nor U41010 (N_41010,N_38503,N_39989);
or U41011 (N_41011,N_38075,N_37918);
and U41012 (N_41012,N_37741,N_38354);
and U41013 (N_41013,N_39670,N_37578);
nor U41014 (N_41014,N_39289,N_37933);
nor U41015 (N_41015,N_39425,N_39012);
or U41016 (N_41016,N_39328,N_39501);
or U41017 (N_41017,N_39840,N_38316);
nor U41018 (N_41018,N_39356,N_39207);
xnor U41019 (N_41019,N_38097,N_37640);
nor U41020 (N_41020,N_38600,N_39031);
or U41021 (N_41021,N_38381,N_38339);
nor U41022 (N_41022,N_39341,N_38636);
or U41023 (N_41023,N_38626,N_39765);
or U41024 (N_41024,N_38913,N_37973);
nand U41025 (N_41025,N_37907,N_37519);
and U41026 (N_41026,N_38586,N_39660);
nand U41027 (N_41027,N_39842,N_39090);
or U41028 (N_41028,N_39687,N_37983);
or U41029 (N_41029,N_39720,N_37849);
or U41030 (N_41030,N_39191,N_38337);
nor U41031 (N_41031,N_37574,N_38616);
nand U41032 (N_41032,N_38396,N_38670);
nand U41033 (N_41033,N_37867,N_39587);
nand U41034 (N_41034,N_39058,N_39684);
nor U41035 (N_41035,N_37797,N_39228);
or U41036 (N_41036,N_39048,N_39941);
nor U41037 (N_41037,N_38973,N_37629);
or U41038 (N_41038,N_37523,N_38310);
nor U41039 (N_41039,N_39478,N_38644);
and U41040 (N_41040,N_37802,N_39340);
nor U41041 (N_41041,N_38461,N_37903);
nand U41042 (N_41042,N_37530,N_39082);
nor U41043 (N_41043,N_39573,N_39431);
or U41044 (N_41044,N_38736,N_39770);
nor U41045 (N_41045,N_39996,N_38298);
or U41046 (N_41046,N_38735,N_39737);
or U41047 (N_41047,N_37861,N_39165);
nor U41048 (N_41048,N_38696,N_37993);
nand U41049 (N_41049,N_37508,N_38026);
nor U41050 (N_41050,N_38049,N_38747);
xor U41051 (N_41051,N_38367,N_39948);
nor U41052 (N_41052,N_38466,N_37844);
xnor U41053 (N_41053,N_38048,N_38934);
nor U41054 (N_41054,N_39476,N_39662);
nand U41055 (N_41055,N_37986,N_38940);
nand U41056 (N_41056,N_38548,N_39294);
nand U41057 (N_41057,N_38051,N_37885);
or U41058 (N_41058,N_38073,N_39359);
and U41059 (N_41059,N_38261,N_39984);
and U41060 (N_41060,N_39523,N_38598);
and U41061 (N_41061,N_37695,N_38288);
or U41062 (N_41062,N_37534,N_39304);
and U41063 (N_41063,N_39985,N_38630);
xor U41064 (N_41064,N_39844,N_37675);
nor U41065 (N_41065,N_38712,N_38356);
nor U41066 (N_41066,N_37539,N_38180);
xor U41067 (N_41067,N_37585,N_39900);
or U41068 (N_41068,N_39360,N_37510);
xnor U41069 (N_41069,N_38305,N_38752);
nor U41070 (N_41070,N_38175,N_37781);
or U41071 (N_41071,N_38498,N_38494);
xnor U41072 (N_41072,N_37779,N_39284);
or U41073 (N_41073,N_39470,N_38118);
and U41074 (N_41074,N_38223,N_39780);
nor U41075 (N_41075,N_38779,N_39296);
and U41076 (N_41076,N_38315,N_39254);
and U41077 (N_41077,N_37676,N_38776);
nand U41078 (N_41078,N_38507,N_39857);
nand U41079 (N_41079,N_39027,N_38898);
and U41080 (N_41080,N_38702,N_38746);
or U41081 (N_41081,N_39795,N_37507);
or U41082 (N_41082,N_37898,N_37860);
nor U41083 (N_41083,N_38631,N_39285);
nor U41084 (N_41084,N_38294,N_38475);
or U41085 (N_41085,N_39286,N_38829);
or U41086 (N_41086,N_37926,N_38024);
nand U41087 (N_41087,N_38386,N_39603);
or U41088 (N_41088,N_37568,N_38762);
and U41089 (N_41089,N_39182,N_38880);
and U41090 (N_41090,N_38908,N_37778);
and U41091 (N_41091,N_39479,N_39162);
nand U41092 (N_41092,N_39146,N_39290);
nor U41093 (N_41093,N_38927,N_38964);
and U41094 (N_41094,N_39266,N_39957);
or U41095 (N_41095,N_38380,N_39156);
and U41096 (N_41096,N_39781,N_38710);
or U41097 (N_41097,N_38966,N_38892);
xnor U41098 (N_41098,N_37654,N_39540);
or U41099 (N_41099,N_37630,N_38447);
nand U41100 (N_41100,N_37794,N_38220);
or U41101 (N_41101,N_37895,N_37858);
nand U41102 (N_41102,N_38041,N_37720);
or U41103 (N_41103,N_37528,N_38176);
xor U41104 (N_41104,N_37690,N_39106);
and U41105 (N_41105,N_37652,N_39287);
nor U41106 (N_41106,N_37626,N_39227);
or U41107 (N_41107,N_37748,N_38190);
xnor U41108 (N_41108,N_38050,N_37892);
nand U41109 (N_41109,N_37735,N_38784);
nor U41110 (N_41110,N_38512,N_39585);
or U41111 (N_41111,N_38623,N_38478);
nor U41112 (N_41112,N_37772,N_38295);
nand U41113 (N_41113,N_38125,N_39190);
and U41114 (N_41114,N_39886,N_37906);
nand U41115 (N_41115,N_37622,N_38378);
nand U41116 (N_41116,N_38232,N_37674);
or U41117 (N_41117,N_37922,N_39803);
and U41118 (N_41118,N_38200,N_37835);
xor U41119 (N_41119,N_39955,N_38486);
nand U41120 (N_41120,N_38578,N_38911);
nand U41121 (N_41121,N_39806,N_39554);
nand U41122 (N_41122,N_38352,N_39168);
or U41123 (N_41123,N_39080,N_38084);
nor U41124 (N_41124,N_39371,N_37980);
or U41125 (N_41125,N_38293,N_39875);
nand U41126 (N_41126,N_37758,N_39882);
nor U41127 (N_41127,N_38490,N_39808);
or U41128 (N_41128,N_38318,N_38555);
or U41129 (N_41129,N_38225,N_38851);
nor U41130 (N_41130,N_39208,N_38088);
nand U41131 (N_41131,N_38650,N_38393);
xor U41132 (N_41132,N_39129,N_39396);
nand U41133 (N_41133,N_39088,N_38664);
or U41134 (N_41134,N_39809,N_39321);
or U41135 (N_41135,N_39045,N_38020);
nand U41136 (N_41136,N_37770,N_37756);
nor U41137 (N_41137,N_37947,N_37598);
or U41138 (N_41138,N_39496,N_37996);
nor U41139 (N_41139,N_37570,N_39534);
nand U41140 (N_41140,N_39256,N_39204);
xnor U41141 (N_41141,N_37671,N_39865);
and U41142 (N_41142,N_38799,N_39459);
or U41143 (N_41143,N_39349,N_38000);
or U41144 (N_41144,N_39280,N_38268);
or U41145 (N_41145,N_39928,N_39612);
nand U41146 (N_41146,N_37745,N_37852);
nor U41147 (N_41147,N_38942,N_38014);
nand U41148 (N_41148,N_39469,N_39143);
nor U41149 (N_41149,N_39432,N_38071);
nor U41150 (N_41150,N_37780,N_39834);
or U41151 (N_41151,N_37761,N_38126);
or U41152 (N_41152,N_39829,N_39338);
nand U41153 (N_41153,N_38362,N_37936);
or U41154 (N_41154,N_38808,N_38033);
or U41155 (N_41155,N_38377,N_38649);
xnor U41156 (N_41156,N_38358,N_39167);
and U41157 (N_41157,N_37765,N_39389);
nand U41158 (N_41158,N_37607,N_38016);
and U41159 (N_41159,N_38159,N_37785);
nor U41160 (N_41160,N_39147,N_38915);
and U41161 (N_41161,N_39300,N_38521);
and U41162 (N_41162,N_38906,N_37522);
or U41163 (N_41163,N_37888,N_37948);
and U41164 (N_41164,N_38825,N_38291);
and U41165 (N_41165,N_39544,N_38154);
nor U41166 (N_41166,N_39807,N_38322);
nand U41167 (N_41167,N_39871,N_39315);
xnor U41168 (N_41168,N_39714,N_37716);
xnor U41169 (N_41169,N_38407,N_38516);
nor U41170 (N_41170,N_38582,N_37939);
nor U41171 (N_41171,N_38039,N_39414);
nor U41172 (N_41172,N_39905,N_39071);
and U41173 (N_41173,N_39261,N_38751);
nand U41174 (N_41174,N_38025,N_39964);
nand U41175 (N_41175,N_39112,N_37573);
or U41176 (N_41176,N_37977,N_37524);
or U41177 (N_41177,N_39913,N_38426);
nand U41178 (N_41178,N_39805,N_38809);
nand U41179 (N_41179,N_39929,N_39592);
nand U41180 (N_41180,N_39137,N_39504);
and U41181 (N_41181,N_39764,N_38009);
nor U41182 (N_41182,N_37800,N_38211);
or U41183 (N_41183,N_38640,N_39068);
or U41184 (N_41184,N_37857,N_37532);
xor U41185 (N_41185,N_37641,N_38347);
and U41186 (N_41186,N_39601,N_37927);
and U41187 (N_41187,N_38960,N_39141);
and U41188 (N_41188,N_37591,N_38491);
nor U41189 (N_41189,N_38775,N_39198);
and U41190 (N_41190,N_39873,N_39253);
or U41191 (N_41191,N_38907,N_39724);
and U41192 (N_41192,N_37869,N_39887);
nor U41193 (N_41193,N_37638,N_39323);
xor U41194 (N_41194,N_39305,N_38379);
or U41195 (N_41195,N_39311,N_37815);
nand U41196 (N_41196,N_39435,N_39408);
nand U41197 (N_41197,N_39270,N_39312);
and U41198 (N_41198,N_39486,N_38693);
or U41199 (N_41199,N_38069,N_37681);
and U41200 (N_41200,N_38274,N_37771);
or U41201 (N_41201,N_39410,N_39157);
and U41202 (N_41202,N_39465,N_38909);
and U41203 (N_41203,N_37991,N_37783);
and U41204 (N_41204,N_37974,N_39621);
and U41205 (N_41205,N_38205,N_37569);
nor U41206 (N_41206,N_39712,N_39965);
or U41207 (N_41207,N_39483,N_39513);
and U41208 (N_41208,N_39111,N_39994);
or U41209 (N_41209,N_37529,N_38247);
nor U41210 (N_41210,N_38359,N_39679);
and U41211 (N_41211,N_38569,N_39762);
or U41212 (N_41212,N_38334,N_37698);
nand U41213 (N_41213,N_38105,N_39238);
or U41214 (N_41214,N_38814,N_37884);
nor U41215 (N_41215,N_38167,N_37729);
nor U41216 (N_41216,N_38832,N_39438);
and U41217 (N_41217,N_37989,N_39052);
or U41218 (N_41218,N_39651,N_39041);
and U41219 (N_41219,N_38258,N_39458);
or U41220 (N_41220,N_39914,N_38057);
and U41221 (N_41221,N_37967,N_38500);
nor U41222 (N_41222,N_38036,N_38716);
nand U41223 (N_41223,N_38525,N_38519);
nand U41224 (N_41224,N_37990,N_38528);
or U41225 (N_41225,N_37957,N_38896);
nand U41226 (N_41226,N_38968,N_39891);
xnor U41227 (N_41227,N_37541,N_39607);
xor U41228 (N_41228,N_38248,N_39858);
or U41229 (N_41229,N_38991,N_37554);
nor U41230 (N_41230,N_37810,N_38529);
and U41231 (N_41231,N_39508,N_37700);
or U41232 (N_41232,N_39214,N_38676);
xnor U41233 (N_41233,N_39931,N_38665);
nand U41234 (N_41234,N_38744,N_39302);
and U41235 (N_41235,N_39382,N_39953);
xnor U41236 (N_41236,N_37746,N_37565);
xnor U41237 (N_41237,N_39412,N_38642);
and U41238 (N_41238,N_37575,N_39236);
or U41239 (N_41239,N_39971,N_37868);
nand U41240 (N_41240,N_39274,N_39810);
nor U41241 (N_41241,N_37599,N_38602);
or U41242 (N_41242,N_38647,N_39881);
and U41243 (N_41243,N_39959,N_39385);
nor U41244 (N_41244,N_37826,N_38080);
nand U41245 (N_41245,N_39134,N_39699);
and U41246 (N_41246,N_37608,N_38965);
or U41247 (N_41247,N_39831,N_39352);
nand U41248 (N_41248,N_39357,N_38564);
nor U41249 (N_41249,N_38662,N_37946);
and U41250 (N_41250,N_38375,N_38021);
and U41251 (N_41251,N_38989,N_39894);
nor U41252 (N_41252,N_39029,N_37633);
and U41253 (N_41253,N_39285,N_38975);
nor U41254 (N_41254,N_39122,N_38307);
nand U41255 (N_41255,N_38467,N_38925);
nand U41256 (N_41256,N_38343,N_37752);
nand U41257 (N_41257,N_37900,N_39736);
nor U41258 (N_41258,N_38253,N_37660);
and U41259 (N_41259,N_37624,N_39950);
nand U41260 (N_41260,N_38051,N_39625);
or U41261 (N_41261,N_38087,N_38615);
nand U41262 (N_41262,N_38318,N_38203);
nand U41263 (N_41263,N_38330,N_38273);
and U41264 (N_41264,N_39764,N_39639);
or U41265 (N_41265,N_39860,N_39523);
xor U41266 (N_41266,N_38734,N_38019);
and U41267 (N_41267,N_38634,N_38808);
xnor U41268 (N_41268,N_38568,N_38439);
or U41269 (N_41269,N_38434,N_37988);
xor U41270 (N_41270,N_39906,N_39358);
nor U41271 (N_41271,N_38349,N_39617);
nand U41272 (N_41272,N_38345,N_38404);
or U41273 (N_41273,N_39168,N_37984);
nand U41274 (N_41274,N_38212,N_37621);
nand U41275 (N_41275,N_37627,N_37819);
and U41276 (N_41276,N_38953,N_38479);
and U41277 (N_41277,N_39484,N_38323);
nand U41278 (N_41278,N_38497,N_38074);
nor U41279 (N_41279,N_37633,N_38572);
or U41280 (N_41280,N_38174,N_39514);
and U41281 (N_41281,N_39068,N_38065);
and U41282 (N_41282,N_39077,N_37718);
and U41283 (N_41283,N_37929,N_37849);
or U41284 (N_41284,N_37719,N_38290);
and U41285 (N_41285,N_38312,N_39624);
and U41286 (N_41286,N_38601,N_39497);
or U41287 (N_41287,N_38564,N_39719);
xor U41288 (N_41288,N_39792,N_38469);
nor U41289 (N_41289,N_38826,N_38048);
nand U41290 (N_41290,N_38071,N_39253);
and U41291 (N_41291,N_37698,N_37545);
and U41292 (N_41292,N_39464,N_39711);
nand U41293 (N_41293,N_39314,N_38236);
nand U41294 (N_41294,N_38806,N_39237);
nor U41295 (N_41295,N_37682,N_38856);
or U41296 (N_41296,N_39801,N_38015);
nor U41297 (N_41297,N_38550,N_38580);
xor U41298 (N_41298,N_39927,N_39967);
or U41299 (N_41299,N_38448,N_37549);
and U41300 (N_41300,N_39751,N_39178);
nand U41301 (N_41301,N_38261,N_38518);
nand U41302 (N_41302,N_38708,N_38956);
and U41303 (N_41303,N_38768,N_37514);
nor U41304 (N_41304,N_38178,N_38834);
nor U41305 (N_41305,N_38335,N_37931);
and U41306 (N_41306,N_39135,N_38684);
nor U41307 (N_41307,N_38869,N_38016);
and U41308 (N_41308,N_39118,N_38705);
nor U41309 (N_41309,N_38356,N_38348);
and U41310 (N_41310,N_39922,N_37546);
or U41311 (N_41311,N_37765,N_37908);
and U41312 (N_41312,N_39840,N_39485);
xor U41313 (N_41313,N_39402,N_37898);
and U41314 (N_41314,N_38872,N_39247);
or U41315 (N_41315,N_38965,N_37709);
and U41316 (N_41316,N_39369,N_38849);
or U41317 (N_41317,N_39802,N_37726);
and U41318 (N_41318,N_39449,N_39534);
nor U41319 (N_41319,N_39542,N_39438);
nand U41320 (N_41320,N_37567,N_38583);
nor U41321 (N_41321,N_39311,N_38623);
and U41322 (N_41322,N_37511,N_38498);
nand U41323 (N_41323,N_37975,N_39834);
nand U41324 (N_41324,N_39254,N_38774);
nand U41325 (N_41325,N_39482,N_37982);
nor U41326 (N_41326,N_38631,N_39432);
xor U41327 (N_41327,N_38855,N_39143);
or U41328 (N_41328,N_39855,N_39892);
or U41329 (N_41329,N_39603,N_37689);
xnor U41330 (N_41330,N_39726,N_39602);
and U41331 (N_41331,N_38705,N_39368);
and U41332 (N_41332,N_39511,N_39853);
nor U41333 (N_41333,N_38866,N_39209);
or U41334 (N_41334,N_38601,N_39651);
nand U41335 (N_41335,N_39401,N_38453);
nor U41336 (N_41336,N_38725,N_39459);
nand U41337 (N_41337,N_39851,N_38441);
nor U41338 (N_41338,N_39036,N_38066);
xnor U41339 (N_41339,N_38710,N_38714);
nor U41340 (N_41340,N_37617,N_37985);
or U41341 (N_41341,N_37563,N_37664);
nor U41342 (N_41342,N_38088,N_38593);
or U41343 (N_41343,N_37647,N_38215);
and U41344 (N_41344,N_37892,N_37760);
or U41345 (N_41345,N_37933,N_39861);
nor U41346 (N_41346,N_37691,N_38323);
nor U41347 (N_41347,N_39429,N_39420);
nor U41348 (N_41348,N_38301,N_39595);
nand U41349 (N_41349,N_38082,N_37533);
nand U41350 (N_41350,N_38211,N_39048);
nand U41351 (N_41351,N_38432,N_39435);
and U41352 (N_41352,N_38582,N_39648);
or U41353 (N_41353,N_39413,N_39654);
or U41354 (N_41354,N_37983,N_38177);
nand U41355 (N_41355,N_38181,N_37573);
nor U41356 (N_41356,N_39378,N_38611);
nor U41357 (N_41357,N_39432,N_38042);
xor U41358 (N_41358,N_38387,N_38253);
nand U41359 (N_41359,N_37916,N_39685);
xnor U41360 (N_41360,N_38505,N_38651);
and U41361 (N_41361,N_39461,N_38862);
and U41362 (N_41362,N_38847,N_38431);
nor U41363 (N_41363,N_38242,N_37902);
or U41364 (N_41364,N_38376,N_39977);
nor U41365 (N_41365,N_37965,N_39613);
nor U41366 (N_41366,N_39753,N_39904);
nand U41367 (N_41367,N_39416,N_39110);
nor U41368 (N_41368,N_38652,N_39802);
nor U41369 (N_41369,N_39640,N_38169);
nor U41370 (N_41370,N_37550,N_37670);
and U41371 (N_41371,N_37699,N_37524);
nand U41372 (N_41372,N_37957,N_37507);
nand U41373 (N_41373,N_39265,N_39184);
xnor U41374 (N_41374,N_39804,N_38003);
or U41375 (N_41375,N_37862,N_38771);
nor U41376 (N_41376,N_38666,N_37698);
and U41377 (N_41377,N_39498,N_38246);
or U41378 (N_41378,N_39409,N_39273);
or U41379 (N_41379,N_39287,N_39953);
or U41380 (N_41380,N_39546,N_38475);
nor U41381 (N_41381,N_37708,N_39718);
and U41382 (N_41382,N_38555,N_38884);
nand U41383 (N_41383,N_38064,N_39694);
or U41384 (N_41384,N_39082,N_39867);
nand U41385 (N_41385,N_37646,N_39180);
and U41386 (N_41386,N_39758,N_39998);
or U41387 (N_41387,N_37790,N_39539);
or U41388 (N_41388,N_37796,N_37516);
nor U41389 (N_41389,N_38849,N_39501);
and U41390 (N_41390,N_37760,N_39995);
nor U41391 (N_41391,N_38158,N_39304);
nand U41392 (N_41392,N_38174,N_38107);
nor U41393 (N_41393,N_37912,N_38257);
nor U41394 (N_41394,N_38916,N_39787);
xnor U41395 (N_41395,N_39246,N_38796);
or U41396 (N_41396,N_39638,N_37920);
nand U41397 (N_41397,N_38118,N_37855);
or U41398 (N_41398,N_38348,N_38002);
nand U41399 (N_41399,N_38083,N_37743);
and U41400 (N_41400,N_39137,N_38285);
or U41401 (N_41401,N_38955,N_37915);
nand U41402 (N_41402,N_38564,N_39897);
nand U41403 (N_41403,N_39940,N_38911);
xor U41404 (N_41404,N_37647,N_38326);
and U41405 (N_41405,N_37794,N_39975);
nor U41406 (N_41406,N_38776,N_38944);
or U41407 (N_41407,N_39509,N_38260);
and U41408 (N_41408,N_38541,N_37965);
nor U41409 (N_41409,N_37649,N_38966);
or U41410 (N_41410,N_39629,N_38581);
nand U41411 (N_41411,N_37675,N_37924);
and U41412 (N_41412,N_38965,N_38935);
nand U41413 (N_41413,N_39915,N_38201);
and U41414 (N_41414,N_38525,N_38586);
and U41415 (N_41415,N_39829,N_38502);
and U41416 (N_41416,N_38899,N_39575);
nand U41417 (N_41417,N_39006,N_38668);
and U41418 (N_41418,N_38634,N_39502);
or U41419 (N_41419,N_37777,N_37986);
or U41420 (N_41420,N_38992,N_38577);
nand U41421 (N_41421,N_37750,N_39206);
nor U41422 (N_41422,N_38514,N_38507);
or U41423 (N_41423,N_39135,N_39111);
xor U41424 (N_41424,N_37518,N_38469);
xnor U41425 (N_41425,N_38168,N_39720);
or U41426 (N_41426,N_39853,N_37535);
and U41427 (N_41427,N_38850,N_39528);
and U41428 (N_41428,N_39927,N_38968);
nand U41429 (N_41429,N_39813,N_39310);
nor U41430 (N_41430,N_38920,N_39231);
nand U41431 (N_41431,N_39014,N_37642);
nand U41432 (N_41432,N_39503,N_37592);
nor U41433 (N_41433,N_37655,N_38646);
or U41434 (N_41434,N_39527,N_39992);
xnor U41435 (N_41435,N_38792,N_38111);
nand U41436 (N_41436,N_37915,N_39276);
nand U41437 (N_41437,N_37588,N_39626);
nor U41438 (N_41438,N_39546,N_39279);
and U41439 (N_41439,N_37673,N_37911);
nor U41440 (N_41440,N_38649,N_39870);
nor U41441 (N_41441,N_39782,N_38447);
and U41442 (N_41442,N_39184,N_38388);
nand U41443 (N_41443,N_39992,N_38553);
and U41444 (N_41444,N_38135,N_39760);
nand U41445 (N_41445,N_37758,N_39155);
or U41446 (N_41446,N_38958,N_37558);
and U41447 (N_41447,N_37523,N_38523);
nor U41448 (N_41448,N_39501,N_38412);
and U41449 (N_41449,N_38677,N_38895);
xor U41450 (N_41450,N_39047,N_38665);
nor U41451 (N_41451,N_38490,N_39472);
and U41452 (N_41452,N_38116,N_38035);
nand U41453 (N_41453,N_38824,N_39785);
or U41454 (N_41454,N_38572,N_39304);
or U41455 (N_41455,N_38351,N_37992);
nand U41456 (N_41456,N_39778,N_39695);
or U41457 (N_41457,N_38976,N_38040);
or U41458 (N_41458,N_37651,N_39933);
or U41459 (N_41459,N_39080,N_38354);
or U41460 (N_41460,N_38116,N_38074);
nor U41461 (N_41461,N_37917,N_39965);
nand U41462 (N_41462,N_37528,N_38386);
nand U41463 (N_41463,N_38285,N_39868);
nand U41464 (N_41464,N_39441,N_38546);
nand U41465 (N_41465,N_38049,N_39706);
or U41466 (N_41466,N_39550,N_38853);
and U41467 (N_41467,N_37558,N_39925);
xnor U41468 (N_41468,N_37586,N_39401);
or U41469 (N_41469,N_38067,N_38838);
nand U41470 (N_41470,N_39000,N_39301);
or U41471 (N_41471,N_39010,N_39062);
and U41472 (N_41472,N_38598,N_39198);
or U41473 (N_41473,N_37988,N_38360);
nand U41474 (N_41474,N_38969,N_39305);
or U41475 (N_41475,N_38768,N_38373);
nor U41476 (N_41476,N_38780,N_38637);
and U41477 (N_41477,N_39447,N_37786);
nand U41478 (N_41478,N_37988,N_38170);
xnor U41479 (N_41479,N_39166,N_39340);
xor U41480 (N_41480,N_38246,N_39683);
or U41481 (N_41481,N_39253,N_38658);
nand U41482 (N_41482,N_39252,N_38755);
nand U41483 (N_41483,N_37786,N_37762);
or U41484 (N_41484,N_38085,N_38401);
nand U41485 (N_41485,N_37520,N_37960);
nand U41486 (N_41486,N_38365,N_38906);
or U41487 (N_41487,N_39164,N_39387);
and U41488 (N_41488,N_39038,N_38441);
nand U41489 (N_41489,N_38664,N_37978);
nor U41490 (N_41490,N_37823,N_37607);
and U41491 (N_41491,N_39722,N_38082);
nand U41492 (N_41492,N_37892,N_38755);
nor U41493 (N_41493,N_38603,N_39521);
or U41494 (N_41494,N_38037,N_39306);
nand U41495 (N_41495,N_37995,N_38356);
or U41496 (N_41496,N_38247,N_38334);
or U41497 (N_41497,N_39745,N_39131);
nor U41498 (N_41498,N_39354,N_39145);
xnor U41499 (N_41499,N_37712,N_37854);
nor U41500 (N_41500,N_38087,N_39453);
and U41501 (N_41501,N_38631,N_38983);
nor U41502 (N_41502,N_38195,N_37865);
xnor U41503 (N_41503,N_37610,N_38275);
and U41504 (N_41504,N_39004,N_37695);
and U41505 (N_41505,N_39533,N_39453);
or U41506 (N_41506,N_37577,N_38033);
or U41507 (N_41507,N_38800,N_38271);
nor U41508 (N_41508,N_38764,N_38787);
or U41509 (N_41509,N_39130,N_39402);
nand U41510 (N_41510,N_39328,N_37730);
xor U41511 (N_41511,N_38566,N_37714);
nor U41512 (N_41512,N_38000,N_39784);
xor U41513 (N_41513,N_39317,N_38998);
or U41514 (N_41514,N_38687,N_39290);
and U41515 (N_41515,N_37626,N_39875);
xor U41516 (N_41516,N_37544,N_38467);
nand U41517 (N_41517,N_37856,N_39473);
nand U41518 (N_41518,N_37656,N_37638);
and U41519 (N_41519,N_38675,N_39296);
nor U41520 (N_41520,N_38677,N_37789);
nand U41521 (N_41521,N_38460,N_38983);
nand U41522 (N_41522,N_39423,N_39910);
or U41523 (N_41523,N_38503,N_37823);
or U41524 (N_41524,N_39044,N_37602);
and U41525 (N_41525,N_37828,N_38057);
xnor U41526 (N_41526,N_39917,N_37537);
or U41527 (N_41527,N_37515,N_38780);
nor U41528 (N_41528,N_38691,N_37890);
nand U41529 (N_41529,N_39032,N_37762);
or U41530 (N_41530,N_37801,N_38138);
nand U41531 (N_41531,N_37807,N_39144);
or U41532 (N_41532,N_38725,N_38594);
nand U41533 (N_41533,N_38708,N_37817);
xnor U41534 (N_41534,N_39511,N_38098);
xnor U41535 (N_41535,N_37751,N_38817);
or U41536 (N_41536,N_38846,N_39948);
nor U41537 (N_41537,N_39245,N_39284);
nor U41538 (N_41538,N_39012,N_39492);
nand U41539 (N_41539,N_39563,N_39008);
nand U41540 (N_41540,N_38761,N_39495);
or U41541 (N_41541,N_37935,N_37857);
and U41542 (N_41542,N_38335,N_38784);
nor U41543 (N_41543,N_38378,N_38195);
nand U41544 (N_41544,N_39673,N_39099);
and U41545 (N_41545,N_38456,N_38419);
and U41546 (N_41546,N_39594,N_39648);
and U41547 (N_41547,N_38745,N_39529);
nand U41548 (N_41548,N_38805,N_39845);
nor U41549 (N_41549,N_38728,N_38111);
or U41550 (N_41550,N_37942,N_38913);
xor U41551 (N_41551,N_38604,N_37712);
nand U41552 (N_41552,N_38662,N_39454);
nor U41553 (N_41553,N_38142,N_37623);
nor U41554 (N_41554,N_38092,N_38965);
and U41555 (N_41555,N_37969,N_37920);
and U41556 (N_41556,N_39442,N_37660);
or U41557 (N_41557,N_38966,N_37762);
nor U41558 (N_41558,N_39359,N_38304);
or U41559 (N_41559,N_39727,N_38241);
nor U41560 (N_41560,N_37512,N_38072);
and U41561 (N_41561,N_38466,N_37574);
nor U41562 (N_41562,N_38442,N_38838);
and U41563 (N_41563,N_37564,N_38926);
nor U41564 (N_41564,N_37648,N_37569);
nand U41565 (N_41565,N_39422,N_37880);
nor U41566 (N_41566,N_39359,N_39266);
and U41567 (N_41567,N_38887,N_38198);
and U41568 (N_41568,N_39393,N_39188);
nor U41569 (N_41569,N_39481,N_38397);
nand U41570 (N_41570,N_38204,N_39743);
or U41571 (N_41571,N_39791,N_39710);
xor U41572 (N_41572,N_38444,N_37799);
nor U41573 (N_41573,N_39889,N_37893);
or U41574 (N_41574,N_38850,N_38898);
and U41575 (N_41575,N_38912,N_38320);
nand U41576 (N_41576,N_39103,N_39928);
nor U41577 (N_41577,N_37700,N_38544);
and U41578 (N_41578,N_39070,N_38928);
nand U41579 (N_41579,N_39422,N_38584);
and U41580 (N_41580,N_38912,N_38815);
nor U41581 (N_41581,N_39046,N_39997);
nor U41582 (N_41582,N_37783,N_39344);
or U41583 (N_41583,N_38218,N_37628);
and U41584 (N_41584,N_39554,N_37542);
nand U41585 (N_41585,N_37643,N_38655);
nor U41586 (N_41586,N_37932,N_39098);
and U41587 (N_41587,N_39557,N_37988);
nand U41588 (N_41588,N_39913,N_39932);
nand U41589 (N_41589,N_39551,N_39215);
and U41590 (N_41590,N_38219,N_38937);
nor U41591 (N_41591,N_38994,N_38117);
and U41592 (N_41592,N_38812,N_39522);
or U41593 (N_41593,N_39803,N_38084);
nor U41594 (N_41594,N_37671,N_39588);
or U41595 (N_41595,N_39396,N_39752);
and U41596 (N_41596,N_39736,N_38170);
nand U41597 (N_41597,N_38900,N_39193);
and U41598 (N_41598,N_39386,N_37547);
nand U41599 (N_41599,N_38048,N_39378);
nor U41600 (N_41600,N_37977,N_39045);
or U41601 (N_41601,N_38304,N_39286);
nor U41602 (N_41602,N_38331,N_38642);
and U41603 (N_41603,N_38393,N_38043);
and U41604 (N_41604,N_38690,N_38518);
or U41605 (N_41605,N_38082,N_39454);
and U41606 (N_41606,N_38329,N_38143);
nor U41607 (N_41607,N_39647,N_38575);
nor U41608 (N_41608,N_39482,N_39292);
and U41609 (N_41609,N_39014,N_39790);
nand U41610 (N_41610,N_38882,N_39760);
nand U41611 (N_41611,N_39829,N_38488);
nand U41612 (N_41612,N_38336,N_38745);
nor U41613 (N_41613,N_39351,N_38769);
and U41614 (N_41614,N_39370,N_38209);
nor U41615 (N_41615,N_37616,N_37976);
or U41616 (N_41616,N_39172,N_37660);
and U41617 (N_41617,N_38079,N_38628);
nor U41618 (N_41618,N_39270,N_39373);
or U41619 (N_41619,N_38406,N_37981);
or U41620 (N_41620,N_39722,N_37942);
and U41621 (N_41621,N_38581,N_39544);
nand U41622 (N_41622,N_39271,N_39711);
nand U41623 (N_41623,N_38083,N_39822);
nor U41624 (N_41624,N_39423,N_38504);
nand U41625 (N_41625,N_38159,N_39837);
or U41626 (N_41626,N_38414,N_38998);
nor U41627 (N_41627,N_39516,N_39870);
nand U41628 (N_41628,N_38996,N_38640);
xnor U41629 (N_41629,N_39274,N_38015);
xor U41630 (N_41630,N_39226,N_37930);
nand U41631 (N_41631,N_39984,N_37844);
nor U41632 (N_41632,N_39605,N_37830);
nor U41633 (N_41633,N_38030,N_39062);
and U41634 (N_41634,N_38304,N_39950);
and U41635 (N_41635,N_39500,N_38415);
or U41636 (N_41636,N_38893,N_38012);
and U41637 (N_41637,N_37885,N_38916);
xor U41638 (N_41638,N_38504,N_38155);
xor U41639 (N_41639,N_39989,N_38285);
nand U41640 (N_41640,N_39824,N_37731);
and U41641 (N_41641,N_37677,N_37974);
nand U41642 (N_41642,N_39552,N_37538);
or U41643 (N_41643,N_39582,N_39692);
xor U41644 (N_41644,N_38715,N_38261);
nand U41645 (N_41645,N_38562,N_38491);
or U41646 (N_41646,N_38228,N_38629);
nand U41647 (N_41647,N_39101,N_39783);
xnor U41648 (N_41648,N_39879,N_38182);
xor U41649 (N_41649,N_39763,N_37690);
xnor U41650 (N_41650,N_38040,N_39226);
and U41651 (N_41651,N_37951,N_37589);
nor U41652 (N_41652,N_37981,N_38687);
and U41653 (N_41653,N_38038,N_39796);
xnor U41654 (N_41654,N_38955,N_38627);
nand U41655 (N_41655,N_39706,N_38093);
and U41656 (N_41656,N_38376,N_37812);
nor U41657 (N_41657,N_38925,N_39514);
or U41658 (N_41658,N_39273,N_38106);
or U41659 (N_41659,N_39090,N_37607);
nand U41660 (N_41660,N_37526,N_39907);
and U41661 (N_41661,N_38573,N_37607);
nand U41662 (N_41662,N_37849,N_38614);
and U41663 (N_41663,N_38241,N_38125);
or U41664 (N_41664,N_37567,N_37578);
nand U41665 (N_41665,N_37700,N_38573);
nor U41666 (N_41666,N_39115,N_39192);
nor U41667 (N_41667,N_37577,N_38834);
nor U41668 (N_41668,N_37537,N_39103);
nand U41669 (N_41669,N_39440,N_38342);
or U41670 (N_41670,N_38072,N_37919);
nor U41671 (N_41671,N_39277,N_38721);
or U41672 (N_41672,N_38686,N_38354);
nand U41673 (N_41673,N_38632,N_39861);
or U41674 (N_41674,N_37545,N_38791);
nand U41675 (N_41675,N_39256,N_38939);
and U41676 (N_41676,N_38440,N_38352);
nand U41677 (N_41677,N_38214,N_38580);
and U41678 (N_41678,N_38739,N_38225);
or U41679 (N_41679,N_39148,N_37648);
xor U41680 (N_41680,N_39182,N_39917);
or U41681 (N_41681,N_39191,N_39743);
nand U41682 (N_41682,N_39039,N_38126);
nor U41683 (N_41683,N_38830,N_39001);
nor U41684 (N_41684,N_39327,N_39271);
nand U41685 (N_41685,N_39662,N_39665);
and U41686 (N_41686,N_39473,N_38753);
nor U41687 (N_41687,N_38312,N_38997);
or U41688 (N_41688,N_38054,N_37986);
or U41689 (N_41689,N_38632,N_38991);
nor U41690 (N_41690,N_38185,N_38796);
or U41691 (N_41691,N_39828,N_38222);
xor U41692 (N_41692,N_39356,N_38498);
nor U41693 (N_41693,N_38394,N_37726);
nor U41694 (N_41694,N_37802,N_39069);
xnor U41695 (N_41695,N_37659,N_38556);
xnor U41696 (N_41696,N_39539,N_38619);
or U41697 (N_41697,N_38095,N_39537);
or U41698 (N_41698,N_38487,N_37879);
or U41699 (N_41699,N_39310,N_38379);
nor U41700 (N_41700,N_37820,N_37753);
and U41701 (N_41701,N_38500,N_38076);
and U41702 (N_41702,N_39050,N_39599);
nor U41703 (N_41703,N_38612,N_39528);
or U41704 (N_41704,N_38035,N_38889);
and U41705 (N_41705,N_38603,N_37599);
nor U41706 (N_41706,N_39939,N_39304);
or U41707 (N_41707,N_38015,N_38544);
nand U41708 (N_41708,N_39673,N_39967);
nand U41709 (N_41709,N_38090,N_37671);
and U41710 (N_41710,N_37956,N_38728);
and U41711 (N_41711,N_38790,N_37876);
xnor U41712 (N_41712,N_39751,N_39986);
xor U41713 (N_41713,N_38874,N_39056);
xnor U41714 (N_41714,N_38947,N_37647);
nor U41715 (N_41715,N_37953,N_37765);
and U41716 (N_41716,N_39132,N_39303);
nand U41717 (N_41717,N_37556,N_39083);
or U41718 (N_41718,N_38233,N_37854);
or U41719 (N_41719,N_38413,N_39563);
nor U41720 (N_41720,N_39512,N_39033);
or U41721 (N_41721,N_39374,N_37665);
or U41722 (N_41722,N_38874,N_38297);
and U41723 (N_41723,N_38174,N_39054);
nand U41724 (N_41724,N_39584,N_38282);
and U41725 (N_41725,N_39382,N_39758);
and U41726 (N_41726,N_39633,N_38783);
or U41727 (N_41727,N_39727,N_39641);
nand U41728 (N_41728,N_39705,N_38232);
or U41729 (N_41729,N_39607,N_37692);
nand U41730 (N_41730,N_38684,N_39808);
nor U41731 (N_41731,N_38266,N_38715);
or U41732 (N_41732,N_38319,N_39781);
and U41733 (N_41733,N_39284,N_39890);
or U41734 (N_41734,N_39135,N_38823);
or U41735 (N_41735,N_38256,N_38048);
nand U41736 (N_41736,N_38126,N_37634);
nor U41737 (N_41737,N_39818,N_38417);
and U41738 (N_41738,N_38216,N_38684);
nand U41739 (N_41739,N_38590,N_37695);
xor U41740 (N_41740,N_37527,N_38008);
nand U41741 (N_41741,N_38426,N_37717);
or U41742 (N_41742,N_38299,N_39259);
nor U41743 (N_41743,N_37748,N_38101);
or U41744 (N_41744,N_38132,N_39598);
nand U41745 (N_41745,N_37696,N_38600);
nor U41746 (N_41746,N_38835,N_37956);
or U41747 (N_41747,N_39753,N_39561);
or U41748 (N_41748,N_38826,N_39601);
or U41749 (N_41749,N_39950,N_37721);
nand U41750 (N_41750,N_38097,N_39883);
or U41751 (N_41751,N_39690,N_38198);
nand U41752 (N_41752,N_37907,N_39747);
nand U41753 (N_41753,N_38031,N_38321);
and U41754 (N_41754,N_38600,N_37825);
and U41755 (N_41755,N_38977,N_39795);
and U41756 (N_41756,N_38181,N_38959);
nor U41757 (N_41757,N_39335,N_38743);
and U41758 (N_41758,N_37756,N_39843);
nand U41759 (N_41759,N_39197,N_37626);
and U41760 (N_41760,N_38156,N_37642);
nand U41761 (N_41761,N_37769,N_37886);
and U41762 (N_41762,N_38456,N_38185);
nor U41763 (N_41763,N_39760,N_39185);
nor U41764 (N_41764,N_37651,N_39482);
xor U41765 (N_41765,N_38303,N_38743);
nand U41766 (N_41766,N_39263,N_38660);
or U41767 (N_41767,N_37780,N_39168);
nor U41768 (N_41768,N_37507,N_39496);
nor U41769 (N_41769,N_39385,N_39287);
or U41770 (N_41770,N_38166,N_39924);
and U41771 (N_41771,N_39278,N_39090);
xnor U41772 (N_41772,N_37824,N_38865);
nor U41773 (N_41773,N_38043,N_38864);
and U41774 (N_41774,N_39200,N_37974);
nand U41775 (N_41775,N_37779,N_38085);
nand U41776 (N_41776,N_37870,N_39962);
and U41777 (N_41777,N_39963,N_39067);
nand U41778 (N_41778,N_38905,N_39269);
or U41779 (N_41779,N_39984,N_38486);
or U41780 (N_41780,N_38368,N_39762);
or U41781 (N_41781,N_39321,N_38152);
or U41782 (N_41782,N_38844,N_39309);
or U41783 (N_41783,N_39419,N_38315);
and U41784 (N_41784,N_39274,N_39593);
nor U41785 (N_41785,N_37644,N_39630);
and U41786 (N_41786,N_37601,N_38982);
and U41787 (N_41787,N_39727,N_38209);
nand U41788 (N_41788,N_39304,N_38050);
nor U41789 (N_41789,N_37993,N_38127);
nor U41790 (N_41790,N_37597,N_38374);
nor U41791 (N_41791,N_39660,N_38349);
nand U41792 (N_41792,N_39253,N_37847);
nor U41793 (N_41793,N_39151,N_38662);
nor U41794 (N_41794,N_38367,N_37700);
nor U41795 (N_41795,N_38627,N_37827);
xnor U41796 (N_41796,N_39068,N_39800);
nand U41797 (N_41797,N_39730,N_39535);
nor U41798 (N_41798,N_38701,N_38502);
and U41799 (N_41799,N_39828,N_39586);
nand U41800 (N_41800,N_39129,N_37530);
or U41801 (N_41801,N_39853,N_38269);
nand U41802 (N_41802,N_39951,N_39189);
xnor U41803 (N_41803,N_38277,N_38865);
nor U41804 (N_41804,N_38892,N_38325);
and U41805 (N_41805,N_37882,N_38619);
or U41806 (N_41806,N_37536,N_39194);
and U41807 (N_41807,N_38725,N_37808);
or U41808 (N_41808,N_39881,N_38766);
or U41809 (N_41809,N_39248,N_38007);
or U41810 (N_41810,N_39846,N_39839);
or U41811 (N_41811,N_38584,N_38543);
xnor U41812 (N_41812,N_38779,N_39733);
nand U41813 (N_41813,N_39897,N_39884);
or U41814 (N_41814,N_38300,N_38791);
and U41815 (N_41815,N_39136,N_38229);
nor U41816 (N_41816,N_37625,N_38902);
xor U41817 (N_41817,N_39137,N_38872);
and U41818 (N_41818,N_38528,N_38028);
and U41819 (N_41819,N_37733,N_39111);
or U41820 (N_41820,N_38716,N_37915);
nand U41821 (N_41821,N_39493,N_37962);
and U41822 (N_41822,N_39827,N_39920);
or U41823 (N_41823,N_39444,N_38519);
nor U41824 (N_41824,N_39487,N_39147);
xor U41825 (N_41825,N_38660,N_38157);
and U41826 (N_41826,N_37717,N_39194);
or U41827 (N_41827,N_38071,N_39843);
nand U41828 (N_41828,N_39081,N_39486);
nor U41829 (N_41829,N_37976,N_39717);
and U41830 (N_41830,N_39840,N_38851);
nor U41831 (N_41831,N_37504,N_37811);
nor U41832 (N_41832,N_39444,N_37549);
nand U41833 (N_41833,N_39133,N_39534);
or U41834 (N_41834,N_37766,N_39565);
and U41835 (N_41835,N_38898,N_38425);
nand U41836 (N_41836,N_38799,N_39742);
or U41837 (N_41837,N_37634,N_37735);
nand U41838 (N_41838,N_38893,N_38689);
and U41839 (N_41839,N_39703,N_38544);
nand U41840 (N_41840,N_37690,N_38078);
nand U41841 (N_41841,N_38328,N_38421);
or U41842 (N_41842,N_37557,N_39661);
nor U41843 (N_41843,N_37878,N_38737);
and U41844 (N_41844,N_39290,N_38515);
and U41845 (N_41845,N_38211,N_38857);
nand U41846 (N_41846,N_38069,N_39067);
nand U41847 (N_41847,N_38294,N_39535);
and U41848 (N_41848,N_38603,N_39352);
nor U41849 (N_41849,N_38267,N_38812);
nor U41850 (N_41850,N_37602,N_39562);
and U41851 (N_41851,N_39300,N_39211);
or U41852 (N_41852,N_38603,N_39921);
and U41853 (N_41853,N_37666,N_38340);
or U41854 (N_41854,N_38082,N_38414);
and U41855 (N_41855,N_39490,N_39731);
xnor U41856 (N_41856,N_39029,N_39693);
and U41857 (N_41857,N_38012,N_38268);
nand U41858 (N_41858,N_37803,N_38685);
xnor U41859 (N_41859,N_39700,N_39936);
and U41860 (N_41860,N_38992,N_37573);
and U41861 (N_41861,N_37880,N_39075);
or U41862 (N_41862,N_39409,N_38669);
nand U41863 (N_41863,N_38068,N_39202);
and U41864 (N_41864,N_37635,N_38751);
and U41865 (N_41865,N_38023,N_38056);
or U41866 (N_41866,N_39922,N_39828);
or U41867 (N_41867,N_38071,N_38618);
nor U41868 (N_41868,N_39227,N_37620);
and U41869 (N_41869,N_38877,N_38303);
xnor U41870 (N_41870,N_37513,N_38449);
xnor U41871 (N_41871,N_38015,N_38552);
or U41872 (N_41872,N_37747,N_38355);
nand U41873 (N_41873,N_37860,N_39739);
nand U41874 (N_41874,N_39691,N_38866);
xor U41875 (N_41875,N_38220,N_39404);
or U41876 (N_41876,N_39315,N_39797);
nor U41877 (N_41877,N_37542,N_39422);
nor U41878 (N_41878,N_38637,N_39016);
nor U41879 (N_41879,N_39119,N_38718);
nor U41880 (N_41880,N_39052,N_39220);
nand U41881 (N_41881,N_39892,N_38798);
nor U41882 (N_41882,N_37661,N_39694);
and U41883 (N_41883,N_37990,N_39446);
nor U41884 (N_41884,N_38407,N_39362);
nor U41885 (N_41885,N_39005,N_37984);
nand U41886 (N_41886,N_38043,N_39014);
nor U41887 (N_41887,N_38662,N_38811);
nand U41888 (N_41888,N_38289,N_37610);
and U41889 (N_41889,N_39985,N_39830);
nor U41890 (N_41890,N_38412,N_38854);
or U41891 (N_41891,N_38261,N_38476);
nand U41892 (N_41892,N_39014,N_37785);
nand U41893 (N_41893,N_38078,N_39164);
and U41894 (N_41894,N_38462,N_38965);
or U41895 (N_41895,N_38349,N_39088);
and U41896 (N_41896,N_39543,N_39402);
and U41897 (N_41897,N_38482,N_39132);
nor U41898 (N_41898,N_39921,N_39404);
nand U41899 (N_41899,N_38770,N_38778);
nand U41900 (N_41900,N_38027,N_39263);
nand U41901 (N_41901,N_37886,N_39039);
and U41902 (N_41902,N_39938,N_39389);
or U41903 (N_41903,N_39245,N_38688);
and U41904 (N_41904,N_38606,N_39007);
xnor U41905 (N_41905,N_37993,N_38838);
or U41906 (N_41906,N_38357,N_39222);
and U41907 (N_41907,N_39310,N_37949);
or U41908 (N_41908,N_38223,N_39392);
nand U41909 (N_41909,N_37885,N_38243);
or U41910 (N_41910,N_38426,N_37639);
nor U41911 (N_41911,N_39673,N_38212);
nand U41912 (N_41912,N_39632,N_38584);
nor U41913 (N_41913,N_39941,N_38547);
nand U41914 (N_41914,N_39893,N_39416);
or U41915 (N_41915,N_38323,N_39588);
xor U41916 (N_41916,N_39822,N_37818);
nand U41917 (N_41917,N_37787,N_38500);
or U41918 (N_41918,N_39832,N_37564);
nand U41919 (N_41919,N_39544,N_39673);
nor U41920 (N_41920,N_39761,N_38475);
nand U41921 (N_41921,N_37681,N_38660);
nor U41922 (N_41922,N_39057,N_39990);
xor U41923 (N_41923,N_38565,N_37778);
and U41924 (N_41924,N_38940,N_39181);
nand U41925 (N_41925,N_39690,N_38150);
and U41926 (N_41926,N_39728,N_38428);
nor U41927 (N_41927,N_38869,N_38203);
nor U41928 (N_41928,N_38737,N_39071);
nand U41929 (N_41929,N_38408,N_39887);
and U41930 (N_41930,N_38081,N_37673);
and U41931 (N_41931,N_39257,N_37523);
and U41932 (N_41932,N_38117,N_39765);
and U41933 (N_41933,N_39778,N_38187);
nand U41934 (N_41934,N_37727,N_38747);
nand U41935 (N_41935,N_38992,N_37690);
and U41936 (N_41936,N_38060,N_38309);
nor U41937 (N_41937,N_38946,N_38789);
nor U41938 (N_41938,N_37507,N_39292);
and U41939 (N_41939,N_37997,N_39080);
nand U41940 (N_41940,N_39839,N_37557);
xor U41941 (N_41941,N_37526,N_39479);
and U41942 (N_41942,N_38832,N_38886);
nand U41943 (N_41943,N_38478,N_39559);
or U41944 (N_41944,N_38610,N_38456);
nand U41945 (N_41945,N_37534,N_37915);
nor U41946 (N_41946,N_38688,N_38618);
nor U41947 (N_41947,N_37843,N_39790);
nor U41948 (N_41948,N_38629,N_39826);
or U41949 (N_41949,N_38649,N_37864);
or U41950 (N_41950,N_37577,N_39196);
nor U41951 (N_41951,N_38955,N_38750);
nand U41952 (N_41952,N_39956,N_39293);
and U41953 (N_41953,N_38280,N_38811);
nand U41954 (N_41954,N_37634,N_39544);
and U41955 (N_41955,N_38774,N_38170);
or U41956 (N_41956,N_39219,N_38609);
xor U41957 (N_41957,N_39879,N_37532);
or U41958 (N_41958,N_39690,N_37582);
nor U41959 (N_41959,N_38775,N_37516);
xnor U41960 (N_41960,N_38392,N_39424);
nand U41961 (N_41961,N_38883,N_39889);
or U41962 (N_41962,N_37587,N_37739);
nor U41963 (N_41963,N_38830,N_39267);
nor U41964 (N_41964,N_38797,N_39887);
or U41965 (N_41965,N_39686,N_37766);
and U41966 (N_41966,N_38249,N_39110);
or U41967 (N_41967,N_37651,N_38450);
or U41968 (N_41968,N_39006,N_38256);
xor U41969 (N_41969,N_38110,N_39728);
xor U41970 (N_41970,N_38993,N_38976);
and U41971 (N_41971,N_39463,N_38346);
nand U41972 (N_41972,N_38122,N_39249);
nor U41973 (N_41973,N_39988,N_39683);
or U41974 (N_41974,N_39184,N_37504);
or U41975 (N_41975,N_37788,N_38926);
or U41976 (N_41976,N_38629,N_38481);
nand U41977 (N_41977,N_39583,N_38232);
nor U41978 (N_41978,N_37861,N_39805);
or U41979 (N_41979,N_38178,N_38323);
nand U41980 (N_41980,N_38145,N_39077);
xor U41981 (N_41981,N_39412,N_39161);
xor U41982 (N_41982,N_38021,N_39841);
nor U41983 (N_41983,N_38851,N_37722);
and U41984 (N_41984,N_37780,N_38259);
or U41985 (N_41985,N_39831,N_37515);
nand U41986 (N_41986,N_39777,N_39586);
or U41987 (N_41987,N_39340,N_38237);
and U41988 (N_41988,N_38322,N_39770);
and U41989 (N_41989,N_37613,N_38487);
and U41990 (N_41990,N_38044,N_38092);
or U41991 (N_41991,N_39134,N_39131);
and U41992 (N_41992,N_38459,N_38952);
nor U41993 (N_41993,N_39378,N_39456);
and U41994 (N_41994,N_39449,N_38205);
nor U41995 (N_41995,N_39629,N_39055);
and U41996 (N_41996,N_39784,N_39398);
or U41997 (N_41997,N_39402,N_38337);
xnor U41998 (N_41998,N_38895,N_37666);
nor U41999 (N_41999,N_39099,N_39024);
xnor U42000 (N_42000,N_37888,N_38232);
xor U42001 (N_42001,N_38808,N_39755);
nor U42002 (N_42002,N_37857,N_38820);
and U42003 (N_42003,N_37689,N_39622);
and U42004 (N_42004,N_37873,N_39498);
and U42005 (N_42005,N_38708,N_38385);
nor U42006 (N_42006,N_38060,N_38086);
and U42007 (N_42007,N_38769,N_39260);
and U42008 (N_42008,N_38541,N_37618);
nor U42009 (N_42009,N_39203,N_38896);
or U42010 (N_42010,N_38820,N_39241);
or U42011 (N_42011,N_38134,N_39013);
nand U42012 (N_42012,N_37786,N_39083);
nand U42013 (N_42013,N_38209,N_38967);
and U42014 (N_42014,N_38794,N_38936);
or U42015 (N_42015,N_38404,N_38556);
or U42016 (N_42016,N_39256,N_39097);
nand U42017 (N_42017,N_37647,N_38133);
xnor U42018 (N_42018,N_39400,N_38912);
nand U42019 (N_42019,N_39107,N_39822);
or U42020 (N_42020,N_39988,N_38341);
nor U42021 (N_42021,N_38846,N_38668);
and U42022 (N_42022,N_39920,N_37815);
nor U42023 (N_42023,N_39411,N_38257);
nand U42024 (N_42024,N_38944,N_38196);
and U42025 (N_42025,N_37627,N_38441);
nand U42026 (N_42026,N_38031,N_39612);
nor U42027 (N_42027,N_37635,N_37822);
nand U42028 (N_42028,N_37682,N_38983);
or U42029 (N_42029,N_38652,N_38670);
nand U42030 (N_42030,N_38257,N_37794);
nor U42031 (N_42031,N_38854,N_37758);
and U42032 (N_42032,N_39564,N_39500);
nor U42033 (N_42033,N_39765,N_38908);
or U42034 (N_42034,N_38275,N_39250);
xor U42035 (N_42035,N_38506,N_38765);
nor U42036 (N_42036,N_37729,N_39672);
and U42037 (N_42037,N_39541,N_39316);
nor U42038 (N_42038,N_38152,N_39873);
or U42039 (N_42039,N_39011,N_38024);
nor U42040 (N_42040,N_39624,N_37877);
nand U42041 (N_42041,N_37604,N_37782);
xor U42042 (N_42042,N_37544,N_38881);
or U42043 (N_42043,N_39407,N_37610);
xor U42044 (N_42044,N_38900,N_37854);
nand U42045 (N_42045,N_39540,N_38314);
and U42046 (N_42046,N_38600,N_39213);
nor U42047 (N_42047,N_37791,N_39248);
nor U42048 (N_42048,N_38414,N_38086);
or U42049 (N_42049,N_39159,N_38096);
nand U42050 (N_42050,N_37835,N_38589);
nand U42051 (N_42051,N_39541,N_39206);
xnor U42052 (N_42052,N_38905,N_37676);
and U42053 (N_42053,N_38275,N_38775);
nor U42054 (N_42054,N_39456,N_38289);
nor U42055 (N_42055,N_38684,N_38310);
nand U42056 (N_42056,N_39338,N_39451);
and U42057 (N_42057,N_39914,N_37901);
or U42058 (N_42058,N_37950,N_38223);
or U42059 (N_42059,N_39730,N_39867);
nor U42060 (N_42060,N_39133,N_37866);
xnor U42061 (N_42061,N_37541,N_37545);
xor U42062 (N_42062,N_39861,N_37770);
and U42063 (N_42063,N_39592,N_38000);
nor U42064 (N_42064,N_38500,N_39302);
xnor U42065 (N_42065,N_38898,N_39852);
nand U42066 (N_42066,N_39791,N_37583);
nand U42067 (N_42067,N_38418,N_37853);
nor U42068 (N_42068,N_37904,N_38022);
or U42069 (N_42069,N_39567,N_39007);
and U42070 (N_42070,N_38297,N_38275);
xor U42071 (N_42071,N_38977,N_38695);
nand U42072 (N_42072,N_39778,N_39831);
or U42073 (N_42073,N_39346,N_39296);
and U42074 (N_42074,N_37750,N_38069);
nor U42075 (N_42075,N_39427,N_37547);
and U42076 (N_42076,N_39371,N_39504);
or U42077 (N_42077,N_37534,N_38248);
nand U42078 (N_42078,N_37531,N_39076);
or U42079 (N_42079,N_38061,N_37785);
nand U42080 (N_42080,N_39605,N_38286);
and U42081 (N_42081,N_38440,N_39713);
xor U42082 (N_42082,N_38813,N_39447);
xor U42083 (N_42083,N_39894,N_39165);
xor U42084 (N_42084,N_39020,N_38169);
or U42085 (N_42085,N_37812,N_39519);
nand U42086 (N_42086,N_39278,N_38916);
xnor U42087 (N_42087,N_38217,N_38461);
or U42088 (N_42088,N_38721,N_38557);
or U42089 (N_42089,N_37647,N_39776);
and U42090 (N_42090,N_38994,N_39459);
nand U42091 (N_42091,N_38851,N_39617);
nand U42092 (N_42092,N_37965,N_38662);
xnor U42093 (N_42093,N_38753,N_37992);
and U42094 (N_42094,N_38595,N_37535);
nor U42095 (N_42095,N_38071,N_38907);
nand U42096 (N_42096,N_39730,N_38878);
nand U42097 (N_42097,N_37556,N_37602);
and U42098 (N_42098,N_38850,N_38770);
nor U42099 (N_42099,N_38459,N_39775);
nor U42100 (N_42100,N_39769,N_38800);
and U42101 (N_42101,N_38163,N_38461);
nand U42102 (N_42102,N_37663,N_39102);
nor U42103 (N_42103,N_39331,N_39195);
and U42104 (N_42104,N_39282,N_38910);
nand U42105 (N_42105,N_38532,N_39086);
xnor U42106 (N_42106,N_38709,N_39341);
or U42107 (N_42107,N_37618,N_39550);
nand U42108 (N_42108,N_37637,N_39368);
and U42109 (N_42109,N_38334,N_39622);
nand U42110 (N_42110,N_38027,N_39708);
xor U42111 (N_42111,N_39187,N_37960);
nand U42112 (N_42112,N_39789,N_39398);
and U42113 (N_42113,N_39276,N_39083);
nand U42114 (N_42114,N_39339,N_39843);
xnor U42115 (N_42115,N_39772,N_38786);
nand U42116 (N_42116,N_39685,N_39298);
nand U42117 (N_42117,N_39049,N_37928);
or U42118 (N_42118,N_39202,N_39624);
nor U42119 (N_42119,N_38492,N_39752);
nor U42120 (N_42120,N_37814,N_39232);
nor U42121 (N_42121,N_38707,N_39357);
nand U42122 (N_42122,N_38654,N_37854);
and U42123 (N_42123,N_39942,N_39526);
nand U42124 (N_42124,N_39743,N_38623);
or U42125 (N_42125,N_39385,N_39312);
or U42126 (N_42126,N_39563,N_37721);
and U42127 (N_42127,N_39421,N_39492);
nor U42128 (N_42128,N_37573,N_37853);
nor U42129 (N_42129,N_38026,N_39606);
nand U42130 (N_42130,N_38792,N_38639);
nand U42131 (N_42131,N_38993,N_39222);
or U42132 (N_42132,N_38728,N_39248);
or U42133 (N_42133,N_39142,N_39888);
and U42134 (N_42134,N_39220,N_39281);
and U42135 (N_42135,N_39898,N_39797);
and U42136 (N_42136,N_39235,N_38805);
and U42137 (N_42137,N_38940,N_39844);
and U42138 (N_42138,N_38987,N_38497);
xor U42139 (N_42139,N_37938,N_37524);
and U42140 (N_42140,N_38731,N_37609);
nand U42141 (N_42141,N_39539,N_38496);
xnor U42142 (N_42142,N_37956,N_38760);
or U42143 (N_42143,N_39523,N_39599);
nor U42144 (N_42144,N_39486,N_39549);
or U42145 (N_42145,N_38446,N_38725);
or U42146 (N_42146,N_39418,N_38143);
nor U42147 (N_42147,N_38388,N_39567);
and U42148 (N_42148,N_39334,N_37683);
nand U42149 (N_42149,N_37782,N_38871);
nor U42150 (N_42150,N_38402,N_37907);
nand U42151 (N_42151,N_39799,N_38067);
or U42152 (N_42152,N_37566,N_39298);
nor U42153 (N_42153,N_38633,N_38115);
nor U42154 (N_42154,N_38934,N_38857);
or U42155 (N_42155,N_39167,N_38995);
xor U42156 (N_42156,N_38296,N_38498);
nor U42157 (N_42157,N_37657,N_38934);
xnor U42158 (N_42158,N_39627,N_39946);
and U42159 (N_42159,N_39299,N_38983);
xor U42160 (N_42160,N_39975,N_39630);
and U42161 (N_42161,N_38967,N_38853);
xor U42162 (N_42162,N_38301,N_38578);
and U42163 (N_42163,N_39871,N_39836);
nand U42164 (N_42164,N_39459,N_38009);
xor U42165 (N_42165,N_38478,N_39928);
and U42166 (N_42166,N_38630,N_37731);
or U42167 (N_42167,N_39924,N_37574);
or U42168 (N_42168,N_38269,N_38033);
and U42169 (N_42169,N_39041,N_37726);
xnor U42170 (N_42170,N_39127,N_39645);
xor U42171 (N_42171,N_37660,N_38395);
xnor U42172 (N_42172,N_39482,N_38755);
nand U42173 (N_42173,N_38374,N_39573);
nand U42174 (N_42174,N_39231,N_39621);
nand U42175 (N_42175,N_37620,N_38005);
or U42176 (N_42176,N_38716,N_38984);
nand U42177 (N_42177,N_37888,N_37767);
nor U42178 (N_42178,N_39106,N_39073);
nand U42179 (N_42179,N_37766,N_37668);
nor U42180 (N_42180,N_38358,N_37636);
nor U42181 (N_42181,N_39284,N_38585);
nor U42182 (N_42182,N_39734,N_38727);
nor U42183 (N_42183,N_38564,N_39938);
or U42184 (N_42184,N_38181,N_37707);
nand U42185 (N_42185,N_39229,N_38444);
and U42186 (N_42186,N_37832,N_38913);
or U42187 (N_42187,N_37551,N_39410);
or U42188 (N_42188,N_38221,N_37896);
or U42189 (N_42189,N_39458,N_39903);
and U42190 (N_42190,N_39164,N_38128);
and U42191 (N_42191,N_38242,N_38381);
nor U42192 (N_42192,N_38428,N_39082);
and U42193 (N_42193,N_38075,N_39071);
nand U42194 (N_42194,N_38486,N_37624);
nand U42195 (N_42195,N_38501,N_39015);
nor U42196 (N_42196,N_38576,N_39368);
or U42197 (N_42197,N_39020,N_39079);
and U42198 (N_42198,N_37606,N_37540);
or U42199 (N_42199,N_39451,N_38317);
xnor U42200 (N_42200,N_37643,N_39293);
nor U42201 (N_42201,N_38327,N_39167);
and U42202 (N_42202,N_38476,N_39204);
and U42203 (N_42203,N_38597,N_38995);
and U42204 (N_42204,N_39135,N_38484);
nand U42205 (N_42205,N_39400,N_38801);
xor U42206 (N_42206,N_39132,N_39158);
and U42207 (N_42207,N_38747,N_37762);
nand U42208 (N_42208,N_38876,N_38705);
and U42209 (N_42209,N_37713,N_37687);
nor U42210 (N_42210,N_38397,N_37882);
nand U42211 (N_42211,N_39372,N_39207);
and U42212 (N_42212,N_39483,N_39411);
and U42213 (N_42213,N_37749,N_37935);
nor U42214 (N_42214,N_39874,N_39031);
and U42215 (N_42215,N_39297,N_38503);
or U42216 (N_42216,N_37963,N_37629);
nor U42217 (N_42217,N_38952,N_39972);
xor U42218 (N_42218,N_37938,N_37926);
or U42219 (N_42219,N_37923,N_37921);
or U42220 (N_42220,N_38040,N_39293);
nand U42221 (N_42221,N_37703,N_38807);
xnor U42222 (N_42222,N_39832,N_38304);
nor U42223 (N_42223,N_38899,N_39184);
nor U42224 (N_42224,N_38960,N_38404);
nand U42225 (N_42225,N_39553,N_37950);
nand U42226 (N_42226,N_39452,N_38287);
nor U42227 (N_42227,N_39527,N_39304);
and U42228 (N_42228,N_38016,N_37500);
xnor U42229 (N_42229,N_39997,N_39679);
or U42230 (N_42230,N_37653,N_39881);
xnor U42231 (N_42231,N_38492,N_39242);
nand U42232 (N_42232,N_38041,N_39708);
or U42233 (N_42233,N_39463,N_37737);
nand U42234 (N_42234,N_38315,N_39869);
or U42235 (N_42235,N_38562,N_39826);
or U42236 (N_42236,N_37777,N_39885);
nor U42237 (N_42237,N_38543,N_39972);
nand U42238 (N_42238,N_38447,N_39985);
nor U42239 (N_42239,N_39127,N_37914);
nand U42240 (N_42240,N_39310,N_39927);
nand U42241 (N_42241,N_37688,N_39413);
nor U42242 (N_42242,N_37888,N_38260);
and U42243 (N_42243,N_38574,N_37854);
or U42244 (N_42244,N_39352,N_37796);
or U42245 (N_42245,N_38815,N_39087);
nand U42246 (N_42246,N_38765,N_39234);
nor U42247 (N_42247,N_37868,N_38232);
nor U42248 (N_42248,N_39195,N_37623);
xnor U42249 (N_42249,N_37504,N_39371);
nor U42250 (N_42250,N_38738,N_39371);
or U42251 (N_42251,N_38053,N_39569);
nor U42252 (N_42252,N_38517,N_38958);
and U42253 (N_42253,N_38526,N_39575);
and U42254 (N_42254,N_39687,N_39891);
nand U42255 (N_42255,N_38342,N_38965);
nand U42256 (N_42256,N_39064,N_39160);
or U42257 (N_42257,N_37622,N_38348);
nand U42258 (N_42258,N_37834,N_39921);
and U42259 (N_42259,N_39554,N_39569);
nand U42260 (N_42260,N_37971,N_38981);
nor U42261 (N_42261,N_39804,N_39677);
nand U42262 (N_42262,N_39192,N_39382);
and U42263 (N_42263,N_37932,N_39020);
and U42264 (N_42264,N_38944,N_39934);
or U42265 (N_42265,N_37761,N_38044);
or U42266 (N_42266,N_37799,N_38490);
and U42267 (N_42267,N_38169,N_39436);
or U42268 (N_42268,N_37913,N_39677);
nor U42269 (N_42269,N_37967,N_39517);
and U42270 (N_42270,N_39044,N_38112);
and U42271 (N_42271,N_37912,N_39160);
or U42272 (N_42272,N_39861,N_37968);
and U42273 (N_42273,N_38296,N_38150);
nand U42274 (N_42274,N_37721,N_38972);
nor U42275 (N_42275,N_37820,N_39085);
and U42276 (N_42276,N_37695,N_38277);
and U42277 (N_42277,N_39865,N_39610);
or U42278 (N_42278,N_38934,N_39994);
nor U42279 (N_42279,N_38540,N_39090);
nor U42280 (N_42280,N_37522,N_39556);
or U42281 (N_42281,N_38614,N_39854);
nor U42282 (N_42282,N_38934,N_38036);
nand U42283 (N_42283,N_38962,N_37515);
or U42284 (N_42284,N_37792,N_37921);
nor U42285 (N_42285,N_38608,N_39823);
and U42286 (N_42286,N_39943,N_39851);
and U42287 (N_42287,N_38309,N_39018);
or U42288 (N_42288,N_38146,N_39492);
nor U42289 (N_42289,N_38641,N_38300);
or U42290 (N_42290,N_38199,N_39268);
nor U42291 (N_42291,N_39900,N_39042);
nor U42292 (N_42292,N_39186,N_39921);
nor U42293 (N_42293,N_38809,N_38129);
and U42294 (N_42294,N_39687,N_38492);
or U42295 (N_42295,N_37991,N_37889);
nor U42296 (N_42296,N_39987,N_39798);
nand U42297 (N_42297,N_38037,N_38798);
nand U42298 (N_42298,N_39370,N_39196);
and U42299 (N_42299,N_38913,N_38457);
nand U42300 (N_42300,N_38581,N_39779);
nand U42301 (N_42301,N_38113,N_38881);
nand U42302 (N_42302,N_39184,N_39550);
nand U42303 (N_42303,N_37910,N_37855);
or U42304 (N_42304,N_38145,N_39360);
xor U42305 (N_42305,N_38271,N_39924);
nand U42306 (N_42306,N_38312,N_37662);
nand U42307 (N_42307,N_39815,N_38745);
and U42308 (N_42308,N_38113,N_39804);
nand U42309 (N_42309,N_37571,N_39830);
xor U42310 (N_42310,N_38385,N_39236);
and U42311 (N_42311,N_37517,N_38197);
nand U42312 (N_42312,N_39144,N_37549);
nand U42313 (N_42313,N_39696,N_38699);
nand U42314 (N_42314,N_38011,N_39940);
and U42315 (N_42315,N_39323,N_37931);
or U42316 (N_42316,N_39889,N_38705);
and U42317 (N_42317,N_38683,N_38028);
and U42318 (N_42318,N_38155,N_37848);
or U42319 (N_42319,N_38626,N_39831);
nand U42320 (N_42320,N_38129,N_37731);
nand U42321 (N_42321,N_38897,N_38068);
xnor U42322 (N_42322,N_38430,N_38407);
nor U42323 (N_42323,N_38198,N_38498);
nor U42324 (N_42324,N_39950,N_38294);
nand U42325 (N_42325,N_38432,N_37560);
or U42326 (N_42326,N_37799,N_38329);
nand U42327 (N_42327,N_39479,N_37734);
nand U42328 (N_42328,N_38503,N_37660);
or U42329 (N_42329,N_37708,N_37669);
nand U42330 (N_42330,N_37827,N_39184);
or U42331 (N_42331,N_39260,N_39805);
nand U42332 (N_42332,N_38905,N_38309);
and U42333 (N_42333,N_39970,N_37516);
xnor U42334 (N_42334,N_39869,N_38199);
nor U42335 (N_42335,N_38893,N_38725);
or U42336 (N_42336,N_39183,N_38677);
and U42337 (N_42337,N_37543,N_37914);
nand U42338 (N_42338,N_37566,N_38104);
and U42339 (N_42339,N_38254,N_38159);
nand U42340 (N_42340,N_37656,N_38291);
or U42341 (N_42341,N_38718,N_39137);
or U42342 (N_42342,N_39001,N_39162);
nor U42343 (N_42343,N_38171,N_37887);
and U42344 (N_42344,N_37790,N_38297);
nand U42345 (N_42345,N_38794,N_38190);
nand U42346 (N_42346,N_39741,N_39917);
nor U42347 (N_42347,N_39389,N_38388);
nand U42348 (N_42348,N_39598,N_39993);
xnor U42349 (N_42349,N_37685,N_38770);
or U42350 (N_42350,N_38700,N_38150);
or U42351 (N_42351,N_37867,N_37998);
nand U42352 (N_42352,N_39912,N_38973);
or U42353 (N_42353,N_38863,N_38168);
nand U42354 (N_42354,N_37638,N_39149);
xor U42355 (N_42355,N_37666,N_38232);
and U42356 (N_42356,N_39270,N_39376);
nor U42357 (N_42357,N_39439,N_38875);
or U42358 (N_42358,N_38551,N_39061);
nor U42359 (N_42359,N_38296,N_39544);
nor U42360 (N_42360,N_37976,N_37661);
or U42361 (N_42361,N_39093,N_38697);
and U42362 (N_42362,N_38851,N_38769);
xnor U42363 (N_42363,N_37850,N_38667);
or U42364 (N_42364,N_39058,N_39939);
or U42365 (N_42365,N_39659,N_39185);
nor U42366 (N_42366,N_39025,N_38479);
xor U42367 (N_42367,N_39743,N_37763);
or U42368 (N_42368,N_37524,N_37671);
and U42369 (N_42369,N_39391,N_39481);
nand U42370 (N_42370,N_38560,N_38326);
and U42371 (N_42371,N_39970,N_39250);
xor U42372 (N_42372,N_39542,N_38128);
and U42373 (N_42373,N_38058,N_37699);
nor U42374 (N_42374,N_39015,N_38998);
xor U42375 (N_42375,N_39521,N_38872);
nor U42376 (N_42376,N_38562,N_38944);
nand U42377 (N_42377,N_39882,N_39864);
or U42378 (N_42378,N_38398,N_37936);
nand U42379 (N_42379,N_37538,N_38615);
and U42380 (N_42380,N_38505,N_38602);
xor U42381 (N_42381,N_39785,N_37720);
nor U42382 (N_42382,N_39863,N_38008);
or U42383 (N_42383,N_39391,N_37824);
nor U42384 (N_42384,N_39259,N_38506);
or U42385 (N_42385,N_39129,N_37911);
or U42386 (N_42386,N_38822,N_37892);
nor U42387 (N_42387,N_38355,N_38155);
and U42388 (N_42388,N_37713,N_39367);
and U42389 (N_42389,N_38878,N_39412);
nor U42390 (N_42390,N_37646,N_39642);
nor U42391 (N_42391,N_37604,N_38753);
nor U42392 (N_42392,N_39027,N_38738);
and U42393 (N_42393,N_39476,N_39196);
or U42394 (N_42394,N_38167,N_38416);
xor U42395 (N_42395,N_37945,N_39554);
and U42396 (N_42396,N_39500,N_38636);
nor U42397 (N_42397,N_39520,N_39438);
nand U42398 (N_42398,N_38807,N_38863);
or U42399 (N_42399,N_39048,N_38779);
and U42400 (N_42400,N_37995,N_39820);
or U42401 (N_42401,N_38015,N_38441);
or U42402 (N_42402,N_37669,N_38035);
or U42403 (N_42403,N_38289,N_39907);
nor U42404 (N_42404,N_38047,N_37731);
and U42405 (N_42405,N_39401,N_38791);
and U42406 (N_42406,N_38595,N_38342);
nand U42407 (N_42407,N_38405,N_39521);
and U42408 (N_42408,N_39063,N_38288);
nand U42409 (N_42409,N_39614,N_38650);
nor U42410 (N_42410,N_39082,N_37701);
nor U42411 (N_42411,N_38337,N_39778);
nand U42412 (N_42412,N_39142,N_39486);
nand U42413 (N_42413,N_37810,N_39071);
nor U42414 (N_42414,N_39192,N_37740);
or U42415 (N_42415,N_39246,N_39405);
or U42416 (N_42416,N_39758,N_39293);
or U42417 (N_42417,N_37968,N_38808);
or U42418 (N_42418,N_38447,N_38012);
xnor U42419 (N_42419,N_39152,N_37695);
xor U42420 (N_42420,N_38012,N_38763);
xor U42421 (N_42421,N_39235,N_39365);
or U42422 (N_42422,N_39182,N_39463);
nand U42423 (N_42423,N_38352,N_39116);
nor U42424 (N_42424,N_38420,N_37857);
and U42425 (N_42425,N_38076,N_37827);
xor U42426 (N_42426,N_37757,N_39473);
or U42427 (N_42427,N_39084,N_38539);
or U42428 (N_42428,N_38782,N_38440);
nor U42429 (N_42429,N_37517,N_39766);
or U42430 (N_42430,N_38743,N_38893);
xor U42431 (N_42431,N_38861,N_39638);
nand U42432 (N_42432,N_39256,N_39185);
or U42433 (N_42433,N_37549,N_37572);
nand U42434 (N_42434,N_39225,N_38181);
and U42435 (N_42435,N_39402,N_39624);
xor U42436 (N_42436,N_38563,N_38368);
or U42437 (N_42437,N_39385,N_38017);
and U42438 (N_42438,N_38772,N_37576);
nor U42439 (N_42439,N_39904,N_38443);
nand U42440 (N_42440,N_39485,N_38869);
nor U42441 (N_42441,N_37602,N_37537);
and U42442 (N_42442,N_39550,N_38325);
and U42443 (N_42443,N_37693,N_39266);
nand U42444 (N_42444,N_38651,N_37752);
nand U42445 (N_42445,N_39498,N_39299);
xnor U42446 (N_42446,N_39995,N_39156);
or U42447 (N_42447,N_39632,N_38434);
nor U42448 (N_42448,N_38477,N_38278);
nor U42449 (N_42449,N_38896,N_39964);
and U42450 (N_42450,N_38451,N_38340);
or U42451 (N_42451,N_37573,N_39491);
and U42452 (N_42452,N_39195,N_37740);
and U42453 (N_42453,N_37786,N_39139);
or U42454 (N_42454,N_38222,N_38508);
or U42455 (N_42455,N_38443,N_37797);
nand U42456 (N_42456,N_39225,N_39086);
nand U42457 (N_42457,N_37783,N_37704);
xnor U42458 (N_42458,N_39634,N_39593);
xnor U42459 (N_42459,N_39324,N_39931);
nor U42460 (N_42460,N_37587,N_38471);
nand U42461 (N_42461,N_39709,N_38633);
and U42462 (N_42462,N_38100,N_37588);
nor U42463 (N_42463,N_38993,N_38587);
nor U42464 (N_42464,N_38683,N_39299);
or U42465 (N_42465,N_37707,N_39607);
or U42466 (N_42466,N_38395,N_37576);
nand U42467 (N_42467,N_39963,N_38266);
xnor U42468 (N_42468,N_39035,N_38175);
nand U42469 (N_42469,N_38665,N_39864);
nand U42470 (N_42470,N_38096,N_39803);
nor U42471 (N_42471,N_39772,N_37774);
nor U42472 (N_42472,N_38928,N_39166);
nand U42473 (N_42473,N_37918,N_39066);
nor U42474 (N_42474,N_39795,N_38849);
nor U42475 (N_42475,N_39783,N_39573);
nand U42476 (N_42476,N_38324,N_38634);
nand U42477 (N_42477,N_39729,N_38237);
nand U42478 (N_42478,N_38815,N_38501);
xnor U42479 (N_42479,N_39888,N_39994);
nand U42480 (N_42480,N_39957,N_38320);
and U42481 (N_42481,N_38327,N_39768);
nand U42482 (N_42482,N_37506,N_38508);
nor U42483 (N_42483,N_38993,N_39672);
or U42484 (N_42484,N_38196,N_38310);
and U42485 (N_42485,N_38635,N_38003);
or U42486 (N_42486,N_38453,N_38709);
nor U42487 (N_42487,N_38944,N_38021);
xnor U42488 (N_42488,N_39236,N_38945);
nand U42489 (N_42489,N_39388,N_39209);
xor U42490 (N_42490,N_38698,N_38611);
and U42491 (N_42491,N_39548,N_39543);
nand U42492 (N_42492,N_39487,N_37650);
nand U42493 (N_42493,N_38655,N_38664);
and U42494 (N_42494,N_38013,N_38501);
nor U42495 (N_42495,N_39011,N_38844);
and U42496 (N_42496,N_39085,N_37800);
nor U42497 (N_42497,N_37511,N_37944);
and U42498 (N_42498,N_39155,N_39097);
nand U42499 (N_42499,N_39800,N_38322);
nor U42500 (N_42500,N_42445,N_42079);
and U42501 (N_42501,N_41829,N_41210);
nor U42502 (N_42502,N_41560,N_41494);
or U42503 (N_42503,N_40578,N_42340);
nor U42504 (N_42504,N_42447,N_41000);
or U42505 (N_42505,N_40406,N_41622);
and U42506 (N_42506,N_40385,N_40835);
and U42507 (N_42507,N_42227,N_41865);
and U42508 (N_42508,N_41596,N_42052);
nor U42509 (N_42509,N_40644,N_40845);
xnor U42510 (N_42510,N_41065,N_40588);
and U42511 (N_42511,N_40408,N_42276);
and U42512 (N_42512,N_42406,N_40494);
and U42513 (N_42513,N_40287,N_41266);
and U42514 (N_42514,N_40358,N_42377);
or U42515 (N_42515,N_40586,N_42464);
nor U42516 (N_42516,N_42026,N_41799);
xor U42517 (N_42517,N_40014,N_41761);
nand U42518 (N_42518,N_40271,N_40770);
or U42519 (N_42519,N_41279,N_41368);
or U42520 (N_42520,N_40846,N_41228);
nor U42521 (N_42521,N_42416,N_41040);
nor U42522 (N_42522,N_41236,N_40104);
and U42523 (N_42523,N_41696,N_41347);
or U42524 (N_42524,N_40660,N_42181);
nor U42525 (N_42525,N_42135,N_40451);
nand U42526 (N_42526,N_41904,N_40830);
or U42527 (N_42527,N_41199,N_41854);
nand U42528 (N_42528,N_41856,N_42129);
and U42529 (N_42529,N_42489,N_40280);
and U42530 (N_42530,N_41974,N_40817);
and U42531 (N_42531,N_42159,N_41863);
nand U42532 (N_42532,N_41657,N_42412);
or U42533 (N_42533,N_41933,N_42485);
nand U42534 (N_42534,N_40158,N_40472);
and U42535 (N_42535,N_41991,N_40464);
and U42536 (N_42536,N_40277,N_41949);
nand U42537 (N_42537,N_40521,N_42278);
and U42538 (N_42538,N_41072,N_40674);
nand U42539 (N_42539,N_41449,N_42338);
nor U42540 (N_42540,N_40795,N_40177);
and U42541 (N_42541,N_40087,N_41101);
or U42542 (N_42542,N_41250,N_40549);
nand U42543 (N_42543,N_42088,N_41203);
or U42544 (N_42544,N_41020,N_40975);
xor U42545 (N_42545,N_41446,N_42454);
nand U42546 (N_42546,N_42097,N_41176);
or U42547 (N_42547,N_40248,N_42323);
xor U42548 (N_42548,N_40194,N_40338);
nor U42549 (N_42549,N_41076,N_42016);
xor U42550 (N_42550,N_40082,N_40354);
and U42551 (N_42551,N_41839,N_41287);
or U42552 (N_42552,N_40321,N_41827);
nor U42553 (N_42553,N_41014,N_41524);
or U42554 (N_42554,N_41993,N_41906);
xnor U42555 (N_42555,N_42066,N_40992);
and U42556 (N_42556,N_40894,N_40422);
xnor U42557 (N_42557,N_41291,N_40323);
nor U42558 (N_42558,N_41424,N_41299);
or U42559 (N_42559,N_40049,N_40524);
nor U42560 (N_42560,N_42253,N_42220);
or U42561 (N_42561,N_42161,N_41378);
nand U42562 (N_42562,N_41788,N_40755);
or U42563 (N_42563,N_41840,N_41721);
and U42564 (N_42564,N_41514,N_40137);
or U42565 (N_42565,N_41711,N_42075);
nand U42566 (N_42566,N_42209,N_41779);
nand U42567 (N_42567,N_41237,N_41284);
xnor U42568 (N_42568,N_40314,N_41166);
or U42569 (N_42569,N_42178,N_40099);
and U42570 (N_42570,N_42341,N_40201);
and U42571 (N_42571,N_41530,N_40802);
or U42572 (N_42572,N_41013,N_40523);
xnor U42573 (N_42573,N_42186,N_42255);
nand U42574 (N_42574,N_41362,N_40225);
and U42575 (N_42575,N_41891,N_42262);
and U42576 (N_42576,N_40142,N_40043);
nand U42577 (N_42577,N_41197,N_41899);
or U42578 (N_42578,N_41874,N_40701);
nor U42579 (N_42579,N_41051,N_41685);
and U42580 (N_42580,N_40138,N_41771);
nand U42581 (N_42581,N_41802,N_40171);
nand U42582 (N_42582,N_40268,N_42003);
nor U42583 (N_42583,N_41443,N_40399);
and U42584 (N_42584,N_42370,N_40032);
nand U42585 (N_42585,N_41884,N_41179);
nor U42586 (N_42586,N_41998,N_42490);
and U42587 (N_42587,N_41147,N_42358);
nand U42588 (N_42588,N_41057,N_42395);
nand U42589 (N_42589,N_41476,N_41457);
nor U42590 (N_42590,N_41777,N_40242);
nand U42591 (N_42591,N_41447,N_42155);
nor U42592 (N_42592,N_42025,N_40543);
nor U42593 (N_42593,N_40526,N_41430);
and U42594 (N_42594,N_41823,N_42472);
nand U42595 (N_42595,N_40959,N_40347);
or U42596 (N_42596,N_41205,N_40196);
nor U42597 (N_42597,N_41209,N_41173);
nand U42598 (N_42598,N_41893,N_41086);
nor U42599 (N_42599,N_41716,N_42420);
nor U42600 (N_42600,N_40286,N_40373);
or U42601 (N_42601,N_40504,N_41545);
xor U42602 (N_42602,N_40465,N_41114);
nand U42603 (N_42603,N_41537,N_41644);
and U42604 (N_42604,N_41329,N_40782);
and U42605 (N_42605,N_42165,N_40890);
nor U42606 (N_42606,N_40355,N_42491);
or U42607 (N_42607,N_41715,N_40348);
nand U42608 (N_42608,N_41178,N_41202);
nand U42609 (N_42609,N_42113,N_42482);
nor U42610 (N_42610,N_41482,N_41499);
or U42611 (N_42611,N_42496,N_41158);
nor U42612 (N_42612,N_40761,N_40346);
nand U42613 (N_42613,N_42099,N_41623);
or U42614 (N_42614,N_40267,N_42004);
and U42615 (N_42615,N_41841,N_40360);
nor U42616 (N_42616,N_42098,N_42304);
xnor U42617 (N_42617,N_41169,N_41328);
nor U42618 (N_42618,N_41693,N_40365);
nand U42619 (N_42619,N_42011,N_40928);
xor U42620 (N_42620,N_40545,N_42419);
nor U42621 (N_42621,N_41023,N_40877);
and U42622 (N_42622,N_42002,N_41774);
xnor U42623 (N_42623,N_40769,N_41433);
and U42624 (N_42624,N_41087,N_40541);
nand U42625 (N_42625,N_40512,N_42204);
nor U42626 (N_42626,N_41379,N_40051);
and U42627 (N_42627,N_42384,N_41872);
and U42628 (N_42628,N_41531,N_40931);
or U42629 (N_42629,N_41533,N_41720);
xnor U42630 (N_42630,N_41021,N_40293);
or U42631 (N_42631,N_41647,N_41832);
or U42632 (N_42632,N_41566,N_41567);
nor U42633 (N_42633,N_40023,N_41763);
and U42634 (N_42634,N_41965,N_40832);
xnor U42635 (N_42635,N_40534,N_42465);
nor U42636 (N_42636,N_41668,N_42145);
or U42637 (N_42637,N_42141,N_42275);
or U42638 (N_42638,N_40468,N_41092);
nor U42639 (N_42639,N_40126,N_40950);
nand U42640 (N_42640,N_40172,N_42417);
xor U42641 (N_42641,N_41978,N_42133);
and U42642 (N_42642,N_40083,N_42134);
or U42643 (N_42643,N_41663,N_42254);
xnor U42644 (N_42644,N_40136,N_40463);
or U42645 (N_42645,N_41935,N_40539);
nand U42646 (N_42646,N_41405,N_40197);
or U42647 (N_42647,N_41645,N_41152);
or U42648 (N_42648,N_40527,N_42261);
nand U42649 (N_42649,N_41425,N_40309);
xor U42650 (N_42650,N_42425,N_40984);
nor U42651 (N_42651,N_40178,N_40934);
or U42652 (N_42652,N_40007,N_41879);
nor U42653 (N_42653,N_40694,N_40506);
xnor U42654 (N_42654,N_41230,N_40658);
nand U42655 (N_42655,N_40706,N_41359);
nor U42656 (N_42656,N_41201,N_41723);
nor U42657 (N_42657,N_42267,N_41925);
nor U42658 (N_42658,N_41670,N_41754);
or U42659 (N_42659,N_41324,N_42245);
nor U42660 (N_42660,N_41646,N_40981);
or U42661 (N_42661,N_42154,N_41049);
or U42662 (N_42662,N_40536,N_40439);
nor U42663 (N_42663,N_41188,N_40907);
nand U42664 (N_42664,N_42208,N_40767);
or U42665 (N_42665,N_40072,N_41349);
nor U42666 (N_42666,N_42424,N_40085);
xor U42667 (N_42667,N_41254,N_41793);
nand U42668 (N_42668,N_41369,N_41756);
nor U42669 (N_42669,N_40969,N_40994);
or U42670 (N_42670,N_40423,N_40038);
and U42671 (N_42671,N_42315,N_40628);
and U42672 (N_42672,N_40115,N_40234);
and U42673 (N_42673,N_41586,N_42012);
or U42674 (N_42674,N_40116,N_40988);
nand U42675 (N_42675,N_40392,N_41038);
nand U42676 (N_42676,N_40731,N_41027);
nor U42677 (N_42677,N_41615,N_41920);
nand U42678 (N_42678,N_40078,N_40317);
and U42679 (N_42679,N_41233,N_40977);
nor U42680 (N_42680,N_42202,N_41616);
xor U42681 (N_42681,N_41019,N_42009);
and U42682 (N_42682,N_40212,N_41985);
nor U42683 (N_42683,N_42122,N_42468);
or U42684 (N_42684,N_40017,N_42118);
nor U42685 (N_42685,N_41298,N_40686);
nor U42686 (N_42686,N_40966,N_40669);
nor U42687 (N_42687,N_42321,N_41951);
xnor U42688 (N_42688,N_40967,N_40488);
and U42689 (N_42689,N_42343,N_41394);
nor U42690 (N_42690,N_42336,N_41707);
and U42691 (N_42691,N_40645,N_40033);
and U42692 (N_42692,N_40489,N_40751);
nor U42693 (N_42693,N_41068,N_41714);
or U42694 (N_42694,N_41932,N_40517);
nor U42695 (N_42695,N_40129,N_40405);
or U42696 (N_42696,N_42397,N_41988);
nor U42697 (N_42697,N_41365,N_41597);
or U42698 (N_42698,N_40409,N_42451);
or U42699 (N_42699,N_40933,N_42110);
nand U42700 (N_42700,N_40379,N_40625);
nand U42701 (N_42701,N_42308,N_40807);
or U42702 (N_42702,N_42277,N_41046);
nand U42703 (N_42703,N_42345,N_41549);
xor U42704 (N_42704,N_41842,N_40161);
nand U42705 (N_42705,N_41052,N_41370);
and U42706 (N_42706,N_42284,N_40233);
and U42707 (N_42707,N_40119,N_41434);
and U42708 (N_42708,N_40842,N_40771);
nand U42709 (N_42709,N_42205,N_42211);
nand U42710 (N_42710,N_42102,N_40105);
nand U42711 (N_42711,N_40389,N_42070);
or U42712 (N_42712,N_41981,N_41061);
nor U42713 (N_42713,N_41285,N_40781);
nand U42714 (N_42714,N_42357,N_40786);
and U42715 (N_42715,N_41706,N_40282);
nand U42716 (N_42716,N_40125,N_41990);
nor U42717 (N_42717,N_40457,N_40708);
and U42718 (N_42718,N_41044,N_41964);
nand U42719 (N_42719,N_40476,N_42034);
xor U42720 (N_42720,N_41372,N_40016);
nor U42721 (N_42721,N_40712,N_41219);
nand U42722 (N_42722,N_41326,N_40165);
nand U42723 (N_42723,N_40011,N_40744);
nor U42724 (N_42724,N_42418,N_41914);
nand U42725 (N_42725,N_40829,N_42303);
nor U42726 (N_42726,N_41913,N_41760);
nor U42727 (N_42727,N_42230,N_41215);
nor U42728 (N_42728,N_42257,N_42317);
nand U42729 (N_42729,N_40444,N_40606);
and U42730 (N_42730,N_40419,N_41193);
nor U42731 (N_42731,N_40329,N_41187);
nor U42732 (N_42732,N_40961,N_40226);
xor U42733 (N_42733,N_40340,N_41684);
and U42734 (N_42734,N_40514,N_41834);
or U42735 (N_42735,N_41374,N_42353);
nand U42736 (N_42736,N_41507,N_41225);
nand U42737 (N_42737,N_41248,N_40434);
and U42738 (N_42738,N_42309,N_40861);
xor U42739 (N_42739,N_40273,N_40491);
nand U42740 (N_42740,N_41744,N_42214);
nor U42741 (N_42741,N_40905,N_41582);
and U42742 (N_42742,N_41541,N_41697);
nand U42743 (N_42743,N_42266,N_41127);
and U42744 (N_42744,N_41729,N_40693);
nand U42745 (N_42745,N_41358,N_42073);
nand U42746 (N_42746,N_41775,N_42189);
nand U42747 (N_42747,N_40054,N_40328);
or U42748 (N_42748,N_40163,N_41082);
nand U42749 (N_42749,N_41278,N_40307);
nand U42750 (N_42750,N_40505,N_41749);
xnor U42751 (N_42751,N_40453,N_40849);
xnor U42752 (N_42752,N_40735,N_40953);
or U42753 (N_42753,N_40486,N_40324);
and U42754 (N_42754,N_42398,N_41815);
nor U42755 (N_42755,N_40983,N_42263);
or U42756 (N_42756,N_40958,N_42362);
nor U42757 (N_42757,N_40583,N_40535);
nand U42758 (N_42758,N_40721,N_41513);
or U42759 (N_42759,N_41239,N_40474);
nand U42760 (N_42760,N_40727,N_41692);
nand U42761 (N_42761,N_42081,N_40508);
nor U42762 (N_42762,N_40519,N_41946);
xnor U42763 (N_42763,N_40264,N_40939);
nor U42764 (N_42764,N_40503,N_40677);
and U42765 (N_42765,N_42044,N_42428);
and U42766 (N_42766,N_40249,N_40942);
nand U42767 (N_42767,N_40777,N_41892);
and U42768 (N_42768,N_42068,N_40613);
nor U42769 (N_42769,N_40112,N_40106);
or U42770 (N_42770,N_40720,N_42125);
nor U42771 (N_42771,N_40438,N_40002);
nor U42772 (N_42772,N_42194,N_40568);
nand U42773 (N_42773,N_40263,N_40008);
or U42774 (N_42774,N_42248,N_41384);
nand U42775 (N_42775,N_40466,N_41496);
nor U42776 (N_42776,N_40925,N_41311);
and U42777 (N_42777,N_40481,N_42020);
nand U42778 (N_42778,N_41901,N_41255);
nand U42779 (N_42779,N_42167,N_41470);
nand U42780 (N_42780,N_40862,N_41383);
nand U42781 (N_42781,N_42055,N_40130);
nor U42782 (N_42782,N_40258,N_41491);
or U42783 (N_42783,N_40809,N_40773);
nor U42784 (N_42784,N_41734,N_42480);
xnor U42785 (N_42785,N_42492,N_40627);
nand U42786 (N_42786,N_41069,N_42136);
or U42787 (N_42787,N_40024,N_41438);
nand U42788 (N_42788,N_42438,N_41363);
nor U42789 (N_42789,N_42059,N_41585);
or U42790 (N_42790,N_40924,N_40614);
xor U42791 (N_42791,N_40956,N_40745);
nand U42792 (N_42792,N_40092,N_40883);
nand U42793 (N_42793,N_40401,N_41241);
nand U42794 (N_42794,N_40823,N_41776);
and U42795 (N_42795,N_41769,N_40326);
nor U42796 (N_42796,N_40923,N_42264);
nor U42797 (N_42797,N_41887,N_41948);
nand U42798 (N_42798,N_41943,N_40580);
or U42799 (N_42799,N_41216,N_42450);
and U42800 (N_42800,N_40272,N_41762);
xor U42801 (N_42801,N_41565,N_42233);
and U42802 (N_42802,N_41752,N_41942);
nor U42803 (N_42803,N_42282,N_41206);
nor U42804 (N_42804,N_42429,N_41157);
nor U42805 (N_42805,N_41428,N_40424);
and U42806 (N_42806,N_41624,N_40045);
nand U42807 (N_42807,N_40801,N_41168);
xnor U42808 (N_42808,N_40122,N_42144);
xor U42809 (N_42809,N_41252,N_40768);
and U42810 (N_42810,N_40251,N_42316);
nor U42811 (N_42811,N_41881,N_41375);
or U42812 (N_42812,N_40921,N_41674);
and U42813 (N_42813,N_40120,N_41970);
or U42814 (N_42814,N_40738,N_40612);
nor U42815 (N_42815,N_42064,N_41796);
nor U42816 (N_42816,N_42393,N_41142);
and U42817 (N_42817,N_41300,N_40775);
nor U42818 (N_42818,N_42077,N_40217);
nand U42819 (N_42819,N_41227,N_41705);
or U42820 (N_42820,N_40626,N_40684);
or U42821 (N_42821,N_40892,N_40396);
or U42822 (N_42822,N_41979,N_42057);
and U42823 (N_42823,N_41969,N_40575);
and U42824 (N_42824,N_40069,N_40029);
or U42825 (N_42825,N_41621,N_40719);
nor U42826 (N_42826,N_40134,N_41410);
or U42827 (N_42827,N_42061,N_40299);
and U42828 (N_42828,N_41850,N_41971);
nor U42829 (N_42829,N_41397,N_41083);
nor U42830 (N_42830,N_42008,N_41824);
or U42831 (N_42831,N_42219,N_42256);
or U42832 (N_42832,N_40790,N_40435);
xor U42833 (N_42833,N_42132,N_40776);
and U42834 (N_42834,N_42448,N_40603);
nor U42835 (N_42835,N_41912,N_41319);
nor U42836 (N_42836,N_41844,N_40009);
nand U42837 (N_42837,N_40943,N_42138);
nand U42838 (N_42838,N_41928,N_40733);
or U42839 (N_42839,N_42101,N_41804);
or U42840 (N_42840,N_42121,N_41195);
or U42841 (N_42841,N_40152,N_40577);
nand U42842 (N_42842,N_40058,N_40715);
nor U42843 (N_42843,N_41515,N_42179);
nor U42844 (N_42844,N_42225,N_42391);
xor U42845 (N_42845,N_40972,N_40840);
and U42846 (N_42846,N_41286,N_40891);
and U42847 (N_42847,N_42191,N_42244);
or U42848 (N_42848,N_40056,N_41024);
nand U42849 (N_42849,N_41973,N_40372);
xnor U42850 (N_42850,N_41118,N_42215);
and U42851 (N_42851,N_42497,N_40441);
and U42852 (N_42852,N_41544,N_40679);
and U42853 (N_42853,N_41699,N_41728);
and U42854 (N_42854,N_41529,N_40525);
nor U42855 (N_42855,N_40368,N_40245);
or U42856 (N_42856,N_41573,N_41427);
nand U42857 (N_42857,N_41355,N_40582);
or U42858 (N_42858,N_42127,N_40863);
and U42859 (N_42859,N_41261,N_41026);
or U42860 (N_42860,N_40095,N_40594);
and U42861 (N_42861,N_42022,N_40900);
nor U42862 (N_42862,N_42476,N_41063);
and U42863 (N_42863,N_42210,N_40602);
or U42864 (N_42864,N_42242,N_40634);
nand U42865 (N_42865,N_41940,N_41032);
nor U42866 (N_42866,N_41121,N_40109);
and U42867 (N_42867,N_42290,N_42457);
and U42868 (N_42868,N_40337,N_40980);
nand U42869 (N_42869,N_41764,N_41648);
xor U42870 (N_42870,N_40901,N_40666);
nor U42871 (N_42871,N_41703,N_40370);
nor U42872 (N_42872,N_40495,N_40652);
or U42873 (N_42873,N_41277,N_40743);
nor U42874 (N_42874,N_42095,N_42301);
or U42875 (N_42875,N_42363,N_40064);
nor U42876 (N_42876,N_42123,N_41005);
nor U42877 (N_42877,N_42330,N_40182);
nand U42878 (N_42878,N_41441,N_42168);
and U42879 (N_42879,N_41126,N_40882);
nor U42880 (N_42880,N_40833,N_42047);
nor U42881 (N_42881,N_42222,N_41709);
and U42882 (N_42882,N_40390,N_40675);
and U42883 (N_42883,N_41478,N_40139);
nand U42884 (N_42884,N_41836,N_42197);
and U42885 (N_42885,N_41497,N_40274);
nor U42886 (N_42886,N_40303,N_42265);
xnor U42887 (N_42887,N_41498,N_40034);
xor U42888 (N_42888,N_40015,N_41325);
or U42889 (N_42889,N_41941,N_40203);
and U42890 (N_42890,N_40607,N_42328);
nand U42891 (N_42891,N_42162,N_42147);
and U42892 (N_42892,N_41308,N_40855);
and U42893 (N_42893,N_41315,N_41518);
or U42894 (N_42894,N_41784,N_42414);
nor U42895 (N_42895,N_41629,N_40055);
nor U42896 (N_42896,N_40920,N_42359);
or U42897 (N_42897,N_40250,N_41245);
nor U42898 (N_42898,N_41382,N_42131);
and U42899 (N_42899,N_40432,N_40713);
or U42900 (N_42900,N_42484,N_42176);
nor U42901 (N_42901,N_42350,N_42394);
or U42902 (N_42902,N_42324,N_40458);
and U42903 (N_42903,N_40787,N_41634);
and U42904 (N_42904,N_42382,N_41407);
or U42905 (N_42905,N_42369,N_41505);
or U42906 (N_42906,N_42349,N_41698);
nand U42907 (N_42907,N_42148,N_40709);
and U42908 (N_42908,N_40803,N_42051);
xor U42909 (N_42909,N_41619,N_40332);
nand U42910 (N_42910,N_41035,N_42031);
and U42911 (N_42911,N_41556,N_40252);
nand U42912 (N_42912,N_40088,N_40825);
nor U42913 (N_42913,N_40334,N_41704);
and U42914 (N_42914,N_40210,N_42335);
nand U42915 (N_42915,N_42030,N_41414);
nand U42916 (N_42916,N_40144,N_41066);
and U42917 (N_42917,N_42106,N_41156);
and U42918 (N_42918,N_40948,N_40620);
and U42919 (N_42919,N_41161,N_40430);
nor U42920 (N_42920,N_41937,N_40828);
xnor U42921 (N_42921,N_41992,N_42319);
nor U42922 (N_42922,N_40382,N_40176);
or U42923 (N_42923,N_40393,N_40499);
and U42924 (N_42924,N_41058,N_42435);
xnor U42925 (N_42925,N_40595,N_42313);
and U42926 (N_42926,N_40622,N_41956);
nor U42927 (N_42927,N_41265,N_41712);
and U42928 (N_42928,N_40698,N_42177);
or U42929 (N_42929,N_40611,N_42413);
or U42930 (N_42930,N_40343,N_40871);
and U42931 (N_42931,N_40223,N_40131);
nor U42932 (N_42932,N_40878,N_40854);
or U42933 (N_42933,N_41594,N_40554);
nor U42934 (N_42934,N_40230,N_41309);
or U42935 (N_42935,N_40780,N_42366);
nand U42936 (N_42936,N_41117,N_41316);
and U42937 (N_42937,N_41364,N_42116);
nand U42938 (N_42938,N_40636,N_42421);
nand U42939 (N_42939,N_42272,N_40367);
nand U42940 (N_42940,N_41732,N_41532);
or U42941 (N_42941,N_40352,N_40522);
nor U42942 (N_42942,N_41520,N_41096);
nand U42943 (N_42943,N_40687,N_41811);
or U42944 (N_42944,N_42183,N_40195);
nand U42945 (N_42945,N_41090,N_41570);
nand U42946 (N_42946,N_40315,N_41898);
nand U42947 (N_42947,N_40736,N_40973);
nor U42948 (N_42948,N_41562,N_42326);
and U42949 (N_42949,N_41831,N_42374);
nand U42950 (N_42950,N_40168,N_40574);
and U42951 (N_42951,N_40560,N_40889);
nor U42952 (N_42952,N_41695,N_42433);
nand U42953 (N_42953,N_41212,N_40822);
and U42954 (N_42954,N_42314,N_40593);
nor U42955 (N_42955,N_41805,N_42458);
or U42956 (N_42956,N_40812,N_41675);
xnor U42957 (N_42957,N_41757,N_41034);
or U42958 (N_42958,N_42249,N_41574);
nor U42959 (N_42959,N_40060,N_42015);
nand U42960 (N_42960,N_40429,N_40440);
nand U42961 (N_42961,N_40487,N_41578);
or U42962 (N_42962,N_42401,N_41897);
xor U42963 (N_42963,N_42234,N_41190);
and U42964 (N_42964,N_40363,N_40552);
xnor U42965 (N_42965,N_41613,N_40659);
or U42966 (N_42966,N_40874,N_41938);
nor U42967 (N_42967,N_41452,N_40123);
nor U42968 (N_42968,N_40717,N_42471);
or U42969 (N_42969,N_42050,N_40623);
and U42970 (N_42970,N_40316,N_40689);
and U42971 (N_42971,N_41817,N_41165);
nor U42972 (N_42972,N_41304,N_40870);
nor U42973 (N_42973,N_41608,N_41852);
nand U42974 (N_42974,N_42446,N_41204);
or U42975 (N_42975,N_41994,N_41639);
xor U42976 (N_42976,N_41396,N_40670);
or U42977 (N_42977,N_42221,N_41876);
and U42978 (N_42978,N_42273,N_41469);
or U42979 (N_42979,N_41381,N_40547);
or U42980 (N_42980,N_41310,N_40885);
or U42981 (N_42981,N_41730,N_41012);
xnor U42982 (N_42982,N_40858,N_41662);
and U42983 (N_42983,N_41883,N_41577);
xor U42984 (N_42984,N_41855,N_42188);
or U42985 (N_42985,N_41004,N_41767);
and U42986 (N_42986,N_40188,N_40414);
xor U42987 (N_42987,N_40053,N_40470);
nor U42988 (N_42988,N_40810,N_40538);
nand U42989 (N_42989,N_40199,N_40661);
nor U42990 (N_42990,N_42185,N_40255);
and U42991 (N_42991,N_40325,N_40847);
nand U42992 (N_42992,N_40425,N_40908);
and U42993 (N_42993,N_41352,N_40797);
and U42994 (N_42994,N_41493,N_40609);
nor U42995 (N_42995,N_41790,N_41847);
nand U42996 (N_42996,N_40851,N_40591);
nand U42997 (N_42997,N_42250,N_42160);
or U42998 (N_42998,N_42207,N_40254);
xor U42999 (N_42999,N_40551,N_42402);
nor U43000 (N_43000,N_40872,N_40193);
and U43001 (N_43001,N_42281,N_42058);
and U43002 (N_43002,N_40540,N_40690);
nand U43003 (N_43003,N_41667,N_40754);
or U43004 (N_43004,N_40906,N_40000);
nor U43005 (N_43005,N_41272,N_42346);
nand U43006 (N_43006,N_40167,N_40986);
xor U43007 (N_43007,N_40362,N_41880);
or U43008 (N_43008,N_41327,N_42403);
or U43009 (N_43009,N_41408,N_41742);
or U43010 (N_43010,N_41361,N_41207);
and U43011 (N_43011,N_40778,N_40615);
nor U43012 (N_43012,N_41314,N_40269);
and U43013 (N_43013,N_41268,N_41385);
and U43014 (N_43014,N_41045,N_40564);
and U43015 (N_43015,N_40221,N_42461);
nor U43016 (N_43016,N_40766,N_40960);
and U43017 (N_43017,N_41139,N_41540);
nor U43018 (N_43018,N_40410,N_40673);
xor U43019 (N_43019,N_42029,N_41910);
and U43020 (N_43020,N_41404,N_40207);
nor U43021 (N_43021,N_41133,N_41183);
nor U43022 (N_43022,N_40198,N_41812);
and U43023 (N_43023,N_41075,N_40443);
and U43024 (N_43024,N_41743,N_41896);
or U43025 (N_43025,N_41751,N_40804);
nor U43026 (N_43026,N_41356,N_41116);
and U43027 (N_43027,N_40876,N_42427);
and U43028 (N_43028,N_40153,N_40556);
nor U43029 (N_43029,N_41043,N_40816);
nor U43030 (N_43030,N_41388,N_42237);
nor U43031 (N_43031,N_42103,N_41801);
nor U43032 (N_43032,N_42013,N_41312);
xnor U43033 (N_43033,N_40955,N_41944);
or U43034 (N_43034,N_42074,N_40159);
nand U43035 (N_43035,N_40298,N_40990);
and U43036 (N_43036,N_41977,N_40218);
and U43037 (N_43037,N_40962,N_40037);
nand U43038 (N_43038,N_41463,N_40837);
nor U43039 (N_43039,N_40655,N_41908);
and U43040 (N_43040,N_40202,N_42296);
or U43041 (N_43041,N_41996,N_41015);
xnor U43042 (N_43042,N_40700,N_41975);
and U43043 (N_43043,N_41922,N_42432);
nor U43044 (N_43044,N_40676,N_42046);
xor U43045 (N_43045,N_40156,N_40827);
nand U43046 (N_43046,N_40544,N_40327);
xnor U43047 (N_43047,N_42119,N_41780);
and U43048 (N_43048,N_42229,N_40289);
or U43049 (N_43049,N_41295,N_41818);
and U43050 (N_43050,N_41568,N_41313);
xor U43051 (N_43051,N_41917,N_40707);
nand U43052 (N_43052,N_41398,N_41345);
nand U43053 (N_43053,N_41002,N_41386);
xor U43054 (N_43054,N_41642,N_40589);
or U43055 (N_43055,N_42224,N_41030);
nor U43056 (N_43056,N_40750,N_41955);
nor U43057 (N_43057,N_40985,N_42067);
and U43058 (N_43058,N_41579,N_40035);
nand U43059 (N_43059,N_40759,N_40621);
nor U43060 (N_43060,N_40187,N_42478);
nor U43061 (N_43061,N_42373,N_40036);
and U43062 (N_43062,N_42364,N_40175);
nor U43063 (N_43063,N_42298,N_40987);
nor U43064 (N_43064,N_42217,N_41828);
xor U43065 (N_43065,N_42322,N_41475);
nand U43066 (N_43066,N_40799,N_41864);
or U43067 (N_43067,N_41708,N_40302);
and U43068 (N_43068,N_41546,N_40572);
nor U43069 (N_43069,N_41590,N_40157);
nand U43070 (N_43070,N_42174,N_40581);
or U43071 (N_43071,N_40141,N_41726);
nand U43072 (N_43072,N_41822,N_41950);
and U43073 (N_43073,N_42201,N_41671);
nand U43074 (N_43074,N_42386,N_41125);
or U43075 (N_43075,N_41104,N_41486);
or U43076 (N_43076,N_40704,N_41957);
nor U43077 (N_43077,N_40420,N_41995);
nand U43078 (N_43078,N_41007,N_40963);
or U43079 (N_43079,N_42071,N_41042);
nand U43080 (N_43080,N_40957,N_40063);
or U43081 (N_43081,N_41354,N_40909);
xor U43082 (N_43082,N_41094,N_41553);
nand U43083 (N_43083,N_40378,N_42005);
or U43084 (N_43084,N_40919,N_40147);
nor U43085 (N_43085,N_41851,N_40412);
nor U43086 (N_43086,N_40844,N_41724);
nor U43087 (N_43087,N_42283,N_40562);
and U43088 (N_43088,N_40654,N_40914);
and U43089 (N_43089,N_41987,N_41343);
nand U43090 (N_43090,N_41921,N_41246);
nand U43091 (N_43091,N_40235,N_42368);
xnor U43092 (N_43092,N_40520,N_42286);
and U43093 (N_43093,N_40947,N_40741);
nor U43094 (N_43094,N_42087,N_42260);
nor U43095 (N_43095,N_41633,N_41819);
nor U43096 (N_43096,N_40301,N_41939);
xor U43097 (N_43097,N_41303,N_41809);
and U43098 (N_43098,N_40737,N_42027);
or U43099 (N_43099,N_41924,N_41797);
and U43100 (N_43100,N_40111,N_40646);
or U43101 (N_43101,N_42259,N_40428);
nand U43102 (N_43102,N_40135,N_40374);
nand U43103 (N_43103,N_42411,N_40240);
xor U43104 (N_43104,N_40490,N_41778);
and U43105 (N_43105,N_40734,N_41650);
nor U43106 (N_43106,N_41517,N_40189);
and U43107 (N_43107,N_41905,N_42238);
nand U43108 (N_43108,N_40529,N_41807);
nand U43109 (N_43109,N_41509,N_41357);
and U43110 (N_43110,N_41640,N_41664);
or U43111 (N_43111,N_41773,N_40573);
nand U43112 (N_43112,N_41412,N_41638);
nor U43113 (N_43113,N_41522,N_42049);
nand U43114 (N_43114,N_40330,N_42376);
and U43115 (N_43115,N_42137,N_42231);
and U43116 (N_43116,N_42470,N_41172);
or U43117 (N_43117,N_41963,N_41947);
and U43118 (N_43118,N_41552,N_41008);
nand U43119 (N_43119,N_40351,N_40387);
and U43120 (N_43120,N_40935,N_42038);
and U43121 (N_43121,N_41067,N_42334);
and U43122 (N_43122,N_41089,N_41909);
xor U43123 (N_43123,N_41402,N_42203);
nor U43124 (N_43124,N_42035,N_41589);
and U43125 (N_43125,N_40515,N_40576);
nor U43126 (N_43126,N_40569,N_40027);
and U43127 (N_43127,N_41198,N_41124);
nor U43128 (N_43128,N_41601,N_40788);
nand U43129 (N_43129,N_40976,N_42043);
and U43130 (N_43130,N_41733,N_41606);
or U43131 (N_43131,N_40046,N_42356);
nor U43132 (N_43132,N_40445,N_42436);
nand U43133 (N_43133,N_40090,N_40021);
and U43134 (N_43134,N_42467,N_40169);
and U43135 (N_43135,N_41466,N_40902);
nor U43136 (N_43136,N_41748,N_42040);
and U43137 (N_43137,N_40079,N_40630);
and U43138 (N_43138,N_40084,N_41062);
or U43139 (N_43139,N_41387,N_41149);
nand U43140 (N_43140,N_40006,N_41317);
or U43141 (N_43141,N_42193,N_40341);
and U43142 (N_43142,N_41442,N_41722);
xnor U43143 (N_43143,N_41334,N_41580);
and U43144 (N_43144,N_41335,N_41502);
and U43145 (N_43145,N_42453,N_41867);
or U43146 (N_43146,N_40208,N_40559);
or U43147 (N_43147,N_42383,N_40665);
and U43148 (N_43148,N_40477,N_40467);
nand U43149 (N_43149,N_41487,N_40710);
and U43150 (N_43150,N_41244,N_41625);
and U43151 (N_43151,N_41945,N_41341);
or U43152 (N_43152,N_40610,N_41416);
nor U43153 (N_43153,N_41554,N_41808);
xnor U43154 (N_43154,N_41563,N_40600);
nor U43155 (N_43155,N_40791,N_41194);
or U43156 (N_43156,N_41274,N_41267);
nand U43157 (N_43157,N_41229,N_40678);
nor U43158 (N_43158,N_41655,N_40604);
xnor U43159 (N_43159,N_41485,N_40200);
and U43160 (N_43160,N_41962,N_40369);
nand U43161 (N_43161,N_42385,N_42289);
nor U43162 (N_43162,N_41677,N_40867);
xor U43163 (N_43163,N_41232,N_41700);
and U43164 (N_43164,N_41857,N_40456);
and U43165 (N_43165,N_41353,N_41710);
nor U43166 (N_43166,N_40730,N_42327);
xor U43167 (N_43167,N_40760,N_41281);
and U43168 (N_43168,N_41064,N_42437);
nor U43169 (N_43169,N_42018,N_41115);
nor U43170 (N_43170,N_40532,N_41571);
nand U43171 (N_43171,N_40567,N_40320);
nor U43172 (N_43172,N_40711,N_41555);
or U43173 (N_43173,N_40074,N_41782);
nand U43174 (N_43174,N_40682,N_41542);
or U43175 (N_43175,N_40296,N_40164);
nor U43176 (N_43176,N_42499,N_41451);
and U43177 (N_43177,N_40398,N_41665);
nor U43178 (N_43178,N_41792,N_40893);
or U43179 (N_43179,N_40146,N_42192);
xor U43180 (N_43180,N_40229,N_42232);
nor U43181 (N_43181,N_40070,N_40256);
and U43182 (N_43182,N_41367,N_40071);
or U43183 (N_43183,N_42228,N_41095);
nor U43184 (N_43184,N_42032,N_40404);
and U43185 (N_43185,N_41474,N_40565);
nor U43186 (N_43186,N_41109,N_41666);
nor U43187 (N_43187,N_41223,N_42111);
and U43188 (N_43188,N_41609,N_40765);
nor U43189 (N_43189,N_41569,N_42422);
xnor U43190 (N_43190,N_42173,N_40062);
nor U43191 (N_43191,N_42409,N_41600);
or U43192 (N_43192,N_40231,N_40391);
and U43193 (N_43193,N_40763,N_40886);
or U43194 (N_43194,N_40501,N_41504);
nor U43195 (N_43195,N_42297,N_42062);
or U43196 (N_43196,N_40026,N_41342);
and U43197 (N_43197,N_40304,N_40815);
nor U43198 (N_43198,N_41907,N_42163);
nor U43199 (N_43199,N_40259,N_40010);
or U43200 (N_43200,N_40705,N_42084);
or U43201 (N_43201,N_40306,N_41462);
and U43202 (N_43202,N_40103,N_42037);
nand U43203 (N_43203,N_40672,N_40018);
and U43204 (N_43204,N_42021,N_40050);
nand U43205 (N_43205,N_42182,N_40852);
nor U43206 (N_43206,N_40794,N_42469);
nand U43207 (N_43207,N_40281,N_40726);
or U43208 (N_43208,N_40896,N_41936);
nand U43209 (N_43209,N_41968,N_40903);
nand U43210 (N_43210,N_41289,N_42400);
and U43211 (N_43211,N_41192,N_41798);
nor U43212 (N_43212,N_40598,N_41806);
and U43213 (N_43213,N_40469,N_40991);
or U43214 (N_43214,N_40566,N_40128);
nor U43215 (N_43215,N_41659,N_41717);
nand U43216 (N_43216,N_42488,N_40528);
xnor U43217 (N_43217,N_41826,N_40459);
nor U43218 (N_43218,N_41725,N_41330);
and U43219 (N_43219,N_41660,N_40318);
nand U43220 (N_43220,N_40542,N_40048);
and U43221 (N_43221,N_41468,N_41348);
or U43222 (N_43222,N_40772,N_40758);
nand U43223 (N_43223,N_40965,N_41795);
and U43224 (N_43224,N_41534,N_42268);
and U43225 (N_43225,N_40149,N_40742);
nand U43226 (N_43226,N_40400,N_41830);
xor U43227 (N_43227,N_41952,N_40848);
nand U43228 (N_43228,N_41911,N_42223);
and U43229 (N_43229,N_41618,N_40025);
nor U43230 (N_43230,N_40998,N_41003);
nand U43231 (N_43231,N_42390,N_40571);
and U43232 (N_43232,N_41878,N_40946);
or U43233 (N_43233,N_40190,N_40285);
nor U43234 (N_43234,N_41459,N_42293);
nor U43235 (N_43235,N_42089,N_41984);
or U43236 (N_43236,N_40498,N_41512);
nand U43237 (N_43237,N_40563,N_41221);
or U43238 (N_43238,N_41678,N_41983);
nor U43239 (N_43239,N_40215,N_40096);
nand U43240 (N_43240,N_40284,N_40898);
and U43241 (N_43241,N_41536,N_40031);
xor U43242 (N_43242,N_42156,N_42387);
nor U43243 (N_43243,N_41243,N_41448);
or U43244 (N_43244,N_40133,N_41132);
nand U43245 (N_43245,N_41886,N_41171);
nor U43246 (N_43246,N_41174,N_40022);
or U43247 (N_43247,N_40283,N_42475);
and U43248 (N_43248,N_40557,N_40294);
nand U43249 (N_43249,N_42006,N_40632);
or U43250 (N_43250,N_40618,N_40642);
or U43251 (N_43251,N_40236,N_40699);
nand U43252 (N_43252,N_42086,N_40297);
nand U43253 (N_43253,N_40004,N_42239);
and U43254 (N_43254,N_41745,N_41269);
nand U43255 (N_43255,N_41612,N_41611);
xnor U43256 (N_43256,N_40356,N_41649);
xnor U43257 (N_43257,N_41406,N_41559);
nor U43258 (N_43258,N_41495,N_42007);
nand U43259 (N_43259,N_41628,N_41120);
or U43260 (N_43260,N_42460,N_41113);
xnor U43261 (N_43261,N_41108,N_40342);
and U43262 (N_43262,N_41750,N_40841);
or U43263 (N_43263,N_41592,N_40811);
nand U43264 (N_43264,N_41894,N_40764);
xnor U43265 (N_43265,N_41143,N_42389);
nand U43266 (N_43266,N_41041,N_41869);
xnor U43267 (N_43267,N_41595,N_41017);
or U43268 (N_43268,N_41997,N_41321);
nor U43269 (N_43269,N_41632,N_40395);
or U43270 (N_43270,N_40478,N_40216);
or U43271 (N_43271,N_42115,N_41288);
and U43272 (N_43272,N_41249,N_40001);
nand U43273 (N_43273,N_42198,N_41653);
and U43274 (N_43274,N_42439,N_40793);
nand U43275 (N_43275,N_40148,N_40880);
nor U43276 (N_43276,N_42473,N_40915);
or U43277 (N_43277,N_40619,N_42126);
nor U43278 (N_43278,N_41794,N_40929);
nor U43279 (N_43279,N_40968,N_41687);
nand U43280 (N_43280,N_42195,N_40380);
nor U43281 (N_43281,N_40426,N_41401);
nand U43282 (N_43282,N_41719,N_40143);
or U43283 (N_43283,N_40729,N_41526);
nor U43284 (N_43284,N_40624,N_40656);
nand U43285 (N_43285,N_42130,N_41181);
nand U43286 (N_43286,N_40114,N_40421);
nor U43287 (N_43287,N_40671,N_42483);
nand U43288 (N_43288,N_42307,N_40941);
nor U43289 (N_43289,N_42442,N_41037);
and U43290 (N_43290,N_40290,N_41050);
nor U43291 (N_43291,N_41755,N_42251);
nor U43292 (N_43292,N_41162,N_41418);
nor U43293 (N_43293,N_40091,N_42477);
nor U43294 (N_43294,N_42033,N_40437);
nand U43295 (N_43295,N_41680,N_41602);
or U43296 (N_43296,N_41079,N_40546);
nand U43297 (N_43297,N_42299,N_42117);
nand U43298 (N_43298,N_40910,N_41803);
nand U43299 (N_43299,N_42092,N_41006);
nor U43300 (N_43300,N_40496,N_41413);
xor U43301 (N_43301,N_42172,N_42128);
nor U43302 (N_43302,N_41868,N_42112);
xor U43303 (N_43303,N_41581,N_40899);
nor U43304 (N_43304,N_40266,N_40930);
nand U43305 (N_43305,N_42380,N_40789);
nand U43306 (N_43306,N_41191,N_41718);
and U43307 (N_43307,N_41163,N_40927);
or U43308 (N_43308,N_40839,N_42190);
or U43309 (N_43309,N_41256,N_40361);
and U43310 (N_43310,N_42440,N_41417);
xor U43311 (N_43311,N_40483,N_40971);
nor U43312 (N_43312,N_42017,N_40997);
nor U43313 (N_43313,N_41954,N_41453);
xnor U43314 (N_43314,N_40663,N_41861);
or U43315 (N_43315,N_42305,N_41376);
nand U43316 (N_43316,N_42039,N_40418);
or U43317 (N_43317,N_40170,N_42295);
or U43318 (N_43318,N_42171,N_42184);
and U43319 (N_43319,N_41322,N_42449);
or U43320 (N_43320,N_41189,N_41242);
xnor U43321 (N_43321,N_41614,N_41890);
or U43322 (N_43322,N_42352,N_41455);
and U43323 (N_43323,N_40785,N_41234);
nand U43324 (N_43324,N_40110,N_40553);
nand U43325 (N_43325,N_40650,N_40639);
and U43326 (N_43326,N_42360,N_41099);
or U43327 (N_43327,N_40319,N_40657);
and U43328 (N_43328,N_41845,N_41766);
xor U43329 (N_43329,N_40692,N_40278);
nand U43330 (N_43330,N_41652,N_41521);
nand U43331 (N_43331,N_41247,N_40066);
and U43332 (N_43332,N_42410,N_40836);
or U43333 (N_43333,N_41182,N_40716);
and U43334 (N_43334,N_40450,N_41631);
xor U43335 (N_43335,N_41643,N_41858);
nand U43336 (N_43336,N_41294,N_40081);
nor U43337 (N_43337,N_41877,N_41055);
and U43338 (N_43338,N_42294,N_41122);
nand U43339 (N_43339,N_40857,N_41539);
nand U43340 (N_43340,N_40860,N_41366);
or U43341 (N_43341,N_41843,N_41888);
xor U43342 (N_43342,N_40019,N_40587);
nor U43343 (N_43343,N_42213,N_41875);
or U43344 (N_43344,N_40295,N_40922);
and U43345 (N_43345,N_40166,N_40897);
nor U43346 (N_43346,N_40637,N_40668);
or U43347 (N_43347,N_40206,N_40649);
nand U43348 (N_43348,N_41186,N_41053);
or U43349 (N_43349,N_40417,N_41253);
xnor U43350 (N_43350,N_41436,N_42365);
or U43351 (N_43351,N_41461,N_41175);
xor U43352 (N_43352,N_40416,N_42287);
and U43353 (N_43353,N_41070,N_40375);
or U43354 (N_43354,N_41025,N_41848);
nand U43355 (N_43355,N_42169,N_41047);
nor U43356 (N_43356,N_42120,N_42375);
and U43357 (N_43357,N_41271,N_41338);
nor U43358 (N_43358,N_41727,N_40974);
or U43359 (N_43359,N_41439,N_40211);
xnor U43360 (N_43360,N_42279,N_42083);
and U43361 (N_43361,N_41078,N_42023);
nand U43362 (N_43362,N_40869,N_42036);
and U43363 (N_43363,N_41576,N_40232);
and U43364 (N_43364,N_42495,N_40511);
or U43365 (N_43365,N_41654,N_40308);
xnor U43366 (N_43366,N_41154,N_41214);
nand U43367 (N_43367,N_42459,N_41488);
and U43368 (N_43368,N_42028,N_40596);
nor U43369 (N_43369,N_41200,N_40411);
and U43370 (N_43370,N_40821,N_41479);
nor U43371 (N_43371,N_40140,N_41337);
nand U43372 (N_43372,N_41658,N_41184);
nand U43373 (N_43373,N_41102,N_41603);
nor U43374 (N_43374,N_41519,N_40643);
or U43375 (N_43375,N_41926,N_40005);
or U43376 (N_43376,N_41141,N_41036);
or U43377 (N_43377,N_42434,N_40774);
nor U43378 (N_43378,N_40185,N_40555);
nand U43379 (N_43379,N_40276,N_41123);
nand U43380 (N_43380,N_40473,N_41435);
and U43381 (N_43381,N_40843,N_42354);
nor U43382 (N_43382,N_40376,N_40270);
nand U43383 (N_43383,N_40680,N_42408);
nand U43384 (N_43384,N_42493,N_41960);
nand U43385 (N_43385,N_41862,N_42166);
nor U43386 (N_43386,N_41501,N_40601);
or U43387 (N_43387,N_40349,N_40866);
xor U43388 (N_43388,N_40331,N_40982);
xor U43389 (N_43389,N_41160,N_41196);
or U43390 (N_43390,N_41208,N_41835);
or U43391 (N_43391,N_41426,N_40228);
nand U43392 (N_43392,N_41465,N_41849);
nand U43393 (N_43393,N_41218,N_42443);
xor U43394 (N_43394,N_41420,N_40204);
nand U43395 (N_43395,N_40089,N_41604);
nand U43396 (N_43396,N_42379,N_41022);
and U43397 (N_43397,N_41953,N_42342);
nand U43398 (N_43398,N_41084,N_41630);
and U43399 (N_43399,N_42216,N_41587);
or U43400 (N_43400,N_41339,N_40641);
xnor U43401 (N_43401,N_40800,N_41982);
nand U43402 (N_43402,N_40237,N_41636);
xnor U43403 (N_43403,N_40502,N_41813);
and U43404 (N_43404,N_40856,N_40599);
or U43405 (N_43405,N_40359,N_41018);
nand U43406 (N_43406,N_40608,N_40640);
and U43407 (N_43407,N_41467,N_40243);
nor U43408 (N_43408,N_40335,N_42226);
and U43409 (N_43409,N_40779,N_42200);
and U43410 (N_43410,N_41033,N_40461);
xnor U43411 (N_43411,N_41525,N_40753);
nor U43412 (N_43412,N_41283,N_40746);
and U43413 (N_43413,N_40403,N_42001);
nand U43414 (N_43414,N_41617,N_40756);
and U43415 (N_43415,N_41185,N_40383);
nand U43416 (N_43416,N_42396,N_42108);
nand U43417 (N_43417,N_41810,N_41136);
nand U43418 (N_43418,N_40484,N_40260);
nand U43419 (N_43419,N_41572,N_40718);
and U43420 (N_43420,N_41758,N_40413);
and U43421 (N_43421,N_40558,N_41275);
nor U43422 (N_43422,N_40073,N_42065);
nor U43423 (N_43423,N_40814,N_40918);
or U43424 (N_43424,N_40460,N_40184);
or U43425 (N_43425,N_40507,N_40020);
and U43426 (N_43426,N_41444,N_40311);
and U43427 (N_43427,N_42302,N_41772);
nor U43428 (N_43428,N_40531,N_41551);
nor U43429 (N_43429,N_42241,N_40605);
or U43430 (N_43430,N_40695,N_42332);
nor U43431 (N_43431,N_41785,N_41377);
nor U43432 (N_43432,N_40057,N_41871);
nor U43433 (N_43433,N_41598,N_41930);
and U43434 (N_43434,N_41490,N_40585);
nor U43435 (N_43435,N_40792,N_41679);
and U43436 (N_43436,N_41736,N_41506);
nor U43437 (N_43437,N_40485,N_42105);
or U43438 (N_43438,N_42311,N_40044);
nor U43439 (N_43439,N_40471,N_40747);
and U43440 (N_43440,N_41610,N_42310);
nor U43441 (N_43441,N_41130,N_40638);
or U43442 (N_43442,N_41231,N_40702);
nor U43443 (N_43443,N_41681,N_41672);
nand U43444 (N_43444,N_40510,N_40344);
and U43445 (N_43445,N_42423,N_42325);
or U43446 (N_43446,N_40214,N_42481);
and U43447 (N_43447,N_41251,N_42157);
nor U43448 (N_43448,N_42218,N_41967);
or U43449 (N_43449,N_40312,N_40030);
and U43450 (N_43450,N_41016,N_42060);
and U43451 (N_43451,N_40068,N_42246);
and U43452 (N_43452,N_41740,N_40310);
nand U43453 (N_43453,N_40292,N_42142);
or U43454 (N_43454,N_40384,N_40313);
xnor U43455 (N_43455,N_40042,N_40397);
and U43456 (N_43456,N_40150,N_41220);
and U43457 (N_43457,N_41787,N_41048);
nand U43458 (N_43458,N_41054,N_40509);
nand U43459 (N_43459,N_40722,N_40749);
nand U43460 (N_43460,N_41923,N_41471);
nand U43461 (N_43461,N_41263,N_42331);
xnor U43462 (N_43462,N_40859,N_40039);
and U43463 (N_43463,N_42288,N_40040);
and U43464 (N_43464,N_40932,N_42076);
xnor U43465 (N_43465,N_40725,N_41391);
or U43466 (N_43466,N_42367,N_41492);
and U43467 (N_43467,N_42270,N_42372);
xor U43468 (N_43468,N_40970,N_42090);
xor U43469 (N_43469,N_40868,N_40584);
nand U43470 (N_43470,N_41895,N_40631);
and U43471 (N_43471,N_41081,N_42212);
or U43472 (N_43472,N_41959,N_41292);
or U43473 (N_43473,N_40683,N_40446);
or U43474 (N_43474,N_41001,N_40550);
nor U43475 (N_43475,N_41085,N_40996);
or U43476 (N_43476,N_41150,N_42348);
nor U43477 (N_43477,N_40592,N_42312);
or U43478 (N_43478,N_41903,N_41535);
xor U43479 (N_43479,N_41464,N_42063);
xor U43480 (N_43480,N_41870,N_42361);
or U43481 (N_43481,N_41833,N_41682);
nand U43482 (N_43482,N_41148,N_40183);
and U43483 (N_43483,N_42355,N_41393);
nor U43484 (N_43484,N_42152,N_40913);
nand U43485 (N_43485,N_41735,N_40940);
and U43486 (N_43486,N_40954,N_40492);
or U43487 (N_43487,N_41332,N_41866);
or U43488 (N_43488,N_40117,N_40813);
nor U43489 (N_43489,N_41686,N_40904);
nand U43490 (N_43490,N_40452,N_41456);
and U43491 (N_43491,N_41814,N_40911);
and U43492 (N_43492,N_41927,N_41656);
xor U43493 (N_43493,N_41528,N_40590);
or U43494 (N_43494,N_40714,N_40887);
nand U43495 (N_43495,N_42019,N_42474);
nand U43496 (N_43496,N_41144,N_41689);
and U43497 (N_43497,N_40864,N_41976);
nor U43498 (N_43498,N_40685,N_40989);
or U43499 (N_43499,N_40875,N_40834);
nor U43500 (N_43500,N_40516,N_42494);
and U43501 (N_43501,N_41135,N_40333);
or U43502 (N_43502,N_40806,N_40696);
or U43503 (N_43503,N_41445,N_41290);
and U43504 (N_43504,N_40648,N_41088);
and U43505 (N_43505,N_41098,N_41472);
nand U43506 (N_43506,N_42096,N_41097);
or U43507 (N_43507,N_42024,N_40180);
nand U43508 (N_43508,N_42206,N_40160);
or U43509 (N_43509,N_41480,N_41889);
nand U43510 (N_43510,N_40796,N_40261);
xnor U43511 (N_43511,N_40191,N_40798);
or U43512 (N_43512,N_40381,N_42180);
or U43513 (N_43513,N_41737,N_42441);
or U43514 (N_43514,N_42247,N_41961);
or U43515 (N_43515,N_40179,N_41783);
nor U43516 (N_43516,N_41543,N_40865);
xnor U43517 (N_43517,N_41558,N_42107);
or U43518 (N_43518,N_40879,N_41637);
and U43519 (N_43519,N_40497,N_41627);
or U43520 (N_43520,N_41919,N_40936);
nor U43521 (N_43521,N_42431,N_41392);
xor U43522 (N_43522,N_41351,N_41473);
and U43523 (N_43523,N_41860,N_41105);
or U43524 (N_43524,N_42292,N_41966);
and U43525 (N_43525,N_41958,N_41273);
and U43526 (N_43526,N_40537,N_40824);
nand U43527 (N_43527,N_42258,N_40533);
nor U43528 (N_43528,N_41741,N_41159);
or U43529 (N_43529,N_40377,N_41885);
nor U43530 (N_43530,N_40238,N_41059);
and U43531 (N_43531,N_41128,N_40740);
xnor U43532 (N_43532,N_42404,N_41235);
and U43533 (N_43533,N_40662,N_40098);
xnor U43534 (N_43534,N_40442,N_41746);
or U43535 (N_43535,N_41713,N_40838);
or U43536 (N_43536,N_41423,N_41825);
and U43537 (N_43537,N_42149,N_40121);
nor U43538 (N_43538,N_41111,N_40579);
nor U43539 (N_43539,N_40691,N_41177);
or U43540 (N_43540,N_41620,N_42378);
nand U43541 (N_43541,N_40482,N_40174);
or U43542 (N_43542,N_41683,N_40061);
nor U43543 (N_43543,N_41297,N_42388);
xnor U43544 (N_43544,N_42339,N_40364);
or U43545 (N_43545,N_41280,N_40762);
nor U43546 (N_43546,N_42042,N_42269);
and U43547 (N_43547,N_41800,N_42318);
nand U43548 (N_43548,N_41583,N_41781);
or U43549 (N_43549,N_41258,N_41934);
xnor U43550 (N_43550,N_42347,N_41134);
nand U43551 (N_43551,N_41838,N_41440);
nand U43552 (N_43552,N_40500,N_40853);
xnor U43553 (N_43553,N_41029,N_40077);
nand U43554 (N_43554,N_40518,N_40227);
and U43555 (N_43555,N_40938,N_40633);
xnor U43556 (N_43556,N_41060,N_41080);
or U43557 (N_43557,N_40475,N_40597);
and U43558 (N_43558,N_40102,N_41422);
nor U43559 (N_43559,N_40253,N_40059);
xnor U43560 (N_43560,N_41131,N_41110);
and U43561 (N_43561,N_40213,N_40186);
nand U43562 (N_43562,N_42069,N_41626);
nand U43563 (N_43563,N_41599,N_41753);
nor U43564 (N_43564,N_41307,N_42455);
nand U43565 (N_43565,N_41731,N_40209);
nor U43566 (N_43566,N_42300,N_40353);
nor U43567 (N_43567,N_40530,N_40076);
xor U43568 (N_43568,N_40052,N_40279);
nor U43569 (N_43569,N_40757,N_41661);
nand U43570 (N_43570,N_41320,N_41489);
nor U43571 (N_43571,N_41765,N_42415);
nand U43572 (N_43572,N_40265,N_41106);
nand U43573 (N_43573,N_41167,N_41484);
or U43574 (N_43574,N_40173,N_40041);
nand U43575 (N_43575,N_41593,N_40831);
or U43576 (N_43576,N_41980,N_40100);
nor U43577 (N_43577,N_42109,N_42048);
nand U43578 (N_43578,N_42124,N_42082);
nand U43579 (N_43579,N_41028,N_41527);
or U43580 (N_43580,N_42274,N_41635);
nor U43581 (N_43581,N_40688,N_42479);
nor U43582 (N_43582,N_40181,N_40732);
xor U43583 (N_43583,N_40826,N_41296);
and U43584 (N_43584,N_41523,N_40222);
and U43585 (N_43585,N_40336,N_40357);
nor U43586 (N_43586,N_40067,N_42010);
and U43587 (N_43587,N_40724,N_40651);
and U43588 (N_43588,N_41301,N_40145);
xor U43589 (N_43589,N_41409,N_40784);
or U43590 (N_43590,N_41119,N_40917);
or U43591 (N_43591,N_40964,N_42452);
or U43592 (N_43592,N_41561,N_40224);
nand U43593 (N_43593,N_41137,N_41074);
xnor U43594 (N_43594,N_42045,N_42094);
and U43595 (N_43595,N_41500,N_42351);
or U43596 (N_43596,N_42456,N_40819);
xor U43597 (N_43597,N_40881,N_42444);
or U43598 (N_43598,N_40241,N_40617);
or U43599 (N_43599,N_41460,N_41429);
nand U43600 (N_43600,N_40244,N_41403);
and U43601 (N_43601,N_40394,N_40220);
and U43602 (N_43602,N_41999,N_40154);
and U43603 (N_43603,N_40415,N_41400);
and U43604 (N_43604,N_41538,N_40262);
nand U43605 (N_43605,N_40937,N_41056);
or U43606 (N_43606,N_42085,N_41211);
xor U43607 (N_43607,N_41009,N_40873);
and U43608 (N_43608,N_40783,N_40107);
or U43609 (N_43609,N_40162,N_41759);
nand U43610 (N_43610,N_41437,N_40065);
nor U43611 (N_43611,N_41103,N_40664);
and U43612 (N_43612,N_41986,N_41222);
nor U43613 (N_43613,N_41346,N_42100);
or U43614 (N_43614,N_40322,N_41146);
and U43615 (N_43615,N_40561,N_40433);
nor U43616 (N_43616,N_42187,N_42271);
or U43617 (N_43617,N_40101,N_40629);
and U43618 (N_43618,N_41318,N_41077);
nand U43619 (N_43619,N_40012,N_41739);
or U43620 (N_43620,N_40075,N_42462);
nand U43621 (N_43621,N_42140,N_41282);
nand U43622 (N_43622,N_41902,N_41972);
and U43623 (N_43623,N_41450,N_42399);
nor U43624 (N_43624,N_41153,N_41107);
nand U43625 (N_43625,N_40449,N_41390);
or U43626 (N_43626,N_40916,N_41415);
xor U43627 (N_43627,N_41931,N_41584);
and U43628 (N_43628,N_40028,N_41270);
and U43629 (N_43629,N_41503,N_41333);
xnor U43630 (N_43630,N_40805,N_41873);
or U43631 (N_43631,N_40086,N_42381);
or U43632 (N_43632,N_42000,N_41900);
or U43633 (N_43633,N_42344,N_41039);
nand U43634 (N_43634,N_41669,N_40402);
nor U43635 (N_43635,N_41170,N_40493);
or U43636 (N_43636,N_42093,N_40739);
and U43637 (N_43637,N_41264,N_40818);
or U43638 (N_43638,N_42164,N_40447);
xor U43639 (N_43639,N_41011,N_41100);
nor U43640 (N_43640,N_41323,N_42146);
nor U43641 (N_43641,N_41164,N_42235);
nand U43642 (N_43642,N_42170,N_41071);
or U43643 (N_43643,N_41454,N_41511);
nand U43644 (N_43644,N_40345,N_41747);
or U43645 (N_43645,N_41350,N_41821);
or U43646 (N_43646,N_42498,N_41557);
nor U43647 (N_43647,N_42014,N_40697);
nand U43648 (N_43648,N_42392,N_40999);
or U43649 (N_43649,N_41257,N_42056);
nand U43650 (N_43650,N_42337,N_40647);
nor U43651 (N_43651,N_41676,N_40748);
nand U43652 (N_43652,N_42054,N_41770);
nand U43653 (N_43653,N_40979,N_41481);
and U43654 (N_43654,N_42114,N_41916);
nand U43655 (N_43655,N_40192,N_42153);
nand U43656 (N_43656,N_41093,N_41702);
and U43657 (N_43657,N_42243,N_40944);
and U43658 (N_43658,N_40978,N_41073);
and U43659 (N_43659,N_42252,N_41673);
and U43660 (N_43660,N_40436,N_40093);
nand U43661 (N_43661,N_41260,N_41421);
or U43662 (N_43662,N_41419,N_41694);
and U43663 (N_43663,N_42143,N_40653);
and U43664 (N_43664,N_41548,N_40239);
and U43665 (N_43665,N_40350,N_40993);
and U43666 (N_43666,N_41360,N_40205);
xnor U43667 (N_43667,N_40888,N_41691);
nor U43668 (N_43668,N_40548,N_40275);
or U43669 (N_43669,N_40371,N_42078);
nor U43670 (N_43670,N_41508,N_40300);
and U43671 (N_43671,N_40462,N_41180);
nor U43672 (N_43672,N_40479,N_41240);
and U43673 (N_43673,N_41738,N_40219);
xor U43674 (N_43674,N_40681,N_42151);
xnor U43675 (N_43675,N_41929,N_42080);
nor U43676 (N_43676,N_40097,N_40047);
nand U43677 (N_43677,N_40155,N_40912);
or U43678 (N_43678,N_41155,N_41853);
xnor U43679 (N_43679,N_41768,N_40752);
and U43680 (N_43680,N_40151,N_41591);
xor U43681 (N_43681,N_41031,N_41820);
or U43682 (N_43682,N_41373,N_41380);
nand U43683 (N_43683,N_40305,N_41458);
nand U43684 (N_43684,N_41399,N_41010);
nand U43685 (N_43685,N_42320,N_41859);
and U43686 (N_43686,N_42150,N_41575);
nand U43687 (N_43687,N_42196,N_41547);
and U43688 (N_43688,N_40513,N_41588);
and U43689 (N_43689,N_40728,N_42041);
and U43690 (N_43690,N_42306,N_40427);
and U43691 (N_43691,N_40952,N_42104);
nand U43692 (N_43692,N_40945,N_41564);
nand U43693 (N_43693,N_42291,N_40288);
nor U43694 (N_43694,N_40667,N_40003);
nand U43695 (N_43695,N_41306,N_41477);
or U43696 (N_43696,N_42463,N_42426);
nor U43697 (N_43697,N_40246,N_41293);
and U43698 (N_43698,N_40013,N_41483);
nor U43699 (N_43699,N_42139,N_42053);
nor U43700 (N_43700,N_41262,N_42285);
or U43701 (N_43701,N_40247,N_41411);
nor U43702 (N_43702,N_42240,N_40570);
or U43703 (N_43703,N_42486,N_41224);
and U43704 (N_43704,N_40480,N_41226);
and U43705 (N_43705,N_41112,N_42405);
nor U43706 (N_43706,N_41837,N_41151);
nor U43707 (N_43707,N_41510,N_42072);
nor U43708 (N_43708,N_42175,N_41340);
nor U43709 (N_43709,N_41431,N_42199);
nor U43710 (N_43710,N_41816,N_42407);
and U43711 (N_43711,N_40257,N_40703);
nor U43712 (N_43712,N_41989,N_40124);
xnor U43713 (N_43713,N_40949,N_41789);
nand U43714 (N_43714,N_40080,N_42466);
nand U43715 (N_43715,N_41915,N_40455);
xor U43716 (N_43716,N_40113,N_41217);
nor U43717 (N_43717,N_42091,N_40339);
nand U43718 (N_43718,N_40951,N_42487);
xnor U43719 (N_43719,N_40094,N_41145);
and U43720 (N_43720,N_40995,N_41432);
and U43721 (N_43721,N_41336,N_41882);
or U43722 (N_43722,N_41605,N_41395);
or U43723 (N_43723,N_40895,N_40291);
and U43724 (N_43724,N_40448,N_41302);
and U43725 (N_43725,N_42329,N_40884);
nand U43726 (N_43726,N_40454,N_41305);
or U43727 (N_43727,N_41344,N_41607);
nand U43728 (N_43728,N_40132,N_40820);
nor U43729 (N_43729,N_41918,N_41238);
xnor U43730 (N_43730,N_42333,N_41331);
nor U43731 (N_43731,N_40431,N_41791);
nand U43732 (N_43732,N_40366,N_40808);
or U43733 (N_43733,N_41786,N_41129);
xnor U43734 (N_43734,N_41138,N_40407);
or U43735 (N_43735,N_40723,N_41259);
and U43736 (N_43736,N_40118,N_41846);
nor U43737 (N_43737,N_42236,N_41091);
nand U43738 (N_43738,N_42371,N_42158);
and U43739 (N_43739,N_42280,N_41276);
nor U43740 (N_43740,N_40127,N_41389);
nor U43741 (N_43741,N_40108,N_41651);
nand U43742 (N_43742,N_41516,N_41371);
nor U43743 (N_43743,N_41550,N_40386);
or U43744 (N_43744,N_41690,N_40635);
nor U43745 (N_43745,N_40850,N_41641);
or U43746 (N_43746,N_41140,N_40388);
nand U43747 (N_43747,N_40616,N_42430);
nand U43748 (N_43748,N_41688,N_40926);
nand U43749 (N_43749,N_41213,N_41701);
nor U43750 (N_43750,N_41813,N_41323);
and U43751 (N_43751,N_42217,N_42057);
xnor U43752 (N_43752,N_41383,N_41618);
nand U43753 (N_43753,N_40309,N_41867);
and U43754 (N_43754,N_40343,N_41777);
nor U43755 (N_43755,N_41201,N_40392);
and U43756 (N_43756,N_40217,N_41062);
or U43757 (N_43757,N_40776,N_41104);
nor U43758 (N_43758,N_42417,N_40242);
or U43759 (N_43759,N_41724,N_41097);
nor U43760 (N_43760,N_40228,N_42482);
or U43761 (N_43761,N_40697,N_40715);
or U43762 (N_43762,N_40295,N_42147);
nor U43763 (N_43763,N_41436,N_40648);
or U43764 (N_43764,N_42284,N_42280);
nand U43765 (N_43765,N_40041,N_40278);
nor U43766 (N_43766,N_41097,N_41277);
and U43767 (N_43767,N_40124,N_40837);
and U43768 (N_43768,N_40198,N_42108);
nor U43769 (N_43769,N_42089,N_40042);
or U43770 (N_43770,N_41301,N_40545);
or U43771 (N_43771,N_42076,N_41386);
xnor U43772 (N_43772,N_40341,N_40800);
or U43773 (N_43773,N_41293,N_40673);
and U43774 (N_43774,N_41926,N_40656);
nor U43775 (N_43775,N_41191,N_40293);
or U43776 (N_43776,N_41147,N_41156);
xor U43777 (N_43777,N_41838,N_40266);
or U43778 (N_43778,N_42371,N_41401);
and U43779 (N_43779,N_41510,N_40574);
nor U43780 (N_43780,N_40489,N_41214);
nor U43781 (N_43781,N_40881,N_41117);
and U43782 (N_43782,N_41362,N_41567);
or U43783 (N_43783,N_41417,N_41157);
or U43784 (N_43784,N_40086,N_42331);
or U43785 (N_43785,N_40597,N_41171);
or U43786 (N_43786,N_41410,N_41232);
nor U43787 (N_43787,N_41277,N_42264);
and U43788 (N_43788,N_42174,N_40045);
nor U43789 (N_43789,N_42281,N_41017);
or U43790 (N_43790,N_41472,N_40991);
and U43791 (N_43791,N_40071,N_41615);
and U43792 (N_43792,N_42255,N_40274);
and U43793 (N_43793,N_40420,N_41808);
or U43794 (N_43794,N_41382,N_41983);
nor U43795 (N_43795,N_40979,N_40003);
xnor U43796 (N_43796,N_40234,N_40104);
or U43797 (N_43797,N_41500,N_41662);
nor U43798 (N_43798,N_40479,N_41666);
nor U43799 (N_43799,N_41756,N_41159);
nand U43800 (N_43800,N_41705,N_40749);
nand U43801 (N_43801,N_42073,N_42252);
nor U43802 (N_43802,N_40806,N_41422);
nand U43803 (N_43803,N_41952,N_40237);
nand U43804 (N_43804,N_41042,N_41811);
and U43805 (N_43805,N_40414,N_41673);
xor U43806 (N_43806,N_40210,N_40036);
and U43807 (N_43807,N_40139,N_40208);
nand U43808 (N_43808,N_41537,N_41733);
nand U43809 (N_43809,N_41670,N_40748);
nand U43810 (N_43810,N_41295,N_41745);
nor U43811 (N_43811,N_41879,N_41600);
nand U43812 (N_43812,N_40902,N_40276);
nand U43813 (N_43813,N_41178,N_40515);
nor U43814 (N_43814,N_41427,N_42264);
and U43815 (N_43815,N_42099,N_42329);
xnor U43816 (N_43816,N_41683,N_41333);
or U43817 (N_43817,N_41702,N_41137);
nand U43818 (N_43818,N_40161,N_41666);
and U43819 (N_43819,N_40437,N_41813);
nand U43820 (N_43820,N_41292,N_40612);
nor U43821 (N_43821,N_41849,N_41111);
and U43822 (N_43822,N_41634,N_40010);
or U43823 (N_43823,N_40847,N_40804);
or U43824 (N_43824,N_40090,N_41987);
xnor U43825 (N_43825,N_40604,N_41671);
xnor U43826 (N_43826,N_40913,N_42072);
or U43827 (N_43827,N_40809,N_41716);
or U43828 (N_43828,N_40064,N_40805);
or U43829 (N_43829,N_42116,N_41430);
nor U43830 (N_43830,N_40084,N_41088);
xor U43831 (N_43831,N_41203,N_41490);
xnor U43832 (N_43832,N_41840,N_40913);
and U43833 (N_43833,N_40892,N_40012);
nand U43834 (N_43834,N_41726,N_42186);
and U43835 (N_43835,N_40301,N_42295);
nor U43836 (N_43836,N_40675,N_40915);
nand U43837 (N_43837,N_41936,N_40647);
or U43838 (N_43838,N_41305,N_40869);
or U43839 (N_43839,N_40080,N_40069);
or U43840 (N_43840,N_42285,N_42250);
or U43841 (N_43841,N_40609,N_40716);
or U43842 (N_43842,N_42408,N_40746);
nand U43843 (N_43843,N_41386,N_42192);
nand U43844 (N_43844,N_41140,N_41662);
nor U43845 (N_43845,N_40921,N_42233);
nor U43846 (N_43846,N_41194,N_40050);
and U43847 (N_43847,N_41264,N_40262);
xnor U43848 (N_43848,N_41783,N_41594);
xor U43849 (N_43849,N_42407,N_41718);
nor U43850 (N_43850,N_41768,N_41017);
nor U43851 (N_43851,N_40160,N_41719);
and U43852 (N_43852,N_40219,N_41930);
nor U43853 (N_43853,N_42122,N_42388);
and U43854 (N_43854,N_42462,N_41874);
and U43855 (N_43855,N_41154,N_42166);
xnor U43856 (N_43856,N_40610,N_40258);
nand U43857 (N_43857,N_41850,N_42250);
or U43858 (N_43858,N_41211,N_41144);
or U43859 (N_43859,N_40689,N_41908);
xnor U43860 (N_43860,N_42259,N_40825);
or U43861 (N_43861,N_41553,N_41295);
and U43862 (N_43862,N_42217,N_41178);
nand U43863 (N_43863,N_41622,N_41544);
and U43864 (N_43864,N_41522,N_40252);
nor U43865 (N_43865,N_42002,N_41921);
xnor U43866 (N_43866,N_40814,N_42384);
nor U43867 (N_43867,N_41585,N_41384);
and U43868 (N_43868,N_40863,N_42348);
nand U43869 (N_43869,N_42316,N_42234);
or U43870 (N_43870,N_40030,N_42162);
xnor U43871 (N_43871,N_41747,N_41628);
or U43872 (N_43872,N_42213,N_41492);
nand U43873 (N_43873,N_42353,N_40303);
and U43874 (N_43874,N_41421,N_41480);
and U43875 (N_43875,N_41383,N_41513);
and U43876 (N_43876,N_40404,N_40138);
nor U43877 (N_43877,N_42066,N_42409);
nand U43878 (N_43878,N_41689,N_40023);
and U43879 (N_43879,N_40777,N_42070);
xor U43880 (N_43880,N_40755,N_41616);
nor U43881 (N_43881,N_41882,N_42128);
nand U43882 (N_43882,N_40677,N_42205);
or U43883 (N_43883,N_41247,N_40036);
nand U43884 (N_43884,N_40586,N_41655);
xor U43885 (N_43885,N_40112,N_41109);
and U43886 (N_43886,N_42140,N_40627);
xor U43887 (N_43887,N_41492,N_41486);
and U43888 (N_43888,N_40046,N_42278);
and U43889 (N_43889,N_41855,N_41609);
or U43890 (N_43890,N_41729,N_40994);
and U43891 (N_43891,N_40965,N_40856);
and U43892 (N_43892,N_41569,N_41430);
xnor U43893 (N_43893,N_42348,N_41831);
nand U43894 (N_43894,N_40103,N_41769);
nand U43895 (N_43895,N_41298,N_41837);
and U43896 (N_43896,N_40980,N_42460);
nand U43897 (N_43897,N_41808,N_42452);
nor U43898 (N_43898,N_41402,N_40049);
or U43899 (N_43899,N_40913,N_41644);
and U43900 (N_43900,N_42263,N_41585);
or U43901 (N_43901,N_40913,N_40229);
xnor U43902 (N_43902,N_40246,N_41639);
xnor U43903 (N_43903,N_40267,N_40337);
nor U43904 (N_43904,N_40373,N_41168);
or U43905 (N_43905,N_40145,N_41057);
xor U43906 (N_43906,N_42244,N_42475);
nand U43907 (N_43907,N_42283,N_41282);
nor U43908 (N_43908,N_40365,N_41261);
nor U43909 (N_43909,N_41803,N_41004);
nand U43910 (N_43910,N_41057,N_40278);
or U43911 (N_43911,N_41489,N_40421);
nand U43912 (N_43912,N_41391,N_41114);
and U43913 (N_43913,N_42131,N_41811);
nand U43914 (N_43914,N_41694,N_40969);
nor U43915 (N_43915,N_40732,N_40617);
and U43916 (N_43916,N_42054,N_41810);
xnor U43917 (N_43917,N_40803,N_40571);
nor U43918 (N_43918,N_41495,N_40097);
xnor U43919 (N_43919,N_41172,N_42344);
nor U43920 (N_43920,N_40718,N_40153);
xnor U43921 (N_43921,N_40239,N_40172);
or U43922 (N_43922,N_40759,N_40725);
nor U43923 (N_43923,N_41393,N_42498);
or U43924 (N_43924,N_40761,N_41865);
and U43925 (N_43925,N_40868,N_40850);
nor U43926 (N_43926,N_41190,N_40889);
and U43927 (N_43927,N_40554,N_41003);
nor U43928 (N_43928,N_40982,N_41166);
or U43929 (N_43929,N_42392,N_41760);
nand U43930 (N_43930,N_40609,N_42374);
nand U43931 (N_43931,N_42405,N_40693);
or U43932 (N_43932,N_40171,N_41982);
and U43933 (N_43933,N_42396,N_40353);
nor U43934 (N_43934,N_40465,N_41343);
nor U43935 (N_43935,N_40790,N_40744);
nand U43936 (N_43936,N_40025,N_41769);
and U43937 (N_43937,N_42091,N_41818);
nand U43938 (N_43938,N_40193,N_41329);
and U43939 (N_43939,N_41574,N_42136);
nor U43940 (N_43940,N_42433,N_41620);
or U43941 (N_43941,N_40252,N_40609);
xnor U43942 (N_43942,N_42015,N_40504);
nor U43943 (N_43943,N_40389,N_40459);
and U43944 (N_43944,N_41716,N_40872);
nor U43945 (N_43945,N_41098,N_42423);
nand U43946 (N_43946,N_41052,N_40044);
xor U43947 (N_43947,N_40140,N_41668);
nor U43948 (N_43948,N_41946,N_40721);
and U43949 (N_43949,N_41769,N_40072);
xnor U43950 (N_43950,N_40981,N_40738);
or U43951 (N_43951,N_41596,N_40995);
nand U43952 (N_43952,N_40442,N_40275);
nor U43953 (N_43953,N_42485,N_41259);
nor U43954 (N_43954,N_42387,N_41112);
or U43955 (N_43955,N_42351,N_40762);
or U43956 (N_43956,N_40071,N_40729);
xnor U43957 (N_43957,N_42358,N_40381);
and U43958 (N_43958,N_41991,N_42179);
nand U43959 (N_43959,N_41993,N_40277);
nor U43960 (N_43960,N_41107,N_40496);
and U43961 (N_43961,N_40046,N_40389);
xor U43962 (N_43962,N_41364,N_40413);
nand U43963 (N_43963,N_40592,N_40940);
nand U43964 (N_43964,N_40468,N_41607);
nand U43965 (N_43965,N_41200,N_40205);
nand U43966 (N_43966,N_42112,N_40320);
nor U43967 (N_43967,N_42172,N_40447);
and U43968 (N_43968,N_40590,N_40365);
nand U43969 (N_43969,N_40815,N_41478);
or U43970 (N_43970,N_41014,N_41971);
xor U43971 (N_43971,N_42098,N_41840);
xor U43972 (N_43972,N_42339,N_41103);
nand U43973 (N_43973,N_42078,N_40132);
nand U43974 (N_43974,N_41606,N_40582);
and U43975 (N_43975,N_40650,N_41924);
or U43976 (N_43976,N_40383,N_40024);
or U43977 (N_43977,N_41516,N_41568);
nand U43978 (N_43978,N_42124,N_41703);
nand U43979 (N_43979,N_40871,N_42308);
nand U43980 (N_43980,N_40768,N_41489);
nand U43981 (N_43981,N_40154,N_41209);
nor U43982 (N_43982,N_42262,N_41124);
or U43983 (N_43983,N_41607,N_40629);
xnor U43984 (N_43984,N_42334,N_42430);
and U43985 (N_43985,N_41350,N_42378);
and U43986 (N_43986,N_41702,N_41913);
nand U43987 (N_43987,N_42231,N_41132);
nand U43988 (N_43988,N_40134,N_40271);
nor U43989 (N_43989,N_40926,N_41013);
or U43990 (N_43990,N_42234,N_41683);
nand U43991 (N_43991,N_40950,N_40369);
and U43992 (N_43992,N_41348,N_41814);
xnor U43993 (N_43993,N_40204,N_41784);
nand U43994 (N_43994,N_40187,N_41335);
or U43995 (N_43995,N_42384,N_42209);
nand U43996 (N_43996,N_40080,N_41214);
or U43997 (N_43997,N_42488,N_41675);
and U43998 (N_43998,N_41807,N_42390);
xnor U43999 (N_43999,N_40284,N_40031);
xor U44000 (N_44000,N_41946,N_42019);
and U44001 (N_44001,N_41123,N_40243);
nand U44002 (N_44002,N_42450,N_41206);
nor U44003 (N_44003,N_42098,N_40287);
nand U44004 (N_44004,N_41403,N_40612);
nor U44005 (N_44005,N_41691,N_42298);
nand U44006 (N_44006,N_40920,N_41672);
nor U44007 (N_44007,N_41442,N_42358);
or U44008 (N_44008,N_41093,N_40213);
or U44009 (N_44009,N_40033,N_40146);
or U44010 (N_44010,N_40788,N_41287);
and U44011 (N_44011,N_40028,N_40440);
nor U44012 (N_44012,N_40576,N_41991);
and U44013 (N_44013,N_41822,N_41621);
nor U44014 (N_44014,N_42355,N_40501);
nand U44015 (N_44015,N_42459,N_42367);
nor U44016 (N_44016,N_41566,N_41147);
nor U44017 (N_44017,N_41760,N_40381);
and U44018 (N_44018,N_40855,N_42410);
xnor U44019 (N_44019,N_42246,N_40942);
or U44020 (N_44020,N_41977,N_40607);
and U44021 (N_44021,N_40873,N_41618);
nand U44022 (N_44022,N_40392,N_42341);
nor U44023 (N_44023,N_41120,N_41770);
or U44024 (N_44024,N_40921,N_42031);
nor U44025 (N_44025,N_40393,N_41787);
and U44026 (N_44026,N_40418,N_41035);
or U44027 (N_44027,N_40925,N_40880);
nand U44028 (N_44028,N_40008,N_40199);
xnor U44029 (N_44029,N_40089,N_40977);
nor U44030 (N_44030,N_41281,N_41274);
and U44031 (N_44031,N_40220,N_41946);
or U44032 (N_44032,N_40243,N_42468);
nor U44033 (N_44033,N_41891,N_41368);
or U44034 (N_44034,N_40127,N_41664);
nand U44035 (N_44035,N_41256,N_40037);
nand U44036 (N_44036,N_40413,N_40261);
xor U44037 (N_44037,N_40371,N_40974);
and U44038 (N_44038,N_40956,N_40997);
nand U44039 (N_44039,N_40970,N_40874);
nor U44040 (N_44040,N_41521,N_40928);
nand U44041 (N_44041,N_41942,N_41943);
or U44042 (N_44042,N_42053,N_40317);
or U44043 (N_44043,N_41443,N_40733);
nand U44044 (N_44044,N_40790,N_42041);
and U44045 (N_44045,N_41764,N_41692);
and U44046 (N_44046,N_41866,N_41649);
xor U44047 (N_44047,N_41957,N_40656);
nor U44048 (N_44048,N_42496,N_40814);
nor U44049 (N_44049,N_40743,N_42163);
nand U44050 (N_44050,N_41615,N_42226);
and U44051 (N_44051,N_40413,N_41732);
xor U44052 (N_44052,N_41414,N_41455);
nand U44053 (N_44053,N_40559,N_40600);
nand U44054 (N_44054,N_40013,N_41755);
nor U44055 (N_44055,N_42134,N_41536);
xnor U44056 (N_44056,N_40670,N_41071);
or U44057 (N_44057,N_40820,N_41211);
xnor U44058 (N_44058,N_41972,N_42349);
nor U44059 (N_44059,N_41269,N_41400);
nand U44060 (N_44060,N_42119,N_40987);
nor U44061 (N_44061,N_42211,N_40260);
and U44062 (N_44062,N_42412,N_42251);
or U44063 (N_44063,N_41462,N_41473);
nand U44064 (N_44064,N_40522,N_42088);
xnor U44065 (N_44065,N_41437,N_40727);
nand U44066 (N_44066,N_41229,N_41591);
nand U44067 (N_44067,N_42336,N_41566);
and U44068 (N_44068,N_40779,N_42246);
xor U44069 (N_44069,N_41072,N_41938);
nor U44070 (N_44070,N_40291,N_40161);
nand U44071 (N_44071,N_40779,N_41620);
and U44072 (N_44072,N_41864,N_41510);
nand U44073 (N_44073,N_41736,N_42160);
nor U44074 (N_44074,N_42427,N_41078);
xor U44075 (N_44075,N_40212,N_41563);
and U44076 (N_44076,N_40015,N_41822);
or U44077 (N_44077,N_40268,N_40961);
nand U44078 (N_44078,N_42275,N_41996);
and U44079 (N_44079,N_41897,N_40452);
or U44080 (N_44080,N_41734,N_41286);
nor U44081 (N_44081,N_40802,N_40804);
nor U44082 (N_44082,N_41767,N_40344);
and U44083 (N_44083,N_41528,N_41558);
or U44084 (N_44084,N_40130,N_41572);
nor U44085 (N_44085,N_40482,N_40416);
nand U44086 (N_44086,N_41795,N_40626);
xor U44087 (N_44087,N_41506,N_41491);
nor U44088 (N_44088,N_40783,N_42017);
or U44089 (N_44089,N_41909,N_40604);
or U44090 (N_44090,N_42040,N_42315);
nand U44091 (N_44091,N_41537,N_41285);
nand U44092 (N_44092,N_40771,N_40473);
nor U44093 (N_44093,N_41670,N_40855);
nor U44094 (N_44094,N_41444,N_41956);
or U44095 (N_44095,N_42026,N_41004);
and U44096 (N_44096,N_40560,N_41170);
or U44097 (N_44097,N_40809,N_41693);
and U44098 (N_44098,N_40240,N_41291);
and U44099 (N_44099,N_40626,N_41073);
nor U44100 (N_44100,N_42194,N_41588);
nor U44101 (N_44101,N_41305,N_41124);
nand U44102 (N_44102,N_41287,N_40099);
and U44103 (N_44103,N_41537,N_40718);
nand U44104 (N_44104,N_41536,N_41952);
nor U44105 (N_44105,N_42153,N_40419);
nor U44106 (N_44106,N_41716,N_40130);
nand U44107 (N_44107,N_41679,N_41896);
nor U44108 (N_44108,N_40542,N_41635);
and U44109 (N_44109,N_42266,N_40081);
nand U44110 (N_44110,N_40515,N_41899);
nand U44111 (N_44111,N_40013,N_41928);
nor U44112 (N_44112,N_40523,N_41466);
nor U44113 (N_44113,N_41758,N_42465);
and U44114 (N_44114,N_41514,N_40728);
nand U44115 (N_44115,N_40711,N_41822);
and U44116 (N_44116,N_41392,N_42236);
xor U44117 (N_44117,N_41221,N_41197);
and U44118 (N_44118,N_42206,N_41848);
nor U44119 (N_44119,N_40638,N_41352);
nand U44120 (N_44120,N_40019,N_40926);
or U44121 (N_44121,N_40945,N_40322);
xor U44122 (N_44122,N_40159,N_42092);
and U44123 (N_44123,N_42026,N_41586);
xor U44124 (N_44124,N_42129,N_42415);
xor U44125 (N_44125,N_41229,N_42083);
or U44126 (N_44126,N_41652,N_42386);
and U44127 (N_44127,N_41940,N_40025);
and U44128 (N_44128,N_41835,N_42125);
nor U44129 (N_44129,N_41863,N_40491);
nor U44130 (N_44130,N_42082,N_41481);
nand U44131 (N_44131,N_41198,N_42287);
or U44132 (N_44132,N_41208,N_41012);
and U44133 (N_44133,N_41963,N_41762);
nand U44134 (N_44134,N_41712,N_42358);
nand U44135 (N_44135,N_42047,N_41783);
or U44136 (N_44136,N_41342,N_40034);
or U44137 (N_44137,N_40757,N_41273);
nor U44138 (N_44138,N_41848,N_40079);
and U44139 (N_44139,N_40646,N_40776);
nand U44140 (N_44140,N_41347,N_42157);
nand U44141 (N_44141,N_41568,N_42318);
and U44142 (N_44142,N_41057,N_41731);
nand U44143 (N_44143,N_40678,N_40139);
nor U44144 (N_44144,N_42265,N_40733);
and U44145 (N_44145,N_40625,N_41350);
or U44146 (N_44146,N_42114,N_40426);
or U44147 (N_44147,N_40112,N_42435);
nor U44148 (N_44148,N_41608,N_40257);
or U44149 (N_44149,N_40714,N_41420);
or U44150 (N_44150,N_40155,N_41561);
and U44151 (N_44151,N_41664,N_42399);
and U44152 (N_44152,N_42377,N_40609);
nor U44153 (N_44153,N_40322,N_40382);
nand U44154 (N_44154,N_42118,N_41242);
and U44155 (N_44155,N_42298,N_41382);
nand U44156 (N_44156,N_41713,N_40128);
nor U44157 (N_44157,N_41404,N_40343);
nand U44158 (N_44158,N_40263,N_42367);
nand U44159 (N_44159,N_41666,N_40430);
xnor U44160 (N_44160,N_40993,N_40641);
or U44161 (N_44161,N_41260,N_40270);
or U44162 (N_44162,N_42371,N_41611);
xnor U44163 (N_44163,N_41690,N_41013);
or U44164 (N_44164,N_40236,N_41818);
nand U44165 (N_44165,N_41965,N_41624);
nor U44166 (N_44166,N_42076,N_41410);
nand U44167 (N_44167,N_41626,N_40301);
nand U44168 (N_44168,N_40679,N_41090);
or U44169 (N_44169,N_42441,N_42391);
and U44170 (N_44170,N_41258,N_40786);
and U44171 (N_44171,N_40540,N_40133);
nand U44172 (N_44172,N_41839,N_41194);
or U44173 (N_44173,N_40839,N_40358);
or U44174 (N_44174,N_41281,N_42492);
nor U44175 (N_44175,N_41598,N_42250);
nand U44176 (N_44176,N_42044,N_41542);
and U44177 (N_44177,N_40574,N_41501);
nor U44178 (N_44178,N_40678,N_40689);
and U44179 (N_44179,N_40028,N_41000);
or U44180 (N_44180,N_41711,N_41145);
nor U44181 (N_44181,N_41310,N_41997);
and U44182 (N_44182,N_40031,N_40707);
or U44183 (N_44183,N_41486,N_41391);
or U44184 (N_44184,N_42282,N_41365);
xor U44185 (N_44185,N_41290,N_40621);
xnor U44186 (N_44186,N_42095,N_40310);
nand U44187 (N_44187,N_41789,N_40551);
xnor U44188 (N_44188,N_41325,N_42172);
xor U44189 (N_44189,N_40952,N_41075);
nor U44190 (N_44190,N_40705,N_41868);
nor U44191 (N_44191,N_41277,N_42029);
and U44192 (N_44192,N_42415,N_42043);
nand U44193 (N_44193,N_40047,N_40793);
nand U44194 (N_44194,N_42460,N_40879);
nand U44195 (N_44195,N_40071,N_40518);
or U44196 (N_44196,N_41869,N_41713);
and U44197 (N_44197,N_40733,N_41315);
xnor U44198 (N_44198,N_40136,N_42107);
nand U44199 (N_44199,N_41966,N_41531);
and U44200 (N_44200,N_42201,N_42224);
nor U44201 (N_44201,N_41128,N_41801);
nand U44202 (N_44202,N_40654,N_40585);
and U44203 (N_44203,N_40126,N_40345);
or U44204 (N_44204,N_41160,N_41664);
nor U44205 (N_44205,N_41197,N_40898);
xor U44206 (N_44206,N_40181,N_42094);
nor U44207 (N_44207,N_40622,N_42146);
xor U44208 (N_44208,N_41624,N_40637);
or U44209 (N_44209,N_41172,N_41779);
nand U44210 (N_44210,N_42271,N_40296);
and U44211 (N_44211,N_42425,N_40798);
nand U44212 (N_44212,N_41306,N_40048);
and U44213 (N_44213,N_40089,N_40264);
nor U44214 (N_44214,N_42047,N_42248);
nor U44215 (N_44215,N_40013,N_40814);
nand U44216 (N_44216,N_41363,N_42265);
and U44217 (N_44217,N_40137,N_42030);
and U44218 (N_44218,N_40530,N_40619);
or U44219 (N_44219,N_42203,N_41593);
nand U44220 (N_44220,N_41098,N_42006);
xor U44221 (N_44221,N_40298,N_40884);
xor U44222 (N_44222,N_41454,N_41530);
nand U44223 (N_44223,N_41884,N_41640);
and U44224 (N_44224,N_40500,N_40010);
or U44225 (N_44225,N_41447,N_40744);
or U44226 (N_44226,N_40698,N_41982);
and U44227 (N_44227,N_40830,N_40918);
nand U44228 (N_44228,N_40216,N_40386);
or U44229 (N_44229,N_40577,N_41576);
nor U44230 (N_44230,N_42064,N_41192);
and U44231 (N_44231,N_41378,N_41260);
nand U44232 (N_44232,N_42040,N_40869);
nand U44233 (N_44233,N_40464,N_40748);
nand U44234 (N_44234,N_41119,N_40088);
nor U44235 (N_44235,N_41202,N_40822);
and U44236 (N_44236,N_42284,N_40956);
or U44237 (N_44237,N_40603,N_40944);
nor U44238 (N_44238,N_40158,N_40823);
nor U44239 (N_44239,N_42012,N_42004);
or U44240 (N_44240,N_41253,N_40638);
nand U44241 (N_44241,N_42203,N_41799);
or U44242 (N_44242,N_40116,N_40110);
and U44243 (N_44243,N_41779,N_42325);
or U44244 (N_44244,N_42405,N_42465);
or U44245 (N_44245,N_40152,N_40113);
or U44246 (N_44246,N_40023,N_42068);
and U44247 (N_44247,N_40607,N_41102);
and U44248 (N_44248,N_41083,N_40155);
nor U44249 (N_44249,N_40538,N_42173);
and U44250 (N_44250,N_41233,N_40530);
nor U44251 (N_44251,N_41971,N_41320);
or U44252 (N_44252,N_42127,N_40121);
nor U44253 (N_44253,N_42143,N_41964);
and U44254 (N_44254,N_41273,N_40177);
nand U44255 (N_44255,N_40426,N_41434);
or U44256 (N_44256,N_41374,N_40706);
nand U44257 (N_44257,N_41739,N_40034);
and U44258 (N_44258,N_40743,N_41414);
or U44259 (N_44259,N_40976,N_41364);
nand U44260 (N_44260,N_42272,N_40751);
nand U44261 (N_44261,N_41444,N_40183);
nor U44262 (N_44262,N_42121,N_41936);
or U44263 (N_44263,N_40293,N_41881);
and U44264 (N_44264,N_41139,N_41174);
nand U44265 (N_44265,N_40280,N_40426);
or U44266 (N_44266,N_41485,N_41114);
nor U44267 (N_44267,N_42225,N_42493);
nand U44268 (N_44268,N_41600,N_42237);
nor U44269 (N_44269,N_40152,N_42482);
and U44270 (N_44270,N_41008,N_41707);
and U44271 (N_44271,N_41413,N_41543);
and U44272 (N_44272,N_42264,N_42115);
nor U44273 (N_44273,N_40617,N_42135);
nand U44274 (N_44274,N_41160,N_41574);
or U44275 (N_44275,N_40636,N_41966);
and U44276 (N_44276,N_40215,N_40717);
nand U44277 (N_44277,N_41431,N_40202);
or U44278 (N_44278,N_40424,N_40897);
nor U44279 (N_44279,N_40521,N_40111);
or U44280 (N_44280,N_40989,N_41588);
nor U44281 (N_44281,N_41155,N_41866);
and U44282 (N_44282,N_41837,N_41974);
and U44283 (N_44283,N_40381,N_41399);
nand U44284 (N_44284,N_42254,N_40363);
nor U44285 (N_44285,N_40820,N_40212);
nor U44286 (N_44286,N_41961,N_41572);
nand U44287 (N_44287,N_40246,N_41976);
nor U44288 (N_44288,N_40157,N_40819);
nor U44289 (N_44289,N_40149,N_40960);
and U44290 (N_44290,N_42076,N_42266);
nand U44291 (N_44291,N_42269,N_40973);
nor U44292 (N_44292,N_40618,N_41118);
xnor U44293 (N_44293,N_40440,N_40781);
nand U44294 (N_44294,N_41994,N_41153);
nand U44295 (N_44295,N_40640,N_41223);
and U44296 (N_44296,N_41512,N_40414);
nand U44297 (N_44297,N_41979,N_40465);
nand U44298 (N_44298,N_40215,N_40186);
nand U44299 (N_44299,N_41783,N_41050);
and U44300 (N_44300,N_42222,N_41617);
or U44301 (N_44301,N_40343,N_40997);
nor U44302 (N_44302,N_40477,N_41892);
or U44303 (N_44303,N_41058,N_40492);
and U44304 (N_44304,N_40783,N_40041);
or U44305 (N_44305,N_41319,N_41167);
nand U44306 (N_44306,N_40220,N_40967);
xnor U44307 (N_44307,N_42289,N_40503);
nand U44308 (N_44308,N_42078,N_41895);
nor U44309 (N_44309,N_41930,N_41934);
nor U44310 (N_44310,N_41221,N_40432);
and U44311 (N_44311,N_40659,N_41860);
xor U44312 (N_44312,N_40922,N_40127);
nor U44313 (N_44313,N_41681,N_41785);
nand U44314 (N_44314,N_41959,N_41634);
xnor U44315 (N_44315,N_41698,N_40628);
nand U44316 (N_44316,N_40888,N_40328);
nand U44317 (N_44317,N_41649,N_40160);
nor U44318 (N_44318,N_41088,N_40913);
nor U44319 (N_44319,N_42134,N_41947);
nor U44320 (N_44320,N_40312,N_42008);
and U44321 (N_44321,N_40700,N_40332);
nand U44322 (N_44322,N_40750,N_42148);
and U44323 (N_44323,N_42497,N_41603);
or U44324 (N_44324,N_40091,N_40304);
nor U44325 (N_44325,N_40876,N_42413);
and U44326 (N_44326,N_41673,N_42295);
nand U44327 (N_44327,N_40456,N_40320);
nor U44328 (N_44328,N_42261,N_40003);
and U44329 (N_44329,N_42150,N_41963);
nand U44330 (N_44330,N_40035,N_41361);
nand U44331 (N_44331,N_40548,N_40989);
and U44332 (N_44332,N_40090,N_40134);
xor U44333 (N_44333,N_40838,N_40762);
and U44334 (N_44334,N_40286,N_41273);
or U44335 (N_44335,N_40063,N_42355);
nor U44336 (N_44336,N_41256,N_42145);
nand U44337 (N_44337,N_40616,N_40373);
or U44338 (N_44338,N_41711,N_41156);
nor U44339 (N_44339,N_41294,N_40910);
and U44340 (N_44340,N_40161,N_40670);
and U44341 (N_44341,N_41799,N_40597);
nor U44342 (N_44342,N_40473,N_40776);
xnor U44343 (N_44343,N_41154,N_40220);
nand U44344 (N_44344,N_41291,N_41399);
nand U44345 (N_44345,N_40829,N_40164);
nand U44346 (N_44346,N_40737,N_42459);
nand U44347 (N_44347,N_40397,N_41406);
or U44348 (N_44348,N_41278,N_40859);
nor U44349 (N_44349,N_40840,N_41858);
nor U44350 (N_44350,N_42399,N_40722);
or U44351 (N_44351,N_41136,N_40532);
or U44352 (N_44352,N_40203,N_40701);
nand U44353 (N_44353,N_41552,N_41120);
nand U44354 (N_44354,N_40948,N_40104);
nor U44355 (N_44355,N_40098,N_41924);
or U44356 (N_44356,N_41271,N_41023);
nor U44357 (N_44357,N_40781,N_40506);
or U44358 (N_44358,N_41399,N_42418);
and U44359 (N_44359,N_40361,N_40789);
or U44360 (N_44360,N_40600,N_40337);
nor U44361 (N_44361,N_40858,N_40491);
nor U44362 (N_44362,N_40554,N_40117);
and U44363 (N_44363,N_42200,N_41237);
and U44364 (N_44364,N_41317,N_42044);
and U44365 (N_44365,N_41686,N_41892);
or U44366 (N_44366,N_41319,N_41342);
or U44367 (N_44367,N_40028,N_41500);
nor U44368 (N_44368,N_42237,N_41313);
or U44369 (N_44369,N_42310,N_40008);
or U44370 (N_44370,N_40535,N_42484);
and U44371 (N_44371,N_40360,N_41213);
xnor U44372 (N_44372,N_40547,N_40030);
nor U44373 (N_44373,N_41400,N_40310);
and U44374 (N_44374,N_40665,N_40892);
or U44375 (N_44375,N_40978,N_40268);
nand U44376 (N_44376,N_40764,N_40224);
nand U44377 (N_44377,N_40451,N_40072);
nor U44378 (N_44378,N_42151,N_41173);
or U44379 (N_44379,N_40758,N_40457);
or U44380 (N_44380,N_40758,N_42314);
xor U44381 (N_44381,N_40103,N_41851);
xnor U44382 (N_44382,N_41525,N_40107);
nand U44383 (N_44383,N_40438,N_40499);
and U44384 (N_44384,N_42090,N_41927);
xor U44385 (N_44385,N_40608,N_40106);
and U44386 (N_44386,N_41610,N_42082);
nand U44387 (N_44387,N_42082,N_42163);
and U44388 (N_44388,N_40005,N_41935);
and U44389 (N_44389,N_40785,N_40541);
nor U44390 (N_44390,N_40668,N_42120);
and U44391 (N_44391,N_41342,N_40075);
and U44392 (N_44392,N_41939,N_41198);
or U44393 (N_44393,N_41736,N_41322);
or U44394 (N_44394,N_42154,N_42001);
or U44395 (N_44395,N_41956,N_40546);
or U44396 (N_44396,N_42280,N_40849);
nor U44397 (N_44397,N_42010,N_40917);
or U44398 (N_44398,N_42221,N_41913);
nand U44399 (N_44399,N_42109,N_42085);
and U44400 (N_44400,N_41105,N_41050);
nor U44401 (N_44401,N_40240,N_42350);
and U44402 (N_44402,N_41592,N_40383);
xnor U44403 (N_44403,N_41150,N_42391);
or U44404 (N_44404,N_42085,N_40692);
xor U44405 (N_44405,N_42113,N_40307);
nor U44406 (N_44406,N_41332,N_42114);
and U44407 (N_44407,N_41407,N_42142);
and U44408 (N_44408,N_42243,N_41369);
nand U44409 (N_44409,N_40657,N_42340);
and U44410 (N_44410,N_41665,N_40531);
nor U44411 (N_44411,N_41697,N_40339);
and U44412 (N_44412,N_41771,N_42279);
or U44413 (N_44413,N_42111,N_42104);
xor U44414 (N_44414,N_42089,N_41639);
and U44415 (N_44415,N_41547,N_40220);
and U44416 (N_44416,N_41321,N_40590);
nand U44417 (N_44417,N_42467,N_41095);
nand U44418 (N_44418,N_41165,N_41005);
or U44419 (N_44419,N_40353,N_40126);
or U44420 (N_44420,N_41275,N_42442);
or U44421 (N_44421,N_41319,N_42382);
and U44422 (N_44422,N_40546,N_41829);
nor U44423 (N_44423,N_41581,N_40792);
or U44424 (N_44424,N_41662,N_41879);
and U44425 (N_44425,N_41043,N_41169);
and U44426 (N_44426,N_41434,N_41284);
nor U44427 (N_44427,N_41325,N_42292);
or U44428 (N_44428,N_40323,N_41076);
or U44429 (N_44429,N_41669,N_40137);
nand U44430 (N_44430,N_41128,N_42366);
and U44431 (N_44431,N_41910,N_40333);
nand U44432 (N_44432,N_40052,N_40059);
or U44433 (N_44433,N_40742,N_40455);
nand U44434 (N_44434,N_42264,N_42242);
and U44435 (N_44435,N_41860,N_41653);
or U44436 (N_44436,N_40638,N_42331);
nand U44437 (N_44437,N_40708,N_42021);
and U44438 (N_44438,N_42049,N_40831);
xor U44439 (N_44439,N_41338,N_42310);
nand U44440 (N_44440,N_41749,N_40881);
nor U44441 (N_44441,N_40297,N_41067);
nand U44442 (N_44442,N_42490,N_42469);
nand U44443 (N_44443,N_40209,N_41028);
or U44444 (N_44444,N_41170,N_41678);
nand U44445 (N_44445,N_40849,N_40560);
xor U44446 (N_44446,N_42180,N_41532);
nand U44447 (N_44447,N_40532,N_40770);
and U44448 (N_44448,N_40223,N_41461);
nand U44449 (N_44449,N_40968,N_41684);
nor U44450 (N_44450,N_40479,N_41677);
or U44451 (N_44451,N_40538,N_41551);
xor U44452 (N_44452,N_42231,N_41052);
or U44453 (N_44453,N_40296,N_40850);
nand U44454 (N_44454,N_40261,N_40678);
xor U44455 (N_44455,N_41589,N_41031);
nor U44456 (N_44456,N_40535,N_40135);
nor U44457 (N_44457,N_40199,N_41571);
nor U44458 (N_44458,N_42112,N_41453);
nand U44459 (N_44459,N_41770,N_42467);
nor U44460 (N_44460,N_40189,N_40782);
and U44461 (N_44461,N_41584,N_40361);
nand U44462 (N_44462,N_41413,N_41633);
or U44463 (N_44463,N_40309,N_41856);
or U44464 (N_44464,N_41307,N_41934);
and U44465 (N_44465,N_40042,N_40421);
nor U44466 (N_44466,N_40646,N_40100);
nor U44467 (N_44467,N_40895,N_40574);
and U44468 (N_44468,N_41196,N_41953);
nand U44469 (N_44469,N_42050,N_40716);
or U44470 (N_44470,N_42421,N_40457);
xnor U44471 (N_44471,N_41539,N_40849);
nor U44472 (N_44472,N_40281,N_42413);
and U44473 (N_44473,N_40061,N_41633);
xor U44474 (N_44474,N_41737,N_41885);
or U44475 (N_44475,N_40874,N_41241);
or U44476 (N_44476,N_41180,N_40827);
xnor U44477 (N_44477,N_42456,N_40506);
nand U44478 (N_44478,N_40851,N_41032);
or U44479 (N_44479,N_40539,N_42422);
and U44480 (N_44480,N_41656,N_41859);
nor U44481 (N_44481,N_41798,N_41575);
and U44482 (N_44482,N_41010,N_42312);
or U44483 (N_44483,N_40122,N_42187);
nor U44484 (N_44484,N_42034,N_40140);
nor U44485 (N_44485,N_41504,N_41514);
or U44486 (N_44486,N_41587,N_40075);
and U44487 (N_44487,N_41077,N_42423);
nand U44488 (N_44488,N_42016,N_41088);
nor U44489 (N_44489,N_41535,N_41858);
nor U44490 (N_44490,N_40657,N_40651);
xor U44491 (N_44491,N_41136,N_40505);
nand U44492 (N_44492,N_41235,N_41744);
nand U44493 (N_44493,N_42328,N_42160);
or U44494 (N_44494,N_40953,N_41972);
and U44495 (N_44495,N_42480,N_40646);
or U44496 (N_44496,N_40986,N_40967);
or U44497 (N_44497,N_41832,N_41397);
or U44498 (N_44498,N_41000,N_41999);
and U44499 (N_44499,N_41626,N_40739);
nand U44500 (N_44500,N_41205,N_41268);
xor U44501 (N_44501,N_40150,N_41464);
nand U44502 (N_44502,N_41277,N_40041);
nand U44503 (N_44503,N_41200,N_41520);
or U44504 (N_44504,N_41865,N_42247);
nor U44505 (N_44505,N_40725,N_41777);
xnor U44506 (N_44506,N_40895,N_40251);
and U44507 (N_44507,N_40411,N_41212);
nor U44508 (N_44508,N_41514,N_41334);
nand U44509 (N_44509,N_42087,N_40501);
nand U44510 (N_44510,N_41253,N_42128);
or U44511 (N_44511,N_41299,N_41901);
nor U44512 (N_44512,N_42305,N_40085);
nor U44513 (N_44513,N_41333,N_42333);
nor U44514 (N_44514,N_40635,N_41319);
xor U44515 (N_44515,N_41261,N_41021);
nor U44516 (N_44516,N_41618,N_40567);
or U44517 (N_44517,N_41507,N_41504);
or U44518 (N_44518,N_40684,N_41968);
or U44519 (N_44519,N_40804,N_41628);
and U44520 (N_44520,N_42178,N_42385);
nor U44521 (N_44521,N_40860,N_40162);
nand U44522 (N_44522,N_41522,N_41166);
nor U44523 (N_44523,N_42355,N_40943);
or U44524 (N_44524,N_42358,N_40201);
nor U44525 (N_44525,N_40346,N_41106);
nand U44526 (N_44526,N_40513,N_41655);
xor U44527 (N_44527,N_41747,N_40093);
nand U44528 (N_44528,N_41999,N_42185);
nand U44529 (N_44529,N_40360,N_40272);
and U44530 (N_44530,N_42104,N_41927);
nand U44531 (N_44531,N_42311,N_42252);
nand U44532 (N_44532,N_40806,N_40539);
nand U44533 (N_44533,N_41766,N_41455);
nand U44534 (N_44534,N_42010,N_41022);
nand U44535 (N_44535,N_41822,N_40619);
or U44536 (N_44536,N_41652,N_42344);
nor U44537 (N_44537,N_41283,N_40846);
or U44538 (N_44538,N_41944,N_41535);
or U44539 (N_44539,N_40080,N_40855);
or U44540 (N_44540,N_41506,N_40385);
nor U44541 (N_44541,N_40184,N_40594);
and U44542 (N_44542,N_40628,N_41818);
or U44543 (N_44543,N_41358,N_42024);
nor U44544 (N_44544,N_40390,N_42151);
nor U44545 (N_44545,N_41760,N_41343);
and U44546 (N_44546,N_40896,N_42111);
xnor U44547 (N_44547,N_41613,N_40658);
xnor U44548 (N_44548,N_40288,N_40170);
nand U44549 (N_44549,N_40304,N_41470);
and U44550 (N_44550,N_41192,N_42046);
xnor U44551 (N_44551,N_41769,N_41496);
xor U44552 (N_44552,N_40984,N_42260);
nor U44553 (N_44553,N_42415,N_41518);
and U44554 (N_44554,N_41544,N_40360);
nor U44555 (N_44555,N_41130,N_40505);
and U44556 (N_44556,N_41348,N_40188);
xor U44557 (N_44557,N_41165,N_40411);
nor U44558 (N_44558,N_41361,N_41429);
xnor U44559 (N_44559,N_41039,N_40553);
and U44560 (N_44560,N_41654,N_42347);
nor U44561 (N_44561,N_40568,N_41337);
nor U44562 (N_44562,N_40520,N_40282);
nand U44563 (N_44563,N_41410,N_40453);
nand U44564 (N_44564,N_40713,N_40498);
or U44565 (N_44565,N_42152,N_41709);
nand U44566 (N_44566,N_41191,N_41547);
or U44567 (N_44567,N_42490,N_42386);
nand U44568 (N_44568,N_40385,N_40856);
or U44569 (N_44569,N_40338,N_41218);
xnor U44570 (N_44570,N_41001,N_40609);
or U44571 (N_44571,N_40017,N_40548);
nor U44572 (N_44572,N_40562,N_40065);
xnor U44573 (N_44573,N_41257,N_40471);
nor U44574 (N_44574,N_41273,N_40844);
or U44575 (N_44575,N_41801,N_41314);
nor U44576 (N_44576,N_40996,N_42049);
nand U44577 (N_44577,N_42191,N_40712);
nand U44578 (N_44578,N_41860,N_41722);
nor U44579 (N_44579,N_41429,N_42231);
nand U44580 (N_44580,N_40765,N_40043);
xnor U44581 (N_44581,N_40381,N_41905);
or U44582 (N_44582,N_40115,N_40981);
nand U44583 (N_44583,N_40062,N_41911);
nor U44584 (N_44584,N_42225,N_40763);
nor U44585 (N_44585,N_42319,N_40645);
and U44586 (N_44586,N_41477,N_40386);
nor U44587 (N_44587,N_42095,N_42362);
or U44588 (N_44588,N_41469,N_41733);
xor U44589 (N_44589,N_40612,N_40987);
or U44590 (N_44590,N_42368,N_41468);
xnor U44591 (N_44591,N_41059,N_41093);
or U44592 (N_44592,N_41203,N_42334);
and U44593 (N_44593,N_40969,N_42309);
and U44594 (N_44594,N_41789,N_42080);
nand U44595 (N_44595,N_40190,N_40427);
and U44596 (N_44596,N_41962,N_42336);
xor U44597 (N_44597,N_40720,N_41927);
or U44598 (N_44598,N_40526,N_41672);
and U44599 (N_44599,N_40141,N_40066);
or U44600 (N_44600,N_40452,N_41331);
nor U44601 (N_44601,N_41521,N_40878);
and U44602 (N_44602,N_41188,N_42373);
xnor U44603 (N_44603,N_41139,N_40839);
nand U44604 (N_44604,N_40331,N_41434);
or U44605 (N_44605,N_42270,N_40566);
or U44606 (N_44606,N_40039,N_40140);
and U44607 (N_44607,N_40870,N_41394);
xor U44608 (N_44608,N_41188,N_41521);
and U44609 (N_44609,N_41719,N_40506);
nor U44610 (N_44610,N_40668,N_40968);
or U44611 (N_44611,N_40627,N_40874);
nor U44612 (N_44612,N_42112,N_41527);
and U44613 (N_44613,N_40401,N_42392);
nor U44614 (N_44614,N_41513,N_40321);
nand U44615 (N_44615,N_42209,N_41595);
and U44616 (N_44616,N_40938,N_41756);
nor U44617 (N_44617,N_41934,N_41381);
nand U44618 (N_44618,N_40808,N_40815);
and U44619 (N_44619,N_40398,N_42007);
nand U44620 (N_44620,N_40283,N_41183);
or U44621 (N_44621,N_41340,N_41615);
and U44622 (N_44622,N_41123,N_40286);
nor U44623 (N_44623,N_41662,N_40698);
nor U44624 (N_44624,N_40296,N_41567);
nor U44625 (N_44625,N_41343,N_41096);
nand U44626 (N_44626,N_42029,N_42378);
nor U44627 (N_44627,N_40205,N_40045);
and U44628 (N_44628,N_41799,N_40066);
nand U44629 (N_44629,N_40808,N_41337);
nand U44630 (N_44630,N_40132,N_42417);
nand U44631 (N_44631,N_40520,N_40973);
xor U44632 (N_44632,N_40728,N_42477);
xnor U44633 (N_44633,N_40457,N_40079);
and U44634 (N_44634,N_40428,N_41529);
or U44635 (N_44635,N_41662,N_42223);
and U44636 (N_44636,N_42306,N_41909);
nand U44637 (N_44637,N_40261,N_41702);
nand U44638 (N_44638,N_40871,N_41671);
nand U44639 (N_44639,N_41462,N_42361);
nand U44640 (N_44640,N_41480,N_41860);
or U44641 (N_44641,N_42029,N_41493);
and U44642 (N_44642,N_42416,N_41865);
or U44643 (N_44643,N_40199,N_41035);
and U44644 (N_44644,N_42129,N_41934);
and U44645 (N_44645,N_41934,N_40968);
xnor U44646 (N_44646,N_40516,N_42260);
nor U44647 (N_44647,N_41866,N_42303);
nand U44648 (N_44648,N_41088,N_42288);
nand U44649 (N_44649,N_41790,N_42112);
nor U44650 (N_44650,N_40237,N_41941);
and U44651 (N_44651,N_42290,N_42134);
and U44652 (N_44652,N_40232,N_41011);
nor U44653 (N_44653,N_42473,N_41759);
and U44654 (N_44654,N_40621,N_40812);
or U44655 (N_44655,N_40676,N_41026);
nor U44656 (N_44656,N_42072,N_42247);
and U44657 (N_44657,N_40838,N_41407);
or U44658 (N_44658,N_41288,N_41730);
xor U44659 (N_44659,N_41135,N_40674);
and U44660 (N_44660,N_40671,N_42455);
nand U44661 (N_44661,N_42002,N_41237);
nand U44662 (N_44662,N_41844,N_42444);
and U44663 (N_44663,N_42154,N_40638);
nand U44664 (N_44664,N_41659,N_41863);
and U44665 (N_44665,N_42280,N_41560);
nor U44666 (N_44666,N_42479,N_41328);
or U44667 (N_44667,N_41769,N_41295);
nand U44668 (N_44668,N_42393,N_40475);
nand U44669 (N_44669,N_41620,N_41665);
nand U44670 (N_44670,N_40763,N_42438);
nand U44671 (N_44671,N_41645,N_41402);
or U44672 (N_44672,N_41588,N_41435);
nand U44673 (N_44673,N_40210,N_41378);
nor U44674 (N_44674,N_40346,N_40614);
or U44675 (N_44675,N_40138,N_40805);
or U44676 (N_44676,N_42474,N_41378);
or U44677 (N_44677,N_40799,N_40460);
or U44678 (N_44678,N_40717,N_42178);
nor U44679 (N_44679,N_41687,N_41734);
nand U44680 (N_44680,N_41090,N_41700);
and U44681 (N_44681,N_41484,N_41999);
or U44682 (N_44682,N_40499,N_40609);
xor U44683 (N_44683,N_42210,N_40366);
and U44684 (N_44684,N_42174,N_42187);
nand U44685 (N_44685,N_41540,N_41170);
nand U44686 (N_44686,N_41348,N_41432);
nor U44687 (N_44687,N_40355,N_40641);
nand U44688 (N_44688,N_40554,N_41669);
or U44689 (N_44689,N_41761,N_41960);
or U44690 (N_44690,N_41653,N_40030);
or U44691 (N_44691,N_40845,N_40656);
nand U44692 (N_44692,N_40469,N_42139);
and U44693 (N_44693,N_41114,N_42439);
nor U44694 (N_44694,N_41101,N_42320);
and U44695 (N_44695,N_40904,N_42362);
and U44696 (N_44696,N_42083,N_41415);
and U44697 (N_44697,N_41361,N_41563);
nand U44698 (N_44698,N_42446,N_40237);
or U44699 (N_44699,N_40133,N_42119);
nand U44700 (N_44700,N_40784,N_41370);
nand U44701 (N_44701,N_41979,N_40306);
and U44702 (N_44702,N_42106,N_40276);
and U44703 (N_44703,N_42282,N_42438);
nand U44704 (N_44704,N_40894,N_41724);
nand U44705 (N_44705,N_41552,N_42361);
nand U44706 (N_44706,N_41368,N_40364);
or U44707 (N_44707,N_41972,N_41973);
nor U44708 (N_44708,N_41389,N_41048);
or U44709 (N_44709,N_42151,N_41736);
and U44710 (N_44710,N_42039,N_40822);
or U44711 (N_44711,N_41866,N_41114);
nand U44712 (N_44712,N_40985,N_41521);
and U44713 (N_44713,N_41809,N_41815);
nor U44714 (N_44714,N_41405,N_41184);
or U44715 (N_44715,N_40636,N_41172);
and U44716 (N_44716,N_40151,N_40828);
nand U44717 (N_44717,N_40810,N_40765);
and U44718 (N_44718,N_40287,N_42429);
nor U44719 (N_44719,N_42379,N_40793);
and U44720 (N_44720,N_41049,N_40175);
and U44721 (N_44721,N_40423,N_41715);
nor U44722 (N_44722,N_42351,N_41196);
and U44723 (N_44723,N_41529,N_40335);
and U44724 (N_44724,N_40647,N_40380);
or U44725 (N_44725,N_42457,N_41089);
nand U44726 (N_44726,N_40728,N_40706);
nor U44727 (N_44727,N_41127,N_40185);
nand U44728 (N_44728,N_42212,N_42047);
nand U44729 (N_44729,N_42470,N_40893);
nor U44730 (N_44730,N_41687,N_41690);
or U44731 (N_44731,N_40352,N_40019);
nor U44732 (N_44732,N_40937,N_40343);
nor U44733 (N_44733,N_40858,N_40232);
nor U44734 (N_44734,N_42388,N_41576);
or U44735 (N_44735,N_41844,N_40182);
and U44736 (N_44736,N_41444,N_41241);
nor U44737 (N_44737,N_40379,N_42145);
or U44738 (N_44738,N_41531,N_41274);
or U44739 (N_44739,N_40635,N_40391);
xnor U44740 (N_44740,N_41399,N_41930);
and U44741 (N_44741,N_42062,N_40537);
and U44742 (N_44742,N_41216,N_41975);
or U44743 (N_44743,N_41514,N_40999);
or U44744 (N_44744,N_41501,N_40845);
xnor U44745 (N_44745,N_41412,N_42315);
nand U44746 (N_44746,N_41496,N_41209);
nor U44747 (N_44747,N_40205,N_41794);
and U44748 (N_44748,N_41920,N_40424);
or U44749 (N_44749,N_41800,N_41598);
and U44750 (N_44750,N_41302,N_40338);
or U44751 (N_44751,N_41310,N_40811);
and U44752 (N_44752,N_40053,N_41615);
and U44753 (N_44753,N_41297,N_42463);
and U44754 (N_44754,N_41708,N_41934);
nand U44755 (N_44755,N_40242,N_40748);
or U44756 (N_44756,N_40343,N_40602);
nor U44757 (N_44757,N_42145,N_41868);
and U44758 (N_44758,N_40087,N_40585);
nand U44759 (N_44759,N_41658,N_42156);
nor U44760 (N_44760,N_40026,N_41785);
or U44761 (N_44761,N_42058,N_41175);
nand U44762 (N_44762,N_42000,N_40640);
nand U44763 (N_44763,N_40348,N_41980);
or U44764 (N_44764,N_40480,N_42481);
nor U44765 (N_44765,N_40822,N_40656);
xor U44766 (N_44766,N_41535,N_41997);
and U44767 (N_44767,N_40014,N_40672);
nor U44768 (N_44768,N_41934,N_40566);
or U44769 (N_44769,N_40563,N_40608);
xnor U44770 (N_44770,N_40969,N_41744);
and U44771 (N_44771,N_40054,N_40681);
or U44772 (N_44772,N_40087,N_40041);
or U44773 (N_44773,N_40131,N_41973);
nor U44774 (N_44774,N_41672,N_40305);
nand U44775 (N_44775,N_40200,N_40712);
nand U44776 (N_44776,N_41406,N_40371);
nor U44777 (N_44777,N_41848,N_40821);
or U44778 (N_44778,N_42132,N_41499);
nor U44779 (N_44779,N_41461,N_40240);
or U44780 (N_44780,N_41640,N_42072);
and U44781 (N_44781,N_42121,N_42034);
xnor U44782 (N_44782,N_40917,N_41431);
or U44783 (N_44783,N_40756,N_42161);
or U44784 (N_44784,N_40512,N_41964);
nand U44785 (N_44785,N_41232,N_41857);
nand U44786 (N_44786,N_41630,N_41178);
xor U44787 (N_44787,N_41574,N_41447);
nor U44788 (N_44788,N_40394,N_41257);
nand U44789 (N_44789,N_40397,N_40897);
and U44790 (N_44790,N_40671,N_41114);
or U44791 (N_44791,N_40446,N_40763);
xor U44792 (N_44792,N_42214,N_42294);
nor U44793 (N_44793,N_41644,N_40157);
nand U44794 (N_44794,N_42049,N_40444);
and U44795 (N_44795,N_41857,N_40600);
and U44796 (N_44796,N_40412,N_40738);
and U44797 (N_44797,N_41347,N_41150);
nor U44798 (N_44798,N_40724,N_41309);
xor U44799 (N_44799,N_40955,N_41872);
nand U44800 (N_44800,N_40515,N_41398);
nor U44801 (N_44801,N_40016,N_42267);
or U44802 (N_44802,N_41325,N_40109);
or U44803 (N_44803,N_41707,N_41781);
or U44804 (N_44804,N_41166,N_42360);
nor U44805 (N_44805,N_41422,N_42326);
and U44806 (N_44806,N_41276,N_41247);
nand U44807 (N_44807,N_40667,N_42207);
or U44808 (N_44808,N_41622,N_40280);
xnor U44809 (N_44809,N_40609,N_41036);
nand U44810 (N_44810,N_40177,N_41299);
nand U44811 (N_44811,N_40837,N_41386);
or U44812 (N_44812,N_41164,N_41627);
nor U44813 (N_44813,N_41367,N_41633);
nor U44814 (N_44814,N_40380,N_40943);
nand U44815 (N_44815,N_41099,N_42017);
and U44816 (N_44816,N_41299,N_40877);
nand U44817 (N_44817,N_41933,N_40459);
nor U44818 (N_44818,N_41136,N_42358);
nand U44819 (N_44819,N_40042,N_40729);
and U44820 (N_44820,N_40954,N_40530);
and U44821 (N_44821,N_40607,N_40020);
or U44822 (N_44822,N_41301,N_41612);
or U44823 (N_44823,N_42470,N_40490);
nor U44824 (N_44824,N_41562,N_40932);
or U44825 (N_44825,N_42134,N_40221);
nand U44826 (N_44826,N_40015,N_40908);
nand U44827 (N_44827,N_40573,N_41333);
and U44828 (N_44828,N_42247,N_42449);
and U44829 (N_44829,N_40671,N_42226);
nand U44830 (N_44830,N_41608,N_41980);
or U44831 (N_44831,N_40172,N_41204);
nor U44832 (N_44832,N_40906,N_40925);
and U44833 (N_44833,N_41225,N_41968);
and U44834 (N_44834,N_40328,N_40064);
or U44835 (N_44835,N_40487,N_42080);
nand U44836 (N_44836,N_42017,N_42157);
and U44837 (N_44837,N_40040,N_40209);
nand U44838 (N_44838,N_40334,N_41651);
or U44839 (N_44839,N_42403,N_41463);
nor U44840 (N_44840,N_41486,N_41501);
nand U44841 (N_44841,N_42489,N_40532);
xor U44842 (N_44842,N_40034,N_42407);
or U44843 (N_44843,N_41332,N_40221);
xor U44844 (N_44844,N_40336,N_41720);
xor U44845 (N_44845,N_42323,N_41177);
or U44846 (N_44846,N_41777,N_41646);
and U44847 (N_44847,N_40879,N_41598);
nor U44848 (N_44848,N_40263,N_40775);
and U44849 (N_44849,N_40288,N_40312);
or U44850 (N_44850,N_42051,N_42477);
nor U44851 (N_44851,N_41714,N_41650);
nand U44852 (N_44852,N_40400,N_40657);
nand U44853 (N_44853,N_41884,N_42092);
or U44854 (N_44854,N_40364,N_40302);
nor U44855 (N_44855,N_40358,N_41561);
xnor U44856 (N_44856,N_42488,N_41999);
or U44857 (N_44857,N_40326,N_41418);
nand U44858 (N_44858,N_40208,N_41400);
nand U44859 (N_44859,N_41888,N_40817);
and U44860 (N_44860,N_42323,N_40566);
xor U44861 (N_44861,N_42486,N_40471);
nor U44862 (N_44862,N_42468,N_40610);
nor U44863 (N_44863,N_42178,N_42077);
and U44864 (N_44864,N_42182,N_41807);
nor U44865 (N_44865,N_42422,N_40232);
and U44866 (N_44866,N_42073,N_40712);
nand U44867 (N_44867,N_41850,N_42332);
xor U44868 (N_44868,N_41485,N_41713);
or U44869 (N_44869,N_40566,N_40513);
nor U44870 (N_44870,N_41629,N_41907);
nor U44871 (N_44871,N_40779,N_42097);
nor U44872 (N_44872,N_41507,N_41932);
nor U44873 (N_44873,N_42000,N_40825);
or U44874 (N_44874,N_40049,N_41405);
nand U44875 (N_44875,N_40929,N_40446);
or U44876 (N_44876,N_42363,N_42108);
nand U44877 (N_44877,N_41978,N_40696);
and U44878 (N_44878,N_41436,N_41259);
or U44879 (N_44879,N_41845,N_41095);
xor U44880 (N_44880,N_40933,N_40666);
nor U44881 (N_44881,N_41163,N_41161);
xor U44882 (N_44882,N_40257,N_41257);
nor U44883 (N_44883,N_42324,N_41378);
and U44884 (N_44884,N_40552,N_41284);
and U44885 (N_44885,N_40715,N_41060);
and U44886 (N_44886,N_42239,N_40317);
nor U44887 (N_44887,N_41887,N_40348);
nand U44888 (N_44888,N_41445,N_40620);
nor U44889 (N_44889,N_41065,N_41648);
nor U44890 (N_44890,N_41485,N_41180);
nand U44891 (N_44891,N_41681,N_40209);
nand U44892 (N_44892,N_40982,N_41386);
nand U44893 (N_44893,N_40133,N_40828);
nand U44894 (N_44894,N_40745,N_42173);
nand U44895 (N_44895,N_41919,N_41292);
or U44896 (N_44896,N_41286,N_40989);
and U44897 (N_44897,N_40287,N_41306);
and U44898 (N_44898,N_40401,N_41467);
or U44899 (N_44899,N_40858,N_41553);
nor U44900 (N_44900,N_40419,N_40656);
and U44901 (N_44901,N_41156,N_40505);
nor U44902 (N_44902,N_42333,N_40949);
and U44903 (N_44903,N_41794,N_40161);
and U44904 (N_44904,N_41409,N_42325);
nor U44905 (N_44905,N_40553,N_41799);
or U44906 (N_44906,N_41018,N_42254);
and U44907 (N_44907,N_40932,N_41184);
nor U44908 (N_44908,N_40195,N_41032);
nor U44909 (N_44909,N_40021,N_41289);
xnor U44910 (N_44910,N_40714,N_42311);
or U44911 (N_44911,N_40545,N_40004);
nor U44912 (N_44912,N_41277,N_40751);
and U44913 (N_44913,N_40327,N_42442);
nand U44914 (N_44914,N_40222,N_40643);
or U44915 (N_44915,N_40369,N_41578);
and U44916 (N_44916,N_40548,N_42395);
nand U44917 (N_44917,N_40710,N_40245);
nand U44918 (N_44918,N_41163,N_41806);
nor U44919 (N_44919,N_41044,N_40950);
nand U44920 (N_44920,N_41195,N_41975);
or U44921 (N_44921,N_40174,N_40623);
and U44922 (N_44922,N_40716,N_40413);
or U44923 (N_44923,N_42019,N_40257);
or U44924 (N_44924,N_41948,N_42107);
nand U44925 (N_44925,N_41833,N_40904);
nand U44926 (N_44926,N_40802,N_41518);
nand U44927 (N_44927,N_40104,N_42259);
and U44928 (N_44928,N_41346,N_40380);
xnor U44929 (N_44929,N_40491,N_40323);
or U44930 (N_44930,N_41136,N_40867);
nor U44931 (N_44931,N_40105,N_40037);
nand U44932 (N_44932,N_40635,N_40583);
and U44933 (N_44933,N_42120,N_40858);
xnor U44934 (N_44934,N_40426,N_40588);
and U44935 (N_44935,N_40586,N_42382);
and U44936 (N_44936,N_41189,N_40706);
nand U44937 (N_44937,N_41106,N_40617);
nor U44938 (N_44938,N_41183,N_40827);
nand U44939 (N_44939,N_42077,N_41139);
or U44940 (N_44940,N_41830,N_40382);
nand U44941 (N_44941,N_40473,N_40136);
nor U44942 (N_44942,N_41325,N_40222);
and U44943 (N_44943,N_41213,N_41115);
nor U44944 (N_44944,N_41519,N_40059);
nor U44945 (N_44945,N_41286,N_40639);
nor U44946 (N_44946,N_40998,N_40626);
nand U44947 (N_44947,N_41556,N_41981);
nand U44948 (N_44948,N_42105,N_41035);
and U44949 (N_44949,N_40977,N_41761);
nor U44950 (N_44950,N_41328,N_41723);
and U44951 (N_44951,N_41331,N_40761);
xnor U44952 (N_44952,N_41027,N_41676);
xor U44953 (N_44953,N_42041,N_40715);
and U44954 (N_44954,N_41607,N_40597);
or U44955 (N_44955,N_40964,N_41751);
nand U44956 (N_44956,N_41840,N_41329);
or U44957 (N_44957,N_40680,N_41170);
nor U44958 (N_44958,N_40026,N_41501);
and U44959 (N_44959,N_42417,N_40281);
xor U44960 (N_44960,N_40702,N_40240);
and U44961 (N_44961,N_40426,N_41554);
or U44962 (N_44962,N_40064,N_40744);
nor U44963 (N_44963,N_41096,N_40459);
nor U44964 (N_44964,N_41849,N_40277);
and U44965 (N_44965,N_41162,N_40147);
nand U44966 (N_44966,N_40433,N_42360);
xnor U44967 (N_44967,N_41370,N_40017);
or U44968 (N_44968,N_42319,N_41990);
and U44969 (N_44969,N_41613,N_42198);
xor U44970 (N_44970,N_42400,N_41878);
nand U44971 (N_44971,N_40002,N_40650);
nor U44972 (N_44972,N_40142,N_40516);
nor U44973 (N_44973,N_42124,N_40595);
and U44974 (N_44974,N_41742,N_42286);
or U44975 (N_44975,N_42461,N_41570);
or U44976 (N_44976,N_41307,N_41609);
or U44977 (N_44977,N_41096,N_40055);
and U44978 (N_44978,N_41146,N_40205);
nand U44979 (N_44979,N_41212,N_41548);
nand U44980 (N_44980,N_40708,N_40256);
or U44981 (N_44981,N_41353,N_42462);
and U44982 (N_44982,N_40639,N_41655);
or U44983 (N_44983,N_42128,N_40801);
nor U44984 (N_44984,N_42441,N_40087);
nand U44985 (N_44985,N_41167,N_42364);
nor U44986 (N_44986,N_41258,N_40198);
nand U44987 (N_44987,N_41610,N_41718);
nand U44988 (N_44988,N_41673,N_41276);
xor U44989 (N_44989,N_40520,N_40158);
or U44990 (N_44990,N_41513,N_42295);
xor U44991 (N_44991,N_41827,N_40106);
nor U44992 (N_44992,N_40512,N_41390);
nor U44993 (N_44993,N_41329,N_40873);
and U44994 (N_44994,N_41886,N_41903);
xor U44995 (N_44995,N_41017,N_41141);
and U44996 (N_44996,N_41131,N_42050);
or U44997 (N_44997,N_41546,N_41978);
nand U44998 (N_44998,N_41875,N_41051);
nor U44999 (N_44999,N_42279,N_42086);
or U45000 (N_45000,N_42864,N_44603);
and U45001 (N_45001,N_43405,N_44743);
or U45002 (N_45002,N_42715,N_43727);
nor U45003 (N_45003,N_43497,N_44087);
and U45004 (N_45004,N_42794,N_44736);
nand U45005 (N_45005,N_43928,N_44651);
xnor U45006 (N_45006,N_44554,N_44486);
nand U45007 (N_45007,N_43155,N_44723);
and U45008 (N_45008,N_44522,N_42703);
or U45009 (N_45009,N_42571,N_44261);
nor U45010 (N_45010,N_44584,N_44403);
and U45011 (N_45011,N_43825,N_43752);
or U45012 (N_45012,N_43474,N_42578);
and U45013 (N_45013,N_44359,N_43258);
or U45014 (N_45014,N_44777,N_43569);
nand U45015 (N_45015,N_43142,N_44582);
nand U45016 (N_45016,N_43080,N_44157);
nand U45017 (N_45017,N_43774,N_42854);
or U45018 (N_45018,N_44558,N_44568);
or U45019 (N_45019,N_44090,N_44181);
nor U45020 (N_45020,N_43366,N_44770);
nand U45021 (N_45021,N_44216,N_43909);
and U45022 (N_45022,N_44659,N_44395);
and U45023 (N_45023,N_43566,N_43183);
xnor U45024 (N_45024,N_42654,N_42754);
nor U45025 (N_45025,N_42580,N_43396);
nor U45026 (N_45026,N_42612,N_44616);
xor U45027 (N_45027,N_44371,N_44705);
or U45028 (N_45028,N_43740,N_44141);
and U45029 (N_45029,N_43586,N_43703);
and U45030 (N_45030,N_43145,N_43284);
or U45031 (N_45031,N_44514,N_43089);
and U45032 (N_45032,N_44009,N_44140);
nor U45033 (N_45033,N_43222,N_44247);
xnor U45034 (N_45034,N_42776,N_43299);
nand U45035 (N_45035,N_42718,N_42641);
and U45036 (N_45036,N_44468,N_43936);
nand U45037 (N_45037,N_43908,N_44585);
or U45038 (N_45038,N_44811,N_42749);
and U45039 (N_45039,N_42515,N_44882);
or U45040 (N_45040,N_43411,N_43522);
nand U45041 (N_45041,N_44117,N_42546);
nand U45042 (N_45042,N_43626,N_44290);
and U45043 (N_45043,N_42604,N_43757);
nand U45044 (N_45044,N_44260,N_43349);
nand U45045 (N_45045,N_44829,N_44146);
nand U45046 (N_45046,N_43961,N_44100);
xnor U45047 (N_45047,N_42652,N_43898);
or U45048 (N_45048,N_44452,N_44861);
nand U45049 (N_45049,N_43565,N_42780);
nand U45050 (N_45050,N_43027,N_44085);
nand U45051 (N_45051,N_44654,N_43718);
xnor U45052 (N_45052,N_44230,N_44111);
xnor U45053 (N_45053,N_43776,N_43841);
nand U45054 (N_45054,N_42885,N_44792);
or U45055 (N_45055,N_44043,N_44560);
xnor U45056 (N_45056,N_44712,N_42672);
nor U45057 (N_45057,N_44674,N_43937);
nand U45058 (N_45058,N_42777,N_43802);
nor U45059 (N_45059,N_44277,N_44800);
and U45060 (N_45060,N_43028,N_42969);
and U45061 (N_45061,N_43094,N_43164);
nor U45062 (N_45062,N_43882,N_43944);
xnor U45063 (N_45063,N_43662,N_44130);
nor U45064 (N_45064,N_42629,N_42511);
nor U45065 (N_45065,N_42665,N_44416);
and U45066 (N_45066,N_43001,N_43714);
xnor U45067 (N_45067,N_43949,N_44205);
and U45068 (N_45068,N_44610,N_43095);
or U45069 (N_45069,N_43933,N_44602);
xnor U45070 (N_45070,N_43584,N_42706);
xor U45071 (N_45071,N_43191,N_44605);
or U45072 (N_45072,N_43036,N_43416);
nand U45073 (N_45073,N_42688,N_42630);
and U45074 (N_45074,N_44653,N_42634);
nor U45075 (N_45075,N_44725,N_42889);
or U45076 (N_45076,N_44940,N_43197);
nand U45077 (N_45077,N_43535,N_43395);
nand U45078 (N_45078,N_42947,N_44912);
nor U45079 (N_45079,N_43336,N_42877);
nor U45080 (N_45080,N_42822,N_43959);
nor U45081 (N_45081,N_43055,N_42748);
and U45082 (N_45082,N_43518,N_42845);
or U45083 (N_45083,N_42853,N_42626);
nor U45084 (N_45084,N_43704,N_44913);
nand U45085 (N_45085,N_43962,N_44187);
xnor U45086 (N_45086,N_42548,N_44017);
xnor U45087 (N_45087,N_44583,N_43005);
and U45088 (N_45088,N_43845,N_43054);
xor U45089 (N_45089,N_43391,N_43086);
or U45090 (N_45090,N_44967,N_42951);
and U45091 (N_45091,N_44224,N_43019);
nor U45092 (N_45092,N_43126,N_44256);
and U45093 (N_45093,N_42576,N_43374);
xnor U45094 (N_45094,N_42646,N_43710);
and U45095 (N_45095,N_44590,N_44986);
or U45096 (N_45096,N_44243,N_42823);
or U45097 (N_45097,N_43975,N_43957);
and U45098 (N_45098,N_44868,N_42613);
or U45099 (N_45099,N_43250,N_43449);
nand U45100 (N_45100,N_43220,N_44565);
and U45101 (N_45101,N_43941,N_43890);
nand U45102 (N_45102,N_42670,N_44380);
nand U45103 (N_45103,N_44000,N_44744);
xor U45104 (N_45104,N_42819,N_42653);
and U45105 (N_45105,N_43448,N_42559);
or U45106 (N_45106,N_44776,N_42940);
nor U45107 (N_45107,N_42751,N_43316);
nor U45108 (N_45108,N_43268,N_43643);
nor U45109 (N_45109,N_44356,N_42659);
nor U45110 (N_45110,N_43397,N_42684);
nand U45111 (N_45111,N_43021,N_44142);
or U45112 (N_45112,N_44608,N_43093);
and U45113 (N_45113,N_42868,N_44992);
and U45114 (N_45114,N_44709,N_44351);
or U45115 (N_45115,N_44499,N_43982);
nand U45116 (N_45116,N_44828,N_44896);
and U45117 (N_45117,N_43153,N_44738);
and U45118 (N_45118,N_42784,N_42887);
or U45119 (N_45119,N_44488,N_43066);
nand U45120 (N_45120,N_42895,N_43043);
or U45121 (N_45121,N_44687,N_43323);
and U45122 (N_45122,N_43230,N_43057);
nand U45123 (N_45123,N_42508,N_42771);
xor U45124 (N_45124,N_42835,N_42957);
and U45125 (N_45125,N_43932,N_43637);
xnor U45126 (N_45126,N_42556,N_42863);
or U45127 (N_45127,N_42640,N_43308);
xor U45128 (N_45128,N_44262,N_42725);
nor U45129 (N_45129,N_44575,N_43798);
and U45130 (N_45130,N_44990,N_44690);
nand U45131 (N_45131,N_44020,N_44268);
nand U45132 (N_45132,N_43623,N_42584);
nor U45133 (N_45133,N_42890,N_43708);
nor U45134 (N_45134,N_44885,N_44657);
nor U45135 (N_45135,N_43294,N_44436);
or U45136 (N_45136,N_42888,N_43223);
nand U45137 (N_45137,N_44075,N_44814);
or U45138 (N_45138,N_42724,N_43796);
xnor U45139 (N_45139,N_43355,N_44822);
or U45140 (N_45140,N_43495,N_42903);
or U45141 (N_45141,N_43510,N_43138);
nand U45142 (N_45142,N_44379,N_43219);
nand U45143 (N_45143,N_42941,N_43891);
nand U45144 (N_45144,N_43827,N_42768);
nor U45145 (N_45145,N_42900,N_43163);
xnor U45146 (N_45146,N_43029,N_44255);
and U45147 (N_45147,N_43666,N_43523);
nand U45148 (N_45148,N_43195,N_42856);
xnor U45149 (N_45149,N_42981,N_43428);
xor U45150 (N_45150,N_44866,N_44597);
and U45151 (N_45151,N_42542,N_44365);
or U45152 (N_45152,N_43635,N_43143);
nand U45153 (N_45153,N_43473,N_44018);
nor U45154 (N_45154,N_44241,N_42717);
nand U45155 (N_45155,N_43023,N_44056);
and U45156 (N_45156,N_44715,N_44831);
nor U45157 (N_45157,N_43877,N_43177);
or U45158 (N_45158,N_44774,N_43152);
nor U45159 (N_45159,N_42944,N_42553);
xnor U45160 (N_45160,N_44340,N_43399);
and U45161 (N_45161,N_43820,N_44294);
or U45162 (N_45162,N_43998,N_42605);
nand U45163 (N_45163,N_44012,N_44806);
and U45164 (N_45164,N_42747,N_44055);
nand U45165 (N_45165,N_44665,N_43656);
nor U45166 (N_45166,N_42860,N_44720);
xnor U45167 (N_45167,N_44646,N_44830);
or U45168 (N_45168,N_44498,N_44617);
and U45169 (N_45169,N_43446,N_43059);
xnor U45170 (N_45170,N_43070,N_42552);
nand U45171 (N_45171,N_44683,N_44004);
and U45172 (N_45172,N_44700,N_43667);
nor U45173 (N_45173,N_44005,N_44221);
or U45174 (N_45174,N_43762,N_43506);
nor U45175 (N_45175,N_43859,N_43289);
xor U45176 (N_45176,N_44483,N_44136);
nand U45177 (N_45177,N_44195,N_43967);
or U45178 (N_45178,N_42818,N_43443);
nor U45179 (N_45179,N_42591,N_44540);
nor U45180 (N_45180,N_43319,N_43713);
or U45181 (N_45181,N_44508,N_44190);
nand U45182 (N_45182,N_43108,N_43300);
nor U45183 (N_45183,N_43646,N_44670);
nor U45184 (N_45184,N_44098,N_44234);
nand U45185 (N_45185,N_44640,N_43022);
or U45186 (N_45186,N_43769,N_43707);
nand U45187 (N_45187,N_43793,N_42529);
nand U45188 (N_45188,N_44444,N_44595);
nand U45189 (N_45189,N_44559,N_43689);
xnor U45190 (N_45190,N_43462,N_42833);
or U45191 (N_45191,N_42943,N_44673);
nand U45192 (N_45192,N_43767,N_42600);
xor U45193 (N_45193,N_43888,N_43334);
nand U45194 (N_45194,N_44629,N_44914);
and U45195 (N_45195,N_44567,N_44675);
or U45196 (N_45196,N_44390,N_42946);
or U45197 (N_45197,N_44387,N_42958);
nor U45198 (N_45198,N_44406,N_43088);
xnor U45199 (N_45199,N_44496,N_42998);
or U45200 (N_45200,N_44834,N_43159);
nand U45201 (N_45201,N_43178,N_44661);
and U45202 (N_45202,N_44202,N_42657);
xor U45203 (N_45203,N_43722,N_43843);
and U45204 (N_45204,N_43678,N_44908);
nor U45205 (N_45205,N_42816,N_44794);
and U45206 (N_45206,N_44721,N_44063);
nor U45207 (N_45207,N_44816,N_44346);
nand U45208 (N_45208,N_43715,N_43842);
nand U45209 (N_45209,N_44501,N_44399);
xor U45210 (N_45210,N_43465,N_44698);
and U45211 (N_45211,N_44276,N_43150);
nor U45212 (N_45212,N_44556,N_43673);
and U45213 (N_45213,N_43161,N_44441);
xor U45214 (N_45214,N_42809,N_43546);
or U45215 (N_45215,N_43075,N_44702);
or U45216 (N_45216,N_44482,N_42583);
or U45217 (N_45217,N_44947,N_44252);
or U45218 (N_45218,N_43551,N_44790);
xnor U45219 (N_45219,N_44587,N_43595);
nand U45220 (N_45220,N_42792,N_44696);
xor U45221 (N_45221,N_42512,N_44102);
nand U45222 (N_45222,N_44311,N_42988);
nor U45223 (N_45223,N_43306,N_43880);
and U45224 (N_45224,N_43658,N_42628);
nor U45225 (N_45225,N_43291,N_44065);
nand U45226 (N_45226,N_43167,N_44415);
xor U45227 (N_45227,N_42732,N_43240);
nand U45228 (N_45228,N_44642,N_44286);
nor U45229 (N_45229,N_44958,N_42638);
and U45230 (N_45230,N_44625,N_43834);
or U45231 (N_45231,N_43298,N_44842);
or U45232 (N_45232,N_43751,N_42907);
nor U45233 (N_45233,N_44166,N_42625);
or U45234 (N_45234,N_43994,N_42610);
or U45235 (N_45235,N_43725,N_43562);
and U45236 (N_45236,N_43854,N_44729);
or U45237 (N_45237,N_44748,N_42622);
nor U45238 (N_45238,N_43192,N_42567);
nand U45239 (N_45239,N_44549,N_42972);
or U45240 (N_45240,N_44758,N_44859);
or U45241 (N_45241,N_44999,N_44572);
xor U45242 (N_45242,N_43753,N_44910);
or U45243 (N_45243,N_43954,N_43369);
and U45244 (N_45244,N_42783,N_43050);
nand U45245 (N_45245,N_42983,N_44152);
and U45246 (N_45246,N_43441,N_44521);
nand U45247 (N_45247,N_43871,N_43971);
xor U45248 (N_45248,N_43594,N_42535);
or U45249 (N_45249,N_43985,N_42793);
and U45250 (N_45250,N_42539,N_42627);
or U45251 (N_45251,N_43322,N_43091);
or U45252 (N_45252,N_44203,N_44228);
nor U45253 (N_45253,N_43368,N_44662);
nand U45254 (N_45254,N_42708,N_42924);
xnor U45255 (N_45255,N_44068,N_44079);
xor U45256 (N_45256,N_43181,N_44529);
and U45257 (N_45257,N_43046,N_44779);
nor U45258 (N_45258,N_44363,N_44123);
nand U45259 (N_45259,N_44167,N_43385);
nand U45260 (N_45260,N_42847,N_43824);
nor U45261 (N_45261,N_43119,N_43477);
and U45262 (N_45262,N_43099,N_43362);
nor U45263 (N_45263,N_44844,N_43568);
nand U45264 (N_45264,N_43668,N_44235);
xnor U45265 (N_45265,N_43582,N_43922);
nand U45266 (N_45266,N_43720,N_44513);
nor U45267 (N_45267,N_42927,N_44706);
nor U45268 (N_45268,N_43453,N_44948);
and U45269 (N_45269,N_44158,N_43672);
and U45270 (N_45270,N_42716,N_43581);
xor U45271 (N_45271,N_43002,N_43614);
or U45272 (N_45272,N_42786,N_44019);
and U45273 (N_45273,N_42753,N_44414);
xnor U45274 (N_45274,N_44377,N_42647);
xor U45275 (N_45275,N_43205,N_44472);
nand U45276 (N_45276,N_43602,N_44088);
and U45277 (N_45277,N_44761,N_44592);
nand U45278 (N_45278,N_42525,N_44516);
or U45279 (N_45279,N_42701,N_44393);
nand U45280 (N_45280,N_42597,N_42541);
nor U45281 (N_45281,N_43135,N_44231);
or U45282 (N_45282,N_43700,N_44957);
nor U45283 (N_45283,N_43400,N_44176);
and U45284 (N_45284,N_44327,N_44765);
or U45285 (N_45285,N_43848,N_42633);
and U45286 (N_45286,N_42516,N_42566);
nor U45287 (N_45287,N_43123,N_44718);
xor U45288 (N_45288,N_43408,N_42862);
or U45289 (N_45289,N_43124,N_43359);
nor U45290 (N_45290,N_44400,N_42668);
xnor U45291 (N_45291,N_44434,N_44192);
or U45292 (N_45292,N_42565,N_42931);
nor U45293 (N_45293,N_44506,N_42857);
and U45294 (N_45294,N_42956,N_42741);
and U45295 (N_45295,N_43206,N_43572);
xnor U45296 (N_45296,N_43243,N_44153);
nand U45297 (N_45297,N_43198,N_43990);
nand U45298 (N_45298,N_42526,N_43147);
nor U45299 (N_45299,N_43730,N_43784);
nand U45300 (N_45300,N_43338,N_43828);
and U45301 (N_45301,N_43530,N_44755);
nand U45302 (N_45302,N_44562,N_43690);
and U45303 (N_45303,N_43879,N_44070);
or U45304 (N_45304,N_43991,N_44366);
or U45305 (N_45305,N_42978,N_44312);
nor U45306 (N_45306,N_42905,N_43134);
and U45307 (N_45307,N_44746,N_44747);
and U45308 (N_45308,N_44808,N_43184);
and U45309 (N_45309,N_42500,N_42593);
nand U45310 (N_45310,N_43232,N_42984);
nand U45311 (N_45311,N_44298,N_44325);
or U45312 (N_45312,N_43846,N_43017);
xnor U45313 (N_45313,N_44451,N_44465);
xor U45314 (N_45314,N_44175,N_43813);
and U45315 (N_45315,N_44108,N_43534);
nor U45316 (N_45316,N_43255,N_44394);
xor U45317 (N_45317,N_44392,N_44784);
nor U45318 (N_45318,N_42585,N_43578);
nand U45319 (N_45319,N_43320,N_42543);
nand U45320 (N_45320,N_44676,N_43978);
xor U45321 (N_45321,N_42966,N_43897);
xnor U45322 (N_45322,N_43615,N_43622);
or U45323 (N_45323,N_44539,N_43218);
nand U45324 (N_45324,N_44291,N_44813);
nor U45325 (N_45325,N_43613,N_43287);
or U45326 (N_45326,N_43025,N_43943);
or U45327 (N_45327,N_44484,N_43296);
and U45328 (N_45328,N_42694,N_43188);
nand U45329 (N_45329,N_43548,N_43141);
and U45330 (N_45330,N_44161,N_42873);
and U45331 (N_45331,N_43940,N_43588);
or U45332 (N_45332,N_43274,N_43372);
nand U45333 (N_45333,N_44273,N_43440);
or U45334 (N_45334,N_44648,N_42642);
nor U45335 (N_45335,N_43144,N_43968);
or U45336 (N_45336,N_44112,N_43857);
and U45337 (N_45337,N_43122,N_44571);
and U45338 (N_45338,N_42899,N_43743);
or U45339 (N_45339,N_44727,N_43194);
nand U45340 (N_45340,N_44898,N_43467);
nand U45341 (N_45341,N_43939,N_44168);
or U45342 (N_45342,N_44271,N_44737);
xnor U45343 (N_45343,N_44149,N_42913);
nor U45344 (N_45344,N_42901,N_43726);
or U45345 (N_45345,N_42648,N_44893);
nor U45346 (N_45346,N_43060,N_42733);
or U45347 (N_45347,N_44427,N_44494);
nor U45348 (N_45348,N_43063,N_43663);
and U45349 (N_45349,N_43648,N_44589);
and U45350 (N_45350,N_43699,N_42573);
nor U45351 (N_45351,N_42719,N_43176);
and U45352 (N_45352,N_44170,N_43868);
nand U45353 (N_45353,N_44352,N_44760);
nand U45354 (N_45354,N_43585,N_43674);
or U45355 (N_45355,N_44109,N_44083);
and U45356 (N_45356,N_43761,N_43992);
xnor U45357 (N_45357,N_44686,N_44825);
and U45358 (N_45358,N_43442,N_44062);
and U45359 (N_45359,N_43280,N_44713);
or U45360 (N_45360,N_44218,N_44671);
nor U45361 (N_45361,N_42547,N_43759);
nand U45362 (N_45362,N_44292,N_42789);
nand U45363 (N_45363,N_43945,N_43335);
nor U45364 (N_45364,N_44970,N_42538);
nand U45365 (N_45365,N_44342,N_43052);
or U45366 (N_45366,N_42821,N_44911);
or U45367 (N_45367,N_44525,N_44080);
nand U45368 (N_45368,N_44734,N_43422);
or U45369 (N_45369,N_43004,N_44222);
or U45370 (N_45370,N_43263,N_43576);
xnor U45371 (N_45371,N_43680,N_44552);
or U45372 (N_45372,N_43779,N_44875);
nand U45373 (N_45373,N_42698,N_42743);
and U45374 (N_45374,N_42985,N_43007);
or U45375 (N_45375,N_43180,N_44201);
nor U45376 (N_45376,N_43640,N_43378);
or U45377 (N_45377,N_43641,N_44133);
or U45378 (N_45378,N_43914,N_43012);
and U45379 (N_45379,N_44778,N_43498);
nand U45380 (N_45380,N_44470,N_43929);
and U45381 (N_45381,N_44909,N_44753);
nor U45382 (N_45382,N_43034,N_43812);
xnor U45383 (N_45383,N_43421,N_44780);
and U45384 (N_45384,N_44066,N_44954);
xor U45385 (N_45385,N_44148,N_44404);
or U45386 (N_45386,N_43304,N_44869);
nor U45387 (N_45387,N_42880,N_44707);
nor U45388 (N_45388,N_44375,N_44313);
nand U45389 (N_45389,N_42611,N_44189);
or U45390 (N_45390,N_43839,N_44607);
and U45391 (N_45391,N_44439,N_43275);
nand U45392 (N_45392,N_43042,N_44071);
and U45393 (N_45393,N_43049,N_44714);
xnor U45394 (N_45394,N_43324,N_44489);
nor U45395 (N_45395,N_43679,N_42699);
nand U45396 (N_45396,N_42620,N_43491);
or U45397 (N_45397,N_44726,N_42680);
nand U45398 (N_45398,N_42902,N_44033);
xor U45399 (N_45399,N_43077,N_43292);
nand U45400 (N_45400,N_42677,N_44469);
or U45401 (N_45401,N_43013,N_44047);
and U45402 (N_45402,N_42769,N_44599);
or U45403 (N_45403,N_42918,N_42832);
nor U45404 (N_45404,N_43329,N_44561);
or U45405 (N_45405,N_43437,N_42679);
xor U45406 (N_45406,N_44953,N_44965);
or U45407 (N_45407,N_42910,N_44384);
and U45408 (N_45408,N_42945,N_44233);
nor U45409 (N_45409,N_43809,N_42550);
and U45410 (N_45410,N_42690,N_44401);
xor U45411 (N_45411,N_44265,N_43283);
and U45412 (N_45412,N_43557,N_42937);
and U45413 (N_45413,N_43352,N_43987);
or U45414 (N_45414,N_44892,N_44807);
and U45415 (N_45415,N_42727,N_42616);
or U45416 (N_45416,N_43763,N_44636);
and U45417 (N_45417,N_42992,N_44178);
and U45418 (N_45418,N_44034,N_44897);
nor U45419 (N_45419,N_43107,N_43958);
and U45420 (N_45420,N_43866,N_43082);
and U45421 (N_45421,N_44338,N_43429);
nor U45422 (N_45422,N_42844,N_43731);
nand U45423 (N_45423,N_44695,N_44775);
xnor U45424 (N_45424,N_43133,N_43424);
or U45425 (N_45425,N_44455,N_43278);
xnor U45426 (N_45426,N_43811,N_44269);
nor U45427 (N_45427,N_43905,N_44889);
and U45428 (N_45428,N_44369,N_42707);
nor U45429 (N_45429,N_44138,N_44491);
xor U45430 (N_45430,N_43310,N_44691);
and U45431 (N_45431,N_44105,N_43203);
xor U45432 (N_45432,N_43386,N_44283);
nand U45433 (N_45433,N_44275,N_43536);
xor U45434 (N_45434,N_43494,N_43047);
and U45435 (N_45435,N_42658,N_42663);
nand U45436 (N_45436,N_43942,N_44735);
xnor U45437 (N_45437,N_43367,N_44282);
nand U45438 (N_45438,N_44998,N_43175);
nor U45439 (N_45439,N_43733,N_43048);
nor U45440 (N_45440,N_43327,N_43382);
nor U45441 (N_45441,N_43317,N_43247);
and U45442 (N_45442,N_42702,N_42935);
nor U45443 (N_45443,N_44523,N_42586);
and U45444 (N_45444,N_42894,N_44824);
or U45445 (N_45445,N_42820,N_43636);
and U45446 (N_45446,N_43960,N_44310);
or U45447 (N_45447,N_44272,N_43709);
nand U45448 (N_45448,N_44076,N_43402);
or U45449 (N_45449,N_44348,N_43267);
nand U45450 (N_45450,N_43480,N_43711);
and U45451 (N_45451,N_44383,N_42848);
nand U45452 (N_45452,N_42623,N_43204);
nand U45453 (N_45453,N_43625,N_44915);
or U45454 (N_45454,N_43930,N_43748);
and U45455 (N_45455,N_42569,N_43865);
and U45456 (N_45456,N_44267,N_44846);
nand U45457 (N_45457,N_44564,N_43547);
or U45458 (N_45458,N_44129,N_44699);
nand U45459 (N_45459,N_44517,N_42834);
and U45460 (N_45460,N_44881,N_44357);
or U45461 (N_45461,N_42510,N_44128);
nand U45462 (N_45462,N_43031,N_43794);
or U45463 (N_45463,N_43861,N_43728);
and U45464 (N_45464,N_43116,N_44320);
and U45465 (N_45465,N_42841,N_42919);
xor U45466 (N_45466,N_43904,N_44308);
nand U45467 (N_45467,N_44923,N_43103);
or U45468 (N_45468,N_44782,N_43593);
xnor U45469 (N_45469,N_42851,N_43035);
or U45470 (N_45470,N_43977,N_44305);
nor U45471 (N_45471,N_42993,N_43910);
and U45472 (N_45472,N_43719,N_42872);
and U45473 (N_45473,N_44028,N_44238);
and U45474 (N_45474,N_43886,N_42979);
and U45475 (N_45475,N_43307,N_43469);
nand U45476 (N_45476,N_44171,N_42831);
xnor U45477 (N_45477,N_43948,N_44025);
and U45478 (N_45478,N_43862,N_43375);
nand U45479 (N_45479,N_43340,N_43540);
or U45480 (N_45480,N_43348,N_43887);
or U45481 (N_45481,N_44754,N_43339);
nor U45482 (N_45482,N_43496,N_43040);
nor U45483 (N_45483,N_44650,N_42869);
nor U45484 (N_45484,N_44941,N_43729);
nand U45485 (N_45485,N_44535,N_43182);
or U45486 (N_45486,N_43587,N_42926);
or U45487 (N_45487,N_43100,N_44643);
or U45488 (N_45488,N_43724,N_42737);
nand U45489 (N_45489,N_44300,N_42810);
nor U45490 (N_45490,N_43235,N_43236);
nor U45491 (N_45491,N_43744,N_44639);
or U45492 (N_45492,N_44096,N_42865);
and U45493 (N_45493,N_44973,N_42660);
and U45494 (N_45494,N_44001,N_44220);
nor U45495 (N_45495,N_44314,N_44658);
or U45496 (N_45496,N_43599,N_42897);
xor U45497 (N_45497,N_44955,N_42893);
nand U45498 (N_45498,N_43445,N_44835);
nand U45499 (N_45499,N_42656,N_43434);
nor U45500 (N_45500,N_44156,N_44126);
and U45501 (N_45501,N_42922,N_44857);
or U45502 (N_45502,N_42961,N_43325);
or U45503 (N_45503,N_44936,N_43808);
or U45504 (N_45504,N_44788,N_42691);
or U45505 (N_45505,N_44870,N_43537);
or U45506 (N_45506,N_44209,N_43528);
or U45507 (N_45507,N_43911,N_44544);
nand U45508 (N_45508,N_43800,N_44173);
or U45509 (N_45509,N_44015,N_43778);
nand U45510 (N_45510,N_42619,N_42728);
xor U45511 (N_45511,N_44550,N_42624);
nor U45512 (N_45512,N_43433,N_43475);
and U45513 (N_45513,N_44939,N_43755);
xor U45514 (N_45514,N_44789,N_42858);
nor U45515 (N_45515,N_44474,N_43447);
xnor U45516 (N_45516,N_42838,N_43190);
and U45517 (N_45517,N_43764,N_43513);
nand U45518 (N_45518,N_44002,N_44880);
xnor U45519 (N_45519,N_43463,N_42962);
nor U45520 (N_45520,N_44854,N_42963);
or U45521 (N_45521,N_43377,N_43716);
or U45522 (N_45522,N_43903,N_43997);
xnor U45523 (N_45523,N_43281,N_42722);
nor U45524 (N_45524,N_43417,N_44449);
nand U45525 (N_45525,N_44988,N_42799);
nor U45526 (N_45526,N_42773,N_44497);
or U45527 (N_45527,N_42517,N_42763);
and U45528 (N_45528,N_43478,N_44211);
and U45529 (N_45529,N_44278,N_43130);
and U45530 (N_45530,N_44966,N_44032);
nor U45531 (N_45531,N_43590,N_44042);
nor U45532 (N_45532,N_44938,N_44791);
nor U45533 (N_45533,N_44891,N_42636);
or U45534 (N_45534,N_43758,N_44219);
xnor U45535 (N_45535,N_43835,N_44551);
xnor U45536 (N_45536,N_43045,N_43693);
nor U45537 (N_45537,N_42867,N_44989);
and U45538 (N_45538,N_42955,N_43900);
and U45539 (N_45539,N_44364,N_44722);
nand U45540 (N_45540,N_43356,N_44345);
or U45541 (N_45541,N_44114,N_43418);
nand U45542 (N_45542,N_44263,N_44959);
and U45543 (N_45543,N_43989,N_44391);
nand U45544 (N_45544,N_42686,N_43030);
and U45545 (N_45545,N_44456,N_44266);
nand U45546 (N_45546,N_44459,N_43394);
and U45547 (N_45547,N_43330,N_42995);
and U45548 (N_45548,N_44037,N_44509);
xor U45549 (N_45549,N_43033,N_42839);
nand U45550 (N_45550,N_44805,N_43723);
or U45551 (N_45551,N_43016,N_42923);
nor U45552 (N_45552,N_43311,N_43884);
nor U45553 (N_45553,N_43605,N_44185);
nor U45554 (N_45554,N_43869,N_44446);
or U45555 (N_45555,N_42681,N_43951);
or U45556 (N_45556,N_43739,N_44058);
nor U45557 (N_45557,N_44604,N_42536);
nand U45558 (N_45558,N_43026,N_42721);
nor U45559 (N_45559,N_43675,N_44903);
nor U45560 (N_45560,N_42667,N_42644);
or U45561 (N_45561,N_43913,N_42965);
or U45562 (N_45562,N_43639,N_44476);
and U45563 (N_45563,N_44095,N_43526);
and U45564 (N_45564,N_44331,N_43878);
nor U45565 (N_45565,N_44878,N_43132);
nand U45566 (N_45566,N_44409,N_44750);
and U45567 (N_45567,N_42800,N_44431);
and U45568 (N_45568,N_44317,N_43101);
or U45569 (N_45569,N_42574,N_42971);
nand U45570 (N_45570,N_43570,N_44086);
and U45571 (N_45571,N_42795,N_44163);
nor U45572 (N_45572,N_43006,N_44930);
nand U45573 (N_45573,N_44628,N_43836);
nor U45574 (N_45574,N_44995,N_43020);
nand U45575 (N_45575,N_44315,N_43251);
and U45576 (N_45576,N_42861,N_43483);
and U45577 (N_45577,N_43917,N_44442);
or U45578 (N_45578,N_44016,N_44905);
xor U45579 (N_45579,N_44570,N_42996);
nor U45580 (N_45580,N_43170,N_43018);
nand U45581 (N_45581,N_44385,N_42932);
nor U45582 (N_45582,N_43269,N_44106);
xor U45583 (N_45583,N_43695,N_43702);
or U45584 (N_45584,N_44024,N_43331);
nor U45585 (N_45585,N_44011,N_44084);
nor U45586 (N_45586,N_42523,N_43476);
and U45587 (N_45587,N_43501,N_42537);
xor U45588 (N_45588,N_43305,N_42598);
nor U45589 (N_45589,N_44367,N_43488);
nand U45590 (N_45590,N_44478,N_43521);
nor U45591 (N_45591,N_42987,N_44901);
and U45592 (N_45592,N_43895,N_42884);
or U45593 (N_45593,N_43371,N_44057);
or U45594 (N_45594,N_42712,N_43136);
or U45595 (N_45595,N_44429,N_44258);
and U45596 (N_45596,N_42524,N_43817);
or U45597 (N_45597,N_43241,N_43067);
and U45598 (N_45598,N_43295,N_42912);
or U45599 (N_45599,N_44902,N_43683);
xnor U45600 (N_45600,N_44081,N_43092);
nand U45601 (N_45601,N_43039,N_44150);
nand U45602 (N_45602,N_44040,N_43775);
nor U45603 (N_45603,N_44165,N_44091);
or U45604 (N_45604,N_43983,N_44799);
nand U45605 (N_45605,N_44143,N_43790);
and U45606 (N_45606,N_43076,N_43254);
nor U45607 (N_45607,N_43343,N_44531);
or U45608 (N_45608,N_43062,N_43872);
and U45609 (N_45609,N_43544,N_44511);
nand U45610 (N_45610,N_43773,N_44756);
xor U45611 (N_45611,N_42505,N_43127);
nor U45612 (N_45612,N_43406,N_43068);
nand U45613 (N_45613,N_44871,N_43456);
nor U45614 (N_45614,N_44144,N_44543);
or U45615 (N_45615,N_43246,N_44664);
or U45616 (N_45616,N_43981,N_42601);
and U45617 (N_45617,N_43550,N_44681);
xnor U45618 (N_45618,N_44981,N_43363);
or U45619 (N_45619,N_44137,N_44010);
or U45620 (N_45620,N_44297,N_44411);
nand U45621 (N_45621,N_44766,N_43517);
or U45622 (N_45622,N_42790,N_43229);
nand U45623 (N_45623,N_42596,N_43721);
or U45624 (N_45624,N_44285,N_44199);
xnor U45625 (N_45625,N_43651,N_43131);
nand U45626 (N_45626,N_44581,N_42632);
nor U45627 (N_45627,N_42886,N_42916);
and U45628 (N_45628,N_43357,N_43174);
nor U45629 (N_45629,N_43392,N_42999);
and U45630 (N_45630,N_43996,N_43556);
or U45631 (N_45631,N_42726,N_43380);
or U45632 (N_45632,N_44576,N_43571);
nor U45633 (N_45633,N_44733,N_43361);
xnor U45634 (N_45634,N_44249,N_44433);
nor U45635 (N_45635,N_42731,N_44860);
and U45636 (N_45636,N_43479,N_43789);
and U45637 (N_45637,N_43925,N_43780);
nor U45638 (N_45638,N_44703,N_42513);
or U45639 (N_45639,N_43657,N_44886);
and U45640 (N_45640,N_44588,N_44716);
nand U45641 (N_45641,N_44669,N_42609);
and U45642 (N_45642,N_43332,N_43965);
xor U45643 (N_45643,N_43976,N_43791);
nor U45644 (N_45644,N_44652,N_44927);
or U45645 (N_45645,N_44280,N_42815);
and U45646 (N_45646,N_42520,N_44630);
and U45647 (N_45647,N_44206,N_42976);
nand U45648 (N_45648,N_44067,N_44026);
and U45649 (N_45649,N_44410,N_43745);
nor U45650 (N_45650,N_42817,N_43677);
or U45651 (N_45651,N_42977,N_43083);
nor U45652 (N_45652,N_44984,N_44350);
nor U45653 (N_45653,N_43567,N_42693);
and U45654 (N_45654,N_44624,N_44319);
nor U45655 (N_45655,N_43297,N_44739);
or U45656 (N_45656,N_44174,N_43829);
and U45657 (N_45657,N_43074,N_43208);
xor U45658 (N_45658,N_44694,N_43113);
and U45659 (N_45659,N_44388,N_43098);
xor U45660 (N_45660,N_44685,N_42791);
nand U45661 (N_45661,N_42934,N_42871);
nand U45662 (N_45662,N_44339,N_44993);
or U45663 (N_45663,N_42645,N_42615);
nand U45664 (N_45664,N_42592,N_42855);
and U45665 (N_45665,N_42814,N_44463);
nor U45666 (N_45666,N_44728,N_43381);
nor U45667 (N_45667,N_44500,N_44477);
or U45668 (N_45668,N_44492,N_43221);
xnor U45669 (N_45669,N_43064,N_43600);
nor U45670 (N_45670,N_43383,N_44125);
or U45671 (N_45671,N_43260,N_43096);
and U45672 (N_45672,N_42949,N_44917);
and U45673 (N_45673,N_42678,N_42802);
or U45674 (N_45674,N_44611,N_44925);
xnor U45675 (N_45675,N_43239,N_43009);
and U45676 (N_45676,N_44536,N_43788);
or U45677 (N_45677,N_42651,N_44719);
nor U45678 (N_45678,N_44935,N_44963);
nand U45679 (N_45679,N_42558,N_44326);
or U45680 (N_45680,N_43634,N_44863);
nor U45681 (N_45681,N_42757,N_42942);
nor U45682 (N_45682,N_44212,N_44155);
and U45683 (N_45683,N_44933,N_43186);
and U45684 (N_45684,N_44647,N_43885);
nand U45685 (N_45685,N_44596,N_44334);
nor U45686 (N_45686,N_43337,N_42772);
nor U45687 (N_45687,N_43867,N_44888);
nor U45688 (N_45688,N_44299,N_42738);
or U45689 (N_45689,N_44372,N_42602);
and U45690 (N_45690,N_44270,N_43815);
nand U45691 (N_45691,N_43468,N_43603);
and U45692 (N_45692,N_43831,N_43655);
or U45693 (N_45693,N_43915,N_44856);
nor U45694 (N_45694,N_43781,N_42696);
or U45695 (N_45695,N_44145,N_44742);
nand U45696 (N_45696,N_42991,N_43552);
nor U45697 (N_45697,N_43771,N_43919);
nand U45698 (N_45698,N_44120,N_42806);
nor U45699 (N_45699,N_44974,N_43249);
and U45700 (N_45700,N_43426,N_44069);
nor U45701 (N_45701,N_44934,N_43664);
nor U45702 (N_45702,N_43489,N_43554);
and U45703 (N_45703,N_44099,N_42579);
or U45704 (N_45704,N_44680,N_43799);
nand U45705 (N_45705,N_43169,N_43492);
nand U45706 (N_45706,N_44621,N_44147);
and U45707 (N_45707,N_42859,N_43532);
and U45708 (N_45708,N_43787,N_43376);
nand U45709 (N_45709,N_43973,N_44773);
nor U45710 (N_45710,N_43003,N_44526);
nand U45711 (N_45711,N_43087,N_43698);
xor U45712 (N_45712,N_42788,N_44920);
or U45713 (N_45713,N_42840,N_42582);
or U45714 (N_45714,N_44578,N_43312);
or U45715 (N_45715,N_42866,N_44107);
and U45716 (N_45716,N_43404,N_42798);
or U45717 (N_45717,N_43580,N_42563);
or U45718 (N_45718,N_43896,N_43644);
nor U45719 (N_45719,N_44772,N_44039);
and U45720 (N_45720,N_44852,N_43899);
nor U45721 (N_45721,N_44645,N_44632);
or U45722 (N_45722,N_44279,N_44402);
xnor U45723 (N_45723,N_44092,N_44593);
or U45724 (N_45724,N_43969,N_43632);
xor U45725 (N_45725,N_44248,N_43326);
and U45726 (N_45726,N_43697,N_44563);
or U45727 (N_45727,N_44932,N_42572);
or U45728 (N_45728,N_43810,N_42635);
or U45729 (N_45729,N_44316,N_44847);
nand U45730 (N_45730,N_44922,N_43259);
nand U45731 (N_45731,N_43756,N_44519);
nand U45732 (N_45732,N_43671,N_43117);
xor U45733 (N_45733,N_43670,N_43207);
nand U45734 (N_45734,N_43515,N_42781);
nor U45735 (N_45735,N_44264,N_42528);
or U45736 (N_45736,N_42687,N_44324);
and U45737 (N_45737,N_44533,N_43747);
nor U45738 (N_45738,N_44838,N_43482);
or U45739 (N_45739,N_43661,N_44877);
or U45740 (N_45740,N_42590,N_42607);
nand U45741 (N_45741,N_42891,N_43607);
nand U45742 (N_45742,N_43875,N_43215);
nor U45743 (N_45743,N_43265,N_42649);
and U45744 (N_45744,N_42664,N_42755);
and U45745 (N_45745,N_44194,N_44851);
nand U45746 (N_45746,N_44493,N_43934);
or U45747 (N_45747,N_42544,N_44064);
or U45748 (N_45748,N_43415,N_44809);
and U45749 (N_45749,N_43742,N_44432);
or U45750 (N_45750,N_43686,N_44381);
xnor U45751 (N_45751,N_43419,N_43665);
or U45752 (N_45752,N_42700,N_42758);
nand U45753 (N_45753,N_44078,N_43874);
xnor U45754 (N_45754,N_44169,N_44022);
or U45755 (N_45755,N_44041,N_44872);
or U45756 (N_45756,N_44803,N_43451);
or U45757 (N_45757,N_44445,N_43065);
and U45758 (N_45758,N_44631,N_44520);
or U45759 (N_45759,N_42994,N_43855);
nor U45760 (N_45760,N_44635,N_44485);
and U45761 (N_45761,N_44412,N_42807);
nand U45762 (N_45762,N_44430,N_44768);
nand U45763 (N_45763,N_44949,N_43350);
or U45764 (N_45764,N_44343,N_42522);
nor U45765 (N_45765,N_43935,N_43782);
nand U45766 (N_45766,N_43455,N_44749);
nand U45767 (N_45767,N_43373,N_43611);
nor U45768 (N_45768,N_43696,N_43227);
or U45769 (N_45769,N_43313,N_43315);
nor U45770 (N_45770,N_43524,N_44546);
nor U45771 (N_45771,N_43110,N_44135);
nor U45772 (N_45772,N_43484,N_44425);
and U45773 (N_45773,N_44244,N_42608);
nand U45774 (N_45774,N_44820,N_44840);
and U45775 (N_45775,N_44188,N_43797);
nand U45776 (N_45776,N_44333,N_42577);
and U45777 (N_45777,N_44060,N_44045);
nor U45778 (N_45778,N_44978,N_42676);
nor U45779 (N_45779,N_42671,N_43950);
and U45780 (N_45780,N_44839,N_42631);
nand U45781 (N_45781,N_44853,N_44336);
or U45782 (N_45782,N_43237,N_44329);
or U45783 (N_45783,N_42805,N_43650);
or U45784 (N_45784,N_42898,N_44887);
xor U45785 (N_45785,N_44036,N_44783);
or U45786 (N_45786,N_43750,N_44355);
or U45787 (N_45787,N_43430,N_44950);
nand U45788 (N_45788,N_43398,N_43341);
or U45789 (N_45789,N_43328,N_43165);
and U45790 (N_45790,N_43228,N_43559);
or U45791 (N_45791,N_42643,N_43792);
and U45792 (N_45792,N_44833,N_43980);
or U45793 (N_45793,N_43529,N_43649);
and U45794 (N_45794,N_43384,N_44752);
nor U45795 (N_45795,N_44217,N_44944);
xnor U45796 (N_45796,N_43078,N_42756);
and U45797 (N_45797,N_44796,N_43162);
and U45798 (N_45798,N_42689,N_44172);
nor U45799 (N_45799,N_43849,N_43706);
nand U45800 (N_45800,N_44253,N_42836);
xor U45801 (N_45801,N_44975,N_43290);
or U45802 (N_45802,N_43112,N_43918);
and U45803 (N_45803,N_44793,N_43257);
or U45804 (N_45804,N_43833,N_43966);
or U45805 (N_45805,N_44089,N_43916);
nand U45806 (N_45806,N_44503,N_44960);
and U45807 (N_45807,N_43248,N_42813);
and U45808 (N_45808,N_42830,N_44795);
nand U45809 (N_45809,N_44462,N_44360);
and U45810 (N_45810,N_44003,N_43072);
and U45811 (N_45811,N_43653,N_44354);
and U45812 (N_45812,N_42618,N_43273);
nor U45813 (N_45813,N_44027,N_44771);
and U45814 (N_45814,N_44845,N_43549);
or U45815 (N_45815,N_43202,N_42531);
and U45816 (N_45816,N_43414,N_42826);
nor U45817 (N_45817,N_44368,N_44295);
nor U45818 (N_45818,N_43850,N_44031);
or U45819 (N_45819,N_44044,N_42764);
and U45820 (N_45820,N_44407,N_44481);
nor U45821 (N_45821,N_44030,N_44119);
nor U45822 (N_45822,N_44541,N_42849);
nand U45823 (N_45823,N_43106,N_44634);
or U45824 (N_45824,N_43105,N_43037);
and U45825 (N_45825,N_43470,N_43407);
nand U45826 (N_45826,N_43795,N_44164);
or U45827 (N_45827,N_43115,N_43746);
nand U45828 (N_45828,N_42904,N_44837);
xor U45829 (N_45829,N_43974,N_44810);
nor U45830 (N_45830,N_43527,N_43705);
nand U45831 (N_45831,N_44302,N_44573);
xor U45832 (N_45832,N_43387,N_44191);
and U45833 (N_45833,N_43597,N_44609);
and U45834 (N_45834,N_42519,N_44038);
or U45835 (N_45835,N_44183,N_44029);
and U45836 (N_45836,N_42990,N_43149);
and U45837 (N_45837,N_43146,N_43420);
nor U45838 (N_45838,N_42774,N_43955);
nor U45839 (N_45839,N_44763,N_43321);
nand U45840 (N_45840,N_44118,N_43947);
and U45841 (N_45841,N_43642,N_43688);
and U45842 (N_45842,N_42669,N_42730);
nor U45843 (N_45843,N_43618,N_43631);
or U45844 (N_45844,N_42551,N_42797);
and U45845 (N_45845,N_44104,N_44553);
xnor U45846 (N_45846,N_43923,N_43596);
or U45847 (N_45847,N_44210,N_43589);
and U45848 (N_45848,N_44428,N_44467);
nand U45849 (N_45849,N_43301,N_44495);
and U45850 (N_45850,N_42796,N_44426);
and U45851 (N_45851,N_44623,N_43993);
nor U45852 (N_45852,N_44767,N_44453);
and U45853 (N_45853,N_43390,N_44122);
nor U45854 (N_45854,N_43608,N_44035);
nand U45855 (N_45855,N_44021,N_44179);
or U45856 (N_45856,N_43681,N_44924);
xnor U45857 (N_45857,N_42570,N_44613);
and U45858 (N_45858,N_43844,N_44656);
xor U45859 (N_45859,N_43620,N_44094);
nor U45860 (N_45860,N_43436,N_44787);
nand U45861 (N_45861,N_44904,N_42532);
nor U45862 (N_45862,N_44906,N_44204);
or U45863 (N_45863,N_43151,N_44962);
and U45864 (N_45864,N_44530,N_43737);
xor U45865 (N_45865,N_44454,N_43754);
and U45866 (N_45866,N_43541,N_43490);
and U45867 (N_45867,N_43601,N_43137);
nor U45868 (N_45868,N_42766,N_43109);
and U45869 (N_45869,N_42697,N_43741);
or U45870 (N_45870,N_42911,N_44884);
nand U45871 (N_45871,N_44196,N_43459);
nand U45872 (N_45872,N_43573,N_43425);
and U45873 (N_45873,N_43216,N_44337);
nand U45874 (N_45874,N_44250,N_44952);
nand U45875 (N_45875,N_43921,N_44855);
nor U45876 (N_45876,N_42892,N_44318);
and U45877 (N_45877,N_43199,N_44579);
or U45878 (N_45878,N_43956,N_42975);
and U45879 (N_45879,N_42557,N_43014);
nand U45880 (N_45880,N_43231,N_43660);
nand U45881 (N_45881,N_42914,N_44193);
xnor U45882 (N_45882,N_44440,N_43279);
nor U45883 (N_45883,N_44619,N_42917);
and U45884 (N_45884,N_44184,N_44448);
nor U45885 (N_45885,N_44418,N_43499);
nor U45886 (N_45886,N_43466,N_42503);
nor U45887 (N_45887,N_44420,N_43125);
and U45888 (N_45888,N_43851,N_43472);
and U45889 (N_45889,N_44223,N_44730);
nor U45890 (N_45890,N_44186,N_43749);
nand U45891 (N_45891,N_43041,N_44207);
nor U45892 (N_45892,N_42746,N_43863);
nor U45893 (N_45893,N_44655,N_43659);
or U45894 (N_45894,N_44574,N_43579);
xor U45895 (N_45895,N_42554,N_43920);
nand U45896 (N_45896,N_44257,N_44867);
and U45897 (N_45897,N_43423,N_43519);
nor U45898 (N_45898,N_44740,N_44361);
nor U45899 (N_45899,N_42506,N_43084);
nand U45900 (N_45900,N_42804,N_44242);
nand U45901 (N_45901,N_43606,N_43187);
and U45902 (N_45902,N_44518,N_42921);
nor U45903 (N_45903,N_44512,N_44227);
nand U45904 (N_45904,N_43458,N_43452);
and U45905 (N_45905,N_42876,N_43893);
and U45906 (N_45906,N_43508,N_43444);
nor U45907 (N_45907,N_44757,N_44490);
nor U45908 (N_45908,N_42533,N_43157);
or U45909 (N_45909,N_43542,N_43073);
and U45910 (N_45910,N_43823,N_43303);
nand U45911 (N_45911,N_43213,N_44979);
xnor U45912 (N_45912,N_44347,N_43111);
or U45913 (N_45913,N_44376,N_43822);
nor U45914 (N_45914,N_44479,N_43520);
nor U45915 (N_45915,N_43069,N_44667);
nand U45916 (N_45916,N_43193,N_44466);
or U45917 (N_45917,N_43225,N_42930);
or U45918 (N_45918,N_44569,N_42762);
or U45919 (N_45919,N_43873,N_44160);
nor U45920 (N_45920,N_43282,N_42639);
and U45921 (N_45921,N_43612,N_44666);
nor U45922 (N_45922,N_42714,N_44421);
nand U45923 (N_45923,N_42742,N_44566);
or U45924 (N_45924,N_44074,N_43765);
and U45925 (N_45925,N_43081,N_44641);
or U45926 (N_45926,N_44547,N_44524);
and U45927 (N_45927,N_44251,N_43261);
nand U45928 (N_45928,N_44689,N_43583);
or U45929 (N_45929,N_44615,N_44931);
xor U45930 (N_45930,N_44626,N_43120);
nand U45931 (N_45931,N_44274,N_43201);
or U45932 (N_45932,N_43346,N_44110);
nand U45933 (N_45933,N_44505,N_44471);
nor U45934 (N_45934,N_42595,N_44332);
nor U45935 (N_45935,N_42775,N_43314);
and U45936 (N_45936,N_43128,N_44423);
nand U45937 (N_45937,N_44557,N_43807);
or U45938 (N_45938,N_42827,N_44007);
nor U45939 (N_45939,N_44097,N_42920);
and U45940 (N_45940,N_43838,N_44344);
xnor U45941 (N_45941,N_44287,N_44873);
nand U45942 (N_45942,N_43172,N_44928);
or U45943 (N_45943,N_44349,N_42734);
nor U45944 (N_45944,N_44598,N_43196);
and U45945 (N_45945,N_44515,N_43351);
nor U45946 (N_45946,N_44821,N_43242);
nor U45947 (N_45947,N_43837,N_43431);
xnor U45948 (N_45948,N_42759,N_42692);
and U45949 (N_45949,N_44386,N_42980);
or U45950 (N_45950,N_44341,N_44054);
and U45951 (N_45951,N_42682,N_44198);
nand U45952 (N_45952,N_42787,N_44994);
xor U45953 (N_45953,N_42617,N_43926);
nor U45954 (N_45954,N_42561,N_44968);
and U45955 (N_45955,N_42808,N_43252);
nand U45956 (N_45956,N_43318,N_44382);
nand U45957 (N_45957,N_44697,N_43840);
or U45958 (N_45958,N_44614,N_43214);
nand U45959 (N_45959,N_44942,N_44213);
and U45960 (N_45960,N_43432,N_43927);
or U45961 (N_45961,N_42530,N_43647);
nand U45962 (N_45962,N_44555,N_42874);
or U45963 (N_45963,N_44049,N_43158);
nand U45964 (N_45964,N_44208,N_43610);
xor U45965 (N_45965,N_43129,N_44502);
or U45966 (N_45966,N_43768,N_44836);
and U45967 (N_45967,N_42655,N_44663);
and U45968 (N_45968,N_43412,N_43370);
nor U45969 (N_45969,N_42908,N_44724);
and U45970 (N_45970,N_44668,N_44151);
and U45971 (N_45971,N_43676,N_43619);
and U45972 (N_45972,N_42744,N_44759);
nand U45973 (N_45973,N_43085,N_43881);
nand U45974 (N_45974,N_42549,N_44850);
and U45975 (N_45975,N_43008,N_44594);
xnor U45976 (N_45976,N_43056,N_43173);
or U45977 (N_45977,N_43293,N_44309);
nor U45978 (N_45978,N_43931,N_43224);
xnor U45979 (N_45979,N_42829,N_43264);
or U45980 (N_45980,N_44545,N_43627);
nor U45981 (N_45981,N_44976,N_42811);
nor U45982 (N_45982,N_43560,N_43717);
xnor U45983 (N_45983,N_44284,N_43500);
and U45984 (N_45984,N_43628,N_44841);
xor U45985 (N_45985,N_42502,N_43938);
or U45986 (N_45986,N_44398,N_43988);
nand U45987 (N_45987,N_44826,N_42852);
nor U45988 (N_45988,N_44818,N_43210);
and U45989 (N_45989,N_44447,N_43814);
or U45990 (N_45990,N_43630,N_43819);
and U45991 (N_45991,N_44289,N_42896);
or U45992 (N_45992,N_43200,N_44649);
and U45993 (N_45993,N_44127,N_44307);
or U45994 (N_45994,N_44618,N_42761);
nand U45995 (N_45995,N_42964,N_43772);
nor U45996 (N_45996,N_42837,N_44082);
and U45997 (N_45997,N_44532,N_42933);
nand U45998 (N_45998,N_43783,N_44051);
xnor U45999 (N_45999,N_42568,N_44577);
and U46000 (N_46000,N_43344,N_43984);
xor U46001 (N_46001,N_43058,N_44961);
nor U46002 (N_46002,N_44926,N_43617);
nand U46003 (N_46003,N_43760,N_44374);
and U46004 (N_46004,N_43806,N_44048);
nand U46005 (N_46005,N_44534,N_44059);
nand U46006 (N_46006,N_43533,N_43450);
and U46007 (N_46007,N_44921,N_44781);
or U46008 (N_46008,N_43234,N_43253);
nor U46009 (N_46009,N_42846,N_44601);
xor U46010 (N_46010,N_44537,N_42739);
nor U46011 (N_46011,N_43156,N_44061);
and U46012 (N_46012,N_42879,N_44510);
xor U46013 (N_46013,N_43277,N_44239);
nor U46014 (N_46014,N_43097,N_44443);
and U46015 (N_46015,N_44865,N_42750);
nor U46016 (N_46016,N_43852,N_44997);
nand U46017 (N_46017,N_44134,N_44843);
nor U46018 (N_46018,N_43609,N_42555);
nor U46019 (N_46019,N_42882,N_43906);
nand U46020 (N_46020,N_42909,N_42870);
and U46021 (N_46021,N_42950,N_44633);
nand U46022 (N_46022,N_44116,N_43276);
nand U46023 (N_46023,N_43061,N_44894);
or U46024 (N_46024,N_44606,N_43413);
nor U46025 (N_46025,N_43577,N_43561);
nor U46026 (N_46026,N_43079,N_43226);
and U46027 (N_46027,N_42606,N_42938);
and U46028 (N_46028,N_43160,N_44895);
or U46029 (N_46029,N_44159,N_44293);
nor U46030 (N_46030,N_42599,N_43734);
xor U46031 (N_46031,N_43354,N_43114);
nor U46032 (N_46032,N_44480,N_43168);
xor U46033 (N_46033,N_43563,N_42928);
nand U46034 (N_46034,N_44475,N_44507);
and U46035 (N_46035,N_42729,N_44797);
or U46036 (N_46036,N_43979,N_43288);
and U46037 (N_46037,N_42953,N_44370);
or U46038 (N_46038,N_43803,N_44457);
nand U46039 (N_46039,N_44132,N_43353);
and U46040 (N_46040,N_43485,N_44548);
and U46041 (N_46041,N_43902,N_43505);
nor U46042 (N_46042,N_44956,N_42986);
nand U46043 (N_46043,N_42801,N_42736);
nand U46044 (N_46044,N_42589,N_43645);
nor U46045 (N_46045,N_44801,N_43952);
and U46046 (N_46046,N_44929,N_43185);
nor U46047 (N_46047,N_44335,N_43493);
and U46048 (N_46048,N_44972,N_42603);
or U46049 (N_46049,N_44162,N_43818);
and U46050 (N_46050,N_43736,N_43735);
or U46051 (N_46051,N_43638,N_43692);
and U46052 (N_46052,N_43245,N_42785);
nor U46053 (N_46053,N_44864,N_42704);
or U46054 (N_46054,N_44919,N_43071);
and U46055 (N_46055,N_43118,N_43687);
xnor U46056 (N_46056,N_43539,N_42545);
xnor U46057 (N_46057,N_42710,N_44113);
nand U46058 (N_46058,N_42752,N_44964);
nor U46059 (N_46059,N_44977,N_44023);
nand U46060 (N_46060,N_43892,N_43256);
nand U46061 (N_46061,N_44812,N_42906);
and U46062 (N_46062,N_44819,N_43770);
and U46063 (N_46063,N_43388,N_44684);
nor U46064 (N_46064,N_44701,N_44214);
and U46065 (N_46065,N_43575,N_44858);
nand U46066 (N_46066,N_44586,N_43912);
or U46067 (N_46067,N_42675,N_43591);
and U46068 (N_46068,N_42765,N_43564);
or U46069 (N_46069,N_43507,N_44996);
and U46070 (N_46070,N_44358,N_42705);
and U46071 (N_46071,N_44259,N_43592);
nand U46072 (N_46072,N_43629,N_44240);
and U46073 (N_46073,N_43669,N_43511);
or U46074 (N_46074,N_43738,N_42842);
or U46075 (N_46075,N_43333,N_44710);
nor U46076 (N_46076,N_44832,N_42915);
or U46077 (N_46077,N_44101,N_43403);
and U46078 (N_46078,N_44154,N_43694);
and U46079 (N_46079,N_43558,N_43342);
or U46080 (N_46080,N_43090,N_44985);
and U46081 (N_46081,N_44879,N_43972);
nand U46082 (N_46082,N_43171,N_43545);
nand U46083 (N_46083,N_43053,N_43986);
nor U46084 (N_46084,N_43907,N_43238);
nor U46085 (N_46085,N_43805,N_42711);
or U46086 (N_46086,N_42661,N_43271);
xnor U46087 (N_46087,N_42564,N_43345);
and U46088 (N_46088,N_43785,N_44378);
or U46089 (N_46089,N_44717,N_44798);
and U46090 (N_46090,N_43946,N_43512);
nand U46091 (N_46091,N_44487,N_43358);
xor U46092 (N_46092,N_44943,N_44762);
nor U46093 (N_46093,N_44301,N_44450);
nand U46094 (N_46094,N_42973,N_44580);
nor U46095 (N_46095,N_43212,N_44991);
nand U46096 (N_46096,N_43286,N_42959);
or U46097 (N_46097,N_44804,N_44731);
or U46098 (N_46098,N_44817,N_44637);
nor U46099 (N_46099,N_44197,N_43409);
or U46100 (N_46100,N_44504,N_43439);
or U46101 (N_46101,N_42674,N_44971);
or U46102 (N_46102,N_43504,N_42828);
nor U46103 (N_46103,N_43531,N_44362);
nand U46104 (N_46104,N_43555,N_44424);
and U46105 (N_46105,N_43104,N_42770);
nor U46106 (N_46106,N_43364,N_44396);
or U46107 (N_46107,N_43502,N_43830);
and U46108 (N_46108,N_43464,N_42709);
and U46109 (N_46109,N_42825,N_43883);
or U46110 (N_46110,N_42881,N_44435);
and U46111 (N_46111,N_44946,N_44693);
nor U46112 (N_46112,N_42713,N_42695);
nand U46113 (N_46113,N_43864,N_42779);
nor U46114 (N_46114,N_43853,N_43652);
nand U46115 (N_46115,N_44918,N_44053);
xor U46116 (N_46116,N_42843,N_44692);
and U46117 (N_46117,N_43684,N_44121);
or U46118 (N_46118,N_44785,N_44177);
and U46119 (N_46119,N_43538,N_44464);
or U46120 (N_46120,N_44093,N_42878);
nor U46121 (N_46121,N_43272,N_42989);
nand U46122 (N_46122,N_44006,N_44591);
nand U46123 (N_46123,N_42507,N_43543);
nor U46124 (N_46124,N_44182,N_43481);
xnor U46125 (N_46125,N_43148,N_42967);
or U46126 (N_46126,N_43365,N_43858);
and U46127 (N_46127,N_44600,N_44708);
nand U46128 (N_46128,N_43461,N_43401);
or U46129 (N_46129,N_44304,N_44232);
nor U46130 (N_46130,N_43209,N_43801);
nand U46131 (N_46131,N_44802,N_44612);
nor U46132 (N_46132,N_44983,N_44848);
or U46133 (N_46133,N_44237,N_42745);
nand U46134 (N_46134,N_44815,N_42740);
and U46135 (N_46135,N_42954,N_43691);
and U46136 (N_46136,N_42974,N_44538);
or U46137 (N_46137,N_43154,N_42581);
or U46138 (N_46138,N_42588,N_42504);
xor U46139 (N_46139,N_42685,N_44682);
nand U46140 (N_46140,N_43389,N_44704);
nand U46141 (N_46141,N_42723,N_44229);
or U46142 (N_46142,N_44627,N_42509);
or U46143 (N_46143,N_43189,N_42782);
nand U46144 (N_46144,N_44620,N_44862);
nand U46145 (N_46145,N_44677,N_42560);
nand U46146 (N_46146,N_44245,N_44982);
and U46147 (N_46147,N_43140,N_43285);
xor U46148 (N_46148,N_43503,N_43553);
and U46149 (N_46149,N_42575,N_43804);
and U46150 (N_46150,N_42997,N_44458);
nand U46151 (N_46151,N_43685,N_44916);
xor U46152 (N_46152,N_43525,N_42735);
and U46153 (N_46153,N_43826,N_44281);
xnor U46154 (N_46154,N_44679,N_44389);
and U46155 (N_46155,N_44900,N_44124);
nand U46156 (N_46156,N_44688,N_44405);
nand U46157 (N_46157,N_44077,N_42720);
nand U46158 (N_46158,N_43616,N_43217);
nor U46159 (N_46159,N_44660,N_42925);
and U46160 (N_46160,N_44225,N_44751);
nand U46161 (N_46161,N_44437,N_44139);
nand U46162 (N_46162,N_42521,N_44422);
nor U46163 (N_46163,N_43410,N_44288);
and U46164 (N_46164,N_44322,N_44052);
nand U46165 (N_46165,N_43970,N_43454);
or U46166 (N_46166,N_42812,N_44823);
nand U46167 (N_46167,N_44745,N_44408);
nand U46168 (N_46168,N_42540,N_42760);
nor U46169 (N_46169,N_44461,N_44328);
or U46170 (N_46170,N_44050,N_42587);
nand U46171 (N_46171,N_44473,N_44226);
or U46172 (N_46172,N_43262,N_44786);
nor U46173 (N_46173,N_43011,N_43266);
or U46174 (N_46174,N_43924,N_43964);
or U46175 (N_46175,N_44827,N_44306);
or U46176 (N_46176,N_43633,N_44907);
or U46177 (N_46177,N_44849,N_44951);
nand U46178 (N_46178,N_44131,N_43766);
and U46179 (N_46179,N_44969,N_42875);
xnor U46180 (N_46180,N_43509,N_42960);
xnor U46181 (N_46181,N_43121,N_44732);
and U46182 (N_46182,N_43777,N_44008);
nor U46183 (N_46183,N_44103,N_44438);
nor U46184 (N_46184,N_42683,N_42514);
xor U46185 (N_46185,N_43270,N_44115);
nor U46186 (N_46186,N_43347,N_42948);
nand U46187 (N_46187,N_44883,N_42621);
or U46188 (N_46188,N_43438,N_44321);
nor U46189 (N_46189,N_44460,N_42534);
nor U46190 (N_46190,N_43244,N_43654);
or U46191 (N_46191,N_44246,N_43486);
nor U46192 (N_46192,N_42594,N_43732);
or U46193 (N_46193,N_43032,N_43487);
xor U46194 (N_46194,N_44987,N_43010);
or U46195 (N_46195,N_43102,N_43460);
and U46196 (N_46196,N_43598,N_42662);
xor U46197 (N_46197,N_43457,N_42637);
and U46198 (N_46198,N_44323,N_44528);
or U46199 (N_46199,N_42673,N_44254);
or U46200 (N_46200,N_44073,N_42803);
or U46201 (N_46201,N_44303,N_44890);
and U46202 (N_46202,N_43963,N_44874);
nand U46203 (N_46203,N_42929,N_43901);
xor U46204 (N_46204,N_43024,N_42767);
or U46205 (N_46205,N_43682,N_44330);
nand U46206 (N_46206,N_44678,N_43309);
nor U46207 (N_46207,N_43139,N_44764);
and U46208 (N_46208,N_43860,N_43786);
and U46209 (N_46209,N_43621,N_44638);
nor U46210 (N_46210,N_44945,N_44527);
nand U46211 (N_46211,N_43471,N_43360);
and U46212 (N_46212,N_43999,N_42968);
nor U46213 (N_46213,N_43821,N_44419);
xnor U46214 (N_46214,N_43870,N_43889);
and U46215 (N_46215,N_44622,N_43302);
or U46216 (N_46216,N_44014,N_44413);
nand U46217 (N_46217,N_42883,N_43894);
xnor U46218 (N_46218,N_42650,N_44644);
and U46219 (N_46219,N_43624,N_44200);
nand U46220 (N_46220,N_42936,N_42614);
or U46221 (N_46221,N_44180,N_44215);
nor U46222 (N_46222,N_44672,N_44072);
nor U46223 (N_46223,N_43876,N_44046);
nand U46224 (N_46224,N_43604,N_43514);
and U46225 (N_46225,N_42527,N_42501);
and U46226 (N_46226,N_43211,N_43051);
nor U46227 (N_46227,N_44236,N_43832);
and U46228 (N_46228,N_44741,N_44769);
nand U46229 (N_46229,N_42824,N_42952);
nand U46230 (N_46230,N_44373,N_43393);
xor U46231 (N_46231,N_43516,N_43379);
or U46232 (N_46232,N_43233,N_43574);
nand U46233 (N_46233,N_42778,N_44980);
or U46234 (N_46234,N_43015,N_43179);
nor U46235 (N_46235,N_44899,N_44296);
or U46236 (N_46236,N_43701,N_44417);
and U46237 (N_46237,N_43038,N_42562);
or U46238 (N_46238,N_42939,N_44937);
and U46239 (N_46239,N_44542,N_44876);
and U46240 (N_46240,N_42518,N_42982);
or U46241 (N_46241,N_44711,N_43847);
and U46242 (N_46242,N_43856,N_43166);
nor U46243 (N_46243,N_43953,N_43044);
nand U46244 (N_46244,N_43995,N_43816);
or U46245 (N_46245,N_43712,N_43435);
and U46246 (N_46246,N_44397,N_42666);
or U46247 (N_46247,N_42970,N_42850);
and U46248 (N_46248,N_43000,N_44353);
or U46249 (N_46249,N_43427,N_44013);
nor U46250 (N_46250,N_44273,N_44795);
and U46251 (N_46251,N_44068,N_44417);
and U46252 (N_46252,N_43127,N_42867);
nor U46253 (N_46253,N_44202,N_43900);
and U46254 (N_46254,N_44563,N_44622);
nand U46255 (N_46255,N_43550,N_43085);
and U46256 (N_46256,N_44464,N_43174);
and U46257 (N_46257,N_44544,N_43778);
nand U46258 (N_46258,N_44504,N_43084);
or U46259 (N_46259,N_44780,N_42617);
nand U46260 (N_46260,N_44807,N_44720);
and U46261 (N_46261,N_44294,N_42599);
xnor U46262 (N_46262,N_44818,N_43022);
nor U46263 (N_46263,N_43283,N_44813);
nor U46264 (N_46264,N_44016,N_44738);
nor U46265 (N_46265,N_44177,N_44533);
and U46266 (N_46266,N_43437,N_42526);
nor U46267 (N_46267,N_43617,N_43908);
or U46268 (N_46268,N_44907,N_43110);
nor U46269 (N_46269,N_44702,N_42859);
nor U46270 (N_46270,N_44939,N_44812);
and U46271 (N_46271,N_44398,N_44482);
nand U46272 (N_46272,N_42582,N_43247);
xor U46273 (N_46273,N_43774,N_42997);
or U46274 (N_46274,N_44600,N_44169);
or U46275 (N_46275,N_43006,N_43615);
or U46276 (N_46276,N_42901,N_43063);
nor U46277 (N_46277,N_44828,N_44352);
or U46278 (N_46278,N_43155,N_44195);
nor U46279 (N_46279,N_43053,N_44439);
and U46280 (N_46280,N_43896,N_43508);
xnor U46281 (N_46281,N_43460,N_43385);
nor U46282 (N_46282,N_42943,N_44654);
nor U46283 (N_46283,N_44754,N_43569);
nor U46284 (N_46284,N_42837,N_44713);
or U46285 (N_46285,N_42710,N_43900);
and U46286 (N_46286,N_44321,N_42737);
nand U46287 (N_46287,N_43982,N_43111);
nor U46288 (N_46288,N_43908,N_44280);
nor U46289 (N_46289,N_43097,N_44148);
nor U46290 (N_46290,N_44127,N_43158);
and U46291 (N_46291,N_42513,N_42701);
or U46292 (N_46292,N_43420,N_42811);
nor U46293 (N_46293,N_43469,N_42656);
nor U46294 (N_46294,N_42680,N_42719);
or U46295 (N_46295,N_44726,N_43414);
or U46296 (N_46296,N_43752,N_43749);
and U46297 (N_46297,N_43838,N_44564);
and U46298 (N_46298,N_43066,N_44542);
nand U46299 (N_46299,N_43722,N_44933);
and U46300 (N_46300,N_44570,N_44503);
nand U46301 (N_46301,N_42542,N_42614);
nand U46302 (N_46302,N_43833,N_43063);
nor U46303 (N_46303,N_44110,N_44661);
nand U46304 (N_46304,N_44105,N_44173);
and U46305 (N_46305,N_44238,N_44044);
and U46306 (N_46306,N_43049,N_43889);
xor U46307 (N_46307,N_44930,N_43236);
or U46308 (N_46308,N_44172,N_43983);
xor U46309 (N_46309,N_42926,N_43664);
nor U46310 (N_46310,N_44659,N_43244);
nor U46311 (N_46311,N_43206,N_44860);
or U46312 (N_46312,N_44191,N_43643);
nor U46313 (N_46313,N_44418,N_43674);
nor U46314 (N_46314,N_42978,N_44455);
or U46315 (N_46315,N_43944,N_44793);
nand U46316 (N_46316,N_43047,N_43427);
or U46317 (N_46317,N_43867,N_44708);
and U46318 (N_46318,N_43931,N_44432);
nor U46319 (N_46319,N_44283,N_43190);
xnor U46320 (N_46320,N_44461,N_43825);
nand U46321 (N_46321,N_44966,N_44324);
xnor U46322 (N_46322,N_44941,N_44329);
or U46323 (N_46323,N_44361,N_44467);
or U46324 (N_46324,N_43016,N_43581);
nor U46325 (N_46325,N_44910,N_43294);
or U46326 (N_46326,N_42756,N_44671);
nand U46327 (N_46327,N_42643,N_44870);
xor U46328 (N_46328,N_43702,N_44079);
or U46329 (N_46329,N_44481,N_43566);
nor U46330 (N_46330,N_44053,N_42744);
nand U46331 (N_46331,N_43597,N_44525);
nand U46332 (N_46332,N_44664,N_44317);
nand U46333 (N_46333,N_43173,N_44476);
or U46334 (N_46334,N_43793,N_44596);
nand U46335 (N_46335,N_42872,N_43912);
nor U46336 (N_46336,N_44295,N_44454);
nor U46337 (N_46337,N_43646,N_42500);
nand U46338 (N_46338,N_44076,N_42804);
and U46339 (N_46339,N_43314,N_42947);
nor U46340 (N_46340,N_43586,N_42647);
or U46341 (N_46341,N_44245,N_44503);
and U46342 (N_46342,N_42909,N_44170);
nand U46343 (N_46343,N_44118,N_44881);
and U46344 (N_46344,N_43654,N_44226);
nor U46345 (N_46345,N_44391,N_44496);
and U46346 (N_46346,N_44280,N_43398);
nand U46347 (N_46347,N_43026,N_43765);
and U46348 (N_46348,N_44750,N_44266);
nand U46349 (N_46349,N_43568,N_43217);
or U46350 (N_46350,N_44615,N_44333);
nor U46351 (N_46351,N_43381,N_44678);
or U46352 (N_46352,N_42554,N_44855);
or U46353 (N_46353,N_43646,N_44708);
and U46354 (N_46354,N_43015,N_43573);
or U46355 (N_46355,N_43187,N_44416);
and U46356 (N_46356,N_44863,N_42732);
xnor U46357 (N_46357,N_42606,N_44133);
and U46358 (N_46358,N_43589,N_43005);
nand U46359 (N_46359,N_43136,N_43765);
nor U46360 (N_46360,N_43272,N_42895);
or U46361 (N_46361,N_44785,N_43547);
nand U46362 (N_46362,N_43092,N_44633);
and U46363 (N_46363,N_43404,N_44535);
nor U46364 (N_46364,N_43610,N_43757);
nor U46365 (N_46365,N_44409,N_43207);
nor U46366 (N_46366,N_43446,N_44241);
nand U46367 (N_46367,N_43455,N_44981);
xor U46368 (N_46368,N_43365,N_43295);
or U46369 (N_46369,N_43839,N_44434);
or U46370 (N_46370,N_44298,N_42766);
nor U46371 (N_46371,N_43058,N_44048);
or U46372 (N_46372,N_42810,N_43523);
or U46373 (N_46373,N_44007,N_44204);
and U46374 (N_46374,N_43461,N_43775);
nand U46375 (N_46375,N_44369,N_43530);
or U46376 (N_46376,N_44369,N_44452);
or U46377 (N_46377,N_43993,N_43546);
nand U46378 (N_46378,N_43779,N_44942);
or U46379 (N_46379,N_44117,N_43748);
nand U46380 (N_46380,N_42787,N_43368);
and U46381 (N_46381,N_44569,N_42982);
xnor U46382 (N_46382,N_44334,N_42520);
nor U46383 (N_46383,N_44387,N_44372);
nand U46384 (N_46384,N_44204,N_43999);
xnor U46385 (N_46385,N_44092,N_43737);
xor U46386 (N_46386,N_43326,N_43225);
nand U46387 (N_46387,N_44827,N_42854);
nor U46388 (N_46388,N_42527,N_44706);
or U46389 (N_46389,N_42714,N_44575);
nor U46390 (N_46390,N_42904,N_44643);
or U46391 (N_46391,N_44827,N_44410);
or U46392 (N_46392,N_44539,N_43736);
or U46393 (N_46393,N_43345,N_42818);
nor U46394 (N_46394,N_43092,N_43194);
and U46395 (N_46395,N_44159,N_42700);
xnor U46396 (N_46396,N_43130,N_44556);
and U46397 (N_46397,N_44111,N_44485);
nor U46398 (N_46398,N_44475,N_42508);
nor U46399 (N_46399,N_44128,N_44957);
nand U46400 (N_46400,N_43636,N_44905);
nand U46401 (N_46401,N_44627,N_44192);
or U46402 (N_46402,N_44785,N_44791);
nand U46403 (N_46403,N_42727,N_43170);
xnor U46404 (N_46404,N_44620,N_43018);
nor U46405 (N_46405,N_42777,N_42557);
and U46406 (N_46406,N_44839,N_44512);
nor U46407 (N_46407,N_42959,N_43525);
and U46408 (N_46408,N_43160,N_44040);
xnor U46409 (N_46409,N_44571,N_44996);
nor U46410 (N_46410,N_42958,N_43898);
nand U46411 (N_46411,N_44308,N_43285);
or U46412 (N_46412,N_44262,N_42549);
and U46413 (N_46413,N_42873,N_44404);
nor U46414 (N_46414,N_42768,N_43208);
nand U46415 (N_46415,N_42528,N_43429);
nor U46416 (N_46416,N_42795,N_42568);
nand U46417 (N_46417,N_44508,N_43405);
or U46418 (N_46418,N_42655,N_43763);
or U46419 (N_46419,N_44343,N_43966);
or U46420 (N_46420,N_44168,N_44473);
nor U46421 (N_46421,N_44544,N_43328);
nand U46422 (N_46422,N_42633,N_43263);
nand U46423 (N_46423,N_43946,N_44767);
or U46424 (N_46424,N_43213,N_43630);
or U46425 (N_46425,N_44062,N_44530);
or U46426 (N_46426,N_44522,N_43281);
nor U46427 (N_46427,N_43247,N_44548);
nor U46428 (N_46428,N_42711,N_44343);
nor U46429 (N_46429,N_43186,N_42873);
and U46430 (N_46430,N_42593,N_44449);
or U46431 (N_46431,N_42955,N_43056);
or U46432 (N_46432,N_44209,N_44324);
nor U46433 (N_46433,N_42869,N_43207);
nor U46434 (N_46434,N_43298,N_43806);
xor U46435 (N_46435,N_44623,N_43600);
and U46436 (N_46436,N_44724,N_43522);
nand U46437 (N_46437,N_42516,N_42630);
xor U46438 (N_46438,N_44555,N_44871);
or U46439 (N_46439,N_44239,N_42732);
or U46440 (N_46440,N_43038,N_43929);
nand U46441 (N_46441,N_44118,N_44230);
nand U46442 (N_46442,N_44150,N_44599);
nor U46443 (N_46443,N_43134,N_43039);
or U46444 (N_46444,N_42737,N_42824);
and U46445 (N_46445,N_43777,N_44073);
nand U46446 (N_46446,N_43469,N_43939);
and U46447 (N_46447,N_44374,N_43057);
or U46448 (N_46448,N_44446,N_42872);
and U46449 (N_46449,N_44568,N_43342);
and U46450 (N_46450,N_43122,N_44678);
nor U46451 (N_46451,N_43209,N_43886);
nand U46452 (N_46452,N_44981,N_42827);
and U46453 (N_46453,N_42926,N_42505);
nand U46454 (N_46454,N_44245,N_44145);
nor U46455 (N_46455,N_43259,N_44849);
and U46456 (N_46456,N_44467,N_42955);
nand U46457 (N_46457,N_43855,N_42971);
xnor U46458 (N_46458,N_44798,N_42512);
and U46459 (N_46459,N_43954,N_43683);
or U46460 (N_46460,N_43507,N_43295);
nor U46461 (N_46461,N_43016,N_44115);
or U46462 (N_46462,N_43177,N_43850);
or U46463 (N_46463,N_44233,N_44622);
nand U46464 (N_46464,N_44177,N_42595);
nand U46465 (N_46465,N_44725,N_44507);
nand U46466 (N_46466,N_43993,N_43698);
or U46467 (N_46467,N_43103,N_44149);
nand U46468 (N_46468,N_43269,N_43934);
xnor U46469 (N_46469,N_42795,N_43719);
nor U46470 (N_46470,N_43767,N_42586);
and U46471 (N_46471,N_44351,N_42797);
nor U46472 (N_46472,N_42506,N_43573);
nor U46473 (N_46473,N_43716,N_42801);
or U46474 (N_46474,N_44478,N_44178);
and U46475 (N_46475,N_44981,N_43873);
and U46476 (N_46476,N_43809,N_44577);
nor U46477 (N_46477,N_43308,N_42508);
and U46478 (N_46478,N_43061,N_44637);
nor U46479 (N_46479,N_43223,N_44503);
nand U46480 (N_46480,N_42567,N_44354);
and U46481 (N_46481,N_44323,N_43389);
or U46482 (N_46482,N_43441,N_44046);
and U46483 (N_46483,N_44408,N_44773);
and U46484 (N_46484,N_43426,N_42709);
or U46485 (N_46485,N_43188,N_43679);
or U46486 (N_46486,N_43881,N_44232);
or U46487 (N_46487,N_42902,N_44110);
xnor U46488 (N_46488,N_44326,N_44956);
xnor U46489 (N_46489,N_44725,N_42592);
and U46490 (N_46490,N_43684,N_44683);
or U46491 (N_46491,N_43621,N_44459);
and U46492 (N_46492,N_43765,N_42882);
and U46493 (N_46493,N_42971,N_43601);
or U46494 (N_46494,N_44702,N_44851);
nand U46495 (N_46495,N_43699,N_44701);
nand U46496 (N_46496,N_44437,N_43546);
nand U46497 (N_46497,N_42513,N_42696);
nor U46498 (N_46498,N_43802,N_42813);
nor U46499 (N_46499,N_43241,N_43257);
nand U46500 (N_46500,N_42927,N_44510);
or U46501 (N_46501,N_44339,N_42531);
and U46502 (N_46502,N_44071,N_43122);
and U46503 (N_46503,N_43906,N_43311);
nor U46504 (N_46504,N_43812,N_44087);
and U46505 (N_46505,N_43656,N_44984);
nand U46506 (N_46506,N_44921,N_43526);
nand U46507 (N_46507,N_44467,N_44906);
nand U46508 (N_46508,N_43536,N_42559);
nor U46509 (N_46509,N_43293,N_43751);
or U46510 (N_46510,N_43561,N_44096);
or U46511 (N_46511,N_44164,N_44471);
and U46512 (N_46512,N_44302,N_43055);
xnor U46513 (N_46513,N_44105,N_43299);
and U46514 (N_46514,N_43859,N_42540);
nand U46515 (N_46515,N_43069,N_43021);
xor U46516 (N_46516,N_44989,N_43446);
and U46517 (N_46517,N_43817,N_43267);
nand U46518 (N_46518,N_44204,N_44579);
nor U46519 (N_46519,N_43899,N_43949);
and U46520 (N_46520,N_43369,N_43874);
nor U46521 (N_46521,N_43306,N_42682);
and U46522 (N_46522,N_42689,N_44747);
or U46523 (N_46523,N_43435,N_43380);
and U46524 (N_46524,N_44240,N_43625);
or U46525 (N_46525,N_44022,N_44628);
nor U46526 (N_46526,N_43788,N_44988);
and U46527 (N_46527,N_44245,N_42904);
or U46528 (N_46528,N_44460,N_43499);
and U46529 (N_46529,N_43055,N_43115);
nand U46530 (N_46530,N_44989,N_44046);
nor U46531 (N_46531,N_42603,N_43988);
nor U46532 (N_46532,N_44507,N_44415);
or U46533 (N_46533,N_42853,N_44839);
nor U46534 (N_46534,N_44680,N_42517);
or U46535 (N_46535,N_42915,N_43098);
xnor U46536 (N_46536,N_44377,N_42952);
or U46537 (N_46537,N_43444,N_43742);
xnor U46538 (N_46538,N_44360,N_44338);
or U46539 (N_46539,N_43376,N_43692);
or U46540 (N_46540,N_44690,N_44553);
xnor U46541 (N_46541,N_43088,N_43184);
or U46542 (N_46542,N_43959,N_44020);
nor U46543 (N_46543,N_43721,N_43359);
and U46544 (N_46544,N_44936,N_44259);
nor U46545 (N_46545,N_43445,N_43354);
nand U46546 (N_46546,N_42959,N_43941);
or U46547 (N_46547,N_43715,N_44467);
nand U46548 (N_46548,N_44005,N_44779);
nand U46549 (N_46549,N_44577,N_44667);
nor U46550 (N_46550,N_44447,N_42651);
nand U46551 (N_46551,N_43108,N_43046);
nand U46552 (N_46552,N_44921,N_42828);
nor U46553 (N_46553,N_43217,N_43215);
nor U46554 (N_46554,N_43139,N_43275);
or U46555 (N_46555,N_44827,N_43697);
and U46556 (N_46556,N_43735,N_42894);
and U46557 (N_46557,N_44094,N_42545);
nor U46558 (N_46558,N_44626,N_43753);
and U46559 (N_46559,N_44328,N_43700);
and U46560 (N_46560,N_44902,N_44908);
nor U46561 (N_46561,N_42522,N_43584);
nand U46562 (N_46562,N_43560,N_44231);
and U46563 (N_46563,N_44821,N_43412);
nand U46564 (N_46564,N_42854,N_43857);
or U46565 (N_46565,N_44184,N_43847);
and U46566 (N_46566,N_42998,N_43716);
nand U46567 (N_46567,N_43039,N_42536);
nand U46568 (N_46568,N_44517,N_44283);
nand U46569 (N_46569,N_43511,N_44848);
nor U46570 (N_46570,N_43915,N_44617);
nor U46571 (N_46571,N_43866,N_42959);
or U46572 (N_46572,N_42841,N_44208);
xnor U46573 (N_46573,N_44929,N_44737);
nor U46574 (N_46574,N_44623,N_43479);
xor U46575 (N_46575,N_43647,N_42835);
nand U46576 (N_46576,N_44655,N_42956);
or U46577 (N_46577,N_44439,N_43573);
nor U46578 (N_46578,N_42814,N_44519);
and U46579 (N_46579,N_43210,N_43193);
and U46580 (N_46580,N_44182,N_44155);
xor U46581 (N_46581,N_44587,N_42838);
nor U46582 (N_46582,N_42968,N_44778);
or U46583 (N_46583,N_44426,N_42656);
and U46584 (N_46584,N_44624,N_43132);
and U46585 (N_46585,N_43359,N_43758);
nand U46586 (N_46586,N_44959,N_42578);
nor U46587 (N_46587,N_44415,N_43943);
nor U46588 (N_46588,N_44384,N_42772);
xnor U46589 (N_46589,N_44224,N_44251);
and U46590 (N_46590,N_43121,N_44697);
xnor U46591 (N_46591,N_43136,N_44318);
nand U46592 (N_46592,N_44122,N_43517);
xnor U46593 (N_46593,N_42837,N_44890);
nand U46594 (N_46594,N_44513,N_43748);
or U46595 (N_46595,N_44246,N_43796);
or U46596 (N_46596,N_43977,N_42549);
or U46597 (N_46597,N_44232,N_42654);
and U46598 (N_46598,N_42512,N_44000);
nand U46599 (N_46599,N_43729,N_44615);
xor U46600 (N_46600,N_42944,N_43801);
and U46601 (N_46601,N_44141,N_43372);
and U46602 (N_46602,N_44376,N_44699);
and U46603 (N_46603,N_44585,N_42788);
nand U46604 (N_46604,N_43722,N_42958);
nor U46605 (N_46605,N_42738,N_42823);
nand U46606 (N_46606,N_42517,N_43844);
nand U46607 (N_46607,N_44663,N_44741);
and U46608 (N_46608,N_42828,N_44530);
and U46609 (N_46609,N_44720,N_43830);
nand U46610 (N_46610,N_43502,N_43985);
or U46611 (N_46611,N_43859,N_44819);
xor U46612 (N_46612,N_43311,N_43982);
or U46613 (N_46613,N_44997,N_44449);
nand U46614 (N_46614,N_44911,N_43990);
xnor U46615 (N_46615,N_43602,N_44525);
nor U46616 (N_46616,N_43684,N_44421);
or U46617 (N_46617,N_42601,N_43698);
or U46618 (N_46618,N_43011,N_44224);
xnor U46619 (N_46619,N_43173,N_43239);
xor U46620 (N_46620,N_44346,N_44045);
and U46621 (N_46621,N_44629,N_43553);
nand U46622 (N_46622,N_42779,N_44639);
nor U46623 (N_46623,N_43627,N_44310);
nor U46624 (N_46624,N_44137,N_43154);
nor U46625 (N_46625,N_42804,N_43109);
and U46626 (N_46626,N_44201,N_43738);
or U46627 (N_46627,N_43441,N_43328);
or U46628 (N_46628,N_42999,N_44365);
or U46629 (N_46629,N_44030,N_43139);
and U46630 (N_46630,N_44034,N_43058);
or U46631 (N_46631,N_43956,N_44457);
xnor U46632 (N_46632,N_44020,N_42615);
or U46633 (N_46633,N_44764,N_44746);
nor U46634 (N_46634,N_44719,N_44226);
nor U46635 (N_46635,N_44579,N_44441);
nand U46636 (N_46636,N_44776,N_43252);
nand U46637 (N_46637,N_42800,N_44898);
nand U46638 (N_46638,N_43894,N_43330);
nor U46639 (N_46639,N_43687,N_44118);
or U46640 (N_46640,N_44591,N_43109);
or U46641 (N_46641,N_43337,N_44004);
or U46642 (N_46642,N_44107,N_44428);
and U46643 (N_46643,N_43619,N_43850);
nand U46644 (N_46644,N_43497,N_43543);
and U46645 (N_46645,N_43721,N_42882);
nor U46646 (N_46646,N_43482,N_42583);
or U46647 (N_46647,N_43342,N_43102);
nand U46648 (N_46648,N_42553,N_44056);
nand U46649 (N_46649,N_43053,N_44595);
nand U46650 (N_46650,N_44176,N_43622);
and U46651 (N_46651,N_43407,N_44677);
nor U46652 (N_46652,N_44328,N_43736);
and U46653 (N_46653,N_44784,N_43716);
and U46654 (N_46654,N_43728,N_44654);
and U46655 (N_46655,N_43235,N_44437);
nor U46656 (N_46656,N_44029,N_42601);
and U46657 (N_46657,N_44087,N_43092);
nor U46658 (N_46658,N_43962,N_43868);
nand U46659 (N_46659,N_44685,N_42889);
or U46660 (N_46660,N_43859,N_44455);
nor U46661 (N_46661,N_42648,N_44028);
nor U46662 (N_46662,N_44188,N_42801);
nand U46663 (N_46663,N_42778,N_43565);
nand U46664 (N_46664,N_42524,N_42510);
nand U46665 (N_46665,N_43526,N_43653);
nor U46666 (N_46666,N_43434,N_44653);
and U46667 (N_46667,N_43904,N_43670);
or U46668 (N_46668,N_43321,N_44081);
nor U46669 (N_46669,N_42549,N_44128);
and U46670 (N_46670,N_44351,N_43056);
nor U46671 (N_46671,N_44742,N_42743);
nand U46672 (N_46672,N_43322,N_43496);
and U46673 (N_46673,N_44230,N_44600);
nand U46674 (N_46674,N_43175,N_44586);
nand U46675 (N_46675,N_44669,N_42784);
nand U46676 (N_46676,N_42970,N_42846);
nand U46677 (N_46677,N_44607,N_43397);
and U46678 (N_46678,N_44976,N_44511);
nand U46679 (N_46679,N_44713,N_43578);
or U46680 (N_46680,N_43326,N_44112);
and U46681 (N_46681,N_44383,N_42535);
or U46682 (N_46682,N_42891,N_44685);
xor U46683 (N_46683,N_42883,N_44361);
or U46684 (N_46684,N_43037,N_44520);
or U46685 (N_46685,N_44342,N_44085);
nor U46686 (N_46686,N_43072,N_44483);
nor U46687 (N_46687,N_42572,N_43335);
nand U46688 (N_46688,N_42969,N_43034);
nor U46689 (N_46689,N_44405,N_44978);
xor U46690 (N_46690,N_43254,N_42860);
or U46691 (N_46691,N_43606,N_43445);
or U46692 (N_46692,N_44129,N_43193);
nor U46693 (N_46693,N_42521,N_44725);
nor U46694 (N_46694,N_42861,N_42836);
or U46695 (N_46695,N_44698,N_43542);
and U46696 (N_46696,N_44630,N_44103);
nor U46697 (N_46697,N_44141,N_44089);
nor U46698 (N_46698,N_44807,N_42953);
nand U46699 (N_46699,N_42882,N_42806);
and U46700 (N_46700,N_43930,N_43016);
nor U46701 (N_46701,N_44951,N_42970);
nand U46702 (N_46702,N_44797,N_42866);
and U46703 (N_46703,N_44854,N_42992);
nand U46704 (N_46704,N_44584,N_43632);
nand U46705 (N_46705,N_43710,N_44932);
nor U46706 (N_46706,N_43243,N_44511);
nor U46707 (N_46707,N_43863,N_43540);
and U46708 (N_46708,N_42709,N_43584);
nand U46709 (N_46709,N_44634,N_43392);
nand U46710 (N_46710,N_44093,N_43536);
xnor U46711 (N_46711,N_43100,N_42746);
nand U46712 (N_46712,N_43434,N_43955);
and U46713 (N_46713,N_42995,N_44121);
and U46714 (N_46714,N_44955,N_42789);
and U46715 (N_46715,N_44732,N_44737);
nor U46716 (N_46716,N_43128,N_42584);
nand U46717 (N_46717,N_44682,N_44560);
nand U46718 (N_46718,N_43152,N_42653);
or U46719 (N_46719,N_43610,N_44415);
and U46720 (N_46720,N_44329,N_44449);
xnor U46721 (N_46721,N_44075,N_44717);
or U46722 (N_46722,N_43426,N_43693);
or U46723 (N_46723,N_44114,N_44061);
and U46724 (N_46724,N_42948,N_44772);
nor U46725 (N_46725,N_44077,N_44214);
nor U46726 (N_46726,N_42611,N_42615);
or U46727 (N_46727,N_44437,N_43190);
and U46728 (N_46728,N_44341,N_44935);
or U46729 (N_46729,N_43511,N_43559);
nand U46730 (N_46730,N_42622,N_44154);
and U46731 (N_46731,N_43642,N_42988);
nand U46732 (N_46732,N_42669,N_43110);
nand U46733 (N_46733,N_44160,N_43943);
or U46734 (N_46734,N_44330,N_42829);
and U46735 (N_46735,N_43214,N_43303);
xnor U46736 (N_46736,N_42781,N_42559);
nand U46737 (N_46737,N_43608,N_44393);
or U46738 (N_46738,N_44716,N_42834);
nor U46739 (N_46739,N_42502,N_43819);
nand U46740 (N_46740,N_44019,N_43895);
or U46741 (N_46741,N_43917,N_42960);
nand U46742 (N_46742,N_43428,N_43618);
nor U46743 (N_46743,N_43000,N_43194);
or U46744 (N_46744,N_44177,N_43319);
and U46745 (N_46745,N_42905,N_44730);
and U46746 (N_46746,N_44243,N_44257);
and U46747 (N_46747,N_44092,N_44049);
nor U46748 (N_46748,N_42527,N_44257);
and U46749 (N_46749,N_43574,N_43304);
xor U46750 (N_46750,N_42840,N_43910);
and U46751 (N_46751,N_43377,N_42561);
nand U46752 (N_46752,N_42874,N_43247);
nand U46753 (N_46753,N_44162,N_44351);
nand U46754 (N_46754,N_44099,N_44447);
xnor U46755 (N_46755,N_43113,N_44788);
or U46756 (N_46756,N_43729,N_43724);
or U46757 (N_46757,N_44653,N_42992);
nor U46758 (N_46758,N_42860,N_42924);
nand U46759 (N_46759,N_44482,N_44412);
nor U46760 (N_46760,N_42643,N_44746);
nor U46761 (N_46761,N_44570,N_43655);
nand U46762 (N_46762,N_42976,N_43467);
or U46763 (N_46763,N_44117,N_42678);
nor U46764 (N_46764,N_44782,N_43287);
or U46765 (N_46765,N_42737,N_43102);
xnor U46766 (N_46766,N_44726,N_43860);
nand U46767 (N_46767,N_43675,N_44106);
or U46768 (N_46768,N_43011,N_44697);
nor U46769 (N_46769,N_43812,N_42522);
nand U46770 (N_46770,N_44808,N_44009);
or U46771 (N_46771,N_44325,N_44391);
nor U46772 (N_46772,N_43210,N_43376);
nand U46773 (N_46773,N_42502,N_44160);
and U46774 (N_46774,N_44568,N_42812);
nor U46775 (N_46775,N_42832,N_43707);
nand U46776 (N_46776,N_42905,N_43997);
or U46777 (N_46777,N_43104,N_43807);
nand U46778 (N_46778,N_42552,N_42666);
nor U46779 (N_46779,N_43532,N_43953);
or U46780 (N_46780,N_42798,N_43704);
nand U46781 (N_46781,N_43051,N_44358);
nor U46782 (N_46782,N_44651,N_42515);
nor U46783 (N_46783,N_44458,N_43882);
or U46784 (N_46784,N_43902,N_43403);
nor U46785 (N_46785,N_43159,N_44832);
and U46786 (N_46786,N_42577,N_43229);
or U46787 (N_46787,N_44581,N_44863);
nand U46788 (N_46788,N_43388,N_42631);
and U46789 (N_46789,N_43424,N_43849);
xnor U46790 (N_46790,N_44083,N_44553);
nor U46791 (N_46791,N_44772,N_44511);
or U46792 (N_46792,N_44784,N_44240);
or U46793 (N_46793,N_43477,N_44674);
or U46794 (N_46794,N_43362,N_43454);
or U46795 (N_46795,N_44583,N_42717);
nand U46796 (N_46796,N_43125,N_44696);
nor U46797 (N_46797,N_44082,N_44962);
nor U46798 (N_46798,N_42929,N_42980);
and U46799 (N_46799,N_43321,N_43969);
xor U46800 (N_46800,N_43223,N_44058);
or U46801 (N_46801,N_43507,N_42687);
or U46802 (N_46802,N_44646,N_43173);
or U46803 (N_46803,N_44425,N_43249);
nor U46804 (N_46804,N_44736,N_44694);
nand U46805 (N_46805,N_43044,N_44755);
and U46806 (N_46806,N_43689,N_43163);
or U46807 (N_46807,N_44688,N_43560);
nand U46808 (N_46808,N_44359,N_43188);
xnor U46809 (N_46809,N_44011,N_43014);
and U46810 (N_46810,N_43365,N_43958);
nand U46811 (N_46811,N_44993,N_44690);
nor U46812 (N_46812,N_43118,N_43680);
or U46813 (N_46813,N_44479,N_43178);
nand U46814 (N_46814,N_44965,N_43866);
or U46815 (N_46815,N_43812,N_44315);
xnor U46816 (N_46816,N_43556,N_43135);
xnor U46817 (N_46817,N_43691,N_42924);
or U46818 (N_46818,N_44654,N_42577);
and U46819 (N_46819,N_42702,N_43580);
or U46820 (N_46820,N_44764,N_44976);
and U46821 (N_46821,N_44096,N_42977);
nand U46822 (N_46822,N_42992,N_44359);
nor U46823 (N_46823,N_42689,N_42788);
and U46824 (N_46824,N_42951,N_43814);
or U46825 (N_46825,N_43825,N_42542);
nor U46826 (N_46826,N_44064,N_44916);
nand U46827 (N_46827,N_44887,N_44064);
nor U46828 (N_46828,N_44538,N_43763);
and U46829 (N_46829,N_43202,N_44989);
nand U46830 (N_46830,N_43045,N_44128);
xor U46831 (N_46831,N_43103,N_44210);
or U46832 (N_46832,N_44103,N_44237);
and U46833 (N_46833,N_44119,N_42816);
nand U46834 (N_46834,N_43554,N_44683);
nor U46835 (N_46835,N_44562,N_44883);
xnor U46836 (N_46836,N_43781,N_44521);
nor U46837 (N_46837,N_42578,N_44794);
nand U46838 (N_46838,N_43902,N_42951);
nand U46839 (N_46839,N_44522,N_42956);
and U46840 (N_46840,N_44671,N_42545);
nor U46841 (N_46841,N_44727,N_42598);
nand U46842 (N_46842,N_42845,N_42531);
nand U46843 (N_46843,N_42926,N_44229);
or U46844 (N_46844,N_42521,N_44380);
nor U46845 (N_46845,N_44244,N_43941);
and U46846 (N_46846,N_43749,N_44057);
nor U46847 (N_46847,N_44751,N_44431);
or U46848 (N_46848,N_43440,N_44074);
and U46849 (N_46849,N_43194,N_44679);
and U46850 (N_46850,N_44786,N_44945);
nor U46851 (N_46851,N_43428,N_44223);
or U46852 (N_46852,N_44710,N_43678);
xor U46853 (N_46853,N_43336,N_44666);
nor U46854 (N_46854,N_43514,N_43826);
nor U46855 (N_46855,N_43462,N_44221);
nand U46856 (N_46856,N_44762,N_44627);
nor U46857 (N_46857,N_44165,N_43256);
or U46858 (N_46858,N_42931,N_44022);
or U46859 (N_46859,N_44731,N_44571);
or U46860 (N_46860,N_43714,N_44724);
or U46861 (N_46861,N_42548,N_42651);
nor U46862 (N_46862,N_43866,N_44311);
nor U46863 (N_46863,N_44370,N_44300);
nand U46864 (N_46864,N_43938,N_43675);
and U46865 (N_46865,N_42597,N_42768);
nand U46866 (N_46866,N_43919,N_44843);
or U46867 (N_46867,N_44994,N_43497);
nor U46868 (N_46868,N_43793,N_44640);
nand U46869 (N_46869,N_43565,N_43758);
nand U46870 (N_46870,N_44376,N_42598);
or U46871 (N_46871,N_43105,N_43586);
xor U46872 (N_46872,N_44429,N_44680);
xnor U46873 (N_46873,N_42945,N_44283);
and U46874 (N_46874,N_42688,N_42761);
or U46875 (N_46875,N_42666,N_44240);
and U46876 (N_46876,N_43859,N_44647);
nor U46877 (N_46877,N_44478,N_44517);
and U46878 (N_46878,N_43790,N_43230);
and U46879 (N_46879,N_44799,N_42581);
and U46880 (N_46880,N_42598,N_44217);
nor U46881 (N_46881,N_43140,N_42594);
nor U46882 (N_46882,N_43319,N_43704);
or U46883 (N_46883,N_43059,N_43691);
and U46884 (N_46884,N_43599,N_44729);
nor U46885 (N_46885,N_44991,N_43893);
and U46886 (N_46886,N_44488,N_43204);
nor U46887 (N_46887,N_44628,N_44203);
xor U46888 (N_46888,N_44557,N_42693);
and U46889 (N_46889,N_44534,N_43973);
and U46890 (N_46890,N_43976,N_43119);
nand U46891 (N_46891,N_44303,N_42857);
or U46892 (N_46892,N_43706,N_43026);
xor U46893 (N_46893,N_44039,N_44603);
and U46894 (N_46894,N_44674,N_43165);
nor U46895 (N_46895,N_43092,N_44336);
nand U46896 (N_46896,N_44950,N_44249);
xnor U46897 (N_46897,N_42580,N_43880);
or U46898 (N_46898,N_44461,N_44577);
or U46899 (N_46899,N_42709,N_44707);
or U46900 (N_46900,N_44395,N_44151);
xnor U46901 (N_46901,N_44659,N_44006);
or U46902 (N_46902,N_43036,N_42785);
nand U46903 (N_46903,N_42590,N_43505);
or U46904 (N_46904,N_42945,N_44827);
and U46905 (N_46905,N_44661,N_44293);
nor U46906 (N_46906,N_43394,N_44444);
and U46907 (N_46907,N_44887,N_43522);
or U46908 (N_46908,N_44136,N_42928);
nor U46909 (N_46909,N_43061,N_43023);
nand U46910 (N_46910,N_44277,N_42879);
xnor U46911 (N_46911,N_43975,N_42681);
xor U46912 (N_46912,N_44890,N_42908);
or U46913 (N_46913,N_44830,N_43708);
or U46914 (N_46914,N_44748,N_43461);
nor U46915 (N_46915,N_42971,N_42635);
or U46916 (N_46916,N_42880,N_44190);
xnor U46917 (N_46917,N_44321,N_44658);
or U46918 (N_46918,N_44849,N_43007);
nor U46919 (N_46919,N_42844,N_43079);
and U46920 (N_46920,N_44804,N_43089);
or U46921 (N_46921,N_42589,N_43898);
and U46922 (N_46922,N_43843,N_44624);
nor U46923 (N_46923,N_44137,N_43558);
or U46924 (N_46924,N_44624,N_43278);
nor U46925 (N_46925,N_43650,N_44453);
nor U46926 (N_46926,N_44819,N_44513);
and U46927 (N_46927,N_42982,N_43935);
nand U46928 (N_46928,N_42557,N_42514);
and U46929 (N_46929,N_43175,N_42586);
or U46930 (N_46930,N_44206,N_43638);
nand U46931 (N_46931,N_43777,N_43593);
and U46932 (N_46932,N_44904,N_44058);
and U46933 (N_46933,N_42882,N_43412);
and U46934 (N_46934,N_44157,N_43797);
xnor U46935 (N_46935,N_43097,N_44408);
nand U46936 (N_46936,N_43125,N_43319);
nand U46937 (N_46937,N_43359,N_42696);
and U46938 (N_46938,N_43124,N_44709);
or U46939 (N_46939,N_42848,N_43895);
or U46940 (N_46940,N_44402,N_42570);
xor U46941 (N_46941,N_43151,N_42649);
nand U46942 (N_46942,N_43859,N_43428);
and U46943 (N_46943,N_42713,N_44487);
or U46944 (N_46944,N_43271,N_43603);
or U46945 (N_46945,N_43299,N_44618);
nor U46946 (N_46946,N_44990,N_44616);
and U46947 (N_46947,N_44527,N_43989);
and U46948 (N_46948,N_43339,N_44722);
and U46949 (N_46949,N_43107,N_44479);
nor U46950 (N_46950,N_44121,N_44571);
and U46951 (N_46951,N_44295,N_43025);
or U46952 (N_46952,N_44454,N_44159);
nor U46953 (N_46953,N_43047,N_44001);
nor U46954 (N_46954,N_44438,N_44560);
and U46955 (N_46955,N_43485,N_43467);
nor U46956 (N_46956,N_42666,N_44002);
nor U46957 (N_46957,N_43879,N_44172);
nor U46958 (N_46958,N_44457,N_44003);
nor U46959 (N_46959,N_43017,N_44228);
or U46960 (N_46960,N_42954,N_44451);
nor U46961 (N_46961,N_44552,N_44520);
nand U46962 (N_46962,N_43409,N_42981);
and U46963 (N_46963,N_44431,N_42517);
nand U46964 (N_46964,N_44886,N_44119);
nand U46965 (N_46965,N_42630,N_43747);
nand U46966 (N_46966,N_43644,N_43237);
nor U46967 (N_46967,N_43133,N_44999);
nand U46968 (N_46968,N_44208,N_42752);
and U46969 (N_46969,N_43998,N_44843);
or U46970 (N_46970,N_44295,N_44017);
or U46971 (N_46971,N_42639,N_42812);
and U46972 (N_46972,N_44576,N_44569);
nor U46973 (N_46973,N_44379,N_44585);
or U46974 (N_46974,N_43633,N_43104);
nor U46975 (N_46975,N_43374,N_44158);
or U46976 (N_46976,N_43094,N_43521);
nand U46977 (N_46977,N_43575,N_43085);
nand U46978 (N_46978,N_44829,N_44367);
nand U46979 (N_46979,N_42722,N_44084);
nand U46980 (N_46980,N_43827,N_44022);
or U46981 (N_46981,N_44407,N_44283);
nor U46982 (N_46982,N_44997,N_44066);
or U46983 (N_46983,N_43990,N_42744);
nand U46984 (N_46984,N_44704,N_42961);
and U46985 (N_46985,N_44765,N_44675);
nor U46986 (N_46986,N_43120,N_43728);
or U46987 (N_46987,N_43879,N_43872);
and U46988 (N_46988,N_44988,N_44632);
and U46989 (N_46989,N_44596,N_42951);
nand U46990 (N_46990,N_44571,N_42763);
and U46991 (N_46991,N_44334,N_43929);
nor U46992 (N_46992,N_43545,N_42662);
or U46993 (N_46993,N_42802,N_44237);
and U46994 (N_46994,N_44288,N_44848);
nand U46995 (N_46995,N_42819,N_44031);
and U46996 (N_46996,N_43896,N_44419);
xor U46997 (N_46997,N_44761,N_43285);
or U46998 (N_46998,N_44031,N_42754);
nor U46999 (N_46999,N_43415,N_43896);
nor U47000 (N_47000,N_42969,N_43279);
nand U47001 (N_47001,N_42690,N_43023);
and U47002 (N_47002,N_44862,N_43985);
and U47003 (N_47003,N_44234,N_44527);
xnor U47004 (N_47004,N_44117,N_44925);
or U47005 (N_47005,N_44970,N_43371);
nand U47006 (N_47006,N_42767,N_44770);
nand U47007 (N_47007,N_43031,N_42840);
and U47008 (N_47008,N_44206,N_44672);
and U47009 (N_47009,N_44655,N_44907);
and U47010 (N_47010,N_43031,N_44340);
or U47011 (N_47011,N_43363,N_42966);
and U47012 (N_47012,N_42521,N_44641);
xor U47013 (N_47013,N_43107,N_43240);
and U47014 (N_47014,N_43312,N_43486);
nand U47015 (N_47015,N_43698,N_44079);
and U47016 (N_47016,N_44549,N_44379);
or U47017 (N_47017,N_43501,N_44671);
nor U47018 (N_47018,N_43532,N_43470);
nand U47019 (N_47019,N_43759,N_44818);
or U47020 (N_47020,N_43467,N_44118);
or U47021 (N_47021,N_43368,N_42944);
nor U47022 (N_47022,N_43193,N_43834);
or U47023 (N_47023,N_44721,N_44710);
nor U47024 (N_47024,N_44998,N_43019);
nor U47025 (N_47025,N_43666,N_44214);
and U47026 (N_47026,N_44408,N_43680);
or U47027 (N_47027,N_44700,N_43894);
or U47028 (N_47028,N_44216,N_42754);
nor U47029 (N_47029,N_43781,N_44888);
xnor U47030 (N_47030,N_42566,N_43119);
or U47031 (N_47031,N_44126,N_44737);
xnor U47032 (N_47032,N_44344,N_43139);
and U47033 (N_47033,N_43037,N_43135);
and U47034 (N_47034,N_43462,N_44393);
or U47035 (N_47035,N_43679,N_44883);
xor U47036 (N_47036,N_43026,N_42639);
and U47037 (N_47037,N_43479,N_43008);
or U47038 (N_47038,N_44681,N_44058);
and U47039 (N_47039,N_44575,N_42781);
xor U47040 (N_47040,N_43885,N_44078);
xnor U47041 (N_47041,N_43218,N_44240);
or U47042 (N_47042,N_43300,N_42689);
xor U47043 (N_47043,N_43187,N_43433);
nor U47044 (N_47044,N_42506,N_44213);
xnor U47045 (N_47045,N_44802,N_44078);
xor U47046 (N_47046,N_42719,N_44953);
nor U47047 (N_47047,N_44483,N_43805);
xnor U47048 (N_47048,N_43882,N_43126);
or U47049 (N_47049,N_43489,N_44924);
xnor U47050 (N_47050,N_44656,N_44598);
xnor U47051 (N_47051,N_43686,N_43627);
nand U47052 (N_47052,N_44243,N_44882);
or U47053 (N_47053,N_44268,N_43345);
or U47054 (N_47054,N_43006,N_44709);
and U47055 (N_47055,N_43945,N_44901);
xor U47056 (N_47056,N_43018,N_43446);
or U47057 (N_47057,N_44812,N_43894);
or U47058 (N_47058,N_43271,N_42761);
and U47059 (N_47059,N_44869,N_44200);
nand U47060 (N_47060,N_43753,N_43781);
nand U47061 (N_47061,N_43188,N_44161);
nor U47062 (N_47062,N_43057,N_43625);
nand U47063 (N_47063,N_43853,N_43882);
and U47064 (N_47064,N_43048,N_42949);
nor U47065 (N_47065,N_43531,N_44532);
and U47066 (N_47066,N_44519,N_44898);
xnor U47067 (N_47067,N_43801,N_44895);
and U47068 (N_47068,N_44289,N_43187);
xnor U47069 (N_47069,N_44070,N_43170);
xor U47070 (N_47070,N_44115,N_42535);
or U47071 (N_47071,N_44659,N_43992);
or U47072 (N_47072,N_44798,N_43465);
nor U47073 (N_47073,N_43791,N_44997);
and U47074 (N_47074,N_44452,N_44119);
nand U47075 (N_47075,N_43830,N_43206);
or U47076 (N_47076,N_44212,N_43609);
nor U47077 (N_47077,N_44626,N_42677);
xnor U47078 (N_47078,N_43939,N_43259);
xnor U47079 (N_47079,N_43064,N_43032);
or U47080 (N_47080,N_43795,N_44062);
nand U47081 (N_47081,N_44656,N_43543);
nor U47082 (N_47082,N_44960,N_42827);
and U47083 (N_47083,N_43695,N_44420);
xnor U47084 (N_47084,N_43675,N_43168);
nor U47085 (N_47085,N_44975,N_43640);
and U47086 (N_47086,N_44989,N_43858);
or U47087 (N_47087,N_44253,N_44073);
nand U47088 (N_47088,N_44687,N_43485);
or U47089 (N_47089,N_43202,N_44325);
or U47090 (N_47090,N_42923,N_42624);
nand U47091 (N_47091,N_42861,N_44571);
nor U47092 (N_47092,N_44727,N_43121);
nand U47093 (N_47093,N_42585,N_44477);
and U47094 (N_47094,N_44857,N_43463);
nand U47095 (N_47095,N_42864,N_44785);
nand U47096 (N_47096,N_42501,N_44717);
nor U47097 (N_47097,N_44116,N_44479);
nor U47098 (N_47098,N_43961,N_42670);
and U47099 (N_47099,N_43798,N_42740);
or U47100 (N_47100,N_44613,N_44825);
and U47101 (N_47101,N_42512,N_43273);
nand U47102 (N_47102,N_43663,N_42741);
or U47103 (N_47103,N_44804,N_43169);
nand U47104 (N_47104,N_44416,N_43159);
and U47105 (N_47105,N_44307,N_44853);
nand U47106 (N_47106,N_44188,N_44996);
nand U47107 (N_47107,N_42541,N_42721);
xor U47108 (N_47108,N_44538,N_43947);
or U47109 (N_47109,N_43277,N_44157);
nand U47110 (N_47110,N_43745,N_44895);
and U47111 (N_47111,N_44901,N_44898);
xnor U47112 (N_47112,N_43080,N_44705);
nor U47113 (N_47113,N_43032,N_42931);
and U47114 (N_47114,N_44942,N_42975);
and U47115 (N_47115,N_44219,N_43034);
or U47116 (N_47116,N_44094,N_43154);
nor U47117 (N_47117,N_44564,N_44570);
and U47118 (N_47118,N_43787,N_42733);
nor U47119 (N_47119,N_43350,N_42532);
and U47120 (N_47120,N_43197,N_43705);
nand U47121 (N_47121,N_44904,N_43509);
or U47122 (N_47122,N_43134,N_43898);
and U47123 (N_47123,N_43432,N_43389);
nor U47124 (N_47124,N_42577,N_44728);
nor U47125 (N_47125,N_43039,N_43967);
nor U47126 (N_47126,N_43687,N_44946);
and U47127 (N_47127,N_44604,N_42849);
nand U47128 (N_47128,N_43434,N_43661);
or U47129 (N_47129,N_43376,N_43641);
nor U47130 (N_47130,N_43079,N_44630);
nand U47131 (N_47131,N_44555,N_44893);
or U47132 (N_47132,N_43020,N_43686);
nand U47133 (N_47133,N_44929,N_43629);
or U47134 (N_47134,N_44031,N_43865);
nor U47135 (N_47135,N_43155,N_44884);
or U47136 (N_47136,N_44182,N_43361);
or U47137 (N_47137,N_43008,N_44353);
or U47138 (N_47138,N_43840,N_43661);
nand U47139 (N_47139,N_42596,N_44586);
nor U47140 (N_47140,N_44768,N_42765);
nand U47141 (N_47141,N_43836,N_43819);
xor U47142 (N_47142,N_44720,N_44717);
nor U47143 (N_47143,N_42978,N_43176);
and U47144 (N_47144,N_43549,N_43024);
or U47145 (N_47145,N_44824,N_44685);
nand U47146 (N_47146,N_44075,N_44356);
or U47147 (N_47147,N_42581,N_43421);
or U47148 (N_47148,N_42794,N_43367);
nor U47149 (N_47149,N_43040,N_42638);
nor U47150 (N_47150,N_42568,N_42555);
and U47151 (N_47151,N_44958,N_44813);
and U47152 (N_47152,N_43996,N_44633);
and U47153 (N_47153,N_43510,N_43896);
and U47154 (N_47154,N_44257,N_42604);
and U47155 (N_47155,N_43431,N_43028);
xor U47156 (N_47156,N_42656,N_43586);
nand U47157 (N_47157,N_43431,N_42935);
xnor U47158 (N_47158,N_43651,N_44487);
nand U47159 (N_47159,N_43403,N_43490);
and U47160 (N_47160,N_43404,N_44872);
or U47161 (N_47161,N_43466,N_44183);
nand U47162 (N_47162,N_44898,N_44293);
or U47163 (N_47163,N_43693,N_44429);
nor U47164 (N_47164,N_43334,N_42606);
or U47165 (N_47165,N_43684,N_43196);
nor U47166 (N_47166,N_44833,N_44497);
or U47167 (N_47167,N_42616,N_43217);
nor U47168 (N_47168,N_43964,N_42715);
xor U47169 (N_47169,N_43911,N_44987);
nor U47170 (N_47170,N_43698,N_44719);
or U47171 (N_47171,N_43674,N_44987);
nor U47172 (N_47172,N_42804,N_43912);
nand U47173 (N_47173,N_43869,N_42625);
xor U47174 (N_47174,N_43943,N_43254);
and U47175 (N_47175,N_43675,N_42516);
or U47176 (N_47176,N_43706,N_43303);
nand U47177 (N_47177,N_42965,N_43997);
or U47178 (N_47178,N_43479,N_42995);
or U47179 (N_47179,N_43307,N_42837);
and U47180 (N_47180,N_43623,N_42650);
or U47181 (N_47181,N_44056,N_43294);
nor U47182 (N_47182,N_44447,N_44278);
or U47183 (N_47183,N_44486,N_44408);
and U47184 (N_47184,N_43549,N_43081);
nor U47185 (N_47185,N_42728,N_42558);
and U47186 (N_47186,N_43970,N_43987);
nand U47187 (N_47187,N_42908,N_44715);
and U47188 (N_47188,N_43904,N_42800);
or U47189 (N_47189,N_43873,N_44937);
and U47190 (N_47190,N_43359,N_43017);
nand U47191 (N_47191,N_43287,N_42559);
nor U47192 (N_47192,N_44231,N_44478);
and U47193 (N_47193,N_43773,N_44876);
nand U47194 (N_47194,N_43878,N_42787);
or U47195 (N_47195,N_42964,N_44354);
nand U47196 (N_47196,N_43541,N_42675);
or U47197 (N_47197,N_42856,N_43409);
or U47198 (N_47198,N_44844,N_44387);
nand U47199 (N_47199,N_44198,N_43908);
and U47200 (N_47200,N_44774,N_42951);
and U47201 (N_47201,N_43121,N_44733);
nand U47202 (N_47202,N_44932,N_43469);
or U47203 (N_47203,N_43326,N_44537);
and U47204 (N_47204,N_44343,N_44620);
or U47205 (N_47205,N_44673,N_44990);
nand U47206 (N_47206,N_43577,N_44781);
or U47207 (N_47207,N_44549,N_42747);
nor U47208 (N_47208,N_43841,N_43638);
nand U47209 (N_47209,N_42596,N_42658);
nand U47210 (N_47210,N_44111,N_42980);
nor U47211 (N_47211,N_42532,N_44776);
xor U47212 (N_47212,N_43615,N_43048);
nor U47213 (N_47213,N_43453,N_43907);
nand U47214 (N_47214,N_44056,N_43236);
or U47215 (N_47215,N_42611,N_42738);
nand U47216 (N_47216,N_43049,N_42959);
and U47217 (N_47217,N_43663,N_43475);
nand U47218 (N_47218,N_44429,N_44775);
nand U47219 (N_47219,N_42592,N_43959);
nand U47220 (N_47220,N_43668,N_43786);
and U47221 (N_47221,N_44776,N_42785);
or U47222 (N_47222,N_44340,N_42976);
nor U47223 (N_47223,N_43152,N_44578);
and U47224 (N_47224,N_44566,N_44825);
or U47225 (N_47225,N_43776,N_42869);
xor U47226 (N_47226,N_43460,N_43649);
nand U47227 (N_47227,N_43467,N_42555);
or U47228 (N_47228,N_44400,N_44483);
or U47229 (N_47229,N_42853,N_42911);
nor U47230 (N_47230,N_43403,N_42645);
nand U47231 (N_47231,N_44636,N_44032);
and U47232 (N_47232,N_42692,N_44599);
nand U47233 (N_47233,N_44533,N_43148);
or U47234 (N_47234,N_42679,N_43249);
or U47235 (N_47235,N_44598,N_43310);
and U47236 (N_47236,N_44103,N_43528);
and U47237 (N_47237,N_44064,N_43733);
and U47238 (N_47238,N_44620,N_43859);
nor U47239 (N_47239,N_44176,N_42843);
nor U47240 (N_47240,N_43452,N_43468);
and U47241 (N_47241,N_43148,N_42932);
and U47242 (N_47242,N_44319,N_42592);
or U47243 (N_47243,N_42932,N_43147);
or U47244 (N_47244,N_44477,N_44816);
nor U47245 (N_47245,N_44605,N_43392);
nor U47246 (N_47246,N_44138,N_42699);
nor U47247 (N_47247,N_43291,N_43155);
nand U47248 (N_47248,N_43359,N_44893);
or U47249 (N_47249,N_43384,N_44363);
nor U47250 (N_47250,N_43945,N_43133);
or U47251 (N_47251,N_43678,N_44492);
nand U47252 (N_47252,N_42644,N_43508);
or U47253 (N_47253,N_43486,N_42552);
or U47254 (N_47254,N_44191,N_44017);
xor U47255 (N_47255,N_44816,N_44206);
or U47256 (N_47256,N_43928,N_43261);
nor U47257 (N_47257,N_42699,N_43936);
and U47258 (N_47258,N_44604,N_43953);
or U47259 (N_47259,N_44501,N_44141);
or U47260 (N_47260,N_43656,N_43003);
nand U47261 (N_47261,N_44322,N_42753);
nor U47262 (N_47262,N_42627,N_42760);
xor U47263 (N_47263,N_43554,N_44250);
and U47264 (N_47264,N_44160,N_43668);
or U47265 (N_47265,N_42705,N_44734);
or U47266 (N_47266,N_44937,N_43272);
xnor U47267 (N_47267,N_44097,N_44315);
and U47268 (N_47268,N_43599,N_43453);
or U47269 (N_47269,N_44715,N_44737);
and U47270 (N_47270,N_43065,N_44342);
nor U47271 (N_47271,N_42857,N_42576);
nand U47272 (N_47272,N_43265,N_43508);
nor U47273 (N_47273,N_43195,N_44685);
nor U47274 (N_47274,N_43013,N_43821);
or U47275 (N_47275,N_43583,N_43703);
nor U47276 (N_47276,N_44170,N_43370);
or U47277 (N_47277,N_44374,N_42887);
nor U47278 (N_47278,N_43459,N_43496);
nand U47279 (N_47279,N_44322,N_44603);
nor U47280 (N_47280,N_43954,N_42625);
nand U47281 (N_47281,N_44730,N_44522);
nand U47282 (N_47282,N_43867,N_44303);
nand U47283 (N_47283,N_43714,N_44850);
nand U47284 (N_47284,N_43501,N_42968);
nand U47285 (N_47285,N_44981,N_43856);
nor U47286 (N_47286,N_44607,N_44280);
nand U47287 (N_47287,N_44315,N_44066);
nor U47288 (N_47288,N_42524,N_42681);
nor U47289 (N_47289,N_43646,N_43913);
or U47290 (N_47290,N_42810,N_43486);
nand U47291 (N_47291,N_43952,N_43261);
and U47292 (N_47292,N_42975,N_44122);
or U47293 (N_47293,N_44775,N_44625);
or U47294 (N_47294,N_44963,N_44033);
nand U47295 (N_47295,N_44749,N_43734);
or U47296 (N_47296,N_44459,N_42683);
nor U47297 (N_47297,N_44403,N_43525);
or U47298 (N_47298,N_44904,N_43957);
nor U47299 (N_47299,N_44348,N_44017);
nor U47300 (N_47300,N_43638,N_42632);
and U47301 (N_47301,N_44662,N_42584);
or U47302 (N_47302,N_44976,N_43379);
nor U47303 (N_47303,N_44223,N_42853);
and U47304 (N_47304,N_43120,N_42890);
or U47305 (N_47305,N_44383,N_43799);
nor U47306 (N_47306,N_42961,N_42519);
nand U47307 (N_47307,N_44719,N_43255);
nand U47308 (N_47308,N_43148,N_43842);
or U47309 (N_47309,N_42624,N_43325);
nand U47310 (N_47310,N_44669,N_44929);
and U47311 (N_47311,N_42735,N_43007);
or U47312 (N_47312,N_44649,N_43451);
or U47313 (N_47313,N_42832,N_43729);
or U47314 (N_47314,N_44705,N_44510);
and U47315 (N_47315,N_44884,N_43407);
nand U47316 (N_47316,N_44659,N_42794);
nand U47317 (N_47317,N_44734,N_43143);
and U47318 (N_47318,N_44177,N_43933);
nor U47319 (N_47319,N_43629,N_43850);
and U47320 (N_47320,N_43469,N_44878);
or U47321 (N_47321,N_43404,N_44408);
and U47322 (N_47322,N_44807,N_43015);
or U47323 (N_47323,N_44274,N_43787);
nand U47324 (N_47324,N_43051,N_44917);
nor U47325 (N_47325,N_44877,N_43321);
nand U47326 (N_47326,N_43297,N_43879);
nor U47327 (N_47327,N_43359,N_44001);
or U47328 (N_47328,N_44532,N_44531);
and U47329 (N_47329,N_43277,N_43846);
or U47330 (N_47330,N_42837,N_44537);
and U47331 (N_47331,N_44614,N_44488);
or U47332 (N_47332,N_44412,N_42797);
or U47333 (N_47333,N_44905,N_43128);
xnor U47334 (N_47334,N_42925,N_42585);
or U47335 (N_47335,N_43854,N_43094);
nand U47336 (N_47336,N_44830,N_44565);
and U47337 (N_47337,N_43418,N_44941);
nor U47338 (N_47338,N_44844,N_44198);
and U47339 (N_47339,N_43035,N_44946);
or U47340 (N_47340,N_44998,N_43230);
nand U47341 (N_47341,N_43966,N_44590);
nor U47342 (N_47342,N_44568,N_43245);
nor U47343 (N_47343,N_44021,N_44281);
nor U47344 (N_47344,N_42688,N_43569);
xor U47345 (N_47345,N_42927,N_44095);
nand U47346 (N_47346,N_44090,N_43684);
or U47347 (N_47347,N_44499,N_43915);
and U47348 (N_47348,N_42640,N_43197);
and U47349 (N_47349,N_44014,N_44994);
nor U47350 (N_47350,N_42791,N_43209);
nor U47351 (N_47351,N_43268,N_42898);
nand U47352 (N_47352,N_44518,N_42655);
nor U47353 (N_47353,N_44705,N_43737);
or U47354 (N_47354,N_42816,N_43518);
or U47355 (N_47355,N_44350,N_42827);
nand U47356 (N_47356,N_43337,N_44824);
nand U47357 (N_47357,N_42889,N_43351);
nand U47358 (N_47358,N_44059,N_43401);
and U47359 (N_47359,N_42965,N_44637);
nand U47360 (N_47360,N_43063,N_42899);
nand U47361 (N_47361,N_42670,N_44453);
nand U47362 (N_47362,N_44897,N_43600);
xnor U47363 (N_47363,N_42790,N_44688);
and U47364 (N_47364,N_44298,N_44211);
nor U47365 (N_47365,N_43318,N_43461);
or U47366 (N_47366,N_42858,N_42649);
nand U47367 (N_47367,N_43591,N_44205);
xnor U47368 (N_47368,N_44345,N_44498);
nor U47369 (N_47369,N_43156,N_43469);
nand U47370 (N_47370,N_43270,N_43776);
nand U47371 (N_47371,N_44506,N_44840);
and U47372 (N_47372,N_42805,N_42673);
and U47373 (N_47373,N_42937,N_42921);
nor U47374 (N_47374,N_44344,N_43855);
and U47375 (N_47375,N_43471,N_44036);
or U47376 (N_47376,N_43861,N_43045);
nor U47377 (N_47377,N_44108,N_44341);
and U47378 (N_47378,N_44460,N_43130);
nor U47379 (N_47379,N_42808,N_44269);
nand U47380 (N_47380,N_43416,N_43727);
and U47381 (N_47381,N_42592,N_44032);
nand U47382 (N_47382,N_43635,N_42791);
nand U47383 (N_47383,N_43969,N_42563);
nand U47384 (N_47384,N_43603,N_44017);
and U47385 (N_47385,N_44659,N_43434);
or U47386 (N_47386,N_42948,N_44519);
and U47387 (N_47387,N_42867,N_44680);
or U47388 (N_47388,N_44189,N_42609);
and U47389 (N_47389,N_42832,N_43146);
xnor U47390 (N_47390,N_44449,N_43291);
nor U47391 (N_47391,N_43818,N_44400);
nand U47392 (N_47392,N_42530,N_44820);
or U47393 (N_47393,N_44299,N_43236);
nor U47394 (N_47394,N_44575,N_44010);
xnor U47395 (N_47395,N_43749,N_42979);
and U47396 (N_47396,N_44549,N_44619);
nor U47397 (N_47397,N_44682,N_43317);
or U47398 (N_47398,N_43357,N_44858);
xnor U47399 (N_47399,N_44270,N_44565);
and U47400 (N_47400,N_44993,N_43198);
or U47401 (N_47401,N_44275,N_44300);
nor U47402 (N_47402,N_42669,N_43705);
nand U47403 (N_47403,N_44031,N_44338);
nand U47404 (N_47404,N_43779,N_42629);
and U47405 (N_47405,N_44157,N_43241);
nand U47406 (N_47406,N_43922,N_43635);
nor U47407 (N_47407,N_43044,N_43931);
nand U47408 (N_47408,N_44094,N_44326);
and U47409 (N_47409,N_44466,N_44598);
xnor U47410 (N_47410,N_43378,N_43480);
and U47411 (N_47411,N_44409,N_44964);
xnor U47412 (N_47412,N_43007,N_44836);
nor U47413 (N_47413,N_44619,N_44601);
nor U47414 (N_47414,N_44686,N_42634);
nand U47415 (N_47415,N_43208,N_43456);
and U47416 (N_47416,N_44777,N_43695);
and U47417 (N_47417,N_43324,N_43945);
nor U47418 (N_47418,N_43253,N_42848);
nor U47419 (N_47419,N_44592,N_42560);
nor U47420 (N_47420,N_43715,N_43334);
and U47421 (N_47421,N_43349,N_42920);
nor U47422 (N_47422,N_44589,N_44992);
or U47423 (N_47423,N_43301,N_44043);
nand U47424 (N_47424,N_44116,N_43691);
or U47425 (N_47425,N_44436,N_43598);
nand U47426 (N_47426,N_44707,N_44589);
and U47427 (N_47427,N_44580,N_44912);
or U47428 (N_47428,N_43725,N_44584);
or U47429 (N_47429,N_44473,N_44850);
or U47430 (N_47430,N_43466,N_43567);
nand U47431 (N_47431,N_43156,N_43688);
or U47432 (N_47432,N_42932,N_43313);
or U47433 (N_47433,N_43869,N_43928);
nand U47434 (N_47434,N_42634,N_44593);
and U47435 (N_47435,N_44793,N_44721);
or U47436 (N_47436,N_42717,N_43159);
nor U47437 (N_47437,N_44966,N_44245);
nand U47438 (N_47438,N_42903,N_43785);
nand U47439 (N_47439,N_44400,N_42808);
or U47440 (N_47440,N_42772,N_44000);
or U47441 (N_47441,N_43146,N_43046);
or U47442 (N_47442,N_44190,N_44433);
and U47443 (N_47443,N_44787,N_42925);
and U47444 (N_47444,N_42605,N_44035);
and U47445 (N_47445,N_43313,N_44241);
and U47446 (N_47446,N_44836,N_44793);
and U47447 (N_47447,N_42860,N_44479);
nand U47448 (N_47448,N_42805,N_44762);
and U47449 (N_47449,N_44401,N_42810);
nand U47450 (N_47450,N_43709,N_44128);
or U47451 (N_47451,N_42578,N_43402);
nand U47452 (N_47452,N_43577,N_42612);
nand U47453 (N_47453,N_42946,N_44045);
and U47454 (N_47454,N_44895,N_43449);
nor U47455 (N_47455,N_43354,N_43052);
xnor U47456 (N_47456,N_42892,N_43925);
or U47457 (N_47457,N_42776,N_43155);
or U47458 (N_47458,N_44134,N_44515);
nor U47459 (N_47459,N_44813,N_44436);
nand U47460 (N_47460,N_44349,N_43375);
nor U47461 (N_47461,N_42554,N_43370);
nor U47462 (N_47462,N_43025,N_44144);
nand U47463 (N_47463,N_42993,N_43307);
xnor U47464 (N_47464,N_42639,N_44863);
xnor U47465 (N_47465,N_43480,N_44406);
nor U47466 (N_47466,N_42813,N_44184);
or U47467 (N_47467,N_44984,N_44498);
and U47468 (N_47468,N_44323,N_43237);
nor U47469 (N_47469,N_44611,N_44398);
nor U47470 (N_47470,N_44286,N_42950);
and U47471 (N_47471,N_42923,N_43851);
nor U47472 (N_47472,N_44694,N_43092);
nor U47473 (N_47473,N_43346,N_43460);
nand U47474 (N_47474,N_44995,N_44008);
xor U47475 (N_47475,N_42924,N_44239);
nor U47476 (N_47476,N_43110,N_44610);
nand U47477 (N_47477,N_43671,N_44290);
nand U47478 (N_47478,N_43169,N_44865);
or U47479 (N_47479,N_44069,N_43853);
nor U47480 (N_47480,N_42724,N_43853);
and U47481 (N_47481,N_43290,N_44158);
xor U47482 (N_47482,N_43029,N_44567);
or U47483 (N_47483,N_43857,N_43830);
nor U47484 (N_47484,N_43809,N_43873);
and U47485 (N_47485,N_43820,N_43282);
nand U47486 (N_47486,N_43132,N_43437);
or U47487 (N_47487,N_43076,N_43270);
or U47488 (N_47488,N_43058,N_43759);
nand U47489 (N_47489,N_43748,N_43069);
or U47490 (N_47490,N_43837,N_43169);
or U47491 (N_47491,N_44848,N_44239);
or U47492 (N_47492,N_44284,N_43244);
nor U47493 (N_47493,N_43224,N_43476);
or U47494 (N_47494,N_43900,N_44303);
nor U47495 (N_47495,N_42629,N_43485);
and U47496 (N_47496,N_44890,N_42625);
and U47497 (N_47497,N_44341,N_43464);
nor U47498 (N_47498,N_44418,N_44819);
or U47499 (N_47499,N_42705,N_42890);
nor U47500 (N_47500,N_46386,N_46274);
and U47501 (N_47501,N_45301,N_46894);
or U47502 (N_47502,N_45224,N_46489);
nand U47503 (N_47503,N_46046,N_45805);
and U47504 (N_47504,N_46311,N_46290);
nand U47505 (N_47505,N_45929,N_46586);
xor U47506 (N_47506,N_47304,N_46638);
or U47507 (N_47507,N_46649,N_45330);
xor U47508 (N_47508,N_46261,N_45140);
nand U47509 (N_47509,N_45773,N_45809);
or U47510 (N_47510,N_47113,N_45179);
nand U47511 (N_47511,N_46068,N_47480);
and U47512 (N_47512,N_47327,N_46527);
and U47513 (N_47513,N_45200,N_46307);
or U47514 (N_47514,N_46763,N_46155);
and U47515 (N_47515,N_45437,N_45495);
or U47516 (N_47516,N_46767,N_46828);
nor U47517 (N_47517,N_47175,N_46922);
and U47518 (N_47518,N_45616,N_46500);
and U47519 (N_47519,N_45125,N_46716);
nand U47520 (N_47520,N_45482,N_45552);
nand U47521 (N_47521,N_46560,N_46698);
nor U47522 (N_47522,N_45696,N_47428);
nand U47523 (N_47523,N_47086,N_46644);
nor U47524 (N_47524,N_46991,N_45409);
nand U47525 (N_47525,N_45303,N_45285);
or U47526 (N_47526,N_46504,N_47207);
xor U47527 (N_47527,N_45941,N_46946);
or U47528 (N_47528,N_45629,N_45671);
nor U47529 (N_47529,N_45857,N_45458);
or U47530 (N_47530,N_45561,N_45212);
and U47531 (N_47531,N_46248,N_47394);
nor U47532 (N_47532,N_46324,N_47254);
or U47533 (N_47533,N_45698,N_46471);
nor U47534 (N_47534,N_46252,N_45311);
xor U47535 (N_47535,N_45227,N_46117);
nand U47536 (N_47536,N_47266,N_46985);
or U47537 (N_47537,N_46693,N_46912);
nor U47538 (N_47538,N_47210,N_47465);
xor U47539 (N_47539,N_45606,N_45540);
nand U47540 (N_47540,N_45995,N_45830);
and U47541 (N_47541,N_45583,N_45176);
and U47542 (N_47542,N_45372,N_46004);
or U47543 (N_47543,N_47366,N_46203);
and U47544 (N_47544,N_46401,N_45849);
nand U47545 (N_47545,N_45317,N_45587);
or U47546 (N_47546,N_45868,N_46986);
or U47547 (N_47547,N_45555,N_45204);
nand U47548 (N_47548,N_45232,N_47371);
and U47549 (N_47549,N_46960,N_45911);
or U47550 (N_47550,N_46949,N_46608);
or U47551 (N_47551,N_47132,N_46734);
and U47552 (N_47552,N_46847,N_47059);
or U47553 (N_47553,N_46498,N_46253);
nor U47554 (N_47554,N_45615,N_46583);
xnor U47555 (N_47555,N_45451,N_46839);
nand U47556 (N_47556,N_47191,N_46926);
nor U47557 (N_47557,N_45948,N_46010);
nor U47558 (N_47558,N_46130,N_45072);
or U47559 (N_47559,N_45353,N_45320);
or U47560 (N_47560,N_45890,N_46310);
or U47561 (N_47561,N_45415,N_46435);
and U47562 (N_47562,N_46948,N_46677);
and U47563 (N_47563,N_47375,N_45340);
nand U47564 (N_47564,N_45380,N_46565);
nor U47565 (N_47565,N_46062,N_46387);
nor U47566 (N_47566,N_46708,N_45876);
nand U47567 (N_47567,N_46662,N_46260);
nor U47568 (N_47568,N_45544,N_46488);
or U47569 (N_47569,N_46600,N_47404);
and U47570 (N_47570,N_45605,N_47115);
nand U47571 (N_47571,N_47449,N_46225);
and U47572 (N_47572,N_46496,N_45993);
nor U47573 (N_47573,N_46047,N_46108);
and U47574 (N_47574,N_45617,N_46786);
nand U47575 (N_47575,N_45196,N_46006);
nand U47576 (N_47576,N_45310,N_45503);
and U47577 (N_47577,N_45289,N_45579);
and U47578 (N_47578,N_46595,N_45553);
and U47579 (N_47579,N_45614,N_45266);
nor U47580 (N_47580,N_45115,N_45172);
nand U47581 (N_47581,N_47152,N_45992);
xor U47582 (N_47582,N_47062,N_45272);
and U47583 (N_47583,N_45977,N_47185);
xor U47584 (N_47584,N_46727,N_45135);
or U47585 (N_47585,N_46074,N_46022);
xnor U47586 (N_47586,N_46367,N_46136);
and U47587 (N_47587,N_46128,N_46439);
or U47588 (N_47588,N_46431,N_45680);
and U47589 (N_47589,N_47451,N_47340);
nor U47590 (N_47590,N_46570,N_45591);
or U47591 (N_47591,N_46483,N_45749);
and U47592 (N_47592,N_45776,N_46011);
or U47593 (N_47593,N_45750,N_46625);
or U47594 (N_47594,N_45539,N_46998);
or U47595 (N_47595,N_45257,N_46393);
nand U47596 (N_47596,N_45510,N_45493);
and U47597 (N_47597,N_47299,N_46701);
nor U47598 (N_47598,N_47282,N_45217);
nor U47599 (N_47599,N_45361,N_45377);
nor U47600 (N_47600,N_46040,N_45011);
or U47601 (N_47601,N_45746,N_46294);
or U47602 (N_47602,N_46369,N_46001);
nor U47603 (N_47603,N_46747,N_47239);
nand U47604 (N_47604,N_47060,N_47281);
and U47605 (N_47605,N_45359,N_46574);
or U47606 (N_47606,N_46609,N_47081);
nor U47607 (N_47607,N_47192,N_47017);
nor U47608 (N_47608,N_46569,N_45085);
nand U47609 (N_47609,N_47102,N_46876);
nand U47610 (N_47610,N_45666,N_47047);
and U47611 (N_47611,N_45633,N_45487);
nor U47612 (N_47612,N_45794,N_46521);
nor U47613 (N_47613,N_47163,N_46928);
xnor U47614 (N_47614,N_45413,N_47172);
xor U47615 (N_47615,N_45659,N_45186);
nand U47616 (N_47616,N_46741,N_46419);
and U47617 (N_47617,N_47349,N_45106);
nand U47618 (N_47618,N_47430,N_47140);
and U47619 (N_47619,N_46650,N_45575);
nor U47620 (N_47620,N_45781,N_45252);
xnor U47621 (N_47621,N_47305,N_45267);
nand U47622 (N_47622,N_45263,N_47408);
or U47623 (N_47623,N_46070,N_45494);
nor U47624 (N_47624,N_45567,N_47258);
or U47625 (N_47625,N_46002,N_47274);
xnor U47626 (N_47626,N_46563,N_45527);
nor U47627 (N_47627,N_46883,N_47129);
nor U47628 (N_47628,N_47149,N_45138);
xor U47629 (N_47629,N_46254,N_46648);
and U47630 (N_47630,N_47079,N_45018);
nor U47631 (N_47631,N_46818,N_47231);
and U47632 (N_47632,N_45463,N_45133);
or U47633 (N_47633,N_46209,N_45914);
nand U47634 (N_47634,N_47442,N_46061);
or U47635 (N_47635,N_46557,N_45348);
nor U47636 (N_47636,N_45128,N_46277);
nor U47637 (N_47637,N_45465,N_45275);
xnor U47638 (N_47638,N_46544,N_46666);
nand U47639 (N_47639,N_45080,N_45058);
nand U47640 (N_47640,N_47436,N_47146);
and U47641 (N_47641,N_46451,N_46753);
nor U47642 (N_47642,N_47409,N_46016);
and U47643 (N_47643,N_46766,N_47443);
xor U47644 (N_47644,N_45077,N_46174);
or U47645 (N_47645,N_46639,N_46581);
or U47646 (N_47646,N_45882,N_46663);
nand U47647 (N_47647,N_46917,N_46309);
or U47648 (N_47648,N_45492,N_46759);
nand U47649 (N_47649,N_45293,N_46775);
nor U47650 (N_47650,N_47325,N_45867);
nor U47651 (N_47651,N_45920,N_46669);
and U47652 (N_47652,N_47201,N_46571);
or U47653 (N_47653,N_47460,N_45811);
or U47654 (N_47654,N_46631,N_46866);
nand U47655 (N_47655,N_46090,N_45020);
nand U47656 (N_47656,N_45417,N_45202);
and U47657 (N_47657,N_46925,N_46719);
or U47658 (N_47658,N_45956,N_46792);
nor U47659 (N_47659,N_47314,N_46194);
and U47660 (N_47660,N_45021,N_47380);
or U47661 (N_47661,N_46954,N_45279);
nor U47662 (N_47662,N_45559,N_45824);
nand U47663 (N_47663,N_45812,N_45858);
and U47664 (N_47664,N_45508,N_47177);
or U47665 (N_47665,N_46402,N_47405);
and U47666 (N_47666,N_45925,N_47120);
or U47667 (N_47667,N_47298,N_45016);
nor U47668 (N_47668,N_46086,N_46983);
nor U47669 (N_47669,N_46167,N_45931);
nand U47670 (N_47670,N_45886,N_45382);
nand U47671 (N_47671,N_45171,N_46906);
nand U47672 (N_47672,N_47472,N_47240);
nand U47673 (N_47673,N_46961,N_45156);
and U47674 (N_47674,N_45891,N_47174);
nand U47675 (N_47675,N_46221,N_46163);
or U47676 (N_47676,N_47348,N_46236);
nor U47677 (N_47677,N_45772,N_45370);
or U47678 (N_47678,N_45490,N_46971);
and U47679 (N_47679,N_46973,N_45641);
nand U47680 (N_47680,N_46826,N_45524);
nor U47681 (N_47681,N_46326,N_46320);
nand U47682 (N_47682,N_45446,N_46603);
or U47683 (N_47683,N_46841,N_46457);
nand U47684 (N_47684,N_47256,N_45919);
nor U47685 (N_47685,N_47234,N_47241);
nand U47686 (N_47686,N_45753,N_46606);
or U47687 (N_47687,N_45439,N_45118);
nand U47688 (N_47688,N_45358,N_46328);
nand U47689 (N_47689,N_45519,N_47243);
nand U47690 (N_47690,N_47013,N_46285);
nand U47691 (N_47691,N_46131,N_46023);
nor U47692 (N_47692,N_46063,N_46373);
nor U47693 (N_47693,N_46887,N_46950);
and U47694 (N_47694,N_47401,N_46640);
nor U47695 (N_47695,N_46758,N_47085);
nor U47696 (N_47696,N_46768,N_46699);
or U47697 (N_47697,N_46377,N_46075);
nor U47698 (N_47698,N_46278,N_47233);
nand U47699 (N_47699,N_46684,N_46342);
nor U47700 (N_47700,N_45057,N_45662);
and U47701 (N_47701,N_46079,N_46980);
xor U47702 (N_47702,N_45197,N_45445);
and U47703 (N_47703,N_45190,N_46143);
nor U47704 (N_47704,N_45274,N_45014);
nor U47705 (N_47705,N_47490,N_45747);
xnor U47706 (N_47706,N_45306,N_45379);
or U47707 (N_47707,N_46739,N_46239);
nand U47708 (N_47708,N_46987,N_46233);
or U47709 (N_47709,N_45887,N_45702);
nor U47710 (N_47710,N_47236,N_46748);
and U47711 (N_47711,N_47058,N_46982);
xnor U47712 (N_47712,N_45572,N_47018);
nand U47713 (N_47713,N_46366,N_46158);
nand U47714 (N_47714,N_47228,N_46978);
or U47715 (N_47715,N_45461,N_45939);
and U47716 (N_47716,N_46548,N_46580);
and U47717 (N_47717,N_45926,N_47462);
and U47718 (N_47718,N_45091,N_47048);
or U47719 (N_47719,N_46802,N_45661);
and U47720 (N_47720,N_46697,N_47082);
and U47721 (N_47721,N_45296,N_45607);
and U47722 (N_47722,N_45184,N_45109);
or U47723 (N_47723,N_47268,N_45449);
or U47724 (N_47724,N_45079,N_45968);
and U47725 (N_47725,N_45239,N_46904);
nor U47726 (N_47726,N_46357,N_45855);
and U47727 (N_47727,N_47347,N_45304);
or U47728 (N_47728,N_46059,N_47306);
nor U47729 (N_47729,N_47414,N_45162);
xor U47730 (N_47730,N_46149,N_45157);
nor U47731 (N_47731,N_47457,N_45143);
nand U47732 (N_47732,N_47135,N_47475);
nand U47733 (N_47733,N_47473,N_45563);
nand U47734 (N_47734,N_46151,N_46966);
nor U47735 (N_47735,N_45679,N_45693);
nand U47736 (N_47736,N_47415,N_46183);
nand U47737 (N_47737,N_47137,N_46341);
nor U47738 (N_47738,N_45716,N_45037);
and U47739 (N_47739,N_45391,N_47288);
or U47740 (N_47740,N_46687,N_47176);
or U47741 (N_47741,N_46354,N_45291);
nor U47742 (N_47742,N_47213,N_47310);
nand U47743 (N_47743,N_46007,N_47464);
nor U47744 (N_47744,N_46453,N_45130);
and U47745 (N_47745,N_45525,N_46737);
nor U47746 (N_47746,N_45342,N_45988);
or U47747 (N_47747,N_46670,N_45093);
nand U47748 (N_47748,N_47131,N_45111);
or U47749 (N_47749,N_46204,N_46125);
or U47750 (N_47750,N_47184,N_47302);
nand U47751 (N_47751,N_46372,N_47158);
or U47752 (N_47752,N_46728,N_46325);
and U47753 (N_47753,N_46654,N_45732);
or U47754 (N_47754,N_46932,N_47063);
nor U47755 (N_47755,N_47211,N_47301);
or U47756 (N_47756,N_45281,N_45959);
or U47757 (N_47757,N_46531,N_47078);
nor U47758 (N_47758,N_47479,N_45778);
or U47759 (N_47759,N_46529,N_46743);
nand U47760 (N_47760,N_46082,N_45308);
nor U47761 (N_47761,N_46497,N_47489);
and U47762 (N_47762,N_46624,N_47484);
nand U47763 (N_47763,N_46682,N_45905);
nand U47764 (N_47764,N_45541,N_45851);
or U47765 (N_47765,N_45282,N_46484);
and U47766 (N_47766,N_47049,N_47220);
and U47767 (N_47767,N_46539,N_45706);
nor U47768 (N_47768,N_45863,N_45460);
or U47769 (N_47769,N_46180,N_46838);
xnor U47770 (N_47770,N_46561,N_47117);
nor U47771 (N_47771,N_45848,N_45218);
nand U47772 (N_47772,N_47030,N_46651);
and U47773 (N_47773,N_45515,N_46340);
or U47774 (N_47774,N_46335,N_45529);
or U47775 (N_47775,N_46875,N_46599);
nor U47776 (N_47776,N_45338,N_45768);
nand U47777 (N_47777,N_45808,N_45964);
nand U47778 (N_47778,N_45721,N_46972);
nor U47779 (N_47779,N_47094,N_45127);
nor U47780 (N_47780,N_47020,N_45268);
nand U47781 (N_47781,N_45334,N_45520);
nor U47782 (N_47782,N_46939,N_46816);
and U47783 (N_47783,N_47046,N_45962);
nor U47784 (N_47784,N_46440,N_45158);
nor U47785 (N_47785,N_46749,N_45825);
and U47786 (N_47786,N_45744,N_45298);
nand U47787 (N_47787,N_47466,N_45895);
nand U47788 (N_47788,N_47204,N_47344);
nor U47789 (N_47789,N_47000,N_47494);
nand U47790 (N_47790,N_46147,N_46406);
nand U47791 (N_47791,N_46746,N_47022);
xnor U47792 (N_47792,N_45767,N_46503);
and U47793 (N_47793,N_46588,N_47364);
xor U47794 (N_47794,N_46013,N_45351);
nor U47795 (N_47795,N_46385,N_45219);
or U47796 (N_47796,N_46189,N_45126);
xnor U47797 (N_47797,N_45346,N_47214);
and U47798 (N_47798,N_47308,N_47315);
nand U47799 (N_47799,N_45793,N_47287);
nor U47800 (N_47800,N_46573,N_45748);
nand U47801 (N_47801,N_45692,N_45728);
xor U47802 (N_47802,N_45104,N_45827);
nor U47803 (N_47803,N_46450,N_45792);
and U47804 (N_47804,N_46423,N_46418);
nor U47805 (N_47805,N_45674,N_46424);
nor U47806 (N_47806,N_45517,N_46282);
or U47807 (N_47807,N_46054,N_45051);
or U47808 (N_47808,N_46733,N_46231);
nand U47809 (N_47809,N_46762,N_45155);
nor U47810 (N_47810,N_46065,N_46618);
nand U47811 (N_47811,N_46868,N_46893);
and U47812 (N_47812,N_46017,N_46592);
nor U47813 (N_47813,N_47379,N_46795);
nand U47814 (N_47814,N_47477,N_47004);
or U47815 (N_47815,N_46105,N_47264);
xnor U47816 (N_47816,N_45713,N_45787);
xnor U47817 (N_47817,N_45250,N_45328);
nand U47818 (N_47818,N_46854,N_45416);
nand U47819 (N_47819,N_47476,N_45972);
xor U47820 (N_47820,N_46159,N_45299);
nor U47821 (N_47821,N_45936,N_46772);
or U47822 (N_47822,N_47067,N_47413);
and U47823 (N_47823,N_45568,N_45230);
nand U47824 (N_47824,N_46752,N_46756);
or U47825 (N_47825,N_45410,N_46232);
or U47826 (N_47826,N_45690,N_45153);
or U47827 (N_47827,N_46635,N_46170);
or U47828 (N_47828,N_45355,N_45352);
or U47829 (N_47829,N_46220,N_45321);
and U47830 (N_47830,N_46929,N_45049);
nor U47831 (N_47831,N_45718,N_46164);
or U47832 (N_47832,N_47119,N_46258);
or U47833 (N_47833,N_46454,N_45996);
and U47834 (N_47834,N_46196,N_46215);
nand U47835 (N_47835,N_47497,N_46956);
and U47836 (N_47836,N_45521,N_45556);
nor U47837 (N_47837,N_45365,N_47411);
and U47838 (N_47838,N_45816,N_46884);
or U47839 (N_47839,N_45782,N_46598);
xor U47840 (N_47840,N_45505,N_45457);
xor U47841 (N_47841,N_47028,N_46653);
or U47842 (N_47842,N_45435,N_45427);
and U47843 (N_47843,N_46053,N_47199);
nand U47844 (N_47844,N_46025,N_46870);
nor U47845 (N_47845,N_45396,N_45287);
nand U47846 (N_47846,N_46229,N_46351);
and U47847 (N_47847,N_45236,N_46878);
nand U47848 (N_47848,N_46725,N_47478);
and U47849 (N_47849,N_46153,N_47026);
nor U47850 (N_47850,N_46553,N_46383);
or U47851 (N_47851,N_47145,N_47461);
nand U47852 (N_47852,N_45625,N_45367);
or U47853 (N_47853,N_46512,N_47105);
nor U47854 (N_47854,N_46099,N_45637);
nand U47855 (N_47855,N_45650,N_45546);
nor U47856 (N_47856,N_46097,N_46869);
nand U47857 (N_47857,N_45994,N_45628);
nor U47858 (N_47858,N_45714,N_46808);
and U47859 (N_47859,N_46764,N_46344);
or U47860 (N_47860,N_45411,N_45198);
or U47861 (N_47861,N_47173,N_45434);
and U47862 (N_47862,N_45678,N_46305);
nor U47863 (N_47863,N_47453,N_47374);
and U47864 (N_47864,N_46886,N_47363);
or U47865 (N_47865,N_46413,N_46318);
or U47866 (N_47866,N_46610,N_45735);
and U47867 (N_47867,N_45665,N_47157);
nor U47868 (N_47868,N_47065,N_46550);
and U47869 (N_47869,N_45842,N_45136);
nand U47870 (N_47870,N_46436,N_45507);
nand U47871 (N_47871,N_46576,N_45086);
or U47872 (N_47872,N_45090,N_47125);
xor U47873 (N_47873,N_46636,N_45804);
xnor U47874 (N_47874,N_46247,N_47057);
or U47875 (N_47875,N_45818,N_46901);
and U47876 (N_47876,N_47104,N_46629);
nor U47877 (N_47877,N_45898,N_45917);
and U47878 (N_47878,N_45976,N_46704);
and U47879 (N_47879,N_45249,N_45548);
and U47880 (N_47880,N_45636,N_47092);
nand U47881 (N_47881,N_46840,N_47037);
nand U47882 (N_47882,N_47181,N_46861);
nor U47883 (N_47883,N_46433,N_47278);
nand U47884 (N_47884,N_46857,N_46460);
nor U47885 (N_47885,N_46617,N_46187);
nor U47886 (N_47886,N_45924,N_46731);
and U47887 (N_47887,N_45549,N_45711);
nand U47888 (N_47888,N_45319,N_45258);
or U47889 (N_47889,N_45089,N_46855);
and U47890 (N_47890,N_46643,N_47360);
nor U47891 (N_47891,N_46992,N_47369);
nand U47892 (N_47892,N_45069,N_45835);
xor U47893 (N_47893,N_45295,N_46999);
nand U47894 (N_47894,N_47147,N_46575);
nand U47895 (N_47895,N_45730,N_45861);
or U47896 (N_47896,N_47008,N_46505);
nor U47897 (N_47897,N_46364,N_47486);
nand U47898 (N_47898,N_46104,N_46447);
nand U47899 (N_47899,N_47196,N_46371);
and U47900 (N_47900,N_46620,N_46522);
and U47901 (N_47901,N_46336,N_46963);
xor U47902 (N_47902,N_45850,N_45623);
or U47903 (N_47903,N_45151,N_45324);
nand U47904 (N_47904,N_45514,N_46438);
nand U47905 (N_47905,N_45468,N_46200);
or U47906 (N_47906,N_46850,N_47332);
or U47907 (N_47907,N_45875,N_47290);
nand U47908 (N_47908,N_45429,N_47109);
xnor U47909 (N_47909,N_45147,N_46323);
nand U47910 (N_47910,N_45425,N_45526);
and U47911 (N_47911,N_45647,N_47316);
and U47912 (N_47912,N_47454,N_45869);
xnor U47913 (N_47913,N_46923,N_47276);
or U47914 (N_47914,N_45677,N_47098);
and U47915 (N_47915,N_47300,N_46888);
nand U47916 (N_47916,N_45283,N_45913);
xor U47917 (N_47917,N_46760,N_45759);
nand U47918 (N_47918,N_45108,N_45065);
nor U47919 (N_47919,N_45044,N_45010);
or U47920 (N_47920,N_45402,N_46686);
or U47921 (N_47921,N_47421,N_46652);
nand U47922 (N_47922,N_46195,N_46833);
nand U47923 (N_47923,N_46129,N_47399);
nand U47924 (N_47924,N_45394,N_45969);
nor U47925 (N_47925,N_46800,N_47367);
or U47926 (N_47926,N_45003,N_47056);
or U47927 (N_47927,N_45054,N_46085);
or U47928 (N_47928,N_46112,N_45512);
nand U47929 (N_47929,N_46420,N_46313);
or U47930 (N_47930,N_46257,N_47225);
and U47931 (N_47931,N_46994,N_45758);
xnor U47932 (N_47932,N_46202,N_45246);
or U47933 (N_47933,N_46027,N_46148);
nor U47934 (N_47934,N_45210,N_46510);
and U47935 (N_47935,N_46138,N_45231);
and U47936 (N_47936,N_45269,N_45984);
xor U47937 (N_47937,N_47356,N_47322);
nand U47938 (N_47938,N_45205,N_46157);
nand U47939 (N_47939,N_46165,N_46896);
or U47940 (N_47940,N_47418,N_46347);
and U47941 (N_47941,N_47025,N_46537);
xnor U47942 (N_47942,N_46156,N_46632);
nand U47943 (N_47943,N_46934,N_45122);
nand U47944 (N_47944,N_45050,N_46846);
and U47945 (N_47945,N_46317,N_45031);
nor U47946 (N_47946,N_46363,N_45648);
or U47947 (N_47947,N_47151,N_46774);
nand U47948 (N_47948,N_46477,N_45879);
and U47949 (N_47949,N_46502,N_46292);
or U47950 (N_47950,N_46616,N_45387);
and U47951 (N_47951,N_46688,N_46547);
xnor U47952 (N_47952,N_47341,N_47474);
or U47953 (N_47953,N_45322,N_46368);
nor U47954 (N_47954,N_46515,N_47051);
or U47955 (N_47955,N_45055,N_46322);
or U47956 (N_47956,N_47128,N_46211);
and U47957 (N_47957,N_45068,N_45194);
and U47958 (N_47958,N_47139,N_47130);
and U47959 (N_47959,N_46559,N_46272);
nand U47960 (N_47960,N_45373,N_46412);
nand U47961 (N_47961,N_45146,N_46582);
xor U47962 (N_47962,N_47010,N_45906);
or U47963 (N_47963,N_46491,N_47377);
nand U47964 (N_47964,N_47331,N_45545);
and U47965 (N_47965,N_46914,N_46283);
nand U47966 (N_47966,N_47354,N_47283);
xor U47967 (N_47967,N_47190,N_46771);
or U47968 (N_47968,N_45096,N_46713);
and U47969 (N_47969,N_45028,N_46037);
nand U47970 (N_47970,N_46181,N_45213);
nor U47971 (N_47971,N_46474,N_47370);
nor U47972 (N_47972,N_45513,N_45004);
nand U47973 (N_47973,N_45347,N_46089);
or U47974 (N_47974,N_47470,N_46429);
and U47975 (N_47975,N_45440,N_46604);
or U47976 (N_47976,N_46829,N_45472);
or U47977 (N_47977,N_46094,N_46102);
nand U47978 (N_47978,N_45916,N_46127);
nand U47979 (N_47979,N_45668,N_47136);
nor U47980 (N_47980,N_46076,N_45958);
and U47981 (N_47981,N_47171,N_46359);
xor U47982 (N_47982,N_45509,N_46607);
nor U47983 (N_47983,N_45700,N_47396);
nor U47984 (N_47984,N_45965,N_46396);
nor U47985 (N_47985,N_45860,N_47438);
or U47986 (N_47986,N_47170,N_45597);
xor U47987 (N_47987,N_45134,N_46793);
nand U47988 (N_47988,N_45901,N_45114);
or U47989 (N_47989,N_47083,N_46584);
nand U47990 (N_47990,N_47335,N_45056);
xnor U47991 (N_47991,N_46877,N_46044);
nand U47992 (N_47992,N_45831,N_46593);
and U47993 (N_47993,N_46192,N_46213);
nor U47994 (N_47994,N_46392,N_46379);
nor U47995 (N_47995,N_45392,N_47485);
xnor U47996 (N_47996,N_45007,N_45598);
nand U47997 (N_47997,N_45585,N_46899);
nand U47998 (N_47998,N_46908,N_47326);
or U47999 (N_47999,N_47277,N_45005);
or U48000 (N_48000,N_45594,N_46427);
nand U48001 (N_48001,N_45586,N_46611);
or U48002 (N_48002,N_46526,N_45182);
nand U48003 (N_48003,N_45316,N_46823);
nor U48004 (N_48004,N_45975,N_46279);
and U48005 (N_48005,N_45253,N_45405);
nand U48006 (N_48006,N_46742,N_47286);
or U48007 (N_48007,N_45286,N_45038);
nor U48008 (N_48008,N_45053,N_47245);
nor U48009 (N_48009,N_46591,N_45061);
nor U48010 (N_48010,N_46664,N_46331);
and U48011 (N_48011,N_45765,N_45626);
and U48012 (N_48012,N_45455,N_45251);
xor U48013 (N_48013,N_46139,N_45538);
nand U48014 (N_48014,N_45954,N_46227);
nor U48015 (N_48015,N_46179,N_46852);
nand U48016 (N_48016,N_45228,N_45593);
nand U48017 (N_48017,N_47361,N_46942);
and U48018 (N_48018,N_45534,N_46809);
or U48019 (N_48019,N_45789,N_46381);
and U48020 (N_48020,N_46564,N_46717);
nor U48021 (N_48021,N_47134,N_46382);
nor U48022 (N_48022,N_45329,N_46135);
nor U48023 (N_48023,N_45588,N_47198);
nand U48024 (N_48024,N_47423,N_46081);
and U48025 (N_48025,N_45543,N_46472);
xnor U48026 (N_48026,N_46375,N_46832);
xor U48027 (N_48027,N_46144,N_46478);
or U48028 (N_48028,N_47471,N_45880);
and U48029 (N_48029,N_45609,N_45012);
or U48030 (N_48030,N_45137,N_45813);
nand U48031 (N_48031,N_46820,N_46009);
xnor U48032 (N_48032,N_47441,N_45999);
nor U48033 (N_48033,N_47116,N_45697);
nor U48034 (N_48034,N_45640,N_47178);
nand U48035 (N_48035,N_46814,N_45675);
and U48036 (N_48036,N_46262,N_45473);
or U48037 (N_48037,N_46405,N_46289);
or U48038 (N_48038,N_45098,N_46974);
or U48039 (N_48039,N_47230,N_46461);
nand U48040 (N_48040,N_46465,N_45378);
nor U48041 (N_48041,N_46018,N_47202);
nand U48042 (N_48042,N_46657,N_45116);
nor U48043 (N_48043,N_47034,N_46633);
nor U48044 (N_48044,N_45945,N_45260);
nand U48045 (N_48045,N_47126,N_47330);
xnor U48046 (N_48046,N_45833,N_47072);
or U48047 (N_48047,N_45256,N_45822);
and U48048 (N_48048,N_45518,N_45979);
and U48049 (N_48049,N_46711,N_46735);
or U48050 (N_48050,N_45986,N_45952);
or U48051 (N_48051,N_47296,N_45261);
and U48052 (N_48052,N_46568,N_45870);
nor U48053 (N_48053,N_47468,N_46738);
nand U48054 (N_48054,N_45297,N_47419);
or U48055 (N_48055,N_45052,N_46810);
nand U48056 (N_48056,N_46041,N_47073);
and U48057 (N_48057,N_46033,N_46676);
and U48058 (N_48058,N_45066,N_46707);
xor U48059 (N_48059,N_45622,N_45166);
and U48060 (N_48060,N_45220,N_45470);
nor U48061 (N_48061,N_45770,N_45381);
and U48062 (N_48062,N_47208,N_47246);
or U48063 (N_48063,N_47142,N_47183);
or U48064 (N_48064,N_45175,N_47154);
and U48065 (N_48065,N_46520,N_46222);
nor U48066 (N_48066,N_46458,N_46172);
nor U48067 (N_48067,N_46957,N_46238);
and U48068 (N_48068,N_46830,N_46880);
and U48069 (N_48069,N_45368,N_46332);
nor U48070 (N_48070,N_45094,N_45922);
nand U48071 (N_48071,N_47160,N_45775);
and U48072 (N_48072,N_46602,N_46691);
nand U48073 (N_48073,N_46043,N_45985);
nand U48074 (N_48074,N_45008,N_46150);
and U48075 (N_48075,N_45845,N_46736);
nor U48076 (N_48076,N_47009,N_47144);
nand U48077 (N_48077,N_46933,N_46732);
and U48078 (N_48078,N_45554,N_47450);
nand U48079 (N_48079,N_45741,N_45479);
or U48080 (N_48080,N_46481,N_45885);
or U48081 (N_48081,N_45337,N_46048);
and U48082 (N_48082,N_45013,N_47089);
nand U48083 (N_48083,N_45300,N_46096);
xor U48084 (N_48084,N_46675,N_46572);
nor U48085 (N_48085,N_46776,N_46791);
and U48086 (N_48086,N_46003,N_46811);
nor U48087 (N_48087,N_46700,N_47339);
nor U48088 (N_48088,N_47249,N_46754);
and U48089 (N_48089,N_47383,N_47123);
nand U48090 (N_48090,N_45025,N_46796);
nor U48091 (N_48091,N_47329,N_45814);
and U48092 (N_48092,N_46920,N_46546);
nor U48093 (N_48093,N_45961,N_46964);
or U48094 (N_48094,N_45292,N_45307);
or U48095 (N_48095,N_45638,N_46995);
or U48096 (N_48096,N_46542,N_47041);
nand U48097 (N_48097,N_47039,N_47312);
nor U48098 (N_48098,N_47070,N_46555);
or U48099 (N_48099,N_45819,N_47493);
and U48100 (N_48100,N_46918,N_46443);
and U48101 (N_48101,N_46803,N_46056);
or U48102 (N_48102,N_45547,N_45935);
and U48103 (N_48103,N_45177,N_46066);
or U48104 (N_48104,N_47499,N_47463);
nor U48105 (N_48105,N_45030,N_46409);
xnor U48106 (N_48106,N_46173,N_46853);
xor U48107 (N_48107,N_45734,N_46398);
nand U48108 (N_48108,N_47093,N_47006);
and U48109 (N_48109,N_46702,N_47141);
xor U48110 (N_48110,N_46249,N_45841);
nand U48111 (N_48111,N_46162,N_46388);
and U48112 (N_48112,N_46511,N_45447);
and U48113 (N_48113,N_47496,N_45834);
nor U48114 (N_48114,N_45273,N_46121);
or U48115 (N_48115,N_45570,N_46293);
or U48116 (N_48116,N_45027,N_47159);
or U48117 (N_48117,N_46988,N_46549);
nand U48118 (N_48118,N_45214,N_46182);
and U48119 (N_48119,N_47311,N_47064);
nor U48120 (N_48120,N_45921,N_46337);
or U48121 (N_48121,N_46781,N_45356);
nand U48122 (N_48122,N_46126,N_45892);
nor U48123 (N_48123,N_46962,N_47481);
nor U48124 (N_48124,N_46724,N_46812);
and U48125 (N_48125,N_47088,N_46273);
and U48126 (N_48126,N_46263,N_46944);
nand U48127 (N_48127,N_46175,N_47218);
and U48128 (N_48128,N_45990,N_47069);
nand U48129 (N_48129,N_45596,N_45474);
and U48130 (N_48130,N_46462,N_45343);
or U48131 (N_48131,N_45738,N_46668);
nor U48132 (N_48132,N_46403,N_46507);
or U48133 (N_48133,N_46851,N_45884);
and U48134 (N_48134,N_47303,N_46067);
nor U48135 (N_48135,N_47498,N_45839);
nand U48136 (N_48136,N_45877,N_46473);
xnor U48137 (N_48137,N_45278,N_46931);
nor U48138 (N_48138,N_45783,N_45497);
nand U48139 (N_48139,N_45737,N_45763);
and U48140 (N_48140,N_46952,N_45270);
nor U48141 (N_48141,N_45523,N_45874);
and U48142 (N_48142,N_45100,N_45412);
nor U48143 (N_48143,N_45684,N_46882);
nand U48144 (N_48144,N_46614,N_46109);
and U48145 (N_48145,N_45344,N_45912);
and U48146 (N_48146,N_46977,N_46224);
nand U48147 (N_48147,N_47324,N_45248);
or U48148 (N_48148,N_45909,N_45397);
nor U48149 (N_48149,N_46452,N_45873);
and U48150 (N_48150,N_45211,N_46286);
nand U48151 (N_48151,N_47032,N_45408);
or U48152 (N_48152,N_45326,N_46967);
nand U48153 (N_48153,N_46740,N_47381);
and U48154 (N_48154,N_45764,N_47259);
or U48155 (N_48155,N_45489,N_45315);
xnor U48156 (N_48156,N_46825,N_46038);
xor U48157 (N_48157,N_46769,N_47043);
and U48158 (N_48158,N_45881,N_46088);
and U48159 (N_48159,N_46411,N_47091);
or U48160 (N_48160,N_45486,N_46597);
xnor U48161 (N_48161,N_45893,N_47227);
or U48162 (N_48162,N_46119,N_46297);
nand U48163 (N_48163,N_45997,N_47054);
or U48164 (N_48164,N_46788,N_45074);
nand U48165 (N_48165,N_45107,N_45902);
nand U48166 (N_48166,N_46223,N_47395);
xor U48167 (N_48167,N_46244,N_46916);
nand U48168 (N_48168,N_46892,N_45309);
and U48169 (N_48169,N_46432,N_45699);
nand U48170 (N_48170,N_46482,N_47036);
or U48171 (N_48171,N_45840,N_45550);
and U48172 (N_48172,N_45192,N_47107);
nor U48173 (N_48173,N_45419,N_45399);
and U48174 (N_48174,N_46142,N_45119);
nand U48175 (N_48175,N_46072,N_45046);
and U48176 (N_48176,N_47487,N_47197);
nor U48177 (N_48177,N_45432,N_45067);
and U48178 (N_48178,N_45847,N_46240);
nor U48179 (N_48179,N_46264,N_45762);
and U48180 (N_48180,N_47206,N_46673);
and U48181 (N_48181,N_45595,N_47293);
nand U48182 (N_48182,N_45159,N_47319);
nand U48183 (N_48183,N_46990,N_45740);
nor U48184 (N_48184,N_46784,N_47272);
xnor U48185 (N_48185,N_47224,N_45371);
or U48186 (N_48186,N_45852,N_47223);
xor U48187 (N_48187,N_45139,N_45888);
or U48188 (N_48188,N_45927,N_47422);
and U48189 (N_48189,N_46801,N_45390);
or U48190 (N_48190,N_46391,N_45488);
and U48191 (N_48191,N_47406,N_46208);
and U48192 (N_48192,N_47402,N_46416);
or U48193 (N_48193,N_46384,N_46804);
and U48194 (N_48194,N_46658,N_45092);
and U48195 (N_48195,N_46596,N_47238);
or U48196 (N_48196,N_45981,N_46069);
and U48197 (N_48197,N_46441,N_45761);
nor U48198 (N_48198,N_46940,N_46308);
and U48199 (N_48199,N_47011,N_46390);
nor U48200 (N_48200,N_45722,N_47292);
or U48201 (N_48201,N_45354,N_46849);
or U48202 (N_48202,N_45817,N_47346);
or U48203 (N_48203,N_45169,N_46216);
or U48204 (N_48204,N_45896,N_45500);
and U48205 (N_48205,N_45838,N_46714);
or U48206 (N_48206,N_46836,N_45105);
nor U48207 (N_48207,N_45632,N_46487);
nand U48208 (N_48208,N_45318,N_45043);
or U48209 (N_48209,N_47267,N_46178);
or U48210 (N_48210,N_47077,N_45456);
and U48211 (N_48211,N_47066,N_46556);
nor U48212 (N_48212,N_46077,N_46137);
and U48213 (N_48213,N_46601,N_46459);
and U48214 (N_48214,N_46408,N_45032);
and U48215 (N_48215,N_46123,N_47189);
or U48216 (N_48216,N_46463,N_45582);
nor U48217 (N_48217,N_45453,N_47045);
or U48218 (N_48218,N_45280,N_45404);
and U48219 (N_48219,N_45469,N_45084);
or U48220 (N_48220,N_46532,N_46578);
nand U48221 (N_48221,N_45654,N_47194);
and U48222 (N_48222,N_45756,N_46087);
nand U48223 (N_48223,N_46184,N_45807);
or U48224 (N_48224,N_47392,N_45889);
and U48225 (N_48225,N_45483,N_45097);
nand U48226 (N_48226,N_45569,N_45953);
and U48227 (N_48227,N_47108,N_45686);
nor U48228 (N_48228,N_47386,N_46678);
nor U48229 (N_48229,N_46630,N_47002);
and U48230 (N_48230,N_45821,N_46304);
xnor U48231 (N_48231,N_47209,N_46345);
nand U48232 (N_48232,N_45099,N_47420);
or U48233 (N_48233,N_45305,N_46268);
and U48234 (N_48234,N_46692,N_47055);
or U48235 (N_48235,N_46060,N_46219);
xnor U48236 (N_48236,N_47221,N_47118);
or U48237 (N_48237,N_46448,N_47337);
or U48238 (N_48238,N_46889,N_45784);
or U48239 (N_48239,N_45095,N_45791);
and U48240 (N_48240,N_45973,N_46807);
nand U48241 (N_48241,N_47382,N_45142);
or U48242 (N_48242,N_45443,N_46193);
nor U48243 (N_48243,N_46480,N_45149);
or U48244 (N_48244,N_45277,N_45599);
and U48245 (N_48245,N_46533,N_45729);
nor U48246 (N_48246,N_46030,N_47257);
nand U48247 (N_48247,N_45612,N_45788);
nand U48248 (N_48248,N_47368,N_45942);
nor U48249 (N_48249,N_46169,N_45314);
nand U48250 (N_48250,N_47150,N_46467);
nand U48251 (N_48251,N_47235,N_47219);
nand U48252 (N_48252,N_45471,N_45535);
or U48253 (N_48253,N_46757,N_46399);
or U48254 (N_48254,N_47050,N_45933);
or U48255 (N_48255,N_47338,N_45573);
or U48256 (N_48256,N_46997,N_46015);
or U48257 (N_48257,N_46778,N_46437);
xor U48258 (N_48258,N_46834,N_46333);
nand U48259 (N_48259,N_47432,N_46538);
and U48260 (N_48260,N_46951,N_45238);
or U48261 (N_48261,N_47095,N_45075);
nor U48262 (N_48262,N_47426,N_46306);
nor U48263 (N_48263,N_47027,N_45694);
xor U48264 (N_48264,N_46005,N_47488);
or U48265 (N_48265,N_46685,N_45477);
or U48266 (N_48266,N_45800,N_45302);
and U48267 (N_48267,N_45400,N_46590);
nand U48268 (N_48268,N_45946,N_45240);
nand U48269 (N_48269,N_46968,N_47237);
nand U48270 (N_48270,N_45047,N_46446);
nor U48271 (N_48271,N_45064,N_45865);
or U48272 (N_48272,N_45780,N_47469);
nor U48273 (N_48273,N_47084,N_46152);
nor U48274 (N_48274,N_47215,N_46185);
and U48275 (N_48275,N_45562,N_45832);
nor U48276 (N_48276,N_47103,N_47265);
and U48277 (N_48277,N_45226,N_46485);
xor U48278 (N_48278,N_46355,N_45271);
or U48279 (N_48279,N_45375,N_47155);
xnor U48280 (N_48280,N_45209,N_45904);
nand U48281 (N_48281,N_45362,N_46585);
nor U48282 (N_48282,N_46523,N_46362);
or U48283 (N_48283,N_46243,N_45872);
nor U48284 (N_48284,N_45323,N_45496);
nand U48285 (N_48285,N_45229,N_47358);
or U48286 (N_48286,N_45769,N_45720);
and U48287 (N_48287,N_46981,N_45284);
and U48288 (N_48288,N_46667,N_45341);
nor U48289 (N_48289,N_45983,N_47143);
nor U48290 (N_48290,N_46897,N_45522);
or U48291 (N_48291,N_45110,N_47053);
nand U48292 (N_48292,N_47068,N_45651);
and U48293 (N_48293,N_45727,N_46468);
and U48294 (N_48294,N_46476,N_46160);
and U48295 (N_48295,N_47024,N_46146);
nand U48296 (N_48296,N_45141,N_45991);
or U48297 (N_48297,N_46250,N_46113);
and U48298 (N_48298,N_46898,N_47351);
or U48299 (N_48299,N_45233,N_46622);
and U48300 (N_48300,N_45856,N_45731);
xor U48301 (N_48301,N_47253,N_47186);
and U48302 (N_48302,N_47029,N_46730);
nand U48303 (N_48303,N_45736,N_46051);
and U48304 (N_48304,N_46092,N_46036);
or U48305 (N_48305,N_45163,N_47393);
nor U48306 (N_48306,N_46696,N_46551);
nor U48307 (N_48307,N_45949,N_45670);
nand U48308 (N_48308,N_45083,N_45918);
nand U48309 (N_48309,N_46111,N_45406);
and U48310 (N_48310,N_46911,N_46358);
nand U48311 (N_48311,N_46513,N_46773);
nand U48312 (N_48312,N_46228,N_45516);
and U48313 (N_48313,N_46770,N_46198);
or U48314 (N_48314,N_47433,N_45613);
and U48315 (N_48315,N_47222,N_46455);
nand U48316 (N_48316,N_46683,N_46824);
or U48317 (N_48317,N_46197,N_46979);
xnor U48318 (N_48318,N_45170,N_46287);
nand U48319 (N_48319,N_46703,N_47096);
and U48320 (N_48320,N_45777,N_45395);
nor U48321 (N_48321,N_47445,N_46494);
nand U48322 (N_48322,N_47333,N_45485);
nand U48323 (N_48323,N_47297,N_46915);
nor U48324 (N_48324,N_47075,N_47439);
nand U48325 (N_48325,N_46177,N_45725);
or U48326 (N_48326,N_46567,N_46837);
nand U48327 (N_48327,N_45121,N_45866);
nand U48328 (N_48328,N_46469,N_46656);
and U48329 (N_48329,N_47416,N_46646);
nand U48330 (N_48330,N_46415,N_47076);
nor U48331 (N_48331,N_46710,N_45459);
nand U48332 (N_48332,N_45774,N_45076);
nor U48333 (N_48333,N_45423,N_45499);
nor U48334 (N_48334,N_47321,N_45798);
nand U48335 (N_48335,N_46937,N_46806);
nand U48336 (N_48336,N_45178,N_45481);
or U48337 (N_48337,N_47101,N_47459);
or U48338 (N_48338,N_47252,N_45235);
or U48339 (N_48339,N_45023,N_45723);
xor U48340 (N_48340,N_47179,N_47226);
or U48341 (N_48341,N_46110,N_47040);
and U48342 (N_48342,N_45349,N_45152);
or U48343 (N_48343,N_47080,N_47180);
nand U48344 (N_48344,N_47313,N_47352);
nand U48345 (N_48345,N_47156,N_46186);
and U48346 (N_48346,N_46891,N_45480);
nor U48347 (N_48347,N_47295,N_45701);
and U48348 (N_48348,N_45183,N_46389);
nand U48349 (N_48349,N_46118,N_45290);
and U48350 (N_48350,N_45683,N_45288);
or U48351 (N_48351,N_45966,N_45760);
xor U48352 (N_48352,N_46965,N_46360);
or U48353 (N_48353,N_47492,N_46034);
and U48354 (N_48354,N_46706,N_47232);
nor U48355 (N_48355,N_45332,N_45828);
nor U48356 (N_48356,N_46241,N_46975);
or U48357 (N_48357,N_46045,N_47188);
or U48358 (N_48358,N_46207,N_46519);
nor U48359 (N_48359,N_46245,N_45589);
nor U48360 (N_48360,N_45689,N_45826);
nor U48361 (N_48361,N_47031,N_46718);
nor U48362 (N_48362,N_46943,N_46035);
nor U48363 (N_48363,N_46647,N_46339);
nor U48364 (N_48364,N_46831,N_47412);
nand U48365 (N_48365,N_46492,N_45653);
and U48366 (N_48366,N_46374,N_45934);
xnor U48367 (N_48367,N_45294,N_47429);
xnor U48368 (N_48368,N_46073,N_45145);
and U48369 (N_48369,N_45766,N_45154);
nor U48370 (N_48370,N_47336,N_45313);
or U48371 (N_48371,N_46380,N_45150);
nand U48372 (N_48372,N_47323,N_45383);
nand U48373 (N_48373,N_46958,N_45103);
nor U48374 (N_48374,N_46534,N_46910);
nor U48375 (N_48375,N_45960,N_47425);
nor U48376 (N_48376,N_46303,N_46445);
xnor U48377 (N_48377,N_46140,N_45846);
nor U48378 (N_48378,N_45073,N_47446);
and U48379 (N_48379,N_45060,N_47090);
nor U48380 (N_48380,N_46536,N_46872);
or U48381 (N_48381,N_46242,N_46970);
nand U48382 (N_48382,N_46428,N_46863);
or U48383 (N_48383,N_47182,N_45366);
or U48384 (N_48384,N_47153,N_46612);
nor U48385 (N_48385,N_45312,N_45719);
or U48386 (N_48386,N_46295,N_45551);
xor U48387 (N_48387,N_45360,N_45797);
nand U48388 (N_48388,N_46490,N_45786);
or U48389 (N_48389,N_46400,N_45646);
nand U48390 (N_48390,N_47165,N_45531);
nor U48391 (N_48391,N_47015,N_46466);
nand U48392 (N_48392,N_45601,N_46579);
nand U48393 (N_48393,N_46346,N_47400);
nor U48394 (N_48394,N_47307,N_46421);
and U48395 (N_48395,N_46765,N_46499);
nor U48396 (N_48396,N_45542,N_47016);
or U48397 (N_48397,N_45712,N_46689);
or U48398 (N_48398,N_45325,N_46516);
and U48399 (N_48399,N_45006,N_45590);
or U48400 (N_48400,N_46410,N_47389);
or U48401 (N_48401,N_46042,N_45181);
and U48402 (N_48402,N_45033,N_46819);
nor U48403 (N_48403,N_46050,N_45967);
and U48404 (N_48404,N_46107,N_46902);
nand U48405 (N_48405,N_45208,N_45630);
or U48406 (N_48406,N_45955,N_45161);
nand U48407 (N_48407,N_46426,N_47491);
and U48408 (N_48408,N_45113,N_46296);
nand U48409 (N_48409,N_46493,N_46545);
nor U48410 (N_48410,N_46314,N_45602);
nor U48411 (N_48411,N_45971,N_46276);
xor U48412 (N_48412,N_46444,N_46230);
or U48413 (N_48413,N_45910,N_45174);
and U48414 (N_48414,N_45908,N_46378);
nand U48415 (N_48415,N_47035,N_45026);
nand U48416 (N_48416,N_47161,N_45600);
nor U48417 (N_48417,N_46842,N_45393);
and U48418 (N_48418,N_45978,N_47397);
or U48419 (N_48419,N_45871,N_47318);
and U48420 (N_48420,N_45426,N_46827);
nand U48421 (N_48421,N_45660,N_46407);
and U48422 (N_48422,N_45036,N_46291);
or U48423 (N_48423,N_46750,N_46251);
nor U48424 (N_48424,N_47133,N_45063);
nor U48425 (N_48425,N_45937,N_46052);
nand U48426 (N_48426,N_46913,N_46080);
or U48427 (N_48427,N_45421,N_45687);
and U48428 (N_48428,N_47260,N_47097);
nand U48429 (N_48429,N_45592,N_45951);
nand U48430 (N_48430,N_45803,N_46751);
nand U48431 (N_48431,N_46848,N_46246);
xor U48432 (N_48432,N_46613,N_45215);
and U48433 (N_48433,N_45484,N_46217);
or U48434 (N_48434,N_45475,N_45581);
and U48435 (N_48435,N_46562,N_46299);
nor U48436 (N_48436,N_45532,N_46032);
nor U48437 (N_48437,N_45160,N_46430);
or U48438 (N_48438,N_46628,N_47285);
and U48439 (N_48439,N_46566,N_47378);
nor U48440 (N_48440,N_47483,N_46256);
and U48441 (N_48441,N_46634,N_47200);
xnor U48442 (N_48442,N_45117,N_47403);
or U48443 (N_48443,N_47279,N_46783);
nor U48444 (N_48444,N_47291,N_47482);
nand U48445 (N_48445,N_46679,N_46316);
nand U48446 (N_48446,N_46014,N_47456);
nor U48447 (N_48447,N_46535,N_46955);
nand U48448 (N_48448,N_45796,N_46864);
and U48449 (N_48449,N_45658,N_45708);
xnor U48450 (N_48450,N_46166,N_45041);
nand U48451 (N_48451,N_46627,N_45673);
nor U48452 (N_48452,N_45088,N_45403);
and U48453 (N_48453,N_47074,N_46422);
or U48454 (N_48454,N_45511,N_45059);
nand U48455 (N_48455,N_46690,N_45566);
xnor U48456 (N_48456,N_46637,N_45441);
nand U48457 (N_48457,N_45565,N_46134);
nand U48458 (N_48458,N_47216,N_45062);
or U48459 (N_48459,N_45448,N_46867);
or U48460 (N_48460,N_45987,N_45862);
and U48461 (N_48461,N_46660,N_45743);
nand U48462 (N_48462,N_45843,N_46984);
or U48463 (N_48463,N_47353,N_45024);
or U48464 (N_48464,N_45963,N_46695);
nand U48465 (N_48465,N_46049,N_47012);
nor U48466 (N_48466,N_46859,N_46936);
and U48467 (N_48467,N_47434,N_47387);
and U48468 (N_48468,N_46205,N_45644);
nor U48469 (N_48469,N_46404,N_46315);
or U48470 (N_48470,N_45462,N_45801);
nand U48471 (N_48471,N_45165,N_46615);
and U48472 (N_48472,N_45221,N_47362);
nand U48473 (N_48473,N_46659,N_46141);
nand U48474 (N_48474,N_45533,N_46903);
or U48475 (N_48475,N_47342,N_45810);
nor U48476 (N_48476,N_47407,N_45045);
nand U48477 (N_48477,N_45502,N_47262);
nand U48478 (N_48478,N_46779,N_46269);
nor U48479 (N_48479,N_46365,N_46031);
nand U48480 (N_48480,N_46927,N_46530);
nor U48481 (N_48481,N_46095,N_47350);
and U48482 (N_48482,N_46199,N_47127);
nand U48483 (N_48483,N_46720,N_45454);
and U48484 (N_48484,N_46275,N_45244);
nand U48485 (N_48485,N_46993,N_46705);
and U48486 (N_48486,N_46237,N_45685);
nand U48487 (N_48487,N_46528,N_46873);
and U48488 (N_48488,N_45019,N_47244);
nor U48489 (N_48489,N_46334,N_46071);
nand U48490 (N_48490,N_46938,N_45385);
or U48491 (N_48491,N_47424,N_46941);
nand U48492 (N_48492,N_46715,N_45844);
nor U48493 (N_48493,N_45262,N_47187);
nor U48494 (N_48494,N_45199,N_45752);
xor U48495 (N_48495,N_47440,N_46996);
and U48496 (N_48496,N_45264,N_45751);
nor U48497 (N_48497,N_46501,N_45571);
and U48498 (N_48498,N_45790,N_46969);
and U48499 (N_48499,N_45336,N_46907);
nor U48500 (N_48500,N_46554,N_47229);
or U48501 (N_48501,N_46552,N_45883);
and U48502 (N_48502,N_46395,N_47410);
nand U48503 (N_48503,N_45333,N_46190);
xnor U48504 (N_48504,N_45189,N_46623);
and U48505 (N_48505,N_47467,N_45430);
nand U48506 (N_48506,N_46361,N_46021);
nor U48507 (N_48507,N_46655,N_45733);
nand U48508 (N_48508,N_46845,N_46201);
nor U48509 (N_48509,N_45537,N_46132);
nor U48510 (N_48510,N_46508,N_45242);
xnor U48511 (N_48511,N_45627,N_47448);
nand U48512 (N_48512,N_45002,N_47111);
nand U48513 (N_48513,N_45682,N_45669);
or U48514 (N_48514,N_46356,N_45265);
or U48515 (N_48515,N_45604,N_46029);
xnor U48516 (N_48516,N_45436,N_45618);
and U48517 (N_48517,N_46641,N_45464);
nand U48518 (N_48518,N_46188,N_46860);
nand U48519 (N_48519,N_46312,N_46486);
or U48520 (N_48520,N_45331,N_47495);
and U48521 (N_48521,N_45837,N_46414);
and U48522 (N_48522,N_45691,N_45915);
nand U48523 (N_48523,N_47317,N_46319);
or U48524 (N_48524,N_46642,N_47343);
and U48525 (N_48525,N_45635,N_46729);
and U48526 (N_48526,N_46680,N_45345);
or U48527 (N_48527,N_46470,N_46349);
nand U48528 (N_48528,N_47269,N_46280);
xor U48529 (N_48529,N_46343,N_45676);
or U48530 (N_48530,N_45899,N_46744);
or U48531 (N_48531,N_45943,N_46924);
and U48532 (N_48532,N_45557,N_47334);
nor U48533 (N_48533,N_45247,N_46154);
and U48534 (N_48534,N_45940,N_45799);
or U48535 (N_48535,N_45854,N_46790);
and U48536 (N_48536,N_46817,N_45364);
nand U48537 (N_48537,N_46794,N_45634);
nand U48538 (N_48538,N_45225,N_45656);
or U48539 (N_48539,N_47357,N_46226);
xnor U48540 (N_48540,N_46723,N_46449);
xor U48541 (N_48541,N_47061,N_46417);
nor U48542 (N_48542,N_45950,N_46558);
xor U48543 (N_48543,N_47458,N_46517);
nor U48544 (N_48544,N_47071,N_46212);
and U48545 (N_48545,N_45576,N_47289);
or U48546 (N_48546,N_46218,N_46514);
xnor U48547 (N_48547,N_45664,N_45414);
xor U48548 (N_48548,N_46301,N_45078);
nand U48549 (N_48549,N_45560,N_46191);
nor U48550 (N_48550,N_47320,N_46039);
or U48551 (N_48551,N_45574,N_46506);
and U48552 (N_48552,N_46509,N_47247);
nor U48553 (N_48553,N_45528,N_45207);
nand U48554 (N_48554,N_46856,N_46265);
and U48555 (N_48555,N_46782,N_45327);
and U48556 (N_48556,N_46058,N_45424);
nor U48557 (N_48557,N_46300,N_47390);
or U48558 (N_48558,N_45923,N_47114);
nand U48559 (N_48559,N_45401,N_45363);
xnor U48560 (N_48560,N_46935,N_46541);
and U48561 (N_48561,N_45771,N_45259);
and U48562 (N_48562,N_46626,N_46712);
xor U48563 (N_48563,N_45970,N_45639);
nor U48564 (N_48564,N_45144,N_45029);
nand U48565 (N_48565,N_46206,N_45823);
nor U48566 (N_48566,N_46797,N_46681);
or U48567 (N_48567,N_46495,N_45580);
nor U48568 (N_48568,N_45384,N_45853);
or U48569 (N_48569,N_46799,N_45255);
and U48570 (N_48570,N_45530,N_46338);
nor U48571 (N_48571,N_45726,N_47447);
or U48572 (N_48572,N_45478,N_45667);
nand U48573 (N_48573,N_46479,N_46425);
and U48574 (N_48574,N_45498,N_45466);
nor U48575 (N_48575,N_46168,N_47255);
nand U48576 (N_48576,N_45082,N_45603);
xnor U48577 (N_48577,N_45859,N_46078);
and U48578 (N_48578,N_45655,N_45042);
nand U48579 (N_48579,N_46101,N_45444);
nand U48580 (N_48580,N_47437,N_45191);
nand U48581 (N_48581,N_45947,N_45820);
and U48582 (N_48582,N_46019,N_46895);
and U48583 (N_48583,N_45944,N_46456);
xor U48584 (N_48584,N_46953,N_45900);
or U48585 (N_48585,N_45501,N_46100);
and U48586 (N_48586,N_47248,N_47372);
nand U48587 (N_48587,N_46284,N_47007);
or U48588 (N_48588,N_45928,N_47261);
or U48589 (N_48589,N_46674,N_47100);
xor U48590 (N_48590,N_46329,N_46115);
nand U48591 (N_48591,N_46844,N_46909);
nor U48592 (N_48592,N_45619,N_45376);
xnor U48593 (N_48593,N_46798,N_45168);
or U48594 (N_48594,N_46921,N_45187);
nor U48595 (N_48595,N_45802,N_45695);
and U48596 (N_48596,N_47005,N_46026);
nor U48597 (N_48597,N_46543,N_46959);
nand U48598 (N_48598,N_46084,N_46645);
xor U48599 (N_48599,N_45932,N_47284);
nor U48600 (N_48600,N_45339,N_47435);
nor U48601 (N_48601,N_45785,N_47391);
or U48602 (N_48602,N_46093,N_45022);
nor U48603 (N_48603,N_47168,N_46671);
nand U48604 (N_48604,N_45034,N_47021);
and U48605 (N_48605,N_45643,N_45180);
nor U48606 (N_48606,N_45864,N_47052);
and U48607 (N_48607,N_46442,N_45407);
nand U48608 (N_48608,N_47273,N_46145);
and U48609 (N_48609,N_46777,N_45491);
nand U48610 (N_48610,N_46376,N_47195);
and U48611 (N_48611,N_46930,N_45742);
xor U48612 (N_48612,N_46976,N_45717);
xor U48613 (N_48613,N_47162,N_46214);
nand U48614 (N_48614,N_47294,N_47169);
nand U48615 (N_48615,N_45584,N_46055);
nor U48616 (N_48616,N_45452,N_47427);
nor U48617 (N_48617,N_46098,N_45389);
and U48618 (N_48618,N_46234,N_45631);
or U48619 (N_48619,N_46858,N_47417);
nor U48620 (N_48620,N_45195,N_46028);
or U48621 (N_48621,N_45188,N_47044);
and U48622 (N_48622,N_45705,N_46475);
nor U48623 (N_48623,N_45657,N_47164);
or U48624 (N_48624,N_45201,N_46885);
xor U48625 (N_48625,N_45124,N_45558);
or U48626 (N_48626,N_46577,N_46270);
nor U48627 (N_48627,N_46843,N_46327);
xor U48628 (N_48628,N_45982,N_45620);
nor U48629 (N_48629,N_45745,N_47099);
nand U48630 (N_48630,N_45704,N_46161);
nand U48631 (N_48631,N_47388,N_46106);
or U48632 (N_48632,N_45071,N_45350);
nor U48633 (N_48633,N_45536,N_45206);
or U48634 (N_48634,N_46890,N_45974);
or U48635 (N_48635,N_45276,N_47270);
or U48636 (N_48636,N_46709,N_45930);
nand U48637 (N_48637,N_45903,N_45223);
nor U48638 (N_48638,N_46302,N_45724);
or U48639 (N_48639,N_45433,N_47112);
xnor U48640 (N_48640,N_45645,N_46353);
or U48641 (N_48641,N_46900,N_46947);
nand U48642 (N_48642,N_47242,N_45611);
nor U48643 (N_48643,N_46298,N_46008);
nand U48644 (N_48644,N_45167,N_45245);
or U48645 (N_48645,N_46024,N_46605);
xor U48646 (N_48646,N_45087,N_46780);
nor U48647 (N_48647,N_47033,N_47452);
and U48648 (N_48648,N_47384,N_47431);
or U48649 (N_48649,N_46787,N_46350);
nor U48650 (N_48650,N_47398,N_45335);
nand U48651 (N_48651,N_46871,N_45709);
nor U48652 (N_48652,N_46835,N_46281);
nand U48653 (N_48653,N_45048,N_46525);
nor U48654 (N_48654,N_46881,N_45795);
and U48655 (N_48655,N_45710,N_47455);
or U48656 (N_48656,N_46524,N_46064);
and U48657 (N_48657,N_46397,N_46665);
or U48658 (N_48658,N_45829,N_45739);
nor U48659 (N_48659,N_45418,N_47166);
and U48660 (N_48660,N_45681,N_47263);
and U48661 (N_48661,N_47193,N_45164);
or U48662 (N_48662,N_47217,N_45398);
and U48663 (N_48663,N_45703,N_45438);
and U48664 (N_48664,N_45035,N_45185);
xor U48665 (N_48665,N_45081,N_46879);
and U48666 (N_48666,N_45754,N_47121);
nand U48667 (N_48667,N_45878,N_45476);
nor U48668 (N_48668,N_45467,N_47042);
or U48669 (N_48669,N_46000,N_47110);
nand U48670 (N_48670,N_46255,N_46267);
nor U48671 (N_48671,N_46171,N_47124);
and U48672 (N_48672,N_46103,N_45608);
xnor U48673 (N_48673,N_46352,N_47309);
xnor U48674 (N_48674,N_45442,N_47271);
and U48675 (N_48675,N_46133,N_46210);
nand U48676 (N_48676,N_45132,N_46330);
or U48677 (N_48677,N_45203,N_47345);
nor U48678 (N_48678,N_45237,N_46761);
xnor U48679 (N_48679,N_45131,N_46120);
and U48680 (N_48680,N_46394,N_45836);
or U48681 (N_48681,N_46589,N_46785);
and U48682 (N_48682,N_47275,N_45907);
and U48683 (N_48683,N_45148,N_45642);
and U48684 (N_48684,N_45241,N_46464);
and U48685 (N_48685,N_45015,N_47167);
and U48686 (N_48686,N_46989,N_46813);
nor U48687 (N_48687,N_46722,N_47205);
nand U48688 (N_48688,N_45755,N_47280);
and U48689 (N_48689,N_46694,N_45388);
nor U48690 (N_48690,N_45894,N_45243);
nor U48691 (N_48691,N_46288,N_47365);
and U48692 (N_48692,N_45652,N_45102);
and U48693 (N_48693,N_47106,N_46370);
nor U48694 (N_48694,N_46116,N_46821);
nor U48695 (N_48695,N_46661,N_47019);
nand U48696 (N_48696,N_45998,N_45374);
nor U48697 (N_48697,N_45254,N_45757);
and U48698 (N_48698,N_47250,N_45129);
nand U48699 (N_48699,N_46266,N_46672);
xor U48700 (N_48700,N_45120,N_46815);
nor U48701 (N_48701,N_46518,N_46862);
and U48702 (N_48702,N_46122,N_47385);
or U48703 (N_48703,N_47023,N_45431);
xor U48704 (N_48704,N_45980,N_46124);
nor U48705 (N_48705,N_47087,N_46805);
nand U48706 (N_48706,N_46057,N_46083);
nand U48707 (N_48707,N_45806,N_45649);
or U48708 (N_48708,N_45112,N_45989);
nor U48709 (N_48709,N_46621,N_45009);
nor U48710 (N_48710,N_45000,N_45564);
nand U48711 (N_48711,N_45578,N_47251);
and U48712 (N_48712,N_45450,N_45222);
nand U48713 (N_48713,N_46235,N_46721);
nand U48714 (N_48714,N_47444,N_45101);
nand U48715 (N_48715,N_45357,N_47328);
or U48716 (N_48716,N_45017,N_45173);
nor U48717 (N_48717,N_46745,N_45193);
xor U48718 (N_48718,N_46822,N_46755);
or U48719 (N_48719,N_45428,N_47373);
xnor U48720 (N_48720,N_45624,N_46348);
nand U48721 (N_48721,N_45715,N_45040);
or U48722 (N_48722,N_46540,N_45688);
nor U48723 (N_48723,N_46587,N_46789);
nand U48724 (N_48724,N_46919,N_45957);
nand U48725 (N_48725,N_45815,N_46434);
and U48726 (N_48726,N_45504,N_47148);
nand U48727 (N_48727,N_47122,N_47001);
nand U48728 (N_48728,N_45369,N_47038);
nand U48729 (N_48729,N_45123,N_46259);
and U48730 (N_48730,N_45577,N_45506);
and U48731 (N_48731,N_46905,N_46114);
nor U48732 (N_48732,N_45234,N_45663);
nand U48733 (N_48733,N_46020,N_46874);
and U48734 (N_48734,N_45707,N_46594);
nand U48735 (N_48735,N_47359,N_46945);
or U48736 (N_48736,N_45039,N_46091);
or U48737 (N_48737,N_46012,N_47003);
xnor U48738 (N_48738,N_45422,N_45779);
nand U48739 (N_48739,N_46726,N_47138);
xnor U48740 (N_48740,N_46321,N_45610);
nor U48741 (N_48741,N_46271,N_46619);
nor U48742 (N_48742,N_47376,N_47355);
nand U48743 (N_48743,N_46865,N_45001);
xnor U48744 (N_48744,N_45897,N_45938);
or U48745 (N_48745,N_47014,N_45070);
xnor U48746 (N_48746,N_45672,N_45621);
and U48747 (N_48747,N_45216,N_45420);
and U48748 (N_48748,N_47203,N_47212);
nor U48749 (N_48749,N_46176,N_45386);
and U48750 (N_48750,N_46551,N_46438);
xnor U48751 (N_48751,N_45197,N_46290);
nor U48752 (N_48752,N_46566,N_45035);
xor U48753 (N_48753,N_45967,N_45420);
xor U48754 (N_48754,N_45712,N_45398);
nand U48755 (N_48755,N_46686,N_47215);
or U48756 (N_48756,N_46178,N_45319);
nor U48757 (N_48757,N_46876,N_45110);
or U48758 (N_48758,N_46631,N_45415);
nand U48759 (N_48759,N_45116,N_46208);
nor U48760 (N_48760,N_46065,N_47397);
nand U48761 (N_48761,N_46377,N_46268);
nand U48762 (N_48762,N_45605,N_45550);
nand U48763 (N_48763,N_46568,N_47243);
or U48764 (N_48764,N_46513,N_46793);
nand U48765 (N_48765,N_45688,N_45282);
xor U48766 (N_48766,N_45293,N_45077);
nand U48767 (N_48767,N_46004,N_47212);
or U48768 (N_48768,N_45900,N_45896);
or U48769 (N_48769,N_45640,N_45738);
nor U48770 (N_48770,N_46656,N_47379);
nand U48771 (N_48771,N_47050,N_45064);
nand U48772 (N_48772,N_46478,N_45818);
or U48773 (N_48773,N_46671,N_46252);
nor U48774 (N_48774,N_46262,N_46036);
nand U48775 (N_48775,N_45531,N_45413);
and U48776 (N_48776,N_45576,N_46421);
and U48777 (N_48777,N_46797,N_47366);
and U48778 (N_48778,N_45234,N_47075);
and U48779 (N_48779,N_46222,N_45991);
nor U48780 (N_48780,N_47047,N_46150);
xor U48781 (N_48781,N_46458,N_46601);
and U48782 (N_48782,N_47193,N_45539);
or U48783 (N_48783,N_47375,N_46166);
nand U48784 (N_48784,N_47042,N_46809);
and U48785 (N_48785,N_47172,N_47443);
xnor U48786 (N_48786,N_45946,N_45295);
nand U48787 (N_48787,N_45574,N_45197);
and U48788 (N_48788,N_45248,N_47491);
xor U48789 (N_48789,N_45758,N_45428);
and U48790 (N_48790,N_46802,N_47151);
nor U48791 (N_48791,N_45253,N_47459);
nand U48792 (N_48792,N_45351,N_47185);
nor U48793 (N_48793,N_46814,N_46004);
and U48794 (N_48794,N_46535,N_45771);
or U48795 (N_48795,N_46085,N_46778);
xor U48796 (N_48796,N_47179,N_46463);
or U48797 (N_48797,N_45139,N_47472);
nand U48798 (N_48798,N_45193,N_45189);
nand U48799 (N_48799,N_45402,N_47473);
nand U48800 (N_48800,N_45936,N_47072);
nor U48801 (N_48801,N_46793,N_45508);
xor U48802 (N_48802,N_45495,N_46467);
and U48803 (N_48803,N_45745,N_45870);
nand U48804 (N_48804,N_47321,N_46289);
xnor U48805 (N_48805,N_46627,N_47363);
nor U48806 (N_48806,N_45256,N_47455);
nand U48807 (N_48807,N_47071,N_45205);
and U48808 (N_48808,N_47314,N_47145);
or U48809 (N_48809,N_45549,N_47493);
nand U48810 (N_48810,N_47457,N_45849);
or U48811 (N_48811,N_46937,N_46462);
nor U48812 (N_48812,N_45404,N_46188);
xnor U48813 (N_48813,N_45903,N_46519);
nand U48814 (N_48814,N_47423,N_47408);
and U48815 (N_48815,N_46661,N_45380);
and U48816 (N_48816,N_45338,N_46007);
and U48817 (N_48817,N_45210,N_45073);
and U48818 (N_48818,N_46225,N_45064);
or U48819 (N_48819,N_46562,N_45917);
and U48820 (N_48820,N_47318,N_45724);
or U48821 (N_48821,N_46516,N_46475);
nand U48822 (N_48822,N_47179,N_46116);
nand U48823 (N_48823,N_45876,N_45924);
xor U48824 (N_48824,N_47444,N_45490);
nand U48825 (N_48825,N_46529,N_45837);
or U48826 (N_48826,N_46522,N_45789);
and U48827 (N_48827,N_46495,N_45980);
nor U48828 (N_48828,N_46930,N_46565);
or U48829 (N_48829,N_47174,N_45158);
and U48830 (N_48830,N_46255,N_46955);
nand U48831 (N_48831,N_46074,N_45787);
xor U48832 (N_48832,N_46729,N_45858);
nor U48833 (N_48833,N_46186,N_47285);
nor U48834 (N_48834,N_46436,N_45115);
nor U48835 (N_48835,N_45908,N_45906);
xor U48836 (N_48836,N_47170,N_46239);
xnor U48837 (N_48837,N_46907,N_45473);
or U48838 (N_48838,N_45415,N_45653);
nand U48839 (N_48839,N_45708,N_45226);
nor U48840 (N_48840,N_45719,N_47021);
nor U48841 (N_48841,N_46159,N_46879);
nor U48842 (N_48842,N_47489,N_45064);
nor U48843 (N_48843,N_46071,N_47418);
and U48844 (N_48844,N_45012,N_46392);
and U48845 (N_48845,N_45966,N_46882);
and U48846 (N_48846,N_46929,N_46597);
or U48847 (N_48847,N_47386,N_45333);
nor U48848 (N_48848,N_45142,N_46630);
nor U48849 (N_48849,N_47186,N_46229);
or U48850 (N_48850,N_46030,N_46214);
xor U48851 (N_48851,N_45477,N_47141);
nand U48852 (N_48852,N_45789,N_46218);
nand U48853 (N_48853,N_46980,N_47450);
nand U48854 (N_48854,N_45634,N_46932);
or U48855 (N_48855,N_45442,N_46556);
and U48856 (N_48856,N_45586,N_46599);
nand U48857 (N_48857,N_46319,N_45247);
nor U48858 (N_48858,N_45440,N_45163);
or U48859 (N_48859,N_45830,N_47350);
nor U48860 (N_48860,N_47194,N_46419);
nor U48861 (N_48861,N_46589,N_47321);
and U48862 (N_48862,N_45042,N_46874);
and U48863 (N_48863,N_47203,N_45811);
or U48864 (N_48864,N_45647,N_46747);
or U48865 (N_48865,N_45157,N_45474);
and U48866 (N_48866,N_46033,N_47290);
xor U48867 (N_48867,N_46272,N_46002);
and U48868 (N_48868,N_47090,N_47363);
nand U48869 (N_48869,N_46072,N_47396);
nor U48870 (N_48870,N_47171,N_46172);
or U48871 (N_48871,N_46343,N_47323);
nor U48872 (N_48872,N_46316,N_46753);
or U48873 (N_48873,N_45231,N_46405);
nand U48874 (N_48874,N_47148,N_47464);
and U48875 (N_48875,N_46394,N_46232);
xnor U48876 (N_48876,N_47226,N_46643);
xnor U48877 (N_48877,N_46039,N_46007);
xnor U48878 (N_48878,N_47072,N_45978);
xor U48879 (N_48879,N_46707,N_46988);
xor U48880 (N_48880,N_45386,N_45823);
and U48881 (N_48881,N_46410,N_45898);
nor U48882 (N_48882,N_45027,N_46669);
and U48883 (N_48883,N_46376,N_45721);
or U48884 (N_48884,N_47328,N_45933);
nor U48885 (N_48885,N_46067,N_45107);
and U48886 (N_48886,N_46281,N_45535);
nand U48887 (N_48887,N_46382,N_45249);
nand U48888 (N_48888,N_46024,N_45141);
and U48889 (N_48889,N_47409,N_46442);
nand U48890 (N_48890,N_45971,N_47063);
or U48891 (N_48891,N_47424,N_46021);
and U48892 (N_48892,N_45594,N_45727);
xnor U48893 (N_48893,N_45151,N_46822);
nor U48894 (N_48894,N_47083,N_47110);
nand U48895 (N_48895,N_46121,N_46767);
nor U48896 (N_48896,N_46029,N_45527);
nor U48897 (N_48897,N_45618,N_47328);
nor U48898 (N_48898,N_45064,N_46838);
or U48899 (N_48899,N_46571,N_45076);
nand U48900 (N_48900,N_45373,N_46723);
nand U48901 (N_48901,N_47304,N_46467);
nor U48902 (N_48902,N_45835,N_46165);
and U48903 (N_48903,N_47397,N_47165);
or U48904 (N_48904,N_46544,N_47181);
nand U48905 (N_48905,N_46211,N_46291);
nor U48906 (N_48906,N_46342,N_45251);
and U48907 (N_48907,N_46755,N_46782);
nand U48908 (N_48908,N_47101,N_46648);
nor U48909 (N_48909,N_47306,N_47392);
and U48910 (N_48910,N_45000,N_45160);
nand U48911 (N_48911,N_45707,N_46068);
nor U48912 (N_48912,N_46066,N_46410);
and U48913 (N_48913,N_45628,N_47499);
or U48914 (N_48914,N_46624,N_46457);
nor U48915 (N_48915,N_45991,N_46508);
nand U48916 (N_48916,N_45860,N_46364);
and U48917 (N_48917,N_45231,N_47487);
nand U48918 (N_48918,N_45778,N_47026);
nor U48919 (N_48919,N_46373,N_45506);
or U48920 (N_48920,N_45474,N_45884);
or U48921 (N_48921,N_45528,N_45598);
or U48922 (N_48922,N_46436,N_45374);
nor U48923 (N_48923,N_45075,N_45274);
nor U48924 (N_48924,N_47034,N_46430);
nand U48925 (N_48925,N_45956,N_45345);
xor U48926 (N_48926,N_46449,N_47393);
or U48927 (N_48927,N_45773,N_47300);
nor U48928 (N_48928,N_46358,N_47336);
nor U48929 (N_48929,N_46684,N_47034);
or U48930 (N_48930,N_46778,N_45485);
or U48931 (N_48931,N_45834,N_46201);
nor U48932 (N_48932,N_47429,N_47246);
nand U48933 (N_48933,N_46278,N_45062);
or U48934 (N_48934,N_47073,N_45224);
and U48935 (N_48935,N_45377,N_45603);
nor U48936 (N_48936,N_46160,N_46482);
and U48937 (N_48937,N_45735,N_45959);
nand U48938 (N_48938,N_46577,N_46114);
nor U48939 (N_48939,N_46006,N_45230);
and U48940 (N_48940,N_45209,N_46065);
nand U48941 (N_48941,N_46916,N_46864);
nand U48942 (N_48942,N_46784,N_45401);
and U48943 (N_48943,N_47196,N_46911);
nor U48944 (N_48944,N_47475,N_47077);
nand U48945 (N_48945,N_46035,N_46378);
nor U48946 (N_48946,N_45963,N_45398);
or U48947 (N_48947,N_45789,N_46737);
nand U48948 (N_48948,N_46507,N_46255);
and U48949 (N_48949,N_46490,N_46428);
nand U48950 (N_48950,N_45253,N_45696);
nor U48951 (N_48951,N_47234,N_46766);
nor U48952 (N_48952,N_45592,N_46099);
nand U48953 (N_48953,N_47073,N_46622);
and U48954 (N_48954,N_45119,N_45189);
and U48955 (N_48955,N_46439,N_46209);
and U48956 (N_48956,N_46454,N_47047);
or U48957 (N_48957,N_47236,N_47162);
xor U48958 (N_48958,N_47013,N_45995);
xor U48959 (N_48959,N_46894,N_45687);
nor U48960 (N_48960,N_46821,N_45724);
nand U48961 (N_48961,N_45288,N_46040);
and U48962 (N_48962,N_45652,N_46298);
or U48963 (N_48963,N_47493,N_46214);
xor U48964 (N_48964,N_45107,N_46878);
nor U48965 (N_48965,N_46243,N_45337);
nor U48966 (N_48966,N_47116,N_46850);
or U48967 (N_48967,N_46491,N_45038);
and U48968 (N_48968,N_46580,N_47443);
nand U48969 (N_48969,N_46079,N_46457);
xor U48970 (N_48970,N_45523,N_45318);
nand U48971 (N_48971,N_46438,N_46818);
or U48972 (N_48972,N_47276,N_45089);
nand U48973 (N_48973,N_45893,N_47446);
nor U48974 (N_48974,N_47342,N_46359);
nand U48975 (N_48975,N_45995,N_45059);
nor U48976 (N_48976,N_45923,N_46480);
and U48977 (N_48977,N_45904,N_45268);
nand U48978 (N_48978,N_47089,N_46047);
or U48979 (N_48979,N_46104,N_47205);
nor U48980 (N_48980,N_45295,N_45552);
nand U48981 (N_48981,N_46327,N_45385);
xor U48982 (N_48982,N_46028,N_46533);
or U48983 (N_48983,N_46104,N_46543);
nand U48984 (N_48984,N_47007,N_47274);
and U48985 (N_48985,N_45472,N_46451);
nor U48986 (N_48986,N_45572,N_45659);
xor U48987 (N_48987,N_47333,N_45305);
nor U48988 (N_48988,N_46277,N_46024);
or U48989 (N_48989,N_47183,N_47468);
or U48990 (N_48990,N_46951,N_45419);
and U48991 (N_48991,N_45732,N_47401);
nor U48992 (N_48992,N_46324,N_45053);
and U48993 (N_48993,N_45985,N_46448);
or U48994 (N_48994,N_46293,N_47318);
nand U48995 (N_48995,N_45574,N_45916);
nand U48996 (N_48996,N_46455,N_46851);
nor U48997 (N_48997,N_46380,N_46152);
and U48998 (N_48998,N_45595,N_45871);
and U48999 (N_48999,N_46496,N_47018);
or U49000 (N_49000,N_45664,N_46141);
nor U49001 (N_49001,N_46401,N_45211);
nand U49002 (N_49002,N_46050,N_45839);
or U49003 (N_49003,N_45031,N_46962);
and U49004 (N_49004,N_45110,N_46516);
or U49005 (N_49005,N_46437,N_47026);
nor U49006 (N_49006,N_45133,N_46128);
nand U49007 (N_49007,N_46992,N_45269);
or U49008 (N_49008,N_46481,N_47173);
nand U49009 (N_49009,N_45491,N_46625);
nor U49010 (N_49010,N_45179,N_46562);
or U49011 (N_49011,N_46951,N_45436);
or U49012 (N_49012,N_45376,N_45146);
nor U49013 (N_49013,N_46304,N_46702);
nor U49014 (N_49014,N_46925,N_46800);
nor U49015 (N_49015,N_45569,N_46519);
nand U49016 (N_49016,N_46470,N_47445);
nand U49017 (N_49017,N_46925,N_47327);
and U49018 (N_49018,N_46177,N_45983);
xor U49019 (N_49019,N_46698,N_46192);
and U49020 (N_49020,N_46103,N_45106);
nor U49021 (N_49021,N_46454,N_47060);
or U49022 (N_49022,N_46038,N_47121);
nor U49023 (N_49023,N_47039,N_45753);
and U49024 (N_49024,N_45386,N_46632);
or U49025 (N_49025,N_47133,N_47079);
nand U49026 (N_49026,N_47480,N_46836);
or U49027 (N_49027,N_47343,N_45985);
or U49028 (N_49028,N_47093,N_46359);
or U49029 (N_49029,N_47162,N_46022);
and U49030 (N_49030,N_45177,N_45847);
nor U49031 (N_49031,N_46021,N_45950);
nor U49032 (N_49032,N_45879,N_45011);
and U49033 (N_49033,N_47495,N_45350);
or U49034 (N_49034,N_45817,N_45017);
nand U49035 (N_49035,N_46941,N_47249);
or U49036 (N_49036,N_46999,N_46671);
and U49037 (N_49037,N_45551,N_45850);
nand U49038 (N_49038,N_46617,N_47444);
nand U49039 (N_49039,N_46556,N_45099);
nand U49040 (N_49040,N_45175,N_45268);
or U49041 (N_49041,N_45185,N_46413);
or U49042 (N_49042,N_45945,N_47493);
nor U49043 (N_49043,N_45022,N_45965);
nor U49044 (N_49044,N_46594,N_45383);
or U49045 (N_49045,N_45788,N_45492);
or U49046 (N_49046,N_45563,N_45181);
and U49047 (N_49047,N_45048,N_46101);
nand U49048 (N_49048,N_46542,N_46780);
nand U49049 (N_49049,N_45897,N_46555);
nand U49050 (N_49050,N_47390,N_45123);
or U49051 (N_49051,N_46487,N_45548);
nor U49052 (N_49052,N_45582,N_46365);
or U49053 (N_49053,N_46108,N_45378);
nor U49054 (N_49054,N_46996,N_46712);
or U49055 (N_49055,N_46419,N_46522);
and U49056 (N_49056,N_46064,N_45859);
nor U49057 (N_49057,N_45265,N_45126);
nor U49058 (N_49058,N_45443,N_46449);
or U49059 (N_49059,N_47047,N_46382);
and U49060 (N_49060,N_47218,N_45602);
nor U49061 (N_49061,N_46567,N_46216);
nand U49062 (N_49062,N_45321,N_46406);
or U49063 (N_49063,N_45085,N_47319);
nor U49064 (N_49064,N_46640,N_45987);
nand U49065 (N_49065,N_45482,N_47123);
and U49066 (N_49066,N_45110,N_45474);
or U49067 (N_49067,N_45502,N_47308);
xnor U49068 (N_49068,N_47452,N_45960);
and U49069 (N_49069,N_45315,N_47359);
nor U49070 (N_49070,N_46765,N_46942);
nand U49071 (N_49071,N_45005,N_46041);
nor U49072 (N_49072,N_45717,N_47230);
nor U49073 (N_49073,N_45759,N_45114);
or U49074 (N_49074,N_47172,N_46249);
nor U49075 (N_49075,N_46698,N_47310);
nand U49076 (N_49076,N_46909,N_46727);
nand U49077 (N_49077,N_47035,N_46248);
xnor U49078 (N_49078,N_46576,N_45030);
xnor U49079 (N_49079,N_45857,N_46388);
and U49080 (N_49080,N_46039,N_45952);
nand U49081 (N_49081,N_47365,N_47308);
and U49082 (N_49082,N_46364,N_45386);
nor U49083 (N_49083,N_45709,N_45122);
or U49084 (N_49084,N_45265,N_46317);
nand U49085 (N_49085,N_46814,N_47471);
xor U49086 (N_49086,N_46342,N_46351);
nand U49087 (N_49087,N_45595,N_47189);
or U49088 (N_49088,N_46872,N_46346);
and U49089 (N_49089,N_46757,N_46065);
or U49090 (N_49090,N_46534,N_47287);
and U49091 (N_49091,N_46256,N_46263);
and U49092 (N_49092,N_45965,N_45805);
nand U49093 (N_49093,N_45811,N_45943);
nand U49094 (N_49094,N_46289,N_46170);
nand U49095 (N_49095,N_47450,N_45514);
nand U49096 (N_49096,N_45527,N_45677);
or U49097 (N_49097,N_46204,N_45586);
and U49098 (N_49098,N_46262,N_46810);
and U49099 (N_49099,N_46352,N_45300);
xnor U49100 (N_49100,N_45365,N_45946);
or U49101 (N_49101,N_47358,N_46042);
nand U49102 (N_49102,N_46358,N_47446);
nand U49103 (N_49103,N_45642,N_47384);
and U49104 (N_49104,N_46309,N_47454);
nor U49105 (N_49105,N_45390,N_45614);
xnor U49106 (N_49106,N_46506,N_45175);
xnor U49107 (N_49107,N_45605,N_45511);
nand U49108 (N_49108,N_47048,N_45938);
nand U49109 (N_49109,N_46053,N_45624);
xor U49110 (N_49110,N_47268,N_46231);
nand U49111 (N_49111,N_47408,N_45976);
and U49112 (N_49112,N_46214,N_45718);
or U49113 (N_49113,N_46508,N_47128);
nand U49114 (N_49114,N_46283,N_46258);
xor U49115 (N_49115,N_46228,N_45354);
and U49116 (N_49116,N_47298,N_45074);
and U49117 (N_49117,N_45695,N_45478);
nor U49118 (N_49118,N_45899,N_46022);
and U49119 (N_49119,N_45761,N_46289);
and U49120 (N_49120,N_45163,N_47296);
or U49121 (N_49121,N_47099,N_46289);
xor U49122 (N_49122,N_46642,N_46527);
nor U49123 (N_49123,N_46169,N_45613);
or U49124 (N_49124,N_45048,N_46489);
nand U49125 (N_49125,N_47235,N_47139);
nand U49126 (N_49126,N_47041,N_46595);
nand U49127 (N_49127,N_46832,N_46341);
nand U49128 (N_49128,N_45921,N_46566);
nand U49129 (N_49129,N_45925,N_46632);
and U49130 (N_49130,N_46619,N_45385);
nor U49131 (N_49131,N_46353,N_46767);
nor U49132 (N_49132,N_47182,N_45136);
nand U49133 (N_49133,N_45758,N_46026);
and U49134 (N_49134,N_45379,N_46637);
or U49135 (N_49135,N_45981,N_47457);
or U49136 (N_49136,N_47335,N_45898);
and U49137 (N_49137,N_45982,N_46986);
or U49138 (N_49138,N_47068,N_46924);
nor U49139 (N_49139,N_45069,N_45539);
nand U49140 (N_49140,N_45472,N_46529);
or U49141 (N_49141,N_45259,N_46006);
nand U49142 (N_49142,N_46893,N_46305);
or U49143 (N_49143,N_45221,N_45069);
and U49144 (N_49144,N_46176,N_46880);
nor U49145 (N_49145,N_46649,N_46045);
nor U49146 (N_49146,N_45454,N_45848);
nor U49147 (N_49147,N_45662,N_45212);
or U49148 (N_49148,N_45175,N_46114);
and U49149 (N_49149,N_46053,N_45143);
and U49150 (N_49150,N_45232,N_47406);
nand U49151 (N_49151,N_46600,N_47124);
and U49152 (N_49152,N_46279,N_46215);
or U49153 (N_49153,N_46421,N_45806);
and U49154 (N_49154,N_46509,N_46654);
or U49155 (N_49155,N_45600,N_45101);
or U49156 (N_49156,N_47374,N_45685);
or U49157 (N_49157,N_47441,N_45831);
or U49158 (N_49158,N_46266,N_46945);
and U49159 (N_49159,N_45480,N_45973);
nand U49160 (N_49160,N_46138,N_45765);
or U49161 (N_49161,N_45410,N_45917);
nand U49162 (N_49162,N_45121,N_45933);
nor U49163 (N_49163,N_46740,N_47311);
nand U49164 (N_49164,N_45855,N_46475);
nor U49165 (N_49165,N_45889,N_45646);
nor U49166 (N_49166,N_46672,N_46811);
nand U49167 (N_49167,N_46199,N_46542);
nor U49168 (N_49168,N_46534,N_47012);
xor U49169 (N_49169,N_47109,N_45724);
nor U49170 (N_49170,N_47355,N_46893);
nand U49171 (N_49171,N_45116,N_47190);
and U49172 (N_49172,N_47446,N_47343);
nor U49173 (N_49173,N_45293,N_47367);
xnor U49174 (N_49174,N_45196,N_47314);
and U49175 (N_49175,N_47410,N_47495);
or U49176 (N_49176,N_46597,N_46576);
nand U49177 (N_49177,N_45961,N_45543);
nor U49178 (N_49178,N_46203,N_45311);
nand U49179 (N_49179,N_46174,N_46567);
and U49180 (N_49180,N_46838,N_45269);
xor U49181 (N_49181,N_45407,N_46364);
and U49182 (N_49182,N_46455,N_47227);
nand U49183 (N_49183,N_45711,N_45881);
xor U49184 (N_49184,N_46282,N_46582);
or U49185 (N_49185,N_45378,N_47249);
nand U49186 (N_49186,N_46352,N_46900);
nor U49187 (N_49187,N_45613,N_46558);
and U49188 (N_49188,N_46299,N_46486);
nor U49189 (N_49189,N_46242,N_45769);
or U49190 (N_49190,N_46874,N_45625);
or U49191 (N_49191,N_46602,N_46367);
nor U49192 (N_49192,N_47152,N_45459);
nand U49193 (N_49193,N_45696,N_45363);
or U49194 (N_49194,N_45883,N_45182);
nor U49195 (N_49195,N_45346,N_47348);
or U49196 (N_49196,N_46644,N_47378);
or U49197 (N_49197,N_45841,N_47376);
nor U49198 (N_49198,N_45565,N_46776);
and U49199 (N_49199,N_46267,N_45821);
and U49200 (N_49200,N_45994,N_46976);
nand U49201 (N_49201,N_46489,N_47125);
nand U49202 (N_49202,N_46688,N_47494);
nor U49203 (N_49203,N_46732,N_47277);
nor U49204 (N_49204,N_46355,N_45159);
xnor U49205 (N_49205,N_45902,N_46576);
or U49206 (N_49206,N_46159,N_45838);
nand U49207 (N_49207,N_46448,N_47214);
nand U49208 (N_49208,N_46420,N_45640);
or U49209 (N_49209,N_46652,N_47298);
or U49210 (N_49210,N_46043,N_47218);
and U49211 (N_49211,N_46834,N_46441);
nor U49212 (N_49212,N_46700,N_45911);
or U49213 (N_49213,N_47248,N_45205);
or U49214 (N_49214,N_47280,N_46196);
nor U49215 (N_49215,N_46489,N_45676);
and U49216 (N_49216,N_47272,N_46630);
xnor U49217 (N_49217,N_46574,N_45026);
nand U49218 (N_49218,N_45548,N_45267);
nand U49219 (N_49219,N_46012,N_46450);
nand U49220 (N_49220,N_45531,N_46594);
nor U49221 (N_49221,N_47470,N_45504);
or U49222 (N_49222,N_45524,N_47474);
nand U49223 (N_49223,N_46573,N_45962);
nor U49224 (N_49224,N_45540,N_45771);
nand U49225 (N_49225,N_46878,N_45242);
nand U49226 (N_49226,N_45002,N_47202);
nand U49227 (N_49227,N_46931,N_46933);
nand U49228 (N_49228,N_45093,N_46281);
nand U49229 (N_49229,N_47004,N_45635);
or U49230 (N_49230,N_47249,N_45747);
and U49231 (N_49231,N_46383,N_46113);
nand U49232 (N_49232,N_46432,N_47472);
xor U49233 (N_49233,N_45603,N_45791);
nand U49234 (N_49234,N_45297,N_45307);
nand U49235 (N_49235,N_45665,N_47271);
xnor U49236 (N_49236,N_46217,N_46425);
nor U49237 (N_49237,N_45757,N_46260);
and U49238 (N_49238,N_47268,N_46523);
and U49239 (N_49239,N_46169,N_46050);
and U49240 (N_49240,N_46682,N_46665);
nor U49241 (N_49241,N_46070,N_45545);
nand U49242 (N_49242,N_46313,N_45819);
nor U49243 (N_49243,N_47221,N_47298);
and U49244 (N_49244,N_47056,N_45083);
and U49245 (N_49245,N_46474,N_46303);
nor U49246 (N_49246,N_46691,N_46224);
and U49247 (N_49247,N_47337,N_47218);
or U49248 (N_49248,N_45422,N_46011);
or U49249 (N_49249,N_47309,N_47171);
and U49250 (N_49250,N_46712,N_46614);
nor U49251 (N_49251,N_45535,N_45500);
xnor U49252 (N_49252,N_45506,N_46665);
nor U49253 (N_49253,N_45406,N_46152);
nor U49254 (N_49254,N_47157,N_46057);
nand U49255 (N_49255,N_45853,N_45376);
or U49256 (N_49256,N_45728,N_45799);
and U49257 (N_49257,N_47104,N_46885);
nand U49258 (N_49258,N_46735,N_45896);
nand U49259 (N_49259,N_45164,N_46336);
nand U49260 (N_49260,N_45712,N_45617);
and U49261 (N_49261,N_46171,N_47210);
nor U49262 (N_49262,N_47120,N_45121);
or U49263 (N_49263,N_45358,N_46140);
and U49264 (N_49264,N_45286,N_46246);
or U49265 (N_49265,N_46061,N_47495);
or U49266 (N_49266,N_46874,N_46960);
or U49267 (N_49267,N_47044,N_45474);
or U49268 (N_49268,N_47338,N_46307);
and U49269 (N_49269,N_45947,N_46206);
nand U49270 (N_49270,N_45637,N_47064);
nand U49271 (N_49271,N_45086,N_46238);
nand U49272 (N_49272,N_47307,N_46546);
nand U49273 (N_49273,N_46455,N_45332);
nor U49274 (N_49274,N_46384,N_45950);
nor U49275 (N_49275,N_46467,N_46902);
nor U49276 (N_49276,N_45426,N_46455);
nand U49277 (N_49277,N_47206,N_45700);
and U49278 (N_49278,N_46136,N_45217);
nor U49279 (N_49279,N_45690,N_46234);
nor U49280 (N_49280,N_47372,N_45960);
and U49281 (N_49281,N_46208,N_45861);
nand U49282 (N_49282,N_45379,N_45162);
or U49283 (N_49283,N_47417,N_45183);
nand U49284 (N_49284,N_46421,N_45981);
nor U49285 (N_49285,N_45811,N_45739);
nor U49286 (N_49286,N_47408,N_46839);
and U49287 (N_49287,N_46611,N_45885);
nor U49288 (N_49288,N_46040,N_45441);
nor U49289 (N_49289,N_45870,N_46848);
and U49290 (N_49290,N_45512,N_45731);
and U49291 (N_49291,N_46089,N_47307);
nor U49292 (N_49292,N_46244,N_47101);
xnor U49293 (N_49293,N_45016,N_46014);
and U49294 (N_49294,N_45181,N_45410);
nand U49295 (N_49295,N_46946,N_47246);
nor U49296 (N_49296,N_46964,N_45068);
and U49297 (N_49297,N_46214,N_46643);
nor U49298 (N_49298,N_46400,N_46967);
xnor U49299 (N_49299,N_46690,N_45600);
and U49300 (N_49300,N_46638,N_46089);
nand U49301 (N_49301,N_46572,N_47091);
nor U49302 (N_49302,N_45902,N_46205);
and U49303 (N_49303,N_47457,N_46282);
or U49304 (N_49304,N_46912,N_45346);
nand U49305 (N_49305,N_45388,N_46510);
or U49306 (N_49306,N_45213,N_45799);
or U49307 (N_49307,N_47496,N_46231);
or U49308 (N_49308,N_45459,N_47328);
nor U49309 (N_49309,N_47157,N_45149);
nand U49310 (N_49310,N_45104,N_46987);
nand U49311 (N_49311,N_47466,N_45085);
nand U49312 (N_49312,N_46867,N_46195);
nor U49313 (N_49313,N_46717,N_47394);
or U49314 (N_49314,N_46411,N_45187);
and U49315 (N_49315,N_46500,N_46356);
or U49316 (N_49316,N_45650,N_46088);
nand U49317 (N_49317,N_45404,N_47460);
nand U49318 (N_49318,N_47110,N_45486);
xor U49319 (N_49319,N_46774,N_46770);
nor U49320 (N_49320,N_46579,N_45646);
nor U49321 (N_49321,N_46161,N_46818);
and U49322 (N_49322,N_46825,N_46854);
or U49323 (N_49323,N_46019,N_45688);
and U49324 (N_49324,N_46644,N_45181);
or U49325 (N_49325,N_47382,N_46260);
nor U49326 (N_49326,N_45522,N_45797);
nor U49327 (N_49327,N_46262,N_46688);
or U49328 (N_49328,N_46255,N_45815);
and U49329 (N_49329,N_45886,N_45362);
xor U49330 (N_49330,N_45443,N_46619);
and U49331 (N_49331,N_45855,N_46525);
xor U49332 (N_49332,N_46133,N_47490);
xnor U49333 (N_49333,N_46073,N_45903);
or U49334 (N_49334,N_47376,N_47006);
nand U49335 (N_49335,N_46259,N_45285);
nand U49336 (N_49336,N_45098,N_47103);
or U49337 (N_49337,N_47118,N_46745);
xor U49338 (N_49338,N_46538,N_45708);
nand U49339 (N_49339,N_46673,N_47450);
and U49340 (N_49340,N_46289,N_45753);
nor U49341 (N_49341,N_45034,N_47115);
or U49342 (N_49342,N_46966,N_46164);
or U49343 (N_49343,N_47161,N_46061);
nand U49344 (N_49344,N_46794,N_45005);
nand U49345 (N_49345,N_47357,N_46016);
or U49346 (N_49346,N_45483,N_45271);
and U49347 (N_49347,N_46134,N_46572);
nand U49348 (N_49348,N_46850,N_46497);
or U49349 (N_49349,N_46557,N_45024);
xnor U49350 (N_49350,N_47488,N_45425);
nor U49351 (N_49351,N_46979,N_45327);
xnor U49352 (N_49352,N_46751,N_46451);
or U49353 (N_49353,N_45085,N_45777);
nand U49354 (N_49354,N_46617,N_46989);
or U49355 (N_49355,N_45539,N_45349);
and U49356 (N_49356,N_47093,N_47324);
and U49357 (N_49357,N_46409,N_45109);
nor U49358 (N_49358,N_46806,N_45632);
nor U49359 (N_49359,N_46357,N_45845);
and U49360 (N_49360,N_46765,N_45332);
or U49361 (N_49361,N_45424,N_45404);
nor U49362 (N_49362,N_46266,N_45248);
nor U49363 (N_49363,N_46256,N_45316);
and U49364 (N_49364,N_46864,N_47344);
or U49365 (N_49365,N_46283,N_46973);
nand U49366 (N_49366,N_46179,N_45185);
nor U49367 (N_49367,N_45700,N_45503);
nand U49368 (N_49368,N_47464,N_47370);
nor U49369 (N_49369,N_46129,N_45931);
or U49370 (N_49370,N_47226,N_46640);
or U49371 (N_49371,N_46257,N_45969);
nor U49372 (N_49372,N_47216,N_45196);
and U49373 (N_49373,N_45998,N_45173);
nor U49374 (N_49374,N_46497,N_46533);
or U49375 (N_49375,N_46274,N_46528);
nand U49376 (N_49376,N_47365,N_45046);
xor U49377 (N_49377,N_45812,N_45448);
xnor U49378 (N_49378,N_46244,N_46557);
and U49379 (N_49379,N_46862,N_46781);
and U49380 (N_49380,N_47327,N_46619);
xor U49381 (N_49381,N_46537,N_46626);
nand U49382 (N_49382,N_47002,N_45947);
nand U49383 (N_49383,N_46847,N_47310);
xor U49384 (N_49384,N_46028,N_46214);
nor U49385 (N_49385,N_45394,N_45829);
or U49386 (N_49386,N_46230,N_47065);
and U49387 (N_49387,N_45708,N_46591);
and U49388 (N_49388,N_46797,N_47041);
and U49389 (N_49389,N_45899,N_46566);
nand U49390 (N_49390,N_45312,N_46572);
or U49391 (N_49391,N_46117,N_46112);
nand U49392 (N_49392,N_45859,N_45789);
nand U49393 (N_49393,N_45942,N_47473);
and U49394 (N_49394,N_45616,N_45222);
nor U49395 (N_49395,N_45033,N_47039);
nand U49396 (N_49396,N_46674,N_45102);
xnor U49397 (N_49397,N_46480,N_47333);
or U49398 (N_49398,N_47482,N_45245);
and U49399 (N_49399,N_45795,N_46734);
or U49400 (N_49400,N_47168,N_45522);
nand U49401 (N_49401,N_45393,N_46870);
nor U49402 (N_49402,N_47448,N_45793);
or U49403 (N_49403,N_45489,N_47134);
or U49404 (N_49404,N_46866,N_45178);
nand U49405 (N_49405,N_46617,N_47367);
or U49406 (N_49406,N_46711,N_45086);
xor U49407 (N_49407,N_46646,N_47390);
and U49408 (N_49408,N_45496,N_46080);
xnor U49409 (N_49409,N_45887,N_46768);
nor U49410 (N_49410,N_47446,N_47157);
or U49411 (N_49411,N_47183,N_47184);
or U49412 (N_49412,N_47463,N_47444);
xor U49413 (N_49413,N_47339,N_46855);
nor U49414 (N_49414,N_45578,N_45220);
or U49415 (N_49415,N_46852,N_45979);
xnor U49416 (N_49416,N_46445,N_45043);
or U49417 (N_49417,N_46833,N_45220);
nand U49418 (N_49418,N_47051,N_46333);
xnor U49419 (N_49419,N_45123,N_45243);
nor U49420 (N_49420,N_46386,N_45188);
xor U49421 (N_49421,N_45432,N_46430);
xor U49422 (N_49422,N_46354,N_45412);
and U49423 (N_49423,N_46367,N_45668);
nor U49424 (N_49424,N_46859,N_46889);
and U49425 (N_49425,N_46663,N_46672);
nor U49426 (N_49426,N_46967,N_46894);
nor U49427 (N_49427,N_46353,N_46203);
xor U49428 (N_49428,N_45432,N_47145);
or U49429 (N_49429,N_45176,N_47373);
and U49430 (N_49430,N_45452,N_46521);
nor U49431 (N_49431,N_46145,N_46423);
and U49432 (N_49432,N_47407,N_47095);
nand U49433 (N_49433,N_45855,N_45200);
nand U49434 (N_49434,N_46220,N_47338);
nand U49435 (N_49435,N_46047,N_46553);
nand U49436 (N_49436,N_45141,N_46372);
nor U49437 (N_49437,N_46064,N_45787);
or U49438 (N_49438,N_47363,N_45998);
nand U49439 (N_49439,N_47295,N_45112);
xnor U49440 (N_49440,N_46746,N_45947);
nor U49441 (N_49441,N_46122,N_45057);
or U49442 (N_49442,N_45736,N_45668);
nor U49443 (N_49443,N_45129,N_47082);
and U49444 (N_49444,N_46762,N_47169);
nor U49445 (N_49445,N_45954,N_45209);
nand U49446 (N_49446,N_47175,N_46183);
nor U49447 (N_49447,N_46313,N_46693);
xnor U49448 (N_49448,N_45093,N_46507);
and U49449 (N_49449,N_45421,N_46604);
and U49450 (N_49450,N_45930,N_46147);
and U49451 (N_49451,N_45545,N_45166);
nand U49452 (N_49452,N_47055,N_46570);
or U49453 (N_49453,N_46317,N_45923);
xnor U49454 (N_49454,N_46246,N_45495);
nand U49455 (N_49455,N_45851,N_46144);
nor U49456 (N_49456,N_46317,N_47252);
nand U49457 (N_49457,N_46301,N_47257);
nand U49458 (N_49458,N_46795,N_45517);
and U49459 (N_49459,N_45192,N_45443);
or U49460 (N_49460,N_47117,N_45910);
nor U49461 (N_49461,N_45953,N_45705);
nor U49462 (N_49462,N_47111,N_46458);
or U49463 (N_49463,N_47426,N_47488);
and U49464 (N_49464,N_46084,N_47094);
nand U49465 (N_49465,N_46647,N_47180);
nand U49466 (N_49466,N_46834,N_45632);
and U49467 (N_49467,N_46868,N_46346);
nor U49468 (N_49468,N_45397,N_46525);
nand U49469 (N_49469,N_47251,N_45417);
nand U49470 (N_49470,N_45482,N_47033);
and U49471 (N_49471,N_45668,N_45253);
nor U49472 (N_49472,N_46316,N_46364);
or U49473 (N_49473,N_46484,N_46261);
nor U49474 (N_49474,N_45165,N_46616);
nand U49475 (N_49475,N_46347,N_46112);
or U49476 (N_49476,N_46644,N_45384);
nand U49477 (N_49477,N_45073,N_47416);
nand U49478 (N_49478,N_46526,N_45420);
or U49479 (N_49479,N_47397,N_47004);
nor U49480 (N_49480,N_45255,N_45100);
nor U49481 (N_49481,N_47322,N_45470);
and U49482 (N_49482,N_45605,N_45487);
nor U49483 (N_49483,N_47110,N_45655);
or U49484 (N_49484,N_45005,N_45361);
nor U49485 (N_49485,N_45668,N_45577);
nand U49486 (N_49486,N_45990,N_45196);
xor U49487 (N_49487,N_46277,N_45126);
and U49488 (N_49488,N_45708,N_46098);
and U49489 (N_49489,N_47235,N_45436);
nor U49490 (N_49490,N_46389,N_46653);
or U49491 (N_49491,N_46307,N_46700);
nand U49492 (N_49492,N_46998,N_46734);
nor U49493 (N_49493,N_46532,N_45482);
nor U49494 (N_49494,N_45697,N_47465);
nor U49495 (N_49495,N_45510,N_45246);
xor U49496 (N_49496,N_46643,N_46078);
or U49497 (N_49497,N_47014,N_47106);
or U49498 (N_49498,N_45858,N_47031);
and U49499 (N_49499,N_46688,N_46222);
and U49500 (N_49500,N_47308,N_47444);
and U49501 (N_49501,N_47017,N_46883);
and U49502 (N_49502,N_46842,N_45658);
or U49503 (N_49503,N_45898,N_47101);
nand U49504 (N_49504,N_46406,N_45089);
xor U49505 (N_49505,N_47459,N_46483);
nor U49506 (N_49506,N_45252,N_45102);
or U49507 (N_49507,N_45069,N_46693);
nor U49508 (N_49508,N_45989,N_46913);
or U49509 (N_49509,N_47420,N_45555);
nor U49510 (N_49510,N_46875,N_45974);
nor U49511 (N_49511,N_46015,N_47476);
or U49512 (N_49512,N_47045,N_46317);
or U49513 (N_49513,N_45953,N_47193);
nor U49514 (N_49514,N_47293,N_47333);
nor U49515 (N_49515,N_47140,N_46906);
nor U49516 (N_49516,N_45131,N_45187);
or U49517 (N_49517,N_46199,N_46038);
xor U49518 (N_49518,N_46504,N_46158);
and U49519 (N_49519,N_47080,N_46188);
nand U49520 (N_49520,N_45947,N_46667);
and U49521 (N_49521,N_45055,N_46180);
nor U49522 (N_49522,N_46379,N_45820);
or U49523 (N_49523,N_46945,N_47262);
and U49524 (N_49524,N_46892,N_47008);
nand U49525 (N_49525,N_46191,N_46702);
nor U49526 (N_49526,N_45300,N_47190);
xor U49527 (N_49527,N_47382,N_46834);
nand U49528 (N_49528,N_45485,N_45298);
or U49529 (N_49529,N_47302,N_47368);
nor U49530 (N_49530,N_46508,N_47297);
or U49531 (N_49531,N_45252,N_45074);
nor U49532 (N_49532,N_45121,N_45608);
nand U49533 (N_49533,N_46491,N_45644);
nand U49534 (N_49534,N_46343,N_47419);
nor U49535 (N_49535,N_46165,N_46208);
nand U49536 (N_49536,N_46514,N_45768);
nand U49537 (N_49537,N_47172,N_46433);
nor U49538 (N_49538,N_45421,N_46289);
nand U49539 (N_49539,N_47024,N_45079);
and U49540 (N_49540,N_46117,N_46807);
nand U49541 (N_49541,N_46132,N_46353);
nand U49542 (N_49542,N_46796,N_47284);
or U49543 (N_49543,N_47114,N_47430);
and U49544 (N_49544,N_47329,N_47420);
nand U49545 (N_49545,N_45099,N_47354);
and U49546 (N_49546,N_46018,N_45876);
nand U49547 (N_49547,N_47451,N_46874);
or U49548 (N_49548,N_45981,N_47052);
or U49549 (N_49549,N_47009,N_45685);
nor U49550 (N_49550,N_45779,N_46732);
nand U49551 (N_49551,N_46542,N_46768);
nor U49552 (N_49552,N_46274,N_46600);
nor U49553 (N_49553,N_47179,N_46598);
or U49554 (N_49554,N_45413,N_47439);
nor U49555 (N_49555,N_47001,N_45872);
xnor U49556 (N_49556,N_47206,N_45531);
nand U49557 (N_49557,N_46469,N_46831);
nand U49558 (N_49558,N_46169,N_46398);
and U49559 (N_49559,N_47108,N_47462);
and U49560 (N_49560,N_46570,N_46490);
or U49561 (N_49561,N_45403,N_46609);
and U49562 (N_49562,N_46397,N_47212);
and U49563 (N_49563,N_46961,N_45078);
or U49564 (N_49564,N_47102,N_47159);
nand U49565 (N_49565,N_47475,N_45824);
and U49566 (N_49566,N_47313,N_46587);
nand U49567 (N_49567,N_45463,N_46087);
xor U49568 (N_49568,N_45913,N_46529);
or U49569 (N_49569,N_46549,N_45986);
nand U49570 (N_49570,N_47475,N_46652);
nor U49571 (N_49571,N_47460,N_45907);
xor U49572 (N_49572,N_47042,N_47326);
nor U49573 (N_49573,N_46998,N_45569);
and U49574 (N_49574,N_45898,N_45993);
and U49575 (N_49575,N_46770,N_45659);
and U49576 (N_49576,N_45367,N_46260);
and U49577 (N_49577,N_46234,N_45463);
and U49578 (N_49578,N_45582,N_46583);
or U49579 (N_49579,N_45445,N_46100);
and U49580 (N_49580,N_46953,N_47058);
nor U49581 (N_49581,N_45598,N_46269);
nand U49582 (N_49582,N_46586,N_46218);
nand U49583 (N_49583,N_47494,N_45046);
xnor U49584 (N_49584,N_45322,N_46000);
nor U49585 (N_49585,N_45732,N_47194);
xnor U49586 (N_49586,N_45852,N_47440);
and U49587 (N_49587,N_45084,N_46658);
or U49588 (N_49588,N_45702,N_47113);
or U49589 (N_49589,N_45187,N_46569);
or U49590 (N_49590,N_47131,N_45440);
xnor U49591 (N_49591,N_45205,N_47240);
and U49592 (N_49592,N_47068,N_45650);
nor U49593 (N_49593,N_45444,N_46397);
nor U49594 (N_49594,N_46405,N_46371);
nand U49595 (N_49595,N_46837,N_45415);
nor U49596 (N_49596,N_46581,N_46570);
or U49597 (N_49597,N_45322,N_46061);
and U49598 (N_49598,N_45855,N_47098);
and U49599 (N_49599,N_46901,N_46209);
nand U49600 (N_49600,N_47331,N_47174);
nand U49601 (N_49601,N_46405,N_46223);
xor U49602 (N_49602,N_46609,N_47475);
xor U49603 (N_49603,N_45465,N_45598);
xnor U49604 (N_49604,N_45265,N_47019);
nand U49605 (N_49605,N_46581,N_45661);
or U49606 (N_49606,N_45996,N_47094);
nor U49607 (N_49607,N_45058,N_46210);
or U49608 (N_49608,N_46441,N_45195);
or U49609 (N_49609,N_45761,N_47052);
nand U49610 (N_49610,N_45305,N_45027);
nor U49611 (N_49611,N_47389,N_45125);
and U49612 (N_49612,N_46268,N_46092);
or U49613 (N_49613,N_45142,N_46619);
or U49614 (N_49614,N_46511,N_47227);
and U49615 (N_49615,N_46767,N_47469);
and U49616 (N_49616,N_46962,N_46531);
or U49617 (N_49617,N_46059,N_47074);
nand U49618 (N_49618,N_45221,N_46585);
or U49619 (N_49619,N_46443,N_46590);
nor U49620 (N_49620,N_47284,N_45039);
and U49621 (N_49621,N_45310,N_46008);
nor U49622 (N_49622,N_46937,N_47491);
nor U49623 (N_49623,N_45510,N_45273);
and U49624 (N_49624,N_46949,N_46908);
nor U49625 (N_49625,N_45510,N_45270);
nor U49626 (N_49626,N_45221,N_45697);
nand U49627 (N_49627,N_47380,N_45224);
nor U49628 (N_49628,N_45871,N_46339);
or U49629 (N_49629,N_45169,N_45541);
or U49630 (N_49630,N_47042,N_47470);
nor U49631 (N_49631,N_45056,N_45299);
nand U49632 (N_49632,N_46111,N_45411);
nand U49633 (N_49633,N_47013,N_47125);
or U49634 (N_49634,N_45265,N_46195);
and U49635 (N_49635,N_47428,N_47394);
nor U49636 (N_49636,N_47176,N_45476);
or U49637 (N_49637,N_47381,N_45261);
nor U49638 (N_49638,N_45303,N_47154);
nor U49639 (N_49639,N_46121,N_46739);
and U49640 (N_49640,N_46788,N_47358);
or U49641 (N_49641,N_45202,N_45986);
xor U49642 (N_49642,N_45630,N_45012);
nor U49643 (N_49643,N_46037,N_47294);
nor U49644 (N_49644,N_46178,N_45903);
xor U49645 (N_49645,N_47137,N_47065);
nor U49646 (N_49646,N_45834,N_46919);
or U49647 (N_49647,N_47491,N_45287);
and U49648 (N_49648,N_47288,N_46492);
or U49649 (N_49649,N_45150,N_46016);
nor U49650 (N_49650,N_47255,N_47357);
or U49651 (N_49651,N_45188,N_45937);
and U49652 (N_49652,N_47100,N_45817);
or U49653 (N_49653,N_46840,N_45793);
nor U49654 (N_49654,N_47048,N_45139);
nor U49655 (N_49655,N_47131,N_45499);
or U49656 (N_49656,N_47190,N_47193);
or U49657 (N_49657,N_47431,N_45790);
and U49658 (N_49658,N_46714,N_45399);
nor U49659 (N_49659,N_47005,N_47229);
nand U49660 (N_49660,N_47467,N_45107);
nor U49661 (N_49661,N_46473,N_45748);
and U49662 (N_49662,N_45510,N_45924);
or U49663 (N_49663,N_46046,N_46555);
nand U49664 (N_49664,N_47329,N_45792);
and U49665 (N_49665,N_47334,N_47060);
and U49666 (N_49666,N_45356,N_45024);
nand U49667 (N_49667,N_45038,N_47201);
xnor U49668 (N_49668,N_46552,N_46722);
and U49669 (N_49669,N_46815,N_47020);
and U49670 (N_49670,N_46814,N_45440);
nor U49671 (N_49671,N_46179,N_46205);
nor U49672 (N_49672,N_46844,N_45608);
xnor U49673 (N_49673,N_46753,N_46213);
and U49674 (N_49674,N_45448,N_45936);
or U49675 (N_49675,N_45889,N_46138);
nor U49676 (N_49676,N_46586,N_45742);
nor U49677 (N_49677,N_46803,N_47489);
nand U49678 (N_49678,N_47123,N_46655);
xor U49679 (N_49679,N_47171,N_46754);
or U49680 (N_49680,N_47297,N_45037);
nand U49681 (N_49681,N_45775,N_46467);
or U49682 (N_49682,N_45876,N_46397);
and U49683 (N_49683,N_45218,N_47108);
nand U49684 (N_49684,N_47382,N_46391);
xnor U49685 (N_49685,N_46776,N_45686);
or U49686 (N_49686,N_45036,N_46013);
nand U49687 (N_49687,N_46238,N_45563);
or U49688 (N_49688,N_47299,N_45038);
nand U49689 (N_49689,N_46807,N_46219);
and U49690 (N_49690,N_46599,N_45516);
nand U49691 (N_49691,N_45461,N_47011);
nand U49692 (N_49692,N_46633,N_45148);
nand U49693 (N_49693,N_47263,N_47291);
xor U49694 (N_49694,N_45307,N_45545);
nand U49695 (N_49695,N_46213,N_46324);
nor U49696 (N_49696,N_46195,N_47097);
nor U49697 (N_49697,N_46428,N_45844);
nor U49698 (N_49698,N_47405,N_46031);
nand U49699 (N_49699,N_47368,N_45284);
xnor U49700 (N_49700,N_45483,N_46720);
nor U49701 (N_49701,N_45712,N_45304);
or U49702 (N_49702,N_47110,N_47481);
and U49703 (N_49703,N_45800,N_47373);
xnor U49704 (N_49704,N_45930,N_47178);
and U49705 (N_49705,N_46661,N_47321);
or U49706 (N_49706,N_46890,N_46831);
xor U49707 (N_49707,N_45438,N_47280);
nor U49708 (N_49708,N_46287,N_46140);
nand U49709 (N_49709,N_46937,N_47439);
nor U49710 (N_49710,N_46654,N_46149);
nand U49711 (N_49711,N_47206,N_45544);
nand U49712 (N_49712,N_45386,N_46964);
or U49713 (N_49713,N_47439,N_46730);
and U49714 (N_49714,N_46344,N_46405);
nand U49715 (N_49715,N_47479,N_47004);
or U49716 (N_49716,N_45933,N_46982);
and U49717 (N_49717,N_46026,N_45271);
nor U49718 (N_49718,N_45645,N_47316);
or U49719 (N_49719,N_46532,N_45149);
nand U49720 (N_49720,N_47306,N_46919);
nand U49721 (N_49721,N_46122,N_45815);
xnor U49722 (N_49722,N_46773,N_45132);
nor U49723 (N_49723,N_46690,N_46484);
and U49724 (N_49724,N_45320,N_47434);
or U49725 (N_49725,N_46159,N_45984);
nor U49726 (N_49726,N_45442,N_47296);
nor U49727 (N_49727,N_46364,N_45426);
nand U49728 (N_49728,N_45925,N_47106);
nand U49729 (N_49729,N_47223,N_45416);
or U49730 (N_49730,N_45781,N_45259);
and U49731 (N_49731,N_46542,N_45427);
xor U49732 (N_49732,N_46303,N_46255);
or U49733 (N_49733,N_46165,N_45087);
nand U49734 (N_49734,N_47265,N_45810);
xor U49735 (N_49735,N_45329,N_45639);
nor U49736 (N_49736,N_45702,N_46492);
nor U49737 (N_49737,N_46043,N_45141);
or U49738 (N_49738,N_45326,N_46629);
and U49739 (N_49739,N_47064,N_45144);
and U49740 (N_49740,N_45426,N_46195);
or U49741 (N_49741,N_45145,N_47001);
and U49742 (N_49742,N_45757,N_45188);
nor U49743 (N_49743,N_46906,N_47226);
nand U49744 (N_49744,N_46012,N_45345);
and U49745 (N_49745,N_46572,N_47287);
nand U49746 (N_49746,N_45510,N_46227);
or U49747 (N_49747,N_45835,N_46119);
and U49748 (N_49748,N_46292,N_47116);
or U49749 (N_49749,N_46960,N_45118);
nand U49750 (N_49750,N_47154,N_45642);
and U49751 (N_49751,N_45949,N_46322);
and U49752 (N_49752,N_46538,N_45801);
xnor U49753 (N_49753,N_46177,N_45641);
nor U49754 (N_49754,N_47039,N_46360);
and U49755 (N_49755,N_46482,N_45923);
nand U49756 (N_49756,N_46923,N_45407);
nand U49757 (N_49757,N_46139,N_46942);
nand U49758 (N_49758,N_47343,N_46261);
nand U49759 (N_49759,N_46362,N_45705);
and U49760 (N_49760,N_45273,N_45487);
or U49761 (N_49761,N_45271,N_45478);
nand U49762 (N_49762,N_45602,N_47292);
xnor U49763 (N_49763,N_45314,N_45192);
nor U49764 (N_49764,N_45911,N_45971);
nand U49765 (N_49765,N_46938,N_45380);
nand U49766 (N_49766,N_46612,N_45890);
or U49767 (N_49767,N_47153,N_46339);
nor U49768 (N_49768,N_46351,N_45416);
nor U49769 (N_49769,N_45764,N_45111);
and U49770 (N_49770,N_47131,N_46739);
or U49771 (N_49771,N_46302,N_46468);
or U49772 (N_49772,N_46248,N_45045);
or U49773 (N_49773,N_47293,N_46703);
and U49774 (N_49774,N_45501,N_47141);
xnor U49775 (N_49775,N_45118,N_47362);
and U49776 (N_49776,N_46056,N_46146);
and U49777 (N_49777,N_46018,N_45797);
and U49778 (N_49778,N_45922,N_45445);
nor U49779 (N_49779,N_46901,N_46555);
and U49780 (N_49780,N_47047,N_46894);
nor U49781 (N_49781,N_46972,N_45238);
nor U49782 (N_49782,N_46070,N_46430);
or U49783 (N_49783,N_46893,N_46929);
xnor U49784 (N_49784,N_45282,N_46432);
nor U49785 (N_49785,N_45343,N_45136);
xor U49786 (N_49786,N_45840,N_45136);
nor U49787 (N_49787,N_46535,N_46132);
nand U49788 (N_49788,N_45209,N_45212);
or U49789 (N_49789,N_46702,N_46550);
and U49790 (N_49790,N_45424,N_46635);
or U49791 (N_49791,N_45656,N_45070);
and U49792 (N_49792,N_46112,N_45316);
nor U49793 (N_49793,N_46937,N_45387);
nor U49794 (N_49794,N_45722,N_45066);
nand U49795 (N_49795,N_45982,N_45759);
xor U49796 (N_49796,N_46415,N_47059);
or U49797 (N_49797,N_46637,N_46508);
nand U49798 (N_49798,N_46260,N_47440);
nand U49799 (N_49799,N_46673,N_45398);
nand U49800 (N_49800,N_45899,N_47334);
or U49801 (N_49801,N_46026,N_47456);
nor U49802 (N_49802,N_45104,N_47176);
nor U49803 (N_49803,N_46493,N_45179);
nand U49804 (N_49804,N_45846,N_47270);
or U49805 (N_49805,N_46030,N_45879);
and U49806 (N_49806,N_47166,N_45350);
and U49807 (N_49807,N_45486,N_47094);
and U49808 (N_49808,N_45157,N_47273);
and U49809 (N_49809,N_46082,N_45369);
or U49810 (N_49810,N_47457,N_45451);
nor U49811 (N_49811,N_46718,N_45401);
and U49812 (N_49812,N_45472,N_45182);
nor U49813 (N_49813,N_46544,N_45049);
or U49814 (N_49814,N_45769,N_46349);
xnor U49815 (N_49815,N_45468,N_45469);
nor U49816 (N_49816,N_45889,N_46590);
and U49817 (N_49817,N_46428,N_45358);
xnor U49818 (N_49818,N_46683,N_45649);
nor U49819 (N_49819,N_45722,N_46964);
and U49820 (N_49820,N_45230,N_46298);
and U49821 (N_49821,N_45660,N_47432);
or U49822 (N_49822,N_47119,N_46176);
and U49823 (N_49823,N_46464,N_47215);
or U49824 (N_49824,N_46329,N_45104);
nand U49825 (N_49825,N_47484,N_46940);
and U49826 (N_49826,N_46555,N_45824);
nand U49827 (N_49827,N_45913,N_46101);
xnor U49828 (N_49828,N_45614,N_46761);
or U49829 (N_49829,N_45281,N_45776);
xor U49830 (N_49830,N_47385,N_45970);
and U49831 (N_49831,N_45398,N_45940);
or U49832 (N_49832,N_45869,N_45623);
and U49833 (N_49833,N_45100,N_46993);
and U49834 (N_49834,N_46330,N_46329);
nand U49835 (N_49835,N_47427,N_45072);
nor U49836 (N_49836,N_45906,N_46751);
nand U49837 (N_49837,N_45492,N_47309);
nand U49838 (N_49838,N_45112,N_45968);
xor U49839 (N_49839,N_45416,N_46840);
or U49840 (N_49840,N_47031,N_47198);
and U49841 (N_49841,N_45409,N_45392);
or U49842 (N_49842,N_45039,N_46228);
nor U49843 (N_49843,N_46775,N_45617);
nor U49844 (N_49844,N_45433,N_46181);
and U49845 (N_49845,N_45566,N_47012);
nand U49846 (N_49846,N_45812,N_45791);
nand U49847 (N_49847,N_45278,N_45629);
xor U49848 (N_49848,N_45556,N_47053);
xor U49849 (N_49849,N_45952,N_47070);
nand U49850 (N_49850,N_45996,N_45601);
nor U49851 (N_49851,N_45472,N_45009);
and U49852 (N_49852,N_46337,N_46281);
nor U49853 (N_49853,N_46523,N_47448);
nand U49854 (N_49854,N_45879,N_47404);
and U49855 (N_49855,N_45421,N_46475);
nor U49856 (N_49856,N_45387,N_46613);
xor U49857 (N_49857,N_45931,N_45519);
nor U49858 (N_49858,N_47214,N_45596);
or U49859 (N_49859,N_46949,N_45955);
and U49860 (N_49860,N_47050,N_46873);
nor U49861 (N_49861,N_46308,N_47419);
or U49862 (N_49862,N_45157,N_46352);
or U49863 (N_49863,N_45115,N_46127);
nand U49864 (N_49864,N_46363,N_46518);
or U49865 (N_49865,N_46601,N_47368);
or U49866 (N_49866,N_46600,N_46062);
and U49867 (N_49867,N_47181,N_45885);
nor U49868 (N_49868,N_45504,N_45851);
nand U49869 (N_49869,N_45351,N_46196);
and U49870 (N_49870,N_45511,N_45034);
or U49871 (N_49871,N_46301,N_47158);
xor U49872 (N_49872,N_46037,N_45760);
nand U49873 (N_49873,N_46421,N_45734);
nand U49874 (N_49874,N_45394,N_45066);
nand U49875 (N_49875,N_45742,N_46185);
and U49876 (N_49876,N_47259,N_46813);
xor U49877 (N_49877,N_47466,N_45977);
nand U49878 (N_49878,N_46484,N_45161);
and U49879 (N_49879,N_46552,N_46434);
nand U49880 (N_49880,N_46614,N_46019);
and U49881 (N_49881,N_46229,N_47488);
nor U49882 (N_49882,N_45644,N_46482);
nor U49883 (N_49883,N_45560,N_46074);
nand U49884 (N_49884,N_45896,N_47076);
and U49885 (N_49885,N_47401,N_45705);
or U49886 (N_49886,N_46985,N_46744);
nand U49887 (N_49887,N_45444,N_47491);
and U49888 (N_49888,N_46543,N_45997);
nor U49889 (N_49889,N_45877,N_47126);
or U49890 (N_49890,N_46645,N_46155);
or U49891 (N_49891,N_46675,N_47393);
xnor U49892 (N_49892,N_46148,N_45250);
and U49893 (N_49893,N_47412,N_45450);
and U49894 (N_49894,N_46740,N_45111);
or U49895 (N_49895,N_45753,N_46019);
nor U49896 (N_49896,N_46314,N_47059);
or U49897 (N_49897,N_46929,N_46017);
and U49898 (N_49898,N_46157,N_46971);
or U49899 (N_49899,N_45095,N_46140);
nor U49900 (N_49900,N_45157,N_46763);
xnor U49901 (N_49901,N_47401,N_47494);
nor U49902 (N_49902,N_46421,N_45815);
and U49903 (N_49903,N_45109,N_45515);
and U49904 (N_49904,N_45527,N_45468);
nor U49905 (N_49905,N_45315,N_46737);
nor U49906 (N_49906,N_46932,N_46777);
nand U49907 (N_49907,N_46254,N_46350);
or U49908 (N_49908,N_46686,N_45736);
nor U49909 (N_49909,N_45265,N_46173);
and U49910 (N_49910,N_45555,N_46186);
nand U49911 (N_49911,N_45368,N_46498);
or U49912 (N_49912,N_46243,N_45513);
nand U49913 (N_49913,N_46585,N_47178);
or U49914 (N_49914,N_47202,N_46807);
and U49915 (N_49915,N_45138,N_46714);
nand U49916 (N_49916,N_47490,N_45553);
nor U49917 (N_49917,N_46954,N_46318);
nand U49918 (N_49918,N_45422,N_47423);
and U49919 (N_49919,N_45939,N_45922);
nor U49920 (N_49920,N_47365,N_47442);
and U49921 (N_49921,N_47125,N_47303);
nand U49922 (N_49922,N_47013,N_46038);
nor U49923 (N_49923,N_45177,N_45159);
and U49924 (N_49924,N_46396,N_46163);
and U49925 (N_49925,N_46293,N_47432);
nor U49926 (N_49926,N_45794,N_46061);
nand U49927 (N_49927,N_45742,N_45637);
nor U49928 (N_49928,N_47346,N_46473);
xnor U49929 (N_49929,N_46173,N_45629);
or U49930 (N_49930,N_46323,N_47040);
or U49931 (N_49931,N_46637,N_45861);
or U49932 (N_49932,N_45421,N_46846);
nand U49933 (N_49933,N_45096,N_47054);
nand U49934 (N_49934,N_47002,N_45442);
nor U49935 (N_49935,N_47125,N_46388);
or U49936 (N_49936,N_45419,N_46557);
nor U49937 (N_49937,N_45744,N_45375);
nor U49938 (N_49938,N_45252,N_47210);
or U49939 (N_49939,N_45083,N_47255);
or U49940 (N_49940,N_46252,N_46056);
nand U49941 (N_49941,N_47274,N_46514);
nor U49942 (N_49942,N_45531,N_47262);
or U49943 (N_49943,N_46674,N_46231);
or U49944 (N_49944,N_45009,N_45334);
xnor U49945 (N_49945,N_45508,N_45829);
xor U49946 (N_49946,N_47423,N_45548);
nand U49947 (N_49947,N_46397,N_46194);
nand U49948 (N_49948,N_45511,N_46744);
nand U49949 (N_49949,N_45482,N_46891);
and U49950 (N_49950,N_46521,N_45115);
nor U49951 (N_49951,N_46926,N_47400);
or U49952 (N_49952,N_46722,N_47330);
or U49953 (N_49953,N_47350,N_45885);
or U49954 (N_49954,N_45705,N_46622);
or U49955 (N_49955,N_45219,N_45538);
or U49956 (N_49956,N_45097,N_45494);
nand U49957 (N_49957,N_46152,N_47059);
nor U49958 (N_49958,N_45661,N_47456);
nand U49959 (N_49959,N_46876,N_46529);
and U49960 (N_49960,N_45526,N_45109);
and U49961 (N_49961,N_45928,N_45187);
nand U49962 (N_49962,N_46562,N_47051);
nor U49963 (N_49963,N_45777,N_45923);
nor U49964 (N_49964,N_45820,N_47188);
or U49965 (N_49965,N_46091,N_46158);
nand U49966 (N_49966,N_46783,N_45351);
and U49967 (N_49967,N_45982,N_47362);
nand U49968 (N_49968,N_47022,N_46876);
or U49969 (N_49969,N_45300,N_46209);
and U49970 (N_49970,N_46784,N_45062);
or U49971 (N_49971,N_46634,N_45699);
nor U49972 (N_49972,N_45132,N_46077);
or U49973 (N_49973,N_45397,N_46509);
or U49974 (N_49974,N_46473,N_45024);
nand U49975 (N_49975,N_45333,N_47383);
and U49976 (N_49976,N_46908,N_46669);
and U49977 (N_49977,N_46056,N_47168);
nand U49978 (N_49978,N_47309,N_46893);
xor U49979 (N_49979,N_47438,N_47174);
and U49980 (N_49980,N_45624,N_45494);
or U49981 (N_49981,N_47186,N_47391);
xor U49982 (N_49982,N_47319,N_47437);
nand U49983 (N_49983,N_47450,N_46377);
nor U49984 (N_49984,N_45058,N_46189);
nor U49985 (N_49985,N_46044,N_46042);
nor U49986 (N_49986,N_45942,N_45768);
and U49987 (N_49987,N_45991,N_45192);
xnor U49988 (N_49988,N_46490,N_45842);
or U49989 (N_49989,N_45013,N_45187);
nor U49990 (N_49990,N_46102,N_45484);
or U49991 (N_49991,N_46389,N_45731);
xor U49992 (N_49992,N_47437,N_46321);
nor U49993 (N_49993,N_47386,N_46055);
nand U49994 (N_49994,N_45151,N_45612);
nor U49995 (N_49995,N_46533,N_46596);
or U49996 (N_49996,N_46391,N_45901);
nand U49997 (N_49997,N_45880,N_45070);
and U49998 (N_49998,N_45860,N_45836);
xor U49999 (N_49999,N_45642,N_46347);
nand UO_0 (O_0,N_48976,N_49038);
nand UO_1 (O_1,N_49680,N_49828);
and UO_2 (O_2,N_47537,N_49530);
nor UO_3 (O_3,N_49989,N_49031);
or UO_4 (O_4,N_48281,N_47611);
nand UO_5 (O_5,N_49830,N_48898);
nand UO_6 (O_6,N_48333,N_49069);
and UO_7 (O_7,N_49938,N_48220);
xnor UO_8 (O_8,N_48454,N_48470);
or UO_9 (O_9,N_47675,N_47962);
and UO_10 (O_10,N_47875,N_49428);
nor UO_11 (O_11,N_49221,N_48244);
nor UO_12 (O_12,N_49350,N_47540);
nor UO_13 (O_13,N_47532,N_48704);
nand UO_14 (O_14,N_49539,N_49956);
nor UO_15 (O_15,N_49771,N_48642);
or UO_16 (O_16,N_48477,N_49160);
nor UO_17 (O_17,N_49168,N_49086);
or UO_18 (O_18,N_48567,N_48628);
nand UO_19 (O_19,N_48964,N_48922);
and UO_20 (O_20,N_49584,N_49367);
nand UO_21 (O_21,N_49731,N_48463);
nand UO_22 (O_22,N_49586,N_48696);
nor UO_23 (O_23,N_47671,N_48757);
nor UO_24 (O_24,N_47708,N_47999);
or UO_25 (O_25,N_47518,N_48969);
or UO_26 (O_26,N_49552,N_48136);
nor UO_27 (O_27,N_47754,N_48232);
nor UO_28 (O_28,N_48049,N_47515);
nor UO_29 (O_29,N_47791,N_49115);
and UO_30 (O_30,N_48042,N_48246);
and UO_31 (O_31,N_48137,N_49833);
or UO_32 (O_32,N_49931,N_49919);
or UO_33 (O_33,N_48574,N_48108);
and UO_34 (O_34,N_47712,N_49492);
and UO_35 (O_35,N_47600,N_47849);
nor UO_36 (O_36,N_48202,N_47822);
and UO_37 (O_37,N_49570,N_48767);
nor UO_38 (O_38,N_48043,N_49531);
and UO_39 (O_39,N_49925,N_48228);
nand UO_40 (O_40,N_49838,N_49276);
and UO_41 (O_41,N_47765,N_49321);
nand UO_42 (O_42,N_49179,N_48818);
nand UO_43 (O_43,N_48159,N_49167);
nand UO_44 (O_44,N_49569,N_47618);
and UO_45 (O_45,N_49389,N_48310);
or UO_46 (O_46,N_47508,N_48441);
or UO_47 (O_47,N_48732,N_48208);
nor UO_48 (O_48,N_49284,N_48100);
and UO_49 (O_49,N_48366,N_48094);
nand UO_50 (O_50,N_48209,N_48096);
or UO_51 (O_51,N_48300,N_49124);
or UO_52 (O_52,N_49161,N_48309);
or UO_53 (O_53,N_49468,N_47858);
nor UO_54 (O_54,N_47805,N_48634);
or UO_55 (O_55,N_48076,N_49968);
or UO_56 (O_56,N_47749,N_48981);
nand UO_57 (O_57,N_49197,N_49722);
and UO_58 (O_58,N_49217,N_47891);
xor UO_59 (O_59,N_48924,N_48806);
xnor UO_60 (O_60,N_48480,N_47677);
and UO_61 (O_61,N_48830,N_48578);
nand UO_62 (O_62,N_48916,N_49690);
or UO_63 (O_63,N_48031,N_49268);
and UO_64 (O_64,N_48793,N_48912);
and UO_65 (O_65,N_47941,N_47715);
and UO_66 (O_66,N_49474,N_48382);
or UO_67 (O_67,N_48637,N_49912);
nand UO_68 (O_68,N_49510,N_47886);
or UO_69 (O_69,N_49053,N_49381);
xnor UO_70 (O_70,N_47978,N_49509);
or UO_71 (O_71,N_48739,N_47757);
nor UO_72 (O_72,N_48845,N_49564);
and UO_73 (O_73,N_49726,N_47780);
or UO_74 (O_74,N_49727,N_49432);
nor UO_75 (O_75,N_48884,N_49274);
nand UO_76 (O_76,N_48283,N_49323);
xor UO_77 (O_77,N_49134,N_49390);
nand UO_78 (O_78,N_47934,N_48458);
or UO_79 (O_79,N_47762,N_48765);
nor UO_80 (O_80,N_48970,N_48685);
and UO_81 (O_81,N_47759,N_49816);
or UO_82 (O_82,N_48059,N_47567);
xor UO_83 (O_83,N_47906,N_49659);
and UO_84 (O_84,N_48038,N_49996);
xnor UO_85 (O_85,N_48760,N_49541);
or UO_86 (O_86,N_49825,N_49252);
or UO_87 (O_87,N_49555,N_47863);
nand UO_88 (O_88,N_49071,N_49653);
nor UO_89 (O_89,N_49739,N_49383);
nand UO_90 (O_90,N_47764,N_49598);
or UO_91 (O_91,N_49412,N_47833);
nand UO_92 (O_92,N_49237,N_48319);
and UO_93 (O_93,N_48506,N_48977);
xor UO_94 (O_94,N_48747,N_49499);
or UO_95 (O_95,N_49190,N_49638);
nand UO_96 (O_96,N_49085,N_48752);
and UO_97 (O_97,N_49880,N_47548);
nor UO_98 (O_98,N_47977,N_48993);
nor UO_99 (O_99,N_48236,N_49758);
xor UO_100 (O_100,N_49741,N_48614);
nor UO_101 (O_101,N_48308,N_49131);
nor UO_102 (O_102,N_48088,N_48329);
nand UO_103 (O_103,N_47761,N_48725);
or UO_104 (O_104,N_49774,N_48180);
and UO_105 (O_105,N_48529,N_49903);
nand UO_106 (O_106,N_47806,N_49534);
or UO_107 (O_107,N_49505,N_47965);
nor UO_108 (O_108,N_49266,N_48770);
or UO_109 (O_109,N_49810,N_48413);
or UO_110 (O_110,N_48412,N_48051);
nand UO_111 (O_111,N_47689,N_49978);
or UO_112 (O_112,N_48996,N_49585);
or UO_113 (O_113,N_48615,N_48937);
or UO_114 (O_114,N_48510,N_49610);
nor UO_115 (O_115,N_48257,N_47866);
nand UO_116 (O_116,N_48841,N_48302);
nand UO_117 (O_117,N_47648,N_48655);
nand UO_118 (O_118,N_47874,N_48758);
xor UO_119 (O_119,N_49821,N_48451);
nor UO_120 (O_120,N_48097,N_48778);
nand UO_121 (O_121,N_48576,N_48691);
nand UO_122 (O_122,N_49720,N_47713);
and UO_123 (O_123,N_49573,N_49634);
nor UO_124 (O_124,N_48876,N_47767);
xnor UO_125 (O_125,N_48086,N_49250);
nor UO_126 (O_126,N_49773,N_49149);
and UO_127 (O_127,N_48870,N_48843);
nand UO_128 (O_128,N_48040,N_48132);
nor UO_129 (O_129,N_47883,N_47629);
and UO_130 (O_130,N_48432,N_47951);
nor UO_131 (O_131,N_47768,N_47572);
nand UO_132 (O_132,N_49713,N_47949);
nor UO_133 (O_133,N_48499,N_48402);
xor UO_134 (O_134,N_48242,N_48552);
nor UO_135 (O_135,N_49769,N_48837);
nor UO_136 (O_136,N_47542,N_48878);
or UO_137 (O_137,N_49300,N_49342);
or UO_138 (O_138,N_47728,N_49138);
or UO_139 (O_139,N_49398,N_48483);
or UO_140 (O_140,N_49861,N_48860);
or UO_141 (O_141,N_48726,N_48507);
or UO_142 (O_142,N_48039,N_48502);
nor UO_143 (O_143,N_48471,N_49910);
nor UO_144 (O_144,N_48145,N_48312);
and UO_145 (O_145,N_49001,N_48724);
xor UO_146 (O_146,N_49642,N_47521);
or UO_147 (O_147,N_49746,N_47651);
nand UO_148 (O_148,N_49316,N_47709);
xor UO_149 (O_149,N_48816,N_48269);
and UO_150 (O_150,N_49035,N_47565);
nand UO_151 (O_151,N_48013,N_48317);
and UO_152 (O_152,N_49278,N_48903);
nand UO_153 (O_153,N_49971,N_49549);
xor UO_154 (O_154,N_47710,N_48178);
nand UO_155 (O_155,N_47993,N_48972);
xnor UO_156 (O_156,N_47606,N_47935);
nand UO_157 (O_157,N_48669,N_48162);
nand UO_158 (O_158,N_49045,N_49074);
or UO_159 (O_159,N_49673,N_48907);
and UO_160 (O_160,N_49106,N_49961);
nor UO_161 (O_161,N_47635,N_49078);
xnor UO_162 (O_162,N_47987,N_48548);
xor UO_163 (O_163,N_47571,N_49789);
and UO_164 (O_164,N_47772,N_47719);
nor UO_165 (O_165,N_48468,N_49360);
or UO_166 (O_166,N_48490,N_49929);
xnor UO_167 (O_167,N_47664,N_48603);
nand UO_168 (O_168,N_48710,N_48360);
nor UO_169 (O_169,N_49027,N_47766);
and UO_170 (O_170,N_47682,N_49139);
nor UO_171 (O_171,N_48868,N_48938);
xnor UO_172 (O_172,N_49671,N_48827);
or UO_173 (O_173,N_47876,N_49437);
or UO_174 (O_174,N_47522,N_47706);
and UO_175 (O_175,N_49332,N_47912);
and UO_176 (O_176,N_49974,N_49211);
nand UO_177 (O_177,N_48847,N_47619);
and UO_178 (O_178,N_48497,N_47793);
and UO_179 (O_179,N_48229,N_48415);
and UO_180 (O_180,N_49275,N_49871);
nor UO_181 (O_181,N_49906,N_49019);
xnor UO_182 (O_182,N_48146,N_49313);
and UO_183 (O_183,N_47528,N_48093);
nand UO_184 (O_184,N_47523,N_47742);
or UO_185 (O_185,N_49459,N_49553);
nand UO_186 (O_186,N_47647,N_48635);
and UO_187 (O_187,N_48619,N_49767);
or UO_188 (O_188,N_48883,N_49756);
or UO_189 (O_189,N_48030,N_48657);
and UO_190 (O_190,N_49312,N_48813);
and UO_191 (O_191,N_49376,N_48745);
xnor UO_192 (O_192,N_47953,N_48945);
or UO_193 (O_193,N_48427,N_48769);
and UO_194 (O_194,N_47847,N_49605);
nand UO_195 (O_195,N_49288,N_47957);
and UO_196 (O_196,N_49839,N_49506);
nand UO_197 (O_197,N_48467,N_49504);
nand UO_198 (O_198,N_48249,N_47992);
nor UO_199 (O_199,N_47788,N_47740);
nand UO_200 (O_200,N_49714,N_47777);
nand UO_201 (O_201,N_48515,N_48825);
nand UO_202 (O_202,N_48905,N_48368);
or UO_203 (O_203,N_48877,N_48929);
or UO_204 (O_204,N_49775,N_49958);
and UO_205 (O_205,N_49556,N_48630);
nor UO_206 (O_206,N_48181,N_47568);
or UO_207 (O_207,N_49467,N_48952);
nor UO_208 (O_208,N_49454,N_47746);
or UO_209 (O_209,N_48150,N_49733);
xnor UO_210 (O_210,N_48340,N_49855);
nand UO_211 (O_211,N_49080,N_47893);
or UO_212 (O_212,N_49719,N_49987);
xor UO_213 (O_213,N_49042,N_48029);
nor UO_214 (O_214,N_49551,N_47990);
nand UO_215 (O_215,N_47673,N_48279);
and UO_216 (O_216,N_47670,N_49725);
nor UO_217 (O_217,N_49473,N_49481);
or UO_218 (O_218,N_48987,N_49574);
nand UO_219 (O_219,N_47760,N_47989);
nor UO_220 (O_220,N_47897,N_49096);
nand UO_221 (O_221,N_47985,N_49755);
nor UO_222 (O_222,N_49753,N_47831);
xor UO_223 (O_223,N_48398,N_48675);
or UO_224 (O_224,N_49923,N_49578);
or UO_225 (O_225,N_49801,N_48528);
nor UO_226 (O_226,N_49147,N_49513);
xor UO_227 (O_227,N_47813,N_48135);
or UO_228 (O_228,N_49976,N_48217);
nor UO_229 (O_229,N_48717,N_49712);
or UO_230 (O_230,N_47937,N_49343);
and UO_231 (O_231,N_49565,N_47633);
nand UO_232 (O_232,N_49143,N_47968);
and UO_233 (O_233,N_49375,N_48580);
nand UO_234 (O_234,N_49365,N_47601);
nor UO_235 (O_235,N_49935,N_48421);
nor UO_236 (O_236,N_49678,N_48826);
and UO_237 (O_237,N_47852,N_48959);
nand UO_238 (O_238,N_48673,N_47845);
and UO_239 (O_239,N_49170,N_49636);
xnor UO_240 (O_240,N_49464,N_47802);
or UO_241 (O_241,N_47610,N_49463);
xor UO_242 (O_242,N_49860,N_47553);
xor UO_243 (O_243,N_48243,N_49227);
nand UO_244 (O_244,N_49180,N_48189);
xor UO_245 (O_245,N_48743,N_48643);
or UO_246 (O_246,N_48064,N_48270);
or UO_247 (O_247,N_47925,N_49255);
xnor UO_248 (O_248,N_49462,N_49583);
nand UO_249 (O_249,N_49141,N_48240);
nand UO_250 (O_250,N_49892,N_48611);
and UO_251 (O_251,N_49701,N_49788);
or UO_252 (O_252,N_47861,N_49595);
or UO_253 (O_253,N_47859,N_49311);
nor UO_254 (O_254,N_49679,N_49715);
xnor UO_255 (O_255,N_49973,N_49178);
and UO_256 (O_256,N_49858,N_48902);
xnor UO_257 (O_257,N_47869,N_48953);
or UO_258 (O_258,N_48605,N_48163);
xnor UO_259 (O_259,N_49740,N_48879);
nand UO_260 (O_260,N_47656,N_48396);
nor UO_261 (O_261,N_49791,N_49814);
or UO_262 (O_262,N_48457,N_48928);
nor UO_263 (O_263,N_47700,N_49859);
and UO_264 (O_264,N_47909,N_48418);
nand UO_265 (O_265,N_48664,N_48335);
nand UO_266 (O_266,N_48728,N_49054);
nor UO_267 (O_267,N_49666,N_47569);
nand UO_268 (O_268,N_49023,N_47860);
xor UO_269 (O_269,N_48046,N_48435);
nor UO_270 (O_270,N_48601,N_49294);
nand UO_271 (O_271,N_48184,N_49682);
xor UO_272 (O_272,N_49614,N_48280);
and UO_273 (O_273,N_49354,N_49808);
or UO_274 (O_274,N_48632,N_49051);
nor UO_275 (O_275,N_47792,N_49851);
nand UO_276 (O_276,N_47870,N_47586);
and UO_277 (O_277,N_47901,N_49724);
and UO_278 (O_278,N_48553,N_48078);
nor UO_279 (O_279,N_48120,N_48535);
nand UO_280 (O_280,N_49271,N_47699);
nor UO_281 (O_281,N_49236,N_48167);
or UO_282 (O_282,N_48289,N_49735);
nor UO_283 (O_283,N_48718,N_49309);
or UO_284 (O_284,N_49108,N_49945);
and UO_285 (O_285,N_48160,N_49022);
nand UO_286 (O_286,N_48836,N_49408);
and UO_287 (O_287,N_49223,N_48484);
nor UO_288 (O_288,N_49994,N_49813);
nor UO_289 (O_289,N_48624,N_48617);
nand UO_290 (O_290,N_49397,N_49544);
and UO_291 (O_291,N_47955,N_47836);
nor UO_292 (O_292,N_48284,N_49199);
nand UO_293 (O_293,N_48800,N_48749);
or UO_294 (O_294,N_49451,N_49920);
nor UO_295 (O_295,N_49647,N_49244);
and UO_296 (O_296,N_48737,N_48720);
xor UO_297 (O_297,N_48833,N_49837);
or UO_298 (O_298,N_49981,N_48095);
nand UO_299 (O_299,N_47686,N_49201);
or UO_300 (O_300,N_48602,N_49441);
nand UO_301 (O_301,N_49356,N_49811);
nor UO_302 (O_302,N_49439,N_48200);
or UO_303 (O_303,N_49848,N_48142);
xnor UO_304 (O_304,N_48393,N_48139);
nand UO_305 (O_305,N_49104,N_49621);
nand UO_306 (O_306,N_48128,N_49533);
and UO_307 (O_307,N_48156,N_48130);
nand UO_308 (O_308,N_47576,N_48526);
or UO_309 (O_309,N_47817,N_48581);
or UO_310 (O_310,N_48835,N_48730);
nand UO_311 (O_311,N_48109,N_47818);
and UO_312 (O_312,N_48362,N_49183);
nand UO_313 (O_313,N_49254,N_49305);
or UO_314 (O_314,N_49664,N_49282);
or UO_315 (O_315,N_48449,N_49650);
nand UO_316 (O_316,N_49964,N_48307);
and UO_317 (O_317,N_49159,N_48384);
or UO_318 (O_318,N_47646,N_47581);
nor UO_319 (O_319,N_49171,N_49602);
and UO_320 (O_320,N_48839,N_49628);
and UO_321 (O_321,N_49029,N_48052);
nor UO_322 (O_322,N_49456,N_48462);
and UO_323 (O_323,N_48460,N_49932);
nand UO_324 (O_324,N_48958,N_49844);
nor UO_325 (O_325,N_48324,N_49803);
nor UO_326 (O_326,N_48067,N_49946);
and UO_327 (O_327,N_48620,N_48895);
xor UO_328 (O_328,N_48684,N_49101);
and UO_329 (O_329,N_48357,N_47920);
and UO_330 (O_330,N_48225,N_47758);
or UO_331 (O_331,N_49818,N_49154);
or UO_332 (O_332,N_49662,N_48399);
or UO_333 (O_333,N_48007,N_48971);
nor UO_334 (O_334,N_48316,N_47520);
nand UO_335 (O_335,N_47782,N_49667);
or UO_336 (O_336,N_49024,N_48985);
or UO_337 (O_337,N_48173,N_48613);
xnor UO_338 (O_338,N_49340,N_49969);
or UO_339 (O_339,N_48320,N_47641);
and UO_340 (O_340,N_48572,N_49301);
and UO_341 (O_341,N_49111,N_48736);
nand UO_342 (O_342,N_48211,N_49654);
nand UO_343 (O_343,N_48414,N_47650);
or UO_344 (O_344,N_49487,N_48161);
nor UO_345 (O_345,N_48858,N_48295);
nor UO_346 (O_346,N_48659,N_49299);
nand UO_347 (O_347,N_47573,N_48573);
xnor UO_348 (O_348,N_47888,N_49500);
or UO_349 (O_349,N_48285,N_47654);
or UO_350 (O_350,N_48666,N_49882);
xor UO_351 (O_351,N_47970,N_49256);
or UO_352 (O_352,N_47778,N_49913);
nor UO_353 (O_353,N_48188,N_49153);
or UO_354 (O_354,N_47819,N_49004);
nand UO_355 (O_355,N_49327,N_48395);
or UO_356 (O_356,N_49224,N_48616);
and UO_357 (O_357,N_47880,N_49387);
and UO_358 (O_358,N_47557,N_48799);
nor UO_359 (O_359,N_49461,N_48492);
nand UO_360 (O_360,N_49623,N_48445);
nor UO_361 (O_361,N_49315,N_49380);
and UO_362 (O_362,N_49422,N_48668);
xor UO_363 (O_363,N_48152,N_49493);
nor UO_364 (O_364,N_48590,N_48822);
nand UO_365 (O_365,N_49264,N_49145);
nand UO_366 (O_366,N_49545,N_48266);
and UO_367 (O_367,N_49942,N_48890);
and UO_368 (O_368,N_48595,N_49070);
and UO_369 (O_369,N_49207,N_49466);
nand UO_370 (O_370,N_48585,N_49607);
nor UO_371 (O_371,N_49182,N_47775);
and UO_372 (O_372,N_48589,N_49377);
nand UO_373 (O_373,N_49874,N_49425);
or UO_374 (O_374,N_48423,N_47716);
nand UO_375 (O_375,N_47517,N_47735);
nand UO_376 (O_376,N_49174,N_48017);
xor UO_377 (O_377,N_48509,N_49943);
nor UO_378 (O_378,N_49802,N_48777);
nand UO_379 (O_379,N_47631,N_49633);
nand UO_380 (O_380,N_48962,N_49897);
or UO_381 (O_381,N_49480,N_49100);
nor UO_382 (O_382,N_48683,N_47628);
nor UO_383 (O_383,N_49829,N_48983);
or UO_384 (O_384,N_49242,N_48562);
nand UO_385 (O_385,N_49547,N_48247);
nand UO_386 (O_386,N_48811,N_49896);
nand UO_387 (O_387,N_49516,N_48627);
nand UO_388 (O_388,N_48230,N_48448);
nor UO_389 (O_389,N_48033,N_48798);
nor UO_390 (O_390,N_48301,N_47695);
nor UO_391 (O_391,N_48450,N_49842);
nor UO_392 (O_392,N_48559,N_47915);
nand UO_393 (O_393,N_49353,N_49857);
nand UO_394 (O_394,N_48154,N_48123);
nor UO_395 (O_395,N_47867,N_47602);
nand UO_396 (O_396,N_49279,N_47707);
nor UO_397 (O_397,N_49296,N_49542);
or UO_398 (O_398,N_47666,N_48795);
or UO_399 (O_399,N_49675,N_48222);
and UO_400 (O_400,N_49947,N_48936);
and UO_401 (O_401,N_49674,N_47913);
nand UO_402 (O_402,N_48420,N_47721);
nand UO_403 (O_403,N_49772,N_49890);
nand UO_404 (O_404,N_47748,N_47835);
or UO_405 (O_405,N_49949,N_48764);
or UO_406 (O_406,N_48610,N_47679);
and UO_407 (O_407,N_49705,N_49091);
nor UO_408 (O_408,N_47687,N_48408);
nand UO_409 (O_409,N_49329,N_47984);
or UO_410 (O_410,N_49099,N_48278);
nand UO_411 (O_411,N_47804,N_48846);
and UO_412 (O_412,N_49637,N_48943);
nand UO_413 (O_413,N_47649,N_49465);
nor UO_414 (O_414,N_48797,N_47585);
nor UO_415 (O_415,N_47637,N_48168);
xnor UO_416 (O_416,N_49780,N_47607);
and UO_417 (O_417,N_49409,N_49962);
xor UO_418 (O_418,N_47956,N_49303);
nor UO_419 (O_419,N_49672,N_49410);
nor UO_420 (O_420,N_47588,N_49436);
nand UO_421 (O_421,N_48688,N_48311);
or UO_422 (O_422,N_47931,N_47959);
and UO_423 (O_423,N_49702,N_48028);
nor UO_424 (O_424,N_49317,N_48264);
nand UO_425 (O_425,N_48794,N_47816);
or UO_426 (O_426,N_48000,N_49326);
nand UO_427 (O_427,N_47640,N_47663);
and UO_428 (O_428,N_48607,N_49611);
nand UO_429 (O_429,N_48920,N_48489);
or UO_430 (O_430,N_49742,N_49140);
nor UO_431 (O_431,N_49191,N_48126);
nor UO_432 (O_432,N_47599,N_49694);
and UO_433 (O_433,N_49215,N_47530);
nand UO_434 (O_434,N_48864,N_49314);
or UO_435 (O_435,N_48367,N_48998);
or UO_436 (O_436,N_48113,N_48862);
xnor UO_437 (O_437,N_49561,N_48260);
or UO_438 (O_438,N_47662,N_48982);
xnor UO_439 (O_439,N_48237,N_48500);
and UO_440 (O_440,N_49229,N_49277);
nand UO_441 (O_441,N_49357,N_47616);
nor UO_442 (O_442,N_49696,N_49900);
and UO_443 (O_443,N_49014,N_48401);
nand UO_444 (O_444,N_47730,N_48694);
xnor UO_445 (O_445,N_48695,N_48119);
and UO_446 (O_446,N_49012,N_47997);
or UO_447 (O_447,N_49990,N_48537);
or UO_448 (O_448,N_49937,N_47979);
xnor UO_449 (O_449,N_47625,N_47604);
or UO_450 (O_450,N_49306,N_48524);
xor UO_451 (O_451,N_48430,N_49185);
nand UO_452 (O_452,N_49895,N_47524);
nor UO_453 (O_453,N_49372,N_47621);
or UO_454 (O_454,N_47502,N_48359);
nand UO_455 (O_455,N_48991,N_48009);
nand UO_456 (O_456,N_48772,N_47794);
nor UO_457 (O_457,N_49033,N_48345);
or UO_458 (O_458,N_49226,N_49563);
nor UO_459 (O_459,N_49495,N_48919);
or UO_460 (O_460,N_48966,N_48873);
nor UO_461 (O_461,N_47595,N_49497);
and UO_462 (O_462,N_49449,N_49339);
nand UO_463 (O_463,N_49512,N_48824);
nor UO_464 (O_464,N_48003,N_47674);
nand UO_465 (O_465,N_49856,N_47832);
nor UO_466 (O_466,N_48901,N_49879);
and UO_467 (O_467,N_48508,N_49386);
or UO_468 (O_468,N_47516,N_49063);
nor UO_469 (O_469,N_49960,N_48298);
and UO_470 (O_470,N_48944,N_48452);
and UO_471 (O_471,N_48440,N_49886);
xor UO_472 (O_472,N_47864,N_48106);
and UO_473 (O_473,N_49572,N_48660);
or UO_474 (O_474,N_49346,N_48804);
nand UO_475 (O_475,N_47653,N_48692);
nor UO_476 (O_476,N_49554,N_49730);
or UO_477 (O_477,N_49006,N_47737);
and UO_478 (O_478,N_47884,N_49194);
or UO_479 (O_479,N_48461,N_49950);
nand UO_480 (O_480,N_47773,N_49576);
nor UO_481 (O_481,N_47552,N_49955);
nor UO_482 (O_482,N_47825,N_48677);
nor UO_483 (O_483,N_49128,N_48556);
nand UO_484 (O_484,N_48428,N_48253);
xor UO_485 (O_485,N_48703,N_48261);
nand UO_486 (O_486,N_48272,N_48582);
or UO_487 (O_487,N_49088,N_48277);
and UO_488 (O_488,N_48874,N_49076);
or UO_489 (O_489,N_49641,N_48789);
xor UO_490 (O_490,N_49447,N_49876);
nor UO_491 (O_491,N_48105,N_49285);
nand UO_492 (O_492,N_49988,N_48872);
or UO_493 (O_493,N_49588,N_48223);
or UO_494 (O_494,N_49807,N_49281);
and UO_495 (O_495,N_48252,N_47842);
and UO_496 (O_496,N_49656,N_48570);
or UO_497 (O_497,N_48075,N_48734);
nor UO_498 (O_498,N_49518,N_49055);
xor UO_499 (O_499,N_49697,N_49385);
or UO_500 (O_500,N_49934,N_49322);
xnor UO_501 (O_501,N_49247,N_48185);
xor UO_502 (O_502,N_49526,N_48338);
and UO_503 (O_503,N_48834,N_49652);
xor UO_504 (O_504,N_48933,N_47535);
nor UO_505 (O_505,N_49157,N_48482);
nor UO_506 (O_506,N_47669,N_48478);
nor UO_507 (O_507,N_49590,N_47905);
and UO_508 (O_508,N_49165,N_48917);
or UO_509 (O_509,N_48554,N_48676);
nand UO_510 (O_510,N_48256,N_49040);
nand UO_511 (O_511,N_49749,N_48424);
nor UO_512 (O_512,N_48687,N_49535);
or UO_513 (O_513,N_48383,N_47509);
nor UO_514 (O_514,N_48783,N_48034);
and UO_515 (O_515,N_48594,N_47902);
nand UO_516 (O_516,N_48848,N_49898);
xnor UO_517 (O_517,N_48274,N_48201);
and UO_518 (O_518,N_49782,N_48979);
nand UO_519 (O_519,N_48176,N_47904);
nand UO_520 (O_520,N_48348,N_48287);
nand UO_521 (O_521,N_49850,N_47636);
nor UO_522 (O_522,N_48918,N_48140);
nor UO_523 (O_523,N_49668,N_47536);
nor UO_524 (O_524,N_47967,N_49348);
nor UO_525 (O_525,N_49328,N_49458);
or UO_526 (O_526,N_49445,N_48784);
nand UO_527 (O_527,N_48775,N_48066);
nand UO_528 (O_528,N_49137,N_49831);
or UO_529 (O_529,N_49234,N_48290);
and UO_530 (O_530,N_49186,N_48378);
nand UO_531 (O_531,N_49995,N_49181);
xnor UO_532 (O_532,N_49762,N_49257);
and UO_533 (O_533,N_49620,N_48861);
or UO_534 (O_534,N_48268,N_48438);
xor UO_535 (O_535,N_47809,N_47879);
nor UO_536 (O_536,N_48195,N_47570);
xnor UO_537 (O_537,N_47652,N_48262);
nor UO_538 (O_538,N_48134,N_49706);
and UO_539 (O_539,N_49496,N_47608);
nor UO_540 (O_540,N_47612,N_47873);
or UO_541 (O_541,N_48851,N_48899);
nand UO_542 (O_542,N_48505,N_49627);
or UO_543 (O_543,N_48215,N_47555);
or UO_544 (O_544,N_48925,N_49424);
nand UO_545 (O_545,N_49954,N_49187);
or UO_546 (O_546,N_47738,N_48361);
nor UO_547 (O_547,N_48942,N_48035);
or UO_548 (O_548,N_48487,N_49832);
and UO_549 (O_549,N_48347,N_48431);
and UO_550 (O_550,N_47890,N_49399);
xor UO_551 (O_551,N_48355,N_49384);
and UO_552 (O_552,N_47741,N_48443);
or UO_553 (O_553,N_47733,N_48464);
or UO_554 (O_554,N_48842,N_48880);
nor UO_555 (O_555,N_48565,N_47854);
or UO_556 (O_556,N_48644,N_48214);
or UO_557 (O_557,N_48372,N_48521);
nor UO_558 (O_558,N_49112,N_49098);
nor UO_559 (O_559,N_48417,N_48349);
nor UO_560 (O_560,N_48711,N_48194);
and UO_561 (O_561,N_47562,N_49822);
and UO_562 (O_562,N_49596,N_49589);
and UO_563 (O_563,N_49097,N_48297);
and UO_564 (O_564,N_49433,N_48885);
or UO_565 (O_565,N_47995,N_48481);
and UO_566 (O_566,N_48085,N_49475);
nand UO_567 (O_567,N_49352,N_48947);
nor UO_568 (O_568,N_48197,N_48315);
nand UO_569 (O_569,N_48286,N_48425);
xnor UO_570 (O_570,N_47892,N_49557);
and UO_571 (O_571,N_49538,N_47948);
and UO_572 (O_572,N_48699,N_47539);
xor UO_573 (O_573,N_48336,N_47501);
nor UO_574 (O_574,N_48473,N_47903);
nand UO_575 (O_575,N_48586,N_48678);
nor UO_576 (O_576,N_49907,N_49738);
and UO_577 (O_577,N_49784,N_49017);
and UO_578 (O_578,N_48271,N_47667);
or UO_579 (O_579,N_47546,N_49093);
nor UO_580 (O_580,N_49366,N_49318);
and UO_581 (O_581,N_47691,N_48318);
nand UO_582 (O_582,N_49765,N_47750);
or UO_583 (O_583,N_49927,N_47739);
nor UO_584 (O_584,N_48558,N_48020);
nand UO_585 (O_585,N_47837,N_48639);
nor UO_586 (O_586,N_47856,N_48817);
xor UO_587 (O_587,N_49616,N_49663);
nor UO_588 (O_588,N_48346,N_48493);
xor UO_589 (O_589,N_49710,N_49952);
nor UO_590 (O_590,N_48263,N_49253);
or UO_591 (O_591,N_49893,N_48867);
nor UO_592 (O_592,N_48205,N_48045);
nor UO_593 (O_593,N_49619,N_48997);
and UO_594 (O_594,N_49241,N_48213);
and UO_595 (O_595,N_48853,N_48314);
nor UO_596 (O_596,N_49026,N_48571);
or UO_597 (O_597,N_47911,N_48053);
nor UO_598 (O_598,N_48875,N_47752);
nand UO_599 (O_599,N_48062,N_48110);
xnor UO_600 (O_600,N_49166,N_48805);
and UO_601 (O_601,N_49273,N_48186);
and UO_602 (O_602,N_49681,N_49047);
nor UO_603 (O_603,N_47507,N_49214);
nand UO_604 (O_604,N_49095,N_48709);
nand UO_605 (O_605,N_49411,N_49013);
or UO_606 (O_606,N_47930,N_47812);
or UO_607 (O_607,N_49151,N_48706);
nand UO_608 (O_608,N_48609,N_49135);
xnor UO_609 (O_609,N_49109,N_48406);
nand UO_610 (O_610,N_48815,N_49362);
nand UO_611 (O_611,N_48474,N_49144);
and UO_612 (O_612,N_49936,N_49593);
nor UO_613 (O_613,N_49905,N_49232);
xnor UO_614 (O_614,N_48596,N_48954);
nand UO_615 (O_615,N_47543,N_49081);
or UO_616 (O_616,N_47789,N_48512);
or UO_617 (O_617,N_48179,N_49037);
or UO_618 (O_618,N_48199,N_49193);
nor UO_619 (O_619,N_48183,N_48658);
or UO_620 (O_620,N_48857,N_48715);
nand UO_621 (O_621,N_48762,N_47729);
nand UO_622 (O_622,N_48077,N_49597);
or UO_623 (O_623,N_49421,N_48363);
xnor UO_624 (O_624,N_48442,N_47587);
xor UO_625 (O_625,N_47942,N_48560);
nand UO_626 (O_626,N_48557,N_49670);
nor UO_627 (O_627,N_48018,N_48790);
and UO_628 (O_628,N_49520,N_47630);
and UO_629 (O_629,N_49817,N_48501);
and UO_630 (O_630,N_47626,N_48723);
nand UO_631 (O_631,N_49122,N_49400);
and UO_632 (O_632,N_49297,N_49172);
and UO_633 (O_633,N_47853,N_47800);
or UO_634 (O_634,N_48436,N_49852);
or UO_635 (O_635,N_48071,N_49687);
xor UO_636 (O_636,N_47960,N_49718);
nor UO_637 (O_637,N_47798,N_48091);
nor UO_638 (O_638,N_47918,N_48713);
or UO_639 (O_639,N_48555,N_48294);
and UO_640 (O_640,N_48148,N_49058);
nor UO_641 (O_641,N_47582,N_48940);
or UO_642 (O_642,N_49537,N_47991);
nand UO_643 (O_643,N_49894,N_49416);
nand UO_644 (O_644,N_47824,N_49501);
and UO_645 (O_645,N_47969,N_49118);
nor UO_646 (O_646,N_47574,N_49862);
nand UO_647 (O_647,N_48542,N_47580);
and UO_648 (O_648,N_48763,N_49543);
xor UO_649 (O_649,N_47963,N_48422);
or UO_650 (O_650,N_48672,N_49635);
and UO_651 (O_651,N_49930,N_48771);
nand UO_652 (O_652,N_47770,N_47694);
or UO_653 (O_653,N_48129,N_48612);
nand UO_654 (O_654,N_48002,N_47790);
nor UO_655 (O_655,N_49815,N_48328);
or UO_656 (O_656,N_49591,N_48303);
or UO_657 (O_657,N_48456,N_48404);
nand UO_658 (O_658,N_49889,N_47623);
nor UO_659 (O_659,N_48494,N_48948);
or UO_660 (O_660,N_47828,N_49373);
nor UO_661 (O_661,N_48177,N_48988);
nor UO_662 (O_662,N_49388,N_49125);
nand UO_663 (O_663,N_49401,N_49524);
or UO_664 (O_664,N_49625,N_48690);
and UO_665 (O_665,N_49016,N_49032);
nor UO_666 (O_666,N_48829,N_49442);
nand UO_667 (O_667,N_48025,N_49594);
nor UO_668 (O_668,N_49034,N_48255);
nor UO_669 (O_669,N_49717,N_48667);
nand UO_670 (O_670,N_49025,N_47510);
and UO_671 (O_671,N_49902,N_48955);
nand UO_672 (O_672,N_47988,N_47921);
xor UO_673 (O_673,N_48759,N_48305);
nand UO_674 (O_674,N_49571,N_48164);
or UO_675 (O_675,N_49909,N_48169);
nand UO_676 (O_676,N_49918,N_47933);
xor UO_677 (O_677,N_48275,N_48840);
nor UO_678 (O_678,N_49688,N_48886);
nand UO_679 (O_679,N_47826,N_47538);
and UO_680 (O_680,N_49310,N_48224);
or UO_681 (O_681,N_48485,N_49146);
nor UO_682 (O_682,N_48859,N_49062);
nor UO_683 (O_683,N_49057,N_49599);
and UO_684 (O_684,N_48522,N_49324);
nor UO_685 (O_685,N_49263,N_47795);
and UO_686 (O_686,N_48549,N_48999);
or UO_687 (O_687,N_49863,N_49854);
or UO_688 (O_688,N_48652,N_49752);
or UO_689 (O_689,N_48079,N_48939);
nor UO_690 (O_690,N_47917,N_48486);
nor UO_691 (O_691,N_48231,N_48661);
and UO_692 (O_692,N_48980,N_47525);
and UO_693 (O_693,N_47658,N_49129);
nand UO_694 (O_694,N_48466,N_48187);
or UO_695 (O_695,N_47895,N_49689);
xnor UO_696 (O_696,N_49626,N_48015);
and UO_697 (O_697,N_47644,N_48496);
and UO_698 (O_698,N_48153,N_47871);
or UO_699 (O_699,N_49676,N_47566);
nand UO_700 (O_700,N_48171,N_49345);
nor UO_701 (O_701,N_48226,N_48103);
nand UO_702 (O_702,N_49846,N_48904);
or UO_703 (O_703,N_49723,N_47850);
nor UO_704 (O_704,N_47797,N_48796);
xor UO_705 (O_705,N_49612,N_49130);
nand UO_706 (O_706,N_49745,N_48591);
or UO_707 (O_707,N_48742,N_49440);
and UO_708 (O_708,N_47513,N_48712);
xor UO_709 (O_709,N_48063,N_49184);
or UO_710 (O_710,N_49420,N_49392);
and UO_711 (O_711,N_49778,N_48563);
and UO_712 (O_712,N_48671,N_47592);
nor UO_713 (O_713,N_47996,N_47511);
and UO_714 (O_714,N_48023,N_48597);
nor UO_715 (O_715,N_47928,N_47534);
or UO_716 (O_716,N_48446,N_49028);
nand UO_717 (O_717,N_48056,N_47878);
nand UO_718 (O_718,N_47862,N_49643);
and UO_719 (O_719,N_47551,N_47556);
nand UO_720 (O_720,N_49716,N_49333);
or UO_721 (O_721,N_47827,N_48910);
nor UO_722 (O_722,N_48083,N_48514);
nand UO_723 (O_723,N_48932,N_48766);
nand UO_724 (O_724,N_48248,N_48994);
or UO_725 (O_725,N_48327,N_47541);
nor UO_726 (O_726,N_49448,N_48854);
nand UO_727 (O_727,N_49246,N_47727);
nor UO_728 (O_728,N_49624,N_48381);
and UO_729 (O_729,N_48894,N_48326);
nor UO_730 (O_730,N_48923,N_49613);
nor UO_731 (O_731,N_49985,N_47946);
nor UO_732 (O_732,N_47983,N_48748);
nand UO_733 (O_733,N_47763,N_49581);
nor UO_734 (O_734,N_49630,N_47944);
xnor UO_735 (O_735,N_48170,N_48869);
or UO_736 (O_736,N_49225,N_49213);
nand UO_737 (O_737,N_47561,N_48437);
nand UO_738 (O_738,N_48014,N_48989);
nand UO_739 (O_739,N_48115,N_49202);
nor UO_740 (O_740,N_48060,N_48935);
xnor UO_741 (O_741,N_49692,N_48027);
or UO_742 (O_742,N_48476,N_49548);
nand UO_743 (O_743,N_49370,N_48058);
and UO_744 (O_744,N_48592,N_47605);
or UO_745 (O_745,N_49188,N_47591);
nor UO_746 (O_746,N_49587,N_49162);
and UO_747 (O_747,N_49498,N_48569);
nor UO_748 (O_748,N_48504,N_49116);
nand UO_749 (O_749,N_49704,N_47681);
nor UO_750 (O_750,N_49517,N_49087);
and UO_751 (O_751,N_48344,N_48037);
or UO_752 (O_752,N_49550,N_48011);
nand UO_753 (O_753,N_48593,N_49864);
or UO_754 (O_754,N_48488,N_49748);
or UO_755 (O_755,N_49640,N_47964);
nor UO_756 (O_756,N_48698,N_49163);
or UO_757 (O_757,N_47945,N_48754);
and UO_758 (O_758,N_49575,N_48267);
nor UO_759 (O_759,N_47657,N_47554);
or UO_760 (O_760,N_48995,N_48965);
nor UO_761 (O_761,N_48331,N_47678);
nand UO_762 (O_762,N_49011,N_47620);
nor UO_763 (O_763,N_48111,N_48598);
and UO_764 (O_764,N_49210,N_49568);
nor UO_765 (O_765,N_49396,N_49413);
and UO_766 (O_766,N_47784,N_48379);
or UO_767 (O_767,N_47560,N_49484);
or UO_768 (O_768,N_47659,N_48479);
nor UO_769 (O_769,N_49812,N_47787);
nor UO_770 (O_770,N_48218,N_49113);
xnor UO_771 (O_771,N_47971,N_48124);
nor UO_772 (O_772,N_48407,N_47590);
or UO_773 (O_773,N_47974,N_49457);
and UO_774 (O_774,N_49683,N_48375);
nand UO_775 (O_775,N_49514,N_48026);
and UO_776 (O_776,N_49827,N_47527);
or UO_777 (O_777,N_49218,N_49270);
and UO_778 (O_778,N_47642,N_47705);
and UO_779 (O_779,N_47688,N_49272);
nor UO_780 (O_780,N_49728,N_49984);
nor UO_781 (O_781,N_48405,N_47952);
nor UO_782 (O_782,N_49494,N_49208);
or UO_783 (O_783,N_49991,N_49754);
or UO_784 (O_784,N_49522,N_48889);
and UO_785 (O_785,N_47732,N_47627);
nor UO_786 (O_786,N_49430,N_49983);
xnor UO_787 (O_787,N_49823,N_47575);
and UO_788 (O_788,N_48656,N_49094);
nor UO_789 (O_789,N_49997,N_49283);
nand UO_790 (O_790,N_49979,N_47731);
nor UO_791 (O_791,N_48566,N_49786);
or UO_792 (O_792,N_49361,N_48741);
nand UO_793 (O_793,N_49404,N_47550);
and UO_794 (O_794,N_49133,N_47982);
nand UO_795 (O_795,N_49750,N_49114);
xnor UO_796 (O_796,N_49503,N_49797);
and UO_797 (O_797,N_49355,N_47865);
or UO_798 (O_798,N_48306,N_49020);
and UO_799 (O_799,N_49941,N_48753);
and UO_800 (O_800,N_48158,N_48016);
nor UO_801 (O_801,N_48400,N_49150);
nand UO_802 (O_802,N_48755,N_47839);
nand UO_803 (O_803,N_48299,N_48934);
xnor UO_804 (O_804,N_49615,N_49426);
or UO_805 (O_805,N_49866,N_48004);
nand UO_806 (O_806,N_48746,N_49721);
nand UO_807 (O_807,N_48721,N_48191);
or UO_808 (O_808,N_49700,N_47981);
or UO_809 (O_809,N_48831,N_48057);
or UO_810 (O_810,N_47718,N_48662);
nor UO_811 (O_811,N_47980,N_49009);
and UO_812 (O_812,N_49155,N_47769);
or UO_813 (O_813,N_49407,N_49922);
nor UO_814 (O_814,N_49546,N_48074);
and UO_815 (O_815,N_48540,N_49779);
nor UO_816 (O_816,N_48047,N_49258);
nor UO_817 (O_817,N_49577,N_48674);
nand UO_818 (O_818,N_48536,N_48444);
and UO_819 (O_819,N_49770,N_49349);
nor UO_820 (O_820,N_49233,N_48838);
or UO_821 (O_821,N_49438,N_49686);
nand UO_822 (O_822,N_49603,N_48370);
nor UO_823 (O_823,N_49230,N_48021);
and UO_824 (O_824,N_48951,N_49911);
or UO_825 (O_825,N_49794,N_47672);
and UO_826 (O_826,N_49540,N_47598);
nand UO_827 (O_827,N_49402,N_49759);
and UO_828 (O_828,N_49986,N_49567);
nand UO_829 (O_829,N_47885,N_49238);
xnor UO_830 (O_830,N_48541,N_47725);
nor UO_831 (O_831,N_49691,N_49368);
xnor UO_832 (O_832,N_48961,N_48700);
nand UO_833 (O_833,N_49793,N_48102);
xor UO_834 (O_834,N_48546,N_48006);
nand UO_835 (O_835,N_47896,N_48744);
nand UO_836 (O_836,N_47848,N_47697);
and UO_837 (O_837,N_49002,N_49046);
and UO_838 (O_838,N_48121,N_49077);
and UO_839 (O_839,N_48334,N_48530);
nand UO_840 (O_840,N_49959,N_48654);
nand UO_841 (O_841,N_49245,N_47645);
nand UO_842 (O_842,N_48012,N_47929);
and UO_843 (O_843,N_49562,N_48358);
and UO_844 (O_844,N_49414,N_48852);
and UO_845 (O_845,N_47665,N_49849);
and UO_846 (O_846,N_48210,N_49039);
or UO_847 (O_847,N_48190,N_49431);
xnor UO_848 (O_848,N_47872,N_47814);
nand UO_849 (O_849,N_48781,N_49049);
and UO_850 (O_850,N_47711,N_49156);
nor UO_851 (O_851,N_48638,N_47834);
nor UO_852 (O_852,N_48321,N_48665);
and UO_853 (O_853,N_49592,N_47734);
and UO_854 (O_854,N_49320,N_49090);
and UO_855 (O_855,N_48527,N_47771);
or UO_856 (O_856,N_48727,N_49734);
or UO_857 (O_857,N_48697,N_49695);
and UO_858 (O_858,N_49806,N_47744);
xor UO_859 (O_859,N_49999,N_47545);
nand UO_860 (O_860,N_47726,N_48192);
or UO_861 (O_861,N_48705,N_48251);
nand UO_862 (O_862,N_49423,N_48495);
and UO_863 (O_863,N_49489,N_49883);
and UO_864 (O_864,N_49371,N_47803);
or UO_865 (O_865,N_47954,N_47811);
nand UO_866 (O_866,N_47881,N_48207);
and UO_867 (O_867,N_49452,N_48821);
nand UO_868 (O_868,N_49865,N_49804);
and UO_869 (O_869,N_47910,N_48882);
nor UO_870 (O_870,N_48551,N_49609);
nand UO_871 (O_871,N_47702,N_48065);
nor UO_872 (O_872,N_48353,N_49977);
nand UO_873 (O_873,N_49403,N_49776);
or UO_874 (O_874,N_49853,N_49527);
or UO_875 (O_875,N_48900,N_48645);
or UO_876 (O_876,N_48072,N_49064);
nor UO_877 (O_877,N_47504,N_48801);
or UO_878 (O_878,N_48282,N_49608);
xor UO_879 (O_879,N_49736,N_47786);
or UO_880 (O_880,N_49631,N_48735);
xnor UO_881 (O_881,N_48089,N_49291);
nor UO_882 (O_882,N_49887,N_48926);
nand UO_883 (O_883,N_49760,N_48702);
and UO_884 (O_884,N_48503,N_48722);
xor UO_885 (O_885,N_48385,N_48024);
nor UO_886 (O_886,N_48532,N_49030);
and UO_887 (O_887,N_48809,N_49737);
nor UO_888 (O_888,N_48693,N_48866);
or UO_889 (O_889,N_47900,N_48157);
nor UO_890 (O_890,N_47855,N_49699);
and UO_891 (O_891,N_48787,N_48606);
xnor UO_892 (O_892,N_49703,N_48774);
or UO_893 (O_893,N_49841,N_48844);
nor UO_894 (O_894,N_49044,N_47584);
or UO_895 (O_895,N_48544,N_48386);
and UO_896 (O_896,N_48101,N_49658);
nor UO_897 (O_897,N_49928,N_48534);
nand UO_898 (O_898,N_49358,N_47751);
or UO_899 (O_899,N_47634,N_49259);
and UO_900 (O_900,N_48127,N_48782);
xor UO_901 (O_901,N_48429,N_49079);
nand UO_902 (O_902,N_48409,N_48410);
and UO_903 (O_903,N_48984,N_49363);
and UO_904 (O_904,N_49405,N_49041);
and UO_905 (O_905,N_48296,N_47851);
nor UO_906 (O_906,N_47958,N_48332);
and UO_907 (O_907,N_47877,N_48908);
nor UO_908 (O_908,N_49127,N_48098);
and UO_909 (O_909,N_48788,N_49970);
nand UO_910 (O_910,N_49507,N_49685);
nand UO_911 (O_911,N_48750,N_49629);
or UO_912 (O_912,N_49231,N_47829);
nor UO_913 (O_913,N_48233,N_48896);
nor UO_914 (O_914,N_47843,N_49820);
and UO_915 (O_915,N_49021,N_49901);
nor UO_916 (O_916,N_49083,N_49477);
or UO_917 (O_917,N_49287,N_49915);
nand UO_918 (O_918,N_47916,N_48863);
nand UO_919 (O_919,N_47815,N_48325);
nand UO_920 (O_920,N_49307,N_48651);
and UO_921 (O_921,N_49528,N_48212);
nor UO_922 (O_922,N_48738,N_49007);
nand UO_923 (O_923,N_48960,N_48193);
nand UO_924 (O_924,N_47519,N_47594);
nand UO_925 (O_925,N_49117,N_49335);
and UO_926 (O_926,N_48791,N_48323);
nand UO_927 (O_927,N_47698,N_48350);
nor UO_928 (O_928,N_48974,N_47638);
or UO_929 (O_929,N_47639,N_48689);
nand UO_930 (O_930,N_48114,N_48629);
and UO_931 (O_931,N_48491,N_47701);
nor UO_932 (O_932,N_49478,N_47807);
xnor UO_933 (O_933,N_48931,N_49073);
nor UO_934 (O_934,N_49617,N_49566);
nor UO_935 (O_935,N_47547,N_49677);
xnor UO_936 (O_936,N_49834,N_48391);
xnor UO_937 (O_937,N_48380,N_48636);
xor UO_938 (O_938,N_48206,N_48584);
and UO_939 (O_939,N_49450,N_49805);
and UO_940 (O_940,N_47745,N_48342);
nor UO_941 (O_941,N_49939,N_48216);
and UO_942 (O_942,N_49651,N_48599);
xnor UO_943 (O_943,N_48856,N_49177);
or UO_944 (O_944,N_47796,N_48914);
or UO_945 (O_945,N_49757,N_49845);
nor UO_946 (O_946,N_49290,N_49665);
nand UO_947 (O_947,N_47943,N_49158);
nand UO_948 (O_948,N_48175,N_49606);
xnor UO_949 (O_949,N_48174,N_49560);
nand UO_950 (O_950,N_48545,N_48373);
nor UO_951 (O_951,N_47961,N_49293);
and UO_952 (O_952,N_48141,N_49600);
and UO_953 (O_953,N_49341,N_48221);
nor UO_954 (O_954,N_47939,N_48949);
and UO_955 (O_955,N_48761,N_47593);
nor UO_956 (O_956,N_49711,N_49873);
or UO_957 (O_957,N_48588,N_49648);
xnor UO_958 (O_958,N_48650,N_49189);
nor UO_959 (O_959,N_48865,N_48087);
nand UO_960 (O_960,N_49847,N_48455);
nand UO_961 (O_961,N_48941,N_48963);
and UO_962 (O_962,N_48390,N_49005);
xnor UO_963 (O_963,N_48968,N_49092);
nor UO_964 (O_964,N_49967,N_49924);
and UO_965 (O_965,N_49884,N_48807);
and UO_966 (O_966,N_49066,N_47696);
and UO_967 (O_967,N_49944,N_49486);
nor UO_968 (O_968,N_49744,N_48068);
or UO_969 (O_969,N_47690,N_47624);
or UO_970 (O_970,N_48147,N_48714);
nor UO_971 (O_971,N_47632,N_48768);
nand UO_972 (O_972,N_48403,N_49195);
nand UO_973 (O_973,N_48776,N_48459);
xnor UO_974 (O_974,N_48099,N_48313);
and UO_975 (O_975,N_49768,N_47596);
and UO_976 (O_976,N_48288,N_48679);
nand UO_977 (O_977,N_49972,N_48921);
or UO_978 (O_978,N_49072,N_49899);
nand UO_979 (O_979,N_48219,N_48516);
or UO_980 (O_980,N_48533,N_48475);
or UO_981 (O_981,N_49824,N_48048);
or UO_982 (O_982,N_47779,N_48054);
or UO_983 (O_983,N_49921,N_49525);
nor UO_984 (O_984,N_48550,N_48234);
and UO_985 (O_985,N_49826,N_47755);
and UO_986 (O_986,N_48055,N_49260);
nand UO_987 (O_987,N_48519,N_47753);
and UO_988 (O_988,N_49075,N_47899);
or UO_989 (O_989,N_48973,N_49836);
xnor UO_990 (O_990,N_47583,N_48649);
or UO_991 (O_991,N_49661,N_49453);
and UO_992 (O_992,N_49120,N_48888);
nor UO_993 (O_993,N_48820,N_47841);
and UO_994 (O_994,N_49331,N_49444);
nor UO_995 (O_995,N_49203,N_48104);
or UO_996 (O_996,N_48392,N_48881);
nand UO_997 (O_997,N_49427,N_48084);
or UO_998 (O_998,N_48273,N_48646);
xor UO_999 (O_999,N_47898,N_49790);
nand UO_1000 (O_1000,N_49337,N_48909);
xor UO_1001 (O_1001,N_49708,N_47781);
xnor UO_1002 (O_1002,N_48733,N_48956);
or UO_1003 (O_1003,N_49216,N_49472);
or UO_1004 (O_1004,N_47919,N_47743);
and UO_1005 (O_1005,N_47966,N_49446);
nor UO_1006 (O_1006,N_49000,N_48819);
or UO_1007 (O_1007,N_48377,N_49251);
nand UO_1008 (O_1008,N_49198,N_49415);
nor UO_1009 (O_1009,N_47703,N_49869);
nand UO_1010 (O_1010,N_49916,N_49751);
and UO_1011 (O_1011,N_48112,N_49119);
nand UO_1012 (O_1012,N_48122,N_49344);
or UO_1013 (O_1013,N_48906,N_48719);
xnor UO_1014 (O_1014,N_47986,N_47559);
and UO_1015 (O_1015,N_47617,N_48849);
nor UO_1016 (O_1016,N_49395,N_47693);
and UO_1017 (O_1017,N_49580,N_48631);
nand UO_1018 (O_1018,N_48036,N_49267);
and UO_1019 (O_1019,N_49660,N_49248);
or UO_1020 (O_1020,N_49173,N_48625);
xor UO_1021 (O_1021,N_48773,N_49835);
nand UO_1022 (O_1022,N_48090,N_49511);
or UO_1023 (O_1023,N_49243,N_48828);
nand UO_1024 (O_1024,N_48050,N_49957);
nand UO_1025 (O_1025,N_48322,N_48080);
nor UO_1026 (O_1026,N_47994,N_48265);
xor UO_1027 (O_1027,N_49084,N_48647);
nor UO_1028 (O_1028,N_48259,N_49292);
nand UO_1029 (O_1029,N_48915,N_48276);
or UO_1030 (O_1030,N_49059,N_49655);
and UO_1031 (O_1031,N_47526,N_49488);
and UO_1032 (O_1032,N_48780,N_48376);
nor UO_1033 (O_1033,N_48621,N_49966);
xnor UO_1034 (O_1034,N_49308,N_48118);
nor UO_1035 (O_1035,N_49523,N_48239);
or UO_1036 (O_1036,N_47613,N_47756);
and UO_1037 (O_1037,N_48871,N_49840);
and UO_1038 (O_1038,N_49993,N_49249);
and UO_1039 (O_1039,N_48138,N_49601);
or UO_1040 (O_1040,N_49036,N_48019);
and UO_1041 (O_1041,N_47808,N_49975);
or UO_1042 (O_1042,N_48241,N_47894);
or UO_1043 (O_1043,N_48618,N_49010);
and UO_1044 (O_1044,N_49239,N_49604);
and UO_1045 (O_1045,N_47868,N_47660);
and UO_1046 (O_1046,N_49766,N_48238);
nor UO_1047 (O_1047,N_48518,N_47975);
and UO_1048 (O_1048,N_48511,N_48538);
and UO_1049 (O_1049,N_47801,N_48081);
nor UO_1050 (O_1050,N_49982,N_48604);
and UO_1051 (O_1051,N_48653,N_47655);
and UO_1052 (O_1052,N_48032,N_48893);
and UO_1053 (O_1053,N_48092,N_47927);
and UO_1054 (O_1054,N_48640,N_47723);
nand UO_1055 (O_1055,N_48892,N_48785);
or UO_1056 (O_1056,N_47720,N_48061);
nand UO_1057 (O_1057,N_49908,N_49286);
nand UO_1058 (O_1058,N_48182,N_49052);
nor UO_1059 (O_1059,N_49374,N_49881);
nand UO_1060 (O_1060,N_49729,N_49369);
and UO_1061 (O_1061,N_49280,N_49639);
nor UO_1062 (O_1062,N_47558,N_48469);
or UO_1063 (O_1063,N_48751,N_49018);
xor UO_1064 (O_1064,N_49558,N_47506);
xnor UO_1065 (O_1065,N_48041,N_49963);
nor UO_1066 (O_1066,N_47932,N_47774);
and UO_1067 (O_1067,N_48583,N_48897);
and UO_1068 (O_1068,N_49519,N_49175);
and UO_1069 (O_1069,N_48887,N_49060);
and UO_1070 (O_1070,N_49043,N_48337);
xnor UO_1071 (O_1071,N_48472,N_48133);
xor UO_1072 (O_1072,N_48707,N_49926);
nand UO_1073 (O_1073,N_48155,N_48670);
nor UO_1074 (O_1074,N_49698,N_49579);
nor UO_1075 (O_1075,N_47882,N_48364);
nor UO_1076 (O_1076,N_49669,N_49136);
nor UO_1077 (O_1077,N_48513,N_47889);
xnor UO_1078 (O_1078,N_47577,N_49645);
or UO_1079 (O_1079,N_49693,N_49212);
nand UO_1080 (O_1080,N_48756,N_49878);
or UO_1081 (O_1081,N_49169,N_47724);
or UO_1082 (O_1082,N_48389,N_47503);
or UO_1083 (O_1083,N_48978,N_47714);
and UO_1084 (O_1084,N_47685,N_49940);
nor UO_1085 (O_1085,N_49261,N_49176);
nand UO_1086 (O_1086,N_47609,N_49056);
nand UO_1087 (O_1087,N_47544,N_47940);
and UO_1088 (O_1088,N_47938,N_48681);
nor UO_1089 (O_1089,N_47505,N_49476);
xnor UO_1090 (O_1090,N_49783,N_48564);
nor UO_1091 (O_1091,N_48950,N_49485);
xor UO_1092 (O_1092,N_49479,N_48547);
nand UO_1093 (O_1093,N_49382,N_49684);
nand UO_1094 (O_1094,N_48001,N_48069);
or UO_1095 (O_1095,N_49269,N_49330);
nor UO_1096 (O_1096,N_47704,N_47844);
or UO_1097 (O_1097,N_48151,N_47692);
nand UO_1098 (O_1098,N_49888,N_49336);
nand UO_1099 (O_1099,N_47643,N_49008);
nand UO_1100 (O_1100,N_48808,N_49219);
nor UO_1101 (O_1101,N_48351,N_49914);
or UO_1102 (O_1102,N_49870,N_48258);
nand UO_1103 (O_1103,N_49364,N_47926);
or UO_1104 (O_1104,N_49003,N_48116);
or UO_1105 (O_1105,N_48245,N_49240);
or UO_1106 (O_1106,N_48731,N_49351);
nor UO_1107 (O_1107,N_48227,N_48369);
nand UO_1108 (O_1108,N_47923,N_48531);
nand UO_1109 (O_1109,N_48166,N_48701);
and UO_1110 (O_1110,N_49508,N_47717);
nor UO_1111 (O_1111,N_48343,N_48005);
xnor UO_1112 (O_1112,N_48465,N_48250);
and UO_1113 (O_1113,N_49295,N_48975);
or UO_1114 (O_1114,N_49378,N_49582);
or UO_1115 (O_1115,N_49434,N_49953);
nor UO_1116 (O_1116,N_49338,N_49325);
or UO_1117 (O_1117,N_49868,N_49298);
nor UO_1118 (O_1118,N_48374,N_48388);
and UO_1119 (O_1119,N_49065,N_47776);
and UO_1120 (O_1120,N_49965,N_48117);
and UO_1121 (O_1121,N_48387,N_47531);
nor UO_1122 (O_1122,N_49809,N_49763);
or UO_1123 (O_1123,N_48832,N_49204);
xor UO_1124 (O_1124,N_48786,N_48165);
and UO_1125 (O_1125,N_49228,N_49419);
nand UO_1126 (O_1126,N_48927,N_47563);
or UO_1127 (O_1127,N_47887,N_47973);
nor UO_1128 (O_1128,N_49200,N_49875);
nor UO_1129 (O_1129,N_48911,N_49262);
xnor UO_1130 (O_1130,N_48439,N_47838);
nand UO_1131 (O_1131,N_48339,N_48913);
nand UO_1132 (O_1132,N_49622,N_49632);
or UO_1133 (O_1133,N_47736,N_49532);
and UO_1134 (O_1134,N_49068,N_49515);
nor UO_1135 (O_1135,N_47799,N_49891);
nand UO_1136 (O_1136,N_47914,N_47500);
and UO_1137 (O_1137,N_48073,N_47840);
and UO_1138 (O_1138,N_49795,N_47783);
xnor UO_1139 (O_1139,N_49867,N_49777);
or UO_1140 (O_1140,N_47821,N_48967);
or UO_1141 (O_1141,N_49709,N_48641);
nand UO_1142 (O_1142,N_48453,N_48992);
nand UO_1143 (O_1143,N_47908,N_47564);
nand UO_1144 (O_1144,N_49792,N_48708);
or UO_1145 (O_1145,N_48716,N_47936);
and UO_1146 (O_1146,N_47597,N_47603);
or UO_1147 (O_1147,N_49800,N_48792);
xor UO_1148 (O_1148,N_47922,N_47668);
nand UO_1149 (O_1149,N_47680,N_47579);
nor UO_1150 (O_1150,N_48203,N_49235);
nand UO_1151 (O_1151,N_48663,N_49192);
and UO_1152 (O_1152,N_47947,N_49393);
or UO_1153 (O_1153,N_48196,N_49359);
and UO_1154 (O_1154,N_49843,N_48575);
nand UO_1155 (O_1155,N_49067,N_48622);
nand UO_1156 (O_1156,N_47661,N_49105);
or UO_1157 (O_1157,N_49142,N_47857);
xnor UO_1158 (O_1158,N_47589,N_47820);
nand UO_1159 (O_1159,N_49435,N_49618);
or UO_1160 (O_1160,N_48682,N_49559);
xor UO_1161 (O_1161,N_48341,N_47514);
or UO_1162 (O_1162,N_48416,N_49644);
nand UO_1163 (O_1163,N_49490,N_48803);
or UO_1164 (O_1164,N_48579,N_49471);
or UO_1165 (O_1165,N_49819,N_48520);
and UO_1166 (O_1166,N_49222,N_49536);
nor UO_1167 (O_1167,N_49334,N_49707);
or UO_1168 (O_1168,N_47614,N_48143);
or UO_1169 (O_1169,N_49491,N_49302);
nand UO_1170 (O_1170,N_48525,N_48539);
or UO_1171 (O_1171,N_49649,N_49089);
xnor UO_1172 (O_1172,N_48022,N_48304);
xnor UO_1173 (O_1173,N_49948,N_49482);
xor UO_1174 (O_1174,N_49152,N_48356);
nand UO_1175 (O_1175,N_49764,N_49126);
xnor UO_1176 (O_1176,N_49732,N_47676);
and UO_1177 (O_1177,N_49379,N_48144);
xor UO_1178 (O_1178,N_49102,N_48812);
and UO_1179 (O_1179,N_48498,N_49521);
and UO_1180 (O_1180,N_48810,N_48814);
or UO_1181 (O_1181,N_47950,N_48823);
and UO_1182 (O_1182,N_49110,N_48517);
nand UO_1183 (O_1183,N_49220,N_47823);
nand UO_1184 (O_1184,N_49265,N_48648);
and UO_1185 (O_1185,N_48623,N_48371);
or UO_1186 (O_1186,N_49998,N_49123);
nand UO_1187 (O_1187,N_48008,N_48397);
xor UO_1188 (O_1188,N_49048,N_47722);
nor UO_1189 (O_1189,N_49904,N_49417);
nor UO_1190 (O_1190,N_48394,N_48740);
xor UO_1191 (O_1191,N_48235,N_49470);
nand UO_1192 (O_1192,N_48986,N_48354);
and UO_1193 (O_1193,N_49429,N_49121);
nor UO_1194 (O_1194,N_48172,N_48125);
nor UO_1195 (O_1195,N_48802,N_48149);
or UO_1196 (O_1196,N_48433,N_48680);
or UO_1197 (O_1197,N_48587,N_49209);
or UO_1198 (O_1198,N_49460,N_48434);
and UO_1199 (O_1199,N_49015,N_47976);
and UO_1200 (O_1200,N_49418,N_47830);
nor UO_1201 (O_1201,N_48729,N_49872);
nor UO_1202 (O_1202,N_49082,N_48891);
or UO_1203 (O_1203,N_47684,N_49761);
nand UO_1204 (O_1204,N_47549,N_47810);
and UO_1205 (O_1205,N_48608,N_47533);
or UO_1206 (O_1206,N_48365,N_48633);
and UO_1207 (O_1207,N_48561,N_47622);
or UO_1208 (O_1208,N_48204,N_47529);
and UO_1209 (O_1209,N_48779,N_48523);
and UO_1210 (O_1210,N_49747,N_48330);
and UO_1211 (O_1211,N_47747,N_49289);
xnor UO_1212 (O_1212,N_49319,N_48010);
nor UO_1213 (O_1213,N_48131,N_47998);
or UO_1214 (O_1214,N_48198,N_48044);
nor UO_1215 (O_1215,N_47785,N_49061);
nor UO_1216 (O_1216,N_47683,N_49391);
and UO_1217 (O_1217,N_49787,N_49799);
nand UO_1218 (O_1218,N_47972,N_47846);
or UO_1219 (O_1219,N_48411,N_47615);
or UO_1220 (O_1220,N_49933,N_48990);
or UO_1221 (O_1221,N_49529,N_48930);
nor UO_1222 (O_1222,N_49206,N_49164);
nor UO_1223 (O_1223,N_47924,N_49483);
or UO_1224 (O_1224,N_48419,N_49980);
nor UO_1225 (O_1225,N_49781,N_48293);
or UO_1226 (O_1226,N_49443,N_48447);
or UO_1227 (O_1227,N_49394,N_48254);
nand UO_1228 (O_1228,N_48082,N_47512);
and UO_1229 (O_1229,N_49196,N_48946);
nor UO_1230 (O_1230,N_49951,N_48850);
nand UO_1231 (O_1231,N_48543,N_49798);
nand UO_1232 (O_1232,N_49132,N_48855);
or UO_1233 (O_1233,N_49050,N_48107);
or UO_1234 (O_1234,N_48426,N_48957);
nor UO_1235 (O_1235,N_49502,N_49103);
nand UO_1236 (O_1236,N_49796,N_49469);
xnor UO_1237 (O_1237,N_49107,N_48070);
nand UO_1238 (O_1238,N_49455,N_48568);
nand UO_1239 (O_1239,N_49917,N_48577);
nor UO_1240 (O_1240,N_49646,N_48292);
nand UO_1241 (O_1241,N_48626,N_48291);
nor UO_1242 (O_1242,N_47578,N_49885);
nand UO_1243 (O_1243,N_49877,N_49148);
or UO_1244 (O_1244,N_49406,N_49657);
nor UO_1245 (O_1245,N_47907,N_49992);
nor UO_1246 (O_1246,N_49743,N_48686);
nand UO_1247 (O_1247,N_48600,N_49785);
xor UO_1248 (O_1248,N_49304,N_49205);
and UO_1249 (O_1249,N_48352,N_49347);
nor UO_1250 (O_1250,N_49182,N_48899);
and UO_1251 (O_1251,N_49803,N_47656);
or UO_1252 (O_1252,N_49177,N_49891);
nand UO_1253 (O_1253,N_49071,N_48594);
and UO_1254 (O_1254,N_49579,N_48284);
or UO_1255 (O_1255,N_48265,N_48474);
or UO_1256 (O_1256,N_48063,N_49177);
xor UO_1257 (O_1257,N_48156,N_48088);
and UO_1258 (O_1258,N_47557,N_48883);
and UO_1259 (O_1259,N_47999,N_49520);
and UO_1260 (O_1260,N_48814,N_48540);
and UO_1261 (O_1261,N_49545,N_47864);
and UO_1262 (O_1262,N_48913,N_49388);
and UO_1263 (O_1263,N_49654,N_48471);
nand UO_1264 (O_1264,N_48637,N_48349);
and UO_1265 (O_1265,N_49820,N_47812);
and UO_1266 (O_1266,N_49796,N_48584);
or UO_1267 (O_1267,N_49619,N_48691);
or UO_1268 (O_1268,N_49673,N_49689);
nand UO_1269 (O_1269,N_47524,N_48651);
or UO_1270 (O_1270,N_48636,N_49393);
and UO_1271 (O_1271,N_48295,N_49422);
or UO_1272 (O_1272,N_48196,N_47754);
and UO_1273 (O_1273,N_49378,N_49478);
and UO_1274 (O_1274,N_47636,N_49160);
or UO_1275 (O_1275,N_49396,N_48632);
nor UO_1276 (O_1276,N_48073,N_47953);
and UO_1277 (O_1277,N_48485,N_48785);
nor UO_1278 (O_1278,N_49371,N_49283);
xnor UO_1279 (O_1279,N_49052,N_47847);
and UO_1280 (O_1280,N_48697,N_48504);
xnor UO_1281 (O_1281,N_49764,N_48118);
xor UO_1282 (O_1282,N_48166,N_48408);
and UO_1283 (O_1283,N_48482,N_48688);
and UO_1284 (O_1284,N_47868,N_49222);
nand UO_1285 (O_1285,N_48726,N_48685);
and UO_1286 (O_1286,N_49802,N_48475);
or UO_1287 (O_1287,N_47805,N_49015);
and UO_1288 (O_1288,N_48647,N_49186);
nor UO_1289 (O_1289,N_49768,N_49322);
nand UO_1290 (O_1290,N_49310,N_48644);
nor UO_1291 (O_1291,N_47624,N_47750);
and UO_1292 (O_1292,N_48668,N_49743);
xnor UO_1293 (O_1293,N_48534,N_48869);
or UO_1294 (O_1294,N_49589,N_49738);
or UO_1295 (O_1295,N_48602,N_48901);
nor UO_1296 (O_1296,N_47786,N_48315);
nor UO_1297 (O_1297,N_49582,N_47578);
xnor UO_1298 (O_1298,N_49848,N_48326);
and UO_1299 (O_1299,N_49608,N_49892);
or UO_1300 (O_1300,N_48599,N_47532);
and UO_1301 (O_1301,N_48560,N_49056);
and UO_1302 (O_1302,N_48113,N_49923);
and UO_1303 (O_1303,N_49170,N_49937);
or UO_1304 (O_1304,N_48114,N_49891);
or UO_1305 (O_1305,N_49233,N_48172);
and UO_1306 (O_1306,N_47935,N_47626);
nor UO_1307 (O_1307,N_49630,N_48691);
or UO_1308 (O_1308,N_47654,N_48447);
or UO_1309 (O_1309,N_48668,N_49466);
nor UO_1310 (O_1310,N_47533,N_48335);
or UO_1311 (O_1311,N_47697,N_49558);
and UO_1312 (O_1312,N_48579,N_48687);
and UO_1313 (O_1313,N_47974,N_47929);
or UO_1314 (O_1314,N_49851,N_48457);
and UO_1315 (O_1315,N_49530,N_47578);
or UO_1316 (O_1316,N_48456,N_49008);
nand UO_1317 (O_1317,N_47887,N_48963);
or UO_1318 (O_1318,N_47997,N_49931);
nand UO_1319 (O_1319,N_49586,N_47603);
and UO_1320 (O_1320,N_49546,N_49715);
and UO_1321 (O_1321,N_49257,N_48224);
and UO_1322 (O_1322,N_48883,N_49513);
nor UO_1323 (O_1323,N_47651,N_47502);
nand UO_1324 (O_1324,N_49236,N_49566);
and UO_1325 (O_1325,N_49887,N_49193);
xor UO_1326 (O_1326,N_49304,N_48205);
and UO_1327 (O_1327,N_47751,N_49892);
or UO_1328 (O_1328,N_49385,N_47787);
nand UO_1329 (O_1329,N_49091,N_48123);
and UO_1330 (O_1330,N_47568,N_47879);
and UO_1331 (O_1331,N_48090,N_48442);
nand UO_1332 (O_1332,N_47711,N_49677);
nand UO_1333 (O_1333,N_49178,N_49243);
nand UO_1334 (O_1334,N_49506,N_49147);
nand UO_1335 (O_1335,N_48841,N_48290);
and UO_1336 (O_1336,N_48262,N_49117);
or UO_1337 (O_1337,N_48196,N_47812);
or UO_1338 (O_1338,N_48430,N_49515);
nand UO_1339 (O_1339,N_49623,N_48582);
or UO_1340 (O_1340,N_47764,N_48663);
nor UO_1341 (O_1341,N_49831,N_47579);
nor UO_1342 (O_1342,N_49623,N_49177);
nand UO_1343 (O_1343,N_49517,N_48827);
xor UO_1344 (O_1344,N_49361,N_47829);
nor UO_1345 (O_1345,N_49060,N_49248);
nand UO_1346 (O_1346,N_48535,N_49220);
nor UO_1347 (O_1347,N_49505,N_49627);
nand UO_1348 (O_1348,N_49662,N_48448);
nor UO_1349 (O_1349,N_47919,N_48465);
nand UO_1350 (O_1350,N_48850,N_49748);
xor UO_1351 (O_1351,N_49288,N_48612);
nor UO_1352 (O_1352,N_48129,N_48809);
and UO_1353 (O_1353,N_49511,N_47733);
xor UO_1354 (O_1354,N_47824,N_49014);
and UO_1355 (O_1355,N_48590,N_49710);
or UO_1356 (O_1356,N_47968,N_48796);
nor UO_1357 (O_1357,N_47885,N_49815);
nand UO_1358 (O_1358,N_49940,N_49478);
or UO_1359 (O_1359,N_47556,N_47824);
and UO_1360 (O_1360,N_49881,N_48957);
and UO_1361 (O_1361,N_49292,N_47556);
nor UO_1362 (O_1362,N_48396,N_48448);
and UO_1363 (O_1363,N_47953,N_48037);
and UO_1364 (O_1364,N_49760,N_49841);
xnor UO_1365 (O_1365,N_49372,N_47656);
and UO_1366 (O_1366,N_48453,N_47924);
nand UO_1367 (O_1367,N_49854,N_49720);
or UO_1368 (O_1368,N_49477,N_49412);
or UO_1369 (O_1369,N_48814,N_48895);
and UO_1370 (O_1370,N_49167,N_48544);
nand UO_1371 (O_1371,N_48418,N_48432);
nor UO_1372 (O_1372,N_47959,N_49882);
nor UO_1373 (O_1373,N_48514,N_49658);
nand UO_1374 (O_1374,N_48752,N_47753);
and UO_1375 (O_1375,N_48133,N_48064);
or UO_1376 (O_1376,N_49029,N_49109);
or UO_1377 (O_1377,N_49157,N_48585);
nor UO_1378 (O_1378,N_47565,N_48929);
nor UO_1379 (O_1379,N_49303,N_49121);
xor UO_1380 (O_1380,N_48369,N_49076);
nand UO_1381 (O_1381,N_48350,N_48750);
xor UO_1382 (O_1382,N_49050,N_48032);
or UO_1383 (O_1383,N_48154,N_48911);
or UO_1384 (O_1384,N_49450,N_49083);
or UO_1385 (O_1385,N_47864,N_48709);
or UO_1386 (O_1386,N_48381,N_49963);
xnor UO_1387 (O_1387,N_49534,N_49306);
nor UO_1388 (O_1388,N_49268,N_48194);
nor UO_1389 (O_1389,N_48620,N_49780);
nor UO_1390 (O_1390,N_48672,N_48548);
and UO_1391 (O_1391,N_49828,N_49127);
or UO_1392 (O_1392,N_47550,N_49513);
nor UO_1393 (O_1393,N_47966,N_47587);
nand UO_1394 (O_1394,N_49634,N_48638);
nor UO_1395 (O_1395,N_47693,N_48923);
or UO_1396 (O_1396,N_49883,N_48401);
nor UO_1397 (O_1397,N_47552,N_49494);
nor UO_1398 (O_1398,N_49941,N_48192);
nor UO_1399 (O_1399,N_48161,N_48227);
nand UO_1400 (O_1400,N_48494,N_49804);
and UO_1401 (O_1401,N_49326,N_49867);
nand UO_1402 (O_1402,N_48664,N_49474);
nor UO_1403 (O_1403,N_49891,N_47602);
or UO_1404 (O_1404,N_49440,N_49029);
nand UO_1405 (O_1405,N_49920,N_49371);
nand UO_1406 (O_1406,N_47588,N_49253);
and UO_1407 (O_1407,N_48352,N_49062);
and UO_1408 (O_1408,N_48259,N_48986);
and UO_1409 (O_1409,N_48727,N_49454);
nor UO_1410 (O_1410,N_49180,N_47600);
xnor UO_1411 (O_1411,N_48639,N_48997);
and UO_1412 (O_1412,N_48740,N_49912);
nand UO_1413 (O_1413,N_49805,N_47722);
nand UO_1414 (O_1414,N_47516,N_48917);
nand UO_1415 (O_1415,N_49954,N_49343);
xnor UO_1416 (O_1416,N_47748,N_49729);
or UO_1417 (O_1417,N_49150,N_49959);
and UO_1418 (O_1418,N_49031,N_47556);
and UO_1419 (O_1419,N_47614,N_48790);
nand UO_1420 (O_1420,N_49662,N_49728);
nand UO_1421 (O_1421,N_47775,N_49091);
or UO_1422 (O_1422,N_49758,N_49500);
nand UO_1423 (O_1423,N_49569,N_48286);
and UO_1424 (O_1424,N_48850,N_49095);
nand UO_1425 (O_1425,N_49223,N_48478);
and UO_1426 (O_1426,N_49826,N_49649);
or UO_1427 (O_1427,N_48444,N_49384);
nor UO_1428 (O_1428,N_49543,N_48857);
nand UO_1429 (O_1429,N_49195,N_49986);
nor UO_1430 (O_1430,N_48919,N_48965);
nor UO_1431 (O_1431,N_48056,N_48384);
and UO_1432 (O_1432,N_49985,N_48443);
nor UO_1433 (O_1433,N_49331,N_48467);
or UO_1434 (O_1434,N_48698,N_47629);
and UO_1435 (O_1435,N_49590,N_47740);
nor UO_1436 (O_1436,N_48676,N_47642);
nand UO_1437 (O_1437,N_48615,N_49341);
and UO_1438 (O_1438,N_48645,N_49428);
and UO_1439 (O_1439,N_49031,N_49601);
nor UO_1440 (O_1440,N_49987,N_49197);
nand UO_1441 (O_1441,N_48636,N_47794);
nor UO_1442 (O_1442,N_47748,N_48326);
or UO_1443 (O_1443,N_49180,N_49381);
or UO_1444 (O_1444,N_49135,N_49940);
nand UO_1445 (O_1445,N_49009,N_49896);
and UO_1446 (O_1446,N_49651,N_48594);
or UO_1447 (O_1447,N_49423,N_49750);
xnor UO_1448 (O_1448,N_49692,N_48249);
and UO_1449 (O_1449,N_49149,N_47872);
nand UO_1450 (O_1450,N_47788,N_49179);
and UO_1451 (O_1451,N_48036,N_47801);
xnor UO_1452 (O_1452,N_49263,N_49765);
and UO_1453 (O_1453,N_47591,N_48129);
nor UO_1454 (O_1454,N_48677,N_47842);
nor UO_1455 (O_1455,N_48429,N_49873);
or UO_1456 (O_1456,N_49023,N_49285);
nand UO_1457 (O_1457,N_47564,N_47575);
xnor UO_1458 (O_1458,N_47529,N_49989);
and UO_1459 (O_1459,N_48513,N_49873);
and UO_1460 (O_1460,N_48497,N_49469);
nand UO_1461 (O_1461,N_47682,N_48429);
and UO_1462 (O_1462,N_47626,N_49622);
and UO_1463 (O_1463,N_48795,N_49607);
nand UO_1464 (O_1464,N_48543,N_49878);
nand UO_1465 (O_1465,N_48647,N_48836);
or UO_1466 (O_1466,N_49540,N_48913);
or UO_1467 (O_1467,N_49462,N_48985);
or UO_1468 (O_1468,N_49180,N_47789);
nor UO_1469 (O_1469,N_49396,N_48573);
and UO_1470 (O_1470,N_48155,N_48055);
xor UO_1471 (O_1471,N_49962,N_48919);
nand UO_1472 (O_1472,N_49417,N_48468);
or UO_1473 (O_1473,N_48943,N_49938);
or UO_1474 (O_1474,N_49531,N_48133);
nand UO_1475 (O_1475,N_49551,N_49810);
nor UO_1476 (O_1476,N_48299,N_48520);
or UO_1477 (O_1477,N_48911,N_47559);
nor UO_1478 (O_1478,N_47890,N_48120);
nor UO_1479 (O_1479,N_48714,N_49600);
and UO_1480 (O_1480,N_49110,N_47582);
nor UO_1481 (O_1481,N_49411,N_47517);
and UO_1482 (O_1482,N_49398,N_48698);
and UO_1483 (O_1483,N_47722,N_47924);
or UO_1484 (O_1484,N_48894,N_47578);
nand UO_1485 (O_1485,N_48434,N_49659);
nor UO_1486 (O_1486,N_47927,N_47852);
or UO_1487 (O_1487,N_49940,N_49668);
or UO_1488 (O_1488,N_49714,N_49349);
or UO_1489 (O_1489,N_48171,N_47598);
nand UO_1490 (O_1490,N_49780,N_47656);
and UO_1491 (O_1491,N_48128,N_49328);
nand UO_1492 (O_1492,N_49314,N_49739);
or UO_1493 (O_1493,N_48888,N_47522);
nor UO_1494 (O_1494,N_49190,N_49968);
nor UO_1495 (O_1495,N_49842,N_49630);
or UO_1496 (O_1496,N_48034,N_48024);
or UO_1497 (O_1497,N_49480,N_49609);
and UO_1498 (O_1498,N_47623,N_48785);
nor UO_1499 (O_1499,N_47617,N_49869);
and UO_1500 (O_1500,N_48146,N_49012);
nor UO_1501 (O_1501,N_48447,N_48970);
nor UO_1502 (O_1502,N_48047,N_47930);
or UO_1503 (O_1503,N_49809,N_48522);
xnor UO_1504 (O_1504,N_49363,N_47842);
or UO_1505 (O_1505,N_48392,N_49589);
or UO_1506 (O_1506,N_48792,N_48330);
nor UO_1507 (O_1507,N_48372,N_48727);
nand UO_1508 (O_1508,N_49348,N_47852);
nor UO_1509 (O_1509,N_47541,N_48680);
and UO_1510 (O_1510,N_49209,N_49191);
and UO_1511 (O_1511,N_49729,N_49379);
and UO_1512 (O_1512,N_48675,N_49652);
or UO_1513 (O_1513,N_49270,N_49226);
nor UO_1514 (O_1514,N_49558,N_48918);
or UO_1515 (O_1515,N_49917,N_48676);
nor UO_1516 (O_1516,N_49357,N_47518);
nand UO_1517 (O_1517,N_49882,N_48538);
or UO_1518 (O_1518,N_49116,N_49820);
xnor UO_1519 (O_1519,N_49403,N_49054);
nor UO_1520 (O_1520,N_49320,N_49008);
nand UO_1521 (O_1521,N_49478,N_49048);
xor UO_1522 (O_1522,N_47591,N_48408);
xnor UO_1523 (O_1523,N_49441,N_48428);
nor UO_1524 (O_1524,N_47625,N_49916);
and UO_1525 (O_1525,N_49184,N_49210);
and UO_1526 (O_1526,N_48522,N_47897);
nor UO_1527 (O_1527,N_49722,N_48512);
and UO_1528 (O_1528,N_49343,N_48617);
nor UO_1529 (O_1529,N_49515,N_49614);
and UO_1530 (O_1530,N_49063,N_49825);
or UO_1531 (O_1531,N_47543,N_48907);
xnor UO_1532 (O_1532,N_47635,N_49130);
nand UO_1533 (O_1533,N_48935,N_49513);
nand UO_1534 (O_1534,N_48494,N_48490);
nor UO_1535 (O_1535,N_49327,N_47840);
nor UO_1536 (O_1536,N_49061,N_48359);
or UO_1537 (O_1537,N_48370,N_49136);
and UO_1538 (O_1538,N_49547,N_49889);
and UO_1539 (O_1539,N_49972,N_49026);
and UO_1540 (O_1540,N_48386,N_48299);
or UO_1541 (O_1541,N_49536,N_49963);
and UO_1542 (O_1542,N_47573,N_48617);
and UO_1543 (O_1543,N_48429,N_48775);
xnor UO_1544 (O_1544,N_49913,N_49943);
nor UO_1545 (O_1545,N_47598,N_47542);
nand UO_1546 (O_1546,N_47957,N_47846);
and UO_1547 (O_1547,N_47674,N_48622);
xnor UO_1548 (O_1548,N_48862,N_49878);
nand UO_1549 (O_1549,N_49412,N_49847);
nand UO_1550 (O_1550,N_49488,N_48823);
or UO_1551 (O_1551,N_48096,N_49907);
nand UO_1552 (O_1552,N_48075,N_48170);
xnor UO_1553 (O_1553,N_47682,N_48381);
and UO_1554 (O_1554,N_48506,N_49913);
nand UO_1555 (O_1555,N_48004,N_49561);
and UO_1556 (O_1556,N_48153,N_48334);
and UO_1557 (O_1557,N_48629,N_48286);
or UO_1558 (O_1558,N_47586,N_48592);
or UO_1559 (O_1559,N_47745,N_48595);
xnor UO_1560 (O_1560,N_49329,N_48160);
nand UO_1561 (O_1561,N_48793,N_49392);
nand UO_1562 (O_1562,N_49825,N_48072);
nand UO_1563 (O_1563,N_48886,N_48747);
nand UO_1564 (O_1564,N_48599,N_48571);
and UO_1565 (O_1565,N_48785,N_47825);
or UO_1566 (O_1566,N_49353,N_48295);
nor UO_1567 (O_1567,N_47636,N_49489);
or UO_1568 (O_1568,N_49373,N_47934);
or UO_1569 (O_1569,N_47930,N_48580);
or UO_1570 (O_1570,N_49303,N_48112);
or UO_1571 (O_1571,N_48592,N_49614);
xnor UO_1572 (O_1572,N_48781,N_49437);
nor UO_1573 (O_1573,N_49070,N_48582);
and UO_1574 (O_1574,N_48514,N_48133);
or UO_1575 (O_1575,N_49951,N_48627);
and UO_1576 (O_1576,N_48919,N_49952);
and UO_1577 (O_1577,N_49858,N_47980);
nand UO_1578 (O_1578,N_47740,N_49508);
xor UO_1579 (O_1579,N_48611,N_48582);
nand UO_1580 (O_1580,N_49650,N_49880);
xnor UO_1581 (O_1581,N_47736,N_48660);
nor UO_1582 (O_1582,N_49086,N_48935);
or UO_1583 (O_1583,N_48291,N_48374);
nor UO_1584 (O_1584,N_49686,N_48697);
and UO_1585 (O_1585,N_49801,N_47767);
and UO_1586 (O_1586,N_48918,N_49145);
nand UO_1587 (O_1587,N_49289,N_48395);
nor UO_1588 (O_1588,N_49932,N_49204);
nor UO_1589 (O_1589,N_47920,N_47894);
and UO_1590 (O_1590,N_48985,N_48778);
nor UO_1591 (O_1591,N_48535,N_49718);
nand UO_1592 (O_1592,N_49291,N_49258);
nor UO_1593 (O_1593,N_48833,N_49955);
xor UO_1594 (O_1594,N_48408,N_49420);
nand UO_1595 (O_1595,N_48120,N_48551);
nand UO_1596 (O_1596,N_49464,N_49612);
and UO_1597 (O_1597,N_48217,N_47861);
nor UO_1598 (O_1598,N_49581,N_49549);
nand UO_1599 (O_1599,N_48382,N_49402);
or UO_1600 (O_1600,N_48170,N_49830);
or UO_1601 (O_1601,N_49812,N_49925);
or UO_1602 (O_1602,N_48642,N_48274);
or UO_1603 (O_1603,N_49321,N_48889);
xor UO_1604 (O_1604,N_49345,N_47691);
or UO_1605 (O_1605,N_48562,N_48798);
xor UO_1606 (O_1606,N_48793,N_49370);
and UO_1607 (O_1607,N_48491,N_49211);
nand UO_1608 (O_1608,N_48851,N_49081);
or UO_1609 (O_1609,N_48194,N_48101);
nor UO_1610 (O_1610,N_47553,N_48067);
xor UO_1611 (O_1611,N_49770,N_48621);
nor UO_1612 (O_1612,N_49509,N_49711);
nor UO_1613 (O_1613,N_49165,N_48971);
and UO_1614 (O_1614,N_49224,N_49858);
and UO_1615 (O_1615,N_49327,N_47999);
and UO_1616 (O_1616,N_48444,N_49438);
or UO_1617 (O_1617,N_49111,N_49033);
xnor UO_1618 (O_1618,N_47966,N_47625);
or UO_1619 (O_1619,N_48912,N_48364);
nor UO_1620 (O_1620,N_48751,N_48651);
nand UO_1621 (O_1621,N_49361,N_49931);
nor UO_1622 (O_1622,N_49273,N_48008);
nor UO_1623 (O_1623,N_48441,N_49038);
nor UO_1624 (O_1624,N_48311,N_48095);
or UO_1625 (O_1625,N_48801,N_48280);
or UO_1626 (O_1626,N_49266,N_49051);
nand UO_1627 (O_1627,N_49375,N_48400);
nand UO_1628 (O_1628,N_48191,N_47627);
nor UO_1629 (O_1629,N_47776,N_49356);
nand UO_1630 (O_1630,N_47504,N_49580);
or UO_1631 (O_1631,N_49430,N_49991);
or UO_1632 (O_1632,N_48534,N_49528);
xnor UO_1633 (O_1633,N_48138,N_48481);
and UO_1634 (O_1634,N_49892,N_49223);
and UO_1635 (O_1635,N_49737,N_49420);
and UO_1636 (O_1636,N_47840,N_48612);
and UO_1637 (O_1637,N_49218,N_47563);
nor UO_1638 (O_1638,N_47620,N_49797);
nor UO_1639 (O_1639,N_48378,N_49895);
nor UO_1640 (O_1640,N_48972,N_49951);
or UO_1641 (O_1641,N_47589,N_48317);
nor UO_1642 (O_1642,N_47660,N_49146);
nor UO_1643 (O_1643,N_49730,N_48176);
nor UO_1644 (O_1644,N_48225,N_49737);
and UO_1645 (O_1645,N_49591,N_48260);
and UO_1646 (O_1646,N_47575,N_49296);
and UO_1647 (O_1647,N_49306,N_48576);
or UO_1648 (O_1648,N_48030,N_47712);
xnor UO_1649 (O_1649,N_48758,N_49880);
nor UO_1650 (O_1650,N_48014,N_49093);
nand UO_1651 (O_1651,N_47907,N_49480);
nand UO_1652 (O_1652,N_48729,N_49987);
xnor UO_1653 (O_1653,N_48769,N_48050);
nor UO_1654 (O_1654,N_49457,N_49327);
nand UO_1655 (O_1655,N_49405,N_48650);
or UO_1656 (O_1656,N_49903,N_48974);
xor UO_1657 (O_1657,N_48681,N_48278);
xnor UO_1658 (O_1658,N_47768,N_47552);
xor UO_1659 (O_1659,N_49416,N_49013);
nor UO_1660 (O_1660,N_48664,N_48389);
xnor UO_1661 (O_1661,N_49414,N_47733);
or UO_1662 (O_1662,N_48675,N_48903);
xnor UO_1663 (O_1663,N_49009,N_48408);
or UO_1664 (O_1664,N_49243,N_47537);
nand UO_1665 (O_1665,N_49854,N_48541);
nand UO_1666 (O_1666,N_49357,N_48384);
nand UO_1667 (O_1667,N_49722,N_49580);
nand UO_1668 (O_1668,N_48906,N_48778);
nand UO_1669 (O_1669,N_49474,N_49016);
xnor UO_1670 (O_1670,N_48408,N_48911);
nand UO_1671 (O_1671,N_48259,N_48270);
nand UO_1672 (O_1672,N_49772,N_48376);
nor UO_1673 (O_1673,N_48540,N_48141);
or UO_1674 (O_1674,N_49472,N_49604);
or UO_1675 (O_1675,N_48102,N_49066);
nor UO_1676 (O_1676,N_47957,N_49974);
xor UO_1677 (O_1677,N_47831,N_49691);
nor UO_1678 (O_1678,N_49997,N_49898);
nor UO_1679 (O_1679,N_49427,N_47591);
or UO_1680 (O_1680,N_49896,N_47693);
xor UO_1681 (O_1681,N_48346,N_49684);
or UO_1682 (O_1682,N_49048,N_49945);
or UO_1683 (O_1683,N_47580,N_49672);
nand UO_1684 (O_1684,N_47917,N_47690);
and UO_1685 (O_1685,N_49071,N_49183);
and UO_1686 (O_1686,N_48563,N_47864);
or UO_1687 (O_1687,N_48697,N_47671);
and UO_1688 (O_1688,N_48243,N_49552);
nor UO_1689 (O_1689,N_47916,N_48447);
or UO_1690 (O_1690,N_47515,N_49463);
and UO_1691 (O_1691,N_48514,N_48943);
nor UO_1692 (O_1692,N_47507,N_48643);
and UO_1693 (O_1693,N_48253,N_49640);
xor UO_1694 (O_1694,N_48851,N_47533);
or UO_1695 (O_1695,N_47523,N_48548);
or UO_1696 (O_1696,N_48983,N_49132);
nor UO_1697 (O_1697,N_49275,N_47930);
and UO_1698 (O_1698,N_47590,N_49309);
nor UO_1699 (O_1699,N_49374,N_49081);
nor UO_1700 (O_1700,N_48069,N_48704);
xnor UO_1701 (O_1701,N_48485,N_48609);
or UO_1702 (O_1702,N_49604,N_48936);
nand UO_1703 (O_1703,N_48591,N_48249);
nand UO_1704 (O_1704,N_48464,N_49256);
and UO_1705 (O_1705,N_47672,N_49561);
xnor UO_1706 (O_1706,N_48104,N_49441);
nand UO_1707 (O_1707,N_47507,N_48309);
nand UO_1708 (O_1708,N_49395,N_48606);
xor UO_1709 (O_1709,N_48652,N_49588);
nand UO_1710 (O_1710,N_49958,N_49223);
nor UO_1711 (O_1711,N_49358,N_49375);
nor UO_1712 (O_1712,N_47794,N_48381);
and UO_1713 (O_1713,N_47529,N_47859);
or UO_1714 (O_1714,N_49193,N_49634);
or UO_1715 (O_1715,N_49572,N_49614);
nand UO_1716 (O_1716,N_48687,N_48296);
xnor UO_1717 (O_1717,N_48196,N_49468);
and UO_1718 (O_1718,N_48787,N_48219);
nand UO_1719 (O_1719,N_47899,N_47698);
nand UO_1720 (O_1720,N_49648,N_48771);
and UO_1721 (O_1721,N_49804,N_49162);
nor UO_1722 (O_1722,N_47810,N_49220);
and UO_1723 (O_1723,N_48156,N_49665);
nand UO_1724 (O_1724,N_49916,N_48434);
or UO_1725 (O_1725,N_49892,N_49568);
and UO_1726 (O_1726,N_49720,N_48814);
and UO_1727 (O_1727,N_48935,N_47884);
or UO_1728 (O_1728,N_47524,N_48508);
nor UO_1729 (O_1729,N_48032,N_49643);
nand UO_1730 (O_1730,N_49938,N_49426);
nor UO_1731 (O_1731,N_48035,N_47621);
nor UO_1732 (O_1732,N_47569,N_49473);
nor UO_1733 (O_1733,N_48538,N_48591);
or UO_1734 (O_1734,N_48920,N_48496);
xnor UO_1735 (O_1735,N_48590,N_49604);
and UO_1736 (O_1736,N_47518,N_49290);
or UO_1737 (O_1737,N_47688,N_49777);
nor UO_1738 (O_1738,N_49487,N_49572);
and UO_1739 (O_1739,N_48869,N_48958);
or UO_1740 (O_1740,N_48793,N_48429);
xnor UO_1741 (O_1741,N_49694,N_49323);
nand UO_1742 (O_1742,N_49623,N_47743);
or UO_1743 (O_1743,N_49514,N_48944);
and UO_1744 (O_1744,N_48650,N_49713);
or UO_1745 (O_1745,N_48207,N_49036);
and UO_1746 (O_1746,N_48642,N_49833);
nand UO_1747 (O_1747,N_47671,N_48874);
or UO_1748 (O_1748,N_49061,N_49245);
or UO_1749 (O_1749,N_47678,N_48714);
nand UO_1750 (O_1750,N_48265,N_48387);
nand UO_1751 (O_1751,N_48614,N_49217);
and UO_1752 (O_1752,N_48668,N_47742);
and UO_1753 (O_1753,N_47525,N_49207);
nand UO_1754 (O_1754,N_49241,N_48747);
nor UO_1755 (O_1755,N_48557,N_49711);
and UO_1756 (O_1756,N_48195,N_47947);
or UO_1757 (O_1757,N_48532,N_49357);
and UO_1758 (O_1758,N_48859,N_49050);
nand UO_1759 (O_1759,N_47836,N_49574);
nor UO_1760 (O_1760,N_49624,N_49161);
or UO_1761 (O_1761,N_48055,N_48604);
and UO_1762 (O_1762,N_47959,N_49342);
nor UO_1763 (O_1763,N_48279,N_49323);
and UO_1764 (O_1764,N_49852,N_49357);
xor UO_1765 (O_1765,N_49913,N_49370);
and UO_1766 (O_1766,N_49385,N_47692);
nand UO_1767 (O_1767,N_48489,N_47882);
nand UO_1768 (O_1768,N_47828,N_48526);
nand UO_1769 (O_1769,N_49153,N_49387);
or UO_1770 (O_1770,N_48393,N_49077);
or UO_1771 (O_1771,N_49300,N_48545);
xor UO_1772 (O_1772,N_49587,N_47793);
and UO_1773 (O_1773,N_47646,N_47971);
nand UO_1774 (O_1774,N_48078,N_49793);
and UO_1775 (O_1775,N_47975,N_49876);
or UO_1776 (O_1776,N_47735,N_49911);
nand UO_1777 (O_1777,N_48025,N_48757);
xor UO_1778 (O_1778,N_48019,N_48662);
nor UO_1779 (O_1779,N_48170,N_49097);
nand UO_1780 (O_1780,N_49907,N_48820);
and UO_1781 (O_1781,N_49661,N_47510);
and UO_1782 (O_1782,N_48002,N_47948);
nand UO_1783 (O_1783,N_48812,N_48095);
and UO_1784 (O_1784,N_49105,N_49181);
and UO_1785 (O_1785,N_47872,N_47604);
nand UO_1786 (O_1786,N_48770,N_48774);
and UO_1787 (O_1787,N_47572,N_49213);
or UO_1788 (O_1788,N_49294,N_47578);
and UO_1789 (O_1789,N_49122,N_48217);
nand UO_1790 (O_1790,N_49817,N_47858);
nor UO_1791 (O_1791,N_49408,N_49248);
nor UO_1792 (O_1792,N_47996,N_48076);
or UO_1793 (O_1793,N_47716,N_49271);
and UO_1794 (O_1794,N_49948,N_48363);
and UO_1795 (O_1795,N_47731,N_48848);
nor UO_1796 (O_1796,N_49722,N_49397);
and UO_1797 (O_1797,N_47720,N_49716);
and UO_1798 (O_1798,N_49343,N_49077);
nand UO_1799 (O_1799,N_47873,N_47956);
and UO_1800 (O_1800,N_49399,N_47840);
nand UO_1801 (O_1801,N_49742,N_49901);
or UO_1802 (O_1802,N_48846,N_49196);
nand UO_1803 (O_1803,N_49690,N_47623);
nand UO_1804 (O_1804,N_48495,N_48982);
nor UO_1805 (O_1805,N_47983,N_49467);
nor UO_1806 (O_1806,N_48348,N_49754);
nor UO_1807 (O_1807,N_49608,N_49125);
nand UO_1808 (O_1808,N_49247,N_49015);
nand UO_1809 (O_1809,N_49152,N_49150);
or UO_1810 (O_1810,N_48801,N_49149);
and UO_1811 (O_1811,N_49921,N_49047);
xnor UO_1812 (O_1812,N_47563,N_47858);
and UO_1813 (O_1813,N_47555,N_49310);
and UO_1814 (O_1814,N_48779,N_49509);
xor UO_1815 (O_1815,N_49010,N_48000);
and UO_1816 (O_1816,N_48654,N_48347);
nand UO_1817 (O_1817,N_47749,N_48997);
or UO_1818 (O_1818,N_48783,N_49189);
xor UO_1819 (O_1819,N_49103,N_49101);
xor UO_1820 (O_1820,N_49236,N_48125);
nor UO_1821 (O_1821,N_47867,N_49365);
and UO_1822 (O_1822,N_48101,N_48463);
and UO_1823 (O_1823,N_48970,N_49272);
or UO_1824 (O_1824,N_47594,N_47743);
and UO_1825 (O_1825,N_47931,N_49017);
or UO_1826 (O_1826,N_49509,N_49025);
nor UO_1827 (O_1827,N_47946,N_48938);
and UO_1828 (O_1828,N_47822,N_49038);
nand UO_1829 (O_1829,N_49470,N_48622);
xor UO_1830 (O_1830,N_49946,N_48079);
nand UO_1831 (O_1831,N_49588,N_47785);
nor UO_1832 (O_1832,N_48519,N_49820);
xor UO_1833 (O_1833,N_48719,N_47961);
nand UO_1834 (O_1834,N_48531,N_48821);
and UO_1835 (O_1835,N_49245,N_49832);
and UO_1836 (O_1836,N_49451,N_49155);
or UO_1837 (O_1837,N_48643,N_48996);
and UO_1838 (O_1838,N_47752,N_49627);
and UO_1839 (O_1839,N_47757,N_47518);
xor UO_1840 (O_1840,N_49665,N_49133);
nor UO_1841 (O_1841,N_48810,N_48831);
or UO_1842 (O_1842,N_49697,N_48906);
xnor UO_1843 (O_1843,N_48256,N_47527);
nor UO_1844 (O_1844,N_49262,N_48083);
or UO_1845 (O_1845,N_48869,N_48777);
or UO_1846 (O_1846,N_49282,N_48538);
xor UO_1847 (O_1847,N_48994,N_48755);
and UO_1848 (O_1848,N_48886,N_49076);
nor UO_1849 (O_1849,N_48820,N_49399);
nand UO_1850 (O_1850,N_49143,N_48057);
and UO_1851 (O_1851,N_49948,N_48103);
nor UO_1852 (O_1852,N_49402,N_49372);
nor UO_1853 (O_1853,N_47825,N_49148);
nand UO_1854 (O_1854,N_47870,N_48188);
and UO_1855 (O_1855,N_49012,N_48008);
or UO_1856 (O_1856,N_49769,N_48387);
xor UO_1857 (O_1857,N_49141,N_49940);
or UO_1858 (O_1858,N_49667,N_48863);
nor UO_1859 (O_1859,N_48912,N_47767);
nor UO_1860 (O_1860,N_48128,N_47887);
nor UO_1861 (O_1861,N_49603,N_47922);
xnor UO_1862 (O_1862,N_49280,N_49330);
xnor UO_1863 (O_1863,N_49305,N_48705);
or UO_1864 (O_1864,N_49969,N_49736);
and UO_1865 (O_1865,N_48855,N_47659);
nor UO_1866 (O_1866,N_49292,N_49223);
and UO_1867 (O_1867,N_49604,N_48632);
nor UO_1868 (O_1868,N_49616,N_48671);
xnor UO_1869 (O_1869,N_47615,N_49043);
xnor UO_1870 (O_1870,N_49254,N_48111);
and UO_1871 (O_1871,N_49133,N_47541);
nand UO_1872 (O_1872,N_49305,N_49042);
and UO_1873 (O_1873,N_49739,N_49964);
and UO_1874 (O_1874,N_48509,N_48787);
nand UO_1875 (O_1875,N_49785,N_48984);
or UO_1876 (O_1876,N_49827,N_49957);
or UO_1877 (O_1877,N_48492,N_49584);
and UO_1878 (O_1878,N_49442,N_48056);
or UO_1879 (O_1879,N_49936,N_47531);
nand UO_1880 (O_1880,N_48237,N_48265);
nor UO_1881 (O_1881,N_48433,N_49707);
or UO_1882 (O_1882,N_48869,N_48693);
and UO_1883 (O_1883,N_49891,N_49809);
nor UO_1884 (O_1884,N_47795,N_48617);
or UO_1885 (O_1885,N_49664,N_49307);
and UO_1886 (O_1886,N_49886,N_48304);
xnor UO_1887 (O_1887,N_48612,N_47704);
nor UO_1888 (O_1888,N_49416,N_49769);
nand UO_1889 (O_1889,N_49762,N_47505);
nand UO_1890 (O_1890,N_48885,N_49522);
and UO_1891 (O_1891,N_49928,N_49273);
nor UO_1892 (O_1892,N_48192,N_48436);
or UO_1893 (O_1893,N_48420,N_49032);
xnor UO_1894 (O_1894,N_47719,N_48085);
nand UO_1895 (O_1895,N_48182,N_48979);
nand UO_1896 (O_1896,N_48379,N_47978);
and UO_1897 (O_1897,N_48407,N_48669);
nor UO_1898 (O_1898,N_49923,N_48849);
or UO_1899 (O_1899,N_49225,N_48722);
or UO_1900 (O_1900,N_48712,N_48738);
or UO_1901 (O_1901,N_48487,N_49761);
nor UO_1902 (O_1902,N_48744,N_47766);
and UO_1903 (O_1903,N_49904,N_49370);
nor UO_1904 (O_1904,N_47662,N_47814);
nand UO_1905 (O_1905,N_49171,N_48885);
and UO_1906 (O_1906,N_48998,N_48618);
or UO_1907 (O_1907,N_48048,N_49526);
or UO_1908 (O_1908,N_48495,N_47996);
and UO_1909 (O_1909,N_49919,N_49654);
nand UO_1910 (O_1910,N_49332,N_47835);
nor UO_1911 (O_1911,N_49203,N_49743);
nand UO_1912 (O_1912,N_48350,N_47571);
or UO_1913 (O_1913,N_47508,N_48518);
and UO_1914 (O_1914,N_47890,N_47984);
and UO_1915 (O_1915,N_47831,N_49814);
nor UO_1916 (O_1916,N_48244,N_49093);
nand UO_1917 (O_1917,N_49522,N_47849);
nand UO_1918 (O_1918,N_47529,N_47525);
or UO_1919 (O_1919,N_49723,N_49146);
and UO_1920 (O_1920,N_49222,N_49203);
xnor UO_1921 (O_1921,N_49411,N_49046);
or UO_1922 (O_1922,N_49654,N_48237);
nor UO_1923 (O_1923,N_49843,N_47697);
nand UO_1924 (O_1924,N_49489,N_48223);
nor UO_1925 (O_1925,N_49320,N_48780);
nor UO_1926 (O_1926,N_47602,N_49045);
nor UO_1927 (O_1927,N_49703,N_47619);
or UO_1928 (O_1928,N_48315,N_48467);
nor UO_1929 (O_1929,N_48448,N_48631);
xor UO_1930 (O_1930,N_47968,N_49659);
and UO_1931 (O_1931,N_47500,N_49545);
xor UO_1932 (O_1932,N_47938,N_48849);
or UO_1933 (O_1933,N_47944,N_49942);
nor UO_1934 (O_1934,N_49477,N_49809);
nand UO_1935 (O_1935,N_49645,N_49468);
and UO_1936 (O_1936,N_49330,N_49691);
nand UO_1937 (O_1937,N_47564,N_48688);
nor UO_1938 (O_1938,N_49945,N_48681);
nand UO_1939 (O_1939,N_48671,N_48119);
or UO_1940 (O_1940,N_48756,N_49414);
or UO_1941 (O_1941,N_47942,N_47568);
nor UO_1942 (O_1942,N_48828,N_49634);
or UO_1943 (O_1943,N_48190,N_49444);
nand UO_1944 (O_1944,N_49797,N_48186);
nor UO_1945 (O_1945,N_48336,N_48131);
nor UO_1946 (O_1946,N_49170,N_48276);
and UO_1947 (O_1947,N_49639,N_48123);
nor UO_1948 (O_1948,N_48962,N_48627);
nor UO_1949 (O_1949,N_48666,N_48426);
or UO_1950 (O_1950,N_49365,N_48859);
nor UO_1951 (O_1951,N_49163,N_48936);
xnor UO_1952 (O_1952,N_49278,N_47764);
nor UO_1953 (O_1953,N_48377,N_48679);
nand UO_1954 (O_1954,N_48561,N_49760);
nor UO_1955 (O_1955,N_49372,N_49824);
nand UO_1956 (O_1956,N_48431,N_48991);
nand UO_1957 (O_1957,N_48843,N_48426);
nor UO_1958 (O_1958,N_49591,N_48404);
nand UO_1959 (O_1959,N_47630,N_47580);
and UO_1960 (O_1960,N_49410,N_47928);
nand UO_1961 (O_1961,N_49636,N_49263);
and UO_1962 (O_1962,N_48552,N_48106);
nor UO_1963 (O_1963,N_49245,N_47984);
or UO_1964 (O_1964,N_49066,N_47699);
and UO_1965 (O_1965,N_49104,N_49626);
nor UO_1966 (O_1966,N_47985,N_48724);
nand UO_1967 (O_1967,N_49964,N_47928);
nor UO_1968 (O_1968,N_49453,N_49820);
and UO_1969 (O_1969,N_49059,N_49688);
or UO_1970 (O_1970,N_48550,N_47505);
or UO_1971 (O_1971,N_49199,N_48260);
or UO_1972 (O_1972,N_48046,N_48995);
and UO_1973 (O_1973,N_48005,N_49800);
nor UO_1974 (O_1974,N_48402,N_49367);
nor UO_1975 (O_1975,N_47953,N_48536);
nor UO_1976 (O_1976,N_49284,N_49134);
or UO_1977 (O_1977,N_49541,N_49143);
and UO_1978 (O_1978,N_49231,N_48326);
nand UO_1979 (O_1979,N_49331,N_49588);
or UO_1980 (O_1980,N_49916,N_49714);
or UO_1981 (O_1981,N_48977,N_48907);
or UO_1982 (O_1982,N_48564,N_48300);
nor UO_1983 (O_1983,N_49314,N_47683);
and UO_1984 (O_1984,N_47802,N_49697);
nor UO_1985 (O_1985,N_48755,N_47536);
or UO_1986 (O_1986,N_48011,N_49312);
nand UO_1987 (O_1987,N_47510,N_49341);
or UO_1988 (O_1988,N_48708,N_48483);
nand UO_1989 (O_1989,N_47541,N_49390);
or UO_1990 (O_1990,N_48374,N_48322);
or UO_1991 (O_1991,N_49502,N_48845);
or UO_1992 (O_1992,N_48766,N_49768);
nand UO_1993 (O_1993,N_47830,N_48607);
or UO_1994 (O_1994,N_48798,N_48605);
nor UO_1995 (O_1995,N_48987,N_48956);
or UO_1996 (O_1996,N_48435,N_49965);
nor UO_1997 (O_1997,N_47873,N_49528);
nand UO_1998 (O_1998,N_48697,N_47611);
nand UO_1999 (O_1999,N_49011,N_47679);
and UO_2000 (O_2000,N_48237,N_47838);
nor UO_2001 (O_2001,N_48940,N_49619);
and UO_2002 (O_2002,N_47614,N_49316);
xor UO_2003 (O_2003,N_49676,N_48202);
and UO_2004 (O_2004,N_48758,N_48770);
xnor UO_2005 (O_2005,N_48089,N_48611);
or UO_2006 (O_2006,N_47808,N_49927);
xor UO_2007 (O_2007,N_49552,N_48514);
or UO_2008 (O_2008,N_48761,N_49322);
nand UO_2009 (O_2009,N_47673,N_49248);
nand UO_2010 (O_2010,N_48625,N_49667);
nor UO_2011 (O_2011,N_47870,N_48021);
nand UO_2012 (O_2012,N_47587,N_47857);
nand UO_2013 (O_2013,N_48102,N_47846);
or UO_2014 (O_2014,N_48451,N_49293);
nand UO_2015 (O_2015,N_48877,N_49985);
nand UO_2016 (O_2016,N_47997,N_47548);
or UO_2017 (O_2017,N_49012,N_49318);
nand UO_2018 (O_2018,N_49920,N_48024);
or UO_2019 (O_2019,N_47529,N_49231);
xor UO_2020 (O_2020,N_49318,N_47574);
and UO_2021 (O_2021,N_48975,N_49163);
nand UO_2022 (O_2022,N_49655,N_48647);
or UO_2023 (O_2023,N_47738,N_49319);
nor UO_2024 (O_2024,N_49324,N_47903);
xnor UO_2025 (O_2025,N_48651,N_47963);
nor UO_2026 (O_2026,N_47994,N_47988);
nor UO_2027 (O_2027,N_48702,N_49308);
nor UO_2028 (O_2028,N_49000,N_48692);
or UO_2029 (O_2029,N_48002,N_48605);
and UO_2030 (O_2030,N_48341,N_49099);
or UO_2031 (O_2031,N_49937,N_47806);
nor UO_2032 (O_2032,N_49758,N_49493);
nor UO_2033 (O_2033,N_48670,N_48704);
xor UO_2034 (O_2034,N_48396,N_48223);
or UO_2035 (O_2035,N_47937,N_47998);
nand UO_2036 (O_2036,N_47728,N_48686);
or UO_2037 (O_2037,N_48921,N_48484);
nor UO_2038 (O_2038,N_47620,N_49611);
or UO_2039 (O_2039,N_48663,N_49385);
or UO_2040 (O_2040,N_48997,N_49439);
nor UO_2041 (O_2041,N_49861,N_49682);
and UO_2042 (O_2042,N_49504,N_48425);
nand UO_2043 (O_2043,N_48935,N_48838);
nand UO_2044 (O_2044,N_48165,N_47824);
xnor UO_2045 (O_2045,N_47634,N_49463);
and UO_2046 (O_2046,N_48090,N_48417);
nor UO_2047 (O_2047,N_49325,N_47605);
nor UO_2048 (O_2048,N_49625,N_47736);
nor UO_2049 (O_2049,N_49409,N_48456);
or UO_2050 (O_2050,N_49609,N_49892);
and UO_2051 (O_2051,N_48073,N_47995);
nor UO_2052 (O_2052,N_47984,N_48330);
nor UO_2053 (O_2053,N_49246,N_49324);
and UO_2054 (O_2054,N_49046,N_49632);
nand UO_2055 (O_2055,N_49026,N_48265);
or UO_2056 (O_2056,N_48170,N_48488);
nand UO_2057 (O_2057,N_49392,N_47793);
nor UO_2058 (O_2058,N_49625,N_49164);
or UO_2059 (O_2059,N_47642,N_48466);
or UO_2060 (O_2060,N_49321,N_47660);
nor UO_2061 (O_2061,N_49356,N_49340);
xnor UO_2062 (O_2062,N_48872,N_47797);
nand UO_2063 (O_2063,N_47856,N_49282);
and UO_2064 (O_2064,N_49791,N_49560);
nor UO_2065 (O_2065,N_49411,N_48263);
and UO_2066 (O_2066,N_49235,N_48024);
xor UO_2067 (O_2067,N_47677,N_49912);
nor UO_2068 (O_2068,N_49781,N_48030);
nand UO_2069 (O_2069,N_49227,N_49906);
or UO_2070 (O_2070,N_49655,N_49980);
nand UO_2071 (O_2071,N_48077,N_49201);
nor UO_2072 (O_2072,N_49342,N_48047);
nor UO_2073 (O_2073,N_49118,N_49254);
or UO_2074 (O_2074,N_49892,N_49416);
nor UO_2075 (O_2075,N_48939,N_48821);
nand UO_2076 (O_2076,N_49991,N_47768);
nand UO_2077 (O_2077,N_47899,N_48066);
and UO_2078 (O_2078,N_49604,N_48682);
and UO_2079 (O_2079,N_48945,N_48314);
nor UO_2080 (O_2080,N_48812,N_47977);
or UO_2081 (O_2081,N_49648,N_48763);
and UO_2082 (O_2082,N_49130,N_49597);
and UO_2083 (O_2083,N_47786,N_48278);
and UO_2084 (O_2084,N_49789,N_47956);
nand UO_2085 (O_2085,N_47929,N_47769);
and UO_2086 (O_2086,N_49593,N_48887);
nand UO_2087 (O_2087,N_47829,N_47524);
nand UO_2088 (O_2088,N_48226,N_49341);
and UO_2089 (O_2089,N_47652,N_48385);
and UO_2090 (O_2090,N_48964,N_49626);
nor UO_2091 (O_2091,N_47570,N_47837);
nor UO_2092 (O_2092,N_48158,N_49554);
or UO_2093 (O_2093,N_49003,N_48750);
and UO_2094 (O_2094,N_48715,N_49290);
nor UO_2095 (O_2095,N_47890,N_49330);
and UO_2096 (O_2096,N_48590,N_48432);
and UO_2097 (O_2097,N_49747,N_47540);
nand UO_2098 (O_2098,N_48462,N_49935);
xnor UO_2099 (O_2099,N_48115,N_48890);
nand UO_2100 (O_2100,N_49698,N_49239);
nand UO_2101 (O_2101,N_48215,N_48424);
nor UO_2102 (O_2102,N_47927,N_48717);
and UO_2103 (O_2103,N_49722,N_48959);
nor UO_2104 (O_2104,N_49368,N_49417);
and UO_2105 (O_2105,N_48754,N_49706);
nand UO_2106 (O_2106,N_48553,N_49486);
or UO_2107 (O_2107,N_48606,N_48137);
and UO_2108 (O_2108,N_48148,N_49557);
nand UO_2109 (O_2109,N_49675,N_47917);
or UO_2110 (O_2110,N_49663,N_49940);
nor UO_2111 (O_2111,N_49082,N_48834);
and UO_2112 (O_2112,N_47837,N_48621);
nand UO_2113 (O_2113,N_49561,N_49557);
or UO_2114 (O_2114,N_47925,N_49890);
or UO_2115 (O_2115,N_49139,N_47974);
nor UO_2116 (O_2116,N_48186,N_49084);
or UO_2117 (O_2117,N_48122,N_48446);
and UO_2118 (O_2118,N_48990,N_48104);
xor UO_2119 (O_2119,N_49014,N_49285);
nor UO_2120 (O_2120,N_47796,N_47746);
and UO_2121 (O_2121,N_48504,N_48038);
or UO_2122 (O_2122,N_49011,N_48062);
nand UO_2123 (O_2123,N_47988,N_49820);
or UO_2124 (O_2124,N_49996,N_48288);
or UO_2125 (O_2125,N_48217,N_48358);
xor UO_2126 (O_2126,N_48665,N_48523);
nor UO_2127 (O_2127,N_48943,N_48039);
and UO_2128 (O_2128,N_47663,N_49534);
nor UO_2129 (O_2129,N_48859,N_49231);
and UO_2130 (O_2130,N_48355,N_47858);
and UO_2131 (O_2131,N_49841,N_49307);
and UO_2132 (O_2132,N_49732,N_47609);
nor UO_2133 (O_2133,N_48238,N_47698);
nor UO_2134 (O_2134,N_48298,N_49019);
and UO_2135 (O_2135,N_47731,N_49687);
and UO_2136 (O_2136,N_48755,N_47746);
nor UO_2137 (O_2137,N_47688,N_47506);
nand UO_2138 (O_2138,N_49301,N_48207);
nand UO_2139 (O_2139,N_49330,N_48802);
or UO_2140 (O_2140,N_48297,N_48138);
nor UO_2141 (O_2141,N_48656,N_47866);
and UO_2142 (O_2142,N_49706,N_47951);
nor UO_2143 (O_2143,N_49549,N_48531);
nand UO_2144 (O_2144,N_48483,N_48527);
nor UO_2145 (O_2145,N_48786,N_49028);
nand UO_2146 (O_2146,N_48982,N_47556);
and UO_2147 (O_2147,N_48951,N_47633);
and UO_2148 (O_2148,N_48585,N_49978);
or UO_2149 (O_2149,N_48069,N_49663);
or UO_2150 (O_2150,N_49450,N_49056);
nand UO_2151 (O_2151,N_49636,N_47883);
nand UO_2152 (O_2152,N_48767,N_48707);
and UO_2153 (O_2153,N_48175,N_48359);
nand UO_2154 (O_2154,N_49687,N_49312);
nor UO_2155 (O_2155,N_48089,N_47682);
or UO_2156 (O_2156,N_47833,N_47543);
and UO_2157 (O_2157,N_48689,N_49103);
xnor UO_2158 (O_2158,N_49676,N_49882);
nor UO_2159 (O_2159,N_48147,N_47743);
and UO_2160 (O_2160,N_48158,N_47654);
or UO_2161 (O_2161,N_49820,N_48228);
and UO_2162 (O_2162,N_48538,N_47505);
or UO_2163 (O_2163,N_49519,N_48129);
and UO_2164 (O_2164,N_49627,N_47589);
or UO_2165 (O_2165,N_48631,N_48418);
or UO_2166 (O_2166,N_49244,N_47934);
and UO_2167 (O_2167,N_49067,N_47537);
xnor UO_2168 (O_2168,N_48952,N_48424);
or UO_2169 (O_2169,N_48560,N_47931);
and UO_2170 (O_2170,N_48767,N_49389);
nor UO_2171 (O_2171,N_48786,N_47768);
nor UO_2172 (O_2172,N_48892,N_48658);
nor UO_2173 (O_2173,N_47705,N_49055);
nand UO_2174 (O_2174,N_47968,N_48678);
nand UO_2175 (O_2175,N_48326,N_48305);
nand UO_2176 (O_2176,N_49274,N_48848);
nor UO_2177 (O_2177,N_49873,N_48449);
nor UO_2178 (O_2178,N_47733,N_49342);
nand UO_2179 (O_2179,N_47715,N_49806);
nor UO_2180 (O_2180,N_49225,N_48966);
xor UO_2181 (O_2181,N_49618,N_47991);
nor UO_2182 (O_2182,N_48539,N_48203);
and UO_2183 (O_2183,N_49568,N_48958);
nor UO_2184 (O_2184,N_48976,N_49072);
or UO_2185 (O_2185,N_48591,N_49927);
nand UO_2186 (O_2186,N_49229,N_49255);
nor UO_2187 (O_2187,N_48260,N_48111);
nor UO_2188 (O_2188,N_47560,N_49657);
nor UO_2189 (O_2189,N_47863,N_47849);
nand UO_2190 (O_2190,N_49674,N_48746);
nor UO_2191 (O_2191,N_49041,N_49462);
nor UO_2192 (O_2192,N_48183,N_48690);
nor UO_2193 (O_2193,N_48158,N_48292);
xnor UO_2194 (O_2194,N_49023,N_48253);
and UO_2195 (O_2195,N_48259,N_47948);
xor UO_2196 (O_2196,N_47706,N_49836);
or UO_2197 (O_2197,N_48510,N_47951);
or UO_2198 (O_2198,N_49789,N_48395);
nand UO_2199 (O_2199,N_48685,N_49209);
or UO_2200 (O_2200,N_48949,N_48108);
xnor UO_2201 (O_2201,N_48326,N_48965);
nor UO_2202 (O_2202,N_48020,N_49010);
or UO_2203 (O_2203,N_49366,N_48909);
nor UO_2204 (O_2204,N_49234,N_49575);
xnor UO_2205 (O_2205,N_49708,N_48484);
and UO_2206 (O_2206,N_48461,N_48270);
nand UO_2207 (O_2207,N_48572,N_47937);
or UO_2208 (O_2208,N_48961,N_48667);
or UO_2209 (O_2209,N_49813,N_47633);
or UO_2210 (O_2210,N_47847,N_49600);
xnor UO_2211 (O_2211,N_47509,N_48631);
xnor UO_2212 (O_2212,N_49298,N_49977);
or UO_2213 (O_2213,N_49125,N_48564);
or UO_2214 (O_2214,N_49367,N_49497);
nor UO_2215 (O_2215,N_48807,N_48258);
and UO_2216 (O_2216,N_47792,N_48869);
or UO_2217 (O_2217,N_48543,N_49710);
nand UO_2218 (O_2218,N_49737,N_48630);
or UO_2219 (O_2219,N_48890,N_49582);
nand UO_2220 (O_2220,N_48304,N_48734);
or UO_2221 (O_2221,N_49070,N_48631);
nand UO_2222 (O_2222,N_47850,N_49794);
or UO_2223 (O_2223,N_48954,N_49129);
nand UO_2224 (O_2224,N_49238,N_49830);
nand UO_2225 (O_2225,N_48590,N_47728);
nand UO_2226 (O_2226,N_49844,N_49597);
and UO_2227 (O_2227,N_49435,N_48911);
and UO_2228 (O_2228,N_48374,N_47803);
and UO_2229 (O_2229,N_48479,N_48775);
and UO_2230 (O_2230,N_49348,N_48400);
nand UO_2231 (O_2231,N_48701,N_48506);
xor UO_2232 (O_2232,N_48348,N_49889);
xnor UO_2233 (O_2233,N_49234,N_48383);
nor UO_2234 (O_2234,N_49275,N_49186);
nand UO_2235 (O_2235,N_48313,N_47520);
or UO_2236 (O_2236,N_49473,N_48463);
xor UO_2237 (O_2237,N_48268,N_49065);
nor UO_2238 (O_2238,N_48995,N_47971);
and UO_2239 (O_2239,N_48802,N_47767);
or UO_2240 (O_2240,N_49390,N_49626);
and UO_2241 (O_2241,N_49287,N_48553);
nor UO_2242 (O_2242,N_48803,N_47797);
xnor UO_2243 (O_2243,N_49541,N_48110);
or UO_2244 (O_2244,N_49217,N_49889);
xnor UO_2245 (O_2245,N_48732,N_49590);
nand UO_2246 (O_2246,N_48893,N_49049);
and UO_2247 (O_2247,N_49328,N_48280);
nor UO_2248 (O_2248,N_48441,N_49308);
nor UO_2249 (O_2249,N_48388,N_48029);
and UO_2250 (O_2250,N_47766,N_47681);
xor UO_2251 (O_2251,N_48520,N_48271);
nand UO_2252 (O_2252,N_48924,N_47577);
nand UO_2253 (O_2253,N_47639,N_48175);
or UO_2254 (O_2254,N_49272,N_49324);
nor UO_2255 (O_2255,N_49375,N_49822);
nand UO_2256 (O_2256,N_49630,N_49004);
and UO_2257 (O_2257,N_49458,N_48262);
or UO_2258 (O_2258,N_49925,N_49858);
or UO_2259 (O_2259,N_48639,N_48729);
nand UO_2260 (O_2260,N_49139,N_48714);
nor UO_2261 (O_2261,N_49909,N_47987);
nand UO_2262 (O_2262,N_48669,N_49120);
or UO_2263 (O_2263,N_48069,N_48974);
nor UO_2264 (O_2264,N_48927,N_49978);
or UO_2265 (O_2265,N_47794,N_48767);
xnor UO_2266 (O_2266,N_47540,N_49692);
and UO_2267 (O_2267,N_49709,N_49394);
nor UO_2268 (O_2268,N_49841,N_49687);
and UO_2269 (O_2269,N_49638,N_48629);
nor UO_2270 (O_2270,N_48797,N_49079);
nand UO_2271 (O_2271,N_48369,N_48865);
nor UO_2272 (O_2272,N_49863,N_48647);
and UO_2273 (O_2273,N_49539,N_47789);
nor UO_2274 (O_2274,N_48447,N_48752);
nand UO_2275 (O_2275,N_47891,N_48821);
nand UO_2276 (O_2276,N_48349,N_47831);
xnor UO_2277 (O_2277,N_48643,N_48151);
or UO_2278 (O_2278,N_48449,N_49636);
xor UO_2279 (O_2279,N_48813,N_48632);
and UO_2280 (O_2280,N_47871,N_49636);
nand UO_2281 (O_2281,N_48385,N_49993);
and UO_2282 (O_2282,N_47611,N_48190);
xor UO_2283 (O_2283,N_48981,N_48013);
nand UO_2284 (O_2284,N_48895,N_48836);
or UO_2285 (O_2285,N_49304,N_48725);
and UO_2286 (O_2286,N_48282,N_48886);
nor UO_2287 (O_2287,N_48426,N_48210);
xnor UO_2288 (O_2288,N_49057,N_49016);
or UO_2289 (O_2289,N_48585,N_48687);
and UO_2290 (O_2290,N_48543,N_48931);
and UO_2291 (O_2291,N_48298,N_47988);
or UO_2292 (O_2292,N_48346,N_49860);
or UO_2293 (O_2293,N_48663,N_47538);
nand UO_2294 (O_2294,N_47545,N_49782);
and UO_2295 (O_2295,N_48191,N_49435);
and UO_2296 (O_2296,N_49406,N_48050);
nor UO_2297 (O_2297,N_48064,N_49374);
and UO_2298 (O_2298,N_48574,N_48697);
and UO_2299 (O_2299,N_48447,N_48432);
and UO_2300 (O_2300,N_49576,N_49891);
nor UO_2301 (O_2301,N_47925,N_49341);
nor UO_2302 (O_2302,N_49947,N_47608);
xnor UO_2303 (O_2303,N_48488,N_47826);
nand UO_2304 (O_2304,N_48642,N_49547);
nand UO_2305 (O_2305,N_49324,N_48807);
and UO_2306 (O_2306,N_47571,N_49481);
nand UO_2307 (O_2307,N_48063,N_47999);
nand UO_2308 (O_2308,N_48922,N_47874);
nor UO_2309 (O_2309,N_48559,N_49098);
nor UO_2310 (O_2310,N_47536,N_47708);
xor UO_2311 (O_2311,N_48391,N_48056);
and UO_2312 (O_2312,N_48785,N_48916);
nand UO_2313 (O_2313,N_48943,N_47605);
or UO_2314 (O_2314,N_48010,N_47539);
nand UO_2315 (O_2315,N_49434,N_48418);
nand UO_2316 (O_2316,N_48630,N_49035);
and UO_2317 (O_2317,N_49820,N_49850);
nor UO_2318 (O_2318,N_49221,N_47820);
nor UO_2319 (O_2319,N_48917,N_48195);
xor UO_2320 (O_2320,N_49984,N_49329);
nand UO_2321 (O_2321,N_48471,N_47740);
nand UO_2322 (O_2322,N_48808,N_47839);
and UO_2323 (O_2323,N_48458,N_47772);
and UO_2324 (O_2324,N_48587,N_49511);
nor UO_2325 (O_2325,N_49556,N_49077);
nor UO_2326 (O_2326,N_48334,N_49946);
nand UO_2327 (O_2327,N_48311,N_47720);
and UO_2328 (O_2328,N_48053,N_48536);
or UO_2329 (O_2329,N_48653,N_49855);
nor UO_2330 (O_2330,N_47839,N_49168);
or UO_2331 (O_2331,N_49841,N_49848);
and UO_2332 (O_2332,N_49482,N_48996);
nor UO_2333 (O_2333,N_48062,N_48294);
and UO_2334 (O_2334,N_48728,N_47833);
or UO_2335 (O_2335,N_49813,N_49485);
nor UO_2336 (O_2336,N_47782,N_48485);
or UO_2337 (O_2337,N_47825,N_49446);
nand UO_2338 (O_2338,N_48491,N_49356);
and UO_2339 (O_2339,N_49381,N_48914);
or UO_2340 (O_2340,N_48924,N_49580);
nor UO_2341 (O_2341,N_47631,N_49788);
nor UO_2342 (O_2342,N_48160,N_49848);
nor UO_2343 (O_2343,N_49288,N_47783);
or UO_2344 (O_2344,N_49509,N_48871);
nand UO_2345 (O_2345,N_48732,N_47779);
or UO_2346 (O_2346,N_47866,N_48347);
nor UO_2347 (O_2347,N_49132,N_47882);
and UO_2348 (O_2348,N_48296,N_48597);
or UO_2349 (O_2349,N_49144,N_48601);
or UO_2350 (O_2350,N_49926,N_48412);
xor UO_2351 (O_2351,N_47596,N_49918);
nor UO_2352 (O_2352,N_48179,N_49507);
nand UO_2353 (O_2353,N_48874,N_49326);
and UO_2354 (O_2354,N_49922,N_48140);
nand UO_2355 (O_2355,N_49771,N_47850);
xor UO_2356 (O_2356,N_48292,N_48987);
or UO_2357 (O_2357,N_48000,N_48367);
nor UO_2358 (O_2358,N_49370,N_47618);
nand UO_2359 (O_2359,N_47663,N_49880);
or UO_2360 (O_2360,N_48255,N_47697);
or UO_2361 (O_2361,N_49161,N_48761);
and UO_2362 (O_2362,N_49262,N_47521);
and UO_2363 (O_2363,N_47740,N_48347);
and UO_2364 (O_2364,N_47519,N_48050);
nor UO_2365 (O_2365,N_49471,N_48927);
or UO_2366 (O_2366,N_49785,N_48693);
nand UO_2367 (O_2367,N_49405,N_48604);
or UO_2368 (O_2368,N_48088,N_48807);
and UO_2369 (O_2369,N_49955,N_48714);
and UO_2370 (O_2370,N_49617,N_48667);
or UO_2371 (O_2371,N_47927,N_48116);
nor UO_2372 (O_2372,N_49081,N_49852);
nand UO_2373 (O_2373,N_48871,N_49940);
nand UO_2374 (O_2374,N_48913,N_49173);
and UO_2375 (O_2375,N_47701,N_49446);
and UO_2376 (O_2376,N_48958,N_49348);
or UO_2377 (O_2377,N_49320,N_47603);
nand UO_2378 (O_2378,N_49325,N_48085);
nand UO_2379 (O_2379,N_48647,N_49395);
nand UO_2380 (O_2380,N_47675,N_48990);
nand UO_2381 (O_2381,N_49668,N_48901);
nand UO_2382 (O_2382,N_48763,N_49145);
or UO_2383 (O_2383,N_48495,N_48152);
nor UO_2384 (O_2384,N_47926,N_49425);
xnor UO_2385 (O_2385,N_49995,N_48703);
nand UO_2386 (O_2386,N_48793,N_48110);
nand UO_2387 (O_2387,N_48346,N_48978);
nand UO_2388 (O_2388,N_48775,N_49380);
nand UO_2389 (O_2389,N_49809,N_48577);
or UO_2390 (O_2390,N_49346,N_49956);
nand UO_2391 (O_2391,N_48950,N_49511);
nor UO_2392 (O_2392,N_49816,N_47993);
nand UO_2393 (O_2393,N_47569,N_49493);
nor UO_2394 (O_2394,N_49679,N_48383);
nor UO_2395 (O_2395,N_47977,N_49843);
nor UO_2396 (O_2396,N_48863,N_48088);
nand UO_2397 (O_2397,N_48868,N_49028);
or UO_2398 (O_2398,N_48855,N_49730);
and UO_2399 (O_2399,N_49566,N_47913);
and UO_2400 (O_2400,N_49357,N_49180);
and UO_2401 (O_2401,N_48049,N_48564);
nor UO_2402 (O_2402,N_49894,N_49759);
or UO_2403 (O_2403,N_48969,N_49310);
nor UO_2404 (O_2404,N_49428,N_48559);
nand UO_2405 (O_2405,N_47584,N_48579);
nand UO_2406 (O_2406,N_48440,N_48992);
or UO_2407 (O_2407,N_49427,N_48178);
xnor UO_2408 (O_2408,N_47554,N_48262);
and UO_2409 (O_2409,N_49590,N_48145);
nor UO_2410 (O_2410,N_47675,N_47696);
nand UO_2411 (O_2411,N_49997,N_49931);
nand UO_2412 (O_2412,N_49893,N_48474);
nor UO_2413 (O_2413,N_48990,N_48964);
or UO_2414 (O_2414,N_48593,N_48624);
nand UO_2415 (O_2415,N_48101,N_48362);
nand UO_2416 (O_2416,N_47623,N_47885);
nand UO_2417 (O_2417,N_48510,N_49586);
nor UO_2418 (O_2418,N_48179,N_47721);
or UO_2419 (O_2419,N_48701,N_49586);
or UO_2420 (O_2420,N_48643,N_48462);
nand UO_2421 (O_2421,N_49394,N_49405);
and UO_2422 (O_2422,N_48612,N_48444);
xnor UO_2423 (O_2423,N_49227,N_47800);
and UO_2424 (O_2424,N_48226,N_49637);
or UO_2425 (O_2425,N_48262,N_47862);
and UO_2426 (O_2426,N_48883,N_49051);
and UO_2427 (O_2427,N_48050,N_49137);
nor UO_2428 (O_2428,N_48977,N_49508);
nand UO_2429 (O_2429,N_48066,N_48121);
and UO_2430 (O_2430,N_48118,N_48381);
xor UO_2431 (O_2431,N_48291,N_49636);
nor UO_2432 (O_2432,N_49222,N_49618);
nor UO_2433 (O_2433,N_48506,N_49071);
or UO_2434 (O_2434,N_47829,N_49755);
nor UO_2435 (O_2435,N_49852,N_48871);
and UO_2436 (O_2436,N_48680,N_48655);
nor UO_2437 (O_2437,N_48574,N_48204);
and UO_2438 (O_2438,N_49784,N_49341);
nand UO_2439 (O_2439,N_47892,N_48453);
nand UO_2440 (O_2440,N_48302,N_49991);
and UO_2441 (O_2441,N_47784,N_47540);
nor UO_2442 (O_2442,N_49189,N_48027);
nor UO_2443 (O_2443,N_47781,N_47872);
nor UO_2444 (O_2444,N_49463,N_49429);
or UO_2445 (O_2445,N_49514,N_48890);
or UO_2446 (O_2446,N_48018,N_49067);
nand UO_2447 (O_2447,N_49722,N_48382);
nor UO_2448 (O_2448,N_49388,N_49568);
or UO_2449 (O_2449,N_47589,N_48557);
nor UO_2450 (O_2450,N_49578,N_47841);
or UO_2451 (O_2451,N_47940,N_49772);
xnor UO_2452 (O_2452,N_49705,N_48719);
nand UO_2453 (O_2453,N_48698,N_49283);
nor UO_2454 (O_2454,N_49646,N_48122);
or UO_2455 (O_2455,N_49799,N_49432);
nor UO_2456 (O_2456,N_49737,N_48214);
nand UO_2457 (O_2457,N_47563,N_49121);
or UO_2458 (O_2458,N_49126,N_48202);
nand UO_2459 (O_2459,N_47793,N_49821);
or UO_2460 (O_2460,N_48242,N_48404);
nand UO_2461 (O_2461,N_49049,N_48942);
nand UO_2462 (O_2462,N_49335,N_49187);
and UO_2463 (O_2463,N_49803,N_47566);
nor UO_2464 (O_2464,N_47933,N_49087);
or UO_2465 (O_2465,N_48825,N_48913);
or UO_2466 (O_2466,N_49046,N_49129);
xnor UO_2467 (O_2467,N_48128,N_47911);
or UO_2468 (O_2468,N_49647,N_47872);
xor UO_2469 (O_2469,N_48534,N_49203);
nand UO_2470 (O_2470,N_49445,N_47859);
or UO_2471 (O_2471,N_48796,N_48239);
nand UO_2472 (O_2472,N_47919,N_49427);
and UO_2473 (O_2473,N_47714,N_48968);
nor UO_2474 (O_2474,N_48193,N_47594);
nor UO_2475 (O_2475,N_49649,N_49122);
nor UO_2476 (O_2476,N_47610,N_49470);
nand UO_2477 (O_2477,N_48529,N_48108);
nor UO_2478 (O_2478,N_49790,N_49789);
xor UO_2479 (O_2479,N_48077,N_49512);
nand UO_2480 (O_2480,N_48925,N_48577);
nor UO_2481 (O_2481,N_47962,N_49338);
nor UO_2482 (O_2482,N_48916,N_49062);
nor UO_2483 (O_2483,N_48142,N_49790);
or UO_2484 (O_2484,N_48154,N_48973);
nand UO_2485 (O_2485,N_49479,N_48246);
nor UO_2486 (O_2486,N_49799,N_49999);
nand UO_2487 (O_2487,N_47713,N_49567);
nand UO_2488 (O_2488,N_47585,N_48415);
or UO_2489 (O_2489,N_48138,N_49829);
or UO_2490 (O_2490,N_48227,N_48511);
and UO_2491 (O_2491,N_49817,N_48671);
xor UO_2492 (O_2492,N_47673,N_49856);
xnor UO_2493 (O_2493,N_47700,N_47846);
nand UO_2494 (O_2494,N_47578,N_48103);
nand UO_2495 (O_2495,N_49628,N_49847);
xnor UO_2496 (O_2496,N_47693,N_48046);
xor UO_2497 (O_2497,N_47868,N_49695);
nor UO_2498 (O_2498,N_48537,N_49004);
or UO_2499 (O_2499,N_47503,N_48537);
and UO_2500 (O_2500,N_49321,N_49386);
or UO_2501 (O_2501,N_49792,N_48858);
and UO_2502 (O_2502,N_48736,N_49457);
or UO_2503 (O_2503,N_47665,N_48106);
nor UO_2504 (O_2504,N_49532,N_49315);
nor UO_2505 (O_2505,N_48044,N_48395);
and UO_2506 (O_2506,N_49913,N_49396);
nand UO_2507 (O_2507,N_49784,N_49670);
or UO_2508 (O_2508,N_49885,N_47616);
and UO_2509 (O_2509,N_49224,N_47717);
and UO_2510 (O_2510,N_48083,N_49567);
and UO_2511 (O_2511,N_47747,N_49658);
or UO_2512 (O_2512,N_47584,N_48301);
nand UO_2513 (O_2513,N_48817,N_48479);
or UO_2514 (O_2514,N_48327,N_48843);
or UO_2515 (O_2515,N_49385,N_48453);
or UO_2516 (O_2516,N_49781,N_47932);
or UO_2517 (O_2517,N_48781,N_49822);
nor UO_2518 (O_2518,N_47829,N_49398);
and UO_2519 (O_2519,N_49281,N_48722);
nor UO_2520 (O_2520,N_48668,N_49980);
and UO_2521 (O_2521,N_49728,N_49207);
xor UO_2522 (O_2522,N_47915,N_49685);
nor UO_2523 (O_2523,N_49890,N_47575);
nor UO_2524 (O_2524,N_49564,N_47871);
nor UO_2525 (O_2525,N_48224,N_48560);
nand UO_2526 (O_2526,N_48373,N_49534);
nor UO_2527 (O_2527,N_49127,N_47565);
and UO_2528 (O_2528,N_49982,N_48117);
and UO_2529 (O_2529,N_48435,N_48815);
nand UO_2530 (O_2530,N_48331,N_49298);
nand UO_2531 (O_2531,N_48764,N_49606);
nand UO_2532 (O_2532,N_49659,N_47777);
and UO_2533 (O_2533,N_49228,N_48648);
xnor UO_2534 (O_2534,N_47731,N_47895);
nand UO_2535 (O_2535,N_47823,N_49825);
or UO_2536 (O_2536,N_48822,N_49604);
nor UO_2537 (O_2537,N_47660,N_49922);
or UO_2538 (O_2538,N_49913,N_49176);
nand UO_2539 (O_2539,N_47953,N_49004);
nor UO_2540 (O_2540,N_48450,N_49661);
or UO_2541 (O_2541,N_48533,N_49789);
nor UO_2542 (O_2542,N_47558,N_49160);
nor UO_2543 (O_2543,N_47886,N_49352);
nand UO_2544 (O_2544,N_49593,N_48415);
or UO_2545 (O_2545,N_49577,N_47908);
and UO_2546 (O_2546,N_48452,N_47564);
nor UO_2547 (O_2547,N_48655,N_48532);
nor UO_2548 (O_2548,N_49144,N_49118);
and UO_2549 (O_2549,N_49655,N_47672);
xnor UO_2550 (O_2550,N_48444,N_48047);
and UO_2551 (O_2551,N_48484,N_49726);
nand UO_2552 (O_2552,N_49270,N_49441);
nor UO_2553 (O_2553,N_47972,N_47848);
and UO_2554 (O_2554,N_48621,N_47737);
nor UO_2555 (O_2555,N_48436,N_49283);
xnor UO_2556 (O_2556,N_48723,N_49592);
xor UO_2557 (O_2557,N_49252,N_48183);
and UO_2558 (O_2558,N_48782,N_49852);
and UO_2559 (O_2559,N_48306,N_48624);
or UO_2560 (O_2560,N_49581,N_49972);
nand UO_2561 (O_2561,N_47607,N_49838);
and UO_2562 (O_2562,N_47994,N_48478);
nand UO_2563 (O_2563,N_47598,N_49052);
nand UO_2564 (O_2564,N_47902,N_48145);
nand UO_2565 (O_2565,N_48297,N_48547);
or UO_2566 (O_2566,N_49018,N_48527);
or UO_2567 (O_2567,N_49870,N_49515);
nand UO_2568 (O_2568,N_47748,N_47992);
or UO_2569 (O_2569,N_47663,N_48758);
nor UO_2570 (O_2570,N_48989,N_47880);
nor UO_2571 (O_2571,N_48516,N_49022);
or UO_2572 (O_2572,N_49296,N_47887);
and UO_2573 (O_2573,N_47934,N_49394);
nand UO_2574 (O_2574,N_48626,N_49807);
and UO_2575 (O_2575,N_48350,N_49914);
nor UO_2576 (O_2576,N_47733,N_49428);
or UO_2577 (O_2577,N_49534,N_49877);
and UO_2578 (O_2578,N_49805,N_48281);
and UO_2579 (O_2579,N_48863,N_49530);
or UO_2580 (O_2580,N_48397,N_49336);
nand UO_2581 (O_2581,N_49631,N_49056);
nand UO_2582 (O_2582,N_47959,N_49730);
nand UO_2583 (O_2583,N_49266,N_48326);
and UO_2584 (O_2584,N_48685,N_47820);
nand UO_2585 (O_2585,N_49143,N_48044);
and UO_2586 (O_2586,N_49583,N_48391);
xnor UO_2587 (O_2587,N_48113,N_49381);
nor UO_2588 (O_2588,N_49026,N_48643);
nor UO_2589 (O_2589,N_49899,N_48270);
nor UO_2590 (O_2590,N_49165,N_47594);
or UO_2591 (O_2591,N_49429,N_48634);
and UO_2592 (O_2592,N_49794,N_49955);
nand UO_2593 (O_2593,N_49946,N_47885);
or UO_2594 (O_2594,N_47925,N_49078);
nor UO_2595 (O_2595,N_47639,N_48954);
or UO_2596 (O_2596,N_49697,N_48970);
nor UO_2597 (O_2597,N_49457,N_48556);
or UO_2598 (O_2598,N_49177,N_47642);
nand UO_2599 (O_2599,N_49356,N_49508);
and UO_2600 (O_2600,N_48263,N_47872);
nor UO_2601 (O_2601,N_49121,N_49060);
xor UO_2602 (O_2602,N_48361,N_48348);
nand UO_2603 (O_2603,N_47537,N_48603);
xnor UO_2604 (O_2604,N_49885,N_47918);
nor UO_2605 (O_2605,N_49351,N_48392);
xor UO_2606 (O_2606,N_49228,N_49374);
nand UO_2607 (O_2607,N_48298,N_49466);
and UO_2608 (O_2608,N_48489,N_48680);
xnor UO_2609 (O_2609,N_48823,N_49569);
or UO_2610 (O_2610,N_48414,N_49431);
and UO_2611 (O_2611,N_49676,N_49085);
and UO_2612 (O_2612,N_49698,N_49236);
or UO_2613 (O_2613,N_49236,N_49751);
nor UO_2614 (O_2614,N_48279,N_49095);
nor UO_2615 (O_2615,N_49378,N_49902);
or UO_2616 (O_2616,N_47929,N_49049);
nand UO_2617 (O_2617,N_47529,N_48646);
nand UO_2618 (O_2618,N_49356,N_48878);
or UO_2619 (O_2619,N_48402,N_49373);
nand UO_2620 (O_2620,N_49041,N_49047);
and UO_2621 (O_2621,N_47973,N_48970);
xnor UO_2622 (O_2622,N_49113,N_49313);
nand UO_2623 (O_2623,N_49110,N_47856);
and UO_2624 (O_2624,N_48571,N_48303);
and UO_2625 (O_2625,N_49715,N_48202);
nand UO_2626 (O_2626,N_49784,N_47664);
xor UO_2627 (O_2627,N_48116,N_48381);
or UO_2628 (O_2628,N_48153,N_47717);
nand UO_2629 (O_2629,N_48483,N_49696);
nand UO_2630 (O_2630,N_47708,N_49172);
nand UO_2631 (O_2631,N_49089,N_49815);
nor UO_2632 (O_2632,N_49778,N_49780);
and UO_2633 (O_2633,N_48315,N_49146);
and UO_2634 (O_2634,N_48780,N_49232);
nor UO_2635 (O_2635,N_49585,N_48157);
xnor UO_2636 (O_2636,N_47673,N_47691);
and UO_2637 (O_2637,N_48397,N_48496);
nor UO_2638 (O_2638,N_48723,N_49106);
xnor UO_2639 (O_2639,N_47508,N_49701);
and UO_2640 (O_2640,N_47894,N_48212);
and UO_2641 (O_2641,N_48461,N_48719);
nor UO_2642 (O_2642,N_49351,N_48636);
nand UO_2643 (O_2643,N_49403,N_49259);
and UO_2644 (O_2644,N_49284,N_48116);
or UO_2645 (O_2645,N_47961,N_49384);
and UO_2646 (O_2646,N_49639,N_49444);
or UO_2647 (O_2647,N_49638,N_48456);
xnor UO_2648 (O_2648,N_49992,N_49053);
nor UO_2649 (O_2649,N_49727,N_49001);
and UO_2650 (O_2650,N_48951,N_48601);
and UO_2651 (O_2651,N_49722,N_49914);
nor UO_2652 (O_2652,N_48517,N_48389);
or UO_2653 (O_2653,N_49212,N_48003);
and UO_2654 (O_2654,N_48575,N_49026);
nand UO_2655 (O_2655,N_48643,N_47733);
nand UO_2656 (O_2656,N_48395,N_47648);
nor UO_2657 (O_2657,N_49627,N_49072);
and UO_2658 (O_2658,N_49307,N_49581);
nand UO_2659 (O_2659,N_48614,N_49699);
nor UO_2660 (O_2660,N_47872,N_49653);
nand UO_2661 (O_2661,N_48735,N_48916);
nor UO_2662 (O_2662,N_49519,N_48762);
nor UO_2663 (O_2663,N_48546,N_48581);
xor UO_2664 (O_2664,N_49136,N_48266);
nor UO_2665 (O_2665,N_47656,N_47647);
nor UO_2666 (O_2666,N_47946,N_47672);
nor UO_2667 (O_2667,N_48935,N_48975);
nand UO_2668 (O_2668,N_48277,N_48046);
xor UO_2669 (O_2669,N_47597,N_47783);
nor UO_2670 (O_2670,N_48157,N_48964);
or UO_2671 (O_2671,N_47684,N_47708);
or UO_2672 (O_2672,N_48411,N_48607);
nor UO_2673 (O_2673,N_48048,N_47993);
or UO_2674 (O_2674,N_47840,N_49075);
nor UO_2675 (O_2675,N_49614,N_48612);
xor UO_2676 (O_2676,N_48889,N_49620);
and UO_2677 (O_2677,N_48982,N_48523);
nand UO_2678 (O_2678,N_49020,N_48901);
and UO_2679 (O_2679,N_48556,N_48701);
nor UO_2680 (O_2680,N_47655,N_49412);
xnor UO_2681 (O_2681,N_49138,N_47595);
xor UO_2682 (O_2682,N_47597,N_49124);
xnor UO_2683 (O_2683,N_48166,N_47822);
nor UO_2684 (O_2684,N_48314,N_49415);
nor UO_2685 (O_2685,N_48435,N_48462);
and UO_2686 (O_2686,N_49990,N_49916);
and UO_2687 (O_2687,N_49469,N_47830);
xor UO_2688 (O_2688,N_49831,N_48193);
xnor UO_2689 (O_2689,N_48755,N_48715);
or UO_2690 (O_2690,N_48635,N_49935);
nor UO_2691 (O_2691,N_47880,N_47581);
or UO_2692 (O_2692,N_47660,N_47936);
nor UO_2693 (O_2693,N_49750,N_49803);
or UO_2694 (O_2694,N_47729,N_47922);
xnor UO_2695 (O_2695,N_49662,N_48351);
nand UO_2696 (O_2696,N_49714,N_49258);
nand UO_2697 (O_2697,N_49911,N_47649);
and UO_2698 (O_2698,N_48351,N_47664);
nor UO_2699 (O_2699,N_48453,N_48607);
nand UO_2700 (O_2700,N_48780,N_48207);
nand UO_2701 (O_2701,N_48239,N_48900);
nor UO_2702 (O_2702,N_47535,N_49796);
nor UO_2703 (O_2703,N_49991,N_49433);
or UO_2704 (O_2704,N_49418,N_49818);
nor UO_2705 (O_2705,N_49388,N_49536);
nor UO_2706 (O_2706,N_49353,N_48828);
nand UO_2707 (O_2707,N_48864,N_49540);
nor UO_2708 (O_2708,N_47590,N_49207);
and UO_2709 (O_2709,N_47993,N_49920);
nor UO_2710 (O_2710,N_47664,N_49066);
nor UO_2711 (O_2711,N_47859,N_47882);
or UO_2712 (O_2712,N_47751,N_47924);
nor UO_2713 (O_2713,N_47737,N_47810);
and UO_2714 (O_2714,N_48253,N_49789);
nand UO_2715 (O_2715,N_48124,N_47556);
or UO_2716 (O_2716,N_47525,N_47857);
nor UO_2717 (O_2717,N_49084,N_49754);
nor UO_2718 (O_2718,N_48681,N_48614);
nor UO_2719 (O_2719,N_48195,N_48030);
or UO_2720 (O_2720,N_49489,N_48645);
and UO_2721 (O_2721,N_48794,N_49008);
and UO_2722 (O_2722,N_47854,N_49909);
and UO_2723 (O_2723,N_48660,N_48724);
or UO_2724 (O_2724,N_49546,N_48134);
or UO_2725 (O_2725,N_49380,N_49780);
and UO_2726 (O_2726,N_48054,N_48779);
and UO_2727 (O_2727,N_49227,N_49002);
nand UO_2728 (O_2728,N_47743,N_49182);
or UO_2729 (O_2729,N_47516,N_49840);
nand UO_2730 (O_2730,N_48157,N_49018);
nor UO_2731 (O_2731,N_48483,N_49511);
and UO_2732 (O_2732,N_47716,N_49853);
and UO_2733 (O_2733,N_49146,N_48190);
and UO_2734 (O_2734,N_49569,N_49058);
nor UO_2735 (O_2735,N_49837,N_48197);
nand UO_2736 (O_2736,N_49141,N_48854);
and UO_2737 (O_2737,N_47851,N_48710);
nand UO_2738 (O_2738,N_48945,N_49537);
nor UO_2739 (O_2739,N_47941,N_49182);
nand UO_2740 (O_2740,N_48253,N_47888);
or UO_2741 (O_2741,N_48343,N_47805);
nor UO_2742 (O_2742,N_47702,N_49565);
and UO_2743 (O_2743,N_49466,N_49846);
nand UO_2744 (O_2744,N_49879,N_49866);
and UO_2745 (O_2745,N_47742,N_49524);
or UO_2746 (O_2746,N_49351,N_48488);
nor UO_2747 (O_2747,N_48733,N_49673);
or UO_2748 (O_2748,N_48064,N_48099);
nor UO_2749 (O_2749,N_49392,N_49560);
nor UO_2750 (O_2750,N_47575,N_48195);
xor UO_2751 (O_2751,N_48636,N_48664);
or UO_2752 (O_2752,N_49213,N_48922);
nand UO_2753 (O_2753,N_48463,N_49990);
nand UO_2754 (O_2754,N_48526,N_47840);
or UO_2755 (O_2755,N_49321,N_49627);
and UO_2756 (O_2756,N_49058,N_49892);
or UO_2757 (O_2757,N_48424,N_49337);
nor UO_2758 (O_2758,N_47859,N_48824);
or UO_2759 (O_2759,N_47647,N_49905);
and UO_2760 (O_2760,N_49787,N_49537);
and UO_2761 (O_2761,N_47677,N_48905);
nand UO_2762 (O_2762,N_48287,N_49352);
nand UO_2763 (O_2763,N_49039,N_49662);
nor UO_2764 (O_2764,N_48415,N_49924);
or UO_2765 (O_2765,N_49151,N_47832);
or UO_2766 (O_2766,N_48407,N_49714);
or UO_2767 (O_2767,N_49747,N_49396);
or UO_2768 (O_2768,N_47988,N_49308);
nand UO_2769 (O_2769,N_49356,N_48245);
nor UO_2770 (O_2770,N_47901,N_48395);
xnor UO_2771 (O_2771,N_48651,N_47978);
xnor UO_2772 (O_2772,N_48511,N_47825);
xnor UO_2773 (O_2773,N_47909,N_49177);
or UO_2774 (O_2774,N_49129,N_48109);
nand UO_2775 (O_2775,N_48006,N_47979);
and UO_2776 (O_2776,N_49367,N_48423);
and UO_2777 (O_2777,N_48696,N_48744);
nor UO_2778 (O_2778,N_48146,N_48518);
xnor UO_2779 (O_2779,N_49668,N_49289);
and UO_2780 (O_2780,N_49326,N_48781);
and UO_2781 (O_2781,N_48895,N_48147);
nor UO_2782 (O_2782,N_47815,N_48529);
and UO_2783 (O_2783,N_47774,N_48735);
and UO_2784 (O_2784,N_48863,N_48313);
or UO_2785 (O_2785,N_47746,N_49512);
and UO_2786 (O_2786,N_48535,N_48868);
nor UO_2787 (O_2787,N_49339,N_49889);
nand UO_2788 (O_2788,N_48694,N_48592);
nand UO_2789 (O_2789,N_49607,N_49089);
xnor UO_2790 (O_2790,N_49365,N_47944);
and UO_2791 (O_2791,N_47568,N_48833);
or UO_2792 (O_2792,N_47606,N_48717);
nor UO_2793 (O_2793,N_47719,N_47872);
nand UO_2794 (O_2794,N_48915,N_47763);
or UO_2795 (O_2795,N_49997,N_48611);
and UO_2796 (O_2796,N_49249,N_48811);
nand UO_2797 (O_2797,N_49882,N_48978);
nor UO_2798 (O_2798,N_48711,N_49301);
nor UO_2799 (O_2799,N_49861,N_48731);
and UO_2800 (O_2800,N_49871,N_49702);
nand UO_2801 (O_2801,N_48965,N_49706);
nor UO_2802 (O_2802,N_47608,N_49618);
and UO_2803 (O_2803,N_47984,N_48531);
nor UO_2804 (O_2804,N_48470,N_49577);
and UO_2805 (O_2805,N_47809,N_48008);
and UO_2806 (O_2806,N_48109,N_49487);
xnor UO_2807 (O_2807,N_47858,N_48035);
or UO_2808 (O_2808,N_49205,N_49548);
or UO_2809 (O_2809,N_48072,N_47784);
nor UO_2810 (O_2810,N_47774,N_48660);
xnor UO_2811 (O_2811,N_49086,N_49492);
and UO_2812 (O_2812,N_47960,N_49371);
and UO_2813 (O_2813,N_47824,N_48908);
nand UO_2814 (O_2814,N_47690,N_49941);
nand UO_2815 (O_2815,N_49800,N_49243);
nor UO_2816 (O_2816,N_49708,N_49467);
or UO_2817 (O_2817,N_48351,N_49939);
or UO_2818 (O_2818,N_48143,N_47633);
nand UO_2819 (O_2819,N_49124,N_48763);
or UO_2820 (O_2820,N_49402,N_47579);
nor UO_2821 (O_2821,N_47591,N_47759);
xor UO_2822 (O_2822,N_49894,N_49502);
xor UO_2823 (O_2823,N_49523,N_48962);
nand UO_2824 (O_2824,N_49605,N_48801);
nor UO_2825 (O_2825,N_47595,N_49355);
nand UO_2826 (O_2826,N_47687,N_49496);
nand UO_2827 (O_2827,N_49865,N_48165);
or UO_2828 (O_2828,N_49477,N_48760);
and UO_2829 (O_2829,N_49964,N_49072);
nand UO_2830 (O_2830,N_49526,N_49473);
or UO_2831 (O_2831,N_47976,N_47987);
nand UO_2832 (O_2832,N_47627,N_49222);
and UO_2833 (O_2833,N_48820,N_49030);
or UO_2834 (O_2834,N_48006,N_48990);
or UO_2835 (O_2835,N_49593,N_47847);
or UO_2836 (O_2836,N_48460,N_49020);
nand UO_2837 (O_2837,N_49594,N_47680);
nor UO_2838 (O_2838,N_49416,N_49104);
xnor UO_2839 (O_2839,N_47520,N_48946);
nor UO_2840 (O_2840,N_48857,N_49038);
nor UO_2841 (O_2841,N_48625,N_49631);
and UO_2842 (O_2842,N_48570,N_47978);
or UO_2843 (O_2843,N_49777,N_49698);
and UO_2844 (O_2844,N_48703,N_47746);
or UO_2845 (O_2845,N_49121,N_48430);
or UO_2846 (O_2846,N_49470,N_48437);
nor UO_2847 (O_2847,N_49330,N_49598);
or UO_2848 (O_2848,N_48078,N_49875);
or UO_2849 (O_2849,N_48475,N_48308);
nor UO_2850 (O_2850,N_49373,N_49187);
nand UO_2851 (O_2851,N_49410,N_47815);
and UO_2852 (O_2852,N_48024,N_49894);
nand UO_2853 (O_2853,N_49936,N_49788);
or UO_2854 (O_2854,N_49422,N_48593);
nor UO_2855 (O_2855,N_49042,N_49451);
and UO_2856 (O_2856,N_49351,N_47742);
and UO_2857 (O_2857,N_47842,N_48663);
and UO_2858 (O_2858,N_48965,N_48517);
and UO_2859 (O_2859,N_47701,N_49939);
nand UO_2860 (O_2860,N_47586,N_49899);
nor UO_2861 (O_2861,N_47573,N_48260);
or UO_2862 (O_2862,N_47573,N_48047);
and UO_2863 (O_2863,N_49156,N_49807);
and UO_2864 (O_2864,N_48431,N_49831);
or UO_2865 (O_2865,N_47635,N_49206);
xnor UO_2866 (O_2866,N_48362,N_47898);
or UO_2867 (O_2867,N_48700,N_47815);
nand UO_2868 (O_2868,N_48829,N_48636);
xor UO_2869 (O_2869,N_48653,N_49179);
nand UO_2870 (O_2870,N_49453,N_47789);
or UO_2871 (O_2871,N_49289,N_48874);
nand UO_2872 (O_2872,N_48563,N_49189);
nor UO_2873 (O_2873,N_48856,N_49598);
and UO_2874 (O_2874,N_48196,N_49353);
nand UO_2875 (O_2875,N_48684,N_49577);
nand UO_2876 (O_2876,N_47552,N_49971);
nand UO_2877 (O_2877,N_49720,N_49759);
nor UO_2878 (O_2878,N_48061,N_48218);
nor UO_2879 (O_2879,N_48536,N_49541);
and UO_2880 (O_2880,N_47733,N_49532);
or UO_2881 (O_2881,N_48904,N_48165);
nand UO_2882 (O_2882,N_48025,N_49768);
xor UO_2883 (O_2883,N_49460,N_48264);
xor UO_2884 (O_2884,N_48950,N_47826);
and UO_2885 (O_2885,N_49800,N_49351);
and UO_2886 (O_2886,N_49126,N_48069);
nor UO_2887 (O_2887,N_48224,N_49535);
xor UO_2888 (O_2888,N_47987,N_49888);
or UO_2889 (O_2889,N_48580,N_49535);
or UO_2890 (O_2890,N_48369,N_48602);
nor UO_2891 (O_2891,N_48444,N_49508);
nor UO_2892 (O_2892,N_48495,N_48095);
or UO_2893 (O_2893,N_49509,N_49602);
or UO_2894 (O_2894,N_49739,N_49206);
nand UO_2895 (O_2895,N_48386,N_48357);
nor UO_2896 (O_2896,N_49618,N_48024);
or UO_2897 (O_2897,N_48484,N_47850);
or UO_2898 (O_2898,N_48930,N_48436);
nor UO_2899 (O_2899,N_47782,N_49918);
xnor UO_2900 (O_2900,N_49354,N_48323);
nor UO_2901 (O_2901,N_48778,N_48731);
nor UO_2902 (O_2902,N_49770,N_48612);
nor UO_2903 (O_2903,N_48032,N_49412);
nand UO_2904 (O_2904,N_49106,N_49569);
nand UO_2905 (O_2905,N_49930,N_49357);
xnor UO_2906 (O_2906,N_48646,N_48919);
nand UO_2907 (O_2907,N_49347,N_49834);
and UO_2908 (O_2908,N_49560,N_48644);
xnor UO_2909 (O_2909,N_48709,N_49542);
nor UO_2910 (O_2910,N_49456,N_49814);
nor UO_2911 (O_2911,N_49245,N_49509);
and UO_2912 (O_2912,N_49194,N_48346);
nand UO_2913 (O_2913,N_49532,N_48912);
nand UO_2914 (O_2914,N_47963,N_49928);
or UO_2915 (O_2915,N_47953,N_49149);
nand UO_2916 (O_2916,N_48092,N_48579);
and UO_2917 (O_2917,N_49197,N_47694);
nor UO_2918 (O_2918,N_47898,N_49288);
and UO_2919 (O_2919,N_49402,N_47788);
or UO_2920 (O_2920,N_47918,N_48679);
nor UO_2921 (O_2921,N_48606,N_49291);
and UO_2922 (O_2922,N_49443,N_49878);
xnor UO_2923 (O_2923,N_48870,N_49966);
or UO_2924 (O_2924,N_48337,N_48010);
and UO_2925 (O_2925,N_48726,N_48246);
nor UO_2926 (O_2926,N_48823,N_49007);
nand UO_2927 (O_2927,N_47674,N_48130);
nor UO_2928 (O_2928,N_49344,N_49981);
and UO_2929 (O_2929,N_48793,N_49055);
xor UO_2930 (O_2930,N_49418,N_48536);
nor UO_2931 (O_2931,N_49681,N_49987);
and UO_2932 (O_2932,N_48330,N_49407);
nor UO_2933 (O_2933,N_47668,N_49967);
and UO_2934 (O_2934,N_48192,N_49150);
and UO_2935 (O_2935,N_48814,N_49453);
nor UO_2936 (O_2936,N_49824,N_49675);
nand UO_2937 (O_2937,N_48605,N_49991);
nor UO_2938 (O_2938,N_48786,N_48887);
nor UO_2939 (O_2939,N_48711,N_49558);
nor UO_2940 (O_2940,N_47978,N_47929);
and UO_2941 (O_2941,N_48988,N_48494);
and UO_2942 (O_2942,N_48620,N_48291);
xor UO_2943 (O_2943,N_49988,N_49966);
nand UO_2944 (O_2944,N_47773,N_49405);
nand UO_2945 (O_2945,N_48584,N_47798);
or UO_2946 (O_2946,N_48166,N_48154);
and UO_2947 (O_2947,N_49701,N_49430);
nor UO_2948 (O_2948,N_47804,N_48197);
or UO_2949 (O_2949,N_48813,N_48595);
nor UO_2950 (O_2950,N_49915,N_48256);
xor UO_2951 (O_2951,N_48873,N_48610);
nand UO_2952 (O_2952,N_47709,N_48629);
and UO_2953 (O_2953,N_49114,N_47732);
or UO_2954 (O_2954,N_49604,N_48984);
and UO_2955 (O_2955,N_49251,N_49987);
nor UO_2956 (O_2956,N_47756,N_47623);
or UO_2957 (O_2957,N_48729,N_47970);
and UO_2958 (O_2958,N_49646,N_47825);
or UO_2959 (O_2959,N_48978,N_48779);
and UO_2960 (O_2960,N_49737,N_49358);
nor UO_2961 (O_2961,N_49858,N_49687);
or UO_2962 (O_2962,N_48506,N_48663);
nor UO_2963 (O_2963,N_47714,N_49705);
or UO_2964 (O_2964,N_47807,N_49742);
nor UO_2965 (O_2965,N_49458,N_48610);
or UO_2966 (O_2966,N_48345,N_47815);
xnor UO_2967 (O_2967,N_47900,N_48114);
nand UO_2968 (O_2968,N_49723,N_48408);
nand UO_2969 (O_2969,N_48209,N_49233);
xor UO_2970 (O_2970,N_47972,N_48801);
nand UO_2971 (O_2971,N_48987,N_48959);
or UO_2972 (O_2972,N_48722,N_48080);
or UO_2973 (O_2973,N_49563,N_47711);
and UO_2974 (O_2974,N_48519,N_49214);
nand UO_2975 (O_2975,N_48907,N_48348);
nand UO_2976 (O_2976,N_49500,N_48347);
and UO_2977 (O_2977,N_48677,N_48953);
nand UO_2978 (O_2978,N_48008,N_49858);
nor UO_2979 (O_2979,N_47510,N_47896);
nand UO_2980 (O_2980,N_48572,N_47544);
nor UO_2981 (O_2981,N_48488,N_49341);
and UO_2982 (O_2982,N_48161,N_48340);
or UO_2983 (O_2983,N_47767,N_48836);
nor UO_2984 (O_2984,N_48354,N_48398);
xor UO_2985 (O_2985,N_47592,N_49319);
nor UO_2986 (O_2986,N_47521,N_48970);
nand UO_2987 (O_2987,N_47708,N_49477);
or UO_2988 (O_2988,N_49000,N_49971);
and UO_2989 (O_2989,N_48005,N_48584);
and UO_2990 (O_2990,N_48314,N_49251);
nand UO_2991 (O_2991,N_47905,N_48638);
and UO_2992 (O_2992,N_49690,N_49263);
or UO_2993 (O_2993,N_49842,N_48543);
or UO_2994 (O_2994,N_49548,N_49849);
nor UO_2995 (O_2995,N_48711,N_49717);
nand UO_2996 (O_2996,N_49160,N_48444);
or UO_2997 (O_2997,N_48169,N_48701);
nand UO_2998 (O_2998,N_49995,N_48654);
or UO_2999 (O_2999,N_48867,N_49498);
or UO_3000 (O_3000,N_47750,N_48019);
nand UO_3001 (O_3001,N_48960,N_48295);
nor UO_3002 (O_3002,N_49088,N_49141);
nor UO_3003 (O_3003,N_48991,N_48160);
nand UO_3004 (O_3004,N_48090,N_47828);
or UO_3005 (O_3005,N_48816,N_48555);
and UO_3006 (O_3006,N_48574,N_48071);
and UO_3007 (O_3007,N_49333,N_48328);
nand UO_3008 (O_3008,N_48819,N_47948);
and UO_3009 (O_3009,N_48211,N_48893);
and UO_3010 (O_3010,N_48795,N_49892);
and UO_3011 (O_3011,N_47590,N_47966);
and UO_3012 (O_3012,N_49203,N_49517);
nand UO_3013 (O_3013,N_48071,N_48883);
and UO_3014 (O_3014,N_49294,N_47898);
nand UO_3015 (O_3015,N_48900,N_49504);
or UO_3016 (O_3016,N_47982,N_47761);
or UO_3017 (O_3017,N_48468,N_48484);
nor UO_3018 (O_3018,N_48801,N_47549);
nand UO_3019 (O_3019,N_48525,N_47711);
or UO_3020 (O_3020,N_47541,N_49437);
or UO_3021 (O_3021,N_49714,N_49726);
and UO_3022 (O_3022,N_49894,N_49694);
nor UO_3023 (O_3023,N_47598,N_49862);
or UO_3024 (O_3024,N_48805,N_49937);
nor UO_3025 (O_3025,N_49860,N_47682);
nor UO_3026 (O_3026,N_49964,N_49598);
or UO_3027 (O_3027,N_49190,N_49087);
nand UO_3028 (O_3028,N_48627,N_48356);
nand UO_3029 (O_3029,N_49890,N_48210);
or UO_3030 (O_3030,N_48681,N_48753);
nor UO_3031 (O_3031,N_49630,N_49045);
and UO_3032 (O_3032,N_47523,N_48279);
and UO_3033 (O_3033,N_48136,N_49084);
nor UO_3034 (O_3034,N_49820,N_47883);
nor UO_3035 (O_3035,N_47842,N_47823);
and UO_3036 (O_3036,N_49228,N_49229);
or UO_3037 (O_3037,N_49911,N_49112);
xor UO_3038 (O_3038,N_49481,N_49511);
and UO_3039 (O_3039,N_49687,N_49444);
or UO_3040 (O_3040,N_48085,N_47758);
and UO_3041 (O_3041,N_49950,N_49458);
nand UO_3042 (O_3042,N_48755,N_48949);
xor UO_3043 (O_3043,N_48778,N_49539);
xnor UO_3044 (O_3044,N_49048,N_48676);
and UO_3045 (O_3045,N_47642,N_49198);
or UO_3046 (O_3046,N_48123,N_49290);
nor UO_3047 (O_3047,N_49197,N_49248);
or UO_3048 (O_3048,N_49591,N_49774);
and UO_3049 (O_3049,N_48117,N_48172);
or UO_3050 (O_3050,N_48652,N_47659);
or UO_3051 (O_3051,N_48442,N_49205);
nand UO_3052 (O_3052,N_48178,N_48242);
nand UO_3053 (O_3053,N_49685,N_49701);
xnor UO_3054 (O_3054,N_49023,N_49953);
and UO_3055 (O_3055,N_49794,N_49176);
and UO_3056 (O_3056,N_47727,N_48488);
and UO_3057 (O_3057,N_48853,N_47801);
xnor UO_3058 (O_3058,N_48806,N_48904);
nor UO_3059 (O_3059,N_48864,N_49400);
xor UO_3060 (O_3060,N_48007,N_48254);
xnor UO_3061 (O_3061,N_47953,N_48036);
nand UO_3062 (O_3062,N_49339,N_48060);
and UO_3063 (O_3063,N_47615,N_48667);
nand UO_3064 (O_3064,N_47627,N_48514);
nor UO_3065 (O_3065,N_49209,N_49993);
or UO_3066 (O_3066,N_48073,N_48994);
xor UO_3067 (O_3067,N_48781,N_48752);
nand UO_3068 (O_3068,N_48278,N_48488);
xor UO_3069 (O_3069,N_47863,N_49417);
nand UO_3070 (O_3070,N_48661,N_47900);
nor UO_3071 (O_3071,N_49512,N_48925);
nor UO_3072 (O_3072,N_47674,N_48172);
nor UO_3073 (O_3073,N_49596,N_48738);
or UO_3074 (O_3074,N_49141,N_47568);
nor UO_3075 (O_3075,N_49989,N_49144);
xor UO_3076 (O_3076,N_48273,N_47810);
and UO_3077 (O_3077,N_49380,N_48349);
or UO_3078 (O_3078,N_48457,N_48753);
and UO_3079 (O_3079,N_48718,N_49680);
nor UO_3080 (O_3080,N_48181,N_48910);
or UO_3081 (O_3081,N_49656,N_49876);
nand UO_3082 (O_3082,N_47520,N_49472);
nand UO_3083 (O_3083,N_49741,N_47744);
and UO_3084 (O_3084,N_48371,N_48549);
or UO_3085 (O_3085,N_48097,N_48138);
nor UO_3086 (O_3086,N_49811,N_48014);
or UO_3087 (O_3087,N_48229,N_49386);
xnor UO_3088 (O_3088,N_49005,N_48584);
or UO_3089 (O_3089,N_49512,N_48662);
nor UO_3090 (O_3090,N_47997,N_48244);
and UO_3091 (O_3091,N_49439,N_48784);
nor UO_3092 (O_3092,N_49978,N_48264);
nand UO_3093 (O_3093,N_49788,N_49822);
xnor UO_3094 (O_3094,N_47952,N_48402);
or UO_3095 (O_3095,N_48457,N_47883);
and UO_3096 (O_3096,N_49132,N_47706);
or UO_3097 (O_3097,N_49198,N_49873);
nand UO_3098 (O_3098,N_49627,N_49551);
and UO_3099 (O_3099,N_47865,N_49791);
or UO_3100 (O_3100,N_48796,N_48649);
nand UO_3101 (O_3101,N_47546,N_49631);
and UO_3102 (O_3102,N_48624,N_48967);
nor UO_3103 (O_3103,N_47999,N_49677);
nor UO_3104 (O_3104,N_49752,N_47854);
nand UO_3105 (O_3105,N_48902,N_48530);
nor UO_3106 (O_3106,N_48768,N_49398);
or UO_3107 (O_3107,N_48942,N_48355);
and UO_3108 (O_3108,N_47992,N_47866);
or UO_3109 (O_3109,N_48465,N_47592);
and UO_3110 (O_3110,N_47539,N_49824);
and UO_3111 (O_3111,N_48755,N_49952);
xor UO_3112 (O_3112,N_47881,N_49638);
or UO_3113 (O_3113,N_48683,N_49852);
nand UO_3114 (O_3114,N_47619,N_47578);
nor UO_3115 (O_3115,N_49129,N_49390);
or UO_3116 (O_3116,N_49608,N_48434);
nor UO_3117 (O_3117,N_48260,N_49835);
nor UO_3118 (O_3118,N_49498,N_47506);
or UO_3119 (O_3119,N_49958,N_48117);
and UO_3120 (O_3120,N_48765,N_49367);
or UO_3121 (O_3121,N_48783,N_47722);
or UO_3122 (O_3122,N_47719,N_49030);
and UO_3123 (O_3123,N_47918,N_49900);
or UO_3124 (O_3124,N_47625,N_48100);
nor UO_3125 (O_3125,N_47959,N_49503);
nand UO_3126 (O_3126,N_48043,N_49124);
or UO_3127 (O_3127,N_47568,N_49057);
or UO_3128 (O_3128,N_49376,N_49070);
nand UO_3129 (O_3129,N_48129,N_48649);
nand UO_3130 (O_3130,N_48597,N_48858);
or UO_3131 (O_3131,N_49204,N_47677);
nor UO_3132 (O_3132,N_47550,N_47690);
nor UO_3133 (O_3133,N_49845,N_49011);
or UO_3134 (O_3134,N_48430,N_48999);
nand UO_3135 (O_3135,N_48105,N_49595);
nand UO_3136 (O_3136,N_47585,N_49988);
nand UO_3137 (O_3137,N_47854,N_48281);
or UO_3138 (O_3138,N_48068,N_48984);
or UO_3139 (O_3139,N_48122,N_49426);
nand UO_3140 (O_3140,N_49116,N_49898);
nand UO_3141 (O_3141,N_47673,N_47893);
and UO_3142 (O_3142,N_49361,N_48397);
and UO_3143 (O_3143,N_49726,N_47946);
xnor UO_3144 (O_3144,N_49085,N_48384);
or UO_3145 (O_3145,N_49571,N_49934);
nor UO_3146 (O_3146,N_48873,N_48082);
nor UO_3147 (O_3147,N_49688,N_49515);
and UO_3148 (O_3148,N_47831,N_48863);
nand UO_3149 (O_3149,N_48099,N_48480);
nand UO_3150 (O_3150,N_47730,N_49699);
xor UO_3151 (O_3151,N_48872,N_48344);
and UO_3152 (O_3152,N_49014,N_48732);
nand UO_3153 (O_3153,N_47642,N_48170);
nand UO_3154 (O_3154,N_49518,N_49884);
and UO_3155 (O_3155,N_48076,N_47805);
or UO_3156 (O_3156,N_47874,N_48775);
nand UO_3157 (O_3157,N_48000,N_47661);
nor UO_3158 (O_3158,N_49105,N_47587);
nor UO_3159 (O_3159,N_48199,N_48879);
and UO_3160 (O_3160,N_48769,N_48355);
nand UO_3161 (O_3161,N_49001,N_48150);
or UO_3162 (O_3162,N_49739,N_49526);
and UO_3163 (O_3163,N_49648,N_47718);
xor UO_3164 (O_3164,N_49003,N_48714);
nand UO_3165 (O_3165,N_48035,N_49482);
and UO_3166 (O_3166,N_49235,N_49268);
nand UO_3167 (O_3167,N_49147,N_48692);
or UO_3168 (O_3168,N_47597,N_47905);
xor UO_3169 (O_3169,N_48385,N_49766);
nor UO_3170 (O_3170,N_48411,N_49421);
xnor UO_3171 (O_3171,N_47679,N_47971);
nand UO_3172 (O_3172,N_48805,N_48701);
and UO_3173 (O_3173,N_47510,N_48238);
or UO_3174 (O_3174,N_49106,N_49867);
nor UO_3175 (O_3175,N_48821,N_49894);
xor UO_3176 (O_3176,N_47649,N_49249);
xnor UO_3177 (O_3177,N_48744,N_48321);
nor UO_3178 (O_3178,N_49111,N_47619);
or UO_3179 (O_3179,N_49343,N_47797);
or UO_3180 (O_3180,N_48546,N_49932);
nand UO_3181 (O_3181,N_47773,N_49066);
nor UO_3182 (O_3182,N_49552,N_48019);
nor UO_3183 (O_3183,N_47874,N_47866);
and UO_3184 (O_3184,N_49914,N_49585);
and UO_3185 (O_3185,N_49943,N_48138);
and UO_3186 (O_3186,N_48325,N_48315);
and UO_3187 (O_3187,N_49959,N_49190);
nand UO_3188 (O_3188,N_48702,N_49365);
and UO_3189 (O_3189,N_48225,N_49049);
nand UO_3190 (O_3190,N_49899,N_48363);
xor UO_3191 (O_3191,N_49259,N_48410);
nor UO_3192 (O_3192,N_48895,N_49239);
and UO_3193 (O_3193,N_48313,N_49183);
nand UO_3194 (O_3194,N_49582,N_49610);
nand UO_3195 (O_3195,N_47884,N_49729);
nor UO_3196 (O_3196,N_49009,N_47713);
nor UO_3197 (O_3197,N_48970,N_48147);
and UO_3198 (O_3198,N_48339,N_49678);
or UO_3199 (O_3199,N_47986,N_48056);
or UO_3200 (O_3200,N_48257,N_48812);
or UO_3201 (O_3201,N_49471,N_48620);
and UO_3202 (O_3202,N_49397,N_49226);
nor UO_3203 (O_3203,N_48970,N_49258);
or UO_3204 (O_3204,N_49942,N_49360);
xnor UO_3205 (O_3205,N_48114,N_48595);
xor UO_3206 (O_3206,N_49504,N_48964);
or UO_3207 (O_3207,N_49175,N_47919);
or UO_3208 (O_3208,N_49542,N_47585);
or UO_3209 (O_3209,N_49410,N_48272);
or UO_3210 (O_3210,N_48994,N_47597);
and UO_3211 (O_3211,N_49039,N_49390);
xnor UO_3212 (O_3212,N_48305,N_49230);
nand UO_3213 (O_3213,N_48670,N_48050);
nor UO_3214 (O_3214,N_49101,N_48349);
and UO_3215 (O_3215,N_48286,N_47588);
nand UO_3216 (O_3216,N_48564,N_47647);
and UO_3217 (O_3217,N_49133,N_48037);
or UO_3218 (O_3218,N_48446,N_48444);
and UO_3219 (O_3219,N_49373,N_49771);
or UO_3220 (O_3220,N_49005,N_48618);
nand UO_3221 (O_3221,N_49623,N_49420);
or UO_3222 (O_3222,N_47787,N_48792);
or UO_3223 (O_3223,N_49102,N_48297);
nand UO_3224 (O_3224,N_47744,N_49240);
xor UO_3225 (O_3225,N_47966,N_47537);
nand UO_3226 (O_3226,N_48850,N_49718);
or UO_3227 (O_3227,N_48537,N_49442);
nand UO_3228 (O_3228,N_49913,N_48405);
nand UO_3229 (O_3229,N_48985,N_48684);
and UO_3230 (O_3230,N_48456,N_49310);
nand UO_3231 (O_3231,N_47579,N_47550);
and UO_3232 (O_3232,N_49739,N_47691);
xor UO_3233 (O_3233,N_49874,N_47764);
nand UO_3234 (O_3234,N_47999,N_47560);
or UO_3235 (O_3235,N_47779,N_47919);
or UO_3236 (O_3236,N_47600,N_49033);
or UO_3237 (O_3237,N_49954,N_47512);
or UO_3238 (O_3238,N_49019,N_49602);
xnor UO_3239 (O_3239,N_49095,N_48327);
nand UO_3240 (O_3240,N_49452,N_49987);
nor UO_3241 (O_3241,N_49552,N_49770);
and UO_3242 (O_3242,N_47589,N_49710);
nand UO_3243 (O_3243,N_49758,N_47799);
nand UO_3244 (O_3244,N_47724,N_47854);
nand UO_3245 (O_3245,N_49208,N_47819);
or UO_3246 (O_3246,N_48164,N_48419);
nand UO_3247 (O_3247,N_49000,N_49180);
nand UO_3248 (O_3248,N_47904,N_49278);
and UO_3249 (O_3249,N_49636,N_49627);
nand UO_3250 (O_3250,N_49417,N_48418);
nor UO_3251 (O_3251,N_49863,N_49985);
or UO_3252 (O_3252,N_49456,N_48940);
nor UO_3253 (O_3253,N_49499,N_49419);
or UO_3254 (O_3254,N_48557,N_49782);
and UO_3255 (O_3255,N_49909,N_47888);
nor UO_3256 (O_3256,N_47518,N_49745);
nand UO_3257 (O_3257,N_48453,N_48405);
and UO_3258 (O_3258,N_48580,N_49705);
nor UO_3259 (O_3259,N_48002,N_48909);
xor UO_3260 (O_3260,N_47935,N_47735);
xnor UO_3261 (O_3261,N_49971,N_49341);
or UO_3262 (O_3262,N_47945,N_49635);
and UO_3263 (O_3263,N_47994,N_48196);
nor UO_3264 (O_3264,N_48676,N_48434);
nand UO_3265 (O_3265,N_47585,N_49162);
nand UO_3266 (O_3266,N_48611,N_49598);
nand UO_3267 (O_3267,N_48149,N_48903);
and UO_3268 (O_3268,N_48964,N_48396);
nand UO_3269 (O_3269,N_49707,N_47856);
nand UO_3270 (O_3270,N_48943,N_49392);
nor UO_3271 (O_3271,N_48717,N_49678);
xor UO_3272 (O_3272,N_49373,N_49643);
nand UO_3273 (O_3273,N_49396,N_48557);
and UO_3274 (O_3274,N_48235,N_48960);
nand UO_3275 (O_3275,N_48463,N_49706);
nor UO_3276 (O_3276,N_48742,N_48177);
nor UO_3277 (O_3277,N_48313,N_47749);
nand UO_3278 (O_3278,N_48683,N_47670);
and UO_3279 (O_3279,N_49822,N_49955);
or UO_3280 (O_3280,N_47755,N_48628);
nor UO_3281 (O_3281,N_49326,N_49125);
or UO_3282 (O_3282,N_48524,N_48136);
nand UO_3283 (O_3283,N_49532,N_48296);
or UO_3284 (O_3284,N_48192,N_49313);
and UO_3285 (O_3285,N_49570,N_47864);
nand UO_3286 (O_3286,N_48834,N_49989);
nand UO_3287 (O_3287,N_48276,N_49042);
nor UO_3288 (O_3288,N_48584,N_49479);
nand UO_3289 (O_3289,N_49744,N_47884);
nor UO_3290 (O_3290,N_48915,N_49264);
and UO_3291 (O_3291,N_47670,N_49950);
nor UO_3292 (O_3292,N_48959,N_48776);
xor UO_3293 (O_3293,N_49292,N_49387);
nor UO_3294 (O_3294,N_48150,N_49456);
or UO_3295 (O_3295,N_48404,N_49144);
nor UO_3296 (O_3296,N_49643,N_49080);
nand UO_3297 (O_3297,N_48926,N_48538);
nor UO_3298 (O_3298,N_47581,N_48952);
and UO_3299 (O_3299,N_47952,N_48669);
nand UO_3300 (O_3300,N_49665,N_48933);
and UO_3301 (O_3301,N_49140,N_48784);
nand UO_3302 (O_3302,N_47803,N_48214);
or UO_3303 (O_3303,N_48521,N_48865);
and UO_3304 (O_3304,N_49729,N_48709);
and UO_3305 (O_3305,N_49257,N_49568);
or UO_3306 (O_3306,N_47734,N_49572);
nor UO_3307 (O_3307,N_49345,N_49986);
xnor UO_3308 (O_3308,N_48730,N_49558);
nand UO_3309 (O_3309,N_49075,N_48919);
and UO_3310 (O_3310,N_49165,N_49889);
nand UO_3311 (O_3311,N_48259,N_49450);
nand UO_3312 (O_3312,N_48118,N_49333);
or UO_3313 (O_3313,N_48687,N_48123);
and UO_3314 (O_3314,N_47780,N_48777);
xnor UO_3315 (O_3315,N_49729,N_49232);
nor UO_3316 (O_3316,N_49372,N_48528);
nand UO_3317 (O_3317,N_49006,N_48212);
or UO_3318 (O_3318,N_47778,N_48903);
or UO_3319 (O_3319,N_48206,N_49601);
nand UO_3320 (O_3320,N_48200,N_49723);
nor UO_3321 (O_3321,N_49420,N_48266);
or UO_3322 (O_3322,N_48981,N_48145);
nand UO_3323 (O_3323,N_49229,N_49609);
nor UO_3324 (O_3324,N_49799,N_47697);
or UO_3325 (O_3325,N_49649,N_49890);
and UO_3326 (O_3326,N_49056,N_48243);
nand UO_3327 (O_3327,N_48164,N_48518);
nor UO_3328 (O_3328,N_47624,N_48790);
and UO_3329 (O_3329,N_48553,N_47776);
or UO_3330 (O_3330,N_48477,N_49053);
and UO_3331 (O_3331,N_49086,N_48999);
or UO_3332 (O_3332,N_47864,N_49500);
nor UO_3333 (O_3333,N_48239,N_49977);
nor UO_3334 (O_3334,N_47763,N_48688);
and UO_3335 (O_3335,N_48296,N_48466);
or UO_3336 (O_3336,N_48487,N_47579);
or UO_3337 (O_3337,N_49433,N_49485);
nand UO_3338 (O_3338,N_49701,N_47733);
xor UO_3339 (O_3339,N_47828,N_49466);
xor UO_3340 (O_3340,N_48365,N_48565);
or UO_3341 (O_3341,N_48846,N_48132);
nand UO_3342 (O_3342,N_48335,N_48534);
xor UO_3343 (O_3343,N_47829,N_47587);
and UO_3344 (O_3344,N_47685,N_49146);
nand UO_3345 (O_3345,N_48797,N_49028);
and UO_3346 (O_3346,N_48101,N_47627);
or UO_3347 (O_3347,N_48213,N_48313);
nor UO_3348 (O_3348,N_47862,N_48118);
or UO_3349 (O_3349,N_48208,N_48564);
nand UO_3350 (O_3350,N_47501,N_48680);
and UO_3351 (O_3351,N_49315,N_47556);
xnor UO_3352 (O_3352,N_49523,N_48451);
and UO_3353 (O_3353,N_48351,N_49096);
and UO_3354 (O_3354,N_49567,N_49593);
xor UO_3355 (O_3355,N_47517,N_48264);
nand UO_3356 (O_3356,N_48834,N_48724);
and UO_3357 (O_3357,N_49302,N_47689);
nand UO_3358 (O_3358,N_48378,N_49270);
xor UO_3359 (O_3359,N_48637,N_48299);
or UO_3360 (O_3360,N_49776,N_48983);
nand UO_3361 (O_3361,N_48151,N_48893);
nor UO_3362 (O_3362,N_49192,N_49277);
nor UO_3363 (O_3363,N_47600,N_48613);
or UO_3364 (O_3364,N_47707,N_48044);
nor UO_3365 (O_3365,N_48323,N_47893);
xnor UO_3366 (O_3366,N_48611,N_49245);
or UO_3367 (O_3367,N_49309,N_48335);
nor UO_3368 (O_3368,N_49129,N_47692);
nand UO_3369 (O_3369,N_48874,N_48071);
and UO_3370 (O_3370,N_48530,N_48570);
or UO_3371 (O_3371,N_49216,N_49800);
nand UO_3372 (O_3372,N_48400,N_49519);
or UO_3373 (O_3373,N_48735,N_48067);
nor UO_3374 (O_3374,N_47570,N_49711);
nand UO_3375 (O_3375,N_47949,N_49522);
nor UO_3376 (O_3376,N_48593,N_48116);
and UO_3377 (O_3377,N_48961,N_48523);
nand UO_3378 (O_3378,N_47673,N_48608);
xor UO_3379 (O_3379,N_49119,N_49171);
nor UO_3380 (O_3380,N_49523,N_49903);
or UO_3381 (O_3381,N_48510,N_48509);
nor UO_3382 (O_3382,N_48723,N_47696);
or UO_3383 (O_3383,N_49960,N_48693);
nor UO_3384 (O_3384,N_49613,N_48381);
xor UO_3385 (O_3385,N_48327,N_49375);
xor UO_3386 (O_3386,N_47570,N_48606);
and UO_3387 (O_3387,N_49073,N_49766);
and UO_3388 (O_3388,N_49878,N_49006);
and UO_3389 (O_3389,N_47926,N_47786);
nor UO_3390 (O_3390,N_49975,N_49456);
nor UO_3391 (O_3391,N_49672,N_49577);
or UO_3392 (O_3392,N_49291,N_48979);
or UO_3393 (O_3393,N_49155,N_48146);
or UO_3394 (O_3394,N_49137,N_47892);
nor UO_3395 (O_3395,N_49220,N_48633);
or UO_3396 (O_3396,N_48400,N_48870);
nor UO_3397 (O_3397,N_47971,N_48927);
nand UO_3398 (O_3398,N_48827,N_47713);
and UO_3399 (O_3399,N_49758,N_48048);
nor UO_3400 (O_3400,N_49701,N_47838);
nor UO_3401 (O_3401,N_49192,N_49339);
or UO_3402 (O_3402,N_49284,N_49182);
and UO_3403 (O_3403,N_47745,N_49436);
nand UO_3404 (O_3404,N_47694,N_48732);
nor UO_3405 (O_3405,N_47662,N_48043);
and UO_3406 (O_3406,N_47941,N_47705);
and UO_3407 (O_3407,N_49949,N_47717);
nand UO_3408 (O_3408,N_47559,N_49584);
nand UO_3409 (O_3409,N_48098,N_48489);
xnor UO_3410 (O_3410,N_48379,N_49462);
xor UO_3411 (O_3411,N_49608,N_49645);
nand UO_3412 (O_3412,N_48875,N_49497);
nand UO_3413 (O_3413,N_47865,N_47698);
or UO_3414 (O_3414,N_49727,N_48615);
and UO_3415 (O_3415,N_48352,N_48281);
and UO_3416 (O_3416,N_47583,N_49985);
and UO_3417 (O_3417,N_48448,N_47726);
or UO_3418 (O_3418,N_48484,N_47502);
nand UO_3419 (O_3419,N_48867,N_48502);
nor UO_3420 (O_3420,N_48128,N_48795);
or UO_3421 (O_3421,N_48404,N_48307);
and UO_3422 (O_3422,N_49629,N_47807);
and UO_3423 (O_3423,N_49117,N_49187);
nor UO_3424 (O_3424,N_49471,N_49426);
nand UO_3425 (O_3425,N_47676,N_48841);
or UO_3426 (O_3426,N_49492,N_49560);
nand UO_3427 (O_3427,N_48193,N_47612);
nand UO_3428 (O_3428,N_48925,N_48976);
nor UO_3429 (O_3429,N_47795,N_47836);
or UO_3430 (O_3430,N_49966,N_47590);
nor UO_3431 (O_3431,N_49939,N_49493);
nand UO_3432 (O_3432,N_49105,N_48305);
nor UO_3433 (O_3433,N_49040,N_49969);
nand UO_3434 (O_3434,N_49049,N_48391);
and UO_3435 (O_3435,N_49433,N_47717);
nor UO_3436 (O_3436,N_49969,N_48381);
and UO_3437 (O_3437,N_47699,N_48772);
nand UO_3438 (O_3438,N_48922,N_48004);
xnor UO_3439 (O_3439,N_49952,N_47788);
nand UO_3440 (O_3440,N_48548,N_49721);
xor UO_3441 (O_3441,N_48102,N_48898);
or UO_3442 (O_3442,N_47829,N_47569);
or UO_3443 (O_3443,N_48043,N_48477);
nor UO_3444 (O_3444,N_48978,N_49910);
and UO_3445 (O_3445,N_49734,N_49934);
or UO_3446 (O_3446,N_48512,N_48390);
nand UO_3447 (O_3447,N_49449,N_47997);
nand UO_3448 (O_3448,N_47874,N_49483);
xnor UO_3449 (O_3449,N_48332,N_49819);
and UO_3450 (O_3450,N_49177,N_49318);
or UO_3451 (O_3451,N_47716,N_49782);
nor UO_3452 (O_3452,N_49683,N_48315);
or UO_3453 (O_3453,N_49333,N_49711);
and UO_3454 (O_3454,N_49451,N_47875);
xor UO_3455 (O_3455,N_47840,N_48781);
or UO_3456 (O_3456,N_48561,N_47752);
nand UO_3457 (O_3457,N_48485,N_49127);
and UO_3458 (O_3458,N_49914,N_47672);
or UO_3459 (O_3459,N_49497,N_49194);
or UO_3460 (O_3460,N_49209,N_47545);
nand UO_3461 (O_3461,N_49107,N_48099);
or UO_3462 (O_3462,N_49359,N_47740);
and UO_3463 (O_3463,N_48056,N_48534);
nor UO_3464 (O_3464,N_49573,N_48448);
nor UO_3465 (O_3465,N_49399,N_49903);
nor UO_3466 (O_3466,N_47817,N_47718);
nand UO_3467 (O_3467,N_48001,N_49281);
nor UO_3468 (O_3468,N_48390,N_48762);
and UO_3469 (O_3469,N_49756,N_49484);
nor UO_3470 (O_3470,N_47987,N_49054);
and UO_3471 (O_3471,N_49110,N_47594);
nand UO_3472 (O_3472,N_48317,N_48445);
xnor UO_3473 (O_3473,N_49855,N_47793);
nand UO_3474 (O_3474,N_48477,N_48355);
nand UO_3475 (O_3475,N_48250,N_48159);
nand UO_3476 (O_3476,N_49857,N_48973);
xnor UO_3477 (O_3477,N_49402,N_48903);
nand UO_3478 (O_3478,N_48566,N_48927);
nand UO_3479 (O_3479,N_49700,N_49177);
nand UO_3480 (O_3480,N_49115,N_48679);
and UO_3481 (O_3481,N_48427,N_49161);
nor UO_3482 (O_3482,N_49805,N_48199);
or UO_3483 (O_3483,N_48134,N_49625);
and UO_3484 (O_3484,N_48661,N_49813);
nand UO_3485 (O_3485,N_49982,N_48057);
nor UO_3486 (O_3486,N_48022,N_49282);
or UO_3487 (O_3487,N_48107,N_47683);
nor UO_3488 (O_3488,N_48304,N_47865);
or UO_3489 (O_3489,N_49501,N_48403);
xnor UO_3490 (O_3490,N_48097,N_49070);
or UO_3491 (O_3491,N_48050,N_47913);
or UO_3492 (O_3492,N_48176,N_48190);
and UO_3493 (O_3493,N_49580,N_48510);
nor UO_3494 (O_3494,N_49297,N_49070);
and UO_3495 (O_3495,N_48893,N_49229);
xnor UO_3496 (O_3496,N_49063,N_48249);
and UO_3497 (O_3497,N_48338,N_49858);
xor UO_3498 (O_3498,N_49687,N_48342);
xnor UO_3499 (O_3499,N_48126,N_48463);
or UO_3500 (O_3500,N_48221,N_49875);
or UO_3501 (O_3501,N_49415,N_48183);
xnor UO_3502 (O_3502,N_48695,N_49164);
and UO_3503 (O_3503,N_49430,N_47815);
nand UO_3504 (O_3504,N_47903,N_49509);
or UO_3505 (O_3505,N_49466,N_47670);
nor UO_3506 (O_3506,N_49650,N_49977);
and UO_3507 (O_3507,N_48286,N_48675);
nor UO_3508 (O_3508,N_48612,N_49918);
and UO_3509 (O_3509,N_47897,N_48223);
nor UO_3510 (O_3510,N_49992,N_49981);
nor UO_3511 (O_3511,N_48969,N_49218);
nand UO_3512 (O_3512,N_47592,N_48375);
or UO_3513 (O_3513,N_47850,N_48144);
xnor UO_3514 (O_3514,N_48682,N_48305);
nand UO_3515 (O_3515,N_49319,N_48404);
or UO_3516 (O_3516,N_49912,N_48276);
or UO_3517 (O_3517,N_48926,N_48678);
or UO_3518 (O_3518,N_48773,N_48792);
nor UO_3519 (O_3519,N_48908,N_48751);
and UO_3520 (O_3520,N_49282,N_48293);
or UO_3521 (O_3521,N_49130,N_49803);
and UO_3522 (O_3522,N_47934,N_49529);
nor UO_3523 (O_3523,N_48808,N_49640);
nor UO_3524 (O_3524,N_48618,N_49547);
and UO_3525 (O_3525,N_47735,N_48505);
or UO_3526 (O_3526,N_48830,N_48855);
or UO_3527 (O_3527,N_49230,N_49312);
nand UO_3528 (O_3528,N_48256,N_49221);
nor UO_3529 (O_3529,N_47921,N_49748);
or UO_3530 (O_3530,N_49200,N_49722);
or UO_3531 (O_3531,N_48103,N_47956);
or UO_3532 (O_3532,N_48784,N_48135);
nor UO_3533 (O_3533,N_47993,N_49523);
nor UO_3534 (O_3534,N_48555,N_49179);
and UO_3535 (O_3535,N_47739,N_49811);
nand UO_3536 (O_3536,N_49142,N_47974);
or UO_3537 (O_3537,N_48362,N_49053);
nand UO_3538 (O_3538,N_47591,N_49320);
nand UO_3539 (O_3539,N_49178,N_48906);
nand UO_3540 (O_3540,N_49690,N_49464);
or UO_3541 (O_3541,N_48688,N_49275);
nand UO_3542 (O_3542,N_47749,N_48254);
nor UO_3543 (O_3543,N_49458,N_47963);
nand UO_3544 (O_3544,N_48341,N_49357);
and UO_3545 (O_3545,N_48489,N_49281);
nor UO_3546 (O_3546,N_48680,N_47870);
xnor UO_3547 (O_3547,N_47521,N_49174);
nor UO_3548 (O_3548,N_47523,N_47818);
nor UO_3549 (O_3549,N_49770,N_47673);
and UO_3550 (O_3550,N_49555,N_48579);
nor UO_3551 (O_3551,N_49441,N_48268);
nand UO_3552 (O_3552,N_48840,N_48947);
or UO_3553 (O_3553,N_47539,N_48160);
xnor UO_3554 (O_3554,N_48274,N_49376);
xor UO_3555 (O_3555,N_48759,N_47856);
nor UO_3556 (O_3556,N_47623,N_48456);
and UO_3557 (O_3557,N_48097,N_49521);
or UO_3558 (O_3558,N_48035,N_48723);
or UO_3559 (O_3559,N_48514,N_48669);
xnor UO_3560 (O_3560,N_47539,N_49890);
and UO_3561 (O_3561,N_47803,N_49889);
nor UO_3562 (O_3562,N_49907,N_49412);
or UO_3563 (O_3563,N_49780,N_49837);
xor UO_3564 (O_3564,N_48140,N_48449);
and UO_3565 (O_3565,N_49345,N_47500);
nand UO_3566 (O_3566,N_48241,N_48877);
or UO_3567 (O_3567,N_48298,N_49151);
nor UO_3568 (O_3568,N_47907,N_49671);
nand UO_3569 (O_3569,N_48576,N_48554);
or UO_3570 (O_3570,N_48582,N_48803);
nand UO_3571 (O_3571,N_49037,N_48311);
or UO_3572 (O_3572,N_48623,N_49996);
and UO_3573 (O_3573,N_49255,N_47545);
nor UO_3574 (O_3574,N_49772,N_48103);
nor UO_3575 (O_3575,N_47695,N_48748);
and UO_3576 (O_3576,N_49589,N_48355);
nand UO_3577 (O_3577,N_48823,N_48658);
nand UO_3578 (O_3578,N_48269,N_48258);
or UO_3579 (O_3579,N_49077,N_48738);
nand UO_3580 (O_3580,N_48245,N_49294);
nor UO_3581 (O_3581,N_47657,N_47587);
and UO_3582 (O_3582,N_49173,N_49229);
nor UO_3583 (O_3583,N_47690,N_48902);
xor UO_3584 (O_3584,N_47869,N_49075);
or UO_3585 (O_3585,N_48723,N_47739);
or UO_3586 (O_3586,N_48936,N_47982);
nor UO_3587 (O_3587,N_48153,N_49073);
nand UO_3588 (O_3588,N_48751,N_49690);
nor UO_3589 (O_3589,N_48546,N_49957);
or UO_3590 (O_3590,N_48385,N_48438);
and UO_3591 (O_3591,N_49570,N_49196);
and UO_3592 (O_3592,N_47978,N_49671);
nand UO_3593 (O_3593,N_48829,N_49059);
nor UO_3594 (O_3594,N_47955,N_49704);
nor UO_3595 (O_3595,N_49694,N_49625);
and UO_3596 (O_3596,N_49271,N_48409);
xnor UO_3597 (O_3597,N_49651,N_47799);
or UO_3598 (O_3598,N_48525,N_48338);
nor UO_3599 (O_3599,N_47903,N_47740);
nor UO_3600 (O_3600,N_48235,N_49952);
nor UO_3601 (O_3601,N_48128,N_49488);
nor UO_3602 (O_3602,N_48687,N_49662);
and UO_3603 (O_3603,N_48646,N_49907);
and UO_3604 (O_3604,N_49714,N_49191);
or UO_3605 (O_3605,N_47865,N_49110);
and UO_3606 (O_3606,N_48270,N_48417);
or UO_3607 (O_3607,N_48884,N_47701);
or UO_3608 (O_3608,N_49545,N_49947);
or UO_3609 (O_3609,N_47678,N_48115);
xnor UO_3610 (O_3610,N_49266,N_49624);
and UO_3611 (O_3611,N_47952,N_49541);
nand UO_3612 (O_3612,N_49917,N_48041);
nor UO_3613 (O_3613,N_49895,N_49738);
nor UO_3614 (O_3614,N_47504,N_47806);
nor UO_3615 (O_3615,N_48050,N_48599);
nand UO_3616 (O_3616,N_48315,N_49199);
nand UO_3617 (O_3617,N_49826,N_49426);
or UO_3618 (O_3618,N_49685,N_49886);
nor UO_3619 (O_3619,N_48894,N_48128);
and UO_3620 (O_3620,N_48868,N_48511);
nor UO_3621 (O_3621,N_49604,N_49573);
nand UO_3622 (O_3622,N_49882,N_49173);
nor UO_3623 (O_3623,N_49961,N_49035);
nand UO_3624 (O_3624,N_48720,N_48164);
nor UO_3625 (O_3625,N_49262,N_47789);
nor UO_3626 (O_3626,N_49150,N_48814);
xnor UO_3627 (O_3627,N_49892,N_47821);
nor UO_3628 (O_3628,N_49424,N_49353);
and UO_3629 (O_3629,N_49947,N_47554);
or UO_3630 (O_3630,N_48531,N_48475);
or UO_3631 (O_3631,N_48785,N_49407);
nor UO_3632 (O_3632,N_47608,N_47649);
nor UO_3633 (O_3633,N_47611,N_49938);
nor UO_3634 (O_3634,N_48742,N_49443);
and UO_3635 (O_3635,N_49966,N_49030);
and UO_3636 (O_3636,N_47950,N_47585);
xor UO_3637 (O_3637,N_48199,N_49125);
nand UO_3638 (O_3638,N_48784,N_49467);
nor UO_3639 (O_3639,N_48251,N_48389);
and UO_3640 (O_3640,N_48328,N_49855);
nand UO_3641 (O_3641,N_49276,N_48811);
nor UO_3642 (O_3642,N_48672,N_48817);
and UO_3643 (O_3643,N_48236,N_49662);
or UO_3644 (O_3644,N_48001,N_48427);
nor UO_3645 (O_3645,N_49312,N_49014);
or UO_3646 (O_3646,N_47503,N_49967);
or UO_3647 (O_3647,N_47520,N_49851);
or UO_3648 (O_3648,N_48745,N_48834);
and UO_3649 (O_3649,N_47794,N_48014);
xnor UO_3650 (O_3650,N_49746,N_48602);
nor UO_3651 (O_3651,N_49831,N_47807);
nand UO_3652 (O_3652,N_48215,N_47952);
or UO_3653 (O_3653,N_48640,N_49674);
nand UO_3654 (O_3654,N_47754,N_47817);
nor UO_3655 (O_3655,N_48812,N_49027);
or UO_3656 (O_3656,N_48242,N_49263);
and UO_3657 (O_3657,N_47561,N_48271);
or UO_3658 (O_3658,N_48474,N_47891);
and UO_3659 (O_3659,N_48259,N_47720);
and UO_3660 (O_3660,N_47834,N_48625);
nor UO_3661 (O_3661,N_47710,N_49968);
or UO_3662 (O_3662,N_48160,N_49425);
or UO_3663 (O_3663,N_49208,N_49284);
nand UO_3664 (O_3664,N_49762,N_48922);
nand UO_3665 (O_3665,N_48336,N_48510);
and UO_3666 (O_3666,N_49823,N_49133);
or UO_3667 (O_3667,N_49339,N_48590);
and UO_3668 (O_3668,N_48355,N_49499);
nor UO_3669 (O_3669,N_49177,N_49952);
and UO_3670 (O_3670,N_49545,N_49103);
nor UO_3671 (O_3671,N_48431,N_47760);
or UO_3672 (O_3672,N_48615,N_48772);
or UO_3673 (O_3673,N_49919,N_47696);
and UO_3674 (O_3674,N_47810,N_48989);
and UO_3675 (O_3675,N_47589,N_48573);
xnor UO_3676 (O_3676,N_48044,N_49240);
nand UO_3677 (O_3677,N_49520,N_48339);
nor UO_3678 (O_3678,N_49790,N_49620);
and UO_3679 (O_3679,N_47799,N_49230);
and UO_3680 (O_3680,N_47615,N_48125);
nand UO_3681 (O_3681,N_47955,N_49356);
nand UO_3682 (O_3682,N_48887,N_47870);
nor UO_3683 (O_3683,N_49107,N_48900);
or UO_3684 (O_3684,N_47814,N_49389);
xor UO_3685 (O_3685,N_49536,N_48277);
nand UO_3686 (O_3686,N_47659,N_48641);
nand UO_3687 (O_3687,N_49269,N_47586);
nor UO_3688 (O_3688,N_48283,N_48165);
nor UO_3689 (O_3689,N_49081,N_49073);
nor UO_3690 (O_3690,N_49564,N_48764);
xnor UO_3691 (O_3691,N_48602,N_49703);
and UO_3692 (O_3692,N_48162,N_47850);
xor UO_3693 (O_3693,N_49457,N_48902);
and UO_3694 (O_3694,N_49227,N_49026);
nand UO_3695 (O_3695,N_47829,N_48550);
and UO_3696 (O_3696,N_48377,N_49215);
or UO_3697 (O_3697,N_47805,N_48788);
nand UO_3698 (O_3698,N_48455,N_49494);
nor UO_3699 (O_3699,N_49268,N_49482);
or UO_3700 (O_3700,N_47843,N_48274);
nor UO_3701 (O_3701,N_48802,N_49048);
nand UO_3702 (O_3702,N_47802,N_49470);
or UO_3703 (O_3703,N_49333,N_48941);
nor UO_3704 (O_3704,N_48455,N_48959);
nand UO_3705 (O_3705,N_48835,N_49333);
or UO_3706 (O_3706,N_47676,N_48289);
or UO_3707 (O_3707,N_48213,N_47846);
nand UO_3708 (O_3708,N_47833,N_48915);
xor UO_3709 (O_3709,N_49467,N_48992);
or UO_3710 (O_3710,N_47900,N_48720);
nor UO_3711 (O_3711,N_48021,N_48889);
and UO_3712 (O_3712,N_47606,N_49225);
and UO_3713 (O_3713,N_49075,N_48607);
or UO_3714 (O_3714,N_47893,N_48804);
nand UO_3715 (O_3715,N_48128,N_48663);
or UO_3716 (O_3716,N_49886,N_49792);
xnor UO_3717 (O_3717,N_48291,N_49400);
nor UO_3718 (O_3718,N_48165,N_49391);
or UO_3719 (O_3719,N_49826,N_47626);
and UO_3720 (O_3720,N_48253,N_47782);
nor UO_3721 (O_3721,N_47693,N_49661);
or UO_3722 (O_3722,N_49082,N_48442);
or UO_3723 (O_3723,N_48562,N_49197);
nand UO_3724 (O_3724,N_48298,N_47950);
or UO_3725 (O_3725,N_48375,N_48051);
or UO_3726 (O_3726,N_47835,N_48481);
nor UO_3727 (O_3727,N_49166,N_48654);
xnor UO_3728 (O_3728,N_47603,N_49742);
nor UO_3729 (O_3729,N_48140,N_48538);
or UO_3730 (O_3730,N_48985,N_48416);
nand UO_3731 (O_3731,N_49712,N_49147);
and UO_3732 (O_3732,N_49026,N_47540);
xnor UO_3733 (O_3733,N_49741,N_47613);
nor UO_3734 (O_3734,N_48731,N_48411);
or UO_3735 (O_3735,N_49605,N_49092);
nor UO_3736 (O_3736,N_48328,N_48155);
xnor UO_3737 (O_3737,N_48147,N_48026);
nor UO_3738 (O_3738,N_49935,N_48542);
and UO_3739 (O_3739,N_49560,N_48416);
xor UO_3740 (O_3740,N_49598,N_49789);
nand UO_3741 (O_3741,N_48748,N_49386);
and UO_3742 (O_3742,N_49157,N_48589);
nand UO_3743 (O_3743,N_48413,N_48589);
xor UO_3744 (O_3744,N_48360,N_48373);
or UO_3745 (O_3745,N_48676,N_47666);
and UO_3746 (O_3746,N_47616,N_47921);
nand UO_3747 (O_3747,N_48034,N_49300);
and UO_3748 (O_3748,N_47774,N_47712);
nor UO_3749 (O_3749,N_47983,N_48566);
and UO_3750 (O_3750,N_47840,N_49149);
nor UO_3751 (O_3751,N_47764,N_47857);
and UO_3752 (O_3752,N_48664,N_48030);
or UO_3753 (O_3753,N_49666,N_49746);
and UO_3754 (O_3754,N_48719,N_48638);
and UO_3755 (O_3755,N_47544,N_48916);
nor UO_3756 (O_3756,N_48509,N_47835);
and UO_3757 (O_3757,N_49784,N_49034);
nand UO_3758 (O_3758,N_48276,N_49058);
nand UO_3759 (O_3759,N_47746,N_47854);
xnor UO_3760 (O_3760,N_48065,N_49753);
or UO_3761 (O_3761,N_49970,N_48743);
nor UO_3762 (O_3762,N_49194,N_48808);
nand UO_3763 (O_3763,N_48905,N_48224);
nand UO_3764 (O_3764,N_49401,N_47559);
and UO_3765 (O_3765,N_48459,N_49747);
or UO_3766 (O_3766,N_49456,N_48484);
and UO_3767 (O_3767,N_48066,N_48194);
nor UO_3768 (O_3768,N_48727,N_48593);
and UO_3769 (O_3769,N_48925,N_48859);
nor UO_3770 (O_3770,N_47880,N_48734);
nand UO_3771 (O_3771,N_49643,N_48826);
or UO_3772 (O_3772,N_48533,N_48744);
or UO_3773 (O_3773,N_48541,N_49095);
nor UO_3774 (O_3774,N_49073,N_48505);
or UO_3775 (O_3775,N_47892,N_49392);
nor UO_3776 (O_3776,N_49011,N_48305);
nand UO_3777 (O_3777,N_49595,N_47957);
nor UO_3778 (O_3778,N_48880,N_49522);
or UO_3779 (O_3779,N_49115,N_49272);
and UO_3780 (O_3780,N_48975,N_49240);
nand UO_3781 (O_3781,N_49181,N_48183);
nor UO_3782 (O_3782,N_49152,N_49271);
nand UO_3783 (O_3783,N_49714,N_48738);
nor UO_3784 (O_3784,N_49220,N_48600);
and UO_3785 (O_3785,N_48970,N_48563);
nor UO_3786 (O_3786,N_48555,N_49318);
and UO_3787 (O_3787,N_48384,N_49952);
nand UO_3788 (O_3788,N_48431,N_47556);
xnor UO_3789 (O_3789,N_49961,N_48362);
nor UO_3790 (O_3790,N_49390,N_49768);
nor UO_3791 (O_3791,N_49362,N_48423);
and UO_3792 (O_3792,N_48542,N_47676);
xnor UO_3793 (O_3793,N_49558,N_49771);
and UO_3794 (O_3794,N_48503,N_48782);
nor UO_3795 (O_3795,N_47618,N_48490);
nor UO_3796 (O_3796,N_48730,N_49712);
and UO_3797 (O_3797,N_48771,N_49516);
nor UO_3798 (O_3798,N_48437,N_48095);
or UO_3799 (O_3799,N_49464,N_47547);
and UO_3800 (O_3800,N_49284,N_49976);
and UO_3801 (O_3801,N_49820,N_48262);
and UO_3802 (O_3802,N_49029,N_47692);
nand UO_3803 (O_3803,N_48029,N_49733);
nand UO_3804 (O_3804,N_49338,N_49360);
and UO_3805 (O_3805,N_49258,N_49369);
nor UO_3806 (O_3806,N_47729,N_49040);
or UO_3807 (O_3807,N_47597,N_47982);
xnor UO_3808 (O_3808,N_49955,N_48099);
xnor UO_3809 (O_3809,N_48521,N_48275);
and UO_3810 (O_3810,N_48942,N_47734);
and UO_3811 (O_3811,N_47833,N_49514);
or UO_3812 (O_3812,N_48383,N_48432);
and UO_3813 (O_3813,N_49956,N_48940);
and UO_3814 (O_3814,N_49615,N_48232);
nor UO_3815 (O_3815,N_49635,N_49702);
nand UO_3816 (O_3816,N_49380,N_49286);
and UO_3817 (O_3817,N_49296,N_49697);
xor UO_3818 (O_3818,N_49730,N_47782);
or UO_3819 (O_3819,N_48356,N_49930);
nor UO_3820 (O_3820,N_47668,N_48081);
and UO_3821 (O_3821,N_48209,N_49461);
and UO_3822 (O_3822,N_48613,N_49226);
and UO_3823 (O_3823,N_48331,N_48151);
and UO_3824 (O_3824,N_48272,N_48240);
nand UO_3825 (O_3825,N_47562,N_47625);
nand UO_3826 (O_3826,N_47569,N_49944);
or UO_3827 (O_3827,N_48800,N_48369);
nor UO_3828 (O_3828,N_49557,N_49823);
or UO_3829 (O_3829,N_48198,N_48851);
nand UO_3830 (O_3830,N_47568,N_49534);
nor UO_3831 (O_3831,N_47721,N_48691);
nor UO_3832 (O_3832,N_49185,N_47529);
nor UO_3833 (O_3833,N_48435,N_48226);
or UO_3834 (O_3834,N_49611,N_49340);
xor UO_3835 (O_3835,N_48076,N_48036);
and UO_3836 (O_3836,N_47836,N_48374);
or UO_3837 (O_3837,N_49437,N_49349);
nand UO_3838 (O_3838,N_49159,N_49727);
xor UO_3839 (O_3839,N_49718,N_48130);
or UO_3840 (O_3840,N_48650,N_47788);
nor UO_3841 (O_3841,N_49516,N_48331);
and UO_3842 (O_3842,N_48183,N_47844);
or UO_3843 (O_3843,N_48214,N_49481);
nor UO_3844 (O_3844,N_49748,N_48069);
or UO_3845 (O_3845,N_49077,N_49942);
and UO_3846 (O_3846,N_47894,N_48744);
nand UO_3847 (O_3847,N_48909,N_47961);
or UO_3848 (O_3848,N_49485,N_49596);
xor UO_3849 (O_3849,N_49409,N_49622);
or UO_3850 (O_3850,N_48065,N_49264);
and UO_3851 (O_3851,N_47964,N_48211);
and UO_3852 (O_3852,N_49748,N_49581);
or UO_3853 (O_3853,N_49171,N_49131);
nor UO_3854 (O_3854,N_48554,N_48003);
or UO_3855 (O_3855,N_48980,N_49862);
xnor UO_3856 (O_3856,N_48786,N_48447);
nand UO_3857 (O_3857,N_48922,N_48852);
and UO_3858 (O_3858,N_48805,N_48047);
nor UO_3859 (O_3859,N_49905,N_48735);
nand UO_3860 (O_3860,N_48097,N_49714);
nor UO_3861 (O_3861,N_49503,N_49822);
nor UO_3862 (O_3862,N_49130,N_49932);
and UO_3863 (O_3863,N_48033,N_48592);
nand UO_3864 (O_3864,N_48419,N_49549);
or UO_3865 (O_3865,N_48472,N_48330);
nor UO_3866 (O_3866,N_48762,N_47766);
and UO_3867 (O_3867,N_49800,N_49132);
and UO_3868 (O_3868,N_48585,N_48749);
nor UO_3869 (O_3869,N_48555,N_47737);
nand UO_3870 (O_3870,N_49438,N_48559);
nor UO_3871 (O_3871,N_47641,N_48280);
or UO_3872 (O_3872,N_48062,N_49210);
nand UO_3873 (O_3873,N_47958,N_48781);
xor UO_3874 (O_3874,N_49268,N_48487);
xnor UO_3875 (O_3875,N_47759,N_47614);
or UO_3876 (O_3876,N_48098,N_49267);
and UO_3877 (O_3877,N_48627,N_49065);
or UO_3878 (O_3878,N_48009,N_48992);
nand UO_3879 (O_3879,N_49104,N_49773);
nand UO_3880 (O_3880,N_49470,N_48356);
nor UO_3881 (O_3881,N_48256,N_49555);
nor UO_3882 (O_3882,N_48373,N_47912);
nor UO_3883 (O_3883,N_49544,N_49260);
and UO_3884 (O_3884,N_47997,N_49675);
or UO_3885 (O_3885,N_48046,N_49815);
nand UO_3886 (O_3886,N_48201,N_47529);
nor UO_3887 (O_3887,N_47877,N_48430);
nand UO_3888 (O_3888,N_48050,N_49873);
nor UO_3889 (O_3889,N_48989,N_47942);
nand UO_3890 (O_3890,N_49449,N_49683);
nor UO_3891 (O_3891,N_48739,N_48673);
nor UO_3892 (O_3892,N_47784,N_48279);
nor UO_3893 (O_3893,N_48516,N_49521);
or UO_3894 (O_3894,N_49884,N_49809);
nor UO_3895 (O_3895,N_48455,N_49745);
or UO_3896 (O_3896,N_48061,N_47665);
or UO_3897 (O_3897,N_47750,N_49761);
nor UO_3898 (O_3898,N_48645,N_48687);
nor UO_3899 (O_3899,N_47979,N_48325);
nand UO_3900 (O_3900,N_48626,N_49638);
or UO_3901 (O_3901,N_48648,N_49145);
nand UO_3902 (O_3902,N_48377,N_49142);
xor UO_3903 (O_3903,N_48710,N_48134);
and UO_3904 (O_3904,N_48360,N_49042);
or UO_3905 (O_3905,N_49052,N_47500);
and UO_3906 (O_3906,N_48170,N_49057);
nand UO_3907 (O_3907,N_47948,N_48354);
nand UO_3908 (O_3908,N_48137,N_48099);
nand UO_3909 (O_3909,N_49081,N_49545);
nand UO_3910 (O_3910,N_48389,N_49129);
nor UO_3911 (O_3911,N_49030,N_48059);
and UO_3912 (O_3912,N_48457,N_49130);
nor UO_3913 (O_3913,N_48801,N_47961);
nand UO_3914 (O_3914,N_49725,N_48869);
and UO_3915 (O_3915,N_48925,N_49898);
nand UO_3916 (O_3916,N_49897,N_49838);
and UO_3917 (O_3917,N_49686,N_47640);
nor UO_3918 (O_3918,N_49954,N_48700);
xnor UO_3919 (O_3919,N_48350,N_48440);
xnor UO_3920 (O_3920,N_48077,N_49821);
and UO_3921 (O_3921,N_49443,N_48179);
and UO_3922 (O_3922,N_48306,N_49122);
or UO_3923 (O_3923,N_47897,N_49838);
and UO_3924 (O_3924,N_47974,N_47933);
nand UO_3925 (O_3925,N_47547,N_48923);
nand UO_3926 (O_3926,N_48335,N_49683);
xnor UO_3927 (O_3927,N_49728,N_48851);
and UO_3928 (O_3928,N_49051,N_48958);
and UO_3929 (O_3929,N_48104,N_49959);
or UO_3930 (O_3930,N_49645,N_48209);
nand UO_3931 (O_3931,N_49959,N_49062);
and UO_3932 (O_3932,N_48025,N_49888);
xnor UO_3933 (O_3933,N_47874,N_49163);
and UO_3934 (O_3934,N_49129,N_47736);
or UO_3935 (O_3935,N_49817,N_48212);
and UO_3936 (O_3936,N_48518,N_47688);
nor UO_3937 (O_3937,N_47860,N_49630);
and UO_3938 (O_3938,N_49911,N_49866);
and UO_3939 (O_3939,N_49852,N_47544);
nand UO_3940 (O_3940,N_48346,N_48105);
and UO_3941 (O_3941,N_48979,N_47741);
and UO_3942 (O_3942,N_47635,N_49352);
and UO_3943 (O_3943,N_48091,N_49856);
and UO_3944 (O_3944,N_48797,N_49385);
and UO_3945 (O_3945,N_48311,N_49831);
xor UO_3946 (O_3946,N_49773,N_48472);
nor UO_3947 (O_3947,N_49454,N_48432);
nor UO_3948 (O_3948,N_48609,N_48513);
or UO_3949 (O_3949,N_48500,N_48496);
nand UO_3950 (O_3950,N_48051,N_47940);
nand UO_3951 (O_3951,N_47659,N_49318);
nor UO_3952 (O_3952,N_49465,N_48530);
nand UO_3953 (O_3953,N_47934,N_49074);
and UO_3954 (O_3954,N_49415,N_48799);
nand UO_3955 (O_3955,N_48968,N_49330);
nand UO_3956 (O_3956,N_47795,N_49417);
or UO_3957 (O_3957,N_48518,N_49545);
nand UO_3958 (O_3958,N_47964,N_48011);
or UO_3959 (O_3959,N_49157,N_49059);
xor UO_3960 (O_3960,N_49424,N_49560);
and UO_3961 (O_3961,N_49354,N_49944);
nand UO_3962 (O_3962,N_49749,N_49189);
nand UO_3963 (O_3963,N_49337,N_48184);
xnor UO_3964 (O_3964,N_47704,N_48672);
or UO_3965 (O_3965,N_49572,N_48929);
nand UO_3966 (O_3966,N_48526,N_48677);
nor UO_3967 (O_3967,N_49553,N_49132);
nand UO_3968 (O_3968,N_48483,N_48533);
and UO_3969 (O_3969,N_47607,N_49617);
nor UO_3970 (O_3970,N_49089,N_49515);
nand UO_3971 (O_3971,N_48065,N_49727);
nor UO_3972 (O_3972,N_49725,N_49702);
nor UO_3973 (O_3973,N_48972,N_48474);
nor UO_3974 (O_3974,N_47776,N_48774);
nor UO_3975 (O_3975,N_49844,N_47902);
nand UO_3976 (O_3976,N_49832,N_48794);
and UO_3977 (O_3977,N_49861,N_49780);
nor UO_3978 (O_3978,N_49754,N_47570);
xor UO_3979 (O_3979,N_47779,N_49321);
nor UO_3980 (O_3980,N_49306,N_48560);
or UO_3981 (O_3981,N_49839,N_48650);
nand UO_3982 (O_3982,N_47664,N_49630);
nand UO_3983 (O_3983,N_47809,N_49448);
nor UO_3984 (O_3984,N_49036,N_48068);
and UO_3985 (O_3985,N_48972,N_48467);
or UO_3986 (O_3986,N_47947,N_47553);
and UO_3987 (O_3987,N_48825,N_47759);
nand UO_3988 (O_3988,N_49611,N_48942);
and UO_3989 (O_3989,N_49775,N_47789);
xnor UO_3990 (O_3990,N_49863,N_49153);
or UO_3991 (O_3991,N_49510,N_48960);
xnor UO_3992 (O_3992,N_49548,N_49906);
nand UO_3993 (O_3993,N_49541,N_49167);
nand UO_3994 (O_3994,N_48845,N_47608);
xor UO_3995 (O_3995,N_49212,N_48814);
xnor UO_3996 (O_3996,N_48574,N_47957);
or UO_3997 (O_3997,N_49877,N_48033);
nor UO_3998 (O_3998,N_48044,N_48137);
nor UO_3999 (O_3999,N_49411,N_48350);
nand UO_4000 (O_4000,N_48513,N_49497);
nor UO_4001 (O_4001,N_48081,N_49548);
nand UO_4002 (O_4002,N_49388,N_48514);
or UO_4003 (O_4003,N_48388,N_49418);
and UO_4004 (O_4004,N_47975,N_49581);
or UO_4005 (O_4005,N_48669,N_47562);
nor UO_4006 (O_4006,N_48642,N_48419);
and UO_4007 (O_4007,N_48464,N_48066);
nand UO_4008 (O_4008,N_48562,N_48560);
or UO_4009 (O_4009,N_48241,N_47900);
nand UO_4010 (O_4010,N_49345,N_48662);
or UO_4011 (O_4011,N_47721,N_47744);
xnor UO_4012 (O_4012,N_48657,N_48302);
nor UO_4013 (O_4013,N_47811,N_49783);
or UO_4014 (O_4014,N_47520,N_48046);
nor UO_4015 (O_4015,N_48781,N_47938);
xor UO_4016 (O_4016,N_48848,N_49411);
nand UO_4017 (O_4017,N_49300,N_47794);
nor UO_4018 (O_4018,N_49396,N_49369);
nand UO_4019 (O_4019,N_49430,N_49947);
nor UO_4020 (O_4020,N_49959,N_47909);
nand UO_4021 (O_4021,N_49871,N_47764);
nor UO_4022 (O_4022,N_48252,N_48106);
and UO_4023 (O_4023,N_49312,N_49032);
nor UO_4024 (O_4024,N_49098,N_48307);
nor UO_4025 (O_4025,N_48783,N_49906);
nand UO_4026 (O_4026,N_48565,N_49255);
nor UO_4027 (O_4027,N_49304,N_48413);
nor UO_4028 (O_4028,N_49514,N_49316);
and UO_4029 (O_4029,N_47767,N_49407);
nor UO_4030 (O_4030,N_47864,N_49892);
nor UO_4031 (O_4031,N_49648,N_49246);
nand UO_4032 (O_4032,N_49785,N_47561);
nand UO_4033 (O_4033,N_48271,N_47551);
xnor UO_4034 (O_4034,N_47732,N_48928);
or UO_4035 (O_4035,N_48711,N_48182);
and UO_4036 (O_4036,N_47989,N_49145);
xor UO_4037 (O_4037,N_49546,N_48280);
and UO_4038 (O_4038,N_47541,N_49023);
and UO_4039 (O_4039,N_49330,N_48582);
or UO_4040 (O_4040,N_49202,N_48965);
or UO_4041 (O_4041,N_48635,N_47561);
and UO_4042 (O_4042,N_47918,N_48180);
nor UO_4043 (O_4043,N_49635,N_47551);
xor UO_4044 (O_4044,N_48479,N_49757);
nor UO_4045 (O_4045,N_48352,N_49162);
nand UO_4046 (O_4046,N_49875,N_48205);
nand UO_4047 (O_4047,N_48534,N_49659);
and UO_4048 (O_4048,N_49013,N_49287);
and UO_4049 (O_4049,N_48505,N_48579);
nand UO_4050 (O_4050,N_49720,N_49443);
nand UO_4051 (O_4051,N_48912,N_48237);
and UO_4052 (O_4052,N_48315,N_49447);
nand UO_4053 (O_4053,N_47745,N_49298);
and UO_4054 (O_4054,N_48924,N_49859);
nor UO_4055 (O_4055,N_48659,N_48938);
or UO_4056 (O_4056,N_48588,N_47882);
nor UO_4057 (O_4057,N_49710,N_47826);
or UO_4058 (O_4058,N_48482,N_47554);
nor UO_4059 (O_4059,N_49220,N_49565);
nand UO_4060 (O_4060,N_48729,N_48618);
or UO_4061 (O_4061,N_48811,N_49032);
xor UO_4062 (O_4062,N_48617,N_49374);
and UO_4063 (O_4063,N_47945,N_48695);
and UO_4064 (O_4064,N_49764,N_47924);
xor UO_4065 (O_4065,N_49640,N_49752);
nand UO_4066 (O_4066,N_48952,N_49905);
and UO_4067 (O_4067,N_49818,N_48140);
nand UO_4068 (O_4068,N_48943,N_47933);
and UO_4069 (O_4069,N_48149,N_47716);
nand UO_4070 (O_4070,N_47815,N_49163);
nand UO_4071 (O_4071,N_48469,N_49434);
or UO_4072 (O_4072,N_48437,N_49745);
and UO_4073 (O_4073,N_49493,N_49047);
or UO_4074 (O_4074,N_49452,N_47503);
or UO_4075 (O_4075,N_48159,N_48642);
nand UO_4076 (O_4076,N_48029,N_49967);
nor UO_4077 (O_4077,N_49051,N_49494);
and UO_4078 (O_4078,N_49463,N_48438);
or UO_4079 (O_4079,N_48308,N_48136);
nand UO_4080 (O_4080,N_47829,N_48761);
xnor UO_4081 (O_4081,N_47668,N_49037);
nor UO_4082 (O_4082,N_49925,N_48003);
nor UO_4083 (O_4083,N_47869,N_49103);
and UO_4084 (O_4084,N_48110,N_49223);
nand UO_4085 (O_4085,N_49489,N_49820);
nor UO_4086 (O_4086,N_49494,N_49982);
and UO_4087 (O_4087,N_49979,N_49525);
nand UO_4088 (O_4088,N_49203,N_48548);
nand UO_4089 (O_4089,N_49731,N_49199);
and UO_4090 (O_4090,N_49344,N_47743);
nor UO_4091 (O_4091,N_49866,N_49969);
or UO_4092 (O_4092,N_49330,N_49018);
nor UO_4093 (O_4093,N_47914,N_48554);
nor UO_4094 (O_4094,N_47563,N_49978);
and UO_4095 (O_4095,N_49981,N_49914);
and UO_4096 (O_4096,N_47893,N_49626);
nand UO_4097 (O_4097,N_47717,N_49454);
nor UO_4098 (O_4098,N_47901,N_47924);
or UO_4099 (O_4099,N_48158,N_47995);
nor UO_4100 (O_4100,N_49604,N_49825);
nand UO_4101 (O_4101,N_48888,N_47609);
nand UO_4102 (O_4102,N_49350,N_48721);
nand UO_4103 (O_4103,N_48127,N_49298);
and UO_4104 (O_4104,N_47662,N_48305);
and UO_4105 (O_4105,N_49876,N_49715);
or UO_4106 (O_4106,N_48480,N_49925);
or UO_4107 (O_4107,N_49700,N_47851);
or UO_4108 (O_4108,N_49860,N_48160);
or UO_4109 (O_4109,N_49930,N_47722);
nand UO_4110 (O_4110,N_48206,N_48574);
nand UO_4111 (O_4111,N_48318,N_48835);
and UO_4112 (O_4112,N_47508,N_49652);
nor UO_4113 (O_4113,N_49115,N_47825);
and UO_4114 (O_4114,N_48509,N_48392);
nor UO_4115 (O_4115,N_49118,N_48078);
and UO_4116 (O_4116,N_49677,N_48845);
or UO_4117 (O_4117,N_49499,N_48830);
xnor UO_4118 (O_4118,N_49081,N_48044);
or UO_4119 (O_4119,N_49392,N_48417);
and UO_4120 (O_4120,N_48620,N_48075);
nand UO_4121 (O_4121,N_49878,N_48836);
and UO_4122 (O_4122,N_49338,N_47695);
xnor UO_4123 (O_4123,N_48287,N_49918);
and UO_4124 (O_4124,N_49840,N_48178);
or UO_4125 (O_4125,N_48201,N_49409);
xnor UO_4126 (O_4126,N_47572,N_48913);
and UO_4127 (O_4127,N_49516,N_49471);
or UO_4128 (O_4128,N_48026,N_47877);
and UO_4129 (O_4129,N_47577,N_49197);
nand UO_4130 (O_4130,N_49425,N_48595);
nor UO_4131 (O_4131,N_49667,N_49943);
nand UO_4132 (O_4132,N_49586,N_49130);
nor UO_4133 (O_4133,N_49212,N_49249);
nor UO_4134 (O_4134,N_49231,N_48581);
and UO_4135 (O_4135,N_49686,N_47736);
and UO_4136 (O_4136,N_48062,N_49984);
nor UO_4137 (O_4137,N_49090,N_49843);
and UO_4138 (O_4138,N_49123,N_48926);
or UO_4139 (O_4139,N_47913,N_49955);
xor UO_4140 (O_4140,N_49352,N_47956);
or UO_4141 (O_4141,N_48790,N_48580);
nand UO_4142 (O_4142,N_48761,N_47755);
or UO_4143 (O_4143,N_49318,N_49964);
xor UO_4144 (O_4144,N_49073,N_49692);
xnor UO_4145 (O_4145,N_49153,N_49536);
nor UO_4146 (O_4146,N_49033,N_48104);
and UO_4147 (O_4147,N_49878,N_48530);
and UO_4148 (O_4148,N_49789,N_48458);
nor UO_4149 (O_4149,N_49567,N_49166);
nand UO_4150 (O_4150,N_49811,N_49411);
nand UO_4151 (O_4151,N_49789,N_49800);
and UO_4152 (O_4152,N_48104,N_48189);
nor UO_4153 (O_4153,N_47968,N_48236);
and UO_4154 (O_4154,N_47933,N_47707);
nor UO_4155 (O_4155,N_48908,N_49127);
nand UO_4156 (O_4156,N_48752,N_48682);
nand UO_4157 (O_4157,N_47985,N_49363);
or UO_4158 (O_4158,N_49530,N_48225);
or UO_4159 (O_4159,N_48048,N_48523);
nand UO_4160 (O_4160,N_48728,N_49394);
and UO_4161 (O_4161,N_49183,N_48181);
xor UO_4162 (O_4162,N_49615,N_48436);
and UO_4163 (O_4163,N_49048,N_47604);
or UO_4164 (O_4164,N_48009,N_49442);
nand UO_4165 (O_4165,N_49941,N_47911);
nor UO_4166 (O_4166,N_48233,N_47852);
and UO_4167 (O_4167,N_49093,N_47608);
nor UO_4168 (O_4168,N_48678,N_48560);
or UO_4169 (O_4169,N_47725,N_48842);
nor UO_4170 (O_4170,N_48963,N_49666);
nand UO_4171 (O_4171,N_49857,N_47752);
and UO_4172 (O_4172,N_47971,N_48974);
and UO_4173 (O_4173,N_49887,N_48835);
nor UO_4174 (O_4174,N_48126,N_49942);
or UO_4175 (O_4175,N_49699,N_49796);
or UO_4176 (O_4176,N_48382,N_47710);
nor UO_4177 (O_4177,N_48210,N_49980);
or UO_4178 (O_4178,N_49861,N_49640);
nand UO_4179 (O_4179,N_47772,N_47522);
nor UO_4180 (O_4180,N_47820,N_47966);
nand UO_4181 (O_4181,N_49502,N_47801);
or UO_4182 (O_4182,N_49455,N_48378);
nor UO_4183 (O_4183,N_49218,N_49919);
nand UO_4184 (O_4184,N_48308,N_49191);
nand UO_4185 (O_4185,N_49333,N_47712);
nor UO_4186 (O_4186,N_47509,N_48312);
nand UO_4187 (O_4187,N_49381,N_49954);
and UO_4188 (O_4188,N_47604,N_49255);
nand UO_4189 (O_4189,N_49805,N_48794);
nor UO_4190 (O_4190,N_49462,N_47990);
and UO_4191 (O_4191,N_48209,N_47554);
or UO_4192 (O_4192,N_47877,N_49230);
or UO_4193 (O_4193,N_49174,N_48211);
nor UO_4194 (O_4194,N_49891,N_49521);
nor UO_4195 (O_4195,N_47923,N_49599);
and UO_4196 (O_4196,N_47752,N_47935);
or UO_4197 (O_4197,N_48330,N_48377);
nor UO_4198 (O_4198,N_48641,N_49919);
and UO_4199 (O_4199,N_48103,N_48290);
xor UO_4200 (O_4200,N_49262,N_48647);
nand UO_4201 (O_4201,N_48376,N_48201);
nand UO_4202 (O_4202,N_49529,N_48710);
nand UO_4203 (O_4203,N_48762,N_47596);
nor UO_4204 (O_4204,N_47948,N_48876);
or UO_4205 (O_4205,N_47711,N_48177);
nand UO_4206 (O_4206,N_48771,N_49639);
xnor UO_4207 (O_4207,N_49279,N_49154);
nand UO_4208 (O_4208,N_48625,N_49999);
or UO_4209 (O_4209,N_49929,N_49369);
and UO_4210 (O_4210,N_49666,N_48739);
nand UO_4211 (O_4211,N_48434,N_48780);
nor UO_4212 (O_4212,N_49729,N_48612);
xnor UO_4213 (O_4213,N_49239,N_48002);
nand UO_4214 (O_4214,N_49298,N_47752);
and UO_4215 (O_4215,N_48068,N_48341);
nand UO_4216 (O_4216,N_48657,N_49552);
and UO_4217 (O_4217,N_49163,N_47980);
and UO_4218 (O_4218,N_49752,N_48424);
or UO_4219 (O_4219,N_47806,N_47629);
and UO_4220 (O_4220,N_48742,N_49941);
nor UO_4221 (O_4221,N_48865,N_47834);
nand UO_4222 (O_4222,N_47834,N_48245);
nand UO_4223 (O_4223,N_49929,N_48808);
or UO_4224 (O_4224,N_47970,N_49345);
nor UO_4225 (O_4225,N_48450,N_48677);
nor UO_4226 (O_4226,N_47686,N_49179);
or UO_4227 (O_4227,N_48025,N_49538);
nor UO_4228 (O_4228,N_48744,N_49783);
nor UO_4229 (O_4229,N_48664,N_48502);
and UO_4230 (O_4230,N_49106,N_49615);
or UO_4231 (O_4231,N_48292,N_49954);
or UO_4232 (O_4232,N_49456,N_49311);
or UO_4233 (O_4233,N_47696,N_49021);
or UO_4234 (O_4234,N_49047,N_49693);
nor UO_4235 (O_4235,N_47583,N_49627);
xor UO_4236 (O_4236,N_47704,N_48857);
or UO_4237 (O_4237,N_48300,N_48849);
or UO_4238 (O_4238,N_48714,N_49193);
and UO_4239 (O_4239,N_49202,N_47627);
and UO_4240 (O_4240,N_48510,N_48148);
or UO_4241 (O_4241,N_49504,N_49830);
or UO_4242 (O_4242,N_49562,N_49966);
nand UO_4243 (O_4243,N_48250,N_49697);
or UO_4244 (O_4244,N_49780,N_49479);
or UO_4245 (O_4245,N_47761,N_48544);
nand UO_4246 (O_4246,N_48872,N_47576);
or UO_4247 (O_4247,N_49196,N_47604);
or UO_4248 (O_4248,N_49304,N_49415);
or UO_4249 (O_4249,N_49954,N_48745);
nand UO_4250 (O_4250,N_47742,N_49688);
nand UO_4251 (O_4251,N_49635,N_49311);
xnor UO_4252 (O_4252,N_48429,N_47763);
nor UO_4253 (O_4253,N_48035,N_48125);
or UO_4254 (O_4254,N_48818,N_48291);
or UO_4255 (O_4255,N_47922,N_48902);
nor UO_4256 (O_4256,N_47669,N_47621);
and UO_4257 (O_4257,N_49938,N_48636);
nor UO_4258 (O_4258,N_47943,N_47684);
nand UO_4259 (O_4259,N_47761,N_48268);
xor UO_4260 (O_4260,N_47725,N_47850);
and UO_4261 (O_4261,N_49004,N_49804);
and UO_4262 (O_4262,N_48043,N_47646);
nand UO_4263 (O_4263,N_47982,N_49072);
or UO_4264 (O_4264,N_48162,N_48968);
nor UO_4265 (O_4265,N_48444,N_48804);
xor UO_4266 (O_4266,N_49968,N_47638);
and UO_4267 (O_4267,N_49934,N_48801);
nand UO_4268 (O_4268,N_47984,N_49488);
or UO_4269 (O_4269,N_48679,N_48962);
nand UO_4270 (O_4270,N_48934,N_47947);
or UO_4271 (O_4271,N_48695,N_47984);
nand UO_4272 (O_4272,N_48091,N_47589);
nand UO_4273 (O_4273,N_49457,N_49289);
or UO_4274 (O_4274,N_49746,N_47998);
nand UO_4275 (O_4275,N_49343,N_49620);
or UO_4276 (O_4276,N_48277,N_49381);
and UO_4277 (O_4277,N_49915,N_48583);
xnor UO_4278 (O_4278,N_48786,N_49288);
nand UO_4279 (O_4279,N_49011,N_48784);
nand UO_4280 (O_4280,N_49900,N_48004);
and UO_4281 (O_4281,N_48737,N_48649);
nand UO_4282 (O_4282,N_48614,N_48214);
nor UO_4283 (O_4283,N_49915,N_48584);
nor UO_4284 (O_4284,N_47525,N_47764);
nor UO_4285 (O_4285,N_48120,N_49666);
nor UO_4286 (O_4286,N_49906,N_49209);
and UO_4287 (O_4287,N_47864,N_48017);
or UO_4288 (O_4288,N_47981,N_47830);
nand UO_4289 (O_4289,N_49172,N_49836);
nand UO_4290 (O_4290,N_48739,N_48218);
or UO_4291 (O_4291,N_48043,N_49952);
or UO_4292 (O_4292,N_48771,N_49775);
xor UO_4293 (O_4293,N_48104,N_49039);
nor UO_4294 (O_4294,N_48513,N_48747);
nand UO_4295 (O_4295,N_49700,N_49927);
nand UO_4296 (O_4296,N_49223,N_48195);
nor UO_4297 (O_4297,N_49189,N_48319);
nand UO_4298 (O_4298,N_49902,N_49816);
and UO_4299 (O_4299,N_47692,N_48696);
or UO_4300 (O_4300,N_48982,N_47613);
and UO_4301 (O_4301,N_48446,N_49392);
and UO_4302 (O_4302,N_49033,N_47780);
xor UO_4303 (O_4303,N_49891,N_49404);
nand UO_4304 (O_4304,N_49959,N_48905);
and UO_4305 (O_4305,N_49548,N_49712);
or UO_4306 (O_4306,N_49797,N_49787);
xor UO_4307 (O_4307,N_48209,N_47719);
nor UO_4308 (O_4308,N_48120,N_47658);
or UO_4309 (O_4309,N_48655,N_48565);
and UO_4310 (O_4310,N_48929,N_49329);
nor UO_4311 (O_4311,N_48807,N_49597);
nor UO_4312 (O_4312,N_48045,N_48028);
nor UO_4313 (O_4313,N_48758,N_49261);
and UO_4314 (O_4314,N_49790,N_49464);
nand UO_4315 (O_4315,N_49425,N_48055);
nand UO_4316 (O_4316,N_47612,N_48699);
and UO_4317 (O_4317,N_47579,N_49535);
xor UO_4318 (O_4318,N_49906,N_48794);
nand UO_4319 (O_4319,N_47756,N_49191);
nor UO_4320 (O_4320,N_47755,N_48881);
nand UO_4321 (O_4321,N_49028,N_49862);
or UO_4322 (O_4322,N_48313,N_47721);
and UO_4323 (O_4323,N_48419,N_48170);
nor UO_4324 (O_4324,N_48733,N_47799);
nand UO_4325 (O_4325,N_48350,N_48467);
nor UO_4326 (O_4326,N_48887,N_48382);
nand UO_4327 (O_4327,N_49372,N_47754);
nor UO_4328 (O_4328,N_48920,N_48121);
or UO_4329 (O_4329,N_48988,N_49775);
and UO_4330 (O_4330,N_49634,N_49922);
xor UO_4331 (O_4331,N_49609,N_49378);
or UO_4332 (O_4332,N_49189,N_49747);
xor UO_4333 (O_4333,N_49775,N_49234);
nand UO_4334 (O_4334,N_49747,N_49179);
nor UO_4335 (O_4335,N_48564,N_49450);
nor UO_4336 (O_4336,N_49438,N_49684);
nand UO_4337 (O_4337,N_48526,N_47743);
nor UO_4338 (O_4338,N_47542,N_48979);
or UO_4339 (O_4339,N_48794,N_49249);
nor UO_4340 (O_4340,N_48946,N_49503);
or UO_4341 (O_4341,N_47605,N_48639);
and UO_4342 (O_4342,N_48864,N_48109);
nand UO_4343 (O_4343,N_49398,N_48237);
and UO_4344 (O_4344,N_49232,N_49724);
and UO_4345 (O_4345,N_47599,N_49371);
nand UO_4346 (O_4346,N_48021,N_47802);
or UO_4347 (O_4347,N_49928,N_48605);
nor UO_4348 (O_4348,N_48486,N_48793);
nand UO_4349 (O_4349,N_48567,N_47821);
nand UO_4350 (O_4350,N_49610,N_49884);
or UO_4351 (O_4351,N_49710,N_48357);
and UO_4352 (O_4352,N_49416,N_49505);
or UO_4353 (O_4353,N_47881,N_47831);
nor UO_4354 (O_4354,N_49955,N_48377);
or UO_4355 (O_4355,N_49113,N_48370);
nand UO_4356 (O_4356,N_49571,N_49726);
or UO_4357 (O_4357,N_49641,N_49710);
nor UO_4358 (O_4358,N_48810,N_49087);
and UO_4359 (O_4359,N_48707,N_49271);
and UO_4360 (O_4360,N_48511,N_47786);
and UO_4361 (O_4361,N_47929,N_48317);
nor UO_4362 (O_4362,N_48873,N_48615);
or UO_4363 (O_4363,N_49997,N_49530);
or UO_4364 (O_4364,N_49062,N_49520);
or UO_4365 (O_4365,N_48152,N_47979);
and UO_4366 (O_4366,N_49997,N_48815);
and UO_4367 (O_4367,N_49771,N_48920);
nand UO_4368 (O_4368,N_47866,N_49118);
and UO_4369 (O_4369,N_49480,N_48674);
xnor UO_4370 (O_4370,N_48960,N_49164);
nor UO_4371 (O_4371,N_48860,N_49782);
or UO_4372 (O_4372,N_49066,N_49445);
xor UO_4373 (O_4373,N_47769,N_48015);
and UO_4374 (O_4374,N_49502,N_48134);
nand UO_4375 (O_4375,N_48234,N_49679);
or UO_4376 (O_4376,N_48881,N_48802);
and UO_4377 (O_4377,N_48489,N_48178);
or UO_4378 (O_4378,N_48200,N_49645);
nor UO_4379 (O_4379,N_49418,N_49840);
nor UO_4380 (O_4380,N_47822,N_48991);
and UO_4381 (O_4381,N_49978,N_49372);
nor UO_4382 (O_4382,N_48438,N_49378);
and UO_4383 (O_4383,N_48288,N_49759);
nor UO_4384 (O_4384,N_48762,N_48005);
and UO_4385 (O_4385,N_48575,N_49479);
nand UO_4386 (O_4386,N_48165,N_48813);
nand UO_4387 (O_4387,N_47713,N_49561);
xnor UO_4388 (O_4388,N_47578,N_49258);
nor UO_4389 (O_4389,N_48755,N_48347);
nand UO_4390 (O_4390,N_48577,N_48793);
nor UO_4391 (O_4391,N_48805,N_48020);
nor UO_4392 (O_4392,N_48695,N_48036);
or UO_4393 (O_4393,N_49152,N_49241);
and UO_4394 (O_4394,N_49962,N_48367);
nor UO_4395 (O_4395,N_48045,N_47810);
nand UO_4396 (O_4396,N_47946,N_49024);
or UO_4397 (O_4397,N_49852,N_47810);
xor UO_4398 (O_4398,N_48197,N_48787);
nand UO_4399 (O_4399,N_48206,N_48297);
nand UO_4400 (O_4400,N_49731,N_48846);
nor UO_4401 (O_4401,N_49790,N_49333);
and UO_4402 (O_4402,N_47862,N_49752);
xnor UO_4403 (O_4403,N_48076,N_49461);
and UO_4404 (O_4404,N_49663,N_48109);
and UO_4405 (O_4405,N_49861,N_47878);
and UO_4406 (O_4406,N_48500,N_49015);
nor UO_4407 (O_4407,N_48725,N_48852);
nor UO_4408 (O_4408,N_49022,N_49116);
nor UO_4409 (O_4409,N_49397,N_49387);
nand UO_4410 (O_4410,N_47824,N_49783);
xor UO_4411 (O_4411,N_47834,N_47556);
and UO_4412 (O_4412,N_49226,N_48324);
nor UO_4413 (O_4413,N_49140,N_49503);
and UO_4414 (O_4414,N_49277,N_47980);
and UO_4415 (O_4415,N_49554,N_49671);
or UO_4416 (O_4416,N_49772,N_48865);
and UO_4417 (O_4417,N_49928,N_49480);
xnor UO_4418 (O_4418,N_49460,N_48176);
and UO_4419 (O_4419,N_48608,N_49908);
or UO_4420 (O_4420,N_48517,N_49016);
or UO_4421 (O_4421,N_48318,N_48280);
or UO_4422 (O_4422,N_48356,N_47855);
or UO_4423 (O_4423,N_48198,N_48620);
and UO_4424 (O_4424,N_48234,N_48634);
or UO_4425 (O_4425,N_47613,N_47985);
nor UO_4426 (O_4426,N_47947,N_49331);
or UO_4427 (O_4427,N_49495,N_48615);
or UO_4428 (O_4428,N_47607,N_48715);
and UO_4429 (O_4429,N_49039,N_47983);
and UO_4430 (O_4430,N_49412,N_48959);
and UO_4431 (O_4431,N_48017,N_49707);
nor UO_4432 (O_4432,N_49313,N_48558);
or UO_4433 (O_4433,N_48784,N_48290);
and UO_4434 (O_4434,N_49531,N_49077);
or UO_4435 (O_4435,N_49317,N_49066);
and UO_4436 (O_4436,N_47910,N_49006);
or UO_4437 (O_4437,N_49481,N_48222);
nor UO_4438 (O_4438,N_49744,N_48260);
or UO_4439 (O_4439,N_48609,N_47547);
nor UO_4440 (O_4440,N_47853,N_49888);
nor UO_4441 (O_4441,N_49809,N_48785);
and UO_4442 (O_4442,N_49741,N_48024);
nor UO_4443 (O_4443,N_47649,N_49781);
or UO_4444 (O_4444,N_48255,N_49991);
nor UO_4445 (O_4445,N_49758,N_49000);
nand UO_4446 (O_4446,N_48495,N_48957);
nand UO_4447 (O_4447,N_49901,N_47991);
and UO_4448 (O_4448,N_48515,N_48919);
nand UO_4449 (O_4449,N_48436,N_49038);
xor UO_4450 (O_4450,N_48404,N_48076);
or UO_4451 (O_4451,N_47703,N_47698);
nor UO_4452 (O_4452,N_47588,N_49292);
xnor UO_4453 (O_4453,N_49023,N_49832);
or UO_4454 (O_4454,N_48968,N_47902);
nand UO_4455 (O_4455,N_49405,N_48277);
or UO_4456 (O_4456,N_48578,N_48860);
or UO_4457 (O_4457,N_47840,N_48933);
nand UO_4458 (O_4458,N_48673,N_48263);
or UO_4459 (O_4459,N_49929,N_49354);
or UO_4460 (O_4460,N_47660,N_48048);
or UO_4461 (O_4461,N_48794,N_47633);
and UO_4462 (O_4462,N_48722,N_49153);
nand UO_4463 (O_4463,N_49511,N_47674);
or UO_4464 (O_4464,N_47618,N_47778);
and UO_4465 (O_4465,N_48431,N_49583);
and UO_4466 (O_4466,N_49229,N_48915);
or UO_4467 (O_4467,N_48730,N_49013);
nand UO_4468 (O_4468,N_48679,N_48409);
nand UO_4469 (O_4469,N_49896,N_48209);
nand UO_4470 (O_4470,N_47920,N_48060);
nor UO_4471 (O_4471,N_48289,N_49265);
or UO_4472 (O_4472,N_49821,N_49956);
nand UO_4473 (O_4473,N_48083,N_49935);
or UO_4474 (O_4474,N_49063,N_49140);
nor UO_4475 (O_4475,N_48909,N_48858);
and UO_4476 (O_4476,N_48092,N_48160);
nor UO_4477 (O_4477,N_49617,N_49090);
nor UO_4478 (O_4478,N_49597,N_48516);
or UO_4479 (O_4479,N_47673,N_48786);
nand UO_4480 (O_4480,N_49802,N_48625);
nor UO_4481 (O_4481,N_49165,N_48914);
or UO_4482 (O_4482,N_48690,N_48320);
or UO_4483 (O_4483,N_47966,N_49645);
and UO_4484 (O_4484,N_49142,N_49497);
xor UO_4485 (O_4485,N_48331,N_47839);
nor UO_4486 (O_4486,N_49933,N_49964);
nand UO_4487 (O_4487,N_48422,N_49924);
nor UO_4488 (O_4488,N_49601,N_49692);
or UO_4489 (O_4489,N_49959,N_49900);
and UO_4490 (O_4490,N_48182,N_48042);
nor UO_4491 (O_4491,N_48347,N_49033);
and UO_4492 (O_4492,N_48292,N_47926);
or UO_4493 (O_4493,N_49642,N_49438);
nand UO_4494 (O_4494,N_47535,N_48689);
nor UO_4495 (O_4495,N_48545,N_47830);
xor UO_4496 (O_4496,N_48981,N_48291);
or UO_4497 (O_4497,N_49547,N_49359);
nor UO_4498 (O_4498,N_48004,N_48054);
or UO_4499 (O_4499,N_48494,N_48597);
nor UO_4500 (O_4500,N_49797,N_48185);
nand UO_4501 (O_4501,N_49710,N_47776);
or UO_4502 (O_4502,N_48746,N_48953);
nand UO_4503 (O_4503,N_48437,N_47736);
or UO_4504 (O_4504,N_49136,N_49487);
and UO_4505 (O_4505,N_49001,N_49229);
nand UO_4506 (O_4506,N_49623,N_49159);
nor UO_4507 (O_4507,N_48406,N_48875);
nand UO_4508 (O_4508,N_49757,N_49622);
and UO_4509 (O_4509,N_49381,N_48523);
and UO_4510 (O_4510,N_49379,N_49567);
xor UO_4511 (O_4511,N_48499,N_48698);
xor UO_4512 (O_4512,N_48200,N_49555);
nand UO_4513 (O_4513,N_49872,N_49630);
nor UO_4514 (O_4514,N_48750,N_49516);
and UO_4515 (O_4515,N_48377,N_48787);
xnor UO_4516 (O_4516,N_47977,N_48743);
nor UO_4517 (O_4517,N_48977,N_48256);
nand UO_4518 (O_4518,N_47727,N_48175);
nand UO_4519 (O_4519,N_48817,N_48946);
nor UO_4520 (O_4520,N_47902,N_49390);
nand UO_4521 (O_4521,N_49707,N_48260);
or UO_4522 (O_4522,N_48701,N_48083);
and UO_4523 (O_4523,N_48680,N_48975);
nor UO_4524 (O_4524,N_49910,N_48974);
or UO_4525 (O_4525,N_48785,N_49907);
nor UO_4526 (O_4526,N_48308,N_49798);
and UO_4527 (O_4527,N_48720,N_47878);
nand UO_4528 (O_4528,N_49500,N_48303);
xor UO_4529 (O_4529,N_49261,N_48647);
or UO_4530 (O_4530,N_48894,N_49962);
or UO_4531 (O_4531,N_49877,N_47638);
nor UO_4532 (O_4532,N_47812,N_49863);
xor UO_4533 (O_4533,N_49445,N_49970);
and UO_4534 (O_4534,N_48483,N_49748);
xor UO_4535 (O_4535,N_49689,N_48213);
and UO_4536 (O_4536,N_48169,N_47840);
nor UO_4537 (O_4537,N_47934,N_49671);
xnor UO_4538 (O_4538,N_47646,N_49834);
xnor UO_4539 (O_4539,N_48683,N_48857);
and UO_4540 (O_4540,N_47868,N_48707);
xor UO_4541 (O_4541,N_47604,N_49256);
or UO_4542 (O_4542,N_48378,N_48865);
or UO_4543 (O_4543,N_48456,N_47609);
xor UO_4544 (O_4544,N_49830,N_48246);
or UO_4545 (O_4545,N_48212,N_47962);
nor UO_4546 (O_4546,N_48736,N_49375);
and UO_4547 (O_4547,N_49969,N_49499);
or UO_4548 (O_4548,N_48547,N_49364);
nand UO_4549 (O_4549,N_47532,N_47731);
or UO_4550 (O_4550,N_48509,N_49866);
or UO_4551 (O_4551,N_49697,N_49725);
and UO_4552 (O_4552,N_49686,N_49573);
or UO_4553 (O_4553,N_48061,N_47990);
nand UO_4554 (O_4554,N_49984,N_48513);
nand UO_4555 (O_4555,N_47792,N_49778);
or UO_4556 (O_4556,N_49318,N_49148);
or UO_4557 (O_4557,N_47512,N_49189);
xor UO_4558 (O_4558,N_49266,N_49090);
nand UO_4559 (O_4559,N_49544,N_47926);
nand UO_4560 (O_4560,N_49537,N_48446);
and UO_4561 (O_4561,N_47863,N_47787);
or UO_4562 (O_4562,N_49426,N_49562);
nand UO_4563 (O_4563,N_47748,N_48490);
or UO_4564 (O_4564,N_47777,N_48189);
or UO_4565 (O_4565,N_48074,N_49916);
and UO_4566 (O_4566,N_48270,N_49688);
nor UO_4567 (O_4567,N_49267,N_47690);
or UO_4568 (O_4568,N_48933,N_47915);
and UO_4569 (O_4569,N_47766,N_49024);
and UO_4570 (O_4570,N_48352,N_49113);
or UO_4571 (O_4571,N_47944,N_48042);
or UO_4572 (O_4572,N_48896,N_48860);
and UO_4573 (O_4573,N_48326,N_47754);
and UO_4574 (O_4574,N_48353,N_48958);
and UO_4575 (O_4575,N_48598,N_48822);
or UO_4576 (O_4576,N_48142,N_47559);
and UO_4577 (O_4577,N_49773,N_48212);
and UO_4578 (O_4578,N_47854,N_47598);
or UO_4579 (O_4579,N_47587,N_48740);
or UO_4580 (O_4580,N_48806,N_49544);
and UO_4581 (O_4581,N_48548,N_47836);
nand UO_4582 (O_4582,N_48717,N_48400);
or UO_4583 (O_4583,N_48066,N_49653);
or UO_4584 (O_4584,N_48186,N_48663);
nand UO_4585 (O_4585,N_49390,N_48923);
nor UO_4586 (O_4586,N_48548,N_49520);
nand UO_4587 (O_4587,N_48214,N_48877);
and UO_4588 (O_4588,N_47972,N_47780);
nor UO_4589 (O_4589,N_47765,N_48354);
or UO_4590 (O_4590,N_48484,N_48272);
and UO_4591 (O_4591,N_49482,N_48878);
and UO_4592 (O_4592,N_48644,N_49415);
or UO_4593 (O_4593,N_47615,N_49710);
or UO_4594 (O_4594,N_49331,N_49590);
or UO_4595 (O_4595,N_48077,N_48918);
xnor UO_4596 (O_4596,N_49352,N_47520);
nand UO_4597 (O_4597,N_48895,N_49714);
nand UO_4598 (O_4598,N_49353,N_49792);
nand UO_4599 (O_4599,N_48715,N_48235);
and UO_4600 (O_4600,N_48423,N_48903);
nand UO_4601 (O_4601,N_49227,N_48416);
nor UO_4602 (O_4602,N_47912,N_48539);
nand UO_4603 (O_4603,N_49742,N_48127);
and UO_4604 (O_4604,N_49809,N_47709);
or UO_4605 (O_4605,N_48392,N_47733);
and UO_4606 (O_4606,N_48034,N_49946);
or UO_4607 (O_4607,N_47824,N_49248);
or UO_4608 (O_4608,N_48228,N_49552);
nand UO_4609 (O_4609,N_48151,N_48492);
and UO_4610 (O_4610,N_48612,N_48701);
and UO_4611 (O_4611,N_49095,N_49933);
and UO_4612 (O_4612,N_48981,N_48937);
nor UO_4613 (O_4613,N_48466,N_47911);
or UO_4614 (O_4614,N_47776,N_48776);
or UO_4615 (O_4615,N_48055,N_48627);
nor UO_4616 (O_4616,N_48336,N_49041);
nand UO_4617 (O_4617,N_49715,N_48268);
xor UO_4618 (O_4618,N_48032,N_49243);
and UO_4619 (O_4619,N_49781,N_48808);
and UO_4620 (O_4620,N_48582,N_48288);
and UO_4621 (O_4621,N_47581,N_49299);
or UO_4622 (O_4622,N_48755,N_49435);
and UO_4623 (O_4623,N_49900,N_49061);
and UO_4624 (O_4624,N_49162,N_48740);
nor UO_4625 (O_4625,N_49784,N_49981);
xnor UO_4626 (O_4626,N_48859,N_48702);
and UO_4627 (O_4627,N_48901,N_49212);
nor UO_4628 (O_4628,N_48888,N_48695);
and UO_4629 (O_4629,N_48778,N_48650);
nand UO_4630 (O_4630,N_49500,N_49643);
or UO_4631 (O_4631,N_48382,N_48495);
or UO_4632 (O_4632,N_48946,N_48952);
or UO_4633 (O_4633,N_49876,N_48869);
or UO_4634 (O_4634,N_49990,N_47904);
nand UO_4635 (O_4635,N_47931,N_49205);
nor UO_4636 (O_4636,N_49479,N_48822);
or UO_4637 (O_4637,N_48526,N_49989);
xnor UO_4638 (O_4638,N_48995,N_49354);
and UO_4639 (O_4639,N_49292,N_49328);
nor UO_4640 (O_4640,N_49683,N_49407);
or UO_4641 (O_4641,N_47681,N_47666);
and UO_4642 (O_4642,N_49544,N_49122);
nand UO_4643 (O_4643,N_47529,N_47949);
nand UO_4644 (O_4644,N_48325,N_49670);
and UO_4645 (O_4645,N_48316,N_48762);
nor UO_4646 (O_4646,N_49434,N_49025);
nand UO_4647 (O_4647,N_48207,N_49950);
nand UO_4648 (O_4648,N_47722,N_47617);
or UO_4649 (O_4649,N_47589,N_48978);
or UO_4650 (O_4650,N_48209,N_47947);
or UO_4651 (O_4651,N_48906,N_48028);
or UO_4652 (O_4652,N_48541,N_48372);
or UO_4653 (O_4653,N_47907,N_47908);
or UO_4654 (O_4654,N_49651,N_47506);
or UO_4655 (O_4655,N_49188,N_49638);
and UO_4656 (O_4656,N_47594,N_49986);
nor UO_4657 (O_4657,N_48547,N_47517);
or UO_4658 (O_4658,N_48241,N_49019);
nand UO_4659 (O_4659,N_49140,N_49797);
or UO_4660 (O_4660,N_48714,N_49522);
nand UO_4661 (O_4661,N_48147,N_49214);
nor UO_4662 (O_4662,N_49116,N_48228);
and UO_4663 (O_4663,N_49126,N_48841);
or UO_4664 (O_4664,N_48740,N_49353);
or UO_4665 (O_4665,N_48057,N_47576);
xnor UO_4666 (O_4666,N_49472,N_49341);
nand UO_4667 (O_4667,N_48756,N_47587);
nand UO_4668 (O_4668,N_48816,N_49391);
xnor UO_4669 (O_4669,N_48821,N_48452);
and UO_4670 (O_4670,N_48875,N_48078);
nor UO_4671 (O_4671,N_48347,N_48580);
nor UO_4672 (O_4672,N_49370,N_48215);
nand UO_4673 (O_4673,N_47969,N_49852);
nor UO_4674 (O_4674,N_49932,N_47919);
and UO_4675 (O_4675,N_49073,N_49638);
and UO_4676 (O_4676,N_48457,N_47858);
nor UO_4677 (O_4677,N_49575,N_48612);
and UO_4678 (O_4678,N_49006,N_48628);
xnor UO_4679 (O_4679,N_49796,N_47944);
and UO_4680 (O_4680,N_48457,N_49187);
and UO_4681 (O_4681,N_48212,N_49345);
nand UO_4682 (O_4682,N_48437,N_49504);
nand UO_4683 (O_4683,N_49014,N_49746);
or UO_4684 (O_4684,N_49212,N_48772);
and UO_4685 (O_4685,N_49669,N_47717);
nor UO_4686 (O_4686,N_49658,N_48891);
or UO_4687 (O_4687,N_48916,N_48887);
xor UO_4688 (O_4688,N_49867,N_48355);
and UO_4689 (O_4689,N_49738,N_49059);
and UO_4690 (O_4690,N_48753,N_48640);
xnor UO_4691 (O_4691,N_47547,N_48824);
nor UO_4692 (O_4692,N_48705,N_48823);
xnor UO_4693 (O_4693,N_49329,N_48136);
nand UO_4694 (O_4694,N_48633,N_47509);
and UO_4695 (O_4695,N_48417,N_47591);
or UO_4696 (O_4696,N_48975,N_49492);
and UO_4697 (O_4697,N_48486,N_49369);
and UO_4698 (O_4698,N_48118,N_49017);
nor UO_4699 (O_4699,N_49241,N_48788);
nor UO_4700 (O_4700,N_49305,N_48884);
nand UO_4701 (O_4701,N_48121,N_48892);
nor UO_4702 (O_4702,N_49491,N_48555);
nand UO_4703 (O_4703,N_49874,N_49440);
nand UO_4704 (O_4704,N_49678,N_49430);
and UO_4705 (O_4705,N_49134,N_48297);
nor UO_4706 (O_4706,N_48073,N_47510);
and UO_4707 (O_4707,N_49542,N_47708);
nand UO_4708 (O_4708,N_49757,N_49867);
or UO_4709 (O_4709,N_48886,N_48026);
and UO_4710 (O_4710,N_49395,N_49320);
nor UO_4711 (O_4711,N_49741,N_48121);
nor UO_4712 (O_4712,N_48603,N_49610);
nor UO_4713 (O_4713,N_47638,N_48792);
or UO_4714 (O_4714,N_48444,N_48516);
and UO_4715 (O_4715,N_48682,N_49200);
nor UO_4716 (O_4716,N_48102,N_47823);
xor UO_4717 (O_4717,N_48147,N_48687);
and UO_4718 (O_4718,N_49627,N_48032);
nor UO_4719 (O_4719,N_48276,N_48659);
xor UO_4720 (O_4720,N_49320,N_49805);
and UO_4721 (O_4721,N_48317,N_49689);
and UO_4722 (O_4722,N_49414,N_48445);
nor UO_4723 (O_4723,N_48077,N_49143);
nand UO_4724 (O_4724,N_49019,N_49074);
and UO_4725 (O_4725,N_47862,N_49135);
nand UO_4726 (O_4726,N_49555,N_48164);
nand UO_4727 (O_4727,N_49819,N_47873);
xnor UO_4728 (O_4728,N_49272,N_48901);
xor UO_4729 (O_4729,N_48072,N_49465);
or UO_4730 (O_4730,N_48725,N_48230);
or UO_4731 (O_4731,N_49049,N_48092);
or UO_4732 (O_4732,N_48521,N_49517);
xor UO_4733 (O_4733,N_49164,N_49728);
or UO_4734 (O_4734,N_49044,N_49575);
nor UO_4735 (O_4735,N_49760,N_48820);
xor UO_4736 (O_4736,N_48939,N_49300);
or UO_4737 (O_4737,N_47989,N_47527);
and UO_4738 (O_4738,N_48269,N_48597);
nand UO_4739 (O_4739,N_49549,N_48013);
nand UO_4740 (O_4740,N_47643,N_48466);
nor UO_4741 (O_4741,N_49915,N_49748);
and UO_4742 (O_4742,N_49145,N_48027);
nor UO_4743 (O_4743,N_47965,N_49861);
nor UO_4744 (O_4744,N_47972,N_48962);
and UO_4745 (O_4745,N_47960,N_48102);
and UO_4746 (O_4746,N_49810,N_48948);
nand UO_4747 (O_4747,N_47667,N_48095);
or UO_4748 (O_4748,N_48306,N_48919);
nor UO_4749 (O_4749,N_48630,N_48096);
and UO_4750 (O_4750,N_48474,N_48054);
or UO_4751 (O_4751,N_49529,N_47729);
nor UO_4752 (O_4752,N_49480,N_49750);
xor UO_4753 (O_4753,N_48539,N_48174);
nand UO_4754 (O_4754,N_49054,N_49181);
and UO_4755 (O_4755,N_48268,N_49501);
nor UO_4756 (O_4756,N_49242,N_49057);
nor UO_4757 (O_4757,N_48406,N_48685);
or UO_4758 (O_4758,N_47764,N_49716);
and UO_4759 (O_4759,N_47982,N_48351);
or UO_4760 (O_4760,N_48622,N_48471);
and UO_4761 (O_4761,N_47769,N_48538);
nor UO_4762 (O_4762,N_49973,N_48601);
nor UO_4763 (O_4763,N_48953,N_48390);
or UO_4764 (O_4764,N_49530,N_49441);
nor UO_4765 (O_4765,N_49291,N_49215);
nor UO_4766 (O_4766,N_48199,N_49719);
nand UO_4767 (O_4767,N_48331,N_48486);
and UO_4768 (O_4768,N_49861,N_49858);
nand UO_4769 (O_4769,N_48633,N_48227);
nor UO_4770 (O_4770,N_49584,N_48376);
nor UO_4771 (O_4771,N_49558,N_49365);
and UO_4772 (O_4772,N_47631,N_48045);
and UO_4773 (O_4773,N_48077,N_48282);
and UO_4774 (O_4774,N_48446,N_47863);
nor UO_4775 (O_4775,N_48041,N_49590);
nand UO_4776 (O_4776,N_49611,N_49625);
or UO_4777 (O_4777,N_49794,N_49392);
or UO_4778 (O_4778,N_49982,N_48125);
and UO_4779 (O_4779,N_47520,N_48403);
xor UO_4780 (O_4780,N_49647,N_48343);
nor UO_4781 (O_4781,N_47737,N_49743);
or UO_4782 (O_4782,N_48410,N_48277);
nor UO_4783 (O_4783,N_48925,N_49493);
nor UO_4784 (O_4784,N_48240,N_49617);
nor UO_4785 (O_4785,N_48062,N_48697);
nor UO_4786 (O_4786,N_49502,N_48823);
and UO_4787 (O_4787,N_49037,N_49775);
or UO_4788 (O_4788,N_48459,N_48568);
nor UO_4789 (O_4789,N_48502,N_49021);
or UO_4790 (O_4790,N_48920,N_49123);
nand UO_4791 (O_4791,N_49577,N_49180);
nor UO_4792 (O_4792,N_48230,N_48789);
or UO_4793 (O_4793,N_49450,N_48794);
and UO_4794 (O_4794,N_49571,N_48450);
nand UO_4795 (O_4795,N_48350,N_49345);
nand UO_4796 (O_4796,N_48764,N_49078);
and UO_4797 (O_4797,N_49630,N_47676);
nand UO_4798 (O_4798,N_48488,N_47597);
and UO_4799 (O_4799,N_49003,N_48686);
nor UO_4800 (O_4800,N_49200,N_49796);
nor UO_4801 (O_4801,N_49689,N_48932);
or UO_4802 (O_4802,N_49634,N_48643);
nor UO_4803 (O_4803,N_47736,N_48558);
and UO_4804 (O_4804,N_47856,N_49349);
nor UO_4805 (O_4805,N_49585,N_48093);
nor UO_4806 (O_4806,N_48358,N_47816);
nor UO_4807 (O_4807,N_48397,N_48498);
nand UO_4808 (O_4808,N_47868,N_48201);
or UO_4809 (O_4809,N_49971,N_49043);
nor UO_4810 (O_4810,N_48828,N_48795);
nand UO_4811 (O_4811,N_49868,N_49943);
xor UO_4812 (O_4812,N_48151,N_49947);
nor UO_4813 (O_4813,N_49554,N_48135);
nand UO_4814 (O_4814,N_48222,N_49007);
and UO_4815 (O_4815,N_49922,N_47943);
and UO_4816 (O_4816,N_47621,N_48089);
and UO_4817 (O_4817,N_48227,N_48722);
nand UO_4818 (O_4818,N_48349,N_49814);
nand UO_4819 (O_4819,N_48082,N_49552);
nor UO_4820 (O_4820,N_49052,N_48170);
nand UO_4821 (O_4821,N_49228,N_47661);
and UO_4822 (O_4822,N_48070,N_48754);
xnor UO_4823 (O_4823,N_49593,N_49440);
and UO_4824 (O_4824,N_49358,N_49035);
or UO_4825 (O_4825,N_48793,N_49574);
and UO_4826 (O_4826,N_48326,N_48479);
nor UO_4827 (O_4827,N_49967,N_49985);
nand UO_4828 (O_4828,N_48200,N_47501);
and UO_4829 (O_4829,N_49616,N_48677);
or UO_4830 (O_4830,N_48397,N_49719);
xnor UO_4831 (O_4831,N_48459,N_47748);
nor UO_4832 (O_4832,N_47836,N_47908);
nor UO_4833 (O_4833,N_49204,N_49274);
or UO_4834 (O_4834,N_48376,N_49586);
and UO_4835 (O_4835,N_49962,N_47813);
nor UO_4836 (O_4836,N_49764,N_47548);
or UO_4837 (O_4837,N_48201,N_48415);
or UO_4838 (O_4838,N_49805,N_47820);
xnor UO_4839 (O_4839,N_49052,N_49874);
and UO_4840 (O_4840,N_48751,N_48269);
or UO_4841 (O_4841,N_47503,N_48147);
xor UO_4842 (O_4842,N_49474,N_48582);
nand UO_4843 (O_4843,N_49589,N_49494);
nor UO_4844 (O_4844,N_49128,N_49337);
xnor UO_4845 (O_4845,N_49639,N_48679);
nor UO_4846 (O_4846,N_48352,N_48197);
or UO_4847 (O_4847,N_47719,N_49093);
or UO_4848 (O_4848,N_49083,N_47956);
nand UO_4849 (O_4849,N_47736,N_47698);
nand UO_4850 (O_4850,N_49831,N_49186);
and UO_4851 (O_4851,N_48462,N_48023);
nand UO_4852 (O_4852,N_48562,N_48548);
or UO_4853 (O_4853,N_47838,N_48140);
or UO_4854 (O_4854,N_49120,N_47901);
nor UO_4855 (O_4855,N_49999,N_48066);
and UO_4856 (O_4856,N_49247,N_48697);
nor UO_4857 (O_4857,N_48757,N_47954);
nor UO_4858 (O_4858,N_49990,N_47741);
nand UO_4859 (O_4859,N_48222,N_48410);
nand UO_4860 (O_4860,N_49382,N_48920);
nor UO_4861 (O_4861,N_48372,N_49552);
nor UO_4862 (O_4862,N_49105,N_48247);
nor UO_4863 (O_4863,N_48872,N_48963);
xor UO_4864 (O_4864,N_49577,N_49919);
nor UO_4865 (O_4865,N_49134,N_47950);
nor UO_4866 (O_4866,N_47542,N_49798);
nor UO_4867 (O_4867,N_49101,N_48641);
or UO_4868 (O_4868,N_49986,N_49851);
nor UO_4869 (O_4869,N_48944,N_48103);
and UO_4870 (O_4870,N_48750,N_48583);
and UO_4871 (O_4871,N_47914,N_49594);
nand UO_4872 (O_4872,N_48785,N_48190);
nand UO_4873 (O_4873,N_49666,N_48632);
nor UO_4874 (O_4874,N_49943,N_48280);
and UO_4875 (O_4875,N_47947,N_48066);
and UO_4876 (O_4876,N_48112,N_47923);
nor UO_4877 (O_4877,N_48014,N_47875);
or UO_4878 (O_4878,N_49591,N_49437);
or UO_4879 (O_4879,N_48480,N_49258);
and UO_4880 (O_4880,N_49978,N_49089);
nand UO_4881 (O_4881,N_48891,N_49108);
nor UO_4882 (O_4882,N_47689,N_47823);
nor UO_4883 (O_4883,N_49841,N_48505);
nor UO_4884 (O_4884,N_48774,N_48150);
or UO_4885 (O_4885,N_48773,N_47565);
nor UO_4886 (O_4886,N_49120,N_47597);
or UO_4887 (O_4887,N_47868,N_48537);
nor UO_4888 (O_4888,N_48531,N_49378);
nor UO_4889 (O_4889,N_48263,N_49109);
nand UO_4890 (O_4890,N_47659,N_48739);
nor UO_4891 (O_4891,N_47701,N_48678);
nand UO_4892 (O_4892,N_49164,N_47500);
xnor UO_4893 (O_4893,N_47669,N_47541);
nand UO_4894 (O_4894,N_49003,N_47661);
or UO_4895 (O_4895,N_47612,N_47984);
xnor UO_4896 (O_4896,N_48177,N_49693);
nand UO_4897 (O_4897,N_47937,N_48306);
and UO_4898 (O_4898,N_47693,N_49351);
nand UO_4899 (O_4899,N_48466,N_49332);
nor UO_4900 (O_4900,N_48626,N_49449);
xnor UO_4901 (O_4901,N_47867,N_49993);
or UO_4902 (O_4902,N_49648,N_49712);
nor UO_4903 (O_4903,N_48731,N_48228);
nor UO_4904 (O_4904,N_48725,N_48607);
xnor UO_4905 (O_4905,N_49415,N_49211);
nand UO_4906 (O_4906,N_49696,N_49574);
xor UO_4907 (O_4907,N_49087,N_47889);
or UO_4908 (O_4908,N_48212,N_47693);
xnor UO_4909 (O_4909,N_49855,N_48215);
xor UO_4910 (O_4910,N_49075,N_48424);
nand UO_4911 (O_4911,N_49249,N_49171);
xor UO_4912 (O_4912,N_48263,N_48821);
and UO_4913 (O_4913,N_49446,N_47815);
xor UO_4914 (O_4914,N_49694,N_48985);
nor UO_4915 (O_4915,N_49675,N_49321);
and UO_4916 (O_4916,N_48312,N_47975);
or UO_4917 (O_4917,N_48344,N_48986);
nor UO_4918 (O_4918,N_49156,N_49867);
nor UO_4919 (O_4919,N_48459,N_49957);
nor UO_4920 (O_4920,N_49319,N_49782);
nand UO_4921 (O_4921,N_49446,N_48310);
and UO_4922 (O_4922,N_48039,N_48587);
xnor UO_4923 (O_4923,N_48503,N_49168);
or UO_4924 (O_4924,N_47882,N_48811);
nand UO_4925 (O_4925,N_48627,N_48763);
or UO_4926 (O_4926,N_48730,N_49881);
xor UO_4927 (O_4927,N_49575,N_49298);
or UO_4928 (O_4928,N_48221,N_48407);
nor UO_4929 (O_4929,N_49041,N_48325);
or UO_4930 (O_4930,N_48874,N_48367);
and UO_4931 (O_4931,N_48575,N_47982);
nor UO_4932 (O_4932,N_48367,N_49785);
and UO_4933 (O_4933,N_48642,N_48130);
nor UO_4934 (O_4934,N_49769,N_47822);
or UO_4935 (O_4935,N_48790,N_49385);
and UO_4936 (O_4936,N_49536,N_47537);
nor UO_4937 (O_4937,N_49357,N_48744);
nand UO_4938 (O_4938,N_47874,N_49451);
and UO_4939 (O_4939,N_47962,N_48071);
nor UO_4940 (O_4940,N_47724,N_48172);
and UO_4941 (O_4941,N_48612,N_49320);
nand UO_4942 (O_4942,N_49300,N_49890);
and UO_4943 (O_4943,N_49701,N_48590);
and UO_4944 (O_4944,N_48817,N_48021);
and UO_4945 (O_4945,N_48116,N_49301);
nand UO_4946 (O_4946,N_48411,N_49652);
or UO_4947 (O_4947,N_47791,N_47675);
or UO_4948 (O_4948,N_49163,N_48824);
nand UO_4949 (O_4949,N_48657,N_48044);
or UO_4950 (O_4950,N_49788,N_48132);
nand UO_4951 (O_4951,N_47716,N_47649);
and UO_4952 (O_4952,N_49900,N_47524);
nor UO_4953 (O_4953,N_48830,N_47647);
nand UO_4954 (O_4954,N_49647,N_48176);
or UO_4955 (O_4955,N_49940,N_49914);
nand UO_4956 (O_4956,N_47553,N_47959);
nand UO_4957 (O_4957,N_48598,N_49685);
nand UO_4958 (O_4958,N_49484,N_48469);
nand UO_4959 (O_4959,N_48357,N_48707);
or UO_4960 (O_4960,N_49686,N_49747);
and UO_4961 (O_4961,N_49715,N_47890);
nand UO_4962 (O_4962,N_48179,N_49681);
or UO_4963 (O_4963,N_48311,N_47971);
and UO_4964 (O_4964,N_47515,N_49552);
nor UO_4965 (O_4965,N_48081,N_48883);
or UO_4966 (O_4966,N_48600,N_48607);
xor UO_4967 (O_4967,N_49243,N_49927);
xor UO_4968 (O_4968,N_49477,N_47903);
nand UO_4969 (O_4969,N_48247,N_48238);
nand UO_4970 (O_4970,N_49583,N_47910);
and UO_4971 (O_4971,N_49616,N_49195);
or UO_4972 (O_4972,N_49691,N_48424);
or UO_4973 (O_4973,N_48785,N_49472);
or UO_4974 (O_4974,N_49141,N_48796);
or UO_4975 (O_4975,N_49377,N_47909);
and UO_4976 (O_4976,N_47644,N_48542);
nand UO_4977 (O_4977,N_48729,N_48949);
xor UO_4978 (O_4978,N_48293,N_48077);
and UO_4979 (O_4979,N_49738,N_47897);
nand UO_4980 (O_4980,N_47539,N_49079);
nor UO_4981 (O_4981,N_49938,N_48060);
or UO_4982 (O_4982,N_47784,N_49949);
nand UO_4983 (O_4983,N_49880,N_48308);
or UO_4984 (O_4984,N_48158,N_48051);
nand UO_4985 (O_4985,N_48380,N_48024);
nand UO_4986 (O_4986,N_49654,N_49206);
nor UO_4987 (O_4987,N_47835,N_49327);
or UO_4988 (O_4988,N_47743,N_48474);
and UO_4989 (O_4989,N_49997,N_49456);
nor UO_4990 (O_4990,N_49067,N_49411);
or UO_4991 (O_4991,N_48709,N_48772);
and UO_4992 (O_4992,N_49416,N_47581);
nor UO_4993 (O_4993,N_49522,N_47579);
nor UO_4994 (O_4994,N_48335,N_48166);
and UO_4995 (O_4995,N_48901,N_49617);
xor UO_4996 (O_4996,N_49214,N_48456);
nor UO_4997 (O_4997,N_49674,N_49913);
nor UO_4998 (O_4998,N_48117,N_48017);
nor UO_4999 (O_4999,N_48387,N_47889);
endmodule