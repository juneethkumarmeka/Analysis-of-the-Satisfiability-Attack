module basic_5000_50000_5000_5_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nor U0 (N_0,In_2017,In_351);
nor U1 (N_1,In_3960,In_3340);
nand U2 (N_2,In_2410,In_4384);
xnor U3 (N_3,In_1082,In_3603);
xnor U4 (N_4,In_1741,In_502);
xnor U5 (N_5,In_449,In_4252);
and U6 (N_6,In_1284,In_14);
and U7 (N_7,In_538,In_3098);
or U8 (N_8,In_1719,In_1476);
nor U9 (N_9,In_2071,In_529);
nand U10 (N_10,In_751,In_4239);
or U11 (N_11,In_4065,In_3396);
or U12 (N_12,In_2494,In_1804);
nor U13 (N_13,In_3195,In_3882);
nand U14 (N_14,In_307,In_1248);
nor U15 (N_15,In_1825,In_3978);
and U16 (N_16,In_3198,In_1515);
nor U17 (N_17,In_1819,In_1483);
nor U18 (N_18,In_1982,In_4025);
and U19 (N_19,In_765,In_2755);
or U20 (N_20,In_2427,In_2531);
and U21 (N_21,In_1312,In_3889);
nand U22 (N_22,In_1875,In_3533);
and U23 (N_23,In_3707,In_3815);
nor U24 (N_24,In_455,In_4807);
and U25 (N_25,In_1184,In_4578);
nor U26 (N_26,In_2969,In_4417);
or U27 (N_27,In_1813,In_1259);
nor U28 (N_28,In_4876,In_3299);
or U29 (N_29,In_717,In_984);
or U30 (N_30,In_2746,In_4776);
or U31 (N_31,In_1932,In_2495);
and U32 (N_32,In_3155,In_3296);
nand U33 (N_33,In_740,In_2174);
and U34 (N_34,In_3138,In_4579);
or U35 (N_35,In_2881,In_3478);
nand U36 (N_36,In_2943,In_2236);
or U37 (N_37,In_677,In_1787);
nand U38 (N_38,In_2005,In_3105);
and U39 (N_39,In_2735,In_924);
and U40 (N_40,In_1058,In_3969);
and U41 (N_41,In_265,In_389);
and U42 (N_42,In_1583,In_4800);
or U43 (N_43,In_1298,In_2786);
nor U44 (N_44,In_4764,In_3315);
xor U45 (N_45,In_22,In_4018);
and U46 (N_46,In_4130,In_4170);
nand U47 (N_47,In_1255,In_3725);
xor U48 (N_48,In_4601,In_4224);
nor U49 (N_49,In_510,In_2161);
xnor U50 (N_50,In_2777,In_1037);
or U51 (N_51,In_4363,In_2973);
and U52 (N_52,In_1480,In_4699);
nor U53 (N_53,In_3568,In_4445);
or U54 (N_54,In_3625,In_746);
or U55 (N_55,In_2854,In_1696);
xor U56 (N_56,In_554,In_4458);
or U57 (N_57,In_3827,In_3481);
and U58 (N_58,In_4533,In_3185);
and U59 (N_59,In_956,In_829);
nor U60 (N_60,In_3559,In_4275);
nand U61 (N_61,In_2576,In_907);
and U62 (N_62,In_4482,In_1160);
and U63 (N_63,In_808,In_382);
or U64 (N_64,In_3666,In_3916);
or U65 (N_65,In_3667,In_4167);
nand U66 (N_66,In_2519,In_4189);
nor U67 (N_67,In_23,In_4113);
and U68 (N_68,In_4325,In_3722);
nand U69 (N_69,In_1580,In_2268);
or U70 (N_70,In_2369,In_50);
nor U71 (N_71,In_3201,In_272);
nor U72 (N_72,In_4432,In_3663);
nor U73 (N_73,In_4536,In_1874);
xor U74 (N_74,In_2074,In_153);
and U75 (N_75,In_4956,In_2364);
nand U76 (N_76,In_4368,In_1214);
and U77 (N_77,In_3131,In_4913);
and U78 (N_78,In_4727,In_3197);
nor U79 (N_79,In_2607,In_4808);
nor U80 (N_80,In_1537,In_3653);
nand U81 (N_81,In_3290,In_711);
xor U82 (N_82,In_1943,In_2840);
or U83 (N_83,In_4382,In_2158);
xor U84 (N_84,In_226,In_4453);
nand U85 (N_85,In_1220,In_3788);
nand U86 (N_86,In_1912,In_1253);
xnor U87 (N_87,In_3675,In_934);
and U88 (N_88,In_4545,In_628);
nand U89 (N_89,In_3780,In_994);
xnor U90 (N_90,In_3638,In_2434);
xnor U91 (N_91,In_2563,In_1050);
or U92 (N_92,In_3819,In_4086);
or U93 (N_93,In_4401,In_42);
and U94 (N_94,In_345,In_1439);
nand U95 (N_95,In_3136,In_2116);
or U96 (N_96,In_1654,In_2716);
and U97 (N_97,In_1520,In_4331);
or U98 (N_98,In_318,In_1285);
xor U99 (N_99,In_173,In_4901);
and U100 (N_100,In_450,In_1780);
nor U101 (N_101,In_965,In_1083);
or U102 (N_102,In_832,In_1022);
nand U103 (N_103,In_3767,In_4833);
nor U104 (N_104,In_4959,In_2258);
or U105 (N_105,In_3432,In_1574);
nand U106 (N_106,In_4046,In_1479);
nor U107 (N_107,In_1901,In_3464);
or U108 (N_108,In_931,In_235);
xor U109 (N_109,In_2053,In_1613);
or U110 (N_110,In_2260,In_1796);
and U111 (N_111,In_192,In_4079);
nor U112 (N_112,In_41,In_1227);
nor U113 (N_113,In_761,In_1842);
nor U114 (N_114,In_3522,In_1935);
xor U115 (N_115,In_1704,In_3879);
and U116 (N_116,In_1258,In_2954);
nand U117 (N_117,In_191,In_4440);
or U118 (N_118,In_3427,In_3945);
nand U119 (N_119,In_4469,In_3293);
nor U120 (N_120,In_511,In_3062);
nand U121 (N_121,In_3918,In_848);
nor U122 (N_122,In_1350,In_1544);
nor U123 (N_123,In_3632,In_4870);
and U124 (N_124,In_1611,In_4400);
xor U125 (N_125,In_1548,In_2029);
and U126 (N_126,In_1824,In_3110);
xor U127 (N_127,In_3554,In_904);
xor U128 (N_128,In_2640,In_1217);
or U129 (N_129,In_3364,In_3965);
or U130 (N_130,In_4675,In_2857);
and U131 (N_131,In_732,In_3408);
nand U132 (N_132,In_4549,In_4403);
nand U133 (N_133,In_2201,In_2220);
xnor U134 (N_134,In_567,In_1942);
xnor U135 (N_135,In_1718,In_3004);
or U136 (N_136,In_3431,In_3567);
xnor U137 (N_137,In_3924,In_424);
nand U138 (N_138,In_3348,In_2899);
nor U139 (N_139,In_2978,In_4017);
nor U140 (N_140,In_1313,In_4567);
xnor U141 (N_141,In_3444,In_653);
nand U142 (N_142,In_2305,In_255);
and U143 (N_143,In_2717,In_1386);
and U144 (N_144,In_4525,In_4067);
nand U145 (N_145,In_1742,In_2023);
nor U146 (N_146,In_301,In_2584);
xor U147 (N_147,In_1535,In_4970);
and U148 (N_148,In_4663,In_3096);
and U149 (N_149,In_2030,In_3613);
and U150 (N_150,In_4611,In_201);
nand U151 (N_151,In_2614,In_2882);
xnor U152 (N_152,In_2965,In_3850);
xnor U153 (N_153,In_3497,In_2350);
nor U154 (N_154,In_327,In_3394);
and U155 (N_155,In_3005,In_2693);
nand U156 (N_156,In_164,In_1713);
nor U157 (N_157,In_1797,In_982);
xor U158 (N_158,In_4635,In_1158);
and U159 (N_159,In_294,In_1534);
nor U160 (N_160,In_2493,In_1146);
or U161 (N_161,In_4791,In_4528);
nand U162 (N_162,In_943,In_2621);
and U163 (N_163,In_3825,In_4514);
nor U164 (N_164,In_2246,In_3515);
nor U165 (N_165,In_3223,In_4850);
nand U166 (N_166,In_4941,In_412);
and U167 (N_167,In_2018,In_2011);
nand U168 (N_168,In_132,In_2467);
and U169 (N_169,In_1044,In_4677);
xnor U170 (N_170,In_3808,In_3082);
and U171 (N_171,In_2183,In_4042);
nand U172 (N_172,In_2935,In_684);
xor U173 (N_173,In_4268,In_3450);
nor U174 (N_174,In_1820,In_2571);
nor U175 (N_175,In_1585,In_3032);
nor U176 (N_176,In_1529,In_1090);
or U177 (N_177,In_702,In_3243);
or U178 (N_178,In_1053,In_0);
xor U179 (N_179,In_3804,In_496);
nor U180 (N_180,In_1474,In_1157);
nand U181 (N_181,In_4561,In_46);
nand U182 (N_182,In_2994,In_1076);
nor U183 (N_183,In_3207,In_3587);
nor U184 (N_184,In_257,In_372);
nor U185 (N_185,In_241,In_1646);
or U186 (N_186,In_331,In_2912);
nor U187 (N_187,In_2413,In_3246);
nor U188 (N_188,In_3038,In_213);
nor U189 (N_189,In_166,In_4124);
xnor U190 (N_190,In_3671,In_264);
nor U191 (N_191,In_3412,In_1377);
and U192 (N_192,In_4883,In_423);
nor U193 (N_193,In_1633,In_2166);
and U194 (N_194,In_4949,In_1149);
nor U195 (N_195,In_2279,In_3742);
or U196 (N_196,In_3120,In_2654);
nand U197 (N_197,In_3174,In_3754);
and U198 (N_198,In_784,In_4947);
or U199 (N_199,In_3764,In_2293);
and U200 (N_200,In_2237,In_1062);
and U201 (N_201,In_2995,In_2468);
nand U202 (N_202,In_663,In_3048);
nor U203 (N_203,In_1635,In_3115);
and U204 (N_204,In_4479,In_3188);
nor U205 (N_205,In_4143,In_2538);
xor U206 (N_206,In_1996,In_769);
or U207 (N_207,In_83,In_2147);
nor U208 (N_208,In_3451,In_851);
or U209 (N_209,In_3205,In_518);
and U210 (N_210,In_3285,In_927);
nor U211 (N_211,In_2918,In_3329);
nand U212 (N_212,In_3463,In_2006);
and U213 (N_213,In_3558,In_3291);
and U214 (N_214,In_4342,In_2356);
or U215 (N_215,In_647,In_3582);
and U216 (N_216,In_2908,In_649);
and U217 (N_217,In_472,In_1614);
nor U218 (N_218,In_200,In_3358);
and U219 (N_219,In_1136,In_1941);
xnor U220 (N_220,In_523,In_3287);
and U221 (N_221,In_11,In_2224);
or U222 (N_222,In_599,In_2856);
and U223 (N_223,In_4010,In_4043);
nand U224 (N_224,In_2322,In_2250);
and U225 (N_225,In_2915,In_707);
xor U226 (N_226,In_4147,In_2172);
nor U227 (N_227,In_3706,In_3523);
nor U228 (N_228,In_1148,In_2781);
nand U229 (N_229,In_1540,In_3061);
nand U230 (N_230,In_2133,In_2405);
nand U231 (N_231,In_3392,In_3413);
nor U232 (N_232,In_1620,In_2221);
and U233 (N_233,In_1594,In_3462);
nand U234 (N_234,In_2437,In_569);
or U235 (N_235,In_3782,In_661);
or U236 (N_236,In_121,In_3863);
nand U237 (N_237,In_959,In_1547);
xor U238 (N_238,In_1222,In_2428);
nand U239 (N_239,In_3772,In_456);
or U240 (N_240,In_857,In_1393);
xnor U241 (N_241,In_1738,In_4412);
or U242 (N_242,In_2546,In_274);
and U243 (N_243,In_2326,In_4072);
or U244 (N_244,In_749,In_1208);
xnor U245 (N_245,In_2549,In_1098);
and U246 (N_246,In_2176,In_1055);
nor U247 (N_247,In_664,In_3307);
nor U248 (N_248,In_2034,In_3812);
and U249 (N_249,In_1297,In_4954);
nor U250 (N_250,In_2970,In_285);
xnor U251 (N_251,In_2265,In_921);
or U252 (N_252,In_2831,In_2698);
and U253 (N_253,In_2270,In_1038);
nor U254 (N_254,In_882,In_4009);
xor U255 (N_255,In_3240,In_4872);
or U256 (N_256,In_4289,In_4311);
or U257 (N_257,In_332,In_4983);
and U258 (N_258,In_3487,In_1555);
or U259 (N_259,In_1325,In_148);
nor U260 (N_260,In_533,In_4217);
and U261 (N_261,In_3901,In_4696);
nand U262 (N_262,In_3502,In_2660);
nand U263 (N_263,In_3360,In_3292);
nand U264 (N_264,In_4308,In_2910);
and U265 (N_265,In_940,In_2163);
nor U266 (N_266,In_2819,In_1133);
and U267 (N_267,In_1884,In_3275);
nand U268 (N_268,In_4165,In_1914);
nand U269 (N_269,In_3775,In_3343);
nand U270 (N_270,In_4612,In_612);
nor U271 (N_271,In_2003,In_1952);
or U272 (N_272,In_3491,In_217);
xor U273 (N_273,In_3622,In_4016);
nand U274 (N_274,In_3732,In_2386);
nand U275 (N_275,In_1968,In_4939);
nor U276 (N_276,In_4175,In_4334);
and U277 (N_277,In_1652,In_1482);
or U278 (N_278,In_308,In_625);
nor U279 (N_279,In_3703,In_3844);
nor U280 (N_280,In_3083,In_1945);
nor U281 (N_281,In_3159,In_3897);
nand U282 (N_282,In_3561,In_2867);
or U283 (N_283,In_2771,In_2475);
xor U284 (N_284,In_1846,In_2838);
nor U285 (N_285,In_4467,In_1166);
nor U286 (N_286,In_1923,In_3849);
xor U287 (N_287,In_3304,In_4407);
nor U288 (N_288,In_4554,In_4837);
nand U289 (N_289,In_4907,In_3893);
nand U290 (N_290,In_4662,In_1992);
or U291 (N_291,In_3002,In_2848);
nand U292 (N_292,In_4874,In_3453);
and U293 (N_293,In_514,In_3847);
xnor U294 (N_294,In_3779,In_2824);
nand U295 (N_295,In_1116,In_1637);
nand U296 (N_296,In_4069,In_913);
nand U297 (N_297,In_4704,In_3405);
xor U298 (N_298,In_2797,In_4212);
or U299 (N_299,In_1930,In_4492);
xnor U300 (N_300,In_4098,In_1740);
xor U301 (N_301,In_1073,In_4512);
nand U302 (N_302,In_2589,In_1273);
nand U303 (N_303,In_4498,In_4793);
nor U304 (N_304,In_3014,In_1957);
or U305 (N_305,In_188,In_4250);
nand U306 (N_306,In_172,In_609);
and U307 (N_307,In_2067,In_1805);
xor U308 (N_308,In_2684,In_555);
or U309 (N_309,In_3132,In_1512);
xnor U310 (N_310,In_1059,In_1697);
and U311 (N_311,In_892,In_2836);
or U312 (N_312,In_4111,In_4355);
and U313 (N_313,In_2573,In_4826);
xor U314 (N_314,In_3086,In_1918);
or U315 (N_315,In_2395,In_2411);
nand U316 (N_316,In_2752,In_2896);
xor U317 (N_317,In_4032,In_3261);
nor U318 (N_318,In_1448,In_798);
nand U319 (N_319,In_905,In_3320);
or U320 (N_320,In_92,In_754);
or U321 (N_321,In_2049,In_2232);
nand U322 (N_322,In_2533,In_2674);
or U323 (N_323,In_4792,In_2566);
xnor U324 (N_324,In_2945,In_1356);
nor U325 (N_325,In_2521,In_592);
nor U326 (N_326,In_1703,In_422);
or U327 (N_327,In_930,In_3127);
or U328 (N_328,In_1997,In_1627);
or U329 (N_329,In_3680,In_3161);
nor U330 (N_330,In_3359,In_2464);
or U331 (N_331,In_3026,In_1553);
nor U332 (N_332,In_708,In_305);
xnor U333 (N_333,In_4877,In_4429);
nor U334 (N_334,In_2630,In_1649);
and U335 (N_335,In_2929,In_1881);
and U336 (N_336,In_2524,In_1488);
and U337 (N_337,In_1127,In_3736);
nor U338 (N_338,In_4955,In_566);
or U339 (N_339,In_3909,In_4166);
or U340 (N_340,In_4026,In_4491);
or U341 (N_341,In_1497,In_16);
nor U342 (N_342,In_1868,In_540);
xor U343 (N_343,In_4716,In_577);
xnor U344 (N_344,In_4717,In_3460);
nand U345 (N_345,In_2765,In_2175);
xor U346 (N_346,In_2466,In_694);
nand U347 (N_347,In_3250,In_3607);
xor U348 (N_348,In_2933,In_2100);
xnor U349 (N_349,In_712,In_1500);
nor U350 (N_350,In_3281,In_1140);
nand U351 (N_351,In_1759,In_6);
or U352 (N_352,In_150,In_838);
xor U353 (N_353,In_3398,In_1833);
xnor U354 (N_354,In_1985,In_1579);
and U355 (N_355,In_2042,In_3573);
xor U356 (N_356,In_452,In_2064);
or U357 (N_357,In_2024,In_219);
xnor U358 (N_358,In_3441,In_4327);
nor U359 (N_359,In_3152,In_2903);
nand U360 (N_360,In_1106,In_2972);
nand U361 (N_361,In_3406,In_4530);
and U362 (N_362,In_1379,In_2155);
xnor U363 (N_363,In_4434,In_4535);
xor U364 (N_364,In_895,In_1145);
nand U365 (N_365,In_4379,In_3309);
or U366 (N_366,In_4868,In_3644);
xor U367 (N_367,In_3410,In_2449);
xnor U368 (N_368,In_1270,In_716);
nor U369 (N_369,In_339,In_3778);
xor U370 (N_370,In_2827,In_64);
and U371 (N_371,In_1773,In_3226);
xor U372 (N_372,In_3721,In_1906);
nor U373 (N_373,In_4692,In_1192);
nand U374 (N_374,In_4348,In_2877);
and U375 (N_375,In_1195,In_742);
nand U376 (N_376,In_1486,In_879);
nor U377 (N_377,In_2188,In_768);
nor U378 (N_378,In_503,In_1089);
or U379 (N_379,In_419,In_2880);
nor U380 (N_380,In_4693,In_2096);
xor U381 (N_381,In_4015,In_850);
nand U382 (N_382,In_1871,In_4701);
nand U383 (N_383,In_1844,In_435);
xor U384 (N_384,In_2715,In_3436);
xnor U385 (N_385,In_1861,In_1563);
nor U386 (N_386,In_120,In_440);
xor U387 (N_387,In_3058,In_3486);
xnor U388 (N_388,In_665,In_4039);
nand U389 (N_389,In_2825,In_3690);
nand U390 (N_390,In_2117,In_3325);
nand U391 (N_391,In_3649,In_3758);
or U392 (N_392,In_4516,In_1228);
xor U393 (N_393,In_3621,In_2196);
nor U394 (N_394,In_2312,In_4673);
and U395 (N_395,In_1523,In_3579);
and U396 (N_396,In_1736,In_1609);
and U397 (N_397,In_2319,In_4511);
and U398 (N_398,In_4084,In_3118);
and U399 (N_399,In_442,In_721);
or U400 (N_400,In_1463,In_4423);
xor U401 (N_401,In_2558,In_506);
nor U402 (N_402,In_2365,In_3683);
or U403 (N_403,In_1802,In_3485);
nand U404 (N_404,In_4919,In_919);
or U405 (N_405,In_2807,In_1444);
xor U406 (N_406,In_1401,In_4085);
nand U407 (N_407,In_3516,In_786);
or U408 (N_408,In_156,In_3387);
and U409 (N_409,In_4182,In_655);
and U410 (N_410,In_4672,In_618);
nand U411 (N_411,In_556,In_1999);
nor U412 (N_412,In_3279,In_3763);
and U413 (N_413,In_1032,In_1416);
nand U414 (N_414,In_643,In_98);
or U415 (N_415,In_73,In_3608);
xnor U416 (N_416,In_2885,In_3113);
nand U417 (N_417,In_4729,In_425);
or U418 (N_418,In_2832,In_4745);
nand U419 (N_419,In_552,In_2636);
and U420 (N_420,In_3762,In_770);
nor U421 (N_421,In_2491,In_4713);
xnor U422 (N_422,In_1645,In_2488);
nand U423 (N_423,In_1408,In_40);
or U424 (N_424,In_4809,In_1114);
nor U425 (N_425,In_4644,In_4075);
xnor U426 (N_426,In_1998,In_1893);
nand U427 (N_427,In_2383,In_18);
or U428 (N_428,In_3941,In_3454);
and U429 (N_429,In_3248,In_2041);
or U430 (N_430,In_3711,In_2271);
nor U431 (N_431,In_2678,In_3739);
and U432 (N_432,In_1684,In_1206);
nor U433 (N_433,In_3846,In_590);
nand U434 (N_434,In_2639,In_2523);
xnor U435 (N_435,In_1698,In_1749);
and U436 (N_436,In_1229,In_194);
nor U437 (N_437,In_2685,In_2381);
or U438 (N_438,In_1430,In_447);
nor U439 (N_439,In_2424,In_1880);
xnor U440 (N_440,In_2105,In_3799);
or U441 (N_441,In_4152,In_4141);
nand U442 (N_442,In_343,In_2429);
nand U443 (N_443,In_3591,In_1245);
and U444 (N_444,In_4569,In_3337);
and U445 (N_445,In_1175,In_3678);
and U446 (N_446,In_3685,In_3407);
nand U447 (N_447,In_2153,In_1337);
xnor U448 (N_448,In_3543,In_4006);
nor U449 (N_449,In_1933,In_3230);
xnor U450 (N_450,In_4125,In_2677);
nand U451 (N_451,In_3121,In_1702);
xor U452 (N_452,In_3416,In_3996);
or U453 (N_453,In_375,In_2726);
and U454 (N_454,In_431,In_3662);
nor U455 (N_455,In_598,In_818);
and U456 (N_456,In_3975,In_312);
xnor U457 (N_457,In_2901,In_3848);
and U458 (N_458,In_4366,In_756);
nor U459 (N_459,In_3595,In_709);
or U460 (N_460,In_3877,In_575);
xnor U461 (N_461,In_2643,In_4736);
nand U462 (N_462,In_4266,In_1276);
or U463 (N_463,In_10,In_2486);
nand U464 (N_464,In_4183,In_3614);
nand U465 (N_465,In_1100,In_3520);
nor U466 (N_466,In_4508,In_3972);
and U467 (N_467,In_380,In_718);
nor U468 (N_468,In_1584,In_1752);
xor U469 (N_469,In_2399,In_2095);
xnor U470 (N_470,In_2472,In_1552);
xor U471 (N_471,In_4587,In_1503);
or U472 (N_472,In_3903,In_1068);
nor U473 (N_473,In_2393,In_320);
nor U474 (N_474,In_1883,In_2559);
and U475 (N_475,In_3075,In_2306);
nor U476 (N_476,In_129,In_2400);
xnor U477 (N_477,In_1168,In_3070);
nand U478 (N_478,In_3245,In_4690);
nor U479 (N_479,In_4679,In_410);
nor U480 (N_480,In_3615,In_3457);
and U481 (N_481,In_2308,In_2724);
nor U482 (N_482,In_189,In_364);
nor U483 (N_483,In_1927,In_427);
nor U484 (N_484,In_1250,In_53);
xor U485 (N_485,In_171,In_4786);
and U486 (N_486,In_386,In_2780);
nand U487 (N_487,In_396,In_2760);
and U488 (N_488,In_757,In_1672);
nor U489 (N_489,In_2782,In_779);
nor U490 (N_490,In_1582,In_4999);
nand U491 (N_491,In_1412,In_1036);
nand U492 (N_492,In_145,In_929);
xor U493 (N_493,In_2477,In_4078);
nor U494 (N_494,In_2079,In_3066);
or U495 (N_495,In_1882,In_898);
nor U496 (N_496,In_3222,In_2567);
nand U497 (N_497,In_1043,In_1021);
xor U498 (N_498,In_1154,In_3040);
or U499 (N_499,In_831,In_3955);
xnor U500 (N_500,In_2154,In_2861);
or U501 (N_501,In_151,In_3802);
nor U502 (N_502,In_3569,In_1256);
xor U503 (N_503,In_2088,In_4639);
and U504 (N_504,In_4652,In_2344);
and U505 (N_505,In_4988,In_4921);
and U506 (N_506,In_3215,In_1224);
or U507 (N_507,In_1319,In_1177);
nor U508 (N_508,In_4742,In_4925);
nand U509 (N_509,In_3344,In_2853);
xnor U510 (N_510,In_2691,In_4159);
nor U511 (N_511,In_2851,In_3545);
or U512 (N_512,In_2507,In_4688);
and U513 (N_513,In_3842,In_2200);
xnor U514 (N_514,In_107,In_1651);
nand U515 (N_515,In_369,In_3947);
and U516 (N_516,In_932,In_492);
or U517 (N_517,In_2921,In_578);
nand U518 (N_518,In_2159,In_522);
and U519 (N_519,In_734,In_1330);
xor U520 (N_520,In_1295,In_4556);
and U521 (N_521,In_1420,In_443);
or U522 (N_522,In_3599,In_3228);
or U523 (N_523,In_4986,In_3570);
nand U524 (N_524,In_976,In_760);
nand U525 (N_525,In_870,In_2700);
nor U526 (N_526,In_4007,In_2961);
or U527 (N_527,In_771,In_571);
or U528 (N_528,In_2846,In_2979);
nor U529 (N_529,In_268,In_2951);
and U530 (N_530,In_4573,In_2906);
nand U531 (N_531,In_3134,In_1054);
or U532 (N_532,In_4433,In_572);
nor U533 (N_533,In_1015,In_4769);
and U534 (N_534,In_112,In_4995);
nand U535 (N_535,In_1783,In_111);
xor U536 (N_536,In_3894,In_4576);
nor U537 (N_537,In_2632,In_1370);
and U538 (N_538,In_3718,In_933);
or U539 (N_539,In_3505,In_293);
nor U540 (N_540,In_1438,In_365);
xor U541 (N_541,In_4819,In_610);
xor U542 (N_542,In_2151,In_2408);
nor U543 (N_543,In_330,In_1744);
nor U544 (N_544,In_2913,In_4409);
and U545 (N_545,In_4276,In_1308);
and U546 (N_546,In_1449,In_204);
nor U547 (N_547,In_3949,In_2645);
or U548 (N_548,In_1770,In_388);
xor U549 (N_549,In_123,In_827);
nor U550 (N_550,In_84,In_1623);
nor U551 (N_551,In_2069,In_2252);
nor U552 (N_552,In_400,In_2865);
nor U553 (N_553,In_4774,In_116);
nand U554 (N_554,In_2438,In_3456);
nand U555 (N_555,In_4201,In_3724);
and U556 (N_556,In_58,In_1834);
and U557 (N_557,In_3748,In_4123);
nor U558 (N_558,In_69,In_3705);
xor U559 (N_559,In_1761,In_4157);
nand U560 (N_560,In_2339,In_3104);
nand U561 (N_561,In_3529,In_570);
xor U562 (N_562,In_1750,In_2606);
and U563 (N_563,In_2214,In_821);
and U564 (N_564,In_4277,In_3571);
nor U565 (N_565,In_3494,In_1953);
xor U566 (N_566,In_1226,In_4711);
xnor U567 (N_567,In_3087,In_3750);
nor U568 (N_568,In_1955,In_4896);
nand U569 (N_569,In_3046,In_4634);
nor U570 (N_570,In_2808,In_2944);
xor U571 (N_571,In_2202,In_2609);
nor U572 (N_572,In_1657,In_4744);
nor U573 (N_573,In_4021,In_4260);
or U574 (N_574,In_3506,In_283);
and U575 (N_575,In_1045,In_3604);
and U576 (N_576,In_1920,In_2812);
nand U577 (N_577,In_4595,In_4647);
or U578 (N_578,In_1959,In_2007);
and U579 (N_579,In_4703,In_2968);
xor U580 (N_580,In_2092,In_2932);
and U581 (N_581,In_1056,In_1292);
xor U582 (N_582,In_4838,In_2770);
xor U583 (N_583,In_77,In_210);
nor U584 (N_584,In_4537,In_167);
nand U585 (N_585,In_1965,In_3578);
nand U586 (N_586,In_4356,In_2757);
or U587 (N_587,In_3154,In_3717);
and U588 (N_588,In_2907,In_723);
or U589 (N_589,In_3274,In_1929);
or U590 (N_590,In_143,In_3146);
and U591 (N_591,In_3759,In_208);
or U592 (N_592,In_476,In_3470);
nand U593 (N_593,In_2705,In_773);
nand U594 (N_594,In_3107,In_2180);
and U595 (N_595,In_544,In_2977);
nor U596 (N_596,In_4979,In_4880);
or U597 (N_597,In_958,In_641);
or U598 (N_598,In_2355,In_1180);
nand U599 (N_599,In_4659,In_3393);
xor U600 (N_600,In_871,In_964);
xor U601 (N_601,In_4628,In_3238);
nand U602 (N_602,In_4044,In_4816);
nand U603 (N_603,In_1691,In_3313);
xnor U604 (N_604,In_1332,In_1267);
and U605 (N_605,In_4349,In_3019);
or U606 (N_606,In_3402,In_4758);
and U607 (N_607,In_3473,In_3824);
xor U608 (N_608,In_693,In_311);
xor U609 (N_609,In_763,In_4169);
xnor U610 (N_610,In_2686,In_2199);
nand U611 (N_611,In_31,In_80);
and U612 (N_612,In_2633,In_2351);
and U613 (N_613,In_4852,In_3791);
or U614 (N_614,In_2320,In_119);
nor U615 (N_615,In_3192,In_4755);
nor U616 (N_616,In_4886,In_2697);
or U617 (N_617,In_4419,In_4242);
or U618 (N_618,In_1341,In_2334);
and U619 (N_619,In_162,In_4884);
or U620 (N_620,In_109,In_2510);
nand U621 (N_621,In_2102,In_1278);
and U622 (N_622,In_3986,In_2616);
and U623 (N_623,In_714,In_849);
or U624 (N_624,In_2459,In_1493);
nor U625 (N_625,In_1794,In_185);
and U626 (N_626,In_774,In_4697);
and U627 (N_627,In_1690,In_4689);
or U628 (N_628,In_4396,In_3106);
xor U629 (N_629,In_3610,In_474);
nand U630 (N_630,In_374,In_3433);
nand U631 (N_631,In_3959,In_4864);
nand U632 (N_632,In_3194,In_3301);
nand U633 (N_633,In_2307,In_4613);
nor U634 (N_634,In_974,In_4293);
or U635 (N_635,In_3179,In_1699);
xnor U636 (N_636,In_4665,In_3713);
and U637 (N_637,In_3227,In_147);
nand U638 (N_638,In_3760,In_1518);
nor U639 (N_639,In_3870,In_2313);
or U640 (N_640,In_2874,In_2718);
and U641 (N_641,In_1171,In_3288);
nor U642 (N_642,In_3422,In_2423);
and U643 (N_643,In_3231,In_4114);
xnor U644 (N_644,In_1357,In_4420);
and U645 (N_645,In_3057,In_3267);
xor U646 (N_646,In_935,In_1000);
nor U647 (N_647,In_2522,In_1095);
and U648 (N_648,In_2646,In_2340);
nor U649 (N_649,In_926,In_4574);
xor U650 (N_650,In_2436,In_1818);
nand U651 (N_651,In_3964,In_3856);
and U652 (N_652,In_2021,In_4917);
or U653 (N_653,In_4814,In_4797);
nor U654 (N_654,In_1215,In_807);
or U655 (N_655,In_519,In_4859);
and U656 (N_656,In_2281,In_1269);
and U657 (N_657,In_3864,In_4763);
xor U658 (N_658,In_1977,In_3974);
xnor U659 (N_659,In_261,In_3388);
or U660 (N_660,In_2253,In_1019);
nor U661 (N_661,In_59,In_3896);
nor U662 (N_662,In_1849,In_4054);
and U663 (N_663,In_4899,In_3813);
nand U664 (N_664,In_1424,In_825);
or U665 (N_665,In_4456,In_1235);
nand U666 (N_666,In_9,In_531);
nand U667 (N_667,In_224,In_2430);
xor U668 (N_668,In_3609,In_1779);
nor U669 (N_669,In_1949,In_2834);
nand U670 (N_670,In_3377,In_405);
xnor U671 (N_671,In_3455,In_4783);
nand U672 (N_672,In_4686,In_1204);
nand U673 (N_673,In_1388,In_4274);
nand U674 (N_674,In_3234,In_3080);
nand U675 (N_675,In_1088,In_2164);
nor U676 (N_676,In_826,In_1924);
nor U677 (N_677,In_3314,In_2348);
nor U678 (N_678,In_3907,In_1628);
and U679 (N_679,In_245,In_1179);
nor U680 (N_680,In_3670,In_4625);
nor U681 (N_681,In_4413,In_4720);
nor U682 (N_682,In_4386,In_1468);
nor U683 (N_683,In_4258,In_1991);
xnor U684 (N_684,In_1491,In_4832);
nand U685 (N_685,In_1018,In_1461);
nor U686 (N_686,In_2963,In_1351);
xor U687 (N_687,In_1169,In_465);
nor U688 (N_688,In_1679,In_1212);
or U689 (N_689,In_3389,In_3043);
nor U690 (N_690,In_3141,In_1134);
nor U691 (N_691,In_4333,In_1971);
nand U692 (N_692,In_2238,In_3646);
and U693 (N_693,In_4847,In_4097);
nand U694 (N_694,In_2012,In_4314);
nand U695 (N_695,In_3961,In_1870);
and U696 (N_696,In_3111,In_2722);
and U697 (N_697,In_2733,In_4952);
nand U698 (N_698,In_2353,In_3731);
xnor U699 (N_699,In_117,In_3629);
nand U700 (N_700,In_2879,In_954);
xor U701 (N_701,In_1233,In_1835);
and U702 (N_702,In_1937,In_3566);
nand U703 (N_703,In_1467,In_781);
nor U704 (N_704,In_3884,In_2863);
xor U705 (N_705,In_4316,In_3880);
nor U706 (N_706,In_88,In_4132);
xnor U707 (N_707,In_4603,In_1119);
xor U708 (N_708,In_4996,In_2296);
or U709 (N_709,In_2261,In_4524);
nor U710 (N_710,In_4892,In_298);
nand U711 (N_711,In_3727,In_2656);
and U712 (N_712,In_3177,In_662);
xnor U713 (N_713,In_2799,In_4139);
xnor U714 (N_714,In_2871,In_315);
nor U715 (N_715,In_4309,In_4653);
nor U716 (N_716,In_1051,In_4813);
nand U717 (N_717,In_206,In_4402);
xnor U718 (N_718,In_1403,In_4888);
nand U719 (N_719,In_1619,In_4991);
nor U720 (N_720,In_1423,In_4609);
nor U721 (N_721,In_4971,In_2694);
or U722 (N_722,In_1610,In_1590);
nor U723 (N_723,In_113,In_1469);
nand U724 (N_724,In_4518,In_3381);
nor U725 (N_725,In_1859,In_4426);
or U726 (N_726,In_4509,In_3593);
and U727 (N_727,In_178,In_2182);
or U728 (N_728,In_2560,In_1550);
xnor U729 (N_729,In_4718,In_4154);
nor U730 (N_730,In_2124,In_2985);
nand U731 (N_731,In_2565,In_353);
nand U732 (N_732,In_1629,In_4782);
nand U733 (N_733,In_3513,In_3490);
and U734 (N_734,In_3940,In_3347);
nor U735 (N_735,In_2998,In_3560);
nor U736 (N_736,In_2000,In_3510);
nor U737 (N_737,In_279,In_1855);
nand U738 (N_738,In_4975,In_2337);
nand U739 (N_739,In_4738,In_3777);
nor U740 (N_740,In_1900,In_2215);
or U741 (N_741,In_4885,In_1693);
xnor U742 (N_742,In_2068,In_134);
nor U743 (N_743,In_1602,In_815);
or U744 (N_744,In_2278,In_4427);
or U745 (N_745,In_1290,In_3446);
and U746 (N_746,In_3468,In_2602);
nand U747 (N_747,In_2803,In_4606);
or U748 (N_748,In_2815,In_1978);
and U749 (N_749,In_2070,In_2373);
nand U750 (N_750,In_3100,In_2942);
or U751 (N_751,In_3531,In_4472);
nor U752 (N_752,In_2756,In_1596);
xor U753 (N_753,In_2625,In_1832);
xor U754 (N_754,In_1631,In_1706);
xnor U755 (N_755,In_4700,In_3994);
or U756 (N_756,In_3800,In_1237);
xnor U757 (N_757,In_4929,In_3442);
nor U758 (N_758,In_4493,In_1108);
and U759 (N_759,In_841,In_230);
and U760 (N_760,In_1790,In_4544);
nand U761 (N_761,In_4712,In_988);
or U762 (N_762,In_2482,In_39);
or U763 (N_763,In_3977,In_1185);
and U764 (N_764,In_1810,In_1315);
nand U765 (N_765,In_4036,In_2764);
nand U766 (N_766,In_3376,In_3429);
nor U767 (N_767,In_2476,In_4616);
or U768 (N_768,In_814,In_1501);
nand U769 (N_769,In_1791,In_2747);
nand U770 (N_770,In_1895,In_229);
or U771 (N_771,In_295,In_2627);
and U772 (N_772,In_3339,In_202);
xor U773 (N_773,In_4617,In_889);
or U774 (N_774,In_918,In_698);
nand U775 (N_775,In_1198,In_1907);
and U776 (N_776,In_1567,In_4047);
nand U777 (N_777,In_3125,In_1183);
or U778 (N_778,In_4449,In_539);
or U779 (N_779,In_2091,In_3374);
nand U780 (N_780,In_4218,In_3836);
nor U781 (N_781,In_1807,In_868);
nand U782 (N_782,In_2592,In_411);
xnor U783 (N_783,In_2108,In_1092);
nand U784 (N_784,In_4927,In_4762);
nand U785 (N_785,In_833,In_3493);
nor U786 (N_786,In_2352,In_1647);
xor U787 (N_787,In_130,In_1006);
or U788 (N_788,In_4008,In_3517);
or U789 (N_789,In_1951,In_3674);
nor U790 (N_790,In_4262,In_634);
nand U791 (N_791,In_1521,In_2775);
nand U792 (N_792,In_2480,In_4073);
xor U793 (N_793,In_3776,In_393);
and U794 (N_794,In_3117,In_2295);
or U795 (N_795,In_3810,In_1422);
or U796 (N_796,In_4138,In_2543);
nor U797 (N_797,In_4570,In_4004);
xor U798 (N_798,In_3160,In_4784);
and U799 (N_799,In_2085,In_68);
or U800 (N_800,In_2409,In_384);
nor U801 (N_801,In_4168,In_49);
and U802 (N_802,In_2131,In_3987);
nand U803 (N_803,In_1575,In_2991);
or U804 (N_804,In_759,In_2924);
nand U805 (N_805,In_2635,In_673);
nand U806 (N_806,In_4360,In_2226);
nand U807 (N_807,In_2368,In_685);
nor U808 (N_808,In_696,In_2010);
nor U809 (N_809,In_886,In_4903);
and U810 (N_810,In_3063,In_2110);
nand U811 (N_811,In_3526,In_809);
and U812 (N_812,In_2759,In_290);
xnor U813 (N_813,In_3773,In_2552);
xor U814 (N_814,In_2455,In_2283);
nor U815 (N_815,In_252,In_817);
xor U816 (N_816,In_2058,In_3126);
and U817 (N_817,In_2890,In_20);
xor U818 (N_818,In_2316,In_3886);
nor U819 (N_819,In_3472,In_4060);
and U820 (N_820,In_1656,In_3867);
nand U821 (N_821,In_4369,In_2629);
nor U822 (N_822,In_4871,In_4630);
and U823 (N_823,In_4261,In_1743);
xnor U824 (N_824,In_4291,In_1668);
and U825 (N_825,In_1241,In_4538);
nand U826 (N_826,In_144,In_4746);
or U827 (N_827,In_3029,In_3375);
or U828 (N_828,In_2833,In_2648);
and U829 (N_829,In_3200,In_3910);
nor U830 (N_830,In_2888,In_475);
nand U831 (N_831,In_2557,In_4594);
nor U832 (N_832,In_2539,In_4622);
xor U833 (N_833,In_4563,In_4708);
nand U834 (N_834,In_1838,In_942);
nor U835 (N_835,In_4362,In_4656);
nand U836 (N_836,In_1346,In_2959);
nor U837 (N_837,In_595,In_4186);
and U838 (N_838,In_3229,In_1748);
and U839 (N_839,In_579,In_1607);
and U840 (N_840,In_3581,In_2448);
and U841 (N_841,In_3575,In_3756);
and U842 (N_842,In_2862,In_1317);
and U843 (N_843,In_660,In_3247);
and U844 (N_844,In_467,In_3984);
and U845 (N_845,In_559,In_3997);
or U846 (N_846,In_1845,In_4893);
nor U847 (N_847,In_1731,In_543);
xnor U848 (N_848,In_277,In_4461);
or U849 (N_849,In_1049,In_4344);
or U850 (N_850,In_854,In_3257);
nand U851 (N_851,In_4685,In_802);
or U852 (N_852,In_482,In_2870);
or U853 (N_853,In_1029,In_2192);
nand U854 (N_854,In_4615,In_4202);
or U855 (N_855,In_3728,In_2389);
and U856 (N_856,In_2778,In_4964);
nor U857 (N_857,In_1514,In_2297);
or U858 (N_858,In_3306,In_344);
or U859 (N_859,In_2086,In_4540);
xor U860 (N_860,In_3242,In_3633);
xnor U861 (N_861,In_966,In_4798);
or U862 (N_862,In_3536,In_2666);
nand U863 (N_863,In_4294,In_2650);
xor U864 (N_864,In_2033,In_4588);
nor U865 (N_865,In_1511,In_1776);
or U866 (N_866,In_4521,In_3166);
and U867 (N_867,In_2442,In_681);
and U868 (N_868,In_2664,In_1326);
xor U869 (N_869,In_299,In_3163);
nor U870 (N_870,In_1903,In_764);
or U871 (N_871,In_4714,In_1873);
or U872 (N_872,In_2976,In_1020);
or U873 (N_873,In_3912,In_2047);
nand U874 (N_874,In_1343,In_2687);
nand U875 (N_875,In_3737,In_4751);
xnor U876 (N_876,In_1969,In_368);
nand U877 (N_877,In_4406,In_48);
or U878 (N_878,In_297,In_2039);
nand U879 (N_879,In_2624,In_1648);
and U880 (N_880,In_669,In_3602);
xor U881 (N_881,In_813,In_3303);
and U882 (N_882,In_4279,In_4121);
and U883 (N_883,In_4878,In_4082);
xor U884 (N_884,In_4297,In_2419);
or U885 (N_885,In_1686,In_819);
nor U886 (N_886,In_3953,In_448);
nor U887 (N_887,In_4526,In_3003);
and U888 (N_888,In_4064,In_3122);
nor U889 (N_889,In_3469,In_269);
nor U890 (N_890,In_244,In_2456);
and U891 (N_891,In_254,In_925);
or U892 (N_892,In_4215,In_4100);
nor U893 (N_893,In_1457,In_2842);
nand U894 (N_894,In_3657,In_484);
or U895 (N_895,In_1928,In_1338);
or U896 (N_896,In_1451,In_176);
or U897 (N_897,In_1425,In_2015);
nor U898 (N_898,In_2119,In_2958);
xor U899 (N_899,In_3740,In_1321);
and U900 (N_900,In_672,In_480);
nor U901 (N_901,In_4338,In_2194);
or U902 (N_902,In_1618,In_2282);
or U903 (N_903,In_381,In_352);
and U904 (N_904,In_1669,In_2801);
or U905 (N_905,In_4306,In_3151);
nand U906 (N_906,In_1390,In_1674);
nand U907 (N_907,In_2138,In_2919);
and U908 (N_908,In_1956,In_2121);
nor U909 (N_909,In_2335,In_2795);
nor U910 (N_910,In_2583,In_3875);
or U911 (N_911,In_4145,In_1887);
nand U912 (N_912,In_4657,In_2481);
nor U913 (N_913,In_75,In_135);
xor U914 (N_914,In_4142,In_568);
xor U915 (N_915,In_1194,In_2287);
and U916 (N_916,In_2130,In_3251);
and U917 (N_917,In_3651,In_704);
or U918 (N_918,In_2662,In_3769);
xnor U919 (N_919,In_887,In_2181);
nor U920 (N_920,In_902,In_4965);
nand U921 (N_921,In_3335,In_1231);
xnor U922 (N_922,In_928,In_3328);
nor U923 (N_923,In_3269,In_3385);
nand U924 (N_924,In_995,In_2371);
xor U925 (N_925,In_3135,In_451);
and U926 (N_926,In_1132,In_1830);
nand U927 (N_927,In_2541,In_1174);
nand U928 (N_928,In_3744,In_2986);
nand U929 (N_929,In_174,In_1879);
nor U930 (N_930,In_2742,In_4370);
xor U931 (N_931,In_1323,In_4933);
xnor U932 (N_932,In_138,In_3710);
nor U933 (N_933,In_990,In_2391);
and U934 (N_934,In_4926,In_4591);
or U935 (N_935,In_391,In_4890);
xor U936 (N_936,In_4352,In_1334);
and U937 (N_937,In_1570,In_2198);
nand U938 (N_938,In_3150,In_992);
and U939 (N_939,In_4916,In_2922);
nand U940 (N_940,In_2048,In_478);
nand U941 (N_941,In_4781,In_720);
and U942 (N_942,In_3009,In_2608);
xnor U943 (N_943,In_4193,In_358);
xnor U944 (N_944,In_2813,In_4920);
nand U945 (N_945,In_3958,In_2556);
and U946 (N_946,In_4473,In_260);
nand U947 (N_947,In_823,In_3642);
nand U948 (N_948,In_894,In_4969);
xor U949 (N_949,In_2983,In_461);
xnor U950 (N_950,In_3798,In_1728);
and U951 (N_951,In_3746,In_2016);
nand U952 (N_952,In_1589,In_1415);
nand U953 (N_953,In_1406,In_2025);
or U954 (N_954,In_1592,In_3101);
nor U955 (N_955,In_890,In_1886);
nand U956 (N_956,In_3224,In_2873);
xor U957 (N_957,In_4505,In_938);
nand U958 (N_958,In_4829,In_4943);
or U959 (N_959,In_1465,In_1533);
nor U960 (N_960,In_2971,In_2542);
and U961 (N_961,In_1435,In_4312);
and U962 (N_962,In_2148,In_154);
xnor U963 (N_963,In_3266,In_3668);
and U964 (N_964,In_2298,In_1296);
nor U965 (N_965,In_1359,In_2738);
xnor U966 (N_966,In_3059,In_668);
xor U967 (N_967,In_4229,In_1200);
xnor U968 (N_968,In_4961,In_3899);
nor U969 (N_969,In_4088,In_3208);
and U970 (N_970,In_3654,In_4757);
xnor U971 (N_971,In_4731,In_2575);
nor U972 (N_972,In_897,In_3322);
nand U973 (N_973,In_2314,In_90);
xnor U974 (N_974,In_81,In_970);
or U975 (N_975,In_957,In_2384);
nor U976 (N_976,In_4869,In_1443);
or U977 (N_977,In_603,In_4255);
xor U978 (N_978,In_3995,In_842);
nor U979 (N_979,In_3682,In_4754);
or U980 (N_980,In_4083,In_2516);
xnor U981 (N_981,In_947,In_4621);
or U982 (N_982,In_347,In_2858);
and U983 (N_983,In_8,In_416);
nor U984 (N_984,In_1121,In_334);
nand U985 (N_985,In_1381,In_866);
or U986 (N_986,In_1163,In_1375);
nor U987 (N_987,In_4735,In_1004);
nand U988 (N_988,In_4364,In_987);
nor U989 (N_989,In_142,In_3199);
or U990 (N_990,In_3428,In_1039);
nand U991 (N_991,In_165,In_891);
or U992 (N_992,In_105,In_1642);
nand U993 (N_993,In_1123,In_4902);
and U994 (N_994,In_747,In_3461);
nor U995 (N_995,In_788,In_650);
nand U996 (N_996,In_3276,In_2241);
and U997 (N_997,In_2680,In_2875);
nand U998 (N_998,In_2822,In_3165);
nand U999 (N_999,In_1275,In_4452);
and U1000 (N_1000,In_4862,In_51);
and U1001 (N_1001,In_4681,In_4393);
and U1002 (N_1002,In_3936,In_4070);
nor U1003 (N_1003,In_546,In_4380);
nor U1004 (N_1004,In_3546,In_2478);
nand U1005 (N_1005,In_3140,In_3130);
nor U1006 (N_1006,In_3641,In_2113);
and U1007 (N_1007,In_4873,In_1111);
nor U1008 (N_1008,In_2515,In_4766);
and U1009 (N_1009,In_376,In_1009);
nor U1010 (N_1010,In_169,In_4843);
nand U1011 (N_1011,In_1970,In_4990);
xnor U1012 (N_1012,In_2610,In_494);
nand U1013 (N_1013,In_2233,In_1453);
and U1014 (N_1014,In_2779,In_3658);
nor U1015 (N_1015,In_2225,In_1339);
and U1016 (N_1016,In_782,In_319);
nand U1017 (N_1017,In_594,In_735);
nor U1018 (N_1018,In_3921,In_1407);
xor U1019 (N_1019,In_4858,In_4454);
and U1020 (N_1020,In_1792,In_3555);
xor U1021 (N_1021,In_4803,In_4394);
nor U1022 (N_1022,In_470,In_909);
and U1023 (N_1023,In_4992,In_4089);
nor U1024 (N_1024,In_3885,In_1694);
nand U1025 (N_1025,In_266,In_3803);
or U1026 (N_1026,In_1564,In_1472);
nor U1027 (N_1027,In_4887,In_1364);
nand U1028 (N_1028,In_4438,In_4317);
nand U1029 (N_1029,In_3049,In_258);
nor U1030 (N_1030,In_3838,In_2111);
nand U1031 (N_1031,In_3187,In_3535);
nor U1032 (N_1032,In_4592,In_824);
nor U1033 (N_1033,In_1509,In_4210);
nor U1034 (N_1034,In_706,In_3056);
nor U1035 (N_1035,In_722,In_949);
or U1036 (N_1036,In_865,In_2044);
nor U1037 (N_1037,In_2157,In_1385);
or U1038 (N_1038,In_3440,In_4496);
and U1039 (N_1039,In_536,In_363);
xor U1040 (N_1040,In_54,In_3249);
xnor U1041 (N_1041,In_3114,In_1244);
nand U1042 (N_1042,In_3418,In_1559);
nor U1043 (N_1043,In_2534,In_1280);
xnor U1044 (N_1044,In_4195,In_454);
nand U1045 (N_1045,In_608,In_1104);
and U1046 (N_1046,In_1661,In_3701);
nand U1047 (N_1047,In_877,In_4749);
or U1048 (N_1048,In_1551,In_3189);
nor U1049 (N_1049,In_3102,In_810);
and U1050 (N_1050,In_205,In_118);
xnor U1051 (N_1051,In_2762,In_2128);
and U1052 (N_1052,In_4226,In_243);
nor U1053 (N_1053,In_2425,In_1925);
and U1054 (N_1054,In_2300,In_3927);
nand U1055 (N_1055,In_1726,In_262);
xnor U1056 (N_1056,In_2905,In_1456);
and U1057 (N_1057,In_4867,In_2235);
xor U1058 (N_1058,In_2421,In_562);
nor U1059 (N_1059,In_2962,In_4940);
nand U1060 (N_1060,In_3297,In_359);
and U1061 (N_1061,In_1432,In_4027);
xor U1062 (N_1062,In_1960,In_3507);
xor U1063 (N_1063,In_3008,In_1101);
and U1064 (N_1064,In_4115,In_3785);
or U1065 (N_1065,In_941,In_2251);
nor U1066 (N_1066,In_2872,In_3183);
and U1067 (N_1067,In_2445,In_4817);
nand U1068 (N_1068,In_528,In_4415);
and U1069 (N_1069,In_35,In_1139);
nor U1070 (N_1070,In_3443,In_4358);
or U1071 (N_1071,In_2753,In_1302);
nand U1072 (N_1072,In_899,In_3382);
nand U1073 (N_1073,In_2382,In_3091);
nor U1074 (N_1074,In_4494,In_3676);
nand U1075 (N_1075,In_211,In_3256);
nor U1076 (N_1076,In_4655,In_2989);
nor U1077 (N_1077,In_1188,In_2280);
nor U1078 (N_1078,In_2349,In_1722);
nor U1079 (N_1079,In_1291,In_597);
nand U1080 (N_1080,In_1349,In_152);
nand U1081 (N_1081,In_1264,In_2139);
nor U1082 (N_1082,In_1897,In_1685);
and U1083 (N_1083,In_3537,In_3051);
nand U1084 (N_1084,In_955,In_910);
nand U1085 (N_1085,In_923,In_3726);
and U1086 (N_1086,In_2730,In_4636);
nor U1087 (N_1087,In_2544,In_1155);
xor U1088 (N_1088,In_1545,In_3645);
nand U1089 (N_1089,In_4739,In_1203);
nand U1090 (N_1090,In_4811,In_1380);
and U1091 (N_1091,In_341,In_3011);
xor U1092 (N_1092,In_3729,In_2767);
nor U1093 (N_1093,In_3316,In_348);
xor U1094 (N_1094,In_3967,In_2537);
and U1095 (N_1095,In_3373,In_3647);
or U1096 (N_1096,In_3547,In_1961);
and U1097 (N_1097,In_322,In_2526);
nand U1098 (N_1098,In_4126,In_4777);
xnor U1099 (N_1099,In_2452,In_4529);
xnor U1100 (N_1100,In_1524,In_1107);
and U1101 (N_1101,In_2343,In_4882);
nor U1102 (N_1102,In_2582,In_3482);
nand U1103 (N_1103,In_2083,In_985);
and U1104 (N_1104,In_1898,In_2420);
and U1105 (N_1105,In_2939,In_488);
nor U1106 (N_1106,In_52,In_1950);
and U1107 (N_1107,In_2136,In_789);
xor U1108 (N_1108,In_3007,In_1196);
nand U1109 (N_1109,In_1615,In_3036);
nor U1110 (N_1110,In_1391,In_4564);
xor U1111 (N_1111,In_1837,In_4828);
nand U1112 (N_1112,In_3635,In_1354);
nor U1113 (N_1113,In_4962,In_2444);
or U1114 (N_1114,In_3853,In_4028);
nor U1115 (N_1115,In_4257,In_1687);
and U1116 (N_1116,In_703,In_3054);
nor U1117 (N_1117,In_1303,In_4441);
nor U1118 (N_1118,In_1355,In_551);
xor U1119 (N_1119,In_2773,In_1274);
nand U1120 (N_1120,In_2276,In_1234);
and U1121 (N_1121,In_403,In_3064);
xnor U1122 (N_1122,In_1398,In_4542);
xnor U1123 (N_1123,In_3911,In_2520);
and U1124 (N_1124,In_516,In_1546);
nand U1125 (N_1125,In_4285,In_2498);
xor U1126 (N_1126,In_1048,In_3273);
and U1127 (N_1127,In_4923,In_2518);
nand U1128 (N_1128,In_2731,In_674);
or U1129 (N_1129,In_2137,In_281);
and U1130 (N_1130,In_4823,In_2628);
and U1131 (N_1131,In_2817,In_1660);
and U1132 (N_1132,In_4728,In_183);
nand U1133 (N_1133,In_1011,In_4179);
or U1134 (N_1134,In_3067,In_1402);
nand U1135 (N_1135,In_1225,In_3795);
or U1136 (N_1136,In_3519,In_799);
or U1137 (N_1137,In_2769,In_4960);
nor U1138 (N_1138,In_1827,In_2170);
xor U1139 (N_1139,In_1641,In_101);
nor U1140 (N_1140,In_1823,In_4190);
and U1141 (N_1141,In_4381,In_4037);
xnor U1142 (N_1142,In_632,In_4254);
nor U1143 (N_1143,In_614,In_78);
and U1144 (N_1144,In_542,In_2499);
nand U1145 (N_1145,In_1671,In_986);
xnor U1146 (N_1146,In_3218,In_4684);
and U1147 (N_1147,In_1757,In_549);
nand U1148 (N_1148,In_4661,In_1392);
nand U1149 (N_1149,In_3181,In_861);
nor U1150 (N_1150,In_3708,In_2707);
nand U1151 (N_1151,In_968,In_2811);
xnor U1152 (N_1152,In_4586,In_4743);
xor U1153 (N_1153,In_908,In_766);
nor U1154 (N_1154,In_3372,In_4894);
xor U1155 (N_1155,In_1543,In_2150);
nor U1156 (N_1156,In_843,In_1621);
nor U1157 (N_1157,In_2277,In_993);
xor U1158 (N_1158,In_3158,In_170);
or U1159 (N_1159,In_3665,In_3258);
and U1160 (N_1160,In_177,In_3898);
nor U1161 (N_1161,In_1427,In_3854);
and U1162 (N_1162,In_803,In_1239);
xor U1163 (N_1163,In_512,In_3605);
and U1164 (N_1164,In_4399,In_3774);
or U1165 (N_1165,In_4059,In_3386);
xnor U1166 (N_1166,In_3000,In_606);
or U1167 (N_1167,In_3540,In_4788);
or U1168 (N_1168,In_4188,In_3068);
nor U1169 (N_1169,In_2931,In_4259);
and U1170 (N_1170,In_3601,In_4033);
nor U1171 (N_1171,In_1368,In_3919);
xor U1172 (N_1172,In_4761,In_4495);
or U1173 (N_1173,In_1872,In_1910);
and U1174 (N_1174,In_3765,In_4733);
and U1175 (N_1175,In_2254,In_4012);
and U1176 (N_1176,In_1681,In_4283);
nand U1177 (N_1177,In_4196,In_3356);
and U1178 (N_1178,In_4341,In_4484);
nand U1179 (N_1179,In_3235,In_1117);
xor U1180 (N_1180,In_541,In_2536);
nand U1181 (N_1181,In_1414,In_2234);
nand U1182 (N_1182,In_1496,In_3116);
nand U1183 (N_1183,In_4103,In_1304);
nor U1184 (N_1184,In_1017,In_4911);
nand U1185 (N_1185,In_3843,In_2605);
nor U1186 (N_1186,In_366,In_4101);
and U1187 (N_1187,In_2403,In_2937);
and U1188 (N_1188,In_1667,In_1360);
or U1189 (N_1189,In_1033,In_4562);
xor U1190 (N_1190,In_2469,In_1653);
nor U1191 (N_1191,In_2227,In_971);
or U1192 (N_1192,In_4559,In_2894);
and U1193 (N_1193,In_1477,In_367);
and U1194 (N_1194,In_1189,In_2720);
nand U1195 (N_1195,In_1087,In_1528);
xnor U1196 (N_1196,In_267,In_2450);
and U1197 (N_1197,In_517,In_1462);
or U1198 (N_1198,In_2231,In_2473);
nand U1199 (N_1199,In_820,In_4678);
or U1200 (N_1200,In_2189,In_743);
xor U1201 (N_1201,In_1899,In_1934);
nor U1202 (N_1202,In_969,In_4773);
and U1203 (N_1203,In_310,In_1588);
xor U1204 (N_1204,In_1600,In_2891);
or U1205 (N_1205,In_4740,In_2876);
or U1206 (N_1206,In_4063,In_362);
or U1207 (N_1207,In_4318,In_2036);
nor U1208 (N_1208,In_4278,In_4804);
or U1209 (N_1209,In_3016,In_3225);
and U1210 (N_1210,In_2597,In_2345);
nand U1211 (N_1211,In_679,In_4230);
xor U1212 (N_1212,In_4785,In_1086);
nand U1213 (N_1213,In_3182,In_97);
nor U1214 (N_1214,In_2835,In_3477);
and U1215 (N_1215,In_3330,In_1190);
or U1216 (N_1216,In_3219,In_3655);
nor U1217 (N_1217,In_2401,In_2019);
xnor U1218 (N_1218,In_1784,In_438);
nand U1219 (N_1219,In_2292,In_2432);
nand U1220 (N_1220,In_4374,In_1441);
or U1221 (N_1221,In_3673,In_2984);
or U1222 (N_1222,In_2020,In_4463);
or U1223 (N_1223,In_221,In_1410);
or U1224 (N_1224,In_3809,In_140);
and U1225 (N_1225,In_12,In_296);
xor U1226 (N_1226,In_212,In_2540);
nand U1227 (N_1227,In_1352,In_3178);
xor U1228 (N_1228,In_3968,In_839);
xor U1229 (N_1229,In_26,In_3797);
nor U1230 (N_1230,In_2783,In_3952);
nor U1231 (N_1231,In_1772,In_944);
xor U1232 (N_1232,In_1164,In_3532);
nand U1233 (N_1233,In_728,In_1078);
and U1234 (N_1234,In_286,In_2204);
xor U1235 (N_1235,In_2247,In_1069);
and U1236 (N_1236,In_306,In_1485);
and U1237 (N_1237,In_3745,In_414);
nor U1238 (N_1238,In_830,In_3286);
or U1239 (N_1239,In_3021,In_3552);
nor U1240 (N_1240,In_4723,In_2657);
nor U1241 (N_1241,In_1829,In_2193);
nand U1242 (N_1242,In_1271,In_3272);
nor U1243 (N_1243,In_3720,In_2887);
or U1244 (N_1244,In_3783,In_1617);
nor U1245 (N_1245,In_2938,In_3241);
xnor U1246 (N_1246,In_3735,In_1219);
and U1247 (N_1247,In_3302,In_3012);
nand U1248 (N_1248,In_4993,In_2506);
xor U1249 (N_1249,In_3890,In_2642);
and U1250 (N_1250,In_1853,In_3881);
and U1251 (N_1251,In_2397,In_3362);
or U1252 (N_1252,In_3129,In_437);
and U1253 (N_1253,In_755,In_4722);
and U1254 (N_1254,In_3088,In_4005);
nand U1255 (N_1255,In_3631,In_2065);
xor U1256 (N_1256,In_4597,In_4435);
nor U1257 (N_1257,In_17,In_4030);
nand U1258 (N_1258,In_4998,In_4050);
xor U1259 (N_1259,In_3217,In_2412);
and U1260 (N_1260,In_3342,In_1193);
and U1261 (N_1261,In_324,In_1677);
or U1262 (N_1262,In_3074,In_1921);
and U1263 (N_1263,In_3597,In_3037);
nor U1264 (N_1264,In_3363,In_1851);
nor U1265 (N_1265,In_379,In_3112);
or U1266 (N_1266,In_4194,In_1847);
and U1267 (N_1267,In_2378,In_1299);
and U1268 (N_1268,In_1946,In_3583);
or U1269 (N_1269,In_3508,In_3488);
or U1270 (N_1270,In_415,In_1399);
or U1271 (N_1271,In_863,In_4627);
nand U1272 (N_1272,In_4371,In_2107);
nor U1273 (N_1273,In_3415,In_4490);
xnor U1274 (N_1274,In_1916,In_4527);
or U1275 (N_1275,In_4637,In_1812);
nor U1276 (N_1276,In_3109,In_3814);
and U1277 (N_1277,In_4058,In_2725);
xor U1278 (N_1278,In_4475,In_1218);
xor U1279 (N_1279,In_1466,In_3081);
or U1280 (N_1280,In_2347,In_3988);
nand U1281 (N_1281,In_187,In_574);
and U1282 (N_1282,In_3395,In_4372);
nor U1283 (N_1283,In_2090,In_4909);
nand U1284 (N_1284,In_4805,In_4918);
or U1285 (N_1285,In_149,In_4499);
xor U1286 (N_1286,In_1151,In_4875);
nand U1287 (N_1287,In_3123,In_2729);
or U1288 (N_1288,In_4534,In_3562);
nor U1289 (N_1289,In_1803,In_2952);
and U1290 (N_1290,In_3693,In_4388);
or U1291 (N_1291,In_4219,In_3925);
nand U1292 (N_1292,In_4149,In_3563);
nand U1293 (N_1293,In_4335,In_233);
nor U1294 (N_1294,In_2084,In_2617);
nor U1295 (N_1295,In_3915,In_3619);
xor U1296 (N_1296,In_1110,In_60);
xor U1297 (N_1297,In_1067,In_4200);
nand U1298 (N_1298,In_4119,In_4223);
and U1299 (N_1299,In_1931,In_3500);
nand U1300 (N_1300,In_4618,In_215);
or U1301 (N_1301,In_4863,In_4243);
xor U1302 (N_1302,In_2611,In_2324);
or U1303 (N_1303,In_3333,In_321);
xor U1304 (N_1304,In_19,In_3752);
and U1305 (N_1305,In_4045,In_133);
xor U1306 (N_1306,In_4906,In_4707);
nor U1307 (N_1307,In_3419,In_4734);
or U1308 (N_1308,In_3577,In_2505);
xor U1309 (N_1309,In_2845,In_2631);
xor U1310 (N_1310,In_534,In_4585);
nand U1311 (N_1311,In_2743,In_3689);
and U1312 (N_1312,In_4806,In_4575);
nand U1313 (N_1313,In_3966,In_3263);
xnor U1314 (N_1314,In_682,In_2547);
or U1315 (N_1315,In_4818,In_4750);
xor U1316 (N_1316,In_2027,In_4502);
or U1317 (N_1317,In_1207,In_4465);
and U1318 (N_1318,In_2554,In_1809);
xnor U1319 (N_1319,In_401,In_2390);
xor U1320 (N_1320,In_3525,In_2223);
nor U1321 (N_1321,In_4228,In_4507);
nor U1322 (N_1322,In_2264,In_2844);
nor U1323 (N_1323,In_1495,In_404);
or U1324 (N_1324,In_3944,In_3001);
nor U1325 (N_1325,In_2471,In_3652);
nor U1326 (N_1326,In_2311,In_695);
nor U1327 (N_1327,In_2892,In_4431);
nor U1328 (N_1328,In_4319,In_3458);
nand U1329 (N_1329,In_2955,In_1475);
xnor U1330 (N_1330,In_1176,In_3938);
and U1331 (N_1331,In_346,In_491);
nand U1332 (N_1332,In_2055,In_4541);
and U1333 (N_1333,In_2089,In_1236);
nand U1334 (N_1334,In_2551,In_3073);
nor U1335 (N_1335,In_2590,In_657);
nor U1336 (N_1336,In_4191,In_3590);
xor U1337 (N_1337,In_4066,In_2816);
xor U1338 (N_1338,In_2031,In_4532);
nand U1339 (N_1339,In_3305,In_724);
xor U1340 (N_1340,In_3369,In_3826);
nand U1341 (N_1341,In_2545,In_4376);
xnor U1342 (N_1342,In_1012,In_2046);
nand U1343 (N_1343,In_3069,In_1345);
nand U1344 (N_1344,In_896,In_3747);
and U1345 (N_1345,In_1286,In_4284);
nor U1346 (N_1346,In_3859,In_3341);
xnor U1347 (N_1347,In_3097,In_2514);
xnor U1348 (N_1348,In_2272,In_3390);
and U1349 (N_1349,In_1786,In_2581);
nand U1350 (N_1350,In_3626,In_2451);
and U1351 (N_1351,In_666,In_76);
nand U1352 (N_1352,In_912,In_2286);
xor U1353 (N_1353,In_2109,In_1138);
and U1354 (N_1354,In_1532,In_3484);
nand U1355 (N_1355,In_3917,In_4944);
and U1356 (N_1356,In_1492,In_168);
and U1357 (N_1357,In_3264,In_3367);
and U1358 (N_1358,In_2548,In_2741);
or U1359 (N_1359,In_936,In_1487);
xor U1360 (N_1360,In_4187,In_3147);
xnor U1361 (N_1361,In_2496,In_3149);
or U1362 (N_1362,In_1120,In_1936);
xor U1363 (N_1363,In_1856,In_1777);
xor U1364 (N_1364,In_4365,In_4470);
and U1365 (N_1365,In_4834,In_4140);
and U1366 (N_1366,In_460,In_3691);
nand U1367 (N_1367,In_811,In_45);
xnor U1368 (N_1368,In_4543,In_3904);
or U1369 (N_1369,In_291,In_4710);
and U1370 (N_1370,In_1944,In_4053);
and U1371 (N_1371,In_3211,In_3501);
xor U1372 (N_1372,In_2993,In_2658);
and U1373 (N_1373,In_2535,In_2001);
xor U1374 (N_1374,In_4510,In_596);
nor U1375 (N_1375,In_4695,In_961);
xnor U1376 (N_1376,In_3860,In_4531);
or U1377 (N_1377,In_2527,In_3868);
nor U1378 (N_1378,In_1209,In_2689);
or U1379 (N_1379,In_4687,In_3861);
nand U1380 (N_1380,In_2054,In_3124);
xor U1381 (N_1381,In_1562,In_3017);
xnor U1382 (N_1382,In_3950,In_1724);
nand U1383 (N_1383,In_2242,In_1605);
nor U1384 (N_1384,In_1789,In_1080);
nor U1385 (N_1385,In_4430,In_4092);
or U1386 (N_1386,In_4506,In_2641);
nor U1387 (N_1387,In_2651,In_91);
nand U1388 (N_1388,In_844,In_3549);
xor U1389 (N_1389,In_2317,In_4821);
nor U1390 (N_1390,In_1876,In_444);
nor U1391 (N_1391,In_626,In_1658);
nor U1392 (N_1392,In_1265,In_2708);
xor U1393 (N_1393,In_4300,In_3326);
or U1394 (N_1394,In_4,In_2165);
xnor U1395 (N_1395,In_2749,In_4448);
or U1396 (N_1396,In_4221,In_4236);
nor U1397 (N_1397,In_4240,In_2402);
nor U1398 (N_1398,In_2790,In_4752);
nor U1399 (N_1399,In_13,In_3699);
nor U1400 (N_1400,In_4246,In_2982);
nand U1401 (N_1401,In_445,In_489);
and U1402 (N_1402,In_729,In_3254);
xnor U1403 (N_1403,In_4270,In_2830);
nand U1404 (N_1404,In_2134,In_3620);
xor U1405 (N_1405,In_675,In_3586);
or U1406 (N_1406,In_797,In_1663);
or U1407 (N_1407,In_2511,In_271);
xnor U1408 (N_1408,In_3806,In_2418);
or U1409 (N_1409,In_122,In_4253);
nor U1410 (N_1410,In_2275,In_4295);
or U1411 (N_1411,In_1904,In_777);
xor U1412 (N_1412,In_4691,In_2751);
and U1413 (N_1413,In_2256,In_1397);
and U1414 (N_1414,In_700,In_2574);
nor U1415 (N_1415,In_4476,In_186);
xnor U1416 (N_1416,In_4945,In_573);
nor U1417 (N_1417,In_3751,In_1287);
nand U1418 (N_1418,In_4566,In_3970);
nor U1419 (N_1419,In_2178,In_1464);
or U1420 (N_1420,In_3895,In_4775);
or U1421 (N_1421,In_648,In_24);
or U1422 (N_1422,In_1257,In_3318);
xnor U1423 (N_1423,In_4129,In_3954);
nand U1424 (N_1424,In_778,In_659);
nand U1425 (N_1425,In_3939,In_1445);
nand U1426 (N_1426,In_1417,In_2814);
nand U1427 (N_1427,In_383,In_4501);
and U1428 (N_1428,In_772,In_3425);
xnor U1429 (N_1429,In_3204,In_203);
nor U1430 (N_1430,In_586,In_4694);
xnor U1431 (N_1431,In_4354,In_1795);
xor U1432 (N_1432,In_4301,In_2082);
and U1433 (N_1433,In_160,In_2099);
nand U1434 (N_1434,In_4957,In_4177);
nand U1435 (N_1435,In_1519,In_417);
or U1436 (N_1436,In_2284,In_2388);
and U1437 (N_1437,In_1826,In_1002);
and U1438 (N_1438,In_4094,In_2638);
or U1439 (N_1439,In_2,In_1554);
or U1440 (N_1440,In_361,In_3771);
or U1441 (N_1441,In_4669,In_2665);
nor U1442 (N_1442,In_4077,In_1729);
nand U1443 (N_1443,In_3922,In_355);
nor U1444 (N_1444,In_1764,In_1378);
nand U1445 (N_1445,In_526,In_4109);
nand U1446 (N_1446,In_2704,In_3233);
nor U1447 (N_1447,In_1367,In_110);
and U1448 (N_1448,In_181,In_1720);
nand U1449 (N_1449,In_4387,In_1850);
or U1450 (N_1450,In_2446,In_1411);
nand U1451 (N_1451,In_1717,In_710);
nand U1452 (N_1452,In_1735,In_2239);
and U1453 (N_1453,In_3015,In_3379);
nand U1454 (N_1454,In_3574,In_2809);
nand U1455 (N_1455,In_2288,In_4181);
xor U1456 (N_1456,In_2637,In_4866);
nand U1457 (N_1457,In_1113,In_1715);
and U1458 (N_1458,In_2050,In_4108);
xor U1459 (N_1459,In_4552,In_2805);
or U1460 (N_1460,In_748,In_4557);
or U1461 (N_1461,In_498,In_524);
nor U1462 (N_1462,In_3817,In_697);
and U1463 (N_1463,In_4520,In_4158);
nand U1464 (N_1464,In_3588,In_249);
xnor U1465 (N_1465,In_3403,In_3600);
and U1466 (N_1466,In_1919,In_3480);
xor U1467 (N_1467,In_1131,In_2745);
nand U1468 (N_1468,In_1622,In_3628);
nor U1469 (N_1469,In_3528,In_2676);
nand U1470 (N_1470,In_2613,In_2263);
and U1471 (N_1471,In_1640,In_2447);
nor U1472 (N_1472,In_507,In_1857);
or U1473 (N_1473,In_619,In_859);
and U1474 (N_1474,In_4329,In_855);
nor U1475 (N_1475,In_3255,In_3232);
or U1476 (N_1476,In_1710,In_1815);
or U1477 (N_1477,In_30,In_2996);
and U1478 (N_1478,In_3259,In_198);
nor U1479 (N_1479,In_4110,In_3686);
nor U1480 (N_1480,In_4350,In_4849);
and U1481 (N_1481,In_2591,In_1561);
nor U1482 (N_1482,In_2123,In_44);
or U1483 (N_1483,In_231,In_2619);
nand U1484 (N_1484,In_390,In_2562);
xnor U1485 (N_1485,In_1801,In_2750);
nand U1486 (N_1486,In_3435,In_1566);
nor U1487 (N_1487,In_1603,In_4014);
or U1488 (N_1488,In_4296,In_3596);
nand U1489 (N_1489,In_2798,In_1967);
or U1490 (N_1490,In_125,In_273);
nor U1491 (N_1491,In_349,In_525);
nor U1492 (N_1492,In_1606,In_4994);
nor U1493 (N_1493,In_775,In_1314);
nand U1494 (N_1494,In_2956,In_1707);
nand U1495 (N_1495,In_1650,In_991);
xor U1496 (N_1496,In_3119,In_2490);
xor U1497 (N_1497,In_4980,In_1137);
or U1498 (N_1498,In_792,In_946);
or U1499 (N_1499,In_1124,In_3370);
and U1500 (N_1500,In_2855,In_3866);
xnor U1501 (N_1501,In_1007,In_3420);
nor U1502 (N_1502,In_4405,In_56);
nand U1503 (N_1503,In_3191,In_1747);
nand U1504 (N_1504,In_1429,In_495);
xor U1505 (N_1505,In_340,In_878);
nand U1506 (N_1506,In_860,In_2301);
and U1507 (N_1507,In_1981,In_4437);
xor U1508 (N_1508,In_2114,In_3010);
and U1509 (N_1509,In_1072,In_407);
nand U1510 (N_1510,In_3467,In_1159);
nand U1511 (N_1511,In_3700,In_2950);
nand U1512 (N_1512,In_3079,In_2190);
nor U1513 (N_1513,In_1766,In_4171);
nor U1514 (N_1514,In_4197,In_3551);
xor U1515 (N_1515,In_3298,In_1186);
and U1516 (N_1516,In_4264,In_1573);
or U1517 (N_1517,In_1167,In_4439);
nand U1518 (N_1518,In_3906,In_4539);
and U1519 (N_1519,In_1821,In_2093);
and U1520 (N_1520,In_2208,In_638);
nand U1521 (N_1521,In_727,In_4789);
nand U1522 (N_1522,In_2240,In_1374);
nand U1523 (N_1523,In_4176,In_3841);
nor U1524 (N_1524,In_4220,In_4481);
nor U1525 (N_1525,In_3424,In_4162);
nand U1526 (N_1526,In_1769,In_4118);
nor U1527 (N_1527,In_584,In_3976);
nand U1528 (N_1528,In_3749,In_939);
and U1529 (N_1529,In_3157,In_497);
or U1530 (N_1530,In_1336,In_4410);
xnor U1531 (N_1531,In_3971,In_4204);
nor U1532 (N_1532,In_1527,In_1093);
nor U1533 (N_1533,In_3214,In_433);
nor U1534 (N_1534,In_623,In_4831);
nor U1535 (N_1535,In_2492,In_4645);
xor U1536 (N_1536,In_2321,In_1989);
nand U1537 (N_1537,In_3715,In_1316);
and U1538 (N_1538,In_256,In_4471);
and U1539 (N_1539,In_2810,In_408);
xnor U1540 (N_1540,In_1558,In_397);
nand U1541 (N_1541,In_3060,In_1711);
xor U1542 (N_1542,In_1361,In_805);
xnor U1543 (N_1543,In_1288,In_3378);
and U1544 (N_1544,In_1572,In_1938);
or U1545 (N_1545,In_1165,In_3041);
or U1546 (N_1546,In_1586,In_1848);
nor U1547 (N_1547,In_137,In_3499);
xor U1548 (N_1548,In_745,In_725);
nor U1549 (N_1549,In_2850,In_1782);
nor U1550 (N_1550,In_1922,In_1156);
xnor U1551 (N_1551,In_3694,In_2672);
xnor U1552 (N_1552,In_1041,In_1440);
nor U1553 (N_1553,In_3999,In_2489);
or U1554 (N_1554,In_3951,In_4444);
and U1555 (N_1555,In_4292,In_4105);
nor U1556 (N_1556,In_1266,In_1843);
xnor U1557 (N_1557,In_4425,In_1289);
nand U1558 (N_1558,In_2487,In_3492);
and U1559 (N_1559,In_3784,In_1122);
and U1560 (N_1560,In_1247,In_3770);
and U1561 (N_1561,In_2504,In_4207);
or U1562 (N_1562,In_1281,In_2462);
xnor U1563 (N_1563,In_2964,In_979);
or U1564 (N_1564,In_4087,In_794);
nand U1565 (N_1565,In_1199,In_3319);
and U1566 (N_1566,In_2776,In_4985);
xnor U1567 (N_1567,In_1419,In_3873);
xnor U1568 (N_1568,In_796,In_2061);
nand U1569 (N_1569,In_2649,In_1995);
or U1570 (N_1570,In_3144,In_4932);
xor U1571 (N_1571,In_3664,In_342);
or U1572 (N_1572,In_2187,In_1081);
xnor U1573 (N_1573,In_2744,In_3616);
or U1574 (N_1574,In_3512,In_4488);
xor U1575 (N_1575,In_874,In_225);
xnor U1576 (N_1576,In_1065,In_1365);
and U1577 (N_1577,In_3572,In_1129);
or U1578 (N_1578,In_4646,In_4610);
and U1579 (N_1579,In_429,In_2396);
xnor U1580 (N_1580,In_284,In_3270);
nand U1581 (N_1581,In_2259,In_2376);
or U1582 (N_1582,In_4760,In_1911);
or U1583 (N_1583,In_3518,In_259);
nor U1584 (N_1584,In_1135,In_67);
nand U1585 (N_1585,In_1261,In_1071);
or U1586 (N_1586,In_2502,In_1371);
and U1587 (N_1587,In_1822,In_1962);
and U1588 (N_1588,In_1984,In_4626);
xor U1589 (N_1589,In_4096,In_2460);
or U1590 (N_1590,In_3153,In_3239);
nand U1591 (N_1591,In_3636,In_1061);
nand U1592 (N_1592,In_688,In_1305);
and U1593 (N_1593,In_66,In_2667);
and U1594 (N_1594,In_3162,In_883);
nor U1595 (N_1595,In_3042,In_1191);
nand U1596 (N_1596,In_4251,In_3437);
nand U1597 (N_1597,In_37,In_209);
or U1598 (N_1598,In_1808,In_1243);
nor U1599 (N_1599,In_3268,In_914);
or U1600 (N_1600,In_1597,In_2653);
nor U1601 (N_1601,In_1734,In_2555);
and U1602 (N_1602,In_2914,In_1077);
or U1603 (N_1603,In_875,In_4287);
xnor U1604 (N_1604,In_3213,In_4322);
or U1605 (N_1605,In_2737,In_128);
xor U1606 (N_1606,In_2868,In_335);
xor U1607 (N_1607,In_108,In_238);
nor U1608 (N_1608,In_3065,In_532);
xnor U1609 (N_1609,In_27,In_3391);
and U1610 (N_1610,In_232,In_2953);
or U1611 (N_1611,In_2228,In_428);
or U1612 (N_1612,In_3702,In_1966);
nor U1613 (N_1613,In_3184,In_3542);
nand U1614 (N_1614,In_4057,In_3942);
and U1615 (N_1615,In_95,In_3835);
xnor U1616 (N_1616,In_3623,In_1249);
nand U1617 (N_1617,In_2948,In_4802);
xnor U1618 (N_1618,In_3796,In_161);
nor U1619 (N_1619,In_2294,In_3022);
nor U1620 (N_1620,In_2186,In_2917);
nor U1621 (N_1621,In_2118,In_2465);
nand U1622 (N_1622,In_2414,In_131);
and U1623 (N_1623,In_1197,In_3327);
nand U1624 (N_1624,In_2245,In_2603);
xor U1625 (N_1625,In_1979,In_4205);
and U1626 (N_1626,In_822,In_558);
xor U1627 (N_1627,In_4137,In_1455);
xor U1628 (N_1628,In_1382,In_3078);
xnor U1629 (N_1629,In_3617,In_1014);
xor U1630 (N_1630,In_338,In_4269);
and U1631 (N_1631,In_1889,In_2184);
nand U1632 (N_1632,In_3821,In_4915);
nand U1633 (N_1633,In_2179,In_4820);
or U1634 (N_1634,In_4671,In_1673);
nand U1635 (N_1635,In_1659,In_2701);
xor U1636 (N_1636,In_535,In_2864);
nor U1637 (N_1637,In_4474,In_3295);
and U1638 (N_1638,In_2377,In_2370);
or U1639 (N_1639,In_4650,In_3353);
nor U1640 (N_1640,In_840,In_1800);
xnor U1641 (N_1641,In_3253,In_3024);
or U1642 (N_1642,In_4001,In_1680);
or U1643 (N_1643,In_1128,In_2570);
nand U1644 (N_1644,In_1541,In_2791);
nand U1645 (N_1645,In_4967,In_82);
or U1646 (N_1646,In_1152,In_2974);
nand U1647 (N_1647,In_247,In_2098);
xor U1648 (N_1648,In_86,In_4582);
xor U1649 (N_1649,In_4464,In_2171);
xnor U1650 (N_1650,In_1499,In_3384);
and U1651 (N_1651,In_2115,In_2529);
xnor U1652 (N_1652,In_2947,In_2739);
nand U1653 (N_1653,In_3351,In_4184);
and U1654 (N_1654,In_3280,In_2222);
and U1655 (N_1655,In_4937,In_4976);
nand U1656 (N_1656,In_1908,In_2062);
nand U1657 (N_1657,In_1678,In_2112);
nand U1658 (N_1658,In_3548,In_635);
or U1659 (N_1659,In_4174,In_4447);
xor U1660 (N_1660,In_317,In_4780);
or U1661 (N_1661,In_4572,In_3612);
nor U1662 (N_1662,In_4922,In_1161);
xnor U1663 (N_1663,In_4392,In_1223);
nor U1664 (N_1664,In_1262,In_3006);
and U1665 (N_1665,In_1282,In_3417);
nor U1666 (N_1666,In_4889,In_644);
nor U1667 (N_1667,In_2497,In_288);
and U1668 (N_1668,In_3076,In_2435);
and U1669 (N_1669,In_3983,In_2142);
nand U1670 (N_1670,In_1023,In_326);
or U1671 (N_1671,In_762,In_2406);
xor U1672 (N_1672,In_2140,In_3430);
nor U1673 (N_1673,In_3175,In_4062);
nand U1674 (N_1674,In_1277,In_3176);
or U1675 (N_1675,In_3434,In_633);
or U1676 (N_1676,In_2732,In_3820);
nor U1677 (N_1677,In_3993,In_4846);
xnor U1678 (N_1678,In_998,In_4767);
or U1679 (N_1679,In_1522,In_582);
xnor U1680 (N_1680,In_4206,In_4272);
and U1681 (N_1681,In_801,In_953);
or U1682 (N_1682,In_1335,In_3209);
or U1683 (N_1683,In_3530,In_246);
nor U1684 (N_1684,In_1767,In_2008);
nand U1685 (N_1685,In_2692,In_1636);
xor U1686 (N_1686,In_1066,In_1531);
and U1687 (N_1687,In_3887,In_2593);
and U1688 (N_1688,In_4247,In_1387);
or U1689 (N_1689,In_3878,In_1506);
nor U1690 (N_1690,In_3143,In_402);
or U1691 (N_1691,In_4772,In_3085);
and U1692 (N_1692,In_2594,In_2859);
nand U1693 (N_1693,In_100,In_972);
or U1694 (N_1694,In_490,In_1625);
or U1695 (N_1695,In_1016,In_915);
or U1696 (N_1696,In_4031,In_2588);
xnor U1697 (N_1697,In_2843,In_806);
nor U1698 (N_1698,In_3156,In_4924);
and U1699 (N_1699,In_1828,In_2975);
and U1700 (N_1700,In_4977,In_2659);
nand U1701 (N_1701,In_1863,In_1404);
nand U1702 (N_1702,In_1394,In_1507);
nor U1703 (N_1703,In_3837,In_3479);
and U1704 (N_1704,In_2167,In_4724);
or U1705 (N_1705,In_1230,In_1141);
nor U1706 (N_1706,In_787,In_4321);
nand U1707 (N_1707,In_515,In_4156);
or U1708 (N_1708,In_3786,In_3757);
nand U1709 (N_1709,In_978,In_4222);
nor U1710 (N_1710,In_4668,In_4074);
nand U1711 (N_1711,In_3594,In_952);
nor U1712 (N_1712,In_1085,In_4854);
xor U1713 (N_1713,In_1172,In_587);
nand U1714 (N_1714,In_3324,In_1450);
and U1715 (N_1715,In_1005,In_1329);
or U1716 (N_1716,In_1762,In_4500);
or U1717 (N_1717,In_4093,In_1601);
and U1718 (N_1718,In_4550,In_3221);
and U1719 (N_1719,In_4856,In_3350);
nor U1720 (N_1720,In_3627,In_2169);
or U1721 (N_1721,In_4323,In_2229);
and U1722 (N_1722,In_4347,In_2997);
nor U1723 (N_1723,In_3908,In_139);
and U1724 (N_1724,In_434,In_3876);
xor U1725 (N_1725,In_2909,In_2604);
or U1726 (N_1726,In_2135,In_639);
nand U1727 (N_1727,In_3338,In_468);
and U1728 (N_1728,In_3793,In_4721);
xor U1729 (N_1729,In_1025,In_2327);
or U1730 (N_1730,In_303,In_4600);
xnor U1731 (N_1731,In_3148,In_4605);
xnor U1732 (N_1732,In_4928,In_3801);
and U1733 (N_1733,In_3445,In_1841);
nor U1734 (N_1734,In_1954,In_2122);
xnor U1735 (N_1735,In_690,In_4825);
xor U1736 (N_1736,In_4339,In_4881);
xnor U1737 (N_1737,In_1608,In_2032);
nand U1738 (N_1738,In_1701,In_4801);
and U1739 (N_1739,In_537,In_645);
and U1740 (N_1740,In_3914,In_3361);
nor U1741 (N_1741,In_2967,In_1437);
or U1742 (N_1742,In_3845,In_3524);
nand U1743 (N_1743,In_4489,In_834);
or U1744 (N_1744,In_4730,In_1758);
xnor U1745 (N_1745,In_4517,In_3943);
or U1746 (N_1746,In_4232,In_72);
or U1747 (N_1747,In_1366,In_4978);
nor U1748 (N_1748,In_471,In_715);
xor U1749 (N_1749,In_4857,In_3252);
nor U1750 (N_1750,In_1309,In_2173);
and U1751 (N_1751,In_94,In_583);
or U1752 (N_1752,In_2710,In_613);
xnor U1753 (N_1753,In_1075,In_4568);
xnor U1754 (N_1754,In_4345,In_2841);
and U1755 (N_1755,In_3283,In_1216);
nor U1756 (N_1756,In_3580,In_4503);
xor U1757 (N_1757,In_2318,In_3565);
nand U1758 (N_1758,In_2706,In_4305);
nand U1759 (N_1759,In_1568,In_1688);
or U1760 (N_1760,In_3935,In_4203);
nor U1761 (N_1761,In_563,In_4748);
and U1762 (N_1762,In_1363,In_4391);
or U1763 (N_1763,In_15,In_4812);
nand U1764 (N_1764,In_2670,In_4861);
nand U1765 (N_1765,In_1251,In_3818);
xnor U1766 (N_1766,In_1556,In_3931);
nand U1767 (N_1767,In_884,In_2620);
xnor U1768 (N_1768,In_159,In_3439);
xnor U1769 (N_1769,In_2679,In_106);
xnor U1770 (N_1770,In_601,In_1240);
nor U1771 (N_1771,In_3180,In_3474);
xor U1772 (N_1772,In_2394,In_1433);
or U1773 (N_1773,In_4898,In_4623);
and U1774 (N_1774,In_1489,In_2766);
and U1775 (N_1775,In_4480,In_1242);
nand U1776 (N_1776,In_2197,In_1490);
xnor U1777 (N_1777,In_1112,In_4660);
and U1778 (N_1778,In_85,In_446);
nor U1779 (N_1779,In_3459,In_4590);
nand U1780 (N_1780,In_33,In_4231);
and U1781 (N_1781,In_1865,In_3696);
and U1782 (N_1782,In_3203,In_3423);
xor U1783 (N_1783,In_2934,In_867);
nor U1784 (N_1784,In_4638,In_1162);
nand U1785 (N_1785,In_4725,In_4198);
nand U1786 (N_1786,In_228,In_1947);
and U1787 (N_1787,In_3466,In_1565);
and U1788 (N_1788,In_3790,In_3816);
nor U1789 (N_1789,In_3805,In_1505);
nor U1790 (N_1790,In_2525,In_1254);
or U1791 (N_1791,In_2040,In_4596);
nor U1792 (N_1792,In_469,In_463);
or U1793 (N_1793,In_547,In_4642);
or U1794 (N_1794,In_4421,In_2243);
nor U1795 (N_1795,In_1798,In_4199);
and U1796 (N_1796,In_1150,In_378);
nor U1797 (N_1797,In_282,In_624);
or U1798 (N_1798,In_2712,In_2209);
or U1799 (N_1799,In_1070,In_466);
nand U1800 (N_1800,In_3311,In_4245);
xnor U1801 (N_1801,In_1890,In_2013);
and U1802 (N_1802,In_3692,In_2669);
nor U1803 (N_1803,In_3448,In_2417);
nor U1804 (N_1804,In_4302,In_1003);
and U1805 (N_1805,In_2893,In_530);
nor U1806 (N_1806,In_3946,In_4102);
xnor U1807 (N_1807,In_2663,In_795);
xnor U1808 (N_1808,In_2077,In_2647);
and U1809 (N_1809,In_1624,In_2763);
xnor U1810 (N_1810,In_3404,In_3857);
nand U1811 (N_1811,In_34,In_3962);
or U1812 (N_1812,In_1409,In_4879);
xor U1813 (N_1813,In_4908,In_687);
or U1814 (N_1814,In_1307,In_3023);
or U1815 (N_1815,In_1712,In_2946);
and U1816 (N_1816,In_4770,In_4698);
nand U1817 (N_1817,In_2800,In_4288);
nand U1818 (N_1818,In_1079,In_2104);
or U1819 (N_1819,In_4237,In_2792);
or U1820 (N_1820,In_767,In_1632);
xor U1821 (N_1821,In_74,In_155);
nand U1822 (N_1822,In_333,In_4104);
or U1823 (N_1823,In_3902,In_2988);
and U1824 (N_1824,In_418,In_705);
and U1825 (N_1825,In_3905,In_4602);
and U1826 (N_1826,In_2508,In_1963);
and U1827 (N_1827,In_3025,In_146);
xor U1828 (N_1828,In_1260,In_1634);
or U1829 (N_1829,In_4061,In_1126);
nor U1830 (N_1830,In_3278,In_4336);
xor U1831 (N_1831,In_3,In_3237);
and U1832 (N_1832,In_4462,In_4958);
xnor U1833 (N_1833,In_3874,In_3679);
nand U1834 (N_1834,In_4106,In_4914);
nor U1835 (N_1835,In_658,In_1604);
xor U1836 (N_1836,In_4756,In_4709);
xor U1837 (N_1837,In_3495,In_4519);
or U1838 (N_1838,In_2028,In_3743);
xor U1839 (N_1839,In_4485,In_1877);
and U1840 (N_1840,In_4310,In_678);
or U1841 (N_1841,In_457,In_2443);
nor U1842 (N_1842,In_3202,In_4604);
or U1843 (N_1843,In_2740,In_4000);
nand U1844 (N_1844,In_550,In_1279);
and U1845 (N_1845,In_1478,In_3930);
nor U1846 (N_1846,In_4487,In_4290);
xor U1847 (N_1847,In_2219,In_2439);
and U1848 (N_1848,In_4648,In_2081);
xor U1849 (N_1849,In_3659,In_4931);
nand U1850 (N_1850,In_3349,In_197);
nor U1851 (N_1851,In_1993,In_2500);
nor U1852 (N_1852,In_4282,In_2453);
xnor U1853 (N_1853,In_4019,In_2902);
nor U1854 (N_1854,In_4326,In_1428);
xnor U1855 (N_1855,In_627,In_739);
nor U1856 (N_1856,In_4631,In_3858);
and U1857 (N_1857,In_4446,In_588);
xnor U1858 (N_1858,In_1915,In_1578);
nand U1859 (N_1859,In_115,In_917);
nor U1860 (N_1860,In_2501,In_3851);
and U1861 (N_1861,In_2774,In_3045);
xnor U1862 (N_1862,In_1396,In_3669);
xor U1863 (N_1863,In_486,In_780);
nor U1864 (N_1864,In_812,In_2618);
nand U1865 (N_1865,In_4664,In_4357);
nand U1866 (N_1866,In_4987,In_1105);
or U1867 (N_1867,In_1263,In_3990);
xor U1868 (N_1868,In_999,In_1130);
nor U1869 (N_1869,In_2579,In_3171);
xor U1870 (N_1870,In_2185,In_4128);
nand U1871 (N_1871,In_1644,In_2060);
and U1872 (N_1872,In_325,In_504);
or U1873 (N_1873,In_4211,In_3606);
and U1874 (N_1874,In_2059,In_1372);
or U1875 (N_1875,In_4936,In_3891);
or U1876 (N_1876,In_2796,In_4164);
and U1877 (N_1877,In_4135,In_3787);
xnor U1878 (N_1878,In_4034,In_2852);
xor U1879 (N_1879,In_223,In_1840);
xor U1880 (N_1880,In_513,In_370);
nor U1881 (N_1881,In_2160,In_3723);
and U1882 (N_1882,In_1010,In_4555);
or U1883 (N_1883,In_1788,In_278);
nor U1884 (N_1884,In_1201,In_4702);
and U1885 (N_1885,In_585,In_1781);
or U1886 (N_1886,In_3072,In_1730);
xnor U1887 (N_1887,In_4038,In_3624);
or U1888 (N_1888,In_1727,In_4256);
nor U1889 (N_1889,In_1310,In_175);
and U1890 (N_1890,In_4003,In_4225);
xor U1891 (N_1891,In_2454,In_4674);
nor U1892 (N_1892,In_4912,In_432);
or U1893 (N_1893,In_360,In_2926);
xnor U1894 (N_1894,In_3426,In_1917);
nand U1895 (N_1895,In_2930,In_2987);
xor U1896 (N_1896,In_3648,In_399);
nand U1897 (N_1897,In_1939,In_4395);
nor U1898 (N_1898,In_462,In_1612);
nand U1899 (N_1899,In_487,In_87);
xor U1900 (N_1900,In_3509,In_2043);
xnor U1901 (N_1901,In_508,In_2285);
or U1902 (N_1902,In_1778,In_2869);
or U1903 (N_1903,In_2904,In_4966);
or U1904 (N_1904,In_1498,In_615);
nor U1905 (N_1905,In_4337,In_1854);
xor U1906 (N_1906,In_3220,In_3807);
or U1907 (N_1907,In_25,In_3366);
nand U1908 (N_1908,In_617,In_1182);
nor U1909 (N_1909,In_4035,In_3738);
nor U1910 (N_1910,In_2094,In_57);
nor U1911 (N_1911,In_2026,In_4968);
and U1912 (N_1912,In_1063,In_2920);
nor U1913 (N_1913,In_3557,In_1756);
and U1914 (N_1914,In_1894,In_4822);
and U1915 (N_1915,In_1210,In_1178);
nor U1916 (N_1916,In_2342,In_3321);
nand U1917 (N_1917,In_4460,In_4233);
nor U1918 (N_1918,In_977,In_3564);
nor U1919 (N_1919,In_790,In_3553);
nor U1920 (N_1920,In_1593,In_2073);
xor U1921 (N_1921,In_1395,In_2359);
nor U1922 (N_1922,In_2754,In_4144);
nand U1923 (N_1923,In_630,In_4307);
and U1924 (N_1924,In_4052,In_4172);
xor U1925 (N_1925,In_667,In_2734);
or U1926 (N_1926,In_3452,In_1454);
nand U1927 (N_1927,In_3556,In_263);
and U1928 (N_1928,In_250,In_207);
nand U1929 (N_1929,In_3681,In_3094);
or U1930 (N_1930,In_1035,In_1060);
nand U1931 (N_1931,In_2248,In_4560);
xor U1932 (N_1932,In_980,In_1670);
xnor U1933 (N_1933,In_4353,In_4905);
and U1934 (N_1934,In_1852,In_3496);
or U1935 (N_1935,In_3913,In_3034);
or U1936 (N_1936,In_292,In_1153);
nor U1937 (N_1937,In_3447,In_3475);
nor U1938 (N_1938,In_4136,In_3397);
or U1939 (N_1939,In_4385,In_1831);
nor U1940 (N_1940,In_2309,In_2362);
or U1941 (N_1941,In_2794,In_1986);
nor U1942 (N_1942,In_3989,In_4938);
nor U1943 (N_1943,In_1516,In_4904);
nand U1944 (N_1944,In_328,In_4436);
or U1945 (N_1945,In_744,In_758);
or U1946 (N_1946,In_2310,In_975);
xor U1947 (N_1947,In_4328,In_2788);
or U1948 (N_1948,In_4483,In_2509);
and U1949 (N_1949,In_21,In_2577);
xnor U1950 (N_1950,In_4608,In_3090);
nor U1951 (N_1951,In_3704,In_4584);
xnor U1952 (N_1952,In_3084,In_1974);
xnor U1953 (N_1953,In_1814,In_2354);
nor U1954 (N_1954,In_2066,In_888);
nand U1955 (N_1955,In_2230,In_1001);
xnor U1956 (N_1956,In_356,In_2244);
xor U1957 (N_1957,In_1751,In_62);
nor U1958 (N_1958,In_4011,In_4629);
or U1959 (N_1959,In_2980,In_4208);
nor U1960 (N_1960,In_607,In_214);
nand U1961 (N_1961,In_670,In_1);
or U1962 (N_1962,In_1695,In_3050);
xnor U1963 (N_1963,In_2379,In_2596);
and U1964 (N_1964,In_1426,In_136);
nand U1965 (N_1965,In_1147,In_4150);
nor U1966 (N_1966,In_4565,In_2218);
or U1967 (N_1967,In_4244,In_2580);
nor U1968 (N_1968,In_1187,In_3768);
nor U1969 (N_1969,In_3598,In_1358);
nand U1970 (N_1970,In_600,In_1892);
nand U1971 (N_1971,In_222,In_4248);
and U1972 (N_1972,In_2035,In_2785);
or U1973 (N_1973,In_4359,In_4910);
nand U1974 (N_1974,In_1723,In_4095);
or U1975 (N_1975,In_4726,In_4607);
or U1976 (N_1976,In_2458,In_1099);
nor U1977 (N_1977,In_4422,In_845);
and U1978 (N_1978,In_1504,In_3716);
xor U1979 (N_1979,In_2304,In_4951);
xor U1980 (N_1980,In_611,In_2826);
and U1981 (N_1981,In_996,In_2255);
nor U1982 (N_1982,In_3352,In_1576);
nand U1983 (N_1983,In_686,In_1926);
and U1984 (N_1984,In_1324,In_2037);
xnor U1985 (N_1985,In_2615,In_4984);
and U1986 (N_1986,In_2900,In_1046);
and U1987 (N_1987,In_406,In_4747);
xor U1988 (N_1988,In_2129,In_1896);
xor U1989 (N_1989,In_622,In_1638);
xnor U1990 (N_1990,In_4478,In_1431);
and U1991 (N_1991,In_3840,In_3312);
or U1992 (N_1992,In_1024,In_3855);
or U1993 (N_1993,In_179,In_989);
nand U1994 (N_1994,In_3028,In_96);
xnor U1995 (N_1995,In_2385,In_4234);
nor U1996 (N_1996,In_4676,In_1013);
or U1997 (N_1997,In_4778,In_4457);
and U1998 (N_1998,In_4361,In_1689);
xnor U1999 (N_1999,In_1913,In_1973);
xnor U2000 (N_2000,In_4513,In_387);
or U2001 (N_2001,In_2461,In_800);
and U2002 (N_2002,In_1400,In_4390);
and U2003 (N_2003,In_2553,In_2703);
nor U2004 (N_2004,In_1459,In_616);
xor U2005 (N_2005,In_3592,In_3956);
or U2006 (N_2006,In_1436,In_2748);
nor U2007 (N_2007,In_2768,In_3476);
nand U2008 (N_2008,In_505,In_2599);
and U2009 (N_2009,In_3828,In_4705);
nand U2010 (N_2010,In_2004,In_719);
nand U2011 (N_2011,In_1143,In_3099);
nor U2012 (N_2012,In_1517,In_394);
nor U2013 (N_2013,In_4213,In_564);
nor U2014 (N_2014,In_3923,In_3980);
nand U2015 (N_2015,In_3128,In_3541);
xor U2016 (N_2016,In_4641,In_3761);
and U2017 (N_2017,In_937,In_3449);
or U2018 (N_2018,In_2360,In_2578);
xnor U2019 (N_2019,In_2380,In_3992);
xor U2020 (N_2020,In_1771,In_3317);
or U2021 (N_2021,In_676,In_2564);
xnor U2022 (N_2022,In_3822,In_4351);
or U2023 (N_2023,In_32,In_4715);
or U2024 (N_2024,In_4753,In_2470);
nor U2025 (N_2025,In_1300,In_3794);
nand U2026 (N_2026,In_4428,In_3730);
nor U2027 (N_2027,In_3829,In_3371);
or U2028 (N_2028,In_426,In_4367);
nor U2029 (N_2029,In_4346,In_3963);
xor U2030 (N_2030,In_3514,In_2056);
nor U2031 (N_2031,In_1102,In_2595);
nand U2032 (N_2032,In_2149,In_3630);
xor U2033 (N_2033,In_63,In_357);
or U2034 (N_2034,In_2696,In_1383);
and U2035 (N_2035,In_1860,In_1725);
nand U2036 (N_2036,In_2106,In_4855);
nand U2037 (N_2037,In_4632,In_2960);
and U2038 (N_2038,In_4161,In_385);
nor U2039 (N_2039,In_4682,In_1320);
and U2040 (N_2040,In_3053,In_3196);
nand U2041 (N_2041,In_2363,In_520);
nor U2042 (N_2042,In_2758,In_651);
or U2043 (N_2043,In_2878,In_47);
and U2044 (N_2044,In_3077,In_4794);
and U2045 (N_2045,In_3308,In_3832);
xor U2046 (N_2046,In_3544,In_1362);
or U2047 (N_2047,In_4599,In_4589);
nor U2048 (N_2048,In_920,In_1581);
nand U2049 (N_2049,In_2828,In_1560);
nor U2050 (N_2050,In_4942,In_1442);
nand U2051 (N_2051,In_4935,In_4160);
nor U2052 (N_2052,In_3684,In_3357);
and U2053 (N_2053,In_336,In_3368);
nand U2054 (N_2054,In_1891,In_3172);
or U2055 (N_2055,In_3399,In_350);
nand U2056 (N_2056,In_3661,In_3489);
nand U2057 (N_2057,In_752,In_2266);
nor U2058 (N_2058,In_1074,In_2484);
and U2059 (N_2059,In_3755,In_479);
nor U2060 (N_2060,In_2291,In_1097);
or U2061 (N_2061,In_836,In_4238);
nand U2062 (N_2062,In_2532,In_2528);
nor U2063 (N_2063,In_2569,In_4973);
xnor U2064 (N_2064,In_3634,In_1530);
nand U2065 (N_2065,In_776,In_1799);
xnor U2066 (N_2066,In_3260,In_3892);
and U2067 (N_2067,In_4214,In_2206);
or U2068 (N_2068,In_1373,In_1318);
or U2069 (N_2069,In_2727,In_4946);
or U2070 (N_2070,In_3933,In_182);
or U2071 (N_2071,In_2675,In_196);
and U2072 (N_2072,In_1494,In_1034);
nand U2073 (N_2073,In_1181,In_4835);
nand U2074 (N_2074,In_962,In_3210);
nor U2075 (N_2075,In_948,In_2440);
nand U2076 (N_2076,In_458,In_2690);
nand U2077 (N_2077,In_1205,In_527);
and U2078 (N_2078,In_3538,In_2981);
and U2079 (N_2079,In_430,In_2143);
nand U2080 (N_2080,In_4553,In_4056);
nor U2081 (N_2081,In_2126,In_1753);
xnor U2082 (N_2082,In_3883,In_3872);
and U2083 (N_2083,In_4051,In_1238);
nand U2084 (N_2084,In_3753,In_1806);
nor U2085 (N_2085,In_713,In_2431);
nor U2086 (N_2086,In_4624,In_4209);
and U2087 (N_2087,In_604,In_791);
nand U2088 (N_2088,In_4614,In_3173);
or U2089 (N_2089,In_2884,In_856);
nor U2090 (N_2090,In_4049,In_2145);
nand U2091 (N_2091,In_4048,In_4651);
and U2092 (N_2092,In_4583,In_1513);
nor U2093 (N_2093,In_227,In_4523);
nand U2094 (N_2094,In_1746,In_1980);
nor U2095 (N_2095,In_4497,In_1598);
and U2096 (N_2096,In_3871,In_309);
nand U2097 (N_2097,In_1064,In_4090);
nor U2098 (N_2098,In_950,In_2661);
xor U2099 (N_2099,In_3035,In_4504);
xor U2100 (N_2100,In_885,In_1760);
nor U2101 (N_2101,In_2051,In_3504);
nand U2102 (N_2102,In_239,In_2688);
nand U2103 (N_2103,In_413,In_1785);
nand U2104 (N_2104,In_3047,In_1683);
xnor U2105 (N_2105,In_2550,In_4787);
nand U2106 (N_2106,In_3937,In_4619);
nand U2107 (N_2107,In_2144,In_3695);
and U2108 (N_2108,In_2923,In_4633);
nor U2109 (N_2109,In_2273,In_4002);
or U2110 (N_2110,In_3345,In_3948);
and U2111 (N_2111,In_3932,In_4765);
nor U2112 (N_2112,In_3133,In_2517);
nand U2113 (N_2113,In_216,In_2210);
and U2114 (N_2114,In_973,In_2847);
xnor U2115 (N_2115,In_377,In_1664);
xnor U2116 (N_2116,In_2474,In_1885);
or U2117 (N_2117,In_2152,In_314);
nand U2118 (N_2118,In_4131,In_4414);
or U2119 (N_2119,In_3282,In_4666);
or U2120 (N_2120,In_692,In_4153);
or U2121 (N_2121,In_4981,In_3284);
xnor U2122 (N_2122,In_2561,In_2207);
xor U2123 (N_2123,In_2191,In_2087);
and U2124 (N_2124,In_4180,In_3503);
nand U2125 (N_2125,In_104,In_4577);
nand U2126 (N_2126,In_3164,In_4024);
nor U2127 (N_2127,In_1591,In_864);
xor U2128 (N_2128,In_4551,In_1972);
nor U2129 (N_2129,In_1405,In_2897);
nand U2130 (N_2130,In_4706,In_4972);
xnor U2131 (N_2131,In_689,In_3852);
xnor U2132 (N_2132,In_4040,In_420);
and U2133 (N_2133,In_963,In_3934);
nor U2134 (N_2134,In_3900,In_3336);
nor U2135 (N_2135,In_2802,In_2303);
nor U2136 (N_2136,In_3781,In_4891);
xor U2137 (N_2137,In_3869,In_1301);
and U2138 (N_2138,In_4404,In_4023);
or U2139 (N_2139,In_793,In_3985);
or U2140 (N_2140,In_242,In_2793);
nand U2141 (N_2141,In_234,In_900);
nor U2142 (N_2142,In_893,In_126);
nand U2143 (N_2143,In_911,In_4068);
xor U2144 (N_2144,In_2156,In_1765);
nor U2145 (N_2145,In_4185,In_3792);
nand U2146 (N_2146,In_2820,In_1763);
nand U2147 (N_2147,In_862,In_4389);
or U2148 (N_2148,In_3511,In_726);
nand U2149 (N_2149,In_3013,In_4486);
or U2150 (N_2150,In_4930,In_4799);
and U2151 (N_2151,In_3033,In_28);
xnor U2152 (N_2152,In_852,In_2695);
nor U2153 (N_2153,In_1976,In_2374);
nand U2154 (N_2154,In_509,In_4383);
nor U2155 (N_2155,In_1754,In_4375);
xnor U2156 (N_2156,In_2586,In_2407);
and U2157 (N_2157,In_4041,In_1470);
and U2158 (N_2158,In_1283,In_253);
and U2159 (N_2159,In_872,In_589);
nor U2160 (N_2160,In_1983,In_1389);
nor U2161 (N_2161,In_1732,In_2289);
nand U2162 (N_2162,In_4466,In_2177);
nor U2163 (N_2163,In_4477,In_2125);
nor U2164 (N_2164,In_3929,In_2375);
and U2165 (N_2165,In_3991,In_4451);
and U2166 (N_2166,In_2990,In_981);
and U2167 (N_2167,In_2302,In_2634);
or U2168 (N_2168,In_2598,In_1452);
and U2169 (N_2169,In_240,In_1333);
and U2170 (N_2170,In_602,In_1052);
and U2171 (N_2171,In_631,In_1047);
or U2172 (N_2172,In_2328,In_3823);
or U2173 (N_2173,In_3383,In_4241);
nand U2174 (N_2174,In_1705,In_2530);
or U2175 (N_2175,In_3103,In_193);
nand U2176 (N_2176,In_3643,In_1538);
xor U2177 (N_2177,In_2889,In_3294);
and U2178 (N_2178,In_4397,In_738);
or U2179 (N_2179,In_3236,In_4558);
and U2180 (N_2180,In_392,In_816);
nor U2181 (N_2181,In_906,In_951);
or U2182 (N_2182,In_4173,In_329);
or U2183 (N_2183,In_1484,In_3139);
xnor U2184 (N_2184,In_3031,In_1662);
nor U2185 (N_2185,In_71,In_636);
nor U2186 (N_2186,In_1458,In_680);
nor U2187 (N_2187,In_4133,In_4844);
or U2188 (N_2188,In_3108,In_4235);
nor U2189 (N_2189,In_3576,In_1173);
xnor U2190 (N_2190,In_4127,In_163);
nand U2191 (N_2191,In_2336,In_4192);
or U2192 (N_2192,In_1709,In_3957);
or U2193 (N_2193,In_1975,In_2761);
or U2194 (N_2194,In_2415,In_2076);
or U2195 (N_2195,In_2392,In_4934);
and U2196 (N_2196,In_2315,In_2849);
and U2197 (N_2197,In_93,In_4340);
nand U2198 (N_2198,In_3979,In_4860);
or U2199 (N_2199,In_876,In_4455);
nor U2200 (N_2200,In_313,In_2728);
or U2201 (N_2201,In_4548,In_2002);
xnor U2202 (N_2202,In_4091,In_2804);
xnor U2203 (N_2203,In_2866,In_4304);
and U2204 (N_2204,In_2387,In_750);
nand U2205 (N_2205,In_1630,In_2101);
and U2206 (N_2206,In_4343,In_557);
and U2207 (N_2207,In_3354,In_565);
nor U2208 (N_2208,In_3186,In_3650);
nand U2209 (N_2209,In_4373,In_901);
xor U2210 (N_2210,In_3265,In_3973);
nor U2211 (N_2211,In_3145,In_1988);
xnor U2212 (N_2212,In_828,In_2568);
xor U2213 (N_2213,In_2652,In_500);
nor U2214 (N_2214,In_2898,In_2072);
nor U2215 (N_2215,In_4680,In_38);
nor U2216 (N_2216,In_1990,In_4029);
and U2217 (N_2217,In_36,In_124);
xnor U2218 (N_2218,In_1481,In_2957);
xor U2219 (N_2219,In_2883,In_3709);
and U2220 (N_2220,In_4810,In_3355);
and U2221 (N_2221,In_2895,In_2358);
or U2222 (N_2222,In_65,In_2513);
and U2223 (N_2223,In_1096,In_1471);
and U2224 (N_2224,In_701,In_545);
nand U2225 (N_2225,In_1745,In_1040);
nor U2226 (N_2226,In_2249,In_3698);
and U2227 (N_2227,In_4571,In_287);
nor U2228 (N_2228,In_1866,In_3400);
and U2229 (N_2229,In_4654,In_4468);
xor U2230 (N_2230,In_873,In_1211);
nand U2231 (N_2231,In_300,In_4741);
xnor U2232 (N_2232,In_4895,In_581);
and U2233 (N_2233,In_4299,In_270);
nor U2234 (N_2234,In_4948,In_1418);
or U2235 (N_2235,In_4768,In_1888);
nand U2236 (N_2236,In_2683,In_4963);
or U2237 (N_2237,In_1311,In_730);
nor U2238 (N_2238,In_4298,In_3766);
and U2239 (N_2239,In_4148,In_3168);
xor U2240 (N_2240,In_2671,In_4249);
xnor U2241 (N_2241,In_916,In_2212);
and U2242 (N_2242,In_731,In_2404);
or U2243 (N_2243,In_1643,In_4116);
or U2244 (N_2244,In_1858,In_2723);
nand U2245 (N_2245,In_3039,In_1774);
or U2246 (N_2246,In_248,In_3142);
nand U2247 (N_2247,In_3137,In_683);
or U2248 (N_2248,In_3811,In_880);
xnor U2249 (N_2249,In_654,In_4851);
and U2250 (N_2250,In_481,In_4146);
nand U2251 (N_2251,In_1094,In_4853);
or U2252 (N_2252,In_2022,In_4227);
nand U2253 (N_2253,In_2341,In_4330);
and U2254 (N_2254,In_1714,In_903);
and U2255 (N_2255,In_3719,In_3438);
nand U2256 (N_2256,In_2195,In_1909);
xnor U2257 (N_2257,In_1306,In_858);
xor U2258 (N_2258,In_3831,In_1525);
and U2259 (N_2259,In_560,In_158);
xor U2260 (N_2260,In_2572,In_236);
nor U2261 (N_2261,In_4271,In_4281);
nand U2262 (N_2262,In_1811,In_2818);
xnor U2263 (N_2263,In_3206,In_2936);
xor U2264 (N_2264,In_2709,In_1616);
or U2265 (N_2265,In_2211,In_2257);
and U2266 (N_2266,In_4790,In_1213);
xnor U2267 (N_2267,In_1733,In_1526);
nand U2268 (N_2268,In_2426,In_441);
or U2269 (N_2269,In_1008,In_3830);
and U2270 (N_2270,In_4795,In_4670);
or U2271 (N_2271,In_4313,In_1595);
nor U2272 (N_2272,In_1170,In_4411);
or U2273 (N_2273,In_2269,In_2702);
nor U2274 (N_2274,In_4546,In_1347);
xnor U2275 (N_2275,In_3697,In_4989);
or U2276 (N_2276,In_1413,In_1816);
xor U2277 (N_2277,In_4117,In_3212);
nand U2278 (N_2278,In_3310,In_2441);
or U2279 (N_2279,In_1344,In_141);
xnor U2280 (N_2280,In_4841,In_2217);
and U2281 (N_2281,In_1905,In_4076);
or U2282 (N_2282,In_1221,In_2213);
or U2283 (N_2283,In_1328,In_4815);
nand U2284 (N_2284,In_1708,In_1682);
nor U2285 (N_2285,In_304,In_3244);
xnor U2286 (N_2286,In_737,In_4547);
xnor U2287 (N_2287,In_2203,In_2057);
xor U2288 (N_2288,In_1836,In_1878);
nor U2289 (N_2289,In_1031,In_2332);
nand U2290 (N_2290,In_1030,In_1675);
nor U2291 (N_2291,In_1026,In_576);
and U2292 (N_2292,In_2806,In_4273);
xnor U2293 (N_2293,In_1144,In_621);
nor U2294 (N_2294,In_3334,In_4827);
nor U2295 (N_2295,In_218,In_1737);
nor U2296 (N_2296,In_99,In_1460);
nand U2297 (N_2297,In_157,In_2216);
and U2298 (N_2298,In_2787,In_2366);
and U2299 (N_2299,In_922,In_127);
and U2300 (N_2300,In_2433,In_3018);
xor U2301 (N_2301,In_3672,In_4112);
nand U2302 (N_2302,In_2361,In_373);
or U2303 (N_2303,In_421,In_1473);
xor U2304 (N_2304,In_3170,In_2699);
nand U2305 (N_2305,In_691,In_2120);
and U2306 (N_2306,In_2457,In_605);
and U2307 (N_2307,In_3414,In_1569);
xor U2308 (N_2308,In_4155,In_2860);
nor U2309 (N_2309,In_4459,In_945);
nand U2310 (N_2310,In_4796,In_4442);
or U2311 (N_2311,In_3527,In_3095);
nor U2312 (N_2312,In_4216,In_4267);
xnor U2313 (N_2313,In_1599,In_835);
nand U2314 (N_2314,In_1665,In_1027);
or U2315 (N_2315,In_2772,In_4378);
and U2316 (N_2316,In_3380,In_2503);
nor U2317 (N_2317,In_4845,In_1958);
nor U2318 (N_2318,In_881,In_4377);
nor U2319 (N_2319,In_1655,In_2290);
nand U2320 (N_2320,In_2463,In_3834);
nor U2321 (N_2321,In_4658,In_2713);
xnor U2322 (N_2322,In_4324,In_1294);
or U2323 (N_2323,In_4974,In_4013);
or U2324 (N_2324,In_2721,In_4265);
and U2325 (N_2325,In_1700,In_967);
nand U2326 (N_2326,In_2928,In_3862);
nor U2327 (N_2327,In_2205,In_464);
nand U2328 (N_2328,In_1384,In_2644);
and U2329 (N_2329,In_3656,In_2299);
and U2330 (N_2330,In_1057,In_276);
nand U2331 (N_2331,In_3409,In_473);
xor U2332 (N_2332,In_2823,In_1142);
and U2333 (N_2333,In_453,In_102);
xnor U2334 (N_2334,In_3734,In_3190);
or U2335 (N_2335,In_2999,In_237);
xor U2336 (N_2336,In_1028,In_2416);
nand U2337 (N_2337,In_3169,In_2333);
nand U2338 (N_2338,In_2127,In_2966);
xor U2339 (N_2339,In_4643,In_3262);
nand U2340 (N_2340,In_2479,In_3833);
nor U2341 (N_2341,In_2274,In_2655);
xnor U2342 (N_2342,In_1502,In_1549);
nor U2343 (N_2343,In_3637,In_4320);
and U2344 (N_2344,In_4055,In_3534);
or U2345 (N_2345,In_3688,In_2367);
or U2346 (N_2346,In_4134,In_3365);
xor U2347 (N_2347,In_2829,In_4779);
nand U2348 (N_2348,In_2346,In_3089);
nor U2349 (N_2349,In_4824,In_4950);
or U2350 (N_2350,In_3498,In_853);
xnor U2351 (N_2351,In_2601,In_1434);
or U2352 (N_2352,In_4771,In_3421);
and U2353 (N_2353,In_114,In_1084);
and U2354 (N_2354,In_3640,In_2168);
nor U2355 (N_2355,In_1340,In_3471);
nor U2356 (N_2356,In_3741,In_3981);
nor U2357 (N_2357,In_3714,In_1272);
nor U2358 (N_2358,In_3483,In_398);
nor U2359 (N_2359,In_485,In_3865);
nor U2360 (N_2360,In_2925,In_459);
or U2361 (N_2361,In_2719,In_1508);
nor U2362 (N_2362,In_4953,In_4022);
xnor U2363 (N_2363,In_3926,In_1768);
nor U2364 (N_2364,In_783,In_3027);
nand U2365 (N_2365,In_1839,In_3331);
and U2366 (N_2366,In_1091,In_2682);
or U2367 (N_2367,In_3584,In_561);
xor U2368 (N_2368,In_1716,In_70);
xor U2369 (N_2369,In_2585,In_1626);
and U2370 (N_2370,In_302,In_1577);
nor U2371 (N_2371,In_1940,In_2483);
nand U2372 (N_2372,In_1232,In_2422);
or U2373 (N_2373,In_4081,In_3277);
nor U2374 (N_2374,In_4842,In_3589);
or U2375 (N_2375,In_2075,In_1252);
xnor U2376 (N_2376,In_2372,In_753);
or U2377 (N_2377,In_2132,In_1817);
xor U2378 (N_2378,In_43,In_436);
or U2379 (N_2379,In_477,In_3712);
and U2380 (N_2380,In_2626,In_2711);
nand U2381 (N_2381,In_4830,In_371);
or U2382 (N_2382,In_29,In_1103);
nor U2383 (N_2383,In_3611,In_3020);
nand U2384 (N_2384,In_4649,In_3193);
and U2385 (N_2385,In_1246,In_4522);
and U2386 (N_2386,In_2009,In_3733);
nor U2387 (N_2387,In_1587,In_2622);
and U2388 (N_2388,In_521,In_1331);
nor U2389 (N_2389,In_1862,In_652);
and U2390 (N_2390,In_3323,In_4515);
and U2391 (N_2391,In_2681,In_337);
xor U2392 (N_2392,In_3839,In_4332);
xor U2393 (N_2393,In_275,In_251);
nor U2394 (N_2394,In_741,In_733);
and U2395 (N_2395,In_3982,In_4398);
and U2396 (N_2396,In_3055,In_4982);
or U2397 (N_2397,In_620,In_4163);
xnor U2398 (N_2398,In_1125,In_184);
nor U2399 (N_2399,In_997,In_2080);
or U2400 (N_2400,In_2612,In_1353);
xnor U2401 (N_2401,In_4737,In_1447);
nand U2402 (N_2402,In_2103,In_847);
nor U2403 (N_2403,In_4620,In_1542);
nand U2404 (N_2404,In_280,In_493);
nand U2405 (N_2405,In_1042,In_3092);
xor U2406 (N_2406,In_3585,In_2325);
or U2407 (N_2407,In_1348,In_2398);
and U2408 (N_2408,In_4416,In_3030);
nor U2409 (N_2409,In_1987,In_846);
nand U2410 (N_2410,In_3332,In_483);
xor U2411 (N_2411,In_2911,In_3521);
nor U2412 (N_2412,In_4263,In_439);
nor U2413 (N_2413,In_3618,In_4151);
and U2414 (N_2414,In_4900,In_1867);
and U2415 (N_2415,In_4178,In_4099);
nand U2416 (N_2416,In_4020,In_2886);
and U2417 (N_2417,In_1864,In_593);
nor U2418 (N_2418,In_2038,In_2162);
xnor U2419 (N_2419,In_983,In_640);
nand U2420 (N_2420,In_4593,In_4286);
or U2421 (N_2421,In_3888,In_1755);
xor U2422 (N_2422,In_1793,In_3920);
nand U2423 (N_2423,In_4280,In_2927);
xor U2424 (N_2424,In_1902,In_4997);
and U2425 (N_2425,In_2141,In_1327);
nand U2426 (N_2426,In_195,In_1118);
nand U2427 (N_2427,In_2329,In_629);
nand U2428 (N_2428,In_2992,In_2485);
xor U2429 (N_2429,In_395,In_4732);
xor U2430 (N_2430,In_1115,In_1376);
or U2431 (N_2431,In_4848,In_4315);
nor U2432 (N_2432,In_2600,In_4424);
or U2433 (N_2433,In_199,In_1869);
nor U2434 (N_2434,In_699,In_2940);
and U2435 (N_2435,In_4865,In_501);
and U2436 (N_2436,In_2331,In_3639);
xnor U2437 (N_2437,In_2097,In_4107);
nor U2438 (N_2438,In_642,In_190);
xnor U2439 (N_2439,In_2323,In_1369);
and U2440 (N_2440,In_4580,In_1639);
xor U2441 (N_2441,In_2078,In_1775);
and U2442 (N_2442,In_4071,In_3677);
and U2443 (N_2443,In_4683,In_3216);
and U2444 (N_2444,In_2267,In_2052);
or U2445 (N_2445,In_3411,In_3052);
xnor U2446 (N_2446,In_79,In_1446);
nor U2447 (N_2447,In_2146,In_1692);
or U2448 (N_2448,In_2338,In_1322);
xor U2449 (N_2449,In_4840,In_3271);
xnor U2450 (N_2450,In_3346,In_837);
and U2451 (N_2451,In_2949,In_3071);
nor U2452 (N_2452,In_1739,In_1964);
or U2453 (N_2453,In_180,In_4667);
nand U2454 (N_2454,In_2045,In_499);
and U2455 (N_2455,In_1676,In_7);
xor U2456 (N_2456,In_869,In_289);
nand U2457 (N_2457,In_804,In_4839);
and U2458 (N_2458,In_354,In_3789);
nor U2459 (N_2459,In_671,In_4408);
xnor U2460 (N_2460,In_323,In_1948);
or U2461 (N_2461,In_55,In_1571);
and U2462 (N_2462,In_2623,In_4418);
or U2463 (N_2463,In_1268,In_2262);
and U2464 (N_2464,In_4080,In_1342);
nor U2465 (N_2465,In_2941,In_2330);
xor U2466 (N_2466,In_4122,In_2916);
nand U2467 (N_2467,In_646,In_1557);
xnor U2468 (N_2468,In_3093,In_1536);
nor U2469 (N_2469,In_4120,In_580);
nand U2470 (N_2470,In_5,In_4303);
nand U2471 (N_2471,In_89,In_3928);
nand U2472 (N_2472,In_1510,In_2587);
and U2473 (N_2473,In_4897,In_3539);
xor U2474 (N_2474,In_4719,In_4450);
nand U2475 (N_2475,In_4581,In_2839);
nand U2476 (N_2476,In_2512,In_2837);
nand U2477 (N_2477,In_3167,In_785);
or U2478 (N_2478,In_2789,In_3465);
xor U2479 (N_2479,In_4598,In_3044);
nand U2480 (N_2480,In_3687,In_2357);
nand U2481 (N_2481,In_1666,In_2673);
and U2482 (N_2482,In_3550,In_3401);
or U2483 (N_2483,In_656,In_2668);
nor U2484 (N_2484,In_1994,In_4640);
nand U2485 (N_2485,In_2736,In_61);
nand U2486 (N_2486,In_637,In_1109);
xor U2487 (N_2487,In_548,In_2014);
and U2488 (N_2488,In_4836,In_736);
nor U2489 (N_2489,In_3660,In_1721);
and U2490 (N_2490,In_591,In_2821);
nand U2491 (N_2491,In_3300,In_1293);
or U2492 (N_2492,In_103,In_2714);
nor U2493 (N_2493,In_960,In_4443);
xnor U2494 (N_2494,In_3998,In_1539);
nand U2495 (N_2495,In_3289,In_2784);
nand U2496 (N_2496,In_4759,In_1421);
xnor U2497 (N_2497,In_553,In_2063);
or U2498 (N_2498,In_409,In_316);
nor U2499 (N_2499,In_220,In_1202);
or U2500 (N_2500,In_1983,In_4668);
xnor U2501 (N_2501,In_3775,In_2493);
or U2502 (N_2502,In_2527,In_3057);
nor U2503 (N_2503,In_4147,In_438);
or U2504 (N_2504,In_2047,In_2380);
and U2505 (N_2505,In_4850,In_2296);
nor U2506 (N_2506,In_3541,In_860);
nand U2507 (N_2507,In_976,In_1146);
or U2508 (N_2508,In_2163,In_2217);
or U2509 (N_2509,In_1053,In_359);
or U2510 (N_2510,In_1326,In_640);
xor U2511 (N_2511,In_323,In_1377);
nand U2512 (N_2512,In_2344,In_2449);
or U2513 (N_2513,In_1076,In_2151);
nand U2514 (N_2514,In_3003,In_2947);
or U2515 (N_2515,In_3157,In_3073);
nor U2516 (N_2516,In_1273,In_3580);
or U2517 (N_2517,In_3253,In_4084);
xor U2518 (N_2518,In_2057,In_1263);
nand U2519 (N_2519,In_496,In_2337);
or U2520 (N_2520,In_3840,In_82);
nand U2521 (N_2521,In_2315,In_2485);
or U2522 (N_2522,In_3911,In_61);
nand U2523 (N_2523,In_551,In_3307);
and U2524 (N_2524,In_4071,In_3507);
xor U2525 (N_2525,In_3296,In_2169);
and U2526 (N_2526,In_4283,In_3999);
and U2527 (N_2527,In_830,In_1822);
nor U2528 (N_2528,In_3303,In_2869);
nor U2529 (N_2529,In_2026,In_1342);
xor U2530 (N_2530,In_4810,In_2814);
or U2531 (N_2531,In_509,In_4373);
xor U2532 (N_2532,In_1354,In_4719);
and U2533 (N_2533,In_1045,In_949);
and U2534 (N_2534,In_4488,In_3265);
and U2535 (N_2535,In_2968,In_2352);
and U2536 (N_2536,In_4202,In_2062);
xor U2537 (N_2537,In_554,In_1470);
nand U2538 (N_2538,In_4075,In_3797);
nor U2539 (N_2539,In_4457,In_3908);
and U2540 (N_2540,In_932,In_2378);
nand U2541 (N_2541,In_2384,In_733);
xor U2542 (N_2542,In_2062,In_1169);
nor U2543 (N_2543,In_2362,In_3097);
nor U2544 (N_2544,In_4976,In_3746);
or U2545 (N_2545,In_487,In_3817);
xnor U2546 (N_2546,In_2724,In_1271);
or U2547 (N_2547,In_1465,In_2185);
nand U2548 (N_2548,In_2838,In_4052);
nor U2549 (N_2549,In_1273,In_4452);
nand U2550 (N_2550,In_3269,In_3230);
nand U2551 (N_2551,In_3252,In_1357);
nand U2552 (N_2552,In_3653,In_870);
or U2553 (N_2553,In_904,In_3166);
and U2554 (N_2554,In_3684,In_4707);
or U2555 (N_2555,In_3955,In_2188);
nor U2556 (N_2556,In_547,In_1436);
nand U2557 (N_2557,In_1057,In_1634);
xor U2558 (N_2558,In_3732,In_1657);
nor U2559 (N_2559,In_574,In_4997);
and U2560 (N_2560,In_2201,In_4676);
and U2561 (N_2561,In_1162,In_3597);
xor U2562 (N_2562,In_608,In_1016);
or U2563 (N_2563,In_1064,In_2370);
and U2564 (N_2564,In_4993,In_1800);
xor U2565 (N_2565,In_3552,In_437);
xnor U2566 (N_2566,In_419,In_3406);
nor U2567 (N_2567,In_3311,In_1148);
nand U2568 (N_2568,In_12,In_686);
or U2569 (N_2569,In_2569,In_4250);
nand U2570 (N_2570,In_1557,In_4714);
and U2571 (N_2571,In_1396,In_4618);
nor U2572 (N_2572,In_3050,In_4700);
or U2573 (N_2573,In_3242,In_3366);
nor U2574 (N_2574,In_2108,In_492);
and U2575 (N_2575,In_3339,In_1697);
nor U2576 (N_2576,In_381,In_3327);
or U2577 (N_2577,In_3173,In_2956);
xor U2578 (N_2578,In_223,In_4723);
nor U2579 (N_2579,In_1079,In_1513);
or U2580 (N_2580,In_4342,In_1716);
nor U2581 (N_2581,In_359,In_1112);
or U2582 (N_2582,In_2117,In_78);
and U2583 (N_2583,In_3452,In_3429);
and U2584 (N_2584,In_3317,In_1249);
nor U2585 (N_2585,In_698,In_3953);
xnor U2586 (N_2586,In_1435,In_4851);
nand U2587 (N_2587,In_1979,In_2935);
xor U2588 (N_2588,In_2162,In_1572);
nor U2589 (N_2589,In_1635,In_2347);
or U2590 (N_2590,In_1453,In_1443);
xnor U2591 (N_2591,In_3520,In_2626);
nor U2592 (N_2592,In_4652,In_772);
or U2593 (N_2593,In_281,In_2103);
nand U2594 (N_2594,In_2390,In_69);
xor U2595 (N_2595,In_271,In_3057);
and U2596 (N_2596,In_3549,In_2798);
nor U2597 (N_2597,In_358,In_3974);
or U2598 (N_2598,In_1279,In_229);
and U2599 (N_2599,In_1098,In_3850);
nor U2600 (N_2600,In_636,In_1945);
nand U2601 (N_2601,In_2927,In_2639);
or U2602 (N_2602,In_3455,In_1018);
and U2603 (N_2603,In_1038,In_3726);
nor U2604 (N_2604,In_3813,In_1842);
nand U2605 (N_2605,In_4928,In_4900);
and U2606 (N_2606,In_2709,In_2136);
and U2607 (N_2607,In_2354,In_1427);
nand U2608 (N_2608,In_3413,In_3246);
and U2609 (N_2609,In_4407,In_1174);
and U2610 (N_2610,In_324,In_1558);
and U2611 (N_2611,In_4421,In_2495);
xor U2612 (N_2612,In_2272,In_3075);
or U2613 (N_2613,In_4952,In_644);
or U2614 (N_2614,In_4782,In_2173);
nand U2615 (N_2615,In_1514,In_412);
nor U2616 (N_2616,In_308,In_3044);
nor U2617 (N_2617,In_4212,In_467);
nand U2618 (N_2618,In_3426,In_2293);
xor U2619 (N_2619,In_3972,In_4615);
xnor U2620 (N_2620,In_4344,In_1838);
and U2621 (N_2621,In_2346,In_1727);
nor U2622 (N_2622,In_1842,In_4780);
and U2623 (N_2623,In_4120,In_1517);
or U2624 (N_2624,In_3488,In_2393);
xor U2625 (N_2625,In_4735,In_4807);
or U2626 (N_2626,In_3977,In_1652);
or U2627 (N_2627,In_3545,In_1461);
or U2628 (N_2628,In_4296,In_4325);
and U2629 (N_2629,In_3621,In_13);
nor U2630 (N_2630,In_2027,In_3361);
xor U2631 (N_2631,In_3210,In_3769);
xor U2632 (N_2632,In_3795,In_2462);
or U2633 (N_2633,In_4732,In_1350);
nor U2634 (N_2634,In_2801,In_3978);
or U2635 (N_2635,In_3175,In_2813);
and U2636 (N_2636,In_4967,In_3657);
or U2637 (N_2637,In_3776,In_2277);
or U2638 (N_2638,In_4703,In_633);
nor U2639 (N_2639,In_3450,In_2261);
and U2640 (N_2640,In_1661,In_1556);
or U2641 (N_2641,In_156,In_606);
nor U2642 (N_2642,In_2319,In_3261);
or U2643 (N_2643,In_4216,In_2635);
nand U2644 (N_2644,In_1528,In_4705);
or U2645 (N_2645,In_3919,In_3252);
and U2646 (N_2646,In_1785,In_2515);
xor U2647 (N_2647,In_4804,In_4282);
and U2648 (N_2648,In_3186,In_4229);
xnor U2649 (N_2649,In_4808,In_2702);
nor U2650 (N_2650,In_2646,In_580);
xnor U2651 (N_2651,In_1094,In_3068);
xor U2652 (N_2652,In_4986,In_2904);
nor U2653 (N_2653,In_4195,In_1811);
or U2654 (N_2654,In_2737,In_2733);
and U2655 (N_2655,In_1240,In_3627);
nand U2656 (N_2656,In_1500,In_2713);
xor U2657 (N_2657,In_4468,In_1907);
and U2658 (N_2658,In_4911,In_753);
nand U2659 (N_2659,In_4909,In_456);
nand U2660 (N_2660,In_887,In_885);
nor U2661 (N_2661,In_4203,In_4065);
nand U2662 (N_2662,In_1588,In_674);
xor U2663 (N_2663,In_2741,In_3793);
xor U2664 (N_2664,In_2775,In_4578);
or U2665 (N_2665,In_1210,In_308);
and U2666 (N_2666,In_189,In_2876);
xnor U2667 (N_2667,In_3016,In_2562);
nand U2668 (N_2668,In_744,In_3399);
xor U2669 (N_2669,In_3930,In_1913);
and U2670 (N_2670,In_2382,In_705);
xor U2671 (N_2671,In_277,In_2617);
or U2672 (N_2672,In_175,In_3511);
xnor U2673 (N_2673,In_1612,In_2206);
nor U2674 (N_2674,In_51,In_1989);
xnor U2675 (N_2675,In_3141,In_543);
or U2676 (N_2676,In_4340,In_1565);
and U2677 (N_2677,In_503,In_1194);
xnor U2678 (N_2678,In_1711,In_3683);
and U2679 (N_2679,In_925,In_2028);
nor U2680 (N_2680,In_2826,In_3475);
or U2681 (N_2681,In_555,In_4097);
and U2682 (N_2682,In_3984,In_3877);
nand U2683 (N_2683,In_2560,In_1920);
nand U2684 (N_2684,In_784,In_711);
nor U2685 (N_2685,In_636,In_3225);
nand U2686 (N_2686,In_4366,In_3776);
or U2687 (N_2687,In_1137,In_4546);
nand U2688 (N_2688,In_2310,In_4263);
or U2689 (N_2689,In_4071,In_697);
xnor U2690 (N_2690,In_1049,In_4325);
nand U2691 (N_2691,In_4997,In_671);
nor U2692 (N_2692,In_3908,In_3576);
xnor U2693 (N_2693,In_3586,In_4955);
xor U2694 (N_2694,In_1592,In_4333);
nor U2695 (N_2695,In_973,In_1744);
nand U2696 (N_2696,In_3811,In_516);
nor U2697 (N_2697,In_2037,In_3078);
xnor U2698 (N_2698,In_329,In_1246);
nor U2699 (N_2699,In_4342,In_3071);
nor U2700 (N_2700,In_2179,In_2344);
xor U2701 (N_2701,In_907,In_1278);
xnor U2702 (N_2702,In_4245,In_2103);
nor U2703 (N_2703,In_3974,In_4096);
and U2704 (N_2704,In_4209,In_2657);
and U2705 (N_2705,In_1802,In_104);
xnor U2706 (N_2706,In_2875,In_2162);
or U2707 (N_2707,In_4824,In_1953);
and U2708 (N_2708,In_3087,In_2849);
and U2709 (N_2709,In_793,In_287);
nor U2710 (N_2710,In_3493,In_2885);
xnor U2711 (N_2711,In_4477,In_4887);
nand U2712 (N_2712,In_3714,In_1883);
xor U2713 (N_2713,In_3778,In_3730);
or U2714 (N_2714,In_1840,In_1639);
and U2715 (N_2715,In_472,In_1436);
nor U2716 (N_2716,In_4830,In_243);
and U2717 (N_2717,In_2340,In_2318);
nand U2718 (N_2718,In_840,In_1406);
or U2719 (N_2719,In_369,In_3593);
nand U2720 (N_2720,In_4125,In_1495);
and U2721 (N_2721,In_1954,In_2333);
nor U2722 (N_2722,In_2384,In_2173);
nand U2723 (N_2723,In_3602,In_1117);
nor U2724 (N_2724,In_1241,In_4568);
and U2725 (N_2725,In_1072,In_4383);
xnor U2726 (N_2726,In_3982,In_1222);
or U2727 (N_2727,In_3858,In_715);
and U2728 (N_2728,In_3665,In_4705);
nor U2729 (N_2729,In_4594,In_4744);
or U2730 (N_2730,In_2289,In_2236);
xor U2731 (N_2731,In_182,In_1173);
nor U2732 (N_2732,In_3477,In_3087);
nand U2733 (N_2733,In_2730,In_2341);
nor U2734 (N_2734,In_3011,In_1476);
or U2735 (N_2735,In_827,In_2113);
and U2736 (N_2736,In_2309,In_1875);
nand U2737 (N_2737,In_4437,In_2648);
nor U2738 (N_2738,In_3189,In_483);
xnor U2739 (N_2739,In_3861,In_4156);
nor U2740 (N_2740,In_2839,In_661);
and U2741 (N_2741,In_4640,In_981);
nand U2742 (N_2742,In_129,In_821);
or U2743 (N_2743,In_3928,In_3259);
nor U2744 (N_2744,In_4585,In_1162);
xor U2745 (N_2745,In_3052,In_3035);
and U2746 (N_2746,In_854,In_2072);
nor U2747 (N_2747,In_484,In_1621);
nor U2748 (N_2748,In_4461,In_3274);
nand U2749 (N_2749,In_368,In_3387);
nor U2750 (N_2750,In_3340,In_3472);
nand U2751 (N_2751,In_2562,In_3900);
nand U2752 (N_2752,In_3656,In_4592);
nor U2753 (N_2753,In_1721,In_509);
and U2754 (N_2754,In_2621,In_2462);
and U2755 (N_2755,In_1031,In_1151);
nand U2756 (N_2756,In_2936,In_841);
nand U2757 (N_2757,In_2958,In_4464);
or U2758 (N_2758,In_2734,In_2160);
xor U2759 (N_2759,In_4271,In_1054);
xor U2760 (N_2760,In_2775,In_3280);
nand U2761 (N_2761,In_1514,In_2353);
nand U2762 (N_2762,In_3717,In_773);
nand U2763 (N_2763,In_3712,In_1337);
nor U2764 (N_2764,In_877,In_568);
and U2765 (N_2765,In_2261,In_4987);
xnor U2766 (N_2766,In_1274,In_186);
xor U2767 (N_2767,In_4312,In_299);
or U2768 (N_2768,In_3386,In_2420);
nand U2769 (N_2769,In_4746,In_4846);
or U2770 (N_2770,In_1067,In_4408);
or U2771 (N_2771,In_2767,In_1894);
or U2772 (N_2772,In_4858,In_3642);
or U2773 (N_2773,In_4438,In_474);
or U2774 (N_2774,In_4588,In_1453);
nand U2775 (N_2775,In_2233,In_2922);
or U2776 (N_2776,In_3899,In_863);
or U2777 (N_2777,In_3973,In_111);
or U2778 (N_2778,In_4227,In_60);
xnor U2779 (N_2779,In_1053,In_4336);
or U2780 (N_2780,In_1260,In_1259);
nor U2781 (N_2781,In_1075,In_954);
nor U2782 (N_2782,In_357,In_92);
and U2783 (N_2783,In_285,In_2754);
or U2784 (N_2784,In_1752,In_1984);
nand U2785 (N_2785,In_4171,In_1953);
and U2786 (N_2786,In_1457,In_4623);
and U2787 (N_2787,In_1628,In_588);
nand U2788 (N_2788,In_4651,In_4867);
xnor U2789 (N_2789,In_3078,In_2571);
xnor U2790 (N_2790,In_3913,In_2226);
xnor U2791 (N_2791,In_2406,In_4714);
and U2792 (N_2792,In_4907,In_2363);
xor U2793 (N_2793,In_3770,In_720);
nand U2794 (N_2794,In_1003,In_4117);
nor U2795 (N_2795,In_111,In_2142);
or U2796 (N_2796,In_4923,In_2880);
or U2797 (N_2797,In_4869,In_2815);
and U2798 (N_2798,In_3634,In_4295);
or U2799 (N_2799,In_4001,In_4772);
nor U2800 (N_2800,In_3998,In_957);
nor U2801 (N_2801,In_1417,In_4034);
and U2802 (N_2802,In_1273,In_3487);
or U2803 (N_2803,In_35,In_2933);
nand U2804 (N_2804,In_1632,In_1727);
nor U2805 (N_2805,In_1425,In_300);
nand U2806 (N_2806,In_694,In_3041);
xor U2807 (N_2807,In_1686,In_1469);
nor U2808 (N_2808,In_864,In_4816);
or U2809 (N_2809,In_2759,In_2775);
xnor U2810 (N_2810,In_1320,In_2951);
nand U2811 (N_2811,In_561,In_4402);
nor U2812 (N_2812,In_2524,In_750);
and U2813 (N_2813,In_263,In_1709);
xor U2814 (N_2814,In_2757,In_1971);
nor U2815 (N_2815,In_4226,In_2875);
or U2816 (N_2816,In_1534,In_4776);
xnor U2817 (N_2817,In_144,In_3548);
or U2818 (N_2818,In_2936,In_2448);
and U2819 (N_2819,In_829,In_3830);
and U2820 (N_2820,In_3524,In_1109);
xor U2821 (N_2821,In_3557,In_852);
nor U2822 (N_2822,In_3008,In_1783);
and U2823 (N_2823,In_4005,In_857);
nand U2824 (N_2824,In_2197,In_1907);
and U2825 (N_2825,In_2172,In_796);
xor U2826 (N_2826,In_1637,In_509);
xor U2827 (N_2827,In_4136,In_2687);
or U2828 (N_2828,In_2665,In_2197);
and U2829 (N_2829,In_1393,In_1854);
or U2830 (N_2830,In_4845,In_3421);
nand U2831 (N_2831,In_2240,In_92);
xor U2832 (N_2832,In_2149,In_4190);
nor U2833 (N_2833,In_1529,In_4770);
nor U2834 (N_2834,In_2350,In_3501);
xor U2835 (N_2835,In_2377,In_3481);
or U2836 (N_2836,In_4366,In_1082);
or U2837 (N_2837,In_4282,In_3402);
nand U2838 (N_2838,In_2869,In_3397);
nand U2839 (N_2839,In_2674,In_655);
xnor U2840 (N_2840,In_1754,In_3136);
nand U2841 (N_2841,In_61,In_181);
nor U2842 (N_2842,In_151,In_1417);
nand U2843 (N_2843,In_4913,In_2636);
xor U2844 (N_2844,In_1128,In_2025);
nand U2845 (N_2845,In_4064,In_1486);
nand U2846 (N_2846,In_3207,In_3837);
and U2847 (N_2847,In_4826,In_1760);
or U2848 (N_2848,In_1649,In_219);
nor U2849 (N_2849,In_4775,In_760);
nor U2850 (N_2850,In_4962,In_2148);
nor U2851 (N_2851,In_821,In_654);
or U2852 (N_2852,In_3656,In_4645);
and U2853 (N_2853,In_1946,In_1637);
or U2854 (N_2854,In_2160,In_1868);
nand U2855 (N_2855,In_1956,In_2124);
xnor U2856 (N_2856,In_1505,In_2481);
and U2857 (N_2857,In_1139,In_4202);
or U2858 (N_2858,In_1895,In_1223);
xor U2859 (N_2859,In_1250,In_2418);
nand U2860 (N_2860,In_4,In_4148);
nor U2861 (N_2861,In_4030,In_3946);
xnor U2862 (N_2862,In_1772,In_377);
nor U2863 (N_2863,In_4663,In_420);
xnor U2864 (N_2864,In_3598,In_3679);
xnor U2865 (N_2865,In_4087,In_1281);
nand U2866 (N_2866,In_4719,In_1137);
and U2867 (N_2867,In_1490,In_3921);
xnor U2868 (N_2868,In_2554,In_991);
nor U2869 (N_2869,In_1253,In_1264);
and U2870 (N_2870,In_650,In_3643);
and U2871 (N_2871,In_1580,In_613);
nand U2872 (N_2872,In_3269,In_1030);
and U2873 (N_2873,In_3625,In_868);
nand U2874 (N_2874,In_3481,In_4684);
nand U2875 (N_2875,In_2386,In_1938);
or U2876 (N_2876,In_1281,In_4026);
nand U2877 (N_2877,In_1211,In_4914);
nand U2878 (N_2878,In_4585,In_3785);
nand U2879 (N_2879,In_238,In_4559);
and U2880 (N_2880,In_1381,In_4771);
and U2881 (N_2881,In_3085,In_1888);
nor U2882 (N_2882,In_4160,In_1227);
and U2883 (N_2883,In_3777,In_3005);
or U2884 (N_2884,In_4734,In_4948);
nand U2885 (N_2885,In_2331,In_4191);
nor U2886 (N_2886,In_124,In_4432);
and U2887 (N_2887,In_4117,In_1025);
xnor U2888 (N_2888,In_2719,In_4315);
nand U2889 (N_2889,In_1377,In_3338);
nand U2890 (N_2890,In_515,In_2054);
nand U2891 (N_2891,In_513,In_2406);
and U2892 (N_2892,In_700,In_831);
or U2893 (N_2893,In_4812,In_2324);
nor U2894 (N_2894,In_2702,In_1986);
nor U2895 (N_2895,In_3100,In_358);
nand U2896 (N_2896,In_2374,In_845);
nor U2897 (N_2897,In_3536,In_1895);
xnor U2898 (N_2898,In_4024,In_459);
nor U2899 (N_2899,In_1210,In_1532);
or U2900 (N_2900,In_3577,In_900);
xnor U2901 (N_2901,In_3445,In_1334);
nor U2902 (N_2902,In_3792,In_3101);
xor U2903 (N_2903,In_2864,In_277);
nand U2904 (N_2904,In_2921,In_144);
and U2905 (N_2905,In_2234,In_1999);
nand U2906 (N_2906,In_4700,In_2362);
and U2907 (N_2907,In_932,In_779);
nor U2908 (N_2908,In_4938,In_3721);
and U2909 (N_2909,In_2859,In_1559);
xnor U2910 (N_2910,In_4336,In_4965);
nand U2911 (N_2911,In_1229,In_3960);
and U2912 (N_2912,In_1651,In_313);
xnor U2913 (N_2913,In_4050,In_114);
nand U2914 (N_2914,In_4098,In_4910);
xnor U2915 (N_2915,In_1991,In_2308);
nor U2916 (N_2916,In_1540,In_3925);
nor U2917 (N_2917,In_4546,In_501);
or U2918 (N_2918,In_3604,In_882);
nand U2919 (N_2919,In_4813,In_3443);
or U2920 (N_2920,In_2624,In_4649);
nand U2921 (N_2921,In_4137,In_3665);
and U2922 (N_2922,In_644,In_1244);
nand U2923 (N_2923,In_4229,In_4710);
and U2924 (N_2924,In_1118,In_777);
or U2925 (N_2925,In_3028,In_1473);
xnor U2926 (N_2926,In_4198,In_992);
nand U2927 (N_2927,In_3869,In_3091);
nand U2928 (N_2928,In_762,In_4963);
nor U2929 (N_2929,In_1961,In_1842);
nand U2930 (N_2930,In_688,In_2006);
and U2931 (N_2931,In_1568,In_4135);
xnor U2932 (N_2932,In_2935,In_4583);
xnor U2933 (N_2933,In_4540,In_1154);
and U2934 (N_2934,In_4483,In_761);
or U2935 (N_2935,In_166,In_2907);
xor U2936 (N_2936,In_1251,In_2097);
or U2937 (N_2937,In_1236,In_3671);
nand U2938 (N_2938,In_2724,In_158);
nor U2939 (N_2939,In_1955,In_2821);
nor U2940 (N_2940,In_1582,In_363);
xor U2941 (N_2941,In_1754,In_756);
nor U2942 (N_2942,In_4072,In_2939);
and U2943 (N_2943,In_1306,In_1561);
nand U2944 (N_2944,In_4964,In_2910);
nor U2945 (N_2945,In_1814,In_1278);
xnor U2946 (N_2946,In_6,In_375);
or U2947 (N_2947,In_4620,In_2373);
nand U2948 (N_2948,In_4228,In_1050);
nand U2949 (N_2949,In_4900,In_141);
xnor U2950 (N_2950,In_629,In_2517);
or U2951 (N_2951,In_1359,In_1668);
xor U2952 (N_2952,In_4959,In_279);
xor U2953 (N_2953,In_517,In_4120);
or U2954 (N_2954,In_1474,In_4301);
xor U2955 (N_2955,In_2464,In_4131);
and U2956 (N_2956,In_4741,In_3774);
or U2957 (N_2957,In_3132,In_756);
nand U2958 (N_2958,In_3730,In_570);
or U2959 (N_2959,In_3104,In_1929);
or U2960 (N_2960,In_3950,In_571);
and U2961 (N_2961,In_278,In_1952);
and U2962 (N_2962,In_2984,In_2601);
or U2963 (N_2963,In_2211,In_3090);
nand U2964 (N_2964,In_1015,In_1822);
nand U2965 (N_2965,In_3428,In_4648);
or U2966 (N_2966,In_932,In_4772);
nand U2967 (N_2967,In_3484,In_200);
nor U2968 (N_2968,In_3905,In_1403);
and U2969 (N_2969,In_1936,In_3181);
and U2970 (N_2970,In_4783,In_1315);
xnor U2971 (N_2971,In_271,In_349);
or U2972 (N_2972,In_1343,In_3477);
nor U2973 (N_2973,In_2781,In_4375);
nor U2974 (N_2974,In_3258,In_4627);
or U2975 (N_2975,In_3642,In_3221);
xnor U2976 (N_2976,In_310,In_824);
and U2977 (N_2977,In_1055,In_542);
xnor U2978 (N_2978,In_2976,In_4618);
nand U2979 (N_2979,In_1753,In_4039);
xnor U2980 (N_2980,In_1208,In_3411);
or U2981 (N_2981,In_927,In_2008);
nand U2982 (N_2982,In_2336,In_4152);
or U2983 (N_2983,In_2663,In_2350);
or U2984 (N_2984,In_2186,In_1599);
nand U2985 (N_2985,In_3846,In_982);
nor U2986 (N_2986,In_1101,In_2971);
nand U2987 (N_2987,In_3397,In_1355);
nand U2988 (N_2988,In_299,In_4244);
or U2989 (N_2989,In_4334,In_1918);
or U2990 (N_2990,In_4620,In_1079);
nor U2991 (N_2991,In_943,In_4956);
nor U2992 (N_2992,In_182,In_2482);
and U2993 (N_2993,In_1856,In_4697);
xor U2994 (N_2994,In_4882,In_4121);
nor U2995 (N_2995,In_696,In_1863);
xor U2996 (N_2996,In_1526,In_772);
or U2997 (N_2997,In_2807,In_2716);
or U2998 (N_2998,In_551,In_3411);
or U2999 (N_2999,In_2939,In_2654);
and U3000 (N_3000,In_3656,In_3007);
xor U3001 (N_3001,In_3730,In_2579);
nor U3002 (N_3002,In_4347,In_1583);
nor U3003 (N_3003,In_1888,In_4588);
xor U3004 (N_3004,In_1855,In_1697);
nand U3005 (N_3005,In_3691,In_704);
or U3006 (N_3006,In_4111,In_2891);
nand U3007 (N_3007,In_1751,In_2454);
or U3008 (N_3008,In_2741,In_162);
and U3009 (N_3009,In_288,In_4814);
nor U3010 (N_3010,In_2205,In_1447);
xnor U3011 (N_3011,In_2686,In_2892);
xnor U3012 (N_3012,In_4976,In_1479);
and U3013 (N_3013,In_244,In_550);
nand U3014 (N_3014,In_2850,In_3814);
and U3015 (N_3015,In_3347,In_1264);
nand U3016 (N_3016,In_3406,In_4721);
nand U3017 (N_3017,In_1904,In_1884);
and U3018 (N_3018,In_2456,In_1048);
and U3019 (N_3019,In_1891,In_4783);
nor U3020 (N_3020,In_83,In_1539);
or U3021 (N_3021,In_595,In_1093);
xor U3022 (N_3022,In_3837,In_2808);
xor U3023 (N_3023,In_329,In_609);
xnor U3024 (N_3024,In_1304,In_1539);
and U3025 (N_3025,In_3314,In_3409);
xor U3026 (N_3026,In_836,In_1814);
nor U3027 (N_3027,In_1352,In_88);
nor U3028 (N_3028,In_3451,In_1107);
xor U3029 (N_3029,In_4396,In_2107);
and U3030 (N_3030,In_1091,In_1221);
xnor U3031 (N_3031,In_3414,In_1583);
nor U3032 (N_3032,In_3100,In_1991);
and U3033 (N_3033,In_3708,In_4212);
nor U3034 (N_3034,In_4039,In_960);
and U3035 (N_3035,In_2856,In_93);
nand U3036 (N_3036,In_114,In_3322);
xnor U3037 (N_3037,In_2024,In_4602);
nand U3038 (N_3038,In_4119,In_1354);
and U3039 (N_3039,In_4548,In_474);
or U3040 (N_3040,In_4005,In_4663);
or U3041 (N_3041,In_195,In_542);
or U3042 (N_3042,In_3489,In_207);
nand U3043 (N_3043,In_3704,In_1871);
or U3044 (N_3044,In_3181,In_960);
nor U3045 (N_3045,In_3678,In_2028);
or U3046 (N_3046,In_4709,In_60);
or U3047 (N_3047,In_3604,In_4774);
xnor U3048 (N_3048,In_3883,In_3770);
xor U3049 (N_3049,In_4533,In_2099);
xnor U3050 (N_3050,In_436,In_1325);
nand U3051 (N_3051,In_1451,In_2205);
nand U3052 (N_3052,In_3036,In_4660);
nand U3053 (N_3053,In_1495,In_1432);
or U3054 (N_3054,In_3879,In_2782);
xor U3055 (N_3055,In_4393,In_314);
or U3056 (N_3056,In_372,In_1291);
nand U3057 (N_3057,In_3176,In_4674);
nor U3058 (N_3058,In_1996,In_2173);
and U3059 (N_3059,In_852,In_1863);
or U3060 (N_3060,In_878,In_133);
xor U3061 (N_3061,In_1402,In_4853);
and U3062 (N_3062,In_2817,In_1455);
and U3063 (N_3063,In_4469,In_1545);
nand U3064 (N_3064,In_811,In_4287);
xnor U3065 (N_3065,In_3047,In_2995);
xnor U3066 (N_3066,In_3669,In_3030);
nand U3067 (N_3067,In_2350,In_3979);
or U3068 (N_3068,In_626,In_712);
and U3069 (N_3069,In_1652,In_2506);
and U3070 (N_3070,In_246,In_521);
nor U3071 (N_3071,In_3615,In_3393);
nor U3072 (N_3072,In_3672,In_1989);
nor U3073 (N_3073,In_1851,In_2162);
or U3074 (N_3074,In_3895,In_3475);
xnor U3075 (N_3075,In_3893,In_2509);
xnor U3076 (N_3076,In_3941,In_665);
nand U3077 (N_3077,In_2970,In_2291);
and U3078 (N_3078,In_2201,In_4961);
or U3079 (N_3079,In_2972,In_3193);
nand U3080 (N_3080,In_4195,In_963);
and U3081 (N_3081,In_4390,In_2888);
and U3082 (N_3082,In_934,In_865);
and U3083 (N_3083,In_4862,In_3900);
or U3084 (N_3084,In_2239,In_1207);
xnor U3085 (N_3085,In_2143,In_3663);
and U3086 (N_3086,In_371,In_1522);
nor U3087 (N_3087,In_1682,In_155);
nand U3088 (N_3088,In_4507,In_2949);
nor U3089 (N_3089,In_4300,In_820);
or U3090 (N_3090,In_2132,In_2766);
nor U3091 (N_3091,In_731,In_1130);
nor U3092 (N_3092,In_4128,In_3842);
xnor U3093 (N_3093,In_628,In_1508);
or U3094 (N_3094,In_4057,In_2820);
nand U3095 (N_3095,In_4719,In_3117);
nor U3096 (N_3096,In_2381,In_2991);
and U3097 (N_3097,In_8,In_4320);
nand U3098 (N_3098,In_1724,In_73);
or U3099 (N_3099,In_3327,In_1875);
nand U3100 (N_3100,In_3026,In_1095);
or U3101 (N_3101,In_3520,In_1311);
nand U3102 (N_3102,In_1212,In_240);
nor U3103 (N_3103,In_2406,In_230);
nand U3104 (N_3104,In_1462,In_1562);
and U3105 (N_3105,In_1595,In_3989);
and U3106 (N_3106,In_2154,In_2350);
and U3107 (N_3107,In_385,In_2175);
or U3108 (N_3108,In_2448,In_3905);
nand U3109 (N_3109,In_591,In_2745);
nor U3110 (N_3110,In_2703,In_283);
xnor U3111 (N_3111,In_4267,In_3417);
nor U3112 (N_3112,In_4178,In_4431);
or U3113 (N_3113,In_1985,In_4899);
or U3114 (N_3114,In_2722,In_753);
and U3115 (N_3115,In_2272,In_4269);
xor U3116 (N_3116,In_3146,In_3849);
nor U3117 (N_3117,In_2228,In_1889);
and U3118 (N_3118,In_2330,In_4316);
nor U3119 (N_3119,In_1201,In_2252);
and U3120 (N_3120,In_3730,In_2776);
xor U3121 (N_3121,In_4210,In_898);
nor U3122 (N_3122,In_947,In_4757);
xor U3123 (N_3123,In_787,In_1734);
or U3124 (N_3124,In_127,In_4244);
nand U3125 (N_3125,In_2889,In_469);
xnor U3126 (N_3126,In_3620,In_4681);
nand U3127 (N_3127,In_3505,In_3061);
xnor U3128 (N_3128,In_1848,In_3756);
nand U3129 (N_3129,In_3835,In_1802);
or U3130 (N_3130,In_835,In_2245);
nor U3131 (N_3131,In_3559,In_873);
nand U3132 (N_3132,In_1098,In_3360);
nor U3133 (N_3133,In_2563,In_2394);
nand U3134 (N_3134,In_3771,In_3453);
or U3135 (N_3135,In_4173,In_2077);
xnor U3136 (N_3136,In_2767,In_1697);
and U3137 (N_3137,In_2479,In_3653);
xor U3138 (N_3138,In_4687,In_3137);
or U3139 (N_3139,In_2811,In_3731);
or U3140 (N_3140,In_3087,In_2400);
nor U3141 (N_3141,In_2384,In_2896);
xor U3142 (N_3142,In_4609,In_1428);
and U3143 (N_3143,In_478,In_2799);
or U3144 (N_3144,In_1561,In_1689);
nand U3145 (N_3145,In_4669,In_1470);
nor U3146 (N_3146,In_2172,In_4172);
nand U3147 (N_3147,In_1192,In_3048);
or U3148 (N_3148,In_4688,In_4054);
nand U3149 (N_3149,In_2272,In_4616);
and U3150 (N_3150,In_4983,In_900);
or U3151 (N_3151,In_3565,In_10);
or U3152 (N_3152,In_814,In_1798);
xor U3153 (N_3153,In_4362,In_4814);
xor U3154 (N_3154,In_1615,In_1894);
nor U3155 (N_3155,In_4959,In_1877);
xnor U3156 (N_3156,In_3092,In_4716);
and U3157 (N_3157,In_61,In_1964);
nor U3158 (N_3158,In_3909,In_3079);
and U3159 (N_3159,In_1357,In_921);
and U3160 (N_3160,In_1436,In_985);
xnor U3161 (N_3161,In_2195,In_4059);
and U3162 (N_3162,In_4595,In_2180);
nor U3163 (N_3163,In_387,In_2670);
nor U3164 (N_3164,In_2075,In_456);
nor U3165 (N_3165,In_3577,In_3781);
or U3166 (N_3166,In_44,In_622);
nor U3167 (N_3167,In_2927,In_4065);
nor U3168 (N_3168,In_1690,In_86);
nand U3169 (N_3169,In_4708,In_2458);
and U3170 (N_3170,In_169,In_4774);
xnor U3171 (N_3171,In_3015,In_3500);
nor U3172 (N_3172,In_316,In_3164);
nor U3173 (N_3173,In_823,In_2523);
and U3174 (N_3174,In_177,In_3212);
nor U3175 (N_3175,In_270,In_2303);
xor U3176 (N_3176,In_3029,In_500);
and U3177 (N_3177,In_4860,In_368);
nor U3178 (N_3178,In_716,In_2567);
xnor U3179 (N_3179,In_3600,In_1178);
nand U3180 (N_3180,In_1370,In_3413);
nor U3181 (N_3181,In_1655,In_1994);
xor U3182 (N_3182,In_4602,In_3051);
or U3183 (N_3183,In_4481,In_163);
nand U3184 (N_3184,In_1546,In_4410);
or U3185 (N_3185,In_695,In_4182);
xor U3186 (N_3186,In_2855,In_956);
nand U3187 (N_3187,In_1951,In_3981);
or U3188 (N_3188,In_4299,In_4717);
nor U3189 (N_3189,In_814,In_863);
xor U3190 (N_3190,In_321,In_2424);
and U3191 (N_3191,In_3506,In_3513);
nor U3192 (N_3192,In_777,In_2263);
nand U3193 (N_3193,In_2060,In_4710);
nor U3194 (N_3194,In_3530,In_198);
and U3195 (N_3195,In_913,In_2844);
nor U3196 (N_3196,In_693,In_4928);
nor U3197 (N_3197,In_3234,In_871);
or U3198 (N_3198,In_422,In_644);
xnor U3199 (N_3199,In_3880,In_3613);
or U3200 (N_3200,In_2576,In_4707);
or U3201 (N_3201,In_3629,In_3599);
nand U3202 (N_3202,In_1141,In_1351);
and U3203 (N_3203,In_3292,In_1937);
xor U3204 (N_3204,In_2815,In_3947);
xnor U3205 (N_3205,In_3994,In_4810);
nor U3206 (N_3206,In_893,In_1916);
nand U3207 (N_3207,In_4794,In_3715);
nor U3208 (N_3208,In_167,In_4466);
or U3209 (N_3209,In_2927,In_2736);
nand U3210 (N_3210,In_4405,In_1808);
or U3211 (N_3211,In_3657,In_4029);
nor U3212 (N_3212,In_415,In_974);
nand U3213 (N_3213,In_3865,In_3007);
and U3214 (N_3214,In_2834,In_4666);
xor U3215 (N_3215,In_79,In_569);
nand U3216 (N_3216,In_2198,In_912);
nor U3217 (N_3217,In_4885,In_3650);
xnor U3218 (N_3218,In_3347,In_1633);
and U3219 (N_3219,In_2183,In_4416);
nor U3220 (N_3220,In_903,In_4858);
and U3221 (N_3221,In_3292,In_684);
nand U3222 (N_3222,In_4652,In_2110);
xor U3223 (N_3223,In_4954,In_3921);
or U3224 (N_3224,In_388,In_3855);
xnor U3225 (N_3225,In_2843,In_1378);
xor U3226 (N_3226,In_4898,In_66);
and U3227 (N_3227,In_4169,In_786);
nand U3228 (N_3228,In_1903,In_4172);
xnor U3229 (N_3229,In_730,In_4886);
nor U3230 (N_3230,In_314,In_1265);
nand U3231 (N_3231,In_616,In_3703);
nor U3232 (N_3232,In_1556,In_1711);
or U3233 (N_3233,In_3770,In_1724);
nand U3234 (N_3234,In_2348,In_1792);
xnor U3235 (N_3235,In_1665,In_2183);
xnor U3236 (N_3236,In_4591,In_325);
nand U3237 (N_3237,In_1313,In_1711);
or U3238 (N_3238,In_4218,In_1629);
or U3239 (N_3239,In_4673,In_2850);
nand U3240 (N_3240,In_4742,In_4921);
and U3241 (N_3241,In_4472,In_1506);
and U3242 (N_3242,In_59,In_1792);
or U3243 (N_3243,In_1589,In_1887);
nand U3244 (N_3244,In_430,In_4361);
and U3245 (N_3245,In_4046,In_2210);
nand U3246 (N_3246,In_3164,In_1489);
nor U3247 (N_3247,In_4823,In_3883);
and U3248 (N_3248,In_3812,In_2682);
xnor U3249 (N_3249,In_2205,In_4010);
or U3250 (N_3250,In_3602,In_3509);
nor U3251 (N_3251,In_3897,In_3041);
nor U3252 (N_3252,In_2441,In_4158);
and U3253 (N_3253,In_3325,In_2446);
xnor U3254 (N_3254,In_2162,In_4859);
or U3255 (N_3255,In_3388,In_4415);
xor U3256 (N_3256,In_1689,In_1647);
or U3257 (N_3257,In_2992,In_4021);
nand U3258 (N_3258,In_667,In_3433);
xnor U3259 (N_3259,In_171,In_3592);
or U3260 (N_3260,In_3556,In_1100);
nand U3261 (N_3261,In_282,In_916);
nor U3262 (N_3262,In_2715,In_3189);
nor U3263 (N_3263,In_2610,In_4254);
nor U3264 (N_3264,In_1413,In_738);
or U3265 (N_3265,In_4443,In_4244);
or U3266 (N_3266,In_411,In_1505);
xnor U3267 (N_3267,In_4973,In_3892);
or U3268 (N_3268,In_2750,In_1891);
nand U3269 (N_3269,In_786,In_1754);
nor U3270 (N_3270,In_3264,In_3666);
and U3271 (N_3271,In_4698,In_344);
and U3272 (N_3272,In_3997,In_4043);
or U3273 (N_3273,In_1846,In_1593);
xor U3274 (N_3274,In_3481,In_2409);
and U3275 (N_3275,In_4245,In_1749);
nand U3276 (N_3276,In_67,In_550);
nand U3277 (N_3277,In_1321,In_1879);
nand U3278 (N_3278,In_920,In_937);
nand U3279 (N_3279,In_4607,In_4647);
and U3280 (N_3280,In_626,In_4403);
or U3281 (N_3281,In_4930,In_636);
or U3282 (N_3282,In_2344,In_3970);
xnor U3283 (N_3283,In_3643,In_25);
nor U3284 (N_3284,In_1892,In_304);
or U3285 (N_3285,In_4853,In_4808);
xnor U3286 (N_3286,In_629,In_2175);
nor U3287 (N_3287,In_614,In_837);
nand U3288 (N_3288,In_4773,In_4992);
and U3289 (N_3289,In_88,In_1894);
nand U3290 (N_3290,In_2982,In_4787);
nor U3291 (N_3291,In_4230,In_3002);
nand U3292 (N_3292,In_3750,In_4765);
and U3293 (N_3293,In_4335,In_3514);
or U3294 (N_3294,In_1134,In_4353);
or U3295 (N_3295,In_4689,In_3652);
and U3296 (N_3296,In_131,In_1624);
nor U3297 (N_3297,In_604,In_1252);
nand U3298 (N_3298,In_1919,In_421);
xor U3299 (N_3299,In_2225,In_4033);
nor U3300 (N_3300,In_3752,In_951);
and U3301 (N_3301,In_261,In_4132);
nand U3302 (N_3302,In_4270,In_1523);
xnor U3303 (N_3303,In_2757,In_4488);
nor U3304 (N_3304,In_632,In_3027);
xnor U3305 (N_3305,In_1906,In_3079);
nand U3306 (N_3306,In_3941,In_3944);
and U3307 (N_3307,In_1046,In_2835);
and U3308 (N_3308,In_1337,In_2323);
or U3309 (N_3309,In_2827,In_4322);
nor U3310 (N_3310,In_1010,In_4798);
xor U3311 (N_3311,In_388,In_4090);
or U3312 (N_3312,In_108,In_1052);
xnor U3313 (N_3313,In_3925,In_77);
nor U3314 (N_3314,In_2807,In_218);
nand U3315 (N_3315,In_2756,In_825);
xnor U3316 (N_3316,In_1389,In_1604);
xor U3317 (N_3317,In_2617,In_4402);
nor U3318 (N_3318,In_4821,In_4319);
or U3319 (N_3319,In_2847,In_1179);
nor U3320 (N_3320,In_4311,In_3285);
xor U3321 (N_3321,In_3772,In_2588);
nor U3322 (N_3322,In_3466,In_3783);
xor U3323 (N_3323,In_4143,In_2170);
nor U3324 (N_3324,In_4485,In_658);
and U3325 (N_3325,In_1964,In_1698);
nor U3326 (N_3326,In_2084,In_173);
or U3327 (N_3327,In_2051,In_2102);
and U3328 (N_3328,In_2549,In_4704);
xnor U3329 (N_3329,In_4369,In_390);
xnor U3330 (N_3330,In_4401,In_1560);
xnor U3331 (N_3331,In_2075,In_1459);
nor U3332 (N_3332,In_674,In_1300);
and U3333 (N_3333,In_4510,In_1121);
or U3334 (N_3334,In_4463,In_1137);
nand U3335 (N_3335,In_1761,In_4360);
or U3336 (N_3336,In_4195,In_4398);
nor U3337 (N_3337,In_3367,In_3609);
or U3338 (N_3338,In_4855,In_643);
nand U3339 (N_3339,In_1486,In_2241);
nand U3340 (N_3340,In_3694,In_2982);
xor U3341 (N_3341,In_436,In_2821);
or U3342 (N_3342,In_1972,In_4877);
xor U3343 (N_3343,In_1593,In_4500);
nand U3344 (N_3344,In_3799,In_3302);
nor U3345 (N_3345,In_3818,In_2834);
nand U3346 (N_3346,In_1591,In_709);
nor U3347 (N_3347,In_4042,In_1140);
or U3348 (N_3348,In_1882,In_2067);
or U3349 (N_3349,In_4321,In_362);
or U3350 (N_3350,In_873,In_2337);
nor U3351 (N_3351,In_1079,In_3161);
nor U3352 (N_3352,In_4125,In_1624);
xnor U3353 (N_3353,In_3754,In_4392);
and U3354 (N_3354,In_2462,In_2247);
and U3355 (N_3355,In_3634,In_3319);
or U3356 (N_3356,In_4889,In_2645);
xnor U3357 (N_3357,In_3963,In_4899);
nand U3358 (N_3358,In_4553,In_4683);
nand U3359 (N_3359,In_651,In_3115);
nor U3360 (N_3360,In_732,In_3989);
nand U3361 (N_3361,In_3382,In_377);
xnor U3362 (N_3362,In_1598,In_4466);
or U3363 (N_3363,In_2720,In_1687);
nor U3364 (N_3364,In_102,In_4377);
or U3365 (N_3365,In_1496,In_1919);
nor U3366 (N_3366,In_1149,In_4156);
xnor U3367 (N_3367,In_3235,In_3743);
and U3368 (N_3368,In_3836,In_3171);
xnor U3369 (N_3369,In_2428,In_1725);
and U3370 (N_3370,In_1911,In_2297);
or U3371 (N_3371,In_589,In_3438);
nand U3372 (N_3372,In_3975,In_4835);
nand U3373 (N_3373,In_2775,In_2908);
xnor U3374 (N_3374,In_4454,In_547);
and U3375 (N_3375,In_2333,In_1416);
and U3376 (N_3376,In_2701,In_306);
xnor U3377 (N_3377,In_2770,In_3105);
xor U3378 (N_3378,In_889,In_4806);
nand U3379 (N_3379,In_861,In_3688);
nor U3380 (N_3380,In_4190,In_1121);
nor U3381 (N_3381,In_895,In_1162);
xnor U3382 (N_3382,In_4736,In_1854);
or U3383 (N_3383,In_4499,In_3899);
nand U3384 (N_3384,In_3841,In_3930);
xnor U3385 (N_3385,In_2333,In_1961);
and U3386 (N_3386,In_4041,In_3473);
xnor U3387 (N_3387,In_1089,In_3288);
nor U3388 (N_3388,In_826,In_3518);
or U3389 (N_3389,In_4598,In_3256);
and U3390 (N_3390,In_4381,In_1992);
nand U3391 (N_3391,In_1210,In_1941);
nand U3392 (N_3392,In_2532,In_4679);
nor U3393 (N_3393,In_1988,In_1400);
xor U3394 (N_3394,In_539,In_2805);
xnor U3395 (N_3395,In_1052,In_4107);
xor U3396 (N_3396,In_4977,In_1581);
or U3397 (N_3397,In_1362,In_2748);
and U3398 (N_3398,In_2399,In_1920);
nand U3399 (N_3399,In_742,In_431);
and U3400 (N_3400,In_945,In_1745);
nor U3401 (N_3401,In_2238,In_4551);
and U3402 (N_3402,In_1640,In_306);
xnor U3403 (N_3403,In_3128,In_1635);
nand U3404 (N_3404,In_2769,In_667);
or U3405 (N_3405,In_4853,In_65);
or U3406 (N_3406,In_4508,In_2432);
xor U3407 (N_3407,In_4029,In_793);
nand U3408 (N_3408,In_4726,In_4740);
nor U3409 (N_3409,In_4176,In_2748);
nand U3410 (N_3410,In_4752,In_48);
nand U3411 (N_3411,In_912,In_3342);
nand U3412 (N_3412,In_593,In_3032);
nor U3413 (N_3413,In_666,In_261);
nor U3414 (N_3414,In_14,In_4861);
xnor U3415 (N_3415,In_952,In_486);
nand U3416 (N_3416,In_696,In_2942);
or U3417 (N_3417,In_2234,In_2010);
and U3418 (N_3418,In_2510,In_259);
nor U3419 (N_3419,In_1225,In_659);
xor U3420 (N_3420,In_2682,In_131);
and U3421 (N_3421,In_3776,In_2257);
nand U3422 (N_3422,In_732,In_853);
nand U3423 (N_3423,In_4390,In_956);
nand U3424 (N_3424,In_1034,In_752);
nor U3425 (N_3425,In_4303,In_3810);
nor U3426 (N_3426,In_3697,In_2712);
or U3427 (N_3427,In_2031,In_4805);
nor U3428 (N_3428,In_1639,In_284);
nand U3429 (N_3429,In_4561,In_82);
nand U3430 (N_3430,In_1521,In_388);
nor U3431 (N_3431,In_1267,In_2633);
and U3432 (N_3432,In_4259,In_3371);
or U3433 (N_3433,In_801,In_313);
or U3434 (N_3434,In_1646,In_3589);
nand U3435 (N_3435,In_4500,In_2149);
nor U3436 (N_3436,In_3999,In_3830);
and U3437 (N_3437,In_4673,In_1504);
nand U3438 (N_3438,In_225,In_4772);
or U3439 (N_3439,In_3878,In_3449);
nor U3440 (N_3440,In_4642,In_3715);
and U3441 (N_3441,In_32,In_4050);
xnor U3442 (N_3442,In_48,In_1607);
and U3443 (N_3443,In_2769,In_3175);
and U3444 (N_3444,In_3130,In_2289);
nand U3445 (N_3445,In_2243,In_2872);
nor U3446 (N_3446,In_3314,In_1436);
nand U3447 (N_3447,In_3878,In_1620);
and U3448 (N_3448,In_4893,In_1536);
or U3449 (N_3449,In_1431,In_3547);
nand U3450 (N_3450,In_392,In_1263);
nand U3451 (N_3451,In_2497,In_4508);
and U3452 (N_3452,In_3966,In_2390);
or U3453 (N_3453,In_2736,In_926);
and U3454 (N_3454,In_1139,In_249);
or U3455 (N_3455,In_1593,In_4412);
xnor U3456 (N_3456,In_1402,In_2489);
and U3457 (N_3457,In_581,In_697);
xor U3458 (N_3458,In_945,In_3113);
nor U3459 (N_3459,In_929,In_3215);
xor U3460 (N_3460,In_1285,In_2604);
and U3461 (N_3461,In_1058,In_2136);
and U3462 (N_3462,In_964,In_4240);
nor U3463 (N_3463,In_3081,In_3545);
and U3464 (N_3464,In_943,In_4792);
xor U3465 (N_3465,In_4195,In_4039);
nor U3466 (N_3466,In_427,In_2989);
or U3467 (N_3467,In_971,In_311);
xnor U3468 (N_3468,In_3208,In_4875);
or U3469 (N_3469,In_1818,In_2121);
nor U3470 (N_3470,In_2561,In_34);
xnor U3471 (N_3471,In_946,In_579);
nor U3472 (N_3472,In_2316,In_322);
and U3473 (N_3473,In_4256,In_1868);
nand U3474 (N_3474,In_2789,In_807);
or U3475 (N_3475,In_2044,In_3874);
and U3476 (N_3476,In_3579,In_3719);
xnor U3477 (N_3477,In_4517,In_4540);
or U3478 (N_3478,In_3198,In_2973);
or U3479 (N_3479,In_1104,In_3146);
nand U3480 (N_3480,In_4126,In_2130);
nor U3481 (N_3481,In_821,In_2316);
or U3482 (N_3482,In_4277,In_2871);
or U3483 (N_3483,In_1499,In_3268);
xnor U3484 (N_3484,In_2872,In_3736);
and U3485 (N_3485,In_3887,In_4377);
nor U3486 (N_3486,In_1621,In_3806);
nand U3487 (N_3487,In_4310,In_1939);
nand U3488 (N_3488,In_3466,In_175);
nor U3489 (N_3489,In_4844,In_2478);
or U3490 (N_3490,In_4106,In_4776);
nor U3491 (N_3491,In_4025,In_3314);
or U3492 (N_3492,In_4298,In_349);
nand U3493 (N_3493,In_3869,In_4307);
xnor U3494 (N_3494,In_746,In_4198);
xnor U3495 (N_3495,In_2151,In_757);
and U3496 (N_3496,In_3773,In_243);
or U3497 (N_3497,In_4992,In_4530);
nor U3498 (N_3498,In_4445,In_3751);
xor U3499 (N_3499,In_2077,In_2119);
nor U3500 (N_3500,In_3388,In_4896);
xor U3501 (N_3501,In_1876,In_171);
and U3502 (N_3502,In_1046,In_3915);
xor U3503 (N_3503,In_1385,In_2820);
or U3504 (N_3504,In_2185,In_4948);
or U3505 (N_3505,In_1056,In_2742);
and U3506 (N_3506,In_859,In_2825);
nand U3507 (N_3507,In_4662,In_3708);
and U3508 (N_3508,In_2213,In_2884);
or U3509 (N_3509,In_652,In_2027);
xnor U3510 (N_3510,In_2822,In_3186);
nor U3511 (N_3511,In_2492,In_505);
nor U3512 (N_3512,In_3022,In_799);
xnor U3513 (N_3513,In_4928,In_2606);
xor U3514 (N_3514,In_2111,In_733);
and U3515 (N_3515,In_1478,In_1462);
xnor U3516 (N_3516,In_3486,In_3056);
and U3517 (N_3517,In_1423,In_2409);
xor U3518 (N_3518,In_3721,In_2358);
or U3519 (N_3519,In_4271,In_1037);
nor U3520 (N_3520,In_2566,In_701);
xnor U3521 (N_3521,In_16,In_4059);
and U3522 (N_3522,In_2761,In_4684);
xnor U3523 (N_3523,In_3208,In_1421);
nand U3524 (N_3524,In_4109,In_3915);
and U3525 (N_3525,In_4851,In_465);
nor U3526 (N_3526,In_2141,In_4607);
xor U3527 (N_3527,In_4935,In_3211);
or U3528 (N_3528,In_3294,In_2861);
xor U3529 (N_3529,In_2628,In_3814);
nand U3530 (N_3530,In_2823,In_1615);
nor U3531 (N_3531,In_2258,In_4396);
and U3532 (N_3532,In_3105,In_3557);
xor U3533 (N_3533,In_3263,In_2638);
and U3534 (N_3534,In_553,In_424);
xor U3535 (N_3535,In_3507,In_4593);
or U3536 (N_3536,In_3061,In_297);
nand U3537 (N_3537,In_581,In_2746);
or U3538 (N_3538,In_3806,In_2251);
or U3539 (N_3539,In_4371,In_3005);
and U3540 (N_3540,In_2693,In_1704);
xnor U3541 (N_3541,In_1586,In_23);
nand U3542 (N_3542,In_3932,In_1667);
and U3543 (N_3543,In_4768,In_1819);
xnor U3544 (N_3544,In_4694,In_3068);
xnor U3545 (N_3545,In_1116,In_2697);
and U3546 (N_3546,In_840,In_3177);
nor U3547 (N_3547,In_3955,In_3387);
or U3548 (N_3548,In_1011,In_2492);
or U3549 (N_3549,In_159,In_1927);
xor U3550 (N_3550,In_2023,In_4975);
nor U3551 (N_3551,In_2405,In_4899);
xor U3552 (N_3552,In_2387,In_1869);
nor U3553 (N_3553,In_236,In_4273);
or U3554 (N_3554,In_1655,In_483);
nor U3555 (N_3555,In_3838,In_4946);
nor U3556 (N_3556,In_649,In_3719);
or U3557 (N_3557,In_2458,In_3166);
nor U3558 (N_3558,In_2914,In_3722);
nor U3559 (N_3559,In_1234,In_234);
xnor U3560 (N_3560,In_2236,In_4687);
nor U3561 (N_3561,In_1573,In_4852);
or U3562 (N_3562,In_320,In_3295);
xor U3563 (N_3563,In_4439,In_383);
nor U3564 (N_3564,In_429,In_2822);
or U3565 (N_3565,In_4695,In_3458);
nor U3566 (N_3566,In_1534,In_557);
and U3567 (N_3567,In_3632,In_1410);
nand U3568 (N_3568,In_2480,In_4201);
xnor U3569 (N_3569,In_943,In_336);
nor U3570 (N_3570,In_2366,In_3148);
nand U3571 (N_3571,In_759,In_3078);
or U3572 (N_3572,In_4100,In_4625);
nor U3573 (N_3573,In_1934,In_2761);
xor U3574 (N_3574,In_4150,In_4752);
xnor U3575 (N_3575,In_2286,In_1205);
or U3576 (N_3576,In_1734,In_4834);
nand U3577 (N_3577,In_154,In_1769);
or U3578 (N_3578,In_145,In_678);
nor U3579 (N_3579,In_1473,In_184);
xor U3580 (N_3580,In_2455,In_2443);
nor U3581 (N_3581,In_1268,In_3098);
and U3582 (N_3582,In_3030,In_3002);
or U3583 (N_3583,In_669,In_4002);
and U3584 (N_3584,In_1325,In_1988);
and U3585 (N_3585,In_3475,In_3455);
or U3586 (N_3586,In_3662,In_4090);
xor U3587 (N_3587,In_3149,In_2599);
xor U3588 (N_3588,In_4524,In_2358);
xor U3589 (N_3589,In_3366,In_4346);
and U3590 (N_3590,In_661,In_2138);
nor U3591 (N_3591,In_2395,In_3650);
or U3592 (N_3592,In_2751,In_2480);
nor U3593 (N_3593,In_4802,In_3885);
xor U3594 (N_3594,In_213,In_3421);
nor U3595 (N_3595,In_4408,In_672);
and U3596 (N_3596,In_4251,In_2632);
or U3597 (N_3597,In_991,In_2253);
nand U3598 (N_3598,In_4457,In_340);
or U3599 (N_3599,In_3058,In_3278);
nand U3600 (N_3600,In_3911,In_572);
or U3601 (N_3601,In_3963,In_3200);
or U3602 (N_3602,In_1346,In_4506);
xor U3603 (N_3603,In_3340,In_289);
or U3604 (N_3604,In_2564,In_2990);
and U3605 (N_3605,In_3698,In_198);
and U3606 (N_3606,In_2032,In_75);
xor U3607 (N_3607,In_2453,In_3905);
xor U3608 (N_3608,In_2509,In_501);
or U3609 (N_3609,In_4499,In_257);
and U3610 (N_3610,In_4899,In_3259);
nor U3611 (N_3611,In_3874,In_3315);
xor U3612 (N_3612,In_4963,In_1692);
xnor U3613 (N_3613,In_233,In_1120);
nor U3614 (N_3614,In_1760,In_3665);
and U3615 (N_3615,In_696,In_447);
or U3616 (N_3616,In_2153,In_2784);
nor U3617 (N_3617,In_1612,In_1056);
and U3618 (N_3618,In_919,In_461);
xnor U3619 (N_3619,In_4494,In_1026);
nand U3620 (N_3620,In_2727,In_4749);
nand U3621 (N_3621,In_4639,In_3609);
xnor U3622 (N_3622,In_2106,In_4364);
or U3623 (N_3623,In_3744,In_1764);
nor U3624 (N_3624,In_4762,In_643);
nor U3625 (N_3625,In_531,In_3382);
xor U3626 (N_3626,In_638,In_3741);
or U3627 (N_3627,In_792,In_1446);
nor U3628 (N_3628,In_610,In_1995);
xnor U3629 (N_3629,In_1720,In_2623);
xnor U3630 (N_3630,In_4284,In_1428);
or U3631 (N_3631,In_520,In_685);
nor U3632 (N_3632,In_1963,In_2384);
nand U3633 (N_3633,In_1698,In_741);
nand U3634 (N_3634,In_2792,In_2346);
and U3635 (N_3635,In_665,In_2130);
and U3636 (N_3636,In_2449,In_4489);
nor U3637 (N_3637,In_36,In_35);
nand U3638 (N_3638,In_3024,In_1346);
nor U3639 (N_3639,In_351,In_817);
nor U3640 (N_3640,In_3009,In_4706);
nor U3641 (N_3641,In_1880,In_2250);
nand U3642 (N_3642,In_1965,In_1641);
and U3643 (N_3643,In_3945,In_1448);
and U3644 (N_3644,In_513,In_4526);
nor U3645 (N_3645,In_2896,In_3878);
nor U3646 (N_3646,In_48,In_761);
nor U3647 (N_3647,In_1674,In_3768);
and U3648 (N_3648,In_4547,In_4962);
xor U3649 (N_3649,In_1386,In_4069);
xor U3650 (N_3650,In_2988,In_3251);
nor U3651 (N_3651,In_3497,In_2756);
nand U3652 (N_3652,In_1275,In_22);
xnor U3653 (N_3653,In_2631,In_2792);
or U3654 (N_3654,In_92,In_1821);
nor U3655 (N_3655,In_1680,In_4572);
and U3656 (N_3656,In_2787,In_1771);
xnor U3657 (N_3657,In_4403,In_1736);
or U3658 (N_3658,In_4804,In_427);
xnor U3659 (N_3659,In_1530,In_3271);
and U3660 (N_3660,In_54,In_4685);
xnor U3661 (N_3661,In_104,In_4935);
xor U3662 (N_3662,In_1723,In_1936);
and U3663 (N_3663,In_3085,In_4841);
nor U3664 (N_3664,In_4044,In_2604);
xor U3665 (N_3665,In_2333,In_2422);
xnor U3666 (N_3666,In_3701,In_1186);
or U3667 (N_3667,In_2360,In_879);
or U3668 (N_3668,In_4395,In_4033);
or U3669 (N_3669,In_4994,In_4522);
nor U3670 (N_3670,In_4912,In_2060);
nand U3671 (N_3671,In_2380,In_4451);
or U3672 (N_3672,In_1098,In_2823);
nor U3673 (N_3673,In_652,In_1612);
or U3674 (N_3674,In_1431,In_2976);
xor U3675 (N_3675,In_797,In_3024);
and U3676 (N_3676,In_3350,In_3595);
or U3677 (N_3677,In_1756,In_2899);
and U3678 (N_3678,In_2382,In_4829);
or U3679 (N_3679,In_2108,In_4977);
or U3680 (N_3680,In_22,In_4771);
nor U3681 (N_3681,In_526,In_1018);
xnor U3682 (N_3682,In_4763,In_4142);
xnor U3683 (N_3683,In_4140,In_2194);
or U3684 (N_3684,In_1542,In_4648);
and U3685 (N_3685,In_1837,In_169);
nor U3686 (N_3686,In_2354,In_1401);
and U3687 (N_3687,In_4701,In_3368);
or U3688 (N_3688,In_3584,In_4831);
and U3689 (N_3689,In_699,In_3477);
and U3690 (N_3690,In_4927,In_135);
or U3691 (N_3691,In_593,In_1928);
xnor U3692 (N_3692,In_4702,In_4078);
nor U3693 (N_3693,In_430,In_2805);
nand U3694 (N_3694,In_2385,In_3718);
or U3695 (N_3695,In_1819,In_3);
or U3696 (N_3696,In_2924,In_1005);
and U3697 (N_3697,In_4675,In_39);
or U3698 (N_3698,In_600,In_4769);
xnor U3699 (N_3699,In_2485,In_834);
nand U3700 (N_3700,In_1497,In_4498);
xnor U3701 (N_3701,In_2632,In_131);
xnor U3702 (N_3702,In_3252,In_3309);
and U3703 (N_3703,In_1793,In_2675);
or U3704 (N_3704,In_2074,In_1397);
nand U3705 (N_3705,In_4528,In_2700);
nand U3706 (N_3706,In_3214,In_3158);
or U3707 (N_3707,In_4176,In_351);
xnor U3708 (N_3708,In_2907,In_1705);
and U3709 (N_3709,In_4008,In_2218);
or U3710 (N_3710,In_2442,In_3525);
xnor U3711 (N_3711,In_2966,In_3432);
and U3712 (N_3712,In_3762,In_1416);
or U3713 (N_3713,In_1033,In_2037);
nand U3714 (N_3714,In_2963,In_4667);
nand U3715 (N_3715,In_4692,In_3229);
nor U3716 (N_3716,In_1594,In_1766);
nor U3717 (N_3717,In_4547,In_4489);
or U3718 (N_3718,In_356,In_4296);
xor U3719 (N_3719,In_2652,In_2712);
nor U3720 (N_3720,In_626,In_3429);
nand U3721 (N_3721,In_2344,In_305);
nand U3722 (N_3722,In_3965,In_3151);
nand U3723 (N_3723,In_3766,In_764);
or U3724 (N_3724,In_1512,In_710);
and U3725 (N_3725,In_1468,In_1521);
or U3726 (N_3726,In_3308,In_1568);
xnor U3727 (N_3727,In_3054,In_154);
and U3728 (N_3728,In_291,In_4610);
and U3729 (N_3729,In_4666,In_2397);
nand U3730 (N_3730,In_1797,In_518);
and U3731 (N_3731,In_1522,In_2043);
or U3732 (N_3732,In_3600,In_1037);
nand U3733 (N_3733,In_1264,In_2854);
nand U3734 (N_3734,In_2985,In_4942);
nand U3735 (N_3735,In_4816,In_2914);
or U3736 (N_3736,In_453,In_22);
or U3737 (N_3737,In_2074,In_4085);
and U3738 (N_3738,In_3834,In_3148);
and U3739 (N_3739,In_4858,In_1218);
or U3740 (N_3740,In_4471,In_2543);
or U3741 (N_3741,In_2963,In_1237);
or U3742 (N_3742,In_187,In_368);
nor U3743 (N_3743,In_2916,In_1568);
nand U3744 (N_3744,In_166,In_4535);
and U3745 (N_3745,In_4508,In_1023);
or U3746 (N_3746,In_2226,In_4692);
or U3747 (N_3747,In_144,In_3166);
and U3748 (N_3748,In_3955,In_4550);
or U3749 (N_3749,In_3334,In_462);
nor U3750 (N_3750,In_3082,In_1406);
or U3751 (N_3751,In_1552,In_4798);
xor U3752 (N_3752,In_97,In_1816);
nor U3753 (N_3753,In_1122,In_1422);
nor U3754 (N_3754,In_1315,In_2856);
nand U3755 (N_3755,In_3781,In_844);
or U3756 (N_3756,In_4456,In_3223);
or U3757 (N_3757,In_3448,In_2524);
nand U3758 (N_3758,In_432,In_1539);
and U3759 (N_3759,In_1145,In_2266);
and U3760 (N_3760,In_2010,In_1639);
and U3761 (N_3761,In_2291,In_4581);
xnor U3762 (N_3762,In_3193,In_4323);
xor U3763 (N_3763,In_2546,In_4967);
nor U3764 (N_3764,In_3314,In_1862);
or U3765 (N_3765,In_1491,In_2941);
and U3766 (N_3766,In_3233,In_2159);
xnor U3767 (N_3767,In_496,In_3028);
xnor U3768 (N_3768,In_4650,In_2229);
nand U3769 (N_3769,In_3321,In_855);
xor U3770 (N_3770,In_2128,In_112);
nor U3771 (N_3771,In_204,In_293);
nand U3772 (N_3772,In_4292,In_960);
nor U3773 (N_3773,In_1620,In_3592);
nand U3774 (N_3774,In_670,In_1704);
and U3775 (N_3775,In_2256,In_4657);
xor U3776 (N_3776,In_666,In_1464);
and U3777 (N_3777,In_1531,In_2009);
nor U3778 (N_3778,In_2215,In_4151);
and U3779 (N_3779,In_2882,In_4082);
xor U3780 (N_3780,In_797,In_2327);
nor U3781 (N_3781,In_3164,In_2192);
or U3782 (N_3782,In_3496,In_3291);
or U3783 (N_3783,In_1825,In_3894);
and U3784 (N_3784,In_2533,In_3938);
xor U3785 (N_3785,In_339,In_1788);
and U3786 (N_3786,In_44,In_1021);
nand U3787 (N_3787,In_3558,In_3356);
or U3788 (N_3788,In_1582,In_155);
or U3789 (N_3789,In_2412,In_3980);
nand U3790 (N_3790,In_1559,In_2363);
nand U3791 (N_3791,In_4115,In_681);
or U3792 (N_3792,In_1154,In_666);
nand U3793 (N_3793,In_1303,In_1430);
xor U3794 (N_3794,In_1684,In_287);
and U3795 (N_3795,In_4568,In_229);
nor U3796 (N_3796,In_2844,In_420);
nor U3797 (N_3797,In_4645,In_2287);
or U3798 (N_3798,In_1239,In_4813);
nor U3799 (N_3799,In_3824,In_1571);
or U3800 (N_3800,In_687,In_425);
nor U3801 (N_3801,In_1894,In_4209);
nand U3802 (N_3802,In_221,In_1186);
and U3803 (N_3803,In_2247,In_1853);
nor U3804 (N_3804,In_1845,In_1017);
nand U3805 (N_3805,In_4062,In_3070);
or U3806 (N_3806,In_2754,In_1052);
nor U3807 (N_3807,In_1067,In_211);
and U3808 (N_3808,In_1688,In_422);
or U3809 (N_3809,In_4350,In_679);
xnor U3810 (N_3810,In_2151,In_3264);
and U3811 (N_3811,In_1618,In_3691);
or U3812 (N_3812,In_1733,In_1270);
xor U3813 (N_3813,In_1457,In_4466);
and U3814 (N_3814,In_2451,In_1678);
nor U3815 (N_3815,In_4518,In_380);
or U3816 (N_3816,In_939,In_3524);
or U3817 (N_3817,In_902,In_2934);
and U3818 (N_3818,In_1752,In_2576);
nand U3819 (N_3819,In_812,In_1813);
nand U3820 (N_3820,In_217,In_3370);
nand U3821 (N_3821,In_3036,In_474);
nand U3822 (N_3822,In_1267,In_874);
nand U3823 (N_3823,In_4304,In_106);
nand U3824 (N_3824,In_3307,In_337);
nor U3825 (N_3825,In_856,In_399);
nand U3826 (N_3826,In_3698,In_2044);
and U3827 (N_3827,In_4919,In_1902);
nor U3828 (N_3828,In_4721,In_4518);
xor U3829 (N_3829,In_4845,In_2491);
nor U3830 (N_3830,In_1413,In_1406);
or U3831 (N_3831,In_4872,In_3268);
or U3832 (N_3832,In_4407,In_642);
nor U3833 (N_3833,In_4772,In_2858);
xnor U3834 (N_3834,In_1479,In_3336);
and U3835 (N_3835,In_3316,In_980);
and U3836 (N_3836,In_4256,In_1924);
and U3837 (N_3837,In_1627,In_3223);
and U3838 (N_3838,In_2671,In_2454);
xnor U3839 (N_3839,In_1551,In_3949);
and U3840 (N_3840,In_27,In_3587);
xnor U3841 (N_3841,In_3572,In_3626);
and U3842 (N_3842,In_200,In_2667);
xnor U3843 (N_3843,In_1158,In_2105);
nand U3844 (N_3844,In_622,In_2855);
nand U3845 (N_3845,In_1688,In_2658);
nor U3846 (N_3846,In_2845,In_534);
and U3847 (N_3847,In_4642,In_4575);
or U3848 (N_3848,In_3586,In_2417);
nand U3849 (N_3849,In_4578,In_2841);
nand U3850 (N_3850,In_2391,In_3322);
xnor U3851 (N_3851,In_819,In_2243);
nand U3852 (N_3852,In_1450,In_906);
nor U3853 (N_3853,In_3578,In_1655);
and U3854 (N_3854,In_2877,In_4623);
or U3855 (N_3855,In_2529,In_4381);
or U3856 (N_3856,In_4282,In_272);
nor U3857 (N_3857,In_2281,In_2242);
and U3858 (N_3858,In_2148,In_2215);
nor U3859 (N_3859,In_1078,In_3585);
nor U3860 (N_3860,In_1928,In_3942);
xor U3861 (N_3861,In_3565,In_4517);
and U3862 (N_3862,In_2476,In_3759);
or U3863 (N_3863,In_4524,In_522);
nand U3864 (N_3864,In_1104,In_1245);
nor U3865 (N_3865,In_1783,In_4730);
nand U3866 (N_3866,In_2396,In_3545);
nor U3867 (N_3867,In_4440,In_241);
and U3868 (N_3868,In_416,In_4616);
or U3869 (N_3869,In_1208,In_2032);
or U3870 (N_3870,In_2695,In_2433);
or U3871 (N_3871,In_950,In_4171);
nor U3872 (N_3872,In_75,In_232);
nand U3873 (N_3873,In_2320,In_3018);
xor U3874 (N_3874,In_2300,In_235);
nor U3875 (N_3875,In_4271,In_4824);
xnor U3876 (N_3876,In_1958,In_4379);
nor U3877 (N_3877,In_3400,In_2724);
xor U3878 (N_3878,In_4854,In_4944);
or U3879 (N_3879,In_3500,In_31);
nand U3880 (N_3880,In_530,In_2714);
and U3881 (N_3881,In_2732,In_2715);
or U3882 (N_3882,In_2023,In_4722);
and U3883 (N_3883,In_3955,In_2684);
and U3884 (N_3884,In_2767,In_3408);
nand U3885 (N_3885,In_793,In_3596);
or U3886 (N_3886,In_3306,In_1843);
and U3887 (N_3887,In_4933,In_3626);
and U3888 (N_3888,In_2288,In_2394);
nand U3889 (N_3889,In_4475,In_4851);
nor U3890 (N_3890,In_441,In_397);
or U3891 (N_3891,In_802,In_1744);
nor U3892 (N_3892,In_3113,In_1580);
nand U3893 (N_3893,In_3112,In_3669);
nor U3894 (N_3894,In_3368,In_4413);
nand U3895 (N_3895,In_4394,In_2652);
and U3896 (N_3896,In_1091,In_3004);
nor U3897 (N_3897,In_1749,In_1312);
xor U3898 (N_3898,In_3559,In_2142);
nor U3899 (N_3899,In_1701,In_4360);
and U3900 (N_3900,In_412,In_1884);
nor U3901 (N_3901,In_1687,In_3263);
xnor U3902 (N_3902,In_2930,In_4511);
and U3903 (N_3903,In_1332,In_3750);
and U3904 (N_3904,In_2814,In_355);
or U3905 (N_3905,In_738,In_1119);
or U3906 (N_3906,In_3755,In_109);
or U3907 (N_3907,In_1162,In_286);
and U3908 (N_3908,In_692,In_558);
nor U3909 (N_3909,In_3914,In_2385);
nor U3910 (N_3910,In_4587,In_2947);
or U3911 (N_3911,In_3348,In_2602);
and U3912 (N_3912,In_3924,In_2515);
or U3913 (N_3913,In_1408,In_3691);
or U3914 (N_3914,In_1352,In_624);
and U3915 (N_3915,In_762,In_920);
or U3916 (N_3916,In_2663,In_376);
xnor U3917 (N_3917,In_2449,In_1033);
xor U3918 (N_3918,In_3842,In_1414);
nand U3919 (N_3919,In_3204,In_2291);
nor U3920 (N_3920,In_623,In_3224);
xnor U3921 (N_3921,In_3581,In_2625);
and U3922 (N_3922,In_613,In_4738);
and U3923 (N_3923,In_4853,In_2407);
nor U3924 (N_3924,In_2050,In_4184);
nor U3925 (N_3925,In_3727,In_1662);
or U3926 (N_3926,In_346,In_4186);
xnor U3927 (N_3927,In_182,In_1527);
and U3928 (N_3928,In_1168,In_3261);
or U3929 (N_3929,In_1097,In_2188);
or U3930 (N_3930,In_9,In_661);
or U3931 (N_3931,In_3862,In_1285);
nand U3932 (N_3932,In_1590,In_1960);
nor U3933 (N_3933,In_482,In_2310);
nand U3934 (N_3934,In_3904,In_3217);
or U3935 (N_3935,In_164,In_3742);
nand U3936 (N_3936,In_4279,In_3244);
and U3937 (N_3937,In_2212,In_1967);
nand U3938 (N_3938,In_4656,In_3234);
and U3939 (N_3939,In_3197,In_1801);
xnor U3940 (N_3940,In_4551,In_3123);
or U3941 (N_3941,In_3819,In_4760);
and U3942 (N_3942,In_3999,In_3279);
or U3943 (N_3943,In_480,In_2334);
or U3944 (N_3944,In_44,In_3961);
and U3945 (N_3945,In_1757,In_2998);
and U3946 (N_3946,In_3532,In_1629);
and U3947 (N_3947,In_3755,In_330);
and U3948 (N_3948,In_4749,In_921);
or U3949 (N_3949,In_750,In_1836);
nand U3950 (N_3950,In_3704,In_984);
or U3951 (N_3951,In_2518,In_4078);
nand U3952 (N_3952,In_4330,In_3237);
nor U3953 (N_3953,In_2238,In_3778);
or U3954 (N_3954,In_3621,In_4207);
nand U3955 (N_3955,In_1418,In_3418);
nor U3956 (N_3956,In_857,In_3648);
xor U3957 (N_3957,In_3059,In_3454);
xnor U3958 (N_3958,In_643,In_155);
xnor U3959 (N_3959,In_2455,In_3700);
xor U3960 (N_3960,In_1738,In_1775);
nand U3961 (N_3961,In_4843,In_3245);
or U3962 (N_3962,In_3779,In_2930);
xnor U3963 (N_3963,In_3490,In_161);
and U3964 (N_3964,In_769,In_3964);
or U3965 (N_3965,In_3304,In_1465);
and U3966 (N_3966,In_3408,In_591);
and U3967 (N_3967,In_3387,In_2646);
or U3968 (N_3968,In_3235,In_2741);
and U3969 (N_3969,In_4415,In_4723);
and U3970 (N_3970,In_4616,In_4333);
nor U3971 (N_3971,In_190,In_2358);
xnor U3972 (N_3972,In_635,In_4885);
nor U3973 (N_3973,In_2227,In_4006);
nand U3974 (N_3974,In_4198,In_891);
or U3975 (N_3975,In_1766,In_3829);
and U3976 (N_3976,In_3719,In_326);
nor U3977 (N_3977,In_2060,In_856);
or U3978 (N_3978,In_55,In_1502);
nor U3979 (N_3979,In_4628,In_4447);
or U3980 (N_3980,In_2171,In_4665);
or U3981 (N_3981,In_1409,In_152);
nand U3982 (N_3982,In_3654,In_2482);
xnor U3983 (N_3983,In_96,In_4804);
or U3984 (N_3984,In_4281,In_4772);
xor U3985 (N_3985,In_741,In_2294);
and U3986 (N_3986,In_3072,In_1143);
nor U3987 (N_3987,In_670,In_3758);
nor U3988 (N_3988,In_436,In_1491);
xnor U3989 (N_3989,In_2458,In_4193);
or U3990 (N_3990,In_3776,In_2417);
xnor U3991 (N_3991,In_2567,In_3868);
and U3992 (N_3992,In_2571,In_2252);
nor U3993 (N_3993,In_4318,In_2629);
xnor U3994 (N_3994,In_478,In_3652);
nand U3995 (N_3995,In_1122,In_768);
and U3996 (N_3996,In_2592,In_1269);
or U3997 (N_3997,In_4323,In_126);
and U3998 (N_3998,In_3957,In_3831);
xor U3999 (N_3999,In_4638,In_3055);
and U4000 (N_4000,In_559,In_2956);
nor U4001 (N_4001,In_1014,In_1259);
nor U4002 (N_4002,In_242,In_4365);
xnor U4003 (N_4003,In_4003,In_3285);
nand U4004 (N_4004,In_1094,In_4204);
nor U4005 (N_4005,In_2293,In_1578);
and U4006 (N_4006,In_792,In_2219);
and U4007 (N_4007,In_2662,In_4957);
xor U4008 (N_4008,In_1985,In_2080);
nand U4009 (N_4009,In_2961,In_2971);
and U4010 (N_4010,In_47,In_3455);
or U4011 (N_4011,In_2778,In_4770);
nor U4012 (N_4012,In_3082,In_4734);
and U4013 (N_4013,In_3614,In_2420);
nand U4014 (N_4014,In_1337,In_3307);
nor U4015 (N_4015,In_3936,In_4634);
or U4016 (N_4016,In_3049,In_1449);
or U4017 (N_4017,In_4904,In_4635);
nand U4018 (N_4018,In_3820,In_1992);
nor U4019 (N_4019,In_1358,In_466);
or U4020 (N_4020,In_1318,In_264);
and U4021 (N_4021,In_2932,In_59);
nand U4022 (N_4022,In_2176,In_1652);
or U4023 (N_4023,In_1931,In_770);
or U4024 (N_4024,In_2179,In_4151);
or U4025 (N_4025,In_748,In_1133);
nand U4026 (N_4026,In_923,In_584);
nor U4027 (N_4027,In_981,In_661);
xor U4028 (N_4028,In_1759,In_4048);
and U4029 (N_4029,In_1211,In_1855);
or U4030 (N_4030,In_3695,In_522);
nand U4031 (N_4031,In_1709,In_3445);
and U4032 (N_4032,In_4788,In_2233);
and U4033 (N_4033,In_4207,In_1966);
xor U4034 (N_4034,In_3393,In_2549);
and U4035 (N_4035,In_4125,In_2003);
nand U4036 (N_4036,In_707,In_516);
nand U4037 (N_4037,In_2310,In_3817);
and U4038 (N_4038,In_3502,In_3356);
nor U4039 (N_4039,In_606,In_4350);
nand U4040 (N_4040,In_4269,In_1044);
and U4041 (N_4041,In_2175,In_3099);
and U4042 (N_4042,In_2533,In_2818);
xor U4043 (N_4043,In_1133,In_619);
xor U4044 (N_4044,In_2164,In_2527);
nand U4045 (N_4045,In_3801,In_3248);
xnor U4046 (N_4046,In_2625,In_3446);
nand U4047 (N_4047,In_4807,In_2585);
xor U4048 (N_4048,In_1782,In_4061);
or U4049 (N_4049,In_2393,In_1765);
nand U4050 (N_4050,In_4853,In_1342);
or U4051 (N_4051,In_3208,In_1439);
nor U4052 (N_4052,In_2862,In_242);
and U4053 (N_4053,In_4651,In_2459);
nor U4054 (N_4054,In_610,In_4168);
and U4055 (N_4055,In_3884,In_1199);
nand U4056 (N_4056,In_2688,In_1504);
and U4057 (N_4057,In_3837,In_121);
nand U4058 (N_4058,In_763,In_1626);
or U4059 (N_4059,In_28,In_4224);
and U4060 (N_4060,In_3003,In_4551);
and U4061 (N_4061,In_2959,In_3153);
nor U4062 (N_4062,In_3725,In_2392);
xor U4063 (N_4063,In_4667,In_2566);
xnor U4064 (N_4064,In_587,In_2398);
xnor U4065 (N_4065,In_1686,In_1956);
or U4066 (N_4066,In_4166,In_4649);
nand U4067 (N_4067,In_2966,In_3898);
or U4068 (N_4068,In_1132,In_1361);
xor U4069 (N_4069,In_1436,In_324);
and U4070 (N_4070,In_592,In_96);
nand U4071 (N_4071,In_2461,In_1833);
or U4072 (N_4072,In_3221,In_2700);
xor U4073 (N_4073,In_2168,In_2200);
nand U4074 (N_4074,In_1947,In_432);
and U4075 (N_4075,In_668,In_680);
and U4076 (N_4076,In_86,In_550);
nor U4077 (N_4077,In_742,In_1989);
nand U4078 (N_4078,In_2173,In_4273);
nand U4079 (N_4079,In_245,In_1517);
xor U4080 (N_4080,In_2913,In_3535);
and U4081 (N_4081,In_1948,In_3266);
and U4082 (N_4082,In_2591,In_784);
nand U4083 (N_4083,In_4036,In_418);
nor U4084 (N_4084,In_2230,In_2892);
nor U4085 (N_4085,In_994,In_3566);
nand U4086 (N_4086,In_2828,In_1169);
or U4087 (N_4087,In_4831,In_4810);
or U4088 (N_4088,In_731,In_198);
nor U4089 (N_4089,In_2590,In_2824);
and U4090 (N_4090,In_3747,In_1890);
xor U4091 (N_4091,In_2329,In_4753);
nand U4092 (N_4092,In_3991,In_3561);
or U4093 (N_4093,In_1092,In_3043);
nand U4094 (N_4094,In_1938,In_1351);
or U4095 (N_4095,In_2016,In_3897);
xor U4096 (N_4096,In_3863,In_1339);
nor U4097 (N_4097,In_231,In_194);
or U4098 (N_4098,In_3531,In_920);
nand U4099 (N_4099,In_597,In_778);
nand U4100 (N_4100,In_2607,In_2007);
and U4101 (N_4101,In_3332,In_3016);
or U4102 (N_4102,In_286,In_3971);
nor U4103 (N_4103,In_900,In_1866);
xnor U4104 (N_4104,In_3448,In_3177);
xnor U4105 (N_4105,In_638,In_3223);
and U4106 (N_4106,In_4582,In_520);
nand U4107 (N_4107,In_3993,In_1089);
xnor U4108 (N_4108,In_3052,In_1673);
or U4109 (N_4109,In_1670,In_4819);
or U4110 (N_4110,In_4005,In_826);
xor U4111 (N_4111,In_4594,In_933);
nand U4112 (N_4112,In_1142,In_4885);
or U4113 (N_4113,In_3042,In_279);
or U4114 (N_4114,In_4748,In_2548);
and U4115 (N_4115,In_2286,In_3528);
nor U4116 (N_4116,In_2304,In_216);
nand U4117 (N_4117,In_4084,In_1868);
or U4118 (N_4118,In_3796,In_3842);
xnor U4119 (N_4119,In_248,In_3786);
nand U4120 (N_4120,In_4726,In_2045);
nand U4121 (N_4121,In_3921,In_1138);
nor U4122 (N_4122,In_1047,In_3774);
and U4123 (N_4123,In_4265,In_2972);
and U4124 (N_4124,In_3823,In_2651);
nor U4125 (N_4125,In_787,In_3696);
nand U4126 (N_4126,In_253,In_4960);
xnor U4127 (N_4127,In_1901,In_1740);
xor U4128 (N_4128,In_4731,In_630);
nand U4129 (N_4129,In_4171,In_2084);
nand U4130 (N_4130,In_1309,In_571);
nand U4131 (N_4131,In_4267,In_4747);
nor U4132 (N_4132,In_4565,In_4298);
nor U4133 (N_4133,In_4257,In_2973);
nor U4134 (N_4134,In_732,In_148);
and U4135 (N_4135,In_1861,In_4436);
and U4136 (N_4136,In_1972,In_3497);
nand U4137 (N_4137,In_1646,In_2405);
nand U4138 (N_4138,In_2289,In_1220);
xnor U4139 (N_4139,In_489,In_400);
nand U4140 (N_4140,In_3673,In_962);
nand U4141 (N_4141,In_2312,In_2462);
nand U4142 (N_4142,In_2277,In_4182);
and U4143 (N_4143,In_2448,In_3781);
xor U4144 (N_4144,In_4136,In_3306);
and U4145 (N_4145,In_3174,In_890);
or U4146 (N_4146,In_404,In_3736);
or U4147 (N_4147,In_1859,In_4234);
nand U4148 (N_4148,In_673,In_2948);
or U4149 (N_4149,In_1823,In_629);
xnor U4150 (N_4150,In_3169,In_1318);
nand U4151 (N_4151,In_2311,In_2117);
nand U4152 (N_4152,In_370,In_2367);
xor U4153 (N_4153,In_1855,In_4252);
and U4154 (N_4154,In_1654,In_3644);
nor U4155 (N_4155,In_2747,In_3202);
nand U4156 (N_4156,In_3130,In_2977);
nand U4157 (N_4157,In_2590,In_2678);
or U4158 (N_4158,In_3244,In_3487);
nor U4159 (N_4159,In_4594,In_465);
nor U4160 (N_4160,In_4292,In_3851);
and U4161 (N_4161,In_541,In_4276);
nand U4162 (N_4162,In_3886,In_1544);
nor U4163 (N_4163,In_1073,In_932);
nand U4164 (N_4164,In_2056,In_3992);
and U4165 (N_4165,In_4763,In_4607);
xor U4166 (N_4166,In_1412,In_2321);
and U4167 (N_4167,In_1777,In_4663);
and U4168 (N_4168,In_4825,In_517);
and U4169 (N_4169,In_3481,In_3479);
or U4170 (N_4170,In_3063,In_40);
nand U4171 (N_4171,In_3276,In_1854);
or U4172 (N_4172,In_858,In_2121);
xnor U4173 (N_4173,In_3657,In_3797);
or U4174 (N_4174,In_2906,In_1509);
nand U4175 (N_4175,In_925,In_3962);
and U4176 (N_4176,In_4299,In_4692);
nor U4177 (N_4177,In_3825,In_4811);
or U4178 (N_4178,In_1908,In_1966);
and U4179 (N_4179,In_337,In_3294);
and U4180 (N_4180,In_490,In_223);
xnor U4181 (N_4181,In_4392,In_3723);
or U4182 (N_4182,In_1811,In_2544);
or U4183 (N_4183,In_3731,In_817);
nand U4184 (N_4184,In_2300,In_4724);
or U4185 (N_4185,In_3635,In_1037);
nand U4186 (N_4186,In_4755,In_623);
and U4187 (N_4187,In_2921,In_2305);
nor U4188 (N_4188,In_4470,In_4635);
nor U4189 (N_4189,In_2279,In_4013);
nand U4190 (N_4190,In_2322,In_327);
or U4191 (N_4191,In_874,In_1608);
nand U4192 (N_4192,In_3543,In_4666);
or U4193 (N_4193,In_2527,In_999);
xnor U4194 (N_4194,In_3146,In_703);
nand U4195 (N_4195,In_773,In_3515);
or U4196 (N_4196,In_2811,In_1803);
or U4197 (N_4197,In_4172,In_2642);
nand U4198 (N_4198,In_2111,In_3153);
and U4199 (N_4199,In_1973,In_952);
xor U4200 (N_4200,In_1335,In_3608);
nor U4201 (N_4201,In_3708,In_928);
nand U4202 (N_4202,In_3141,In_1351);
nand U4203 (N_4203,In_2268,In_953);
nand U4204 (N_4204,In_992,In_2281);
and U4205 (N_4205,In_3337,In_1038);
nor U4206 (N_4206,In_1833,In_3861);
nor U4207 (N_4207,In_2955,In_1045);
nand U4208 (N_4208,In_2528,In_4434);
xor U4209 (N_4209,In_761,In_2097);
nand U4210 (N_4210,In_1006,In_2823);
xor U4211 (N_4211,In_4271,In_447);
nor U4212 (N_4212,In_4495,In_381);
nor U4213 (N_4213,In_47,In_2447);
or U4214 (N_4214,In_223,In_2210);
xor U4215 (N_4215,In_4731,In_3159);
nor U4216 (N_4216,In_836,In_737);
and U4217 (N_4217,In_257,In_4375);
and U4218 (N_4218,In_3168,In_257);
or U4219 (N_4219,In_4692,In_3376);
nor U4220 (N_4220,In_3607,In_3552);
and U4221 (N_4221,In_4576,In_1759);
xnor U4222 (N_4222,In_2005,In_3841);
and U4223 (N_4223,In_4492,In_1927);
nand U4224 (N_4224,In_1994,In_3782);
nor U4225 (N_4225,In_866,In_1589);
and U4226 (N_4226,In_4211,In_1828);
nand U4227 (N_4227,In_4916,In_3292);
nor U4228 (N_4228,In_1194,In_4625);
nor U4229 (N_4229,In_1959,In_1260);
nand U4230 (N_4230,In_2017,In_3975);
xor U4231 (N_4231,In_1084,In_21);
nand U4232 (N_4232,In_2159,In_2245);
and U4233 (N_4233,In_4753,In_4192);
and U4234 (N_4234,In_889,In_863);
or U4235 (N_4235,In_1854,In_3909);
and U4236 (N_4236,In_2840,In_3993);
xor U4237 (N_4237,In_418,In_90);
nor U4238 (N_4238,In_191,In_4618);
nor U4239 (N_4239,In_3185,In_4244);
or U4240 (N_4240,In_3676,In_2593);
xnor U4241 (N_4241,In_2833,In_1409);
or U4242 (N_4242,In_3265,In_2853);
xor U4243 (N_4243,In_2789,In_4233);
xor U4244 (N_4244,In_2995,In_4040);
or U4245 (N_4245,In_1442,In_2356);
or U4246 (N_4246,In_2315,In_1972);
xor U4247 (N_4247,In_3613,In_4809);
and U4248 (N_4248,In_1594,In_1086);
or U4249 (N_4249,In_1746,In_4979);
nor U4250 (N_4250,In_3290,In_2243);
xnor U4251 (N_4251,In_3619,In_616);
nor U4252 (N_4252,In_560,In_2460);
and U4253 (N_4253,In_2638,In_2598);
and U4254 (N_4254,In_2835,In_3366);
nand U4255 (N_4255,In_55,In_2784);
nand U4256 (N_4256,In_4970,In_2395);
and U4257 (N_4257,In_1042,In_2621);
xor U4258 (N_4258,In_1928,In_3547);
or U4259 (N_4259,In_3,In_1711);
xnor U4260 (N_4260,In_2662,In_2371);
nand U4261 (N_4261,In_4264,In_3363);
and U4262 (N_4262,In_3755,In_451);
nand U4263 (N_4263,In_4714,In_1052);
nor U4264 (N_4264,In_1925,In_1800);
and U4265 (N_4265,In_1136,In_246);
nand U4266 (N_4266,In_345,In_745);
xnor U4267 (N_4267,In_52,In_3240);
and U4268 (N_4268,In_821,In_3091);
nor U4269 (N_4269,In_4662,In_169);
or U4270 (N_4270,In_4605,In_4861);
or U4271 (N_4271,In_2788,In_1902);
nor U4272 (N_4272,In_4339,In_733);
nand U4273 (N_4273,In_2783,In_4);
and U4274 (N_4274,In_2284,In_2368);
and U4275 (N_4275,In_679,In_570);
xor U4276 (N_4276,In_3328,In_2123);
nand U4277 (N_4277,In_2074,In_2473);
nor U4278 (N_4278,In_3519,In_1915);
and U4279 (N_4279,In_1150,In_4396);
nand U4280 (N_4280,In_4149,In_1029);
or U4281 (N_4281,In_4158,In_3150);
or U4282 (N_4282,In_2678,In_3792);
and U4283 (N_4283,In_2011,In_3773);
and U4284 (N_4284,In_3580,In_2189);
or U4285 (N_4285,In_1636,In_2184);
and U4286 (N_4286,In_1679,In_2906);
and U4287 (N_4287,In_2612,In_4638);
nand U4288 (N_4288,In_1892,In_3981);
nor U4289 (N_4289,In_4521,In_1622);
xor U4290 (N_4290,In_119,In_1417);
and U4291 (N_4291,In_2249,In_3288);
nor U4292 (N_4292,In_1086,In_1461);
or U4293 (N_4293,In_3876,In_1419);
or U4294 (N_4294,In_4080,In_4402);
xor U4295 (N_4295,In_3378,In_1125);
or U4296 (N_4296,In_2616,In_64);
nand U4297 (N_4297,In_3651,In_2317);
xnor U4298 (N_4298,In_4066,In_3644);
xnor U4299 (N_4299,In_4964,In_2066);
or U4300 (N_4300,In_1486,In_4463);
or U4301 (N_4301,In_144,In_1058);
or U4302 (N_4302,In_995,In_915);
nor U4303 (N_4303,In_380,In_1885);
nand U4304 (N_4304,In_2732,In_1086);
or U4305 (N_4305,In_3284,In_4206);
nor U4306 (N_4306,In_4278,In_1344);
or U4307 (N_4307,In_1100,In_4513);
xnor U4308 (N_4308,In_4830,In_3987);
and U4309 (N_4309,In_173,In_4537);
and U4310 (N_4310,In_2967,In_1250);
nand U4311 (N_4311,In_240,In_3326);
nand U4312 (N_4312,In_2584,In_3258);
nand U4313 (N_4313,In_2057,In_2176);
nand U4314 (N_4314,In_111,In_372);
and U4315 (N_4315,In_4483,In_3635);
or U4316 (N_4316,In_3369,In_1111);
and U4317 (N_4317,In_3499,In_4698);
nor U4318 (N_4318,In_3713,In_2752);
or U4319 (N_4319,In_2170,In_579);
and U4320 (N_4320,In_379,In_2691);
or U4321 (N_4321,In_986,In_793);
and U4322 (N_4322,In_1160,In_846);
xnor U4323 (N_4323,In_4007,In_1572);
xor U4324 (N_4324,In_918,In_4680);
and U4325 (N_4325,In_2390,In_692);
nand U4326 (N_4326,In_655,In_4051);
and U4327 (N_4327,In_4007,In_2481);
xnor U4328 (N_4328,In_392,In_1855);
nand U4329 (N_4329,In_4871,In_3145);
nor U4330 (N_4330,In_4547,In_2869);
and U4331 (N_4331,In_364,In_2228);
xnor U4332 (N_4332,In_839,In_274);
nor U4333 (N_4333,In_376,In_378);
nand U4334 (N_4334,In_2198,In_4438);
nor U4335 (N_4335,In_2509,In_2327);
or U4336 (N_4336,In_4575,In_1693);
and U4337 (N_4337,In_2781,In_3091);
nand U4338 (N_4338,In_2266,In_3319);
xnor U4339 (N_4339,In_586,In_537);
nor U4340 (N_4340,In_4436,In_4101);
nor U4341 (N_4341,In_214,In_482);
or U4342 (N_4342,In_4916,In_1181);
and U4343 (N_4343,In_1249,In_2762);
or U4344 (N_4344,In_3442,In_1534);
nand U4345 (N_4345,In_4335,In_4263);
nor U4346 (N_4346,In_4549,In_3160);
or U4347 (N_4347,In_982,In_1995);
or U4348 (N_4348,In_3367,In_113);
nor U4349 (N_4349,In_123,In_626);
nor U4350 (N_4350,In_2099,In_2159);
nand U4351 (N_4351,In_4906,In_488);
nor U4352 (N_4352,In_3127,In_4931);
nor U4353 (N_4353,In_4317,In_1984);
nand U4354 (N_4354,In_1462,In_1545);
nand U4355 (N_4355,In_1425,In_524);
nor U4356 (N_4356,In_1086,In_2355);
nor U4357 (N_4357,In_3355,In_449);
nor U4358 (N_4358,In_1876,In_121);
and U4359 (N_4359,In_481,In_673);
and U4360 (N_4360,In_337,In_561);
and U4361 (N_4361,In_4977,In_2061);
xnor U4362 (N_4362,In_1672,In_4831);
nand U4363 (N_4363,In_2517,In_3075);
or U4364 (N_4364,In_3866,In_1110);
nand U4365 (N_4365,In_1996,In_165);
nor U4366 (N_4366,In_1870,In_4304);
nor U4367 (N_4367,In_4555,In_2424);
xor U4368 (N_4368,In_1847,In_173);
xnor U4369 (N_4369,In_4023,In_4210);
and U4370 (N_4370,In_823,In_4716);
nand U4371 (N_4371,In_1768,In_48);
and U4372 (N_4372,In_1066,In_3334);
or U4373 (N_4373,In_3045,In_3237);
xor U4374 (N_4374,In_2607,In_4103);
and U4375 (N_4375,In_4478,In_119);
xnor U4376 (N_4376,In_1950,In_331);
and U4377 (N_4377,In_4909,In_749);
nor U4378 (N_4378,In_689,In_2725);
nor U4379 (N_4379,In_2040,In_135);
or U4380 (N_4380,In_1341,In_273);
and U4381 (N_4381,In_1919,In_1481);
nor U4382 (N_4382,In_2706,In_3854);
nand U4383 (N_4383,In_2810,In_1493);
and U4384 (N_4384,In_547,In_3484);
and U4385 (N_4385,In_981,In_2212);
nor U4386 (N_4386,In_4340,In_2612);
nand U4387 (N_4387,In_4982,In_4053);
nand U4388 (N_4388,In_3470,In_1686);
xnor U4389 (N_4389,In_1751,In_3726);
nand U4390 (N_4390,In_2441,In_3467);
or U4391 (N_4391,In_564,In_4515);
nor U4392 (N_4392,In_4800,In_2804);
or U4393 (N_4393,In_3784,In_1125);
and U4394 (N_4394,In_2366,In_2584);
and U4395 (N_4395,In_1199,In_420);
and U4396 (N_4396,In_2199,In_442);
and U4397 (N_4397,In_2795,In_4384);
nand U4398 (N_4398,In_4596,In_193);
nor U4399 (N_4399,In_2001,In_620);
and U4400 (N_4400,In_1740,In_4223);
xor U4401 (N_4401,In_3338,In_910);
or U4402 (N_4402,In_3229,In_4984);
nor U4403 (N_4403,In_650,In_413);
xor U4404 (N_4404,In_3456,In_3604);
or U4405 (N_4405,In_4514,In_1079);
or U4406 (N_4406,In_4860,In_3099);
nor U4407 (N_4407,In_3209,In_1178);
nand U4408 (N_4408,In_2024,In_125);
nand U4409 (N_4409,In_4307,In_4148);
xnor U4410 (N_4410,In_3631,In_2326);
or U4411 (N_4411,In_1291,In_1886);
nor U4412 (N_4412,In_4415,In_1436);
xnor U4413 (N_4413,In_3590,In_983);
and U4414 (N_4414,In_413,In_1364);
xnor U4415 (N_4415,In_1239,In_3075);
and U4416 (N_4416,In_895,In_3860);
nor U4417 (N_4417,In_1416,In_1670);
xnor U4418 (N_4418,In_3752,In_2764);
xor U4419 (N_4419,In_4522,In_2048);
xnor U4420 (N_4420,In_1733,In_4419);
or U4421 (N_4421,In_2704,In_2891);
nor U4422 (N_4422,In_3,In_1577);
nor U4423 (N_4423,In_3037,In_3859);
nor U4424 (N_4424,In_2708,In_2273);
nand U4425 (N_4425,In_3592,In_2118);
or U4426 (N_4426,In_3148,In_4718);
nand U4427 (N_4427,In_2084,In_3363);
or U4428 (N_4428,In_114,In_4817);
xor U4429 (N_4429,In_3437,In_4053);
xnor U4430 (N_4430,In_1576,In_1987);
nand U4431 (N_4431,In_3261,In_1999);
and U4432 (N_4432,In_4538,In_2415);
or U4433 (N_4433,In_2177,In_746);
nand U4434 (N_4434,In_3597,In_1813);
and U4435 (N_4435,In_3642,In_633);
and U4436 (N_4436,In_4771,In_2119);
and U4437 (N_4437,In_1724,In_3483);
xor U4438 (N_4438,In_1279,In_2492);
nor U4439 (N_4439,In_2892,In_185);
nor U4440 (N_4440,In_2991,In_1431);
nor U4441 (N_4441,In_315,In_3057);
nor U4442 (N_4442,In_4700,In_0);
or U4443 (N_4443,In_2793,In_923);
and U4444 (N_4444,In_2064,In_1988);
and U4445 (N_4445,In_3713,In_3606);
nand U4446 (N_4446,In_1171,In_556);
nor U4447 (N_4447,In_4345,In_523);
and U4448 (N_4448,In_2491,In_946);
nor U4449 (N_4449,In_1499,In_2694);
or U4450 (N_4450,In_1685,In_2661);
xnor U4451 (N_4451,In_19,In_3844);
xnor U4452 (N_4452,In_2541,In_1867);
and U4453 (N_4453,In_3196,In_683);
xor U4454 (N_4454,In_3774,In_2523);
xor U4455 (N_4455,In_3302,In_3231);
nor U4456 (N_4456,In_2647,In_2245);
xnor U4457 (N_4457,In_1793,In_4455);
nand U4458 (N_4458,In_2006,In_294);
or U4459 (N_4459,In_3251,In_767);
and U4460 (N_4460,In_2788,In_3027);
xnor U4461 (N_4461,In_1160,In_3311);
or U4462 (N_4462,In_2769,In_149);
nand U4463 (N_4463,In_1013,In_4816);
nor U4464 (N_4464,In_4595,In_1333);
and U4465 (N_4465,In_2741,In_4173);
nor U4466 (N_4466,In_4290,In_4486);
and U4467 (N_4467,In_238,In_1002);
or U4468 (N_4468,In_2504,In_1671);
nand U4469 (N_4469,In_2630,In_2603);
nand U4470 (N_4470,In_469,In_2694);
nand U4471 (N_4471,In_1154,In_2016);
nand U4472 (N_4472,In_3248,In_1954);
and U4473 (N_4473,In_806,In_3951);
nor U4474 (N_4474,In_4940,In_1182);
xor U4475 (N_4475,In_4125,In_2076);
or U4476 (N_4476,In_2061,In_4211);
nor U4477 (N_4477,In_2717,In_1305);
nand U4478 (N_4478,In_4362,In_1138);
or U4479 (N_4479,In_520,In_564);
nand U4480 (N_4480,In_1240,In_3525);
or U4481 (N_4481,In_1749,In_4355);
nand U4482 (N_4482,In_1555,In_2598);
nand U4483 (N_4483,In_2030,In_4519);
or U4484 (N_4484,In_2243,In_1702);
nor U4485 (N_4485,In_3040,In_1428);
nand U4486 (N_4486,In_3673,In_2634);
and U4487 (N_4487,In_859,In_4288);
and U4488 (N_4488,In_529,In_2485);
and U4489 (N_4489,In_2631,In_782);
nor U4490 (N_4490,In_3080,In_3665);
nor U4491 (N_4491,In_851,In_972);
nand U4492 (N_4492,In_782,In_2110);
nor U4493 (N_4493,In_2084,In_483);
and U4494 (N_4494,In_2609,In_2476);
and U4495 (N_4495,In_2854,In_262);
nand U4496 (N_4496,In_4793,In_221);
xor U4497 (N_4497,In_1009,In_3388);
or U4498 (N_4498,In_226,In_4041);
nand U4499 (N_4499,In_685,In_4507);
nor U4500 (N_4500,In_433,In_2308);
nand U4501 (N_4501,In_3396,In_425);
or U4502 (N_4502,In_4489,In_2152);
and U4503 (N_4503,In_2939,In_4815);
nand U4504 (N_4504,In_3881,In_1750);
xor U4505 (N_4505,In_1476,In_3645);
and U4506 (N_4506,In_3604,In_794);
or U4507 (N_4507,In_439,In_1118);
nor U4508 (N_4508,In_3739,In_1676);
and U4509 (N_4509,In_905,In_4108);
nor U4510 (N_4510,In_3714,In_637);
xnor U4511 (N_4511,In_4963,In_2384);
nor U4512 (N_4512,In_2022,In_1447);
nand U4513 (N_4513,In_2865,In_1199);
and U4514 (N_4514,In_1485,In_2363);
or U4515 (N_4515,In_476,In_3221);
or U4516 (N_4516,In_76,In_3812);
nor U4517 (N_4517,In_4888,In_179);
or U4518 (N_4518,In_2579,In_2943);
nand U4519 (N_4519,In_799,In_1767);
and U4520 (N_4520,In_1400,In_3750);
xnor U4521 (N_4521,In_3868,In_1848);
xnor U4522 (N_4522,In_3373,In_715);
nand U4523 (N_4523,In_4640,In_1839);
nor U4524 (N_4524,In_2339,In_2533);
or U4525 (N_4525,In_583,In_2018);
xor U4526 (N_4526,In_3802,In_1894);
xor U4527 (N_4527,In_4915,In_1509);
nand U4528 (N_4528,In_4800,In_2002);
and U4529 (N_4529,In_915,In_2432);
and U4530 (N_4530,In_1408,In_3636);
nand U4531 (N_4531,In_4760,In_39);
xnor U4532 (N_4532,In_4876,In_1755);
xor U4533 (N_4533,In_1984,In_3904);
nor U4534 (N_4534,In_4869,In_4803);
and U4535 (N_4535,In_748,In_3327);
xor U4536 (N_4536,In_4827,In_1894);
nand U4537 (N_4537,In_844,In_956);
and U4538 (N_4538,In_3557,In_3617);
or U4539 (N_4539,In_884,In_305);
nor U4540 (N_4540,In_3009,In_2221);
nand U4541 (N_4541,In_3082,In_640);
and U4542 (N_4542,In_2770,In_748);
nand U4543 (N_4543,In_4028,In_1631);
and U4544 (N_4544,In_299,In_342);
nand U4545 (N_4545,In_3048,In_4614);
and U4546 (N_4546,In_4185,In_2423);
xor U4547 (N_4547,In_3167,In_4016);
and U4548 (N_4548,In_756,In_2599);
nor U4549 (N_4549,In_3544,In_3765);
nor U4550 (N_4550,In_1104,In_3538);
or U4551 (N_4551,In_4315,In_451);
or U4552 (N_4552,In_4996,In_2814);
or U4553 (N_4553,In_807,In_285);
and U4554 (N_4554,In_2175,In_1171);
or U4555 (N_4555,In_2749,In_4935);
xnor U4556 (N_4556,In_1992,In_416);
nand U4557 (N_4557,In_98,In_3081);
xnor U4558 (N_4558,In_869,In_816);
or U4559 (N_4559,In_902,In_2551);
xnor U4560 (N_4560,In_2219,In_458);
nor U4561 (N_4561,In_3899,In_625);
nor U4562 (N_4562,In_1953,In_216);
xor U4563 (N_4563,In_1643,In_1180);
and U4564 (N_4564,In_3040,In_237);
xnor U4565 (N_4565,In_3382,In_247);
nand U4566 (N_4566,In_2102,In_2785);
nor U4567 (N_4567,In_3276,In_383);
or U4568 (N_4568,In_2801,In_3748);
nor U4569 (N_4569,In_2719,In_2272);
nand U4570 (N_4570,In_4107,In_731);
and U4571 (N_4571,In_2058,In_4321);
or U4572 (N_4572,In_3781,In_2391);
and U4573 (N_4573,In_4873,In_4514);
and U4574 (N_4574,In_2730,In_3596);
nor U4575 (N_4575,In_4832,In_4734);
nor U4576 (N_4576,In_4566,In_4990);
or U4577 (N_4577,In_3231,In_3263);
xor U4578 (N_4578,In_3380,In_3396);
or U4579 (N_4579,In_2190,In_2546);
xor U4580 (N_4580,In_1879,In_3241);
and U4581 (N_4581,In_3485,In_368);
or U4582 (N_4582,In_1562,In_2762);
nand U4583 (N_4583,In_4760,In_2996);
and U4584 (N_4584,In_147,In_4296);
nand U4585 (N_4585,In_1644,In_4366);
nor U4586 (N_4586,In_1319,In_4421);
and U4587 (N_4587,In_3460,In_2518);
nor U4588 (N_4588,In_425,In_4984);
xor U4589 (N_4589,In_8,In_4401);
or U4590 (N_4590,In_3390,In_1559);
nand U4591 (N_4591,In_959,In_1076);
or U4592 (N_4592,In_132,In_421);
or U4593 (N_4593,In_895,In_2981);
nor U4594 (N_4594,In_1268,In_1776);
xnor U4595 (N_4595,In_2337,In_1471);
nor U4596 (N_4596,In_2623,In_1770);
nor U4597 (N_4597,In_1436,In_1289);
nand U4598 (N_4598,In_3777,In_4346);
nand U4599 (N_4599,In_970,In_2252);
nor U4600 (N_4600,In_2387,In_4696);
and U4601 (N_4601,In_2176,In_4889);
or U4602 (N_4602,In_3132,In_1626);
nor U4603 (N_4603,In_1812,In_2107);
xnor U4604 (N_4604,In_2036,In_595);
nand U4605 (N_4605,In_935,In_3004);
nand U4606 (N_4606,In_267,In_2697);
xor U4607 (N_4607,In_3606,In_4393);
and U4608 (N_4608,In_4646,In_3720);
xnor U4609 (N_4609,In_1445,In_4335);
xor U4610 (N_4610,In_2529,In_1188);
nand U4611 (N_4611,In_2006,In_1306);
or U4612 (N_4612,In_1784,In_3876);
nand U4613 (N_4613,In_2267,In_4377);
xnor U4614 (N_4614,In_624,In_1717);
or U4615 (N_4615,In_2931,In_43);
xnor U4616 (N_4616,In_899,In_774);
and U4617 (N_4617,In_1726,In_1600);
xor U4618 (N_4618,In_1841,In_4733);
xnor U4619 (N_4619,In_883,In_22);
or U4620 (N_4620,In_2228,In_3947);
or U4621 (N_4621,In_2208,In_2657);
or U4622 (N_4622,In_3909,In_2629);
and U4623 (N_4623,In_2345,In_2558);
nand U4624 (N_4624,In_318,In_4152);
or U4625 (N_4625,In_1858,In_4842);
xor U4626 (N_4626,In_2120,In_2748);
or U4627 (N_4627,In_4357,In_1758);
and U4628 (N_4628,In_1374,In_1055);
xor U4629 (N_4629,In_26,In_1123);
nand U4630 (N_4630,In_527,In_2283);
and U4631 (N_4631,In_4768,In_1777);
nor U4632 (N_4632,In_4046,In_3341);
and U4633 (N_4633,In_4477,In_1020);
and U4634 (N_4634,In_857,In_1411);
nand U4635 (N_4635,In_2237,In_3607);
nand U4636 (N_4636,In_1286,In_3495);
nand U4637 (N_4637,In_2400,In_2254);
nand U4638 (N_4638,In_1514,In_1350);
xor U4639 (N_4639,In_2623,In_1104);
and U4640 (N_4640,In_3143,In_1733);
or U4641 (N_4641,In_3607,In_4118);
nand U4642 (N_4642,In_1999,In_4353);
and U4643 (N_4643,In_3727,In_4486);
or U4644 (N_4644,In_3327,In_4831);
xnor U4645 (N_4645,In_2382,In_409);
nor U4646 (N_4646,In_1154,In_2802);
nor U4647 (N_4647,In_3413,In_663);
or U4648 (N_4648,In_1588,In_1322);
or U4649 (N_4649,In_264,In_2175);
nand U4650 (N_4650,In_1731,In_3255);
and U4651 (N_4651,In_1116,In_4351);
nor U4652 (N_4652,In_3949,In_2034);
and U4653 (N_4653,In_551,In_190);
xnor U4654 (N_4654,In_1357,In_4558);
xnor U4655 (N_4655,In_4306,In_626);
nand U4656 (N_4656,In_3375,In_3423);
and U4657 (N_4657,In_4441,In_906);
nand U4658 (N_4658,In_1157,In_1964);
nand U4659 (N_4659,In_216,In_422);
nand U4660 (N_4660,In_1353,In_871);
or U4661 (N_4661,In_4667,In_1877);
nand U4662 (N_4662,In_4578,In_3581);
nand U4663 (N_4663,In_526,In_4093);
xnor U4664 (N_4664,In_960,In_2993);
and U4665 (N_4665,In_2552,In_3277);
or U4666 (N_4666,In_1233,In_301);
and U4667 (N_4667,In_1830,In_3656);
xor U4668 (N_4668,In_2998,In_372);
nand U4669 (N_4669,In_2056,In_2221);
and U4670 (N_4670,In_2171,In_628);
nor U4671 (N_4671,In_418,In_1738);
nor U4672 (N_4672,In_2143,In_314);
nor U4673 (N_4673,In_2929,In_1810);
or U4674 (N_4674,In_4540,In_3056);
nor U4675 (N_4675,In_1164,In_4785);
nor U4676 (N_4676,In_70,In_2962);
or U4677 (N_4677,In_647,In_101);
nand U4678 (N_4678,In_2065,In_389);
and U4679 (N_4679,In_1871,In_3520);
and U4680 (N_4680,In_3322,In_825);
or U4681 (N_4681,In_3693,In_2070);
nand U4682 (N_4682,In_2104,In_861);
and U4683 (N_4683,In_1499,In_1904);
and U4684 (N_4684,In_4360,In_863);
nor U4685 (N_4685,In_1292,In_114);
nor U4686 (N_4686,In_3465,In_3245);
or U4687 (N_4687,In_2038,In_1621);
nor U4688 (N_4688,In_2094,In_2851);
and U4689 (N_4689,In_1007,In_280);
or U4690 (N_4690,In_4818,In_3756);
and U4691 (N_4691,In_1689,In_3347);
nor U4692 (N_4692,In_4142,In_2037);
nor U4693 (N_4693,In_1632,In_2366);
nand U4694 (N_4694,In_3793,In_1381);
nand U4695 (N_4695,In_4868,In_3169);
or U4696 (N_4696,In_1817,In_4598);
or U4697 (N_4697,In_2564,In_1359);
or U4698 (N_4698,In_1333,In_647);
xnor U4699 (N_4699,In_1779,In_4071);
nor U4700 (N_4700,In_4315,In_743);
or U4701 (N_4701,In_2634,In_2814);
xnor U4702 (N_4702,In_677,In_4119);
or U4703 (N_4703,In_3252,In_1206);
or U4704 (N_4704,In_221,In_1038);
nand U4705 (N_4705,In_1191,In_257);
and U4706 (N_4706,In_2572,In_2739);
nor U4707 (N_4707,In_1623,In_661);
nor U4708 (N_4708,In_3561,In_4230);
and U4709 (N_4709,In_4019,In_3162);
nand U4710 (N_4710,In_4274,In_888);
nand U4711 (N_4711,In_2114,In_3372);
xor U4712 (N_4712,In_2461,In_3611);
and U4713 (N_4713,In_3816,In_4263);
nand U4714 (N_4714,In_2327,In_542);
nor U4715 (N_4715,In_1997,In_338);
nand U4716 (N_4716,In_3190,In_732);
and U4717 (N_4717,In_980,In_1818);
or U4718 (N_4718,In_1727,In_769);
and U4719 (N_4719,In_713,In_4612);
or U4720 (N_4720,In_3544,In_458);
nor U4721 (N_4721,In_1154,In_4931);
nor U4722 (N_4722,In_3080,In_2485);
nor U4723 (N_4723,In_2168,In_1510);
and U4724 (N_4724,In_2856,In_4286);
nand U4725 (N_4725,In_2387,In_4197);
nand U4726 (N_4726,In_1770,In_239);
nor U4727 (N_4727,In_3886,In_2669);
or U4728 (N_4728,In_232,In_3018);
nor U4729 (N_4729,In_4931,In_2147);
nor U4730 (N_4730,In_134,In_664);
and U4731 (N_4731,In_3537,In_3960);
or U4732 (N_4732,In_4493,In_529);
nor U4733 (N_4733,In_3447,In_4108);
nor U4734 (N_4734,In_280,In_4205);
nor U4735 (N_4735,In_4145,In_2175);
xor U4736 (N_4736,In_751,In_1337);
or U4737 (N_4737,In_3603,In_639);
or U4738 (N_4738,In_1752,In_4490);
nand U4739 (N_4739,In_4541,In_2150);
nor U4740 (N_4740,In_3375,In_693);
or U4741 (N_4741,In_1362,In_924);
nand U4742 (N_4742,In_2252,In_142);
nand U4743 (N_4743,In_2918,In_1957);
xor U4744 (N_4744,In_1424,In_4930);
xnor U4745 (N_4745,In_1148,In_1322);
or U4746 (N_4746,In_4070,In_4562);
nand U4747 (N_4747,In_530,In_659);
nor U4748 (N_4748,In_381,In_2534);
and U4749 (N_4749,In_4780,In_1125);
nor U4750 (N_4750,In_4943,In_1845);
xnor U4751 (N_4751,In_230,In_2739);
xnor U4752 (N_4752,In_4080,In_1091);
xor U4753 (N_4753,In_2973,In_2437);
nand U4754 (N_4754,In_2370,In_2430);
xnor U4755 (N_4755,In_309,In_3271);
nand U4756 (N_4756,In_1692,In_52);
xor U4757 (N_4757,In_4955,In_3698);
nand U4758 (N_4758,In_4681,In_1491);
nand U4759 (N_4759,In_4038,In_3616);
nand U4760 (N_4760,In_1031,In_3352);
and U4761 (N_4761,In_4762,In_1896);
xnor U4762 (N_4762,In_2919,In_4315);
or U4763 (N_4763,In_1779,In_620);
nor U4764 (N_4764,In_4847,In_2074);
and U4765 (N_4765,In_2184,In_255);
or U4766 (N_4766,In_3626,In_3606);
and U4767 (N_4767,In_1427,In_2801);
and U4768 (N_4768,In_1151,In_4574);
and U4769 (N_4769,In_3862,In_4278);
or U4770 (N_4770,In_4277,In_4333);
or U4771 (N_4771,In_1874,In_1698);
and U4772 (N_4772,In_1470,In_4774);
or U4773 (N_4773,In_1495,In_253);
nand U4774 (N_4774,In_2693,In_3546);
nand U4775 (N_4775,In_924,In_493);
or U4776 (N_4776,In_705,In_4148);
and U4777 (N_4777,In_2800,In_1121);
xor U4778 (N_4778,In_2312,In_2654);
xor U4779 (N_4779,In_491,In_421);
nand U4780 (N_4780,In_2807,In_280);
or U4781 (N_4781,In_1963,In_3500);
nor U4782 (N_4782,In_4822,In_3471);
xnor U4783 (N_4783,In_403,In_502);
nor U4784 (N_4784,In_3798,In_94);
and U4785 (N_4785,In_3451,In_2781);
nor U4786 (N_4786,In_2244,In_4079);
nor U4787 (N_4787,In_3329,In_4614);
or U4788 (N_4788,In_4129,In_502);
or U4789 (N_4789,In_1557,In_4040);
nor U4790 (N_4790,In_734,In_1847);
or U4791 (N_4791,In_168,In_708);
xor U4792 (N_4792,In_3924,In_3353);
nor U4793 (N_4793,In_1829,In_739);
nor U4794 (N_4794,In_1330,In_1829);
or U4795 (N_4795,In_1097,In_1967);
xnor U4796 (N_4796,In_2512,In_2437);
nor U4797 (N_4797,In_48,In_4313);
or U4798 (N_4798,In_4555,In_4634);
nor U4799 (N_4799,In_3090,In_1310);
and U4800 (N_4800,In_3704,In_1857);
nor U4801 (N_4801,In_862,In_4109);
nand U4802 (N_4802,In_4074,In_4421);
nand U4803 (N_4803,In_4692,In_4827);
or U4804 (N_4804,In_3343,In_1779);
xor U4805 (N_4805,In_2902,In_2914);
xor U4806 (N_4806,In_219,In_2470);
or U4807 (N_4807,In_1797,In_3326);
or U4808 (N_4808,In_3470,In_1222);
nand U4809 (N_4809,In_2514,In_3298);
or U4810 (N_4810,In_940,In_396);
and U4811 (N_4811,In_3145,In_2393);
xor U4812 (N_4812,In_3035,In_2211);
nand U4813 (N_4813,In_1780,In_3670);
nor U4814 (N_4814,In_3067,In_3638);
or U4815 (N_4815,In_204,In_4648);
or U4816 (N_4816,In_2672,In_2663);
or U4817 (N_4817,In_2102,In_3595);
nand U4818 (N_4818,In_335,In_3023);
and U4819 (N_4819,In_805,In_4584);
and U4820 (N_4820,In_1221,In_2016);
nand U4821 (N_4821,In_3071,In_3068);
xnor U4822 (N_4822,In_4843,In_1011);
nor U4823 (N_4823,In_1761,In_2575);
and U4824 (N_4824,In_1223,In_2979);
nor U4825 (N_4825,In_2773,In_4158);
and U4826 (N_4826,In_3581,In_4628);
or U4827 (N_4827,In_3286,In_1212);
xnor U4828 (N_4828,In_3735,In_673);
and U4829 (N_4829,In_4889,In_2806);
or U4830 (N_4830,In_2999,In_4778);
nand U4831 (N_4831,In_2409,In_4415);
and U4832 (N_4832,In_2917,In_168);
nor U4833 (N_4833,In_199,In_1308);
and U4834 (N_4834,In_4040,In_3204);
nand U4835 (N_4835,In_4825,In_4142);
or U4836 (N_4836,In_479,In_843);
xor U4837 (N_4837,In_2413,In_3953);
nand U4838 (N_4838,In_3319,In_3149);
nor U4839 (N_4839,In_65,In_1246);
nor U4840 (N_4840,In_2660,In_2646);
or U4841 (N_4841,In_1929,In_328);
or U4842 (N_4842,In_3895,In_1976);
or U4843 (N_4843,In_3892,In_465);
or U4844 (N_4844,In_926,In_3122);
or U4845 (N_4845,In_176,In_2789);
or U4846 (N_4846,In_2689,In_1194);
and U4847 (N_4847,In_2957,In_2116);
or U4848 (N_4848,In_2646,In_117);
nand U4849 (N_4849,In_4441,In_1871);
nand U4850 (N_4850,In_1646,In_3915);
and U4851 (N_4851,In_3113,In_944);
nand U4852 (N_4852,In_4689,In_3045);
xnor U4853 (N_4853,In_3344,In_633);
nand U4854 (N_4854,In_4650,In_3258);
and U4855 (N_4855,In_4930,In_2135);
or U4856 (N_4856,In_124,In_4893);
and U4857 (N_4857,In_3621,In_4646);
and U4858 (N_4858,In_1696,In_799);
or U4859 (N_4859,In_4013,In_2285);
nand U4860 (N_4860,In_4709,In_1192);
and U4861 (N_4861,In_2898,In_1958);
nand U4862 (N_4862,In_2184,In_2816);
or U4863 (N_4863,In_1957,In_3644);
nand U4864 (N_4864,In_2488,In_511);
or U4865 (N_4865,In_4060,In_4894);
nor U4866 (N_4866,In_1166,In_4614);
nand U4867 (N_4867,In_3732,In_4975);
nor U4868 (N_4868,In_2309,In_4309);
or U4869 (N_4869,In_1577,In_688);
or U4870 (N_4870,In_3837,In_4266);
nand U4871 (N_4871,In_2276,In_3963);
or U4872 (N_4872,In_616,In_706);
and U4873 (N_4873,In_2243,In_3586);
and U4874 (N_4874,In_4567,In_2073);
and U4875 (N_4875,In_4043,In_3361);
xnor U4876 (N_4876,In_2581,In_2442);
nor U4877 (N_4877,In_4724,In_4716);
or U4878 (N_4878,In_3918,In_387);
xnor U4879 (N_4879,In_3676,In_442);
or U4880 (N_4880,In_1179,In_3206);
and U4881 (N_4881,In_4157,In_2425);
nand U4882 (N_4882,In_829,In_3120);
and U4883 (N_4883,In_3729,In_1642);
nor U4884 (N_4884,In_2280,In_4934);
or U4885 (N_4885,In_871,In_3795);
and U4886 (N_4886,In_2734,In_4750);
nand U4887 (N_4887,In_4984,In_913);
or U4888 (N_4888,In_68,In_4762);
and U4889 (N_4889,In_4762,In_4446);
or U4890 (N_4890,In_3138,In_3301);
nand U4891 (N_4891,In_2351,In_3472);
and U4892 (N_4892,In_1509,In_3942);
xnor U4893 (N_4893,In_2967,In_4217);
and U4894 (N_4894,In_3109,In_3644);
nand U4895 (N_4895,In_3352,In_674);
nor U4896 (N_4896,In_4481,In_2758);
nor U4897 (N_4897,In_3566,In_1346);
and U4898 (N_4898,In_2071,In_4070);
and U4899 (N_4899,In_2591,In_1533);
nor U4900 (N_4900,In_2317,In_3376);
and U4901 (N_4901,In_80,In_1020);
xor U4902 (N_4902,In_4722,In_3575);
xnor U4903 (N_4903,In_4581,In_4484);
and U4904 (N_4904,In_1385,In_4403);
or U4905 (N_4905,In_1208,In_585);
and U4906 (N_4906,In_29,In_707);
xnor U4907 (N_4907,In_3953,In_4906);
xnor U4908 (N_4908,In_4410,In_2568);
xnor U4909 (N_4909,In_3375,In_4601);
and U4910 (N_4910,In_1448,In_455);
xor U4911 (N_4911,In_1697,In_4052);
nand U4912 (N_4912,In_1983,In_1889);
or U4913 (N_4913,In_3610,In_879);
or U4914 (N_4914,In_1103,In_3464);
or U4915 (N_4915,In_731,In_247);
xnor U4916 (N_4916,In_2209,In_2718);
xnor U4917 (N_4917,In_349,In_760);
or U4918 (N_4918,In_2573,In_1323);
xor U4919 (N_4919,In_1031,In_4568);
or U4920 (N_4920,In_4442,In_4983);
xor U4921 (N_4921,In_4331,In_474);
nand U4922 (N_4922,In_2378,In_4512);
nand U4923 (N_4923,In_4526,In_4246);
xor U4924 (N_4924,In_3660,In_269);
or U4925 (N_4925,In_4007,In_314);
and U4926 (N_4926,In_3340,In_4175);
xnor U4927 (N_4927,In_3008,In_2317);
and U4928 (N_4928,In_4838,In_2764);
nand U4929 (N_4929,In_2587,In_702);
nor U4930 (N_4930,In_3645,In_4293);
xor U4931 (N_4931,In_4047,In_1947);
or U4932 (N_4932,In_1573,In_1932);
or U4933 (N_4933,In_374,In_2209);
nand U4934 (N_4934,In_2677,In_1389);
or U4935 (N_4935,In_1412,In_3330);
or U4936 (N_4936,In_4624,In_1371);
nand U4937 (N_4937,In_2758,In_2805);
nor U4938 (N_4938,In_1876,In_4509);
xnor U4939 (N_4939,In_3185,In_4688);
nor U4940 (N_4940,In_1913,In_601);
nand U4941 (N_4941,In_459,In_737);
nand U4942 (N_4942,In_2335,In_4815);
or U4943 (N_4943,In_2467,In_276);
nand U4944 (N_4944,In_2621,In_4886);
nand U4945 (N_4945,In_3360,In_2406);
nor U4946 (N_4946,In_4680,In_720);
or U4947 (N_4947,In_1613,In_3468);
xor U4948 (N_4948,In_1685,In_1455);
and U4949 (N_4949,In_4534,In_4314);
nand U4950 (N_4950,In_1563,In_2033);
or U4951 (N_4951,In_2263,In_3131);
or U4952 (N_4952,In_1866,In_3516);
nor U4953 (N_4953,In_2932,In_1529);
nand U4954 (N_4954,In_667,In_2828);
and U4955 (N_4955,In_4393,In_3910);
nand U4956 (N_4956,In_2218,In_1504);
or U4957 (N_4957,In_2102,In_4315);
and U4958 (N_4958,In_3213,In_1664);
nand U4959 (N_4959,In_2141,In_1158);
or U4960 (N_4960,In_2268,In_1786);
nand U4961 (N_4961,In_76,In_1147);
xnor U4962 (N_4962,In_3670,In_2081);
nor U4963 (N_4963,In_1291,In_3905);
and U4964 (N_4964,In_1720,In_3699);
nand U4965 (N_4965,In_3247,In_2238);
nand U4966 (N_4966,In_2312,In_2491);
nor U4967 (N_4967,In_2423,In_4616);
or U4968 (N_4968,In_3545,In_559);
and U4969 (N_4969,In_4363,In_708);
and U4970 (N_4970,In_4476,In_2430);
xnor U4971 (N_4971,In_3516,In_627);
or U4972 (N_4972,In_1299,In_3161);
xnor U4973 (N_4973,In_638,In_1208);
nor U4974 (N_4974,In_2833,In_1672);
nand U4975 (N_4975,In_2642,In_163);
or U4976 (N_4976,In_1301,In_4773);
nand U4977 (N_4977,In_868,In_4246);
nand U4978 (N_4978,In_3971,In_3011);
or U4979 (N_4979,In_2300,In_2454);
and U4980 (N_4980,In_1644,In_3759);
xor U4981 (N_4981,In_4196,In_983);
and U4982 (N_4982,In_980,In_3369);
nor U4983 (N_4983,In_489,In_4585);
xor U4984 (N_4984,In_3855,In_2033);
and U4985 (N_4985,In_2043,In_4457);
xnor U4986 (N_4986,In_2727,In_1505);
and U4987 (N_4987,In_2924,In_1279);
and U4988 (N_4988,In_4191,In_4967);
nor U4989 (N_4989,In_2380,In_301);
or U4990 (N_4990,In_4350,In_298);
nor U4991 (N_4991,In_2630,In_2343);
nand U4992 (N_4992,In_4356,In_2349);
and U4993 (N_4993,In_533,In_915);
xor U4994 (N_4994,In_3512,In_4864);
nor U4995 (N_4995,In_435,In_3850);
nand U4996 (N_4996,In_1290,In_456);
nand U4997 (N_4997,In_115,In_3948);
or U4998 (N_4998,In_1518,In_2836);
nand U4999 (N_4999,In_1293,In_4992);
or U5000 (N_5000,In_85,In_1482);
or U5001 (N_5001,In_566,In_4853);
or U5002 (N_5002,In_3011,In_3243);
or U5003 (N_5003,In_70,In_3822);
xnor U5004 (N_5004,In_710,In_4029);
xor U5005 (N_5005,In_1591,In_2291);
nand U5006 (N_5006,In_3628,In_1798);
or U5007 (N_5007,In_4987,In_3599);
or U5008 (N_5008,In_3022,In_3217);
or U5009 (N_5009,In_1208,In_523);
nand U5010 (N_5010,In_257,In_3835);
or U5011 (N_5011,In_4964,In_1523);
nor U5012 (N_5012,In_2644,In_862);
xor U5013 (N_5013,In_49,In_249);
and U5014 (N_5014,In_3491,In_432);
nand U5015 (N_5015,In_2475,In_30);
and U5016 (N_5016,In_1919,In_1810);
nor U5017 (N_5017,In_412,In_1043);
or U5018 (N_5018,In_858,In_2764);
nand U5019 (N_5019,In_56,In_4466);
nand U5020 (N_5020,In_642,In_3546);
and U5021 (N_5021,In_603,In_302);
nor U5022 (N_5022,In_2323,In_1735);
xor U5023 (N_5023,In_424,In_109);
and U5024 (N_5024,In_926,In_3658);
nor U5025 (N_5025,In_2779,In_2463);
nand U5026 (N_5026,In_322,In_2407);
nor U5027 (N_5027,In_3259,In_4960);
or U5028 (N_5028,In_2461,In_2957);
nand U5029 (N_5029,In_666,In_472);
nand U5030 (N_5030,In_810,In_496);
nor U5031 (N_5031,In_4804,In_140);
nand U5032 (N_5032,In_4896,In_4413);
or U5033 (N_5033,In_4872,In_3123);
nand U5034 (N_5034,In_1940,In_2710);
nor U5035 (N_5035,In_3472,In_1357);
xor U5036 (N_5036,In_2017,In_3960);
nand U5037 (N_5037,In_1334,In_3229);
or U5038 (N_5038,In_1464,In_370);
nor U5039 (N_5039,In_1068,In_1532);
or U5040 (N_5040,In_4649,In_990);
and U5041 (N_5041,In_3000,In_3376);
nand U5042 (N_5042,In_4247,In_4342);
nand U5043 (N_5043,In_1610,In_2617);
xor U5044 (N_5044,In_2154,In_1516);
nor U5045 (N_5045,In_973,In_1759);
or U5046 (N_5046,In_4754,In_658);
nand U5047 (N_5047,In_1806,In_2718);
nor U5048 (N_5048,In_415,In_3983);
and U5049 (N_5049,In_1301,In_3149);
nor U5050 (N_5050,In_1847,In_4376);
nor U5051 (N_5051,In_1782,In_62);
or U5052 (N_5052,In_2366,In_790);
nand U5053 (N_5053,In_3661,In_3335);
xor U5054 (N_5054,In_4345,In_1437);
and U5055 (N_5055,In_4934,In_507);
xnor U5056 (N_5056,In_1010,In_1154);
and U5057 (N_5057,In_3176,In_4329);
nand U5058 (N_5058,In_459,In_578);
and U5059 (N_5059,In_4199,In_2096);
xor U5060 (N_5060,In_3051,In_3678);
or U5061 (N_5061,In_1085,In_2435);
xor U5062 (N_5062,In_92,In_1417);
nor U5063 (N_5063,In_438,In_571);
xnor U5064 (N_5064,In_3829,In_2546);
xor U5065 (N_5065,In_4692,In_2990);
nor U5066 (N_5066,In_2534,In_3985);
nor U5067 (N_5067,In_2843,In_490);
xnor U5068 (N_5068,In_19,In_3802);
nor U5069 (N_5069,In_1874,In_438);
xor U5070 (N_5070,In_3523,In_2420);
nand U5071 (N_5071,In_1748,In_4026);
xor U5072 (N_5072,In_684,In_4110);
or U5073 (N_5073,In_900,In_693);
nor U5074 (N_5074,In_2566,In_4166);
nand U5075 (N_5075,In_1680,In_4506);
nand U5076 (N_5076,In_4705,In_2742);
nand U5077 (N_5077,In_2792,In_3142);
xor U5078 (N_5078,In_3864,In_504);
xnor U5079 (N_5079,In_4347,In_3438);
xnor U5080 (N_5080,In_3679,In_3552);
or U5081 (N_5081,In_38,In_2510);
nor U5082 (N_5082,In_3900,In_1704);
nand U5083 (N_5083,In_3246,In_58);
nor U5084 (N_5084,In_2124,In_1089);
nand U5085 (N_5085,In_1957,In_469);
xor U5086 (N_5086,In_3490,In_1258);
nor U5087 (N_5087,In_4003,In_4183);
or U5088 (N_5088,In_282,In_690);
and U5089 (N_5089,In_2508,In_2229);
and U5090 (N_5090,In_107,In_1372);
and U5091 (N_5091,In_724,In_411);
and U5092 (N_5092,In_1796,In_1221);
nand U5093 (N_5093,In_244,In_4944);
xor U5094 (N_5094,In_16,In_3682);
and U5095 (N_5095,In_3655,In_3833);
nand U5096 (N_5096,In_1080,In_635);
xnor U5097 (N_5097,In_1332,In_4878);
or U5098 (N_5098,In_223,In_3219);
xnor U5099 (N_5099,In_4683,In_618);
nor U5100 (N_5100,In_3893,In_1241);
xor U5101 (N_5101,In_4173,In_4909);
nand U5102 (N_5102,In_4959,In_4775);
or U5103 (N_5103,In_1268,In_4023);
xor U5104 (N_5104,In_529,In_3979);
xor U5105 (N_5105,In_4108,In_321);
or U5106 (N_5106,In_4682,In_1706);
and U5107 (N_5107,In_1873,In_2297);
nand U5108 (N_5108,In_3377,In_3948);
and U5109 (N_5109,In_2568,In_1564);
nor U5110 (N_5110,In_2943,In_4563);
nand U5111 (N_5111,In_4988,In_3334);
nand U5112 (N_5112,In_1069,In_1746);
xnor U5113 (N_5113,In_1617,In_2693);
or U5114 (N_5114,In_876,In_1040);
or U5115 (N_5115,In_635,In_664);
nand U5116 (N_5116,In_3798,In_2211);
or U5117 (N_5117,In_866,In_4012);
xnor U5118 (N_5118,In_4845,In_1703);
and U5119 (N_5119,In_2095,In_1209);
xnor U5120 (N_5120,In_3984,In_958);
xor U5121 (N_5121,In_1297,In_2776);
xnor U5122 (N_5122,In_3597,In_3687);
nand U5123 (N_5123,In_2020,In_726);
or U5124 (N_5124,In_183,In_1004);
and U5125 (N_5125,In_2815,In_4610);
and U5126 (N_5126,In_2236,In_2561);
and U5127 (N_5127,In_1466,In_3900);
xnor U5128 (N_5128,In_3460,In_2803);
xor U5129 (N_5129,In_4405,In_2804);
nor U5130 (N_5130,In_2281,In_4131);
nor U5131 (N_5131,In_1564,In_46);
or U5132 (N_5132,In_3188,In_2322);
or U5133 (N_5133,In_3752,In_874);
nor U5134 (N_5134,In_616,In_537);
nand U5135 (N_5135,In_3264,In_2598);
nor U5136 (N_5136,In_4436,In_923);
or U5137 (N_5137,In_3409,In_3230);
xor U5138 (N_5138,In_1573,In_2661);
xor U5139 (N_5139,In_3656,In_2621);
nand U5140 (N_5140,In_1430,In_50);
nand U5141 (N_5141,In_3346,In_1184);
xnor U5142 (N_5142,In_3276,In_3187);
nor U5143 (N_5143,In_1171,In_4625);
or U5144 (N_5144,In_1821,In_4078);
and U5145 (N_5145,In_4847,In_4991);
or U5146 (N_5146,In_4871,In_2115);
nand U5147 (N_5147,In_2181,In_3965);
nand U5148 (N_5148,In_1955,In_4221);
nand U5149 (N_5149,In_2181,In_40);
and U5150 (N_5150,In_1343,In_1999);
nand U5151 (N_5151,In_4862,In_2737);
xnor U5152 (N_5152,In_1480,In_2353);
or U5153 (N_5153,In_1454,In_857);
or U5154 (N_5154,In_226,In_697);
nand U5155 (N_5155,In_2491,In_1829);
xor U5156 (N_5156,In_861,In_3286);
or U5157 (N_5157,In_2313,In_541);
or U5158 (N_5158,In_1685,In_2697);
xor U5159 (N_5159,In_4658,In_1795);
and U5160 (N_5160,In_1773,In_3786);
nand U5161 (N_5161,In_4750,In_4145);
xor U5162 (N_5162,In_4845,In_2816);
xor U5163 (N_5163,In_1209,In_1564);
nand U5164 (N_5164,In_3783,In_2346);
xnor U5165 (N_5165,In_402,In_2685);
nor U5166 (N_5166,In_2816,In_995);
xnor U5167 (N_5167,In_3272,In_4112);
nor U5168 (N_5168,In_4851,In_1871);
and U5169 (N_5169,In_3231,In_4911);
xor U5170 (N_5170,In_2265,In_2942);
and U5171 (N_5171,In_1072,In_3558);
xnor U5172 (N_5172,In_1172,In_1368);
nor U5173 (N_5173,In_2444,In_1348);
and U5174 (N_5174,In_403,In_2608);
xor U5175 (N_5175,In_259,In_2539);
or U5176 (N_5176,In_3377,In_1757);
and U5177 (N_5177,In_4379,In_2032);
xnor U5178 (N_5178,In_4022,In_3943);
xor U5179 (N_5179,In_2725,In_4709);
nand U5180 (N_5180,In_2303,In_3714);
or U5181 (N_5181,In_1375,In_3767);
or U5182 (N_5182,In_378,In_3275);
nor U5183 (N_5183,In_2340,In_1060);
xor U5184 (N_5184,In_345,In_4385);
nand U5185 (N_5185,In_3617,In_3488);
nand U5186 (N_5186,In_4441,In_35);
and U5187 (N_5187,In_1846,In_507);
and U5188 (N_5188,In_248,In_3503);
xor U5189 (N_5189,In_3801,In_3784);
and U5190 (N_5190,In_4782,In_1664);
and U5191 (N_5191,In_75,In_2570);
or U5192 (N_5192,In_2905,In_2885);
xor U5193 (N_5193,In_653,In_275);
nor U5194 (N_5194,In_2738,In_1414);
xor U5195 (N_5195,In_767,In_1025);
xor U5196 (N_5196,In_504,In_2003);
nand U5197 (N_5197,In_557,In_456);
xnor U5198 (N_5198,In_4358,In_2083);
nor U5199 (N_5199,In_3615,In_2011);
and U5200 (N_5200,In_1418,In_1106);
and U5201 (N_5201,In_1832,In_2471);
xor U5202 (N_5202,In_4608,In_4844);
nor U5203 (N_5203,In_4193,In_2925);
nor U5204 (N_5204,In_4632,In_513);
and U5205 (N_5205,In_4203,In_3722);
and U5206 (N_5206,In_374,In_1528);
nand U5207 (N_5207,In_4577,In_4266);
xor U5208 (N_5208,In_373,In_239);
or U5209 (N_5209,In_1692,In_3038);
nor U5210 (N_5210,In_4831,In_2904);
or U5211 (N_5211,In_571,In_548);
or U5212 (N_5212,In_4087,In_876);
xor U5213 (N_5213,In_1225,In_3157);
nand U5214 (N_5214,In_1984,In_4540);
or U5215 (N_5215,In_4051,In_1766);
xnor U5216 (N_5216,In_3116,In_3963);
nand U5217 (N_5217,In_3299,In_2142);
nand U5218 (N_5218,In_608,In_2277);
xor U5219 (N_5219,In_3762,In_4631);
xnor U5220 (N_5220,In_4142,In_4799);
nor U5221 (N_5221,In_2674,In_1676);
and U5222 (N_5222,In_2053,In_2608);
nand U5223 (N_5223,In_4016,In_4205);
and U5224 (N_5224,In_2639,In_4067);
nand U5225 (N_5225,In_151,In_720);
nand U5226 (N_5226,In_2564,In_3572);
xnor U5227 (N_5227,In_3308,In_4224);
xor U5228 (N_5228,In_580,In_3993);
xor U5229 (N_5229,In_753,In_2493);
and U5230 (N_5230,In_460,In_3984);
nand U5231 (N_5231,In_1581,In_3900);
or U5232 (N_5232,In_2564,In_3735);
or U5233 (N_5233,In_4400,In_3415);
nand U5234 (N_5234,In_3173,In_2204);
nor U5235 (N_5235,In_4651,In_275);
and U5236 (N_5236,In_4087,In_2030);
xor U5237 (N_5237,In_1041,In_4756);
nand U5238 (N_5238,In_1450,In_2583);
nor U5239 (N_5239,In_4068,In_4391);
or U5240 (N_5240,In_2305,In_1338);
and U5241 (N_5241,In_3141,In_3015);
and U5242 (N_5242,In_3101,In_2751);
and U5243 (N_5243,In_3074,In_3049);
nor U5244 (N_5244,In_3183,In_3035);
nand U5245 (N_5245,In_4682,In_1747);
xnor U5246 (N_5246,In_3127,In_2668);
nor U5247 (N_5247,In_1510,In_1674);
nor U5248 (N_5248,In_3513,In_2076);
nand U5249 (N_5249,In_4739,In_601);
nor U5250 (N_5250,In_2614,In_1878);
nor U5251 (N_5251,In_3483,In_2031);
or U5252 (N_5252,In_4379,In_4684);
and U5253 (N_5253,In_2203,In_4589);
xor U5254 (N_5254,In_3058,In_1411);
or U5255 (N_5255,In_91,In_3725);
and U5256 (N_5256,In_4143,In_681);
xnor U5257 (N_5257,In_4777,In_3521);
and U5258 (N_5258,In_1159,In_1679);
or U5259 (N_5259,In_831,In_80);
nand U5260 (N_5260,In_3859,In_2492);
nand U5261 (N_5261,In_746,In_1441);
nor U5262 (N_5262,In_4209,In_94);
and U5263 (N_5263,In_1422,In_952);
xor U5264 (N_5264,In_2657,In_4734);
nor U5265 (N_5265,In_1659,In_927);
nand U5266 (N_5266,In_1304,In_281);
or U5267 (N_5267,In_2046,In_3599);
nor U5268 (N_5268,In_935,In_1901);
nand U5269 (N_5269,In_4975,In_486);
or U5270 (N_5270,In_3236,In_3313);
nand U5271 (N_5271,In_1467,In_53);
and U5272 (N_5272,In_422,In_3987);
or U5273 (N_5273,In_4354,In_334);
xnor U5274 (N_5274,In_1907,In_2010);
and U5275 (N_5275,In_1196,In_4394);
xnor U5276 (N_5276,In_2829,In_2730);
xnor U5277 (N_5277,In_4339,In_4756);
xor U5278 (N_5278,In_2176,In_534);
nor U5279 (N_5279,In_2533,In_4465);
or U5280 (N_5280,In_2897,In_883);
and U5281 (N_5281,In_3459,In_2891);
nand U5282 (N_5282,In_2058,In_2505);
nor U5283 (N_5283,In_661,In_4108);
nand U5284 (N_5284,In_2676,In_4673);
or U5285 (N_5285,In_4821,In_87);
or U5286 (N_5286,In_2060,In_4629);
and U5287 (N_5287,In_2455,In_3924);
or U5288 (N_5288,In_500,In_4700);
nand U5289 (N_5289,In_4730,In_128);
xnor U5290 (N_5290,In_3426,In_124);
or U5291 (N_5291,In_547,In_1989);
nor U5292 (N_5292,In_3134,In_1593);
and U5293 (N_5293,In_3556,In_2577);
and U5294 (N_5294,In_1936,In_2382);
xor U5295 (N_5295,In_1238,In_4729);
nor U5296 (N_5296,In_1917,In_1527);
xor U5297 (N_5297,In_1398,In_2340);
xnor U5298 (N_5298,In_422,In_3225);
and U5299 (N_5299,In_3883,In_633);
nor U5300 (N_5300,In_89,In_2261);
xor U5301 (N_5301,In_3240,In_795);
or U5302 (N_5302,In_4299,In_1102);
nand U5303 (N_5303,In_3761,In_41);
nand U5304 (N_5304,In_3608,In_2123);
nor U5305 (N_5305,In_3694,In_157);
nor U5306 (N_5306,In_2516,In_4627);
xnor U5307 (N_5307,In_4061,In_2850);
nor U5308 (N_5308,In_3595,In_3985);
and U5309 (N_5309,In_3692,In_3936);
and U5310 (N_5310,In_1483,In_3089);
and U5311 (N_5311,In_2761,In_2175);
or U5312 (N_5312,In_960,In_4872);
or U5313 (N_5313,In_3603,In_3441);
nor U5314 (N_5314,In_4861,In_1789);
xnor U5315 (N_5315,In_1846,In_1778);
xor U5316 (N_5316,In_237,In_2468);
nand U5317 (N_5317,In_3111,In_1225);
and U5318 (N_5318,In_3367,In_1525);
nand U5319 (N_5319,In_509,In_3898);
nand U5320 (N_5320,In_1495,In_4905);
or U5321 (N_5321,In_4143,In_1482);
or U5322 (N_5322,In_2733,In_887);
or U5323 (N_5323,In_2515,In_1685);
nor U5324 (N_5324,In_2904,In_2778);
nand U5325 (N_5325,In_763,In_2878);
nor U5326 (N_5326,In_3436,In_244);
xor U5327 (N_5327,In_4792,In_4916);
xnor U5328 (N_5328,In_2990,In_779);
nand U5329 (N_5329,In_1542,In_428);
and U5330 (N_5330,In_2374,In_338);
nor U5331 (N_5331,In_4836,In_312);
or U5332 (N_5332,In_1603,In_3242);
and U5333 (N_5333,In_3529,In_3493);
and U5334 (N_5334,In_2958,In_1418);
and U5335 (N_5335,In_3026,In_4625);
nand U5336 (N_5336,In_4534,In_3387);
nand U5337 (N_5337,In_1157,In_4412);
xor U5338 (N_5338,In_2550,In_4551);
nand U5339 (N_5339,In_4042,In_1900);
nand U5340 (N_5340,In_1199,In_947);
xor U5341 (N_5341,In_829,In_4815);
nor U5342 (N_5342,In_3231,In_2024);
or U5343 (N_5343,In_2600,In_4126);
xor U5344 (N_5344,In_2993,In_3564);
xor U5345 (N_5345,In_881,In_2967);
nor U5346 (N_5346,In_1735,In_4619);
nor U5347 (N_5347,In_961,In_826);
xor U5348 (N_5348,In_2941,In_2404);
and U5349 (N_5349,In_3735,In_4722);
or U5350 (N_5350,In_2239,In_684);
or U5351 (N_5351,In_3871,In_4895);
or U5352 (N_5352,In_1188,In_4845);
nand U5353 (N_5353,In_3729,In_2318);
nor U5354 (N_5354,In_3871,In_2416);
xor U5355 (N_5355,In_2040,In_3976);
nor U5356 (N_5356,In_2507,In_2052);
or U5357 (N_5357,In_1134,In_855);
nor U5358 (N_5358,In_248,In_1171);
nor U5359 (N_5359,In_3021,In_3312);
and U5360 (N_5360,In_2566,In_1772);
or U5361 (N_5361,In_2756,In_1442);
xor U5362 (N_5362,In_4393,In_3640);
or U5363 (N_5363,In_836,In_723);
xnor U5364 (N_5364,In_4409,In_1814);
or U5365 (N_5365,In_1231,In_2491);
nor U5366 (N_5366,In_770,In_3884);
and U5367 (N_5367,In_3609,In_1739);
nor U5368 (N_5368,In_28,In_4185);
and U5369 (N_5369,In_3874,In_1816);
nand U5370 (N_5370,In_3790,In_124);
or U5371 (N_5371,In_2106,In_880);
and U5372 (N_5372,In_4627,In_939);
nor U5373 (N_5373,In_2966,In_4007);
and U5374 (N_5374,In_2757,In_3056);
nor U5375 (N_5375,In_1836,In_4088);
or U5376 (N_5376,In_2460,In_64);
nor U5377 (N_5377,In_2076,In_1121);
or U5378 (N_5378,In_4894,In_1030);
nand U5379 (N_5379,In_4096,In_18);
or U5380 (N_5380,In_4929,In_1289);
xnor U5381 (N_5381,In_1682,In_52);
or U5382 (N_5382,In_872,In_3068);
xnor U5383 (N_5383,In_1083,In_294);
nor U5384 (N_5384,In_1202,In_3406);
nor U5385 (N_5385,In_4666,In_1927);
nand U5386 (N_5386,In_3431,In_367);
xnor U5387 (N_5387,In_4072,In_3032);
nand U5388 (N_5388,In_1690,In_2048);
or U5389 (N_5389,In_238,In_3571);
and U5390 (N_5390,In_2887,In_2669);
or U5391 (N_5391,In_2421,In_2831);
nand U5392 (N_5392,In_3248,In_3756);
nand U5393 (N_5393,In_1911,In_3951);
nand U5394 (N_5394,In_3361,In_3372);
and U5395 (N_5395,In_4626,In_3981);
nor U5396 (N_5396,In_4566,In_3092);
xnor U5397 (N_5397,In_1925,In_3873);
nand U5398 (N_5398,In_4531,In_1756);
nand U5399 (N_5399,In_2741,In_2098);
and U5400 (N_5400,In_3486,In_2016);
nor U5401 (N_5401,In_4792,In_2228);
nor U5402 (N_5402,In_1366,In_2219);
nor U5403 (N_5403,In_4836,In_1208);
xor U5404 (N_5404,In_4047,In_3044);
xor U5405 (N_5405,In_1554,In_3792);
xor U5406 (N_5406,In_3565,In_4438);
nand U5407 (N_5407,In_2962,In_1236);
nor U5408 (N_5408,In_2133,In_3279);
nand U5409 (N_5409,In_3261,In_1965);
xor U5410 (N_5410,In_47,In_1641);
nand U5411 (N_5411,In_1168,In_3951);
nand U5412 (N_5412,In_1226,In_1136);
nand U5413 (N_5413,In_3859,In_457);
and U5414 (N_5414,In_3985,In_2860);
and U5415 (N_5415,In_335,In_3332);
or U5416 (N_5416,In_1611,In_4959);
or U5417 (N_5417,In_2269,In_2828);
nand U5418 (N_5418,In_4908,In_4652);
and U5419 (N_5419,In_4653,In_2113);
nor U5420 (N_5420,In_899,In_1286);
and U5421 (N_5421,In_188,In_1135);
xor U5422 (N_5422,In_63,In_4910);
xor U5423 (N_5423,In_4071,In_4965);
nor U5424 (N_5424,In_4248,In_3633);
nor U5425 (N_5425,In_3948,In_2788);
xor U5426 (N_5426,In_485,In_1161);
or U5427 (N_5427,In_2156,In_327);
or U5428 (N_5428,In_3955,In_102);
xor U5429 (N_5429,In_2823,In_4596);
and U5430 (N_5430,In_3831,In_2377);
and U5431 (N_5431,In_1268,In_2412);
nor U5432 (N_5432,In_1628,In_3540);
nand U5433 (N_5433,In_4255,In_4437);
or U5434 (N_5434,In_1734,In_3617);
nor U5435 (N_5435,In_2886,In_2672);
nor U5436 (N_5436,In_2963,In_705);
and U5437 (N_5437,In_4887,In_1589);
or U5438 (N_5438,In_771,In_3521);
or U5439 (N_5439,In_828,In_2976);
nor U5440 (N_5440,In_2209,In_1868);
nor U5441 (N_5441,In_2404,In_783);
nor U5442 (N_5442,In_4378,In_86);
xor U5443 (N_5443,In_2286,In_2403);
nor U5444 (N_5444,In_4404,In_4478);
nor U5445 (N_5445,In_4266,In_2880);
nor U5446 (N_5446,In_1614,In_4070);
and U5447 (N_5447,In_4513,In_182);
xor U5448 (N_5448,In_3052,In_4596);
or U5449 (N_5449,In_3273,In_0);
xor U5450 (N_5450,In_1924,In_1821);
nand U5451 (N_5451,In_3944,In_4943);
xor U5452 (N_5452,In_2620,In_3980);
nand U5453 (N_5453,In_3925,In_4420);
nor U5454 (N_5454,In_2518,In_3297);
and U5455 (N_5455,In_132,In_2043);
nor U5456 (N_5456,In_1986,In_2116);
nand U5457 (N_5457,In_4654,In_4180);
or U5458 (N_5458,In_1182,In_3923);
nor U5459 (N_5459,In_4170,In_4393);
and U5460 (N_5460,In_906,In_998);
or U5461 (N_5461,In_4399,In_2278);
xor U5462 (N_5462,In_147,In_3413);
and U5463 (N_5463,In_4164,In_1648);
and U5464 (N_5464,In_714,In_3015);
nand U5465 (N_5465,In_3378,In_3973);
nand U5466 (N_5466,In_3205,In_1489);
or U5467 (N_5467,In_81,In_926);
or U5468 (N_5468,In_3668,In_3427);
or U5469 (N_5469,In_42,In_572);
nand U5470 (N_5470,In_2367,In_1413);
and U5471 (N_5471,In_2639,In_1186);
and U5472 (N_5472,In_905,In_3475);
or U5473 (N_5473,In_2489,In_4858);
xnor U5474 (N_5474,In_3256,In_3490);
xor U5475 (N_5475,In_3561,In_3869);
and U5476 (N_5476,In_751,In_4006);
and U5477 (N_5477,In_3074,In_906);
nand U5478 (N_5478,In_1236,In_526);
and U5479 (N_5479,In_4641,In_1877);
nand U5480 (N_5480,In_418,In_3929);
nor U5481 (N_5481,In_3265,In_2288);
nand U5482 (N_5482,In_3488,In_4134);
and U5483 (N_5483,In_889,In_395);
nand U5484 (N_5484,In_1472,In_1365);
nand U5485 (N_5485,In_2050,In_997);
nand U5486 (N_5486,In_4880,In_1034);
xnor U5487 (N_5487,In_4401,In_4878);
nand U5488 (N_5488,In_976,In_623);
and U5489 (N_5489,In_3875,In_2);
nor U5490 (N_5490,In_2279,In_1347);
and U5491 (N_5491,In_2755,In_471);
and U5492 (N_5492,In_1658,In_1010);
nor U5493 (N_5493,In_647,In_3133);
or U5494 (N_5494,In_3880,In_1488);
or U5495 (N_5495,In_3700,In_424);
and U5496 (N_5496,In_1659,In_4350);
and U5497 (N_5497,In_2927,In_1724);
nand U5498 (N_5498,In_4619,In_4776);
and U5499 (N_5499,In_460,In_2111);
and U5500 (N_5500,In_4404,In_1626);
xor U5501 (N_5501,In_4104,In_3120);
xnor U5502 (N_5502,In_4789,In_1924);
and U5503 (N_5503,In_1437,In_4526);
and U5504 (N_5504,In_1465,In_3737);
or U5505 (N_5505,In_1332,In_4425);
and U5506 (N_5506,In_4809,In_4741);
xnor U5507 (N_5507,In_4056,In_698);
or U5508 (N_5508,In_180,In_1564);
and U5509 (N_5509,In_4072,In_2502);
xor U5510 (N_5510,In_2075,In_53);
nor U5511 (N_5511,In_4823,In_4471);
and U5512 (N_5512,In_2318,In_1147);
xnor U5513 (N_5513,In_323,In_1150);
nor U5514 (N_5514,In_2968,In_3970);
xor U5515 (N_5515,In_3387,In_1979);
and U5516 (N_5516,In_1169,In_3770);
or U5517 (N_5517,In_228,In_39);
or U5518 (N_5518,In_3427,In_229);
or U5519 (N_5519,In_2979,In_1678);
xor U5520 (N_5520,In_4784,In_1547);
nor U5521 (N_5521,In_421,In_4796);
nand U5522 (N_5522,In_4627,In_3721);
and U5523 (N_5523,In_3822,In_3878);
xnor U5524 (N_5524,In_1109,In_2718);
xor U5525 (N_5525,In_4882,In_4226);
and U5526 (N_5526,In_2123,In_2168);
nor U5527 (N_5527,In_4252,In_1579);
nand U5528 (N_5528,In_2195,In_2137);
or U5529 (N_5529,In_4726,In_620);
and U5530 (N_5530,In_4139,In_4005);
and U5531 (N_5531,In_27,In_3240);
or U5532 (N_5532,In_4337,In_4052);
and U5533 (N_5533,In_2970,In_2283);
xnor U5534 (N_5534,In_3674,In_599);
nand U5535 (N_5535,In_1794,In_3347);
or U5536 (N_5536,In_4538,In_2803);
nand U5537 (N_5537,In_2461,In_168);
xor U5538 (N_5538,In_1610,In_133);
nand U5539 (N_5539,In_2075,In_4828);
and U5540 (N_5540,In_2149,In_513);
xor U5541 (N_5541,In_3208,In_4643);
nor U5542 (N_5542,In_2787,In_898);
nand U5543 (N_5543,In_3453,In_4420);
and U5544 (N_5544,In_1794,In_4264);
xor U5545 (N_5545,In_145,In_1998);
or U5546 (N_5546,In_2875,In_472);
nand U5547 (N_5547,In_3397,In_4929);
nor U5548 (N_5548,In_1182,In_4345);
nor U5549 (N_5549,In_1670,In_1700);
xor U5550 (N_5550,In_1949,In_1803);
or U5551 (N_5551,In_1761,In_4073);
and U5552 (N_5552,In_4025,In_1937);
or U5553 (N_5553,In_4280,In_472);
xnor U5554 (N_5554,In_4156,In_1603);
xnor U5555 (N_5555,In_989,In_4653);
or U5556 (N_5556,In_1316,In_3918);
nand U5557 (N_5557,In_456,In_1543);
nand U5558 (N_5558,In_2074,In_2572);
xnor U5559 (N_5559,In_4826,In_816);
xnor U5560 (N_5560,In_565,In_1611);
or U5561 (N_5561,In_4279,In_3417);
and U5562 (N_5562,In_375,In_4665);
xnor U5563 (N_5563,In_469,In_3061);
nand U5564 (N_5564,In_4981,In_4027);
nor U5565 (N_5565,In_1207,In_238);
and U5566 (N_5566,In_893,In_481);
nor U5567 (N_5567,In_577,In_3581);
and U5568 (N_5568,In_4735,In_3204);
or U5569 (N_5569,In_56,In_307);
nor U5570 (N_5570,In_715,In_2223);
nor U5571 (N_5571,In_2039,In_4140);
nand U5572 (N_5572,In_1045,In_669);
and U5573 (N_5573,In_3842,In_3733);
or U5574 (N_5574,In_2872,In_4113);
nor U5575 (N_5575,In_4917,In_3913);
or U5576 (N_5576,In_362,In_107);
nor U5577 (N_5577,In_3750,In_454);
nand U5578 (N_5578,In_1893,In_2001);
nand U5579 (N_5579,In_3511,In_2590);
or U5580 (N_5580,In_496,In_4120);
or U5581 (N_5581,In_2781,In_3760);
nor U5582 (N_5582,In_972,In_157);
and U5583 (N_5583,In_946,In_1149);
nand U5584 (N_5584,In_4972,In_1969);
or U5585 (N_5585,In_4918,In_1269);
or U5586 (N_5586,In_1995,In_3779);
or U5587 (N_5587,In_3665,In_4277);
and U5588 (N_5588,In_1880,In_1779);
and U5589 (N_5589,In_156,In_2218);
or U5590 (N_5590,In_513,In_4266);
xnor U5591 (N_5591,In_4693,In_2886);
xnor U5592 (N_5592,In_4413,In_3014);
nand U5593 (N_5593,In_4475,In_4988);
xor U5594 (N_5594,In_510,In_2596);
xor U5595 (N_5595,In_2712,In_743);
nor U5596 (N_5596,In_3538,In_4404);
nand U5597 (N_5597,In_1349,In_700);
xor U5598 (N_5598,In_461,In_4318);
nor U5599 (N_5599,In_1905,In_4354);
and U5600 (N_5600,In_3931,In_325);
and U5601 (N_5601,In_468,In_1317);
nor U5602 (N_5602,In_536,In_1953);
nor U5603 (N_5603,In_3272,In_3373);
nor U5604 (N_5604,In_4570,In_3817);
nand U5605 (N_5605,In_4634,In_4895);
nor U5606 (N_5606,In_2193,In_2386);
nand U5607 (N_5607,In_1285,In_4067);
xor U5608 (N_5608,In_1957,In_2949);
nor U5609 (N_5609,In_1349,In_2829);
nor U5610 (N_5610,In_4033,In_4896);
or U5611 (N_5611,In_3421,In_114);
and U5612 (N_5612,In_3656,In_4359);
xnor U5613 (N_5613,In_4204,In_1275);
nand U5614 (N_5614,In_816,In_4267);
or U5615 (N_5615,In_967,In_593);
nor U5616 (N_5616,In_659,In_3600);
xor U5617 (N_5617,In_1839,In_2326);
xor U5618 (N_5618,In_2652,In_2920);
or U5619 (N_5619,In_1044,In_3415);
nand U5620 (N_5620,In_1902,In_1327);
nand U5621 (N_5621,In_413,In_4499);
nand U5622 (N_5622,In_3102,In_4436);
nand U5623 (N_5623,In_4499,In_3215);
xnor U5624 (N_5624,In_3971,In_3714);
nand U5625 (N_5625,In_3437,In_386);
xnor U5626 (N_5626,In_4198,In_1768);
or U5627 (N_5627,In_1418,In_3504);
nand U5628 (N_5628,In_819,In_254);
nand U5629 (N_5629,In_3203,In_3290);
or U5630 (N_5630,In_2014,In_2638);
xor U5631 (N_5631,In_2472,In_1291);
or U5632 (N_5632,In_1809,In_4564);
and U5633 (N_5633,In_1339,In_3384);
xor U5634 (N_5634,In_4879,In_4818);
xor U5635 (N_5635,In_924,In_177);
and U5636 (N_5636,In_3594,In_1122);
nand U5637 (N_5637,In_1776,In_287);
and U5638 (N_5638,In_3255,In_1116);
nor U5639 (N_5639,In_3740,In_3614);
or U5640 (N_5640,In_2446,In_1564);
xnor U5641 (N_5641,In_1374,In_1523);
nand U5642 (N_5642,In_2562,In_3598);
nand U5643 (N_5643,In_3608,In_1293);
or U5644 (N_5644,In_2974,In_76);
xor U5645 (N_5645,In_189,In_4209);
or U5646 (N_5646,In_3104,In_331);
nand U5647 (N_5647,In_4296,In_4596);
and U5648 (N_5648,In_208,In_4409);
xor U5649 (N_5649,In_1619,In_2262);
nand U5650 (N_5650,In_4743,In_2195);
or U5651 (N_5651,In_2489,In_4746);
and U5652 (N_5652,In_807,In_3630);
nor U5653 (N_5653,In_202,In_2959);
nand U5654 (N_5654,In_4951,In_3998);
or U5655 (N_5655,In_2627,In_3026);
nand U5656 (N_5656,In_419,In_932);
or U5657 (N_5657,In_2359,In_2951);
nand U5658 (N_5658,In_630,In_1511);
or U5659 (N_5659,In_4526,In_4253);
nand U5660 (N_5660,In_3939,In_4727);
nor U5661 (N_5661,In_3711,In_3078);
and U5662 (N_5662,In_2672,In_2185);
nor U5663 (N_5663,In_1412,In_2144);
xor U5664 (N_5664,In_1411,In_248);
and U5665 (N_5665,In_4075,In_521);
nand U5666 (N_5666,In_2526,In_4224);
and U5667 (N_5667,In_309,In_751);
xnor U5668 (N_5668,In_3670,In_4359);
xnor U5669 (N_5669,In_4488,In_862);
or U5670 (N_5670,In_2082,In_740);
nor U5671 (N_5671,In_16,In_4696);
nor U5672 (N_5672,In_680,In_173);
or U5673 (N_5673,In_52,In_565);
nor U5674 (N_5674,In_13,In_965);
or U5675 (N_5675,In_2607,In_3782);
xnor U5676 (N_5676,In_748,In_1579);
nor U5677 (N_5677,In_4526,In_3466);
nor U5678 (N_5678,In_4584,In_1129);
nand U5679 (N_5679,In_850,In_2325);
and U5680 (N_5680,In_951,In_3042);
and U5681 (N_5681,In_4207,In_3087);
nor U5682 (N_5682,In_1756,In_1874);
nor U5683 (N_5683,In_1098,In_884);
and U5684 (N_5684,In_1552,In_1307);
xnor U5685 (N_5685,In_2260,In_4799);
nor U5686 (N_5686,In_1047,In_1855);
and U5687 (N_5687,In_3812,In_137);
and U5688 (N_5688,In_3667,In_803);
or U5689 (N_5689,In_597,In_3307);
xor U5690 (N_5690,In_1444,In_2139);
or U5691 (N_5691,In_3054,In_676);
and U5692 (N_5692,In_2646,In_2497);
or U5693 (N_5693,In_3738,In_1335);
nor U5694 (N_5694,In_59,In_4115);
or U5695 (N_5695,In_4774,In_4859);
xnor U5696 (N_5696,In_3768,In_4917);
and U5697 (N_5697,In_3167,In_1052);
xor U5698 (N_5698,In_4038,In_752);
and U5699 (N_5699,In_375,In_2656);
xor U5700 (N_5700,In_189,In_577);
and U5701 (N_5701,In_3917,In_3984);
and U5702 (N_5702,In_2791,In_3321);
nor U5703 (N_5703,In_3849,In_318);
and U5704 (N_5704,In_1422,In_258);
xnor U5705 (N_5705,In_2011,In_3071);
xnor U5706 (N_5706,In_4076,In_3402);
nand U5707 (N_5707,In_3001,In_1387);
nor U5708 (N_5708,In_267,In_3236);
and U5709 (N_5709,In_1606,In_1118);
nor U5710 (N_5710,In_2715,In_3861);
and U5711 (N_5711,In_4849,In_3003);
and U5712 (N_5712,In_19,In_2303);
xnor U5713 (N_5713,In_3447,In_4719);
nor U5714 (N_5714,In_299,In_4124);
nand U5715 (N_5715,In_4832,In_3659);
xor U5716 (N_5716,In_2060,In_4238);
nor U5717 (N_5717,In_2975,In_500);
nand U5718 (N_5718,In_4122,In_3869);
nand U5719 (N_5719,In_3399,In_768);
xnor U5720 (N_5720,In_1795,In_1889);
nor U5721 (N_5721,In_3632,In_2664);
and U5722 (N_5722,In_77,In_2404);
nand U5723 (N_5723,In_4498,In_4579);
and U5724 (N_5724,In_4744,In_3589);
or U5725 (N_5725,In_1845,In_1175);
nor U5726 (N_5726,In_311,In_1292);
nor U5727 (N_5727,In_4838,In_4052);
or U5728 (N_5728,In_3453,In_1886);
nand U5729 (N_5729,In_4978,In_3501);
or U5730 (N_5730,In_2450,In_2214);
nor U5731 (N_5731,In_1547,In_520);
xor U5732 (N_5732,In_3801,In_3680);
or U5733 (N_5733,In_1025,In_2320);
and U5734 (N_5734,In_574,In_1596);
nor U5735 (N_5735,In_3490,In_4806);
or U5736 (N_5736,In_3482,In_1035);
xor U5737 (N_5737,In_2733,In_867);
nor U5738 (N_5738,In_4175,In_1199);
or U5739 (N_5739,In_4501,In_4548);
xnor U5740 (N_5740,In_632,In_3387);
nand U5741 (N_5741,In_1992,In_1600);
or U5742 (N_5742,In_4083,In_4655);
xor U5743 (N_5743,In_287,In_2714);
or U5744 (N_5744,In_1431,In_4968);
nor U5745 (N_5745,In_4619,In_4910);
nor U5746 (N_5746,In_1545,In_168);
and U5747 (N_5747,In_2760,In_122);
and U5748 (N_5748,In_2745,In_2043);
or U5749 (N_5749,In_1741,In_2434);
or U5750 (N_5750,In_1147,In_3977);
and U5751 (N_5751,In_3254,In_3374);
nand U5752 (N_5752,In_3145,In_2504);
xnor U5753 (N_5753,In_1517,In_2910);
nand U5754 (N_5754,In_4067,In_2700);
and U5755 (N_5755,In_2138,In_1008);
nand U5756 (N_5756,In_2372,In_4036);
nand U5757 (N_5757,In_1585,In_2293);
nand U5758 (N_5758,In_2220,In_1660);
nand U5759 (N_5759,In_85,In_1577);
nor U5760 (N_5760,In_3382,In_38);
nand U5761 (N_5761,In_2965,In_2854);
or U5762 (N_5762,In_150,In_3186);
xnor U5763 (N_5763,In_836,In_3310);
and U5764 (N_5764,In_3453,In_3971);
nand U5765 (N_5765,In_1068,In_1209);
and U5766 (N_5766,In_1349,In_1285);
nor U5767 (N_5767,In_3673,In_386);
and U5768 (N_5768,In_870,In_2483);
or U5769 (N_5769,In_2053,In_1142);
nand U5770 (N_5770,In_1571,In_4183);
or U5771 (N_5771,In_588,In_1479);
or U5772 (N_5772,In_1198,In_791);
nand U5773 (N_5773,In_4080,In_1323);
nand U5774 (N_5774,In_1139,In_2436);
xor U5775 (N_5775,In_649,In_2457);
nand U5776 (N_5776,In_1613,In_2118);
or U5777 (N_5777,In_1650,In_2872);
and U5778 (N_5778,In_1271,In_3081);
or U5779 (N_5779,In_2628,In_1714);
nand U5780 (N_5780,In_1738,In_1182);
or U5781 (N_5781,In_2833,In_1518);
nor U5782 (N_5782,In_3214,In_2165);
xor U5783 (N_5783,In_3570,In_1066);
and U5784 (N_5784,In_3534,In_1522);
and U5785 (N_5785,In_2546,In_430);
and U5786 (N_5786,In_3900,In_1891);
nor U5787 (N_5787,In_1321,In_1916);
and U5788 (N_5788,In_1596,In_4963);
xor U5789 (N_5789,In_2210,In_2869);
nand U5790 (N_5790,In_3988,In_4674);
nor U5791 (N_5791,In_2337,In_3483);
nor U5792 (N_5792,In_3281,In_3897);
and U5793 (N_5793,In_4067,In_202);
nor U5794 (N_5794,In_4348,In_2700);
or U5795 (N_5795,In_4253,In_3100);
nand U5796 (N_5796,In_205,In_1240);
xnor U5797 (N_5797,In_2684,In_1890);
or U5798 (N_5798,In_1578,In_2607);
and U5799 (N_5799,In_2592,In_3255);
or U5800 (N_5800,In_2676,In_42);
nand U5801 (N_5801,In_1919,In_3098);
nor U5802 (N_5802,In_4918,In_4453);
and U5803 (N_5803,In_2004,In_4864);
nor U5804 (N_5804,In_3150,In_3168);
xor U5805 (N_5805,In_3467,In_1951);
and U5806 (N_5806,In_1333,In_3789);
xor U5807 (N_5807,In_2315,In_2216);
nand U5808 (N_5808,In_2516,In_642);
nor U5809 (N_5809,In_1216,In_4094);
and U5810 (N_5810,In_2989,In_1975);
nand U5811 (N_5811,In_2108,In_1543);
xor U5812 (N_5812,In_747,In_4298);
xnor U5813 (N_5813,In_3007,In_4429);
nor U5814 (N_5814,In_3488,In_1370);
nand U5815 (N_5815,In_3926,In_1307);
nand U5816 (N_5816,In_1117,In_2440);
nand U5817 (N_5817,In_2193,In_509);
xnor U5818 (N_5818,In_121,In_2990);
nand U5819 (N_5819,In_951,In_3788);
and U5820 (N_5820,In_795,In_2761);
and U5821 (N_5821,In_1457,In_3421);
and U5822 (N_5822,In_4652,In_2141);
and U5823 (N_5823,In_1280,In_197);
xnor U5824 (N_5824,In_3193,In_1266);
and U5825 (N_5825,In_2439,In_4187);
nor U5826 (N_5826,In_3188,In_3044);
and U5827 (N_5827,In_3029,In_4642);
xnor U5828 (N_5828,In_357,In_4354);
xnor U5829 (N_5829,In_1197,In_4650);
nand U5830 (N_5830,In_617,In_1411);
xnor U5831 (N_5831,In_3020,In_2913);
or U5832 (N_5832,In_3782,In_3280);
and U5833 (N_5833,In_3162,In_4692);
xor U5834 (N_5834,In_739,In_2824);
or U5835 (N_5835,In_4168,In_3028);
xnor U5836 (N_5836,In_760,In_1459);
nor U5837 (N_5837,In_808,In_4887);
nand U5838 (N_5838,In_3425,In_249);
and U5839 (N_5839,In_394,In_3636);
nand U5840 (N_5840,In_4180,In_1459);
and U5841 (N_5841,In_2808,In_3845);
nor U5842 (N_5842,In_3230,In_1005);
and U5843 (N_5843,In_3039,In_854);
nand U5844 (N_5844,In_3666,In_4038);
xor U5845 (N_5845,In_3308,In_762);
and U5846 (N_5846,In_2003,In_4471);
xor U5847 (N_5847,In_3144,In_3627);
and U5848 (N_5848,In_2703,In_4208);
xor U5849 (N_5849,In_241,In_1844);
or U5850 (N_5850,In_499,In_4115);
xor U5851 (N_5851,In_486,In_4876);
nand U5852 (N_5852,In_1132,In_4875);
or U5853 (N_5853,In_4232,In_1873);
or U5854 (N_5854,In_300,In_2534);
nor U5855 (N_5855,In_1628,In_2776);
xnor U5856 (N_5856,In_4316,In_4768);
and U5857 (N_5857,In_2547,In_9);
xor U5858 (N_5858,In_144,In_600);
nand U5859 (N_5859,In_1639,In_4899);
nand U5860 (N_5860,In_1082,In_1976);
and U5861 (N_5861,In_560,In_2669);
and U5862 (N_5862,In_487,In_3171);
nor U5863 (N_5863,In_4093,In_642);
and U5864 (N_5864,In_3326,In_4792);
and U5865 (N_5865,In_1870,In_218);
xor U5866 (N_5866,In_3710,In_1311);
or U5867 (N_5867,In_1557,In_1382);
and U5868 (N_5868,In_3965,In_1007);
xor U5869 (N_5869,In_3187,In_2734);
xnor U5870 (N_5870,In_4195,In_3381);
and U5871 (N_5871,In_3359,In_4289);
nor U5872 (N_5872,In_2614,In_1347);
nor U5873 (N_5873,In_3730,In_3291);
nand U5874 (N_5874,In_99,In_4847);
xor U5875 (N_5875,In_1907,In_69);
nand U5876 (N_5876,In_1420,In_3580);
nor U5877 (N_5877,In_205,In_1632);
xnor U5878 (N_5878,In_2309,In_817);
nand U5879 (N_5879,In_825,In_3461);
or U5880 (N_5880,In_4431,In_4744);
or U5881 (N_5881,In_1288,In_2803);
nor U5882 (N_5882,In_3344,In_1450);
xor U5883 (N_5883,In_1292,In_1102);
nor U5884 (N_5884,In_2324,In_1241);
or U5885 (N_5885,In_2301,In_1998);
nor U5886 (N_5886,In_1618,In_4155);
or U5887 (N_5887,In_616,In_2198);
nand U5888 (N_5888,In_1892,In_1359);
nand U5889 (N_5889,In_2160,In_1990);
and U5890 (N_5890,In_349,In_1154);
nand U5891 (N_5891,In_3490,In_3291);
xnor U5892 (N_5892,In_1876,In_1680);
nand U5893 (N_5893,In_1998,In_2154);
or U5894 (N_5894,In_4059,In_972);
and U5895 (N_5895,In_4678,In_1644);
and U5896 (N_5896,In_2235,In_4235);
xnor U5897 (N_5897,In_3917,In_2711);
or U5898 (N_5898,In_2497,In_3783);
nand U5899 (N_5899,In_979,In_2993);
nor U5900 (N_5900,In_1781,In_4901);
or U5901 (N_5901,In_4057,In_2847);
nand U5902 (N_5902,In_4742,In_1443);
and U5903 (N_5903,In_3633,In_3961);
or U5904 (N_5904,In_4415,In_2478);
nor U5905 (N_5905,In_2653,In_2998);
xor U5906 (N_5906,In_4176,In_3567);
nand U5907 (N_5907,In_988,In_3035);
or U5908 (N_5908,In_4451,In_1652);
xor U5909 (N_5909,In_4916,In_1709);
xor U5910 (N_5910,In_588,In_376);
nand U5911 (N_5911,In_4460,In_2097);
or U5912 (N_5912,In_1945,In_1564);
nand U5913 (N_5913,In_2423,In_4665);
nor U5914 (N_5914,In_4354,In_2053);
and U5915 (N_5915,In_365,In_194);
nor U5916 (N_5916,In_2403,In_1074);
nand U5917 (N_5917,In_349,In_1875);
nand U5918 (N_5918,In_72,In_3405);
xor U5919 (N_5919,In_3904,In_2215);
xor U5920 (N_5920,In_4787,In_588);
or U5921 (N_5921,In_3190,In_4475);
xor U5922 (N_5922,In_829,In_3368);
or U5923 (N_5923,In_3416,In_4342);
xnor U5924 (N_5924,In_3700,In_2027);
xor U5925 (N_5925,In_4975,In_3458);
nor U5926 (N_5926,In_2632,In_1492);
and U5927 (N_5927,In_2759,In_215);
xnor U5928 (N_5928,In_4704,In_4632);
nor U5929 (N_5929,In_2070,In_1145);
and U5930 (N_5930,In_3054,In_1710);
xor U5931 (N_5931,In_551,In_2727);
and U5932 (N_5932,In_3964,In_3596);
or U5933 (N_5933,In_931,In_2535);
and U5934 (N_5934,In_1547,In_4877);
xnor U5935 (N_5935,In_442,In_887);
and U5936 (N_5936,In_3388,In_541);
nand U5937 (N_5937,In_1336,In_2006);
and U5938 (N_5938,In_4739,In_3831);
nand U5939 (N_5939,In_3179,In_1881);
and U5940 (N_5940,In_4794,In_3643);
nand U5941 (N_5941,In_17,In_2286);
nand U5942 (N_5942,In_106,In_3155);
nand U5943 (N_5943,In_1920,In_236);
xnor U5944 (N_5944,In_2486,In_3445);
xnor U5945 (N_5945,In_188,In_4621);
and U5946 (N_5946,In_38,In_2582);
nor U5947 (N_5947,In_3347,In_3348);
xor U5948 (N_5948,In_1550,In_1541);
nand U5949 (N_5949,In_1305,In_1679);
and U5950 (N_5950,In_3771,In_1234);
nor U5951 (N_5951,In_775,In_399);
nand U5952 (N_5952,In_2651,In_4959);
or U5953 (N_5953,In_4426,In_307);
and U5954 (N_5954,In_712,In_2111);
nand U5955 (N_5955,In_2537,In_710);
and U5956 (N_5956,In_3057,In_4399);
xnor U5957 (N_5957,In_1592,In_1317);
or U5958 (N_5958,In_2944,In_4577);
nor U5959 (N_5959,In_3318,In_4760);
xor U5960 (N_5960,In_272,In_1272);
xor U5961 (N_5961,In_4040,In_3994);
and U5962 (N_5962,In_4601,In_4371);
and U5963 (N_5963,In_3450,In_4959);
nand U5964 (N_5964,In_4720,In_293);
nor U5965 (N_5965,In_2023,In_1494);
nand U5966 (N_5966,In_1940,In_670);
nand U5967 (N_5967,In_4767,In_862);
xor U5968 (N_5968,In_2703,In_3497);
nand U5969 (N_5969,In_1531,In_3169);
nor U5970 (N_5970,In_2806,In_3724);
and U5971 (N_5971,In_2370,In_593);
nand U5972 (N_5972,In_3254,In_3234);
nand U5973 (N_5973,In_4511,In_4088);
nand U5974 (N_5974,In_2430,In_4359);
nand U5975 (N_5975,In_935,In_3314);
xor U5976 (N_5976,In_3771,In_4470);
or U5977 (N_5977,In_4092,In_1431);
nor U5978 (N_5978,In_3293,In_4425);
xor U5979 (N_5979,In_1989,In_1032);
nor U5980 (N_5980,In_3,In_511);
nand U5981 (N_5981,In_810,In_2490);
xnor U5982 (N_5982,In_2372,In_3254);
or U5983 (N_5983,In_4688,In_2667);
or U5984 (N_5984,In_3361,In_3575);
nand U5985 (N_5985,In_2384,In_316);
or U5986 (N_5986,In_4392,In_3210);
nor U5987 (N_5987,In_3723,In_4618);
nor U5988 (N_5988,In_1809,In_3829);
nor U5989 (N_5989,In_980,In_4634);
and U5990 (N_5990,In_4461,In_3555);
and U5991 (N_5991,In_2486,In_1815);
or U5992 (N_5992,In_2834,In_2093);
and U5993 (N_5993,In_1906,In_2757);
xor U5994 (N_5994,In_4355,In_2186);
nand U5995 (N_5995,In_122,In_1076);
and U5996 (N_5996,In_692,In_417);
and U5997 (N_5997,In_1885,In_1742);
nor U5998 (N_5998,In_4340,In_4648);
nor U5999 (N_5999,In_2417,In_4820);
xor U6000 (N_6000,In_2383,In_3017);
and U6001 (N_6001,In_2723,In_3349);
xor U6002 (N_6002,In_3043,In_2325);
nor U6003 (N_6003,In_1458,In_573);
and U6004 (N_6004,In_463,In_4243);
nor U6005 (N_6005,In_3914,In_305);
nor U6006 (N_6006,In_2314,In_4149);
xor U6007 (N_6007,In_3246,In_3014);
nor U6008 (N_6008,In_4186,In_779);
nor U6009 (N_6009,In_978,In_1290);
or U6010 (N_6010,In_2979,In_1979);
or U6011 (N_6011,In_1220,In_3685);
xor U6012 (N_6012,In_3061,In_2605);
nor U6013 (N_6013,In_3613,In_374);
nand U6014 (N_6014,In_1041,In_2137);
and U6015 (N_6015,In_3119,In_1009);
and U6016 (N_6016,In_889,In_996);
nor U6017 (N_6017,In_2175,In_2141);
xor U6018 (N_6018,In_807,In_2068);
and U6019 (N_6019,In_1313,In_3430);
and U6020 (N_6020,In_2228,In_3356);
nand U6021 (N_6021,In_3407,In_2326);
nor U6022 (N_6022,In_840,In_1131);
nor U6023 (N_6023,In_1629,In_4971);
and U6024 (N_6024,In_4208,In_2694);
nor U6025 (N_6025,In_925,In_3161);
nor U6026 (N_6026,In_2611,In_840);
xor U6027 (N_6027,In_3318,In_3313);
nor U6028 (N_6028,In_116,In_3038);
and U6029 (N_6029,In_4610,In_4668);
xnor U6030 (N_6030,In_2741,In_3621);
xor U6031 (N_6031,In_1280,In_641);
nand U6032 (N_6032,In_3664,In_2321);
nor U6033 (N_6033,In_4756,In_2434);
nand U6034 (N_6034,In_3645,In_1877);
and U6035 (N_6035,In_3444,In_3659);
or U6036 (N_6036,In_1858,In_1812);
nor U6037 (N_6037,In_3913,In_575);
xnor U6038 (N_6038,In_3576,In_643);
nor U6039 (N_6039,In_1165,In_1878);
and U6040 (N_6040,In_1651,In_3242);
nor U6041 (N_6041,In_3666,In_519);
nor U6042 (N_6042,In_854,In_2800);
xor U6043 (N_6043,In_4311,In_4895);
or U6044 (N_6044,In_4359,In_3677);
and U6045 (N_6045,In_601,In_1914);
or U6046 (N_6046,In_414,In_3723);
nor U6047 (N_6047,In_364,In_3166);
nor U6048 (N_6048,In_1998,In_1006);
nand U6049 (N_6049,In_3966,In_3824);
or U6050 (N_6050,In_3433,In_1607);
nor U6051 (N_6051,In_1194,In_1555);
nor U6052 (N_6052,In_310,In_1785);
xnor U6053 (N_6053,In_2904,In_3609);
or U6054 (N_6054,In_4537,In_2337);
nand U6055 (N_6055,In_620,In_736);
or U6056 (N_6056,In_523,In_2357);
nor U6057 (N_6057,In_3396,In_4875);
and U6058 (N_6058,In_4380,In_3222);
and U6059 (N_6059,In_1504,In_4297);
nor U6060 (N_6060,In_1187,In_4113);
xor U6061 (N_6061,In_4104,In_62);
xor U6062 (N_6062,In_3905,In_2341);
nand U6063 (N_6063,In_1483,In_4914);
xor U6064 (N_6064,In_1767,In_938);
nand U6065 (N_6065,In_455,In_2476);
and U6066 (N_6066,In_1283,In_3983);
nor U6067 (N_6067,In_4174,In_337);
or U6068 (N_6068,In_2254,In_4550);
nor U6069 (N_6069,In_1834,In_3166);
xor U6070 (N_6070,In_833,In_3949);
nand U6071 (N_6071,In_3537,In_304);
and U6072 (N_6072,In_21,In_898);
nor U6073 (N_6073,In_2015,In_4061);
and U6074 (N_6074,In_1809,In_3614);
nand U6075 (N_6075,In_3652,In_73);
xnor U6076 (N_6076,In_553,In_4292);
or U6077 (N_6077,In_4260,In_2049);
nand U6078 (N_6078,In_2679,In_2216);
nor U6079 (N_6079,In_1184,In_1986);
or U6080 (N_6080,In_4401,In_671);
and U6081 (N_6081,In_4303,In_2109);
nand U6082 (N_6082,In_232,In_610);
nor U6083 (N_6083,In_274,In_3836);
nand U6084 (N_6084,In_1110,In_2795);
nor U6085 (N_6085,In_4390,In_4724);
or U6086 (N_6086,In_2562,In_417);
and U6087 (N_6087,In_1304,In_1343);
nor U6088 (N_6088,In_1008,In_1041);
xor U6089 (N_6089,In_599,In_566);
nand U6090 (N_6090,In_4819,In_1643);
xor U6091 (N_6091,In_2454,In_1);
xnor U6092 (N_6092,In_1871,In_1120);
or U6093 (N_6093,In_1342,In_4435);
or U6094 (N_6094,In_548,In_3924);
or U6095 (N_6095,In_4832,In_3246);
nor U6096 (N_6096,In_3444,In_1437);
nor U6097 (N_6097,In_1898,In_1344);
nor U6098 (N_6098,In_3515,In_4913);
xor U6099 (N_6099,In_2193,In_4746);
nand U6100 (N_6100,In_945,In_4500);
xnor U6101 (N_6101,In_2544,In_859);
nor U6102 (N_6102,In_531,In_667);
or U6103 (N_6103,In_312,In_30);
nor U6104 (N_6104,In_1924,In_4035);
nand U6105 (N_6105,In_3099,In_3717);
xor U6106 (N_6106,In_1039,In_242);
and U6107 (N_6107,In_4396,In_3582);
nand U6108 (N_6108,In_3638,In_4688);
and U6109 (N_6109,In_2207,In_893);
nor U6110 (N_6110,In_4486,In_940);
nand U6111 (N_6111,In_2629,In_1712);
nor U6112 (N_6112,In_3289,In_4343);
nor U6113 (N_6113,In_4633,In_2130);
nand U6114 (N_6114,In_4530,In_4095);
nor U6115 (N_6115,In_4226,In_681);
xor U6116 (N_6116,In_2535,In_2539);
nor U6117 (N_6117,In_2314,In_201);
or U6118 (N_6118,In_4249,In_2513);
nand U6119 (N_6119,In_4986,In_3216);
xor U6120 (N_6120,In_1180,In_2607);
and U6121 (N_6121,In_4608,In_574);
and U6122 (N_6122,In_222,In_4633);
nand U6123 (N_6123,In_1467,In_4651);
xor U6124 (N_6124,In_412,In_2622);
nand U6125 (N_6125,In_3330,In_545);
nand U6126 (N_6126,In_4212,In_656);
xor U6127 (N_6127,In_132,In_3983);
xnor U6128 (N_6128,In_2049,In_1418);
xor U6129 (N_6129,In_1329,In_4786);
or U6130 (N_6130,In_3644,In_3816);
or U6131 (N_6131,In_4356,In_1708);
xor U6132 (N_6132,In_1465,In_2107);
nand U6133 (N_6133,In_3691,In_3651);
and U6134 (N_6134,In_4664,In_4867);
or U6135 (N_6135,In_1845,In_1434);
and U6136 (N_6136,In_3565,In_1351);
or U6137 (N_6137,In_3287,In_900);
xor U6138 (N_6138,In_609,In_4247);
nand U6139 (N_6139,In_4893,In_2340);
nor U6140 (N_6140,In_4105,In_4325);
and U6141 (N_6141,In_3624,In_3360);
nor U6142 (N_6142,In_3243,In_626);
or U6143 (N_6143,In_3519,In_2999);
xnor U6144 (N_6144,In_25,In_524);
and U6145 (N_6145,In_45,In_123);
and U6146 (N_6146,In_1814,In_1350);
nor U6147 (N_6147,In_3248,In_4446);
nand U6148 (N_6148,In_1006,In_391);
xnor U6149 (N_6149,In_2411,In_2534);
nor U6150 (N_6150,In_3248,In_484);
and U6151 (N_6151,In_4031,In_1218);
and U6152 (N_6152,In_323,In_2493);
and U6153 (N_6153,In_471,In_608);
and U6154 (N_6154,In_1032,In_3172);
or U6155 (N_6155,In_3408,In_2287);
nor U6156 (N_6156,In_1098,In_160);
and U6157 (N_6157,In_604,In_2004);
nor U6158 (N_6158,In_4916,In_2060);
nand U6159 (N_6159,In_3236,In_593);
nand U6160 (N_6160,In_4147,In_774);
nand U6161 (N_6161,In_2114,In_4760);
or U6162 (N_6162,In_507,In_185);
or U6163 (N_6163,In_696,In_1346);
or U6164 (N_6164,In_4274,In_2073);
or U6165 (N_6165,In_2242,In_4832);
and U6166 (N_6166,In_3328,In_3519);
or U6167 (N_6167,In_2028,In_282);
nand U6168 (N_6168,In_3553,In_1911);
and U6169 (N_6169,In_646,In_1729);
nand U6170 (N_6170,In_3293,In_4002);
and U6171 (N_6171,In_2240,In_4506);
nor U6172 (N_6172,In_1495,In_4765);
and U6173 (N_6173,In_3985,In_4271);
xnor U6174 (N_6174,In_203,In_3668);
nor U6175 (N_6175,In_4968,In_1385);
nand U6176 (N_6176,In_1613,In_3942);
or U6177 (N_6177,In_2847,In_2092);
xnor U6178 (N_6178,In_2762,In_3721);
and U6179 (N_6179,In_4837,In_1467);
and U6180 (N_6180,In_321,In_3627);
nor U6181 (N_6181,In_4187,In_4173);
xnor U6182 (N_6182,In_3251,In_3152);
nor U6183 (N_6183,In_3610,In_4317);
xor U6184 (N_6184,In_792,In_2728);
xor U6185 (N_6185,In_392,In_2772);
nor U6186 (N_6186,In_4122,In_2288);
nand U6187 (N_6187,In_3405,In_2897);
xor U6188 (N_6188,In_2697,In_588);
nor U6189 (N_6189,In_4088,In_166);
nor U6190 (N_6190,In_2009,In_3538);
nor U6191 (N_6191,In_336,In_19);
nor U6192 (N_6192,In_135,In_803);
xor U6193 (N_6193,In_870,In_778);
nand U6194 (N_6194,In_1459,In_2283);
xor U6195 (N_6195,In_625,In_1080);
nand U6196 (N_6196,In_4310,In_2431);
nand U6197 (N_6197,In_4187,In_3739);
nand U6198 (N_6198,In_4886,In_4367);
nand U6199 (N_6199,In_935,In_201);
or U6200 (N_6200,In_940,In_3893);
nand U6201 (N_6201,In_3798,In_4668);
or U6202 (N_6202,In_1525,In_818);
nor U6203 (N_6203,In_1084,In_810);
or U6204 (N_6204,In_2804,In_2537);
nor U6205 (N_6205,In_2226,In_1287);
nand U6206 (N_6206,In_320,In_2359);
or U6207 (N_6207,In_3086,In_4895);
nand U6208 (N_6208,In_1924,In_3425);
nor U6209 (N_6209,In_1860,In_2363);
and U6210 (N_6210,In_3278,In_4950);
xnor U6211 (N_6211,In_1259,In_4551);
or U6212 (N_6212,In_542,In_386);
or U6213 (N_6213,In_2005,In_3010);
nor U6214 (N_6214,In_2829,In_2337);
and U6215 (N_6215,In_3902,In_1293);
or U6216 (N_6216,In_1649,In_4052);
xor U6217 (N_6217,In_258,In_3649);
or U6218 (N_6218,In_2449,In_496);
and U6219 (N_6219,In_553,In_3770);
nor U6220 (N_6220,In_641,In_2962);
and U6221 (N_6221,In_3331,In_1876);
or U6222 (N_6222,In_1275,In_3343);
nand U6223 (N_6223,In_4669,In_938);
and U6224 (N_6224,In_2622,In_3060);
xor U6225 (N_6225,In_665,In_2393);
nand U6226 (N_6226,In_4413,In_946);
or U6227 (N_6227,In_2418,In_2462);
nand U6228 (N_6228,In_4769,In_2671);
or U6229 (N_6229,In_1665,In_3953);
nor U6230 (N_6230,In_2929,In_2963);
xor U6231 (N_6231,In_2935,In_3493);
or U6232 (N_6232,In_3836,In_3239);
xor U6233 (N_6233,In_3510,In_1551);
xor U6234 (N_6234,In_2996,In_1405);
nor U6235 (N_6235,In_1347,In_4761);
nor U6236 (N_6236,In_828,In_3875);
xnor U6237 (N_6237,In_3591,In_995);
or U6238 (N_6238,In_2411,In_4922);
nor U6239 (N_6239,In_4378,In_227);
nand U6240 (N_6240,In_3932,In_3675);
nor U6241 (N_6241,In_4772,In_4075);
or U6242 (N_6242,In_1920,In_3764);
nand U6243 (N_6243,In_2833,In_1768);
and U6244 (N_6244,In_932,In_3656);
nor U6245 (N_6245,In_661,In_3805);
nand U6246 (N_6246,In_2845,In_172);
nor U6247 (N_6247,In_4612,In_627);
nand U6248 (N_6248,In_1461,In_2559);
nand U6249 (N_6249,In_4936,In_4368);
xor U6250 (N_6250,In_3342,In_4133);
xor U6251 (N_6251,In_4575,In_33);
xnor U6252 (N_6252,In_1858,In_4390);
xor U6253 (N_6253,In_1572,In_4293);
xor U6254 (N_6254,In_857,In_2916);
or U6255 (N_6255,In_4292,In_4230);
xnor U6256 (N_6256,In_881,In_738);
xnor U6257 (N_6257,In_1423,In_3499);
xor U6258 (N_6258,In_125,In_2385);
or U6259 (N_6259,In_4660,In_360);
or U6260 (N_6260,In_1318,In_1947);
or U6261 (N_6261,In_1060,In_2482);
nor U6262 (N_6262,In_388,In_1201);
xor U6263 (N_6263,In_335,In_2810);
and U6264 (N_6264,In_81,In_1655);
nand U6265 (N_6265,In_1039,In_1020);
nor U6266 (N_6266,In_2264,In_4391);
nor U6267 (N_6267,In_1795,In_4828);
nand U6268 (N_6268,In_1536,In_1431);
or U6269 (N_6269,In_3546,In_2587);
or U6270 (N_6270,In_1246,In_4706);
nand U6271 (N_6271,In_1575,In_1904);
nor U6272 (N_6272,In_40,In_3822);
nor U6273 (N_6273,In_4464,In_4412);
nand U6274 (N_6274,In_4199,In_1488);
nand U6275 (N_6275,In_2431,In_651);
nand U6276 (N_6276,In_3186,In_220);
nor U6277 (N_6277,In_3799,In_4249);
nand U6278 (N_6278,In_3426,In_580);
and U6279 (N_6279,In_2687,In_4985);
or U6280 (N_6280,In_1328,In_4816);
and U6281 (N_6281,In_3613,In_3140);
nand U6282 (N_6282,In_4699,In_1690);
nand U6283 (N_6283,In_4130,In_4670);
and U6284 (N_6284,In_2507,In_2755);
nand U6285 (N_6285,In_1288,In_215);
xnor U6286 (N_6286,In_4128,In_4765);
nand U6287 (N_6287,In_3783,In_4869);
nor U6288 (N_6288,In_3736,In_4544);
or U6289 (N_6289,In_3422,In_528);
and U6290 (N_6290,In_920,In_4243);
nand U6291 (N_6291,In_1838,In_745);
xor U6292 (N_6292,In_23,In_313);
nor U6293 (N_6293,In_1651,In_4463);
or U6294 (N_6294,In_2255,In_3382);
xnor U6295 (N_6295,In_2935,In_4494);
nor U6296 (N_6296,In_1545,In_1773);
and U6297 (N_6297,In_3312,In_3318);
xor U6298 (N_6298,In_4791,In_2484);
xor U6299 (N_6299,In_4610,In_2970);
and U6300 (N_6300,In_2305,In_4322);
nor U6301 (N_6301,In_1916,In_3520);
nand U6302 (N_6302,In_1492,In_4107);
and U6303 (N_6303,In_3740,In_1395);
nor U6304 (N_6304,In_3056,In_3947);
or U6305 (N_6305,In_3074,In_1391);
nand U6306 (N_6306,In_3001,In_3102);
nor U6307 (N_6307,In_2996,In_1698);
and U6308 (N_6308,In_3986,In_3098);
nand U6309 (N_6309,In_4499,In_2324);
xnor U6310 (N_6310,In_4547,In_426);
or U6311 (N_6311,In_4100,In_3412);
and U6312 (N_6312,In_2896,In_1983);
or U6313 (N_6313,In_2550,In_1518);
and U6314 (N_6314,In_555,In_419);
xnor U6315 (N_6315,In_2663,In_4134);
xnor U6316 (N_6316,In_3493,In_2283);
xor U6317 (N_6317,In_773,In_2346);
xnor U6318 (N_6318,In_2634,In_1247);
nor U6319 (N_6319,In_3784,In_1374);
and U6320 (N_6320,In_1457,In_4315);
or U6321 (N_6321,In_4585,In_52);
or U6322 (N_6322,In_2700,In_4532);
nand U6323 (N_6323,In_1824,In_3867);
nand U6324 (N_6324,In_4301,In_3075);
xor U6325 (N_6325,In_2643,In_1732);
nand U6326 (N_6326,In_3529,In_4202);
or U6327 (N_6327,In_2578,In_3263);
or U6328 (N_6328,In_4437,In_3422);
xor U6329 (N_6329,In_2727,In_1144);
nor U6330 (N_6330,In_2599,In_1723);
or U6331 (N_6331,In_3626,In_3811);
nand U6332 (N_6332,In_3482,In_748);
xnor U6333 (N_6333,In_3812,In_3649);
or U6334 (N_6334,In_4553,In_1003);
nor U6335 (N_6335,In_3516,In_300);
xor U6336 (N_6336,In_324,In_4497);
or U6337 (N_6337,In_269,In_3238);
xor U6338 (N_6338,In_876,In_4186);
or U6339 (N_6339,In_4254,In_4024);
and U6340 (N_6340,In_4708,In_1674);
or U6341 (N_6341,In_922,In_2230);
nand U6342 (N_6342,In_4832,In_1948);
nor U6343 (N_6343,In_4825,In_544);
xor U6344 (N_6344,In_1602,In_2872);
nand U6345 (N_6345,In_642,In_2027);
and U6346 (N_6346,In_1507,In_1137);
or U6347 (N_6347,In_3856,In_1992);
and U6348 (N_6348,In_4744,In_1282);
nor U6349 (N_6349,In_828,In_503);
or U6350 (N_6350,In_3084,In_14);
nor U6351 (N_6351,In_1286,In_474);
xnor U6352 (N_6352,In_1149,In_4418);
or U6353 (N_6353,In_1680,In_915);
xnor U6354 (N_6354,In_562,In_2912);
and U6355 (N_6355,In_136,In_1511);
and U6356 (N_6356,In_4036,In_4287);
xnor U6357 (N_6357,In_4949,In_3442);
nand U6358 (N_6358,In_1876,In_4011);
nand U6359 (N_6359,In_736,In_474);
or U6360 (N_6360,In_2173,In_2163);
nor U6361 (N_6361,In_279,In_435);
or U6362 (N_6362,In_231,In_4848);
nand U6363 (N_6363,In_3283,In_1285);
or U6364 (N_6364,In_4411,In_3075);
or U6365 (N_6365,In_440,In_3777);
or U6366 (N_6366,In_449,In_4983);
nor U6367 (N_6367,In_2802,In_3119);
or U6368 (N_6368,In_4006,In_1655);
nand U6369 (N_6369,In_2203,In_569);
or U6370 (N_6370,In_2098,In_1315);
nor U6371 (N_6371,In_4144,In_3600);
nor U6372 (N_6372,In_1881,In_4672);
nor U6373 (N_6373,In_4370,In_4264);
xor U6374 (N_6374,In_3180,In_1339);
nand U6375 (N_6375,In_274,In_3951);
nor U6376 (N_6376,In_3288,In_105);
xnor U6377 (N_6377,In_1510,In_3723);
nand U6378 (N_6378,In_2685,In_2189);
nor U6379 (N_6379,In_4266,In_1217);
and U6380 (N_6380,In_2195,In_967);
and U6381 (N_6381,In_4350,In_2615);
nor U6382 (N_6382,In_1182,In_3614);
or U6383 (N_6383,In_2372,In_2182);
nand U6384 (N_6384,In_979,In_613);
and U6385 (N_6385,In_2534,In_315);
and U6386 (N_6386,In_2009,In_2993);
nand U6387 (N_6387,In_1434,In_1962);
nor U6388 (N_6388,In_415,In_1594);
nor U6389 (N_6389,In_2164,In_4851);
xnor U6390 (N_6390,In_3020,In_4833);
and U6391 (N_6391,In_1519,In_490);
or U6392 (N_6392,In_907,In_2966);
nand U6393 (N_6393,In_3120,In_935);
nand U6394 (N_6394,In_2443,In_2424);
xor U6395 (N_6395,In_15,In_1363);
nand U6396 (N_6396,In_3577,In_3949);
or U6397 (N_6397,In_4795,In_428);
and U6398 (N_6398,In_166,In_4637);
nand U6399 (N_6399,In_1756,In_2988);
or U6400 (N_6400,In_1110,In_3722);
and U6401 (N_6401,In_1266,In_3010);
or U6402 (N_6402,In_3705,In_4808);
xnor U6403 (N_6403,In_4480,In_0);
xor U6404 (N_6404,In_2016,In_1996);
or U6405 (N_6405,In_599,In_1817);
xnor U6406 (N_6406,In_4422,In_873);
nand U6407 (N_6407,In_4568,In_1197);
nand U6408 (N_6408,In_2325,In_989);
or U6409 (N_6409,In_754,In_4491);
nor U6410 (N_6410,In_457,In_913);
xnor U6411 (N_6411,In_276,In_517);
and U6412 (N_6412,In_4235,In_1545);
nand U6413 (N_6413,In_1263,In_3101);
and U6414 (N_6414,In_1500,In_2298);
nor U6415 (N_6415,In_868,In_1271);
and U6416 (N_6416,In_4031,In_1159);
and U6417 (N_6417,In_4576,In_4813);
nand U6418 (N_6418,In_4220,In_3934);
nor U6419 (N_6419,In_3030,In_246);
and U6420 (N_6420,In_3203,In_710);
nor U6421 (N_6421,In_4688,In_2118);
nor U6422 (N_6422,In_1446,In_87);
or U6423 (N_6423,In_92,In_3215);
or U6424 (N_6424,In_3141,In_1858);
xnor U6425 (N_6425,In_4518,In_2490);
nand U6426 (N_6426,In_2078,In_2450);
xor U6427 (N_6427,In_2090,In_4686);
nand U6428 (N_6428,In_2155,In_3178);
and U6429 (N_6429,In_194,In_3962);
and U6430 (N_6430,In_730,In_579);
nand U6431 (N_6431,In_3136,In_423);
nand U6432 (N_6432,In_1471,In_3677);
and U6433 (N_6433,In_4966,In_1988);
and U6434 (N_6434,In_82,In_851);
and U6435 (N_6435,In_3737,In_4941);
xnor U6436 (N_6436,In_2363,In_2522);
or U6437 (N_6437,In_2648,In_3782);
nand U6438 (N_6438,In_606,In_2873);
nand U6439 (N_6439,In_3526,In_806);
nand U6440 (N_6440,In_3147,In_1519);
xnor U6441 (N_6441,In_3378,In_475);
xnor U6442 (N_6442,In_2900,In_252);
xor U6443 (N_6443,In_3901,In_2347);
xor U6444 (N_6444,In_4536,In_2028);
xor U6445 (N_6445,In_2956,In_4234);
and U6446 (N_6446,In_3440,In_600);
nor U6447 (N_6447,In_4994,In_4629);
nor U6448 (N_6448,In_4558,In_82);
nor U6449 (N_6449,In_3793,In_4266);
and U6450 (N_6450,In_3938,In_831);
and U6451 (N_6451,In_2409,In_1436);
and U6452 (N_6452,In_4572,In_2973);
nand U6453 (N_6453,In_3307,In_4090);
nor U6454 (N_6454,In_3313,In_4632);
and U6455 (N_6455,In_1136,In_4025);
and U6456 (N_6456,In_536,In_3540);
and U6457 (N_6457,In_2451,In_3743);
xnor U6458 (N_6458,In_1937,In_1569);
and U6459 (N_6459,In_1530,In_3517);
and U6460 (N_6460,In_4748,In_127);
and U6461 (N_6461,In_1659,In_676);
xor U6462 (N_6462,In_3796,In_229);
nand U6463 (N_6463,In_848,In_309);
nor U6464 (N_6464,In_1550,In_574);
nand U6465 (N_6465,In_3964,In_1117);
or U6466 (N_6466,In_749,In_1769);
and U6467 (N_6467,In_1242,In_120);
nor U6468 (N_6468,In_602,In_3394);
nand U6469 (N_6469,In_1250,In_2002);
nand U6470 (N_6470,In_374,In_2621);
nand U6471 (N_6471,In_3703,In_3103);
xor U6472 (N_6472,In_3686,In_1002);
xor U6473 (N_6473,In_1959,In_534);
xor U6474 (N_6474,In_4348,In_2121);
nand U6475 (N_6475,In_1047,In_3458);
nand U6476 (N_6476,In_2195,In_3372);
xor U6477 (N_6477,In_391,In_3655);
or U6478 (N_6478,In_3102,In_4527);
or U6479 (N_6479,In_3273,In_1595);
nand U6480 (N_6480,In_1979,In_3643);
and U6481 (N_6481,In_3092,In_1269);
xor U6482 (N_6482,In_663,In_2500);
xnor U6483 (N_6483,In_1877,In_2962);
and U6484 (N_6484,In_2671,In_4361);
and U6485 (N_6485,In_3769,In_927);
or U6486 (N_6486,In_1597,In_4133);
xor U6487 (N_6487,In_2109,In_2402);
nand U6488 (N_6488,In_1655,In_3797);
nand U6489 (N_6489,In_3134,In_2010);
xnor U6490 (N_6490,In_4925,In_2690);
nor U6491 (N_6491,In_3519,In_3638);
nor U6492 (N_6492,In_155,In_1685);
and U6493 (N_6493,In_4045,In_2529);
and U6494 (N_6494,In_902,In_3710);
and U6495 (N_6495,In_1877,In_3391);
xnor U6496 (N_6496,In_2080,In_1341);
or U6497 (N_6497,In_391,In_1414);
and U6498 (N_6498,In_323,In_2372);
and U6499 (N_6499,In_3770,In_27);
nand U6500 (N_6500,In_3678,In_3903);
or U6501 (N_6501,In_697,In_3944);
and U6502 (N_6502,In_2268,In_4090);
and U6503 (N_6503,In_2098,In_1267);
xnor U6504 (N_6504,In_1314,In_1568);
or U6505 (N_6505,In_4164,In_247);
and U6506 (N_6506,In_2742,In_1935);
nor U6507 (N_6507,In_363,In_4522);
nand U6508 (N_6508,In_115,In_4193);
and U6509 (N_6509,In_1114,In_2049);
and U6510 (N_6510,In_2350,In_4556);
nand U6511 (N_6511,In_2097,In_1103);
nand U6512 (N_6512,In_2341,In_2309);
xor U6513 (N_6513,In_80,In_1819);
xor U6514 (N_6514,In_1332,In_2318);
nand U6515 (N_6515,In_3677,In_1008);
nor U6516 (N_6516,In_4273,In_2496);
and U6517 (N_6517,In_3883,In_1236);
nand U6518 (N_6518,In_2966,In_3389);
nor U6519 (N_6519,In_405,In_695);
and U6520 (N_6520,In_3771,In_3221);
xor U6521 (N_6521,In_3501,In_3339);
nand U6522 (N_6522,In_3139,In_2725);
xnor U6523 (N_6523,In_4,In_178);
nor U6524 (N_6524,In_739,In_2879);
nor U6525 (N_6525,In_2845,In_1733);
or U6526 (N_6526,In_1119,In_3125);
xnor U6527 (N_6527,In_257,In_4312);
and U6528 (N_6528,In_2900,In_1209);
or U6529 (N_6529,In_4341,In_3207);
and U6530 (N_6530,In_2679,In_4210);
nand U6531 (N_6531,In_4663,In_4363);
nand U6532 (N_6532,In_4114,In_4940);
xor U6533 (N_6533,In_4929,In_1305);
or U6534 (N_6534,In_2862,In_3503);
and U6535 (N_6535,In_2513,In_3237);
nor U6536 (N_6536,In_445,In_4577);
nand U6537 (N_6537,In_1077,In_4073);
nand U6538 (N_6538,In_4080,In_1193);
and U6539 (N_6539,In_2778,In_3943);
xnor U6540 (N_6540,In_2507,In_4265);
nand U6541 (N_6541,In_742,In_2797);
nor U6542 (N_6542,In_3203,In_4586);
and U6543 (N_6543,In_4229,In_1715);
and U6544 (N_6544,In_3776,In_329);
nor U6545 (N_6545,In_990,In_795);
or U6546 (N_6546,In_3948,In_2600);
or U6547 (N_6547,In_3424,In_2214);
and U6548 (N_6548,In_2597,In_3817);
xnor U6549 (N_6549,In_2054,In_4285);
nor U6550 (N_6550,In_839,In_4644);
and U6551 (N_6551,In_4831,In_763);
xnor U6552 (N_6552,In_765,In_1063);
nand U6553 (N_6553,In_1852,In_1249);
or U6554 (N_6554,In_232,In_2570);
nor U6555 (N_6555,In_2015,In_2633);
nor U6556 (N_6556,In_3812,In_2340);
or U6557 (N_6557,In_332,In_2100);
and U6558 (N_6558,In_3080,In_3666);
and U6559 (N_6559,In_1662,In_794);
and U6560 (N_6560,In_2820,In_3687);
xor U6561 (N_6561,In_1974,In_2331);
nand U6562 (N_6562,In_2356,In_3800);
nor U6563 (N_6563,In_4798,In_1443);
xnor U6564 (N_6564,In_2778,In_3623);
nand U6565 (N_6565,In_743,In_1769);
or U6566 (N_6566,In_2531,In_106);
nand U6567 (N_6567,In_2946,In_1967);
and U6568 (N_6568,In_2705,In_3088);
or U6569 (N_6569,In_1794,In_2328);
and U6570 (N_6570,In_4887,In_3495);
and U6571 (N_6571,In_897,In_562);
or U6572 (N_6572,In_560,In_3678);
and U6573 (N_6573,In_1520,In_1911);
or U6574 (N_6574,In_352,In_3413);
and U6575 (N_6575,In_4744,In_4138);
xnor U6576 (N_6576,In_2108,In_2803);
nor U6577 (N_6577,In_4243,In_4080);
and U6578 (N_6578,In_2017,In_1353);
or U6579 (N_6579,In_2839,In_2223);
or U6580 (N_6580,In_4134,In_3516);
nor U6581 (N_6581,In_2219,In_3787);
and U6582 (N_6582,In_2027,In_2847);
nand U6583 (N_6583,In_556,In_1441);
or U6584 (N_6584,In_1120,In_1862);
nor U6585 (N_6585,In_2971,In_506);
nor U6586 (N_6586,In_437,In_312);
xor U6587 (N_6587,In_2350,In_3399);
or U6588 (N_6588,In_1970,In_4306);
nor U6589 (N_6589,In_3251,In_1489);
xor U6590 (N_6590,In_1578,In_4284);
nor U6591 (N_6591,In_4897,In_2866);
and U6592 (N_6592,In_3585,In_2502);
nand U6593 (N_6593,In_3507,In_915);
xnor U6594 (N_6594,In_595,In_754);
xnor U6595 (N_6595,In_4742,In_1477);
and U6596 (N_6596,In_4879,In_485);
or U6597 (N_6597,In_2170,In_4937);
nor U6598 (N_6598,In_2777,In_2499);
and U6599 (N_6599,In_1622,In_4084);
or U6600 (N_6600,In_280,In_4678);
and U6601 (N_6601,In_716,In_1934);
nand U6602 (N_6602,In_4067,In_4534);
nand U6603 (N_6603,In_4074,In_2530);
nand U6604 (N_6604,In_4497,In_4816);
xnor U6605 (N_6605,In_1774,In_4241);
xnor U6606 (N_6606,In_582,In_4851);
nor U6607 (N_6607,In_771,In_12);
or U6608 (N_6608,In_2694,In_1233);
or U6609 (N_6609,In_4552,In_4407);
nor U6610 (N_6610,In_260,In_2989);
nand U6611 (N_6611,In_2077,In_4047);
xnor U6612 (N_6612,In_3345,In_3302);
nor U6613 (N_6613,In_107,In_1054);
nor U6614 (N_6614,In_2323,In_4523);
and U6615 (N_6615,In_4492,In_364);
and U6616 (N_6616,In_3581,In_4072);
and U6617 (N_6617,In_3230,In_4245);
nor U6618 (N_6618,In_4229,In_4848);
and U6619 (N_6619,In_646,In_2052);
nor U6620 (N_6620,In_1478,In_2793);
xnor U6621 (N_6621,In_1400,In_592);
nand U6622 (N_6622,In_645,In_516);
nand U6623 (N_6623,In_3198,In_3947);
xor U6624 (N_6624,In_4649,In_3136);
and U6625 (N_6625,In_1693,In_3375);
or U6626 (N_6626,In_3711,In_4280);
xor U6627 (N_6627,In_4931,In_856);
and U6628 (N_6628,In_1326,In_434);
xnor U6629 (N_6629,In_10,In_2311);
xor U6630 (N_6630,In_4842,In_4937);
nand U6631 (N_6631,In_4642,In_1938);
xnor U6632 (N_6632,In_891,In_3181);
and U6633 (N_6633,In_1572,In_4881);
xor U6634 (N_6634,In_2811,In_2341);
and U6635 (N_6635,In_2767,In_2725);
or U6636 (N_6636,In_4991,In_747);
xnor U6637 (N_6637,In_4991,In_2114);
xor U6638 (N_6638,In_3683,In_4647);
and U6639 (N_6639,In_4217,In_3838);
nand U6640 (N_6640,In_2358,In_1922);
nand U6641 (N_6641,In_4589,In_4650);
xor U6642 (N_6642,In_3999,In_3951);
xor U6643 (N_6643,In_1481,In_572);
and U6644 (N_6644,In_1843,In_4325);
and U6645 (N_6645,In_571,In_4741);
or U6646 (N_6646,In_4376,In_3671);
and U6647 (N_6647,In_3192,In_1469);
or U6648 (N_6648,In_599,In_306);
nand U6649 (N_6649,In_4385,In_3820);
and U6650 (N_6650,In_3925,In_2034);
or U6651 (N_6651,In_3371,In_3996);
nor U6652 (N_6652,In_3585,In_2205);
or U6653 (N_6653,In_294,In_2159);
and U6654 (N_6654,In_2172,In_577);
nor U6655 (N_6655,In_4032,In_4572);
and U6656 (N_6656,In_3979,In_2576);
nand U6657 (N_6657,In_1653,In_4747);
or U6658 (N_6658,In_361,In_1060);
xnor U6659 (N_6659,In_3059,In_4915);
xor U6660 (N_6660,In_2571,In_950);
and U6661 (N_6661,In_4599,In_2969);
nand U6662 (N_6662,In_1468,In_4602);
and U6663 (N_6663,In_4953,In_2713);
and U6664 (N_6664,In_1901,In_27);
nor U6665 (N_6665,In_1490,In_369);
xnor U6666 (N_6666,In_164,In_1202);
or U6667 (N_6667,In_2866,In_390);
nor U6668 (N_6668,In_1467,In_1249);
nor U6669 (N_6669,In_2820,In_2665);
xor U6670 (N_6670,In_2806,In_1618);
nor U6671 (N_6671,In_2731,In_4634);
xnor U6672 (N_6672,In_190,In_1829);
nor U6673 (N_6673,In_2151,In_669);
and U6674 (N_6674,In_2454,In_727);
or U6675 (N_6675,In_1712,In_12);
nor U6676 (N_6676,In_465,In_1008);
nor U6677 (N_6677,In_109,In_1560);
nand U6678 (N_6678,In_2888,In_4629);
nand U6679 (N_6679,In_2762,In_884);
or U6680 (N_6680,In_1877,In_3014);
and U6681 (N_6681,In_2956,In_2360);
nor U6682 (N_6682,In_3225,In_4844);
nand U6683 (N_6683,In_1190,In_3006);
nand U6684 (N_6684,In_3155,In_2029);
or U6685 (N_6685,In_193,In_55);
nor U6686 (N_6686,In_1404,In_2718);
or U6687 (N_6687,In_4794,In_404);
or U6688 (N_6688,In_2550,In_3801);
xor U6689 (N_6689,In_2277,In_3233);
nand U6690 (N_6690,In_1978,In_3168);
or U6691 (N_6691,In_143,In_2031);
xnor U6692 (N_6692,In_4371,In_3023);
nand U6693 (N_6693,In_923,In_2490);
and U6694 (N_6694,In_1753,In_1165);
or U6695 (N_6695,In_3231,In_613);
xnor U6696 (N_6696,In_2554,In_246);
nor U6697 (N_6697,In_165,In_1698);
nor U6698 (N_6698,In_2137,In_716);
nor U6699 (N_6699,In_1767,In_1582);
nand U6700 (N_6700,In_3041,In_273);
and U6701 (N_6701,In_4182,In_3254);
xnor U6702 (N_6702,In_3989,In_4477);
nand U6703 (N_6703,In_2067,In_143);
or U6704 (N_6704,In_2310,In_878);
and U6705 (N_6705,In_2182,In_2686);
nand U6706 (N_6706,In_4338,In_171);
nor U6707 (N_6707,In_2218,In_4101);
nand U6708 (N_6708,In_462,In_2214);
nand U6709 (N_6709,In_3241,In_3119);
xnor U6710 (N_6710,In_3736,In_935);
and U6711 (N_6711,In_2058,In_615);
nand U6712 (N_6712,In_224,In_3455);
nand U6713 (N_6713,In_280,In_3311);
and U6714 (N_6714,In_3615,In_1284);
nor U6715 (N_6715,In_174,In_492);
and U6716 (N_6716,In_2920,In_844);
or U6717 (N_6717,In_582,In_484);
and U6718 (N_6718,In_3639,In_2650);
nor U6719 (N_6719,In_4077,In_1629);
xnor U6720 (N_6720,In_3489,In_1876);
nand U6721 (N_6721,In_4741,In_1042);
nor U6722 (N_6722,In_2162,In_3617);
nand U6723 (N_6723,In_1451,In_1251);
xnor U6724 (N_6724,In_2803,In_941);
xor U6725 (N_6725,In_2503,In_4309);
nor U6726 (N_6726,In_1448,In_1853);
and U6727 (N_6727,In_4904,In_3929);
or U6728 (N_6728,In_4152,In_1445);
xor U6729 (N_6729,In_38,In_3695);
nor U6730 (N_6730,In_3060,In_4529);
nand U6731 (N_6731,In_1397,In_851);
nor U6732 (N_6732,In_3961,In_2888);
nand U6733 (N_6733,In_618,In_2711);
and U6734 (N_6734,In_28,In_1574);
xor U6735 (N_6735,In_3713,In_3431);
xor U6736 (N_6736,In_2435,In_2340);
nand U6737 (N_6737,In_3630,In_1728);
nand U6738 (N_6738,In_4369,In_1331);
nor U6739 (N_6739,In_785,In_1306);
or U6740 (N_6740,In_4417,In_4882);
xor U6741 (N_6741,In_4821,In_958);
or U6742 (N_6742,In_2206,In_4180);
nor U6743 (N_6743,In_3687,In_420);
or U6744 (N_6744,In_1697,In_2831);
nand U6745 (N_6745,In_4497,In_3435);
and U6746 (N_6746,In_1637,In_469);
nand U6747 (N_6747,In_829,In_2946);
nor U6748 (N_6748,In_214,In_4446);
nand U6749 (N_6749,In_3573,In_514);
or U6750 (N_6750,In_698,In_260);
nand U6751 (N_6751,In_3407,In_3413);
nand U6752 (N_6752,In_2775,In_3704);
nand U6753 (N_6753,In_3713,In_1965);
nor U6754 (N_6754,In_4422,In_4073);
nand U6755 (N_6755,In_4118,In_3011);
nand U6756 (N_6756,In_2165,In_1616);
or U6757 (N_6757,In_4104,In_2621);
xor U6758 (N_6758,In_47,In_1524);
xnor U6759 (N_6759,In_4859,In_4632);
xnor U6760 (N_6760,In_3865,In_4683);
or U6761 (N_6761,In_2169,In_1627);
or U6762 (N_6762,In_2617,In_3891);
nor U6763 (N_6763,In_2346,In_3571);
or U6764 (N_6764,In_3778,In_2469);
xnor U6765 (N_6765,In_2175,In_1938);
nor U6766 (N_6766,In_1918,In_1048);
and U6767 (N_6767,In_2548,In_3607);
nor U6768 (N_6768,In_3518,In_2816);
xor U6769 (N_6769,In_4576,In_3648);
and U6770 (N_6770,In_2900,In_1387);
and U6771 (N_6771,In_3128,In_1569);
nor U6772 (N_6772,In_4694,In_2027);
and U6773 (N_6773,In_3196,In_1762);
and U6774 (N_6774,In_246,In_2380);
xor U6775 (N_6775,In_968,In_4767);
xnor U6776 (N_6776,In_3052,In_1247);
nand U6777 (N_6777,In_637,In_3704);
or U6778 (N_6778,In_4906,In_2292);
nor U6779 (N_6779,In_1407,In_1235);
nor U6780 (N_6780,In_2199,In_472);
nor U6781 (N_6781,In_4702,In_1152);
or U6782 (N_6782,In_4931,In_2444);
xor U6783 (N_6783,In_1422,In_3870);
xor U6784 (N_6784,In_4432,In_4749);
nor U6785 (N_6785,In_3136,In_2493);
xnor U6786 (N_6786,In_955,In_4330);
xor U6787 (N_6787,In_3757,In_4100);
xnor U6788 (N_6788,In_586,In_4222);
xor U6789 (N_6789,In_4096,In_4825);
nand U6790 (N_6790,In_3511,In_846);
nand U6791 (N_6791,In_4548,In_1094);
or U6792 (N_6792,In_2618,In_2836);
and U6793 (N_6793,In_953,In_4057);
nor U6794 (N_6794,In_3610,In_3499);
nor U6795 (N_6795,In_2382,In_3730);
or U6796 (N_6796,In_987,In_1183);
nor U6797 (N_6797,In_972,In_223);
nand U6798 (N_6798,In_4350,In_2338);
and U6799 (N_6799,In_2920,In_339);
nand U6800 (N_6800,In_989,In_2973);
and U6801 (N_6801,In_4170,In_551);
or U6802 (N_6802,In_4589,In_2377);
nand U6803 (N_6803,In_3229,In_1579);
or U6804 (N_6804,In_4983,In_3328);
xor U6805 (N_6805,In_2255,In_3264);
or U6806 (N_6806,In_2340,In_1129);
nor U6807 (N_6807,In_1299,In_2490);
nand U6808 (N_6808,In_2471,In_2739);
or U6809 (N_6809,In_2713,In_1851);
or U6810 (N_6810,In_1433,In_3302);
nor U6811 (N_6811,In_2313,In_43);
nand U6812 (N_6812,In_2729,In_1123);
nor U6813 (N_6813,In_236,In_2587);
or U6814 (N_6814,In_4324,In_429);
nand U6815 (N_6815,In_2096,In_1639);
nand U6816 (N_6816,In_2090,In_2103);
and U6817 (N_6817,In_3593,In_1458);
nand U6818 (N_6818,In_3416,In_2709);
and U6819 (N_6819,In_3588,In_222);
and U6820 (N_6820,In_1556,In_943);
nand U6821 (N_6821,In_3637,In_4053);
xor U6822 (N_6822,In_1883,In_2944);
and U6823 (N_6823,In_2516,In_204);
xnor U6824 (N_6824,In_4576,In_4982);
nor U6825 (N_6825,In_4946,In_3008);
or U6826 (N_6826,In_3112,In_1435);
nand U6827 (N_6827,In_2642,In_854);
nand U6828 (N_6828,In_4379,In_1045);
nand U6829 (N_6829,In_1564,In_3707);
xnor U6830 (N_6830,In_4735,In_3116);
nand U6831 (N_6831,In_4302,In_4152);
nand U6832 (N_6832,In_3045,In_4873);
and U6833 (N_6833,In_2413,In_4880);
nand U6834 (N_6834,In_4063,In_2155);
and U6835 (N_6835,In_2296,In_1617);
and U6836 (N_6836,In_3291,In_1052);
xnor U6837 (N_6837,In_252,In_907);
or U6838 (N_6838,In_3852,In_1510);
or U6839 (N_6839,In_1860,In_1881);
and U6840 (N_6840,In_654,In_3202);
nand U6841 (N_6841,In_4690,In_4812);
nand U6842 (N_6842,In_2514,In_2174);
or U6843 (N_6843,In_2170,In_2212);
or U6844 (N_6844,In_4518,In_3088);
and U6845 (N_6845,In_2277,In_1212);
or U6846 (N_6846,In_4432,In_1870);
xor U6847 (N_6847,In_1208,In_836);
xnor U6848 (N_6848,In_1941,In_910);
and U6849 (N_6849,In_3936,In_4005);
nor U6850 (N_6850,In_3508,In_3964);
and U6851 (N_6851,In_175,In_2568);
and U6852 (N_6852,In_2772,In_3287);
xnor U6853 (N_6853,In_706,In_472);
and U6854 (N_6854,In_1758,In_3326);
nand U6855 (N_6855,In_370,In_2020);
nor U6856 (N_6856,In_2085,In_1414);
nor U6857 (N_6857,In_891,In_1008);
nor U6858 (N_6858,In_4270,In_4066);
nand U6859 (N_6859,In_910,In_4066);
nor U6860 (N_6860,In_4238,In_874);
xnor U6861 (N_6861,In_4412,In_1584);
xnor U6862 (N_6862,In_1916,In_3368);
nor U6863 (N_6863,In_818,In_4417);
or U6864 (N_6864,In_3537,In_2605);
nand U6865 (N_6865,In_223,In_3053);
or U6866 (N_6866,In_1925,In_891);
nor U6867 (N_6867,In_3849,In_2084);
or U6868 (N_6868,In_4090,In_3251);
or U6869 (N_6869,In_4001,In_930);
or U6870 (N_6870,In_3280,In_1009);
or U6871 (N_6871,In_3142,In_4637);
and U6872 (N_6872,In_1389,In_4020);
xor U6873 (N_6873,In_4207,In_4547);
and U6874 (N_6874,In_1361,In_1164);
and U6875 (N_6875,In_966,In_1812);
nand U6876 (N_6876,In_2886,In_2359);
or U6877 (N_6877,In_2443,In_1210);
or U6878 (N_6878,In_2936,In_4447);
nor U6879 (N_6879,In_764,In_1829);
xnor U6880 (N_6880,In_2509,In_746);
xnor U6881 (N_6881,In_939,In_1928);
and U6882 (N_6882,In_2796,In_3531);
and U6883 (N_6883,In_3709,In_32);
or U6884 (N_6884,In_951,In_2470);
xnor U6885 (N_6885,In_661,In_4346);
nand U6886 (N_6886,In_4139,In_1179);
xnor U6887 (N_6887,In_4879,In_2506);
nand U6888 (N_6888,In_833,In_1450);
or U6889 (N_6889,In_3601,In_3683);
nor U6890 (N_6890,In_258,In_4317);
nand U6891 (N_6891,In_4216,In_1308);
or U6892 (N_6892,In_723,In_1863);
nor U6893 (N_6893,In_3566,In_1045);
xor U6894 (N_6894,In_3038,In_1263);
nor U6895 (N_6895,In_2488,In_784);
or U6896 (N_6896,In_4304,In_1434);
nor U6897 (N_6897,In_3656,In_893);
nand U6898 (N_6898,In_546,In_2859);
nand U6899 (N_6899,In_2584,In_3585);
xnor U6900 (N_6900,In_1988,In_4143);
nor U6901 (N_6901,In_2444,In_4728);
xnor U6902 (N_6902,In_2052,In_354);
nor U6903 (N_6903,In_1063,In_2284);
or U6904 (N_6904,In_1945,In_3167);
nand U6905 (N_6905,In_4979,In_2802);
nor U6906 (N_6906,In_1017,In_3464);
or U6907 (N_6907,In_1550,In_3122);
and U6908 (N_6908,In_4862,In_3301);
or U6909 (N_6909,In_1996,In_2469);
nor U6910 (N_6910,In_3425,In_1126);
xor U6911 (N_6911,In_2455,In_3250);
xor U6912 (N_6912,In_2713,In_2439);
and U6913 (N_6913,In_1024,In_1580);
and U6914 (N_6914,In_4883,In_4618);
and U6915 (N_6915,In_2837,In_1930);
nor U6916 (N_6916,In_840,In_395);
nor U6917 (N_6917,In_1006,In_485);
and U6918 (N_6918,In_615,In_2817);
or U6919 (N_6919,In_3607,In_1994);
nor U6920 (N_6920,In_1841,In_446);
nand U6921 (N_6921,In_1480,In_4);
xor U6922 (N_6922,In_120,In_4783);
or U6923 (N_6923,In_4705,In_2305);
nor U6924 (N_6924,In_3928,In_4172);
nand U6925 (N_6925,In_1343,In_3715);
nor U6926 (N_6926,In_2057,In_2000);
nand U6927 (N_6927,In_4358,In_3750);
nand U6928 (N_6928,In_1536,In_3251);
or U6929 (N_6929,In_4759,In_3766);
xnor U6930 (N_6930,In_1728,In_3647);
and U6931 (N_6931,In_4861,In_92);
nand U6932 (N_6932,In_2624,In_2584);
or U6933 (N_6933,In_4787,In_2135);
nor U6934 (N_6934,In_470,In_3660);
nand U6935 (N_6935,In_2543,In_4029);
nor U6936 (N_6936,In_2963,In_2063);
nand U6937 (N_6937,In_298,In_377);
or U6938 (N_6938,In_4378,In_2253);
nand U6939 (N_6939,In_779,In_4421);
nor U6940 (N_6940,In_2291,In_824);
or U6941 (N_6941,In_1526,In_329);
nor U6942 (N_6942,In_4636,In_2248);
or U6943 (N_6943,In_4479,In_2171);
xor U6944 (N_6944,In_3365,In_1393);
or U6945 (N_6945,In_4580,In_1849);
or U6946 (N_6946,In_3890,In_464);
or U6947 (N_6947,In_3588,In_4317);
xor U6948 (N_6948,In_794,In_3437);
nor U6949 (N_6949,In_1006,In_4689);
nor U6950 (N_6950,In_4565,In_423);
and U6951 (N_6951,In_686,In_4363);
nor U6952 (N_6952,In_3461,In_611);
nor U6953 (N_6953,In_4645,In_2460);
nor U6954 (N_6954,In_4694,In_2784);
nand U6955 (N_6955,In_1087,In_4958);
nor U6956 (N_6956,In_3850,In_2593);
nand U6957 (N_6957,In_3682,In_4082);
or U6958 (N_6958,In_1804,In_4901);
nor U6959 (N_6959,In_2263,In_1853);
xnor U6960 (N_6960,In_2449,In_3283);
nor U6961 (N_6961,In_3814,In_1200);
or U6962 (N_6962,In_603,In_1055);
nand U6963 (N_6963,In_4606,In_1695);
or U6964 (N_6964,In_2162,In_1690);
xnor U6965 (N_6965,In_3044,In_310);
nor U6966 (N_6966,In_3266,In_1035);
or U6967 (N_6967,In_4225,In_1541);
nand U6968 (N_6968,In_814,In_4988);
and U6969 (N_6969,In_565,In_2233);
xor U6970 (N_6970,In_4294,In_4816);
xnor U6971 (N_6971,In_2398,In_4297);
nor U6972 (N_6972,In_2997,In_4961);
or U6973 (N_6973,In_3010,In_4430);
xor U6974 (N_6974,In_1009,In_4242);
or U6975 (N_6975,In_3721,In_272);
and U6976 (N_6976,In_4232,In_2969);
nand U6977 (N_6977,In_1192,In_2323);
nand U6978 (N_6978,In_2883,In_17);
xor U6979 (N_6979,In_4446,In_3362);
or U6980 (N_6980,In_1187,In_453);
nand U6981 (N_6981,In_3666,In_1320);
and U6982 (N_6982,In_3768,In_3076);
nor U6983 (N_6983,In_4975,In_128);
nand U6984 (N_6984,In_4864,In_4939);
xnor U6985 (N_6985,In_3703,In_1039);
and U6986 (N_6986,In_1681,In_190);
and U6987 (N_6987,In_2013,In_1996);
and U6988 (N_6988,In_4989,In_3905);
nor U6989 (N_6989,In_2022,In_3220);
nand U6990 (N_6990,In_2072,In_3165);
or U6991 (N_6991,In_2524,In_4247);
and U6992 (N_6992,In_1080,In_4371);
nor U6993 (N_6993,In_715,In_2416);
and U6994 (N_6994,In_2608,In_4783);
nor U6995 (N_6995,In_2414,In_3276);
or U6996 (N_6996,In_3640,In_975);
or U6997 (N_6997,In_3412,In_4946);
xor U6998 (N_6998,In_39,In_2364);
and U6999 (N_6999,In_4076,In_3394);
or U7000 (N_7000,In_2808,In_3347);
or U7001 (N_7001,In_4083,In_2467);
nand U7002 (N_7002,In_85,In_4568);
nand U7003 (N_7003,In_399,In_535);
and U7004 (N_7004,In_3287,In_2795);
nor U7005 (N_7005,In_60,In_2876);
and U7006 (N_7006,In_1909,In_3608);
nand U7007 (N_7007,In_199,In_3097);
xnor U7008 (N_7008,In_3203,In_1083);
nand U7009 (N_7009,In_4602,In_3774);
nand U7010 (N_7010,In_789,In_2869);
nand U7011 (N_7011,In_497,In_1931);
nand U7012 (N_7012,In_3213,In_824);
nor U7013 (N_7013,In_4514,In_3290);
and U7014 (N_7014,In_4781,In_782);
xor U7015 (N_7015,In_2141,In_3818);
and U7016 (N_7016,In_3963,In_1882);
and U7017 (N_7017,In_1993,In_4865);
and U7018 (N_7018,In_2649,In_3155);
and U7019 (N_7019,In_2910,In_3131);
xor U7020 (N_7020,In_465,In_2969);
or U7021 (N_7021,In_1322,In_303);
and U7022 (N_7022,In_1838,In_1609);
or U7023 (N_7023,In_1683,In_1182);
nor U7024 (N_7024,In_3047,In_3014);
xnor U7025 (N_7025,In_646,In_3445);
and U7026 (N_7026,In_2005,In_1685);
nor U7027 (N_7027,In_4657,In_2911);
xor U7028 (N_7028,In_1579,In_4362);
nor U7029 (N_7029,In_2422,In_572);
and U7030 (N_7030,In_4275,In_2740);
or U7031 (N_7031,In_4415,In_4314);
or U7032 (N_7032,In_3115,In_2388);
or U7033 (N_7033,In_2079,In_3821);
nor U7034 (N_7034,In_3186,In_4341);
xnor U7035 (N_7035,In_4234,In_4983);
nand U7036 (N_7036,In_2768,In_2140);
nor U7037 (N_7037,In_4800,In_3597);
nand U7038 (N_7038,In_1550,In_4080);
xnor U7039 (N_7039,In_1958,In_2822);
or U7040 (N_7040,In_572,In_3876);
nand U7041 (N_7041,In_1192,In_2139);
or U7042 (N_7042,In_2467,In_1187);
and U7043 (N_7043,In_4628,In_516);
and U7044 (N_7044,In_2029,In_458);
and U7045 (N_7045,In_1669,In_2598);
or U7046 (N_7046,In_225,In_1512);
xor U7047 (N_7047,In_4527,In_1729);
nor U7048 (N_7048,In_437,In_787);
nand U7049 (N_7049,In_3146,In_508);
nor U7050 (N_7050,In_4319,In_3760);
and U7051 (N_7051,In_594,In_2546);
and U7052 (N_7052,In_2936,In_35);
nor U7053 (N_7053,In_2737,In_4322);
nand U7054 (N_7054,In_4109,In_2399);
xor U7055 (N_7055,In_3121,In_4355);
nand U7056 (N_7056,In_1401,In_478);
nand U7057 (N_7057,In_633,In_1507);
xor U7058 (N_7058,In_3723,In_1776);
and U7059 (N_7059,In_4450,In_1369);
and U7060 (N_7060,In_998,In_4611);
xnor U7061 (N_7061,In_3725,In_2886);
nor U7062 (N_7062,In_3302,In_264);
or U7063 (N_7063,In_2608,In_4162);
nor U7064 (N_7064,In_3435,In_468);
nor U7065 (N_7065,In_1279,In_706);
nand U7066 (N_7066,In_199,In_1827);
nor U7067 (N_7067,In_734,In_4478);
nor U7068 (N_7068,In_2429,In_3582);
or U7069 (N_7069,In_3866,In_144);
nand U7070 (N_7070,In_226,In_2617);
and U7071 (N_7071,In_1114,In_17);
nand U7072 (N_7072,In_2711,In_2331);
and U7073 (N_7073,In_2194,In_3214);
nor U7074 (N_7074,In_1213,In_4228);
or U7075 (N_7075,In_4226,In_4496);
nor U7076 (N_7076,In_3886,In_3524);
and U7077 (N_7077,In_3794,In_951);
nand U7078 (N_7078,In_4053,In_2255);
nor U7079 (N_7079,In_4948,In_584);
and U7080 (N_7080,In_4232,In_2645);
nand U7081 (N_7081,In_1545,In_1168);
and U7082 (N_7082,In_377,In_4351);
nand U7083 (N_7083,In_455,In_3968);
nand U7084 (N_7084,In_1389,In_3605);
and U7085 (N_7085,In_4196,In_179);
and U7086 (N_7086,In_3479,In_3894);
or U7087 (N_7087,In_3394,In_4538);
or U7088 (N_7088,In_3451,In_2040);
xnor U7089 (N_7089,In_3481,In_4423);
or U7090 (N_7090,In_3899,In_3301);
nor U7091 (N_7091,In_3095,In_2996);
and U7092 (N_7092,In_2307,In_3900);
nand U7093 (N_7093,In_236,In_4115);
xnor U7094 (N_7094,In_4330,In_3862);
nand U7095 (N_7095,In_724,In_881);
xnor U7096 (N_7096,In_2832,In_3502);
nand U7097 (N_7097,In_2171,In_3248);
xnor U7098 (N_7098,In_3322,In_2663);
xnor U7099 (N_7099,In_3952,In_50);
nor U7100 (N_7100,In_181,In_3393);
and U7101 (N_7101,In_4172,In_3000);
nand U7102 (N_7102,In_3796,In_1735);
nor U7103 (N_7103,In_111,In_377);
and U7104 (N_7104,In_4029,In_2934);
and U7105 (N_7105,In_1911,In_4601);
nor U7106 (N_7106,In_3370,In_1315);
nor U7107 (N_7107,In_4139,In_3573);
or U7108 (N_7108,In_4095,In_2726);
or U7109 (N_7109,In_2267,In_593);
and U7110 (N_7110,In_625,In_3484);
and U7111 (N_7111,In_2183,In_3414);
nand U7112 (N_7112,In_3374,In_4534);
nand U7113 (N_7113,In_3087,In_137);
and U7114 (N_7114,In_4769,In_2347);
and U7115 (N_7115,In_728,In_3078);
and U7116 (N_7116,In_1827,In_3368);
or U7117 (N_7117,In_902,In_448);
or U7118 (N_7118,In_187,In_3086);
nor U7119 (N_7119,In_1540,In_4985);
xor U7120 (N_7120,In_3035,In_2755);
xnor U7121 (N_7121,In_4230,In_3149);
or U7122 (N_7122,In_2208,In_332);
nor U7123 (N_7123,In_2207,In_2168);
or U7124 (N_7124,In_483,In_4207);
or U7125 (N_7125,In_2490,In_3752);
nand U7126 (N_7126,In_1633,In_3711);
or U7127 (N_7127,In_93,In_999);
or U7128 (N_7128,In_4169,In_3924);
xnor U7129 (N_7129,In_1331,In_1790);
nand U7130 (N_7130,In_3245,In_2869);
nand U7131 (N_7131,In_4921,In_533);
nor U7132 (N_7132,In_115,In_4900);
or U7133 (N_7133,In_2023,In_1830);
nand U7134 (N_7134,In_3017,In_1989);
nand U7135 (N_7135,In_2805,In_15);
nand U7136 (N_7136,In_525,In_2893);
or U7137 (N_7137,In_2714,In_237);
or U7138 (N_7138,In_2304,In_3425);
and U7139 (N_7139,In_2114,In_3222);
or U7140 (N_7140,In_4278,In_32);
nand U7141 (N_7141,In_779,In_3617);
nand U7142 (N_7142,In_1131,In_2046);
nor U7143 (N_7143,In_568,In_1201);
or U7144 (N_7144,In_2502,In_1860);
xor U7145 (N_7145,In_1570,In_3583);
nor U7146 (N_7146,In_1025,In_3093);
or U7147 (N_7147,In_2411,In_2671);
xnor U7148 (N_7148,In_1500,In_3955);
nand U7149 (N_7149,In_3019,In_1640);
nand U7150 (N_7150,In_1554,In_1532);
nand U7151 (N_7151,In_4446,In_300);
or U7152 (N_7152,In_4837,In_534);
nand U7153 (N_7153,In_476,In_4815);
nor U7154 (N_7154,In_425,In_4067);
xor U7155 (N_7155,In_3414,In_262);
xnor U7156 (N_7156,In_4865,In_4905);
xnor U7157 (N_7157,In_1212,In_4610);
nor U7158 (N_7158,In_1029,In_3930);
xnor U7159 (N_7159,In_300,In_1914);
nor U7160 (N_7160,In_574,In_3507);
xnor U7161 (N_7161,In_687,In_4084);
nor U7162 (N_7162,In_3656,In_1863);
nand U7163 (N_7163,In_4376,In_3586);
and U7164 (N_7164,In_2703,In_2775);
nand U7165 (N_7165,In_1864,In_3498);
xnor U7166 (N_7166,In_2520,In_1288);
nor U7167 (N_7167,In_1003,In_2188);
and U7168 (N_7168,In_4682,In_4069);
and U7169 (N_7169,In_3102,In_3029);
nand U7170 (N_7170,In_44,In_3888);
nand U7171 (N_7171,In_202,In_1167);
and U7172 (N_7172,In_3032,In_4546);
nand U7173 (N_7173,In_1289,In_459);
and U7174 (N_7174,In_4188,In_2026);
nand U7175 (N_7175,In_4585,In_4147);
nand U7176 (N_7176,In_3716,In_1789);
and U7177 (N_7177,In_1831,In_2237);
and U7178 (N_7178,In_4943,In_1468);
nor U7179 (N_7179,In_4222,In_3381);
and U7180 (N_7180,In_1242,In_1946);
nand U7181 (N_7181,In_1797,In_1380);
or U7182 (N_7182,In_2046,In_4162);
xnor U7183 (N_7183,In_2321,In_347);
and U7184 (N_7184,In_24,In_1368);
or U7185 (N_7185,In_1243,In_214);
and U7186 (N_7186,In_3132,In_1151);
nand U7187 (N_7187,In_2151,In_277);
xor U7188 (N_7188,In_1288,In_2435);
nor U7189 (N_7189,In_4773,In_697);
xor U7190 (N_7190,In_2991,In_1889);
and U7191 (N_7191,In_2749,In_894);
or U7192 (N_7192,In_3836,In_40);
nor U7193 (N_7193,In_1748,In_2847);
or U7194 (N_7194,In_1655,In_1548);
nor U7195 (N_7195,In_2232,In_3860);
nor U7196 (N_7196,In_1587,In_4997);
or U7197 (N_7197,In_543,In_3683);
nor U7198 (N_7198,In_135,In_4584);
and U7199 (N_7199,In_1786,In_3996);
nor U7200 (N_7200,In_3356,In_1979);
xnor U7201 (N_7201,In_2272,In_2196);
and U7202 (N_7202,In_2219,In_825);
nor U7203 (N_7203,In_1846,In_3357);
nand U7204 (N_7204,In_1076,In_4598);
or U7205 (N_7205,In_4528,In_3014);
xnor U7206 (N_7206,In_2556,In_4821);
xor U7207 (N_7207,In_2055,In_1357);
and U7208 (N_7208,In_3603,In_69);
xnor U7209 (N_7209,In_82,In_2370);
xor U7210 (N_7210,In_4541,In_2131);
xor U7211 (N_7211,In_817,In_2045);
or U7212 (N_7212,In_1899,In_597);
xor U7213 (N_7213,In_1331,In_1547);
or U7214 (N_7214,In_3795,In_1986);
or U7215 (N_7215,In_3344,In_1475);
nor U7216 (N_7216,In_331,In_335);
nor U7217 (N_7217,In_2080,In_1108);
or U7218 (N_7218,In_2103,In_4635);
nand U7219 (N_7219,In_2050,In_2035);
nand U7220 (N_7220,In_3675,In_2084);
xor U7221 (N_7221,In_4170,In_2377);
nor U7222 (N_7222,In_2216,In_3234);
or U7223 (N_7223,In_314,In_1449);
nand U7224 (N_7224,In_469,In_3147);
nand U7225 (N_7225,In_2075,In_2743);
xor U7226 (N_7226,In_2785,In_1019);
xnor U7227 (N_7227,In_3625,In_2422);
nand U7228 (N_7228,In_2331,In_1256);
xnor U7229 (N_7229,In_3025,In_4576);
nor U7230 (N_7230,In_1481,In_4531);
nand U7231 (N_7231,In_4107,In_447);
and U7232 (N_7232,In_4144,In_2144);
xor U7233 (N_7233,In_2766,In_701);
and U7234 (N_7234,In_3984,In_894);
nor U7235 (N_7235,In_3505,In_3496);
and U7236 (N_7236,In_1872,In_557);
nor U7237 (N_7237,In_1476,In_2000);
or U7238 (N_7238,In_835,In_2166);
nor U7239 (N_7239,In_3102,In_4477);
nand U7240 (N_7240,In_112,In_909);
nand U7241 (N_7241,In_1798,In_2705);
xnor U7242 (N_7242,In_3259,In_3900);
nand U7243 (N_7243,In_4766,In_1882);
or U7244 (N_7244,In_734,In_156);
nand U7245 (N_7245,In_656,In_151);
xor U7246 (N_7246,In_1796,In_4333);
xor U7247 (N_7247,In_2709,In_521);
or U7248 (N_7248,In_492,In_3905);
xor U7249 (N_7249,In_4047,In_2069);
xnor U7250 (N_7250,In_1393,In_1959);
and U7251 (N_7251,In_3253,In_2793);
nand U7252 (N_7252,In_4935,In_1126);
nor U7253 (N_7253,In_1763,In_963);
nor U7254 (N_7254,In_2831,In_4883);
or U7255 (N_7255,In_4363,In_4536);
nand U7256 (N_7256,In_535,In_193);
nand U7257 (N_7257,In_1085,In_1617);
or U7258 (N_7258,In_1352,In_4058);
xor U7259 (N_7259,In_3571,In_1541);
or U7260 (N_7260,In_723,In_768);
and U7261 (N_7261,In_1496,In_2383);
nor U7262 (N_7262,In_4321,In_2028);
xnor U7263 (N_7263,In_3835,In_4585);
nor U7264 (N_7264,In_4107,In_3305);
nand U7265 (N_7265,In_2877,In_4910);
nand U7266 (N_7266,In_3621,In_1064);
and U7267 (N_7267,In_3690,In_1663);
xor U7268 (N_7268,In_902,In_4801);
xor U7269 (N_7269,In_1383,In_4934);
nor U7270 (N_7270,In_4669,In_980);
nor U7271 (N_7271,In_3318,In_2048);
and U7272 (N_7272,In_2742,In_922);
and U7273 (N_7273,In_4954,In_3548);
xnor U7274 (N_7274,In_725,In_2906);
nand U7275 (N_7275,In_3416,In_3244);
nor U7276 (N_7276,In_620,In_1211);
and U7277 (N_7277,In_1047,In_4601);
nor U7278 (N_7278,In_1822,In_817);
nand U7279 (N_7279,In_921,In_4518);
nor U7280 (N_7280,In_795,In_1650);
xor U7281 (N_7281,In_1902,In_2753);
and U7282 (N_7282,In_3125,In_1945);
and U7283 (N_7283,In_850,In_2509);
nand U7284 (N_7284,In_2955,In_1957);
nand U7285 (N_7285,In_317,In_2571);
and U7286 (N_7286,In_205,In_3200);
nand U7287 (N_7287,In_1712,In_1865);
or U7288 (N_7288,In_2446,In_4014);
and U7289 (N_7289,In_2288,In_508);
xnor U7290 (N_7290,In_2165,In_2900);
and U7291 (N_7291,In_1940,In_859);
or U7292 (N_7292,In_962,In_3912);
nor U7293 (N_7293,In_1638,In_3150);
nor U7294 (N_7294,In_2583,In_4727);
and U7295 (N_7295,In_591,In_1117);
and U7296 (N_7296,In_1684,In_2682);
or U7297 (N_7297,In_4865,In_4209);
and U7298 (N_7298,In_3815,In_2773);
xor U7299 (N_7299,In_588,In_3234);
xor U7300 (N_7300,In_630,In_1231);
or U7301 (N_7301,In_3919,In_4938);
nor U7302 (N_7302,In_3825,In_2957);
nor U7303 (N_7303,In_2286,In_392);
and U7304 (N_7304,In_4772,In_3821);
nand U7305 (N_7305,In_2413,In_3002);
nand U7306 (N_7306,In_1417,In_1808);
xnor U7307 (N_7307,In_3416,In_3716);
xor U7308 (N_7308,In_317,In_4030);
nand U7309 (N_7309,In_3546,In_1852);
xnor U7310 (N_7310,In_3775,In_2259);
xnor U7311 (N_7311,In_634,In_3478);
nand U7312 (N_7312,In_3033,In_660);
xnor U7313 (N_7313,In_2445,In_4438);
nand U7314 (N_7314,In_2562,In_2274);
or U7315 (N_7315,In_872,In_4907);
and U7316 (N_7316,In_2131,In_3410);
xnor U7317 (N_7317,In_3531,In_339);
or U7318 (N_7318,In_2265,In_3928);
and U7319 (N_7319,In_53,In_3412);
xnor U7320 (N_7320,In_3587,In_392);
nand U7321 (N_7321,In_2269,In_2301);
nor U7322 (N_7322,In_4891,In_505);
xor U7323 (N_7323,In_1407,In_1972);
or U7324 (N_7324,In_3037,In_716);
xnor U7325 (N_7325,In_4466,In_490);
or U7326 (N_7326,In_3052,In_1698);
and U7327 (N_7327,In_3100,In_2833);
xnor U7328 (N_7328,In_3292,In_60);
xor U7329 (N_7329,In_1173,In_2540);
or U7330 (N_7330,In_3606,In_4617);
nand U7331 (N_7331,In_2053,In_888);
nand U7332 (N_7332,In_652,In_1994);
or U7333 (N_7333,In_3240,In_822);
nor U7334 (N_7334,In_4788,In_2930);
or U7335 (N_7335,In_352,In_4979);
xor U7336 (N_7336,In_4342,In_4253);
xnor U7337 (N_7337,In_2650,In_444);
nand U7338 (N_7338,In_117,In_1092);
nor U7339 (N_7339,In_1750,In_280);
nor U7340 (N_7340,In_1518,In_2949);
xnor U7341 (N_7341,In_501,In_4413);
and U7342 (N_7342,In_2795,In_1008);
nor U7343 (N_7343,In_4601,In_1060);
nand U7344 (N_7344,In_609,In_564);
and U7345 (N_7345,In_1045,In_994);
and U7346 (N_7346,In_4023,In_1893);
nand U7347 (N_7347,In_563,In_2727);
nand U7348 (N_7348,In_139,In_541);
xor U7349 (N_7349,In_2821,In_718);
or U7350 (N_7350,In_37,In_4990);
or U7351 (N_7351,In_2004,In_3318);
nand U7352 (N_7352,In_3374,In_3367);
nor U7353 (N_7353,In_4229,In_2636);
nand U7354 (N_7354,In_1997,In_2314);
and U7355 (N_7355,In_4038,In_3785);
nand U7356 (N_7356,In_652,In_4985);
or U7357 (N_7357,In_546,In_2930);
nor U7358 (N_7358,In_468,In_4933);
or U7359 (N_7359,In_2898,In_2128);
nor U7360 (N_7360,In_3641,In_166);
xnor U7361 (N_7361,In_1942,In_2665);
or U7362 (N_7362,In_3088,In_2424);
nand U7363 (N_7363,In_4862,In_4211);
xor U7364 (N_7364,In_4693,In_3879);
or U7365 (N_7365,In_4956,In_4264);
nor U7366 (N_7366,In_3676,In_759);
nand U7367 (N_7367,In_2413,In_4861);
xnor U7368 (N_7368,In_2919,In_523);
xnor U7369 (N_7369,In_186,In_1995);
xnor U7370 (N_7370,In_1586,In_4958);
nor U7371 (N_7371,In_3936,In_3886);
and U7372 (N_7372,In_2985,In_76);
and U7373 (N_7373,In_1676,In_1883);
xor U7374 (N_7374,In_3695,In_606);
and U7375 (N_7375,In_2700,In_4424);
nand U7376 (N_7376,In_1930,In_511);
nand U7377 (N_7377,In_1810,In_325);
xnor U7378 (N_7378,In_3764,In_4131);
or U7379 (N_7379,In_1370,In_501);
or U7380 (N_7380,In_4694,In_466);
or U7381 (N_7381,In_1577,In_29);
and U7382 (N_7382,In_3404,In_4737);
and U7383 (N_7383,In_3852,In_730);
xnor U7384 (N_7384,In_752,In_3166);
nand U7385 (N_7385,In_280,In_1875);
nand U7386 (N_7386,In_4228,In_1755);
or U7387 (N_7387,In_4953,In_361);
and U7388 (N_7388,In_4338,In_1446);
and U7389 (N_7389,In_4700,In_879);
and U7390 (N_7390,In_917,In_4802);
or U7391 (N_7391,In_1042,In_4469);
and U7392 (N_7392,In_1360,In_2950);
xnor U7393 (N_7393,In_1202,In_1781);
nor U7394 (N_7394,In_2896,In_2091);
and U7395 (N_7395,In_4301,In_4426);
or U7396 (N_7396,In_4238,In_1338);
or U7397 (N_7397,In_2972,In_530);
xor U7398 (N_7398,In_4837,In_3350);
and U7399 (N_7399,In_1603,In_686);
nor U7400 (N_7400,In_3968,In_1770);
nand U7401 (N_7401,In_1013,In_1222);
nor U7402 (N_7402,In_3599,In_2920);
nor U7403 (N_7403,In_4523,In_1263);
xnor U7404 (N_7404,In_3097,In_4760);
or U7405 (N_7405,In_4634,In_383);
nand U7406 (N_7406,In_3138,In_1401);
or U7407 (N_7407,In_1185,In_102);
and U7408 (N_7408,In_2430,In_3729);
xor U7409 (N_7409,In_845,In_541);
nand U7410 (N_7410,In_1347,In_104);
nand U7411 (N_7411,In_2482,In_2348);
or U7412 (N_7412,In_57,In_3190);
nor U7413 (N_7413,In_3180,In_4511);
and U7414 (N_7414,In_3492,In_4401);
nor U7415 (N_7415,In_4005,In_712);
or U7416 (N_7416,In_158,In_4538);
xnor U7417 (N_7417,In_4622,In_1882);
nor U7418 (N_7418,In_4904,In_1747);
or U7419 (N_7419,In_1418,In_1100);
xnor U7420 (N_7420,In_701,In_2868);
xor U7421 (N_7421,In_4314,In_4071);
and U7422 (N_7422,In_1784,In_2866);
nor U7423 (N_7423,In_1059,In_407);
and U7424 (N_7424,In_2921,In_34);
or U7425 (N_7425,In_2523,In_141);
or U7426 (N_7426,In_4210,In_389);
and U7427 (N_7427,In_1299,In_3124);
xnor U7428 (N_7428,In_3949,In_587);
xnor U7429 (N_7429,In_4491,In_862);
or U7430 (N_7430,In_3466,In_2524);
nor U7431 (N_7431,In_4819,In_111);
nor U7432 (N_7432,In_2218,In_1837);
xnor U7433 (N_7433,In_2536,In_4012);
nand U7434 (N_7434,In_104,In_4893);
or U7435 (N_7435,In_2459,In_4924);
nor U7436 (N_7436,In_545,In_2502);
and U7437 (N_7437,In_4179,In_4198);
or U7438 (N_7438,In_614,In_2979);
nand U7439 (N_7439,In_4057,In_815);
xor U7440 (N_7440,In_2963,In_4677);
nand U7441 (N_7441,In_2623,In_4728);
nor U7442 (N_7442,In_2555,In_2528);
xnor U7443 (N_7443,In_3072,In_870);
or U7444 (N_7444,In_1643,In_4681);
nand U7445 (N_7445,In_1147,In_589);
nor U7446 (N_7446,In_254,In_4153);
nand U7447 (N_7447,In_4333,In_3654);
or U7448 (N_7448,In_4857,In_1402);
nor U7449 (N_7449,In_515,In_1934);
and U7450 (N_7450,In_922,In_3614);
xor U7451 (N_7451,In_3711,In_2256);
nand U7452 (N_7452,In_1877,In_3180);
xor U7453 (N_7453,In_2771,In_925);
nor U7454 (N_7454,In_363,In_1739);
xor U7455 (N_7455,In_3334,In_3013);
nand U7456 (N_7456,In_309,In_4397);
or U7457 (N_7457,In_1967,In_4869);
nand U7458 (N_7458,In_4595,In_727);
xor U7459 (N_7459,In_4659,In_1235);
or U7460 (N_7460,In_2400,In_4064);
or U7461 (N_7461,In_3419,In_1072);
nand U7462 (N_7462,In_2072,In_2367);
nand U7463 (N_7463,In_32,In_1159);
xor U7464 (N_7464,In_1678,In_2271);
xor U7465 (N_7465,In_3991,In_3628);
and U7466 (N_7466,In_3956,In_1462);
and U7467 (N_7467,In_321,In_3926);
and U7468 (N_7468,In_3668,In_1624);
nand U7469 (N_7469,In_3560,In_1);
nor U7470 (N_7470,In_4686,In_3664);
and U7471 (N_7471,In_4561,In_70);
nor U7472 (N_7472,In_2284,In_242);
nor U7473 (N_7473,In_2879,In_4031);
xnor U7474 (N_7474,In_2337,In_2264);
nand U7475 (N_7475,In_547,In_2601);
xor U7476 (N_7476,In_2051,In_2113);
nand U7477 (N_7477,In_3816,In_4763);
nand U7478 (N_7478,In_4845,In_3235);
nand U7479 (N_7479,In_786,In_897);
nor U7480 (N_7480,In_127,In_2308);
nor U7481 (N_7481,In_3127,In_1288);
nor U7482 (N_7482,In_3657,In_2524);
nand U7483 (N_7483,In_2958,In_2129);
or U7484 (N_7484,In_4425,In_3735);
nor U7485 (N_7485,In_3871,In_1822);
nand U7486 (N_7486,In_1657,In_90);
nor U7487 (N_7487,In_2995,In_1151);
or U7488 (N_7488,In_3971,In_1568);
nand U7489 (N_7489,In_222,In_2850);
and U7490 (N_7490,In_3812,In_1953);
nor U7491 (N_7491,In_3740,In_2487);
xnor U7492 (N_7492,In_1782,In_2288);
and U7493 (N_7493,In_1035,In_2224);
nor U7494 (N_7494,In_617,In_772);
and U7495 (N_7495,In_2510,In_789);
and U7496 (N_7496,In_1362,In_4032);
or U7497 (N_7497,In_544,In_4567);
and U7498 (N_7498,In_3384,In_4909);
and U7499 (N_7499,In_984,In_1254);
and U7500 (N_7500,In_2231,In_1280);
nand U7501 (N_7501,In_1999,In_4772);
nand U7502 (N_7502,In_3425,In_1660);
and U7503 (N_7503,In_3820,In_3958);
nand U7504 (N_7504,In_2783,In_10);
nor U7505 (N_7505,In_4689,In_2568);
xnor U7506 (N_7506,In_293,In_3805);
xnor U7507 (N_7507,In_4708,In_599);
or U7508 (N_7508,In_4896,In_3395);
or U7509 (N_7509,In_375,In_3847);
nand U7510 (N_7510,In_3081,In_2847);
or U7511 (N_7511,In_4511,In_1503);
or U7512 (N_7512,In_1237,In_3421);
xnor U7513 (N_7513,In_4258,In_3556);
or U7514 (N_7514,In_3048,In_3526);
and U7515 (N_7515,In_3308,In_2880);
xnor U7516 (N_7516,In_4716,In_4837);
nor U7517 (N_7517,In_3728,In_3990);
or U7518 (N_7518,In_3855,In_628);
nor U7519 (N_7519,In_4478,In_3893);
nor U7520 (N_7520,In_431,In_1139);
nand U7521 (N_7521,In_3825,In_4868);
or U7522 (N_7522,In_1664,In_664);
nand U7523 (N_7523,In_1893,In_1405);
and U7524 (N_7524,In_1107,In_2059);
xor U7525 (N_7525,In_1419,In_2235);
and U7526 (N_7526,In_538,In_3695);
and U7527 (N_7527,In_1695,In_3378);
and U7528 (N_7528,In_4150,In_4765);
nor U7529 (N_7529,In_3962,In_4205);
and U7530 (N_7530,In_1133,In_3529);
xnor U7531 (N_7531,In_2232,In_811);
and U7532 (N_7532,In_733,In_4200);
xnor U7533 (N_7533,In_3197,In_4572);
nor U7534 (N_7534,In_540,In_690);
nor U7535 (N_7535,In_712,In_3269);
nor U7536 (N_7536,In_70,In_2074);
nand U7537 (N_7537,In_2292,In_4466);
nor U7538 (N_7538,In_4702,In_1599);
and U7539 (N_7539,In_801,In_2651);
xor U7540 (N_7540,In_2328,In_601);
or U7541 (N_7541,In_880,In_1060);
xnor U7542 (N_7542,In_835,In_448);
or U7543 (N_7543,In_2828,In_155);
or U7544 (N_7544,In_4928,In_729);
xor U7545 (N_7545,In_1204,In_3965);
nor U7546 (N_7546,In_1025,In_3161);
nand U7547 (N_7547,In_3981,In_1031);
nand U7548 (N_7548,In_3357,In_1776);
nand U7549 (N_7549,In_1504,In_3392);
xnor U7550 (N_7550,In_3217,In_1954);
or U7551 (N_7551,In_3607,In_4875);
or U7552 (N_7552,In_2467,In_3205);
nor U7553 (N_7553,In_3933,In_1725);
nor U7554 (N_7554,In_713,In_4257);
or U7555 (N_7555,In_3447,In_4579);
xor U7556 (N_7556,In_4742,In_2140);
and U7557 (N_7557,In_4693,In_875);
nor U7558 (N_7558,In_2806,In_2714);
nor U7559 (N_7559,In_4697,In_4605);
nor U7560 (N_7560,In_342,In_3036);
or U7561 (N_7561,In_2003,In_3383);
nand U7562 (N_7562,In_2847,In_2492);
or U7563 (N_7563,In_3980,In_801);
nand U7564 (N_7564,In_3384,In_1470);
xnor U7565 (N_7565,In_1254,In_3663);
xor U7566 (N_7566,In_1026,In_859);
nand U7567 (N_7567,In_146,In_120);
and U7568 (N_7568,In_3059,In_833);
nor U7569 (N_7569,In_3601,In_3795);
and U7570 (N_7570,In_4919,In_2096);
and U7571 (N_7571,In_1991,In_1519);
nand U7572 (N_7572,In_757,In_235);
nand U7573 (N_7573,In_4192,In_3507);
nor U7574 (N_7574,In_471,In_2397);
xnor U7575 (N_7575,In_4261,In_2929);
or U7576 (N_7576,In_1637,In_779);
xnor U7577 (N_7577,In_4654,In_152);
nor U7578 (N_7578,In_3468,In_3502);
or U7579 (N_7579,In_644,In_2934);
nor U7580 (N_7580,In_4393,In_2090);
xnor U7581 (N_7581,In_4704,In_3781);
and U7582 (N_7582,In_571,In_736);
nor U7583 (N_7583,In_700,In_1256);
nor U7584 (N_7584,In_4001,In_3046);
nor U7585 (N_7585,In_349,In_3176);
xnor U7586 (N_7586,In_45,In_161);
nand U7587 (N_7587,In_4013,In_4007);
nor U7588 (N_7588,In_2514,In_3625);
nand U7589 (N_7589,In_299,In_2870);
nand U7590 (N_7590,In_198,In_1656);
nand U7591 (N_7591,In_323,In_2141);
nor U7592 (N_7592,In_234,In_632);
and U7593 (N_7593,In_1974,In_360);
or U7594 (N_7594,In_2925,In_3043);
xnor U7595 (N_7595,In_4956,In_4686);
or U7596 (N_7596,In_484,In_3801);
nand U7597 (N_7597,In_698,In_1928);
nor U7598 (N_7598,In_844,In_3335);
and U7599 (N_7599,In_4207,In_114);
nor U7600 (N_7600,In_1427,In_2113);
nand U7601 (N_7601,In_909,In_2405);
nor U7602 (N_7602,In_19,In_905);
nand U7603 (N_7603,In_3165,In_1965);
nor U7604 (N_7604,In_3506,In_181);
or U7605 (N_7605,In_3914,In_2703);
xor U7606 (N_7606,In_3786,In_3130);
and U7607 (N_7607,In_610,In_1670);
and U7608 (N_7608,In_4391,In_2909);
or U7609 (N_7609,In_2713,In_2972);
or U7610 (N_7610,In_464,In_430);
nand U7611 (N_7611,In_4601,In_1362);
nor U7612 (N_7612,In_2810,In_3274);
or U7613 (N_7613,In_4161,In_1080);
xnor U7614 (N_7614,In_4816,In_3395);
xor U7615 (N_7615,In_1932,In_1261);
xor U7616 (N_7616,In_4118,In_4714);
and U7617 (N_7617,In_1941,In_952);
and U7618 (N_7618,In_812,In_3106);
nand U7619 (N_7619,In_4676,In_4698);
and U7620 (N_7620,In_252,In_4693);
and U7621 (N_7621,In_2932,In_4452);
nor U7622 (N_7622,In_237,In_2729);
nor U7623 (N_7623,In_1342,In_4073);
nand U7624 (N_7624,In_3050,In_531);
xor U7625 (N_7625,In_1896,In_1478);
and U7626 (N_7626,In_4350,In_3658);
nand U7627 (N_7627,In_1031,In_424);
and U7628 (N_7628,In_1911,In_2411);
nand U7629 (N_7629,In_3371,In_1414);
or U7630 (N_7630,In_241,In_1393);
nand U7631 (N_7631,In_439,In_4154);
nand U7632 (N_7632,In_3887,In_4907);
and U7633 (N_7633,In_1250,In_3270);
or U7634 (N_7634,In_4421,In_1603);
xor U7635 (N_7635,In_4708,In_2886);
nand U7636 (N_7636,In_1254,In_3527);
and U7637 (N_7637,In_109,In_2589);
or U7638 (N_7638,In_4659,In_4395);
nand U7639 (N_7639,In_330,In_1680);
xnor U7640 (N_7640,In_3558,In_4074);
nand U7641 (N_7641,In_3925,In_2418);
nor U7642 (N_7642,In_3818,In_2403);
xnor U7643 (N_7643,In_1218,In_2381);
xor U7644 (N_7644,In_4480,In_2750);
nor U7645 (N_7645,In_583,In_4221);
xnor U7646 (N_7646,In_2572,In_3015);
and U7647 (N_7647,In_4436,In_4007);
nand U7648 (N_7648,In_2250,In_103);
nor U7649 (N_7649,In_4818,In_2246);
and U7650 (N_7650,In_4508,In_1048);
and U7651 (N_7651,In_1743,In_4188);
nand U7652 (N_7652,In_459,In_4467);
and U7653 (N_7653,In_2043,In_150);
nand U7654 (N_7654,In_525,In_213);
and U7655 (N_7655,In_8,In_3173);
and U7656 (N_7656,In_4055,In_4815);
and U7657 (N_7657,In_3598,In_3200);
or U7658 (N_7658,In_4340,In_3702);
or U7659 (N_7659,In_4723,In_176);
xnor U7660 (N_7660,In_1803,In_1882);
nand U7661 (N_7661,In_1638,In_1560);
nand U7662 (N_7662,In_1758,In_1441);
and U7663 (N_7663,In_2808,In_3046);
nand U7664 (N_7664,In_3514,In_7);
and U7665 (N_7665,In_374,In_3040);
nor U7666 (N_7666,In_1454,In_4157);
and U7667 (N_7667,In_669,In_1406);
xnor U7668 (N_7668,In_3359,In_3255);
xor U7669 (N_7669,In_2426,In_4696);
or U7670 (N_7670,In_1700,In_1925);
nand U7671 (N_7671,In_1645,In_3438);
nor U7672 (N_7672,In_2900,In_4993);
and U7673 (N_7673,In_4101,In_4611);
nor U7674 (N_7674,In_4360,In_3302);
and U7675 (N_7675,In_4960,In_3275);
and U7676 (N_7676,In_1587,In_3292);
nor U7677 (N_7677,In_4221,In_3727);
nand U7678 (N_7678,In_243,In_633);
and U7679 (N_7679,In_1698,In_1941);
nand U7680 (N_7680,In_3552,In_430);
nor U7681 (N_7681,In_167,In_2247);
and U7682 (N_7682,In_1690,In_2909);
xnor U7683 (N_7683,In_3257,In_1248);
xor U7684 (N_7684,In_350,In_3921);
xor U7685 (N_7685,In_818,In_766);
nand U7686 (N_7686,In_3290,In_277);
nand U7687 (N_7687,In_283,In_2891);
xor U7688 (N_7688,In_4968,In_4191);
or U7689 (N_7689,In_2624,In_547);
nand U7690 (N_7690,In_342,In_2002);
nand U7691 (N_7691,In_2722,In_4743);
nor U7692 (N_7692,In_4541,In_1088);
nor U7693 (N_7693,In_1517,In_3894);
and U7694 (N_7694,In_3242,In_1473);
xnor U7695 (N_7695,In_866,In_1188);
or U7696 (N_7696,In_2675,In_4852);
nor U7697 (N_7697,In_4927,In_832);
and U7698 (N_7698,In_3831,In_1829);
or U7699 (N_7699,In_1134,In_2368);
nor U7700 (N_7700,In_3803,In_4495);
nand U7701 (N_7701,In_1342,In_846);
xnor U7702 (N_7702,In_4833,In_3037);
and U7703 (N_7703,In_550,In_3721);
or U7704 (N_7704,In_3316,In_2547);
and U7705 (N_7705,In_4031,In_4214);
nand U7706 (N_7706,In_1760,In_1271);
nor U7707 (N_7707,In_2627,In_509);
and U7708 (N_7708,In_2258,In_2185);
or U7709 (N_7709,In_2367,In_156);
or U7710 (N_7710,In_976,In_1925);
nand U7711 (N_7711,In_2445,In_2336);
or U7712 (N_7712,In_3253,In_101);
xor U7713 (N_7713,In_1666,In_4806);
nand U7714 (N_7714,In_3031,In_324);
nor U7715 (N_7715,In_4212,In_1150);
xnor U7716 (N_7716,In_2230,In_1883);
nand U7717 (N_7717,In_1584,In_3190);
nor U7718 (N_7718,In_3275,In_396);
xnor U7719 (N_7719,In_1155,In_3860);
or U7720 (N_7720,In_236,In_4405);
nand U7721 (N_7721,In_1237,In_118);
xor U7722 (N_7722,In_927,In_895);
nor U7723 (N_7723,In_1230,In_4131);
and U7724 (N_7724,In_2262,In_1635);
nand U7725 (N_7725,In_3901,In_2503);
or U7726 (N_7726,In_311,In_4517);
and U7727 (N_7727,In_1802,In_4205);
xnor U7728 (N_7728,In_3286,In_2202);
nor U7729 (N_7729,In_1714,In_1993);
xor U7730 (N_7730,In_2316,In_2928);
xor U7731 (N_7731,In_1179,In_1361);
xor U7732 (N_7732,In_2809,In_4489);
xnor U7733 (N_7733,In_2117,In_2749);
nor U7734 (N_7734,In_3980,In_3841);
nor U7735 (N_7735,In_3554,In_968);
xnor U7736 (N_7736,In_2281,In_685);
nand U7737 (N_7737,In_404,In_2296);
nor U7738 (N_7738,In_1435,In_1010);
nor U7739 (N_7739,In_226,In_2769);
or U7740 (N_7740,In_2753,In_3606);
or U7741 (N_7741,In_214,In_817);
and U7742 (N_7742,In_202,In_2043);
nand U7743 (N_7743,In_2999,In_3182);
or U7744 (N_7744,In_1465,In_1694);
xnor U7745 (N_7745,In_3773,In_1562);
or U7746 (N_7746,In_3875,In_947);
nand U7747 (N_7747,In_751,In_4155);
and U7748 (N_7748,In_4544,In_2316);
nand U7749 (N_7749,In_1048,In_4326);
and U7750 (N_7750,In_1287,In_4971);
and U7751 (N_7751,In_3162,In_3157);
nor U7752 (N_7752,In_1535,In_481);
nand U7753 (N_7753,In_3724,In_1594);
nor U7754 (N_7754,In_2560,In_2450);
xor U7755 (N_7755,In_2955,In_292);
or U7756 (N_7756,In_1212,In_162);
xor U7757 (N_7757,In_3609,In_3523);
or U7758 (N_7758,In_2165,In_1464);
nand U7759 (N_7759,In_3827,In_4239);
nor U7760 (N_7760,In_2211,In_945);
and U7761 (N_7761,In_1549,In_1535);
nand U7762 (N_7762,In_4562,In_3603);
nand U7763 (N_7763,In_2308,In_125);
xnor U7764 (N_7764,In_3192,In_3044);
and U7765 (N_7765,In_3262,In_4454);
nor U7766 (N_7766,In_2068,In_1043);
nor U7767 (N_7767,In_1682,In_338);
nand U7768 (N_7768,In_3743,In_4441);
nand U7769 (N_7769,In_3887,In_2174);
nor U7770 (N_7770,In_4336,In_4852);
xnor U7771 (N_7771,In_236,In_290);
and U7772 (N_7772,In_3517,In_2537);
and U7773 (N_7773,In_710,In_2855);
and U7774 (N_7774,In_264,In_3434);
and U7775 (N_7775,In_3860,In_3923);
nand U7776 (N_7776,In_1996,In_882);
nor U7777 (N_7777,In_1083,In_510);
xnor U7778 (N_7778,In_4702,In_2502);
nor U7779 (N_7779,In_2351,In_3928);
and U7780 (N_7780,In_2890,In_124);
nor U7781 (N_7781,In_134,In_4357);
and U7782 (N_7782,In_4698,In_2158);
or U7783 (N_7783,In_4481,In_110);
nand U7784 (N_7784,In_1499,In_1886);
nand U7785 (N_7785,In_2154,In_3881);
and U7786 (N_7786,In_4675,In_1662);
nor U7787 (N_7787,In_110,In_3804);
and U7788 (N_7788,In_1325,In_1346);
nor U7789 (N_7789,In_4298,In_936);
nand U7790 (N_7790,In_748,In_4044);
nor U7791 (N_7791,In_2606,In_589);
or U7792 (N_7792,In_4298,In_1520);
or U7793 (N_7793,In_20,In_2685);
nor U7794 (N_7794,In_2522,In_3102);
and U7795 (N_7795,In_2111,In_992);
nand U7796 (N_7796,In_1559,In_3786);
nand U7797 (N_7797,In_158,In_3252);
xor U7798 (N_7798,In_1836,In_4879);
xnor U7799 (N_7799,In_4042,In_238);
nor U7800 (N_7800,In_628,In_81);
nor U7801 (N_7801,In_2731,In_777);
xnor U7802 (N_7802,In_4230,In_1022);
and U7803 (N_7803,In_1519,In_2880);
nor U7804 (N_7804,In_3391,In_2160);
or U7805 (N_7805,In_4474,In_2640);
xor U7806 (N_7806,In_4928,In_4410);
and U7807 (N_7807,In_4993,In_1045);
nand U7808 (N_7808,In_4987,In_2987);
xor U7809 (N_7809,In_3590,In_3777);
nand U7810 (N_7810,In_1822,In_3688);
or U7811 (N_7811,In_4981,In_468);
or U7812 (N_7812,In_2693,In_1545);
nor U7813 (N_7813,In_3056,In_3957);
and U7814 (N_7814,In_1455,In_3373);
or U7815 (N_7815,In_4891,In_1896);
xnor U7816 (N_7816,In_3497,In_4430);
nand U7817 (N_7817,In_2666,In_4759);
nor U7818 (N_7818,In_3565,In_4458);
and U7819 (N_7819,In_406,In_1399);
xnor U7820 (N_7820,In_313,In_3179);
or U7821 (N_7821,In_546,In_4414);
and U7822 (N_7822,In_3118,In_3522);
or U7823 (N_7823,In_3561,In_3032);
nand U7824 (N_7824,In_2662,In_83);
xnor U7825 (N_7825,In_1341,In_1182);
and U7826 (N_7826,In_4754,In_2158);
nor U7827 (N_7827,In_215,In_4547);
nor U7828 (N_7828,In_1520,In_2242);
nand U7829 (N_7829,In_1443,In_1352);
nand U7830 (N_7830,In_3819,In_833);
nor U7831 (N_7831,In_1290,In_2626);
xnor U7832 (N_7832,In_225,In_1218);
and U7833 (N_7833,In_1615,In_983);
and U7834 (N_7834,In_1543,In_4181);
nand U7835 (N_7835,In_4646,In_1102);
nand U7836 (N_7836,In_1529,In_189);
nand U7837 (N_7837,In_2429,In_353);
nand U7838 (N_7838,In_3724,In_3797);
or U7839 (N_7839,In_104,In_3753);
nand U7840 (N_7840,In_2904,In_2413);
or U7841 (N_7841,In_1213,In_1413);
nor U7842 (N_7842,In_642,In_1753);
nor U7843 (N_7843,In_4589,In_2108);
nand U7844 (N_7844,In_1147,In_2502);
or U7845 (N_7845,In_2612,In_2869);
nand U7846 (N_7846,In_573,In_635);
and U7847 (N_7847,In_1890,In_899);
or U7848 (N_7848,In_963,In_2952);
nand U7849 (N_7849,In_3305,In_3185);
xnor U7850 (N_7850,In_2983,In_2804);
and U7851 (N_7851,In_1991,In_1008);
nor U7852 (N_7852,In_2904,In_528);
and U7853 (N_7853,In_4967,In_3335);
or U7854 (N_7854,In_3503,In_2709);
and U7855 (N_7855,In_2026,In_1721);
or U7856 (N_7856,In_1672,In_852);
and U7857 (N_7857,In_4747,In_3283);
xnor U7858 (N_7858,In_3956,In_739);
xnor U7859 (N_7859,In_358,In_1797);
xor U7860 (N_7860,In_4993,In_4302);
nor U7861 (N_7861,In_2836,In_2940);
xor U7862 (N_7862,In_984,In_519);
or U7863 (N_7863,In_2585,In_1126);
nor U7864 (N_7864,In_4621,In_3474);
or U7865 (N_7865,In_4739,In_3410);
or U7866 (N_7866,In_3974,In_623);
xor U7867 (N_7867,In_293,In_999);
nor U7868 (N_7868,In_4445,In_4834);
nor U7869 (N_7869,In_1647,In_4967);
xnor U7870 (N_7870,In_2456,In_2577);
or U7871 (N_7871,In_2761,In_76);
nand U7872 (N_7872,In_4864,In_2362);
and U7873 (N_7873,In_2686,In_3374);
nand U7874 (N_7874,In_2344,In_4633);
nand U7875 (N_7875,In_16,In_4691);
nor U7876 (N_7876,In_1162,In_2243);
xor U7877 (N_7877,In_768,In_4959);
and U7878 (N_7878,In_797,In_1322);
xor U7879 (N_7879,In_39,In_3955);
xor U7880 (N_7880,In_1576,In_2253);
nand U7881 (N_7881,In_2073,In_2290);
or U7882 (N_7882,In_3846,In_2318);
or U7883 (N_7883,In_1774,In_3897);
nand U7884 (N_7884,In_1458,In_971);
nand U7885 (N_7885,In_175,In_2008);
nor U7886 (N_7886,In_2403,In_3361);
or U7887 (N_7887,In_1472,In_1541);
nand U7888 (N_7888,In_1636,In_956);
or U7889 (N_7889,In_3133,In_3538);
and U7890 (N_7890,In_1048,In_998);
and U7891 (N_7891,In_4754,In_3962);
nand U7892 (N_7892,In_1103,In_2823);
xor U7893 (N_7893,In_716,In_1558);
or U7894 (N_7894,In_4352,In_1476);
or U7895 (N_7895,In_4025,In_3561);
or U7896 (N_7896,In_1844,In_1334);
xnor U7897 (N_7897,In_3015,In_3997);
xnor U7898 (N_7898,In_2400,In_3544);
nand U7899 (N_7899,In_4699,In_3352);
nor U7900 (N_7900,In_3882,In_1774);
nor U7901 (N_7901,In_4516,In_875);
xor U7902 (N_7902,In_4700,In_3452);
nor U7903 (N_7903,In_1589,In_1768);
xor U7904 (N_7904,In_4292,In_2334);
nand U7905 (N_7905,In_4642,In_4641);
nand U7906 (N_7906,In_2668,In_2006);
nor U7907 (N_7907,In_2897,In_2345);
or U7908 (N_7908,In_1958,In_901);
nand U7909 (N_7909,In_4151,In_2846);
nand U7910 (N_7910,In_201,In_1774);
nand U7911 (N_7911,In_248,In_1484);
nor U7912 (N_7912,In_482,In_1310);
nand U7913 (N_7913,In_3645,In_639);
xnor U7914 (N_7914,In_4122,In_850);
nand U7915 (N_7915,In_1570,In_2735);
nor U7916 (N_7916,In_55,In_4628);
and U7917 (N_7917,In_4087,In_2752);
xnor U7918 (N_7918,In_3976,In_1538);
or U7919 (N_7919,In_2001,In_1428);
nand U7920 (N_7920,In_1904,In_3594);
or U7921 (N_7921,In_332,In_3554);
xor U7922 (N_7922,In_1978,In_1669);
xor U7923 (N_7923,In_535,In_1271);
nor U7924 (N_7924,In_2792,In_4281);
nand U7925 (N_7925,In_3935,In_2676);
nor U7926 (N_7926,In_4564,In_1913);
or U7927 (N_7927,In_3970,In_2119);
nor U7928 (N_7928,In_4798,In_3044);
xnor U7929 (N_7929,In_4029,In_607);
nor U7930 (N_7930,In_3271,In_4946);
nor U7931 (N_7931,In_3909,In_2176);
nand U7932 (N_7932,In_2155,In_834);
or U7933 (N_7933,In_1435,In_3649);
xor U7934 (N_7934,In_859,In_2664);
and U7935 (N_7935,In_601,In_405);
and U7936 (N_7936,In_2981,In_1697);
or U7937 (N_7937,In_3975,In_1929);
xor U7938 (N_7938,In_3718,In_1646);
nand U7939 (N_7939,In_1909,In_2094);
and U7940 (N_7940,In_4605,In_3843);
nor U7941 (N_7941,In_3257,In_1518);
xor U7942 (N_7942,In_3856,In_1233);
and U7943 (N_7943,In_4766,In_4902);
and U7944 (N_7944,In_4950,In_2505);
nand U7945 (N_7945,In_1962,In_19);
and U7946 (N_7946,In_569,In_2550);
xor U7947 (N_7947,In_4168,In_3846);
nand U7948 (N_7948,In_892,In_10);
and U7949 (N_7949,In_1002,In_2039);
or U7950 (N_7950,In_2117,In_4866);
nor U7951 (N_7951,In_194,In_2542);
and U7952 (N_7952,In_1730,In_2447);
or U7953 (N_7953,In_2128,In_1572);
xnor U7954 (N_7954,In_4859,In_1201);
or U7955 (N_7955,In_1029,In_2045);
nor U7956 (N_7956,In_3765,In_3242);
nor U7957 (N_7957,In_3067,In_1828);
nand U7958 (N_7958,In_396,In_166);
or U7959 (N_7959,In_3438,In_3590);
and U7960 (N_7960,In_4655,In_4682);
nor U7961 (N_7961,In_3674,In_4194);
or U7962 (N_7962,In_2688,In_622);
or U7963 (N_7963,In_2018,In_364);
nand U7964 (N_7964,In_2755,In_2164);
xnor U7965 (N_7965,In_4738,In_2484);
nor U7966 (N_7966,In_4061,In_1136);
nand U7967 (N_7967,In_1753,In_479);
nand U7968 (N_7968,In_3339,In_1727);
nand U7969 (N_7969,In_4448,In_4940);
xnor U7970 (N_7970,In_1224,In_3390);
and U7971 (N_7971,In_2147,In_3871);
nor U7972 (N_7972,In_1613,In_3640);
nand U7973 (N_7973,In_4265,In_1686);
nor U7974 (N_7974,In_1945,In_3138);
xnor U7975 (N_7975,In_4267,In_3596);
nand U7976 (N_7976,In_4705,In_3312);
nor U7977 (N_7977,In_3070,In_378);
xnor U7978 (N_7978,In_1038,In_64);
nor U7979 (N_7979,In_4788,In_3034);
nand U7980 (N_7980,In_1795,In_24);
and U7981 (N_7981,In_3148,In_2821);
xnor U7982 (N_7982,In_3623,In_4510);
nand U7983 (N_7983,In_4555,In_2664);
or U7984 (N_7984,In_2613,In_3831);
and U7985 (N_7985,In_923,In_1692);
xor U7986 (N_7986,In_3786,In_2819);
nor U7987 (N_7987,In_1308,In_4704);
nor U7988 (N_7988,In_800,In_2279);
or U7989 (N_7989,In_843,In_2211);
and U7990 (N_7990,In_1189,In_3077);
and U7991 (N_7991,In_629,In_4892);
xor U7992 (N_7992,In_3604,In_2718);
xnor U7993 (N_7993,In_4269,In_3287);
or U7994 (N_7994,In_3214,In_4287);
or U7995 (N_7995,In_3398,In_4377);
nand U7996 (N_7996,In_1893,In_1503);
xnor U7997 (N_7997,In_2777,In_1023);
nor U7998 (N_7998,In_3315,In_1934);
or U7999 (N_7999,In_1232,In_1356);
and U8000 (N_8000,In_140,In_2819);
xnor U8001 (N_8001,In_3509,In_1783);
nand U8002 (N_8002,In_3891,In_888);
xor U8003 (N_8003,In_1821,In_2836);
and U8004 (N_8004,In_4758,In_3934);
or U8005 (N_8005,In_2268,In_1653);
or U8006 (N_8006,In_1118,In_3671);
nand U8007 (N_8007,In_1383,In_3490);
and U8008 (N_8008,In_1040,In_363);
or U8009 (N_8009,In_2717,In_625);
and U8010 (N_8010,In_3484,In_3696);
and U8011 (N_8011,In_4148,In_1736);
and U8012 (N_8012,In_2821,In_4612);
and U8013 (N_8013,In_662,In_2509);
xor U8014 (N_8014,In_1423,In_3374);
xor U8015 (N_8015,In_3979,In_2285);
nand U8016 (N_8016,In_4173,In_780);
xor U8017 (N_8017,In_2561,In_2339);
nand U8018 (N_8018,In_1896,In_1450);
or U8019 (N_8019,In_1512,In_3167);
xor U8020 (N_8020,In_4146,In_3743);
nor U8021 (N_8021,In_4717,In_3394);
nor U8022 (N_8022,In_480,In_3746);
or U8023 (N_8023,In_3392,In_4017);
and U8024 (N_8024,In_3029,In_4615);
nor U8025 (N_8025,In_3478,In_4634);
nor U8026 (N_8026,In_838,In_3959);
or U8027 (N_8027,In_4765,In_3106);
nor U8028 (N_8028,In_1582,In_4114);
and U8029 (N_8029,In_621,In_48);
nand U8030 (N_8030,In_1420,In_3360);
or U8031 (N_8031,In_545,In_3174);
nand U8032 (N_8032,In_2981,In_1022);
or U8033 (N_8033,In_117,In_146);
and U8034 (N_8034,In_1227,In_2218);
nor U8035 (N_8035,In_3988,In_2527);
nor U8036 (N_8036,In_3183,In_1213);
xor U8037 (N_8037,In_4829,In_1527);
xor U8038 (N_8038,In_373,In_3747);
nand U8039 (N_8039,In_3142,In_3712);
xnor U8040 (N_8040,In_4149,In_3486);
or U8041 (N_8041,In_324,In_1628);
nand U8042 (N_8042,In_4195,In_4738);
nor U8043 (N_8043,In_3625,In_2095);
nor U8044 (N_8044,In_4330,In_4954);
or U8045 (N_8045,In_1459,In_4034);
nor U8046 (N_8046,In_4474,In_749);
and U8047 (N_8047,In_877,In_2551);
xor U8048 (N_8048,In_2916,In_1879);
xor U8049 (N_8049,In_4833,In_3817);
nor U8050 (N_8050,In_3565,In_45);
nand U8051 (N_8051,In_281,In_3159);
and U8052 (N_8052,In_4084,In_4735);
or U8053 (N_8053,In_1633,In_2485);
nand U8054 (N_8054,In_2516,In_892);
or U8055 (N_8055,In_4430,In_4060);
nor U8056 (N_8056,In_4270,In_1444);
xnor U8057 (N_8057,In_2573,In_2444);
or U8058 (N_8058,In_4582,In_4952);
nand U8059 (N_8059,In_1962,In_4957);
nand U8060 (N_8060,In_2584,In_3739);
nand U8061 (N_8061,In_3457,In_2565);
xor U8062 (N_8062,In_2110,In_2660);
xor U8063 (N_8063,In_2735,In_34);
nand U8064 (N_8064,In_2178,In_1334);
and U8065 (N_8065,In_4940,In_4650);
xor U8066 (N_8066,In_4229,In_2546);
nand U8067 (N_8067,In_1089,In_253);
or U8068 (N_8068,In_4411,In_1348);
xnor U8069 (N_8069,In_4217,In_1653);
nor U8070 (N_8070,In_3838,In_2363);
or U8071 (N_8071,In_3521,In_659);
nand U8072 (N_8072,In_3970,In_1378);
or U8073 (N_8073,In_1783,In_4939);
xor U8074 (N_8074,In_2921,In_1390);
or U8075 (N_8075,In_826,In_1589);
nand U8076 (N_8076,In_4284,In_4778);
nor U8077 (N_8077,In_2759,In_4871);
xor U8078 (N_8078,In_4260,In_3077);
or U8079 (N_8079,In_4676,In_3430);
nor U8080 (N_8080,In_2032,In_3759);
xor U8081 (N_8081,In_1811,In_4689);
xor U8082 (N_8082,In_4293,In_4641);
nor U8083 (N_8083,In_1175,In_476);
xor U8084 (N_8084,In_4994,In_2561);
xnor U8085 (N_8085,In_785,In_3209);
nand U8086 (N_8086,In_1337,In_3683);
or U8087 (N_8087,In_2869,In_1627);
xor U8088 (N_8088,In_3185,In_4178);
and U8089 (N_8089,In_25,In_4671);
nor U8090 (N_8090,In_3862,In_3750);
nand U8091 (N_8091,In_4847,In_1940);
or U8092 (N_8092,In_1424,In_1266);
xor U8093 (N_8093,In_3394,In_2894);
nor U8094 (N_8094,In_2017,In_901);
nand U8095 (N_8095,In_3077,In_2967);
and U8096 (N_8096,In_4649,In_2471);
nand U8097 (N_8097,In_3483,In_4075);
xnor U8098 (N_8098,In_670,In_4856);
xor U8099 (N_8099,In_2534,In_2096);
and U8100 (N_8100,In_883,In_4099);
or U8101 (N_8101,In_3170,In_3252);
nand U8102 (N_8102,In_383,In_3968);
or U8103 (N_8103,In_3435,In_1536);
or U8104 (N_8104,In_4095,In_3991);
nor U8105 (N_8105,In_261,In_288);
and U8106 (N_8106,In_1004,In_4019);
nand U8107 (N_8107,In_4380,In_268);
nand U8108 (N_8108,In_745,In_3586);
nor U8109 (N_8109,In_1249,In_918);
or U8110 (N_8110,In_3749,In_3293);
nor U8111 (N_8111,In_4018,In_4856);
xor U8112 (N_8112,In_249,In_4325);
nand U8113 (N_8113,In_265,In_613);
nand U8114 (N_8114,In_4878,In_2666);
xor U8115 (N_8115,In_1011,In_3622);
xor U8116 (N_8116,In_1736,In_3799);
nand U8117 (N_8117,In_3734,In_1149);
nand U8118 (N_8118,In_1083,In_341);
nand U8119 (N_8119,In_1491,In_2464);
nand U8120 (N_8120,In_3000,In_4525);
or U8121 (N_8121,In_3319,In_4518);
and U8122 (N_8122,In_155,In_4481);
nand U8123 (N_8123,In_696,In_3961);
and U8124 (N_8124,In_328,In_2790);
and U8125 (N_8125,In_4628,In_980);
and U8126 (N_8126,In_1328,In_4033);
nand U8127 (N_8127,In_4098,In_3801);
nand U8128 (N_8128,In_3949,In_4284);
or U8129 (N_8129,In_4031,In_1579);
or U8130 (N_8130,In_353,In_4880);
xnor U8131 (N_8131,In_2828,In_2294);
or U8132 (N_8132,In_290,In_337);
nor U8133 (N_8133,In_4581,In_2114);
nand U8134 (N_8134,In_4701,In_1236);
xor U8135 (N_8135,In_2463,In_27);
or U8136 (N_8136,In_3136,In_719);
nand U8137 (N_8137,In_3106,In_2288);
or U8138 (N_8138,In_4704,In_1509);
nand U8139 (N_8139,In_1842,In_1433);
nand U8140 (N_8140,In_725,In_1400);
nor U8141 (N_8141,In_3175,In_330);
nor U8142 (N_8142,In_4116,In_3194);
or U8143 (N_8143,In_1265,In_3057);
xor U8144 (N_8144,In_3709,In_1028);
and U8145 (N_8145,In_2188,In_4375);
xnor U8146 (N_8146,In_4557,In_3619);
and U8147 (N_8147,In_1551,In_2921);
and U8148 (N_8148,In_3546,In_2855);
nand U8149 (N_8149,In_4422,In_1750);
nor U8150 (N_8150,In_3708,In_4237);
or U8151 (N_8151,In_3647,In_4135);
or U8152 (N_8152,In_4484,In_1708);
xnor U8153 (N_8153,In_720,In_2587);
nor U8154 (N_8154,In_3328,In_3332);
or U8155 (N_8155,In_2412,In_2029);
or U8156 (N_8156,In_4229,In_3288);
and U8157 (N_8157,In_3201,In_4953);
and U8158 (N_8158,In_2997,In_4474);
nand U8159 (N_8159,In_1324,In_3957);
and U8160 (N_8160,In_2288,In_4345);
xor U8161 (N_8161,In_3373,In_4418);
or U8162 (N_8162,In_1385,In_983);
nor U8163 (N_8163,In_4483,In_3086);
xnor U8164 (N_8164,In_2554,In_2658);
xor U8165 (N_8165,In_3933,In_948);
nand U8166 (N_8166,In_2587,In_3841);
or U8167 (N_8167,In_4857,In_1852);
xor U8168 (N_8168,In_1226,In_3646);
or U8169 (N_8169,In_4952,In_41);
nor U8170 (N_8170,In_1653,In_523);
or U8171 (N_8171,In_3791,In_2930);
xnor U8172 (N_8172,In_4350,In_2140);
nand U8173 (N_8173,In_3673,In_1056);
or U8174 (N_8174,In_4633,In_4157);
nand U8175 (N_8175,In_3304,In_4124);
nor U8176 (N_8176,In_4064,In_1740);
nor U8177 (N_8177,In_4431,In_2848);
nand U8178 (N_8178,In_2242,In_3143);
or U8179 (N_8179,In_2119,In_3192);
nor U8180 (N_8180,In_1337,In_4052);
nand U8181 (N_8181,In_4645,In_2675);
nand U8182 (N_8182,In_4611,In_1402);
xor U8183 (N_8183,In_3578,In_2508);
xor U8184 (N_8184,In_694,In_4312);
nand U8185 (N_8185,In_321,In_1334);
and U8186 (N_8186,In_318,In_697);
and U8187 (N_8187,In_4934,In_2123);
nor U8188 (N_8188,In_1824,In_796);
nor U8189 (N_8189,In_3295,In_2723);
and U8190 (N_8190,In_3541,In_3787);
and U8191 (N_8191,In_4971,In_4049);
xor U8192 (N_8192,In_749,In_2385);
and U8193 (N_8193,In_4215,In_180);
and U8194 (N_8194,In_3478,In_4177);
nand U8195 (N_8195,In_1703,In_3749);
xnor U8196 (N_8196,In_4005,In_4847);
nor U8197 (N_8197,In_3865,In_2474);
or U8198 (N_8198,In_3393,In_1270);
nor U8199 (N_8199,In_1087,In_4649);
xor U8200 (N_8200,In_4183,In_731);
or U8201 (N_8201,In_4727,In_950);
nand U8202 (N_8202,In_3596,In_2589);
and U8203 (N_8203,In_2299,In_3413);
nand U8204 (N_8204,In_49,In_1482);
nor U8205 (N_8205,In_3161,In_3479);
or U8206 (N_8206,In_46,In_4680);
and U8207 (N_8207,In_1786,In_311);
nand U8208 (N_8208,In_4164,In_3903);
nand U8209 (N_8209,In_2423,In_2747);
or U8210 (N_8210,In_1682,In_948);
nand U8211 (N_8211,In_939,In_3418);
nand U8212 (N_8212,In_3543,In_18);
nor U8213 (N_8213,In_678,In_3492);
xor U8214 (N_8214,In_858,In_4860);
xnor U8215 (N_8215,In_4415,In_2172);
and U8216 (N_8216,In_4788,In_3057);
xnor U8217 (N_8217,In_4099,In_11);
or U8218 (N_8218,In_167,In_670);
and U8219 (N_8219,In_4812,In_1562);
nand U8220 (N_8220,In_1965,In_141);
nand U8221 (N_8221,In_935,In_2687);
or U8222 (N_8222,In_3035,In_2591);
nor U8223 (N_8223,In_579,In_4621);
or U8224 (N_8224,In_4479,In_2920);
nor U8225 (N_8225,In_4097,In_4088);
nor U8226 (N_8226,In_2975,In_1852);
and U8227 (N_8227,In_4183,In_3473);
nor U8228 (N_8228,In_1506,In_2067);
nor U8229 (N_8229,In_2544,In_2842);
nor U8230 (N_8230,In_2708,In_4432);
nand U8231 (N_8231,In_4365,In_4326);
xnor U8232 (N_8232,In_1818,In_4301);
xor U8233 (N_8233,In_1457,In_4651);
nor U8234 (N_8234,In_4779,In_1609);
nor U8235 (N_8235,In_1219,In_1373);
and U8236 (N_8236,In_1450,In_207);
or U8237 (N_8237,In_292,In_1161);
xor U8238 (N_8238,In_1886,In_1220);
xnor U8239 (N_8239,In_1398,In_3689);
xor U8240 (N_8240,In_1376,In_4917);
nand U8241 (N_8241,In_1323,In_3456);
or U8242 (N_8242,In_3880,In_1143);
and U8243 (N_8243,In_170,In_766);
or U8244 (N_8244,In_322,In_2013);
nand U8245 (N_8245,In_1384,In_1809);
nor U8246 (N_8246,In_1214,In_4410);
or U8247 (N_8247,In_800,In_4086);
nor U8248 (N_8248,In_3752,In_2986);
and U8249 (N_8249,In_4219,In_3009);
nand U8250 (N_8250,In_264,In_4616);
xnor U8251 (N_8251,In_2418,In_4835);
or U8252 (N_8252,In_65,In_1642);
and U8253 (N_8253,In_1603,In_4829);
nand U8254 (N_8254,In_767,In_3891);
and U8255 (N_8255,In_3416,In_4661);
or U8256 (N_8256,In_556,In_3812);
xor U8257 (N_8257,In_2768,In_4799);
and U8258 (N_8258,In_4118,In_4502);
xnor U8259 (N_8259,In_3090,In_4706);
xnor U8260 (N_8260,In_3540,In_3744);
and U8261 (N_8261,In_3541,In_2956);
nand U8262 (N_8262,In_3591,In_4298);
nand U8263 (N_8263,In_2616,In_397);
nor U8264 (N_8264,In_3428,In_619);
xnor U8265 (N_8265,In_4081,In_3806);
or U8266 (N_8266,In_3230,In_2081);
or U8267 (N_8267,In_2098,In_4050);
xnor U8268 (N_8268,In_4944,In_1763);
xnor U8269 (N_8269,In_2033,In_2233);
xnor U8270 (N_8270,In_2196,In_1834);
xnor U8271 (N_8271,In_3046,In_971);
nor U8272 (N_8272,In_2438,In_3500);
nor U8273 (N_8273,In_2564,In_1709);
or U8274 (N_8274,In_3568,In_1640);
nand U8275 (N_8275,In_2199,In_2181);
and U8276 (N_8276,In_4488,In_3835);
nor U8277 (N_8277,In_1385,In_4175);
xor U8278 (N_8278,In_2979,In_1436);
or U8279 (N_8279,In_60,In_1649);
or U8280 (N_8280,In_4137,In_4549);
or U8281 (N_8281,In_3397,In_1959);
nor U8282 (N_8282,In_3680,In_94);
nor U8283 (N_8283,In_3788,In_1360);
and U8284 (N_8284,In_2632,In_1598);
and U8285 (N_8285,In_3223,In_4551);
xnor U8286 (N_8286,In_4749,In_1257);
xnor U8287 (N_8287,In_1628,In_3622);
xnor U8288 (N_8288,In_3864,In_4901);
or U8289 (N_8289,In_417,In_4207);
or U8290 (N_8290,In_259,In_2153);
and U8291 (N_8291,In_489,In_2015);
xnor U8292 (N_8292,In_2149,In_2927);
nand U8293 (N_8293,In_4701,In_2955);
or U8294 (N_8294,In_592,In_1817);
xnor U8295 (N_8295,In_1368,In_3130);
nor U8296 (N_8296,In_2798,In_4775);
and U8297 (N_8297,In_1735,In_846);
nor U8298 (N_8298,In_193,In_1049);
and U8299 (N_8299,In_4296,In_1373);
nand U8300 (N_8300,In_2016,In_4760);
and U8301 (N_8301,In_3040,In_3486);
nand U8302 (N_8302,In_4622,In_598);
or U8303 (N_8303,In_2805,In_2769);
or U8304 (N_8304,In_849,In_2165);
nor U8305 (N_8305,In_2967,In_2811);
xor U8306 (N_8306,In_1194,In_180);
nand U8307 (N_8307,In_2592,In_437);
nor U8308 (N_8308,In_1609,In_341);
nor U8309 (N_8309,In_2587,In_264);
and U8310 (N_8310,In_1357,In_4636);
or U8311 (N_8311,In_4982,In_4230);
nor U8312 (N_8312,In_2234,In_436);
nor U8313 (N_8313,In_1001,In_3895);
xnor U8314 (N_8314,In_599,In_1239);
xor U8315 (N_8315,In_2522,In_554);
or U8316 (N_8316,In_3938,In_4411);
or U8317 (N_8317,In_650,In_4466);
or U8318 (N_8318,In_3002,In_3211);
xor U8319 (N_8319,In_2253,In_3003);
and U8320 (N_8320,In_4961,In_3583);
and U8321 (N_8321,In_4703,In_898);
nand U8322 (N_8322,In_1892,In_1039);
xor U8323 (N_8323,In_3972,In_1862);
xor U8324 (N_8324,In_2876,In_2157);
nor U8325 (N_8325,In_1889,In_2794);
and U8326 (N_8326,In_2,In_1841);
nor U8327 (N_8327,In_545,In_1420);
nand U8328 (N_8328,In_2418,In_2904);
or U8329 (N_8329,In_1799,In_2693);
or U8330 (N_8330,In_3209,In_4361);
xor U8331 (N_8331,In_268,In_914);
and U8332 (N_8332,In_4835,In_1903);
nor U8333 (N_8333,In_4137,In_2524);
nor U8334 (N_8334,In_4053,In_984);
xnor U8335 (N_8335,In_2591,In_3987);
nand U8336 (N_8336,In_874,In_969);
nand U8337 (N_8337,In_413,In_3949);
and U8338 (N_8338,In_1229,In_3631);
xnor U8339 (N_8339,In_3141,In_4913);
and U8340 (N_8340,In_3036,In_1483);
nor U8341 (N_8341,In_3645,In_1386);
nor U8342 (N_8342,In_4430,In_147);
nor U8343 (N_8343,In_1519,In_1884);
nand U8344 (N_8344,In_4657,In_4568);
or U8345 (N_8345,In_1717,In_1869);
nor U8346 (N_8346,In_2301,In_2021);
and U8347 (N_8347,In_2771,In_2959);
nor U8348 (N_8348,In_2358,In_1820);
xnor U8349 (N_8349,In_1833,In_869);
xnor U8350 (N_8350,In_2248,In_2516);
nor U8351 (N_8351,In_3638,In_2043);
or U8352 (N_8352,In_4698,In_2333);
xor U8353 (N_8353,In_4186,In_2572);
and U8354 (N_8354,In_4837,In_631);
xnor U8355 (N_8355,In_4233,In_3149);
nor U8356 (N_8356,In_1982,In_659);
xnor U8357 (N_8357,In_1801,In_4783);
or U8358 (N_8358,In_519,In_1091);
or U8359 (N_8359,In_4616,In_2943);
nand U8360 (N_8360,In_244,In_3543);
xor U8361 (N_8361,In_641,In_3282);
and U8362 (N_8362,In_4944,In_3800);
or U8363 (N_8363,In_3893,In_166);
and U8364 (N_8364,In_862,In_240);
and U8365 (N_8365,In_2953,In_4620);
and U8366 (N_8366,In_320,In_2927);
nor U8367 (N_8367,In_1604,In_127);
nor U8368 (N_8368,In_1764,In_4728);
xor U8369 (N_8369,In_3035,In_3852);
or U8370 (N_8370,In_2614,In_1772);
nor U8371 (N_8371,In_890,In_4163);
and U8372 (N_8372,In_2132,In_3441);
xor U8373 (N_8373,In_4699,In_3266);
nor U8374 (N_8374,In_3348,In_32);
and U8375 (N_8375,In_3949,In_1206);
xor U8376 (N_8376,In_2195,In_822);
nand U8377 (N_8377,In_2935,In_453);
nor U8378 (N_8378,In_2607,In_2479);
and U8379 (N_8379,In_2106,In_4122);
and U8380 (N_8380,In_2587,In_4387);
and U8381 (N_8381,In_4218,In_2981);
or U8382 (N_8382,In_233,In_562);
nor U8383 (N_8383,In_4952,In_974);
nor U8384 (N_8384,In_1620,In_450);
xnor U8385 (N_8385,In_3458,In_583);
and U8386 (N_8386,In_225,In_4265);
or U8387 (N_8387,In_3156,In_3195);
nor U8388 (N_8388,In_2520,In_1393);
and U8389 (N_8389,In_4720,In_3068);
and U8390 (N_8390,In_2672,In_663);
or U8391 (N_8391,In_389,In_771);
and U8392 (N_8392,In_377,In_2223);
xor U8393 (N_8393,In_4691,In_4186);
nand U8394 (N_8394,In_140,In_2230);
xor U8395 (N_8395,In_2401,In_3393);
nor U8396 (N_8396,In_3958,In_974);
or U8397 (N_8397,In_2173,In_2277);
nand U8398 (N_8398,In_284,In_3053);
or U8399 (N_8399,In_3869,In_541);
nor U8400 (N_8400,In_2590,In_4606);
xor U8401 (N_8401,In_131,In_833);
nor U8402 (N_8402,In_4884,In_4659);
nand U8403 (N_8403,In_4253,In_671);
and U8404 (N_8404,In_1256,In_657);
or U8405 (N_8405,In_3838,In_4785);
or U8406 (N_8406,In_4147,In_1447);
and U8407 (N_8407,In_4115,In_643);
xor U8408 (N_8408,In_2448,In_1535);
and U8409 (N_8409,In_165,In_2999);
xnor U8410 (N_8410,In_3618,In_3848);
nor U8411 (N_8411,In_2663,In_4894);
xor U8412 (N_8412,In_1466,In_4730);
nor U8413 (N_8413,In_4605,In_3346);
xnor U8414 (N_8414,In_3805,In_4980);
nand U8415 (N_8415,In_1668,In_3153);
or U8416 (N_8416,In_2153,In_394);
nand U8417 (N_8417,In_966,In_2994);
nand U8418 (N_8418,In_3642,In_2481);
nand U8419 (N_8419,In_1289,In_1166);
or U8420 (N_8420,In_4949,In_1503);
xor U8421 (N_8421,In_4215,In_4207);
nand U8422 (N_8422,In_4776,In_532);
or U8423 (N_8423,In_3631,In_4034);
and U8424 (N_8424,In_4745,In_4997);
and U8425 (N_8425,In_4421,In_2533);
nor U8426 (N_8426,In_2834,In_3952);
nand U8427 (N_8427,In_4564,In_2894);
and U8428 (N_8428,In_4499,In_1833);
and U8429 (N_8429,In_840,In_3559);
or U8430 (N_8430,In_365,In_1233);
xor U8431 (N_8431,In_218,In_2849);
and U8432 (N_8432,In_1246,In_422);
and U8433 (N_8433,In_2448,In_1900);
xnor U8434 (N_8434,In_4658,In_336);
nor U8435 (N_8435,In_2326,In_2827);
and U8436 (N_8436,In_4789,In_4013);
or U8437 (N_8437,In_1982,In_4138);
nor U8438 (N_8438,In_385,In_4676);
or U8439 (N_8439,In_1107,In_2734);
and U8440 (N_8440,In_458,In_4518);
nand U8441 (N_8441,In_3336,In_3574);
nand U8442 (N_8442,In_2169,In_756);
nor U8443 (N_8443,In_4717,In_2681);
xor U8444 (N_8444,In_1067,In_2343);
and U8445 (N_8445,In_1135,In_4043);
nor U8446 (N_8446,In_2552,In_3710);
xor U8447 (N_8447,In_4716,In_3142);
nand U8448 (N_8448,In_2957,In_4146);
xor U8449 (N_8449,In_1149,In_37);
xnor U8450 (N_8450,In_3717,In_3287);
or U8451 (N_8451,In_3137,In_3294);
nor U8452 (N_8452,In_685,In_4849);
or U8453 (N_8453,In_3907,In_3250);
xor U8454 (N_8454,In_476,In_2897);
or U8455 (N_8455,In_2252,In_4504);
xor U8456 (N_8456,In_370,In_3208);
nor U8457 (N_8457,In_75,In_2051);
or U8458 (N_8458,In_228,In_2547);
xor U8459 (N_8459,In_4526,In_1796);
nor U8460 (N_8460,In_3440,In_2539);
nand U8461 (N_8461,In_1901,In_2307);
nor U8462 (N_8462,In_3744,In_3882);
nor U8463 (N_8463,In_1843,In_565);
nand U8464 (N_8464,In_798,In_785);
nand U8465 (N_8465,In_4381,In_865);
and U8466 (N_8466,In_848,In_3876);
nand U8467 (N_8467,In_612,In_514);
and U8468 (N_8468,In_749,In_1841);
and U8469 (N_8469,In_2391,In_4623);
or U8470 (N_8470,In_2065,In_4310);
or U8471 (N_8471,In_775,In_603);
xnor U8472 (N_8472,In_1099,In_2281);
and U8473 (N_8473,In_3485,In_3830);
xnor U8474 (N_8474,In_3168,In_2017);
or U8475 (N_8475,In_491,In_926);
and U8476 (N_8476,In_2865,In_4002);
nor U8477 (N_8477,In_2241,In_2560);
and U8478 (N_8478,In_4146,In_3717);
or U8479 (N_8479,In_168,In_2943);
xnor U8480 (N_8480,In_4621,In_1637);
and U8481 (N_8481,In_4463,In_1335);
and U8482 (N_8482,In_4231,In_3467);
nand U8483 (N_8483,In_2356,In_541);
nand U8484 (N_8484,In_2364,In_586);
nand U8485 (N_8485,In_156,In_4746);
nor U8486 (N_8486,In_3446,In_44);
nor U8487 (N_8487,In_4683,In_1316);
or U8488 (N_8488,In_3732,In_1915);
and U8489 (N_8489,In_746,In_1489);
or U8490 (N_8490,In_1855,In_2021);
nand U8491 (N_8491,In_3582,In_4903);
nor U8492 (N_8492,In_2613,In_1230);
or U8493 (N_8493,In_3502,In_4736);
and U8494 (N_8494,In_2662,In_317);
nor U8495 (N_8495,In_3601,In_4196);
or U8496 (N_8496,In_18,In_725);
or U8497 (N_8497,In_1421,In_2678);
xnor U8498 (N_8498,In_1107,In_649);
and U8499 (N_8499,In_2488,In_639);
nand U8500 (N_8500,In_2033,In_50);
xnor U8501 (N_8501,In_4835,In_1889);
xnor U8502 (N_8502,In_2764,In_2990);
xnor U8503 (N_8503,In_3414,In_2255);
nor U8504 (N_8504,In_3125,In_1681);
nand U8505 (N_8505,In_2132,In_1684);
or U8506 (N_8506,In_2090,In_2958);
and U8507 (N_8507,In_1906,In_4118);
nand U8508 (N_8508,In_3925,In_4397);
and U8509 (N_8509,In_3014,In_2301);
xor U8510 (N_8510,In_2188,In_3300);
or U8511 (N_8511,In_3936,In_1842);
nand U8512 (N_8512,In_298,In_2479);
nor U8513 (N_8513,In_2353,In_2523);
nand U8514 (N_8514,In_2050,In_1289);
xnor U8515 (N_8515,In_4892,In_4729);
or U8516 (N_8516,In_1374,In_1522);
xnor U8517 (N_8517,In_1689,In_2686);
and U8518 (N_8518,In_198,In_2985);
nor U8519 (N_8519,In_3051,In_1424);
and U8520 (N_8520,In_3665,In_979);
nor U8521 (N_8521,In_3778,In_3887);
xnor U8522 (N_8522,In_1753,In_2887);
nor U8523 (N_8523,In_3529,In_2920);
and U8524 (N_8524,In_510,In_4269);
xor U8525 (N_8525,In_3718,In_3434);
and U8526 (N_8526,In_4940,In_343);
nand U8527 (N_8527,In_3480,In_1011);
or U8528 (N_8528,In_3424,In_1060);
nor U8529 (N_8529,In_2080,In_2194);
nand U8530 (N_8530,In_4743,In_2964);
xor U8531 (N_8531,In_3145,In_1775);
nor U8532 (N_8532,In_2603,In_2440);
xor U8533 (N_8533,In_4250,In_3461);
xor U8534 (N_8534,In_54,In_2225);
nand U8535 (N_8535,In_1028,In_4513);
xor U8536 (N_8536,In_3692,In_3382);
or U8537 (N_8537,In_975,In_2318);
xnor U8538 (N_8538,In_2624,In_4342);
xnor U8539 (N_8539,In_1781,In_891);
xnor U8540 (N_8540,In_371,In_2817);
and U8541 (N_8541,In_4332,In_3615);
nor U8542 (N_8542,In_4093,In_3665);
nand U8543 (N_8543,In_320,In_3546);
xnor U8544 (N_8544,In_3773,In_1313);
or U8545 (N_8545,In_2946,In_1627);
and U8546 (N_8546,In_549,In_3268);
nand U8547 (N_8547,In_21,In_3812);
or U8548 (N_8548,In_2485,In_858);
nor U8549 (N_8549,In_2444,In_1329);
and U8550 (N_8550,In_3712,In_68);
nor U8551 (N_8551,In_3219,In_3472);
xnor U8552 (N_8552,In_2285,In_788);
nand U8553 (N_8553,In_1124,In_2769);
and U8554 (N_8554,In_4192,In_4679);
and U8555 (N_8555,In_3941,In_2964);
nor U8556 (N_8556,In_4909,In_4296);
and U8557 (N_8557,In_1715,In_4949);
or U8558 (N_8558,In_2487,In_294);
or U8559 (N_8559,In_3570,In_2859);
nor U8560 (N_8560,In_4763,In_3322);
xnor U8561 (N_8561,In_2050,In_3470);
nor U8562 (N_8562,In_3849,In_3497);
nand U8563 (N_8563,In_2081,In_2748);
nor U8564 (N_8564,In_1579,In_3727);
or U8565 (N_8565,In_63,In_2198);
nand U8566 (N_8566,In_4084,In_2735);
nor U8567 (N_8567,In_2921,In_363);
and U8568 (N_8568,In_1452,In_586);
xnor U8569 (N_8569,In_2781,In_2619);
or U8570 (N_8570,In_2468,In_1390);
xnor U8571 (N_8571,In_2927,In_362);
xnor U8572 (N_8572,In_2118,In_1026);
or U8573 (N_8573,In_103,In_2046);
nor U8574 (N_8574,In_2500,In_2854);
xor U8575 (N_8575,In_4997,In_4607);
xor U8576 (N_8576,In_3949,In_3480);
nand U8577 (N_8577,In_614,In_105);
xnor U8578 (N_8578,In_1734,In_4020);
nand U8579 (N_8579,In_4301,In_3713);
and U8580 (N_8580,In_4938,In_794);
nor U8581 (N_8581,In_2075,In_3335);
nor U8582 (N_8582,In_2768,In_416);
xnor U8583 (N_8583,In_3868,In_2077);
nand U8584 (N_8584,In_1690,In_2190);
or U8585 (N_8585,In_3026,In_3692);
and U8586 (N_8586,In_553,In_3089);
xnor U8587 (N_8587,In_1124,In_280);
nand U8588 (N_8588,In_3887,In_561);
or U8589 (N_8589,In_2038,In_4779);
and U8590 (N_8590,In_2817,In_2539);
nor U8591 (N_8591,In_3204,In_3425);
or U8592 (N_8592,In_2196,In_4632);
nor U8593 (N_8593,In_3848,In_4783);
and U8594 (N_8594,In_746,In_1363);
xor U8595 (N_8595,In_3491,In_2446);
and U8596 (N_8596,In_3930,In_3663);
nor U8597 (N_8597,In_1906,In_4099);
nor U8598 (N_8598,In_431,In_4234);
nor U8599 (N_8599,In_3303,In_35);
xnor U8600 (N_8600,In_2584,In_4499);
nor U8601 (N_8601,In_4266,In_151);
xor U8602 (N_8602,In_487,In_2414);
xor U8603 (N_8603,In_3998,In_1285);
xor U8604 (N_8604,In_2311,In_1583);
xor U8605 (N_8605,In_2472,In_337);
nor U8606 (N_8606,In_1435,In_1386);
and U8607 (N_8607,In_4922,In_3872);
nor U8608 (N_8608,In_559,In_1053);
nor U8609 (N_8609,In_245,In_4440);
and U8610 (N_8610,In_198,In_1979);
nor U8611 (N_8611,In_188,In_3497);
and U8612 (N_8612,In_4034,In_1264);
and U8613 (N_8613,In_2581,In_431);
nor U8614 (N_8614,In_3146,In_3308);
nor U8615 (N_8615,In_4971,In_4702);
nand U8616 (N_8616,In_3588,In_1224);
and U8617 (N_8617,In_1274,In_4004);
nor U8618 (N_8618,In_2891,In_1958);
and U8619 (N_8619,In_291,In_2342);
and U8620 (N_8620,In_3709,In_1773);
nand U8621 (N_8621,In_856,In_141);
and U8622 (N_8622,In_3665,In_4234);
and U8623 (N_8623,In_1670,In_737);
xor U8624 (N_8624,In_2932,In_3630);
and U8625 (N_8625,In_2283,In_2391);
and U8626 (N_8626,In_2739,In_1221);
or U8627 (N_8627,In_4004,In_4223);
nand U8628 (N_8628,In_2643,In_4712);
and U8629 (N_8629,In_1723,In_1817);
nor U8630 (N_8630,In_1414,In_1473);
nor U8631 (N_8631,In_3905,In_2451);
or U8632 (N_8632,In_2204,In_2301);
nor U8633 (N_8633,In_3520,In_562);
or U8634 (N_8634,In_3922,In_3938);
xnor U8635 (N_8635,In_1140,In_806);
and U8636 (N_8636,In_2856,In_4810);
and U8637 (N_8637,In_3048,In_1745);
or U8638 (N_8638,In_2348,In_1385);
or U8639 (N_8639,In_398,In_1550);
nor U8640 (N_8640,In_4108,In_1263);
nand U8641 (N_8641,In_805,In_4241);
xor U8642 (N_8642,In_2910,In_2095);
or U8643 (N_8643,In_4505,In_944);
nand U8644 (N_8644,In_1775,In_1408);
nand U8645 (N_8645,In_1926,In_3508);
xor U8646 (N_8646,In_1892,In_1178);
xnor U8647 (N_8647,In_3444,In_174);
nand U8648 (N_8648,In_4074,In_2917);
nor U8649 (N_8649,In_1991,In_1132);
nor U8650 (N_8650,In_4903,In_629);
nor U8651 (N_8651,In_1280,In_4414);
and U8652 (N_8652,In_2097,In_4811);
xnor U8653 (N_8653,In_2461,In_8);
or U8654 (N_8654,In_165,In_4230);
or U8655 (N_8655,In_1628,In_1992);
nand U8656 (N_8656,In_4348,In_4734);
nor U8657 (N_8657,In_3459,In_2074);
nor U8658 (N_8658,In_4021,In_3933);
nand U8659 (N_8659,In_2226,In_341);
or U8660 (N_8660,In_4786,In_1224);
xor U8661 (N_8661,In_267,In_1555);
and U8662 (N_8662,In_4778,In_4535);
or U8663 (N_8663,In_3350,In_2075);
or U8664 (N_8664,In_4519,In_2693);
or U8665 (N_8665,In_1786,In_2236);
xor U8666 (N_8666,In_651,In_1984);
and U8667 (N_8667,In_1934,In_3099);
nor U8668 (N_8668,In_3195,In_1443);
nor U8669 (N_8669,In_2664,In_2773);
nand U8670 (N_8670,In_200,In_2002);
xnor U8671 (N_8671,In_196,In_3698);
and U8672 (N_8672,In_1836,In_4766);
nand U8673 (N_8673,In_1473,In_3384);
and U8674 (N_8674,In_3093,In_851);
nand U8675 (N_8675,In_1475,In_270);
xor U8676 (N_8676,In_3759,In_988);
nand U8677 (N_8677,In_183,In_1237);
nor U8678 (N_8678,In_2292,In_4923);
or U8679 (N_8679,In_4334,In_2043);
nor U8680 (N_8680,In_1128,In_3455);
nor U8681 (N_8681,In_2306,In_2657);
and U8682 (N_8682,In_3350,In_3324);
nand U8683 (N_8683,In_2649,In_2887);
or U8684 (N_8684,In_2004,In_4287);
nand U8685 (N_8685,In_3947,In_2104);
or U8686 (N_8686,In_4536,In_3599);
and U8687 (N_8687,In_1569,In_2270);
or U8688 (N_8688,In_4759,In_4463);
nand U8689 (N_8689,In_4328,In_238);
nor U8690 (N_8690,In_3995,In_4268);
nand U8691 (N_8691,In_1228,In_1838);
nand U8692 (N_8692,In_1453,In_883);
nand U8693 (N_8693,In_2764,In_2721);
and U8694 (N_8694,In_3487,In_3195);
nand U8695 (N_8695,In_758,In_548);
nand U8696 (N_8696,In_4128,In_4447);
or U8697 (N_8697,In_1537,In_2246);
nor U8698 (N_8698,In_3122,In_982);
or U8699 (N_8699,In_4377,In_1367);
nand U8700 (N_8700,In_721,In_720);
or U8701 (N_8701,In_32,In_3195);
nand U8702 (N_8702,In_1268,In_2286);
or U8703 (N_8703,In_335,In_2352);
xor U8704 (N_8704,In_4272,In_821);
nand U8705 (N_8705,In_3510,In_4607);
nor U8706 (N_8706,In_4064,In_3716);
xnor U8707 (N_8707,In_2326,In_3691);
or U8708 (N_8708,In_3361,In_4104);
or U8709 (N_8709,In_3993,In_670);
nor U8710 (N_8710,In_4407,In_2766);
nor U8711 (N_8711,In_165,In_4895);
nor U8712 (N_8712,In_1966,In_2782);
or U8713 (N_8713,In_4588,In_3482);
nand U8714 (N_8714,In_18,In_295);
and U8715 (N_8715,In_3904,In_1609);
or U8716 (N_8716,In_963,In_2924);
xnor U8717 (N_8717,In_3990,In_3877);
xor U8718 (N_8718,In_3743,In_4799);
nand U8719 (N_8719,In_2301,In_1822);
or U8720 (N_8720,In_1297,In_1561);
nand U8721 (N_8721,In_3653,In_4573);
nand U8722 (N_8722,In_2532,In_3938);
and U8723 (N_8723,In_4344,In_1462);
nand U8724 (N_8724,In_667,In_2070);
nand U8725 (N_8725,In_865,In_1827);
and U8726 (N_8726,In_996,In_1239);
or U8727 (N_8727,In_4432,In_3201);
nand U8728 (N_8728,In_3213,In_3198);
nand U8729 (N_8729,In_3973,In_4774);
or U8730 (N_8730,In_39,In_3116);
nor U8731 (N_8731,In_1575,In_2035);
or U8732 (N_8732,In_3273,In_1037);
nand U8733 (N_8733,In_4666,In_2808);
or U8734 (N_8734,In_345,In_485);
nand U8735 (N_8735,In_2792,In_2439);
or U8736 (N_8736,In_874,In_1070);
and U8737 (N_8737,In_4185,In_1150);
nor U8738 (N_8738,In_2250,In_3375);
and U8739 (N_8739,In_67,In_4129);
and U8740 (N_8740,In_2289,In_1040);
nand U8741 (N_8741,In_3696,In_2348);
and U8742 (N_8742,In_2921,In_2145);
and U8743 (N_8743,In_3396,In_3342);
xnor U8744 (N_8744,In_978,In_2940);
and U8745 (N_8745,In_4476,In_1280);
and U8746 (N_8746,In_578,In_3814);
xor U8747 (N_8747,In_3527,In_4023);
or U8748 (N_8748,In_2161,In_3279);
nand U8749 (N_8749,In_3064,In_3928);
nor U8750 (N_8750,In_2849,In_868);
nor U8751 (N_8751,In_2595,In_1574);
or U8752 (N_8752,In_1909,In_919);
xor U8753 (N_8753,In_1052,In_3919);
or U8754 (N_8754,In_2180,In_745);
nand U8755 (N_8755,In_275,In_3328);
xor U8756 (N_8756,In_850,In_1342);
nor U8757 (N_8757,In_3763,In_1954);
nor U8758 (N_8758,In_1103,In_3874);
or U8759 (N_8759,In_1702,In_3094);
nor U8760 (N_8760,In_4801,In_4154);
nand U8761 (N_8761,In_1822,In_4240);
xnor U8762 (N_8762,In_300,In_3676);
nand U8763 (N_8763,In_1244,In_967);
and U8764 (N_8764,In_3517,In_4921);
and U8765 (N_8765,In_2248,In_1737);
and U8766 (N_8766,In_1127,In_1338);
nand U8767 (N_8767,In_28,In_3062);
xor U8768 (N_8768,In_976,In_3427);
and U8769 (N_8769,In_537,In_3169);
xnor U8770 (N_8770,In_2322,In_4638);
nand U8771 (N_8771,In_254,In_979);
and U8772 (N_8772,In_2699,In_4412);
nand U8773 (N_8773,In_3176,In_1756);
and U8774 (N_8774,In_434,In_4011);
or U8775 (N_8775,In_942,In_757);
xor U8776 (N_8776,In_3666,In_1330);
nor U8777 (N_8777,In_120,In_819);
nor U8778 (N_8778,In_121,In_4223);
or U8779 (N_8779,In_92,In_2109);
nand U8780 (N_8780,In_4938,In_3698);
nor U8781 (N_8781,In_183,In_1595);
xnor U8782 (N_8782,In_4877,In_805);
xnor U8783 (N_8783,In_4181,In_2004);
nor U8784 (N_8784,In_4489,In_517);
xor U8785 (N_8785,In_3131,In_3640);
nor U8786 (N_8786,In_1355,In_3494);
nand U8787 (N_8787,In_1874,In_1483);
and U8788 (N_8788,In_4448,In_345);
or U8789 (N_8789,In_2000,In_4585);
nor U8790 (N_8790,In_4506,In_3278);
and U8791 (N_8791,In_4594,In_3643);
and U8792 (N_8792,In_4016,In_1643);
nor U8793 (N_8793,In_1880,In_269);
or U8794 (N_8794,In_1393,In_4052);
nor U8795 (N_8795,In_1435,In_4893);
nor U8796 (N_8796,In_3524,In_1991);
and U8797 (N_8797,In_4641,In_3113);
xnor U8798 (N_8798,In_4354,In_4072);
nand U8799 (N_8799,In_438,In_3896);
nand U8800 (N_8800,In_820,In_4915);
nand U8801 (N_8801,In_33,In_1951);
or U8802 (N_8802,In_4326,In_785);
nor U8803 (N_8803,In_1658,In_1406);
nor U8804 (N_8804,In_4554,In_1770);
xor U8805 (N_8805,In_2281,In_3636);
or U8806 (N_8806,In_1899,In_4735);
nor U8807 (N_8807,In_4749,In_4808);
or U8808 (N_8808,In_512,In_4090);
nand U8809 (N_8809,In_3388,In_4511);
nand U8810 (N_8810,In_1866,In_2666);
or U8811 (N_8811,In_543,In_1120);
nor U8812 (N_8812,In_3052,In_2861);
nor U8813 (N_8813,In_565,In_825);
or U8814 (N_8814,In_2686,In_732);
or U8815 (N_8815,In_3669,In_2626);
and U8816 (N_8816,In_355,In_3841);
nor U8817 (N_8817,In_3760,In_1255);
nor U8818 (N_8818,In_2982,In_2955);
nor U8819 (N_8819,In_3996,In_4818);
and U8820 (N_8820,In_2723,In_4507);
xnor U8821 (N_8821,In_2227,In_3152);
nor U8822 (N_8822,In_3501,In_1240);
and U8823 (N_8823,In_1929,In_3331);
xor U8824 (N_8824,In_4423,In_4517);
xnor U8825 (N_8825,In_2038,In_3436);
xnor U8826 (N_8826,In_4595,In_3407);
xor U8827 (N_8827,In_3983,In_1145);
nand U8828 (N_8828,In_1983,In_3247);
and U8829 (N_8829,In_4494,In_2117);
nand U8830 (N_8830,In_390,In_1284);
and U8831 (N_8831,In_1391,In_2540);
nor U8832 (N_8832,In_1501,In_577);
and U8833 (N_8833,In_751,In_116);
nand U8834 (N_8834,In_3457,In_1576);
nand U8835 (N_8835,In_1474,In_1256);
nand U8836 (N_8836,In_4829,In_3175);
nand U8837 (N_8837,In_880,In_4032);
nand U8838 (N_8838,In_2528,In_2974);
xor U8839 (N_8839,In_1472,In_2921);
xnor U8840 (N_8840,In_1898,In_2079);
or U8841 (N_8841,In_4429,In_136);
xor U8842 (N_8842,In_4795,In_3342);
nor U8843 (N_8843,In_1466,In_4857);
nor U8844 (N_8844,In_29,In_4714);
and U8845 (N_8845,In_1411,In_3935);
and U8846 (N_8846,In_91,In_4141);
xnor U8847 (N_8847,In_1634,In_4030);
xor U8848 (N_8848,In_4331,In_206);
nand U8849 (N_8849,In_4334,In_145);
and U8850 (N_8850,In_1376,In_2414);
nand U8851 (N_8851,In_4029,In_1581);
and U8852 (N_8852,In_3527,In_2594);
and U8853 (N_8853,In_90,In_1332);
nand U8854 (N_8854,In_1259,In_2557);
xor U8855 (N_8855,In_1236,In_633);
nor U8856 (N_8856,In_3927,In_2277);
or U8857 (N_8857,In_4815,In_1905);
nand U8858 (N_8858,In_2817,In_2918);
nor U8859 (N_8859,In_27,In_4406);
and U8860 (N_8860,In_802,In_858);
or U8861 (N_8861,In_3463,In_1130);
nand U8862 (N_8862,In_4753,In_4924);
xnor U8863 (N_8863,In_2603,In_70);
nand U8864 (N_8864,In_885,In_2494);
nand U8865 (N_8865,In_2408,In_1631);
and U8866 (N_8866,In_3073,In_4833);
or U8867 (N_8867,In_793,In_2068);
or U8868 (N_8868,In_1695,In_3776);
nand U8869 (N_8869,In_1363,In_1592);
nor U8870 (N_8870,In_658,In_2492);
nor U8871 (N_8871,In_3044,In_4664);
or U8872 (N_8872,In_1376,In_2966);
xnor U8873 (N_8873,In_3747,In_534);
or U8874 (N_8874,In_3138,In_2729);
nor U8875 (N_8875,In_4029,In_3313);
and U8876 (N_8876,In_1204,In_679);
and U8877 (N_8877,In_92,In_298);
nor U8878 (N_8878,In_3454,In_4998);
or U8879 (N_8879,In_2709,In_1164);
and U8880 (N_8880,In_1413,In_4720);
or U8881 (N_8881,In_1908,In_2126);
and U8882 (N_8882,In_4981,In_1330);
and U8883 (N_8883,In_28,In_4058);
or U8884 (N_8884,In_3037,In_3596);
xor U8885 (N_8885,In_4188,In_1686);
and U8886 (N_8886,In_2011,In_1630);
nand U8887 (N_8887,In_2887,In_3841);
or U8888 (N_8888,In_4831,In_852);
or U8889 (N_8889,In_2205,In_4948);
nor U8890 (N_8890,In_1295,In_470);
and U8891 (N_8891,In_3216,In_1076);
and U8892 (N_8892,In_990,In_4309);
nor U8893 (N_8893,In_1314,In_1200);
nor U8894 (N_8894,In_4565,In_2041);
xor U8895 (N_8895,In_3067,In_4741);
nor U8896 (N_8896,In_2889,In_1724);
and U8897 (N_8897,In_4835,In_2488);
nor U8898 (N_8898,In_3922,In_2646);
and U8899 (N_8899,In_556,In_1385);
xor U8900 (N_8900,In_2933,In_3249);
xor U8901 (N_8901,In_174,In_591);
or U8902 (N_8902,In_4554,In_4927);
and U8903 (N_8903,In_3582,In_4567);
nor U8904 (N_8904,In_217,In_1834);
nor U8905 (N_8905,In_159,In_2368);
nand U8906 (N_8906,In_3890,In_1137);
and U8907 (N_8907,In_2048,In_2022);
nand U8908 (N_8908,In_245,In_1075);
and U8909 (N_8909,In_4818,In_2632);
nor U8910 (N_8910,In_3444,In_1068);
xnor U8911 (N_8911,In_1290,In_3428);
xnor U8912 (N_8912,In_2767,In_1991);
xor U8913 (N_8913,In_2917,In_3189);
xor U8914 (N_8914,In_1083,In_2310);
or U8915 (N_8915,In_4834,In_1749);
nand U8916 (N_8916,In_1980,In_977);
xnor U8917 (N_8917,In_2030,In_1672);
nor U8918 (N_8918,In_2325,In_4165);
nor U8919 (N_8919,In_2170,In_2683);
nand U8920 (N_8920,In_4328,In_114);
nand U8921 (N_8921,In_1693,In_3209);
xor U8922 (N_8922,In_1700,In_1649);
nor U8923 (N_8923,In_897,In_2847);
xnor U8924 (N_8924,In_1652,In_4730);
or U8925 (N_8925,In_705,In_788);
xnor U8926 (N_8926,In_1276,In_2796);
xnor U8927 (N_8927,In_1953,In_4367);
or U8928 (N_8928,In_3234,In_4362);
xnor U8929 (N_8929,In_3730,In_600);
nor U8930 (N_8930,In_1558,In_3291);
nor U8931 (N_8931,In_527,In_1866);
and U8932 (N_8932,In_4915,In_4890);
and U8933 (N_8933,In_3426,In_2898);
xnor U8934 (N_8934,In_3625,In_4507);
xnor U8935 (N_8935,In_4750,In_1174);
and U8936 (N_8936,In_3873,In_2184);
nor U8937 (N_8937,In_3730,In_4108);
nand U8938 (N_8938,In_2545,In_3840);
nand U8939 (N_8939,In_3530,In_1816);
or U8940 (N_8940,In_997,In_851);
nand U8941 (N_8941,In_4858,In_3622);
nor U8942 (N_8942,In_3268,In_169);
nand U8943 (N_8943,In_771,In_333);
or U8944 (N_8944,In_4512,In_3256);
or U8945 (N_8945,In_3461,In_4836);
nand U8946 (N_8946,In_827,In_2208);
xor U8947 (N_8947,In_175,In_3811);
and U8948 (N_8948,In_2936,In_1120);
nor U8949 (N_8949,In_4171,In_3038);
nand U8950 (N_8950,In_4011,In_4001);
xnor U8951 (N_8951,In_512,In_3188);
nand U8952 (N_8952,In_3837,In_787);
and U8953 (N_8953,In_1868,In_4121);
xor U8954 (N_8954,In_2659,In_381);
xnor U8955 (N_8955,In_1750,In_3805);
xnor U8956 (N_8956,In_2985,In_2371);
or U8957 (N_8957,In_264,In_706);
or U8958 (N_8958,In_4500,In_3172);
or U8959 (N_8959,In_464,In_3789);
and U8960 (N_8960,In_3316,In_1324);
xnor U8961 (N_8961,In_1706,In_3088);
and U8962 (N_8962,In_3950,In_4084);
and U8963 (N_8963,In_2423,In_1153);
nand U8964 (N_8964,In_1296,In_583);
xnor U8965 (N_8965,In_4612,In_595);
xor U8966 (N_8966,In_1859,In_995);
or U8967 (N_8967,In_330,In_3459);
and U8968 (N_8968,In_2418,In_73);
nor U8969 (N_8969,In_2078,In_269);
xor U8970 (N_8970,In_2326,In_1043);
and U8971 (N_8971,In_1417,In_1486);
nand U8972 (N_8972,In_834,In_1765);
xor U8973 (N_8973,In_360,In_1274);
nand U8974 (N_8974,In_4120,In_2510);
or U8975 (N_8975,In_3220,In_252);
xor U8976 (N_8976,In_4521,In_860);
and U8977 (N_8977,In_2443,In_3042);
nand U8978 (N_8978,In_4589,In_150);
xor U8979 (N_8979,In_1493,In_1415);
nor U8980 (N_8980,In_2633,In_308);
nor U8981 (N_8981,In_701,In_233);
xnor U8982 (N_8982,In_383,In_2976);
nand U8983 (N_8983,In_4060,In_3909);
and U8984 (N_8984,In_1666,In_976);
nor U8985 (N_8985,In_3724,In_310);
nor U8986 (N_8986,In_4018,In_3049);
nand U8987 (N_8987,In_2599,In_239);
nor U8988 (N_8988,In_1166,In_2852);
xor U8989 (N_8989,In_1465,In_3971);
and U8990 (N_8990,In_2892,In_3287);
xor U8991 (N_8991,In_2186,In_3618);
nand U8992 (N_8992,In_142,In_758);
nand U8993 (N_8993,In_1709,In_2171);
nor U8994 (N_8994,In_3047,In_4856);
xor U8995 (N_8995,In_3803,In_2016);
xnor U8996 (N_8996,In_4789,In_1740);
nand U8997 (N_8997,In_3461,In_3417);
xnor U8998 (N_8998,In_4891,In_4664);
nor U8999 (N_8999,In_1750,In_2327);
xor U9000 (N_9000,In_2118,In_3372);
xor U9001 (N_9001,In_1418,In_823);
nand U9002 (N_9002,In_3547,In_1903);
xnor U9003 (N_9003,In_3647,In_3009);
nand U9004 (N_9004,In_4350,In_1836);
or U9005 (N_9005,In_3107,In_3454);
and U9006 (N_9006,In_3273,In_684);
and U9007 (N_9007,In_1527,In_3381);
nand U9008 (N_9008,In_339,In_3606);
or U9009 (N_9009,In_2388,In_3349);
and U9010 (N_9010,In_2670,In_2545);
or U9011 (N_9011,In_3945,In_1999);
nand U9012 (N_9012,In_3966,In_1693);
or U9013 (N_9013,In_979,In_4934);
and U9014 (N_9014,In_13,In_44);
xor U9015 (N_9015,In_2155,In_12);
and U9016 (N_9016,In_2429,In_3354);
and U9017 (N_9017,In_2683,In_4227);
nor U9018 (N_9018,In_2926,In_3574);
xnor U9019 (N_9019,In_1878,In_4700);
nor U9020 (N_9020,In_4505,In_2115);
xor U9021 (N_9021,In_3731,In_4481);
nor U9022 (N_9022,In_1265,In_123);
xnor U9023 (N_9023,In_2055,In_2186);
nand U9024 (N_9024,In_4551,In_3599);
and U9025 (N_9025,In_4163,In_804);
nand U9026 (N_9026,In_234,In_1706);
or U9027 (N_9027,In_1007,In_3269);
nand U9028 (N_9028,In_4484,In_3129);
xnor U9029 (N_9029,In_3358,In_2916);
nand U9030 (N_9030,In_2482,In_1055);
nand U9031 (N_9031,In_1480,In_3630);
xnor U9032 (N_9032,In_3365,In_4414);
xnor U9033 (N_9033,In_4665,In_4197);
xor U9034 (N_9034,In_3364,In_2651);
and U9035 (N_9035,In_1238,In_3070);
or U9036 (N_9036,In_3688,In_2874);
nand U9037 (N_9037,In_4207,In_764);
and U9038 (N_9038,In_855,In_3850);
or U9039 (N_9039,In_1094,In_1142);
or U9040 (N_9040,In_24,In_2581);
xor U9041 (N_9041,In_2114,In_2853);
nand U9042 (N_9042,In_417,In_4901);
and U9043 (N_9043,In_4707,In_3000);
xnor U9044 (N_9044,In_510,In_1642);
and U9045 (N_9045,In_3912,In_4612);
and U9046 (N_9046,In_1022,In_2740);
xnor U9047 (N_9047,In_1053,In_2522);
xnor U9048 (N_9048,In_3957,In_2698);
or U9049 (N_9049,In_1899,In_3420);
nor U9050 (N_9050,In_1027,In_3465);
nor U9051 (N_9051,In_1125,In_639);
nor U9052 (N_9052,In_4112,In_1833);
and U9053 (N_9053,In_1369,In_1929);
nor U9054 (N_9054,In_4932,In_628);
and U9055 (N_9055,In_2148,In_2482);
or U9056 (N_9056,In_1484,In_2044);
and U9057 (N_9057,In_816,In_170);
or U9058 (N_9058,In_955,In_681);
nor U9059 (N_9059,In_50,In_4248);
xnor U9060 (N_9060,In_3634,In_558);
or U9061 (N_9061,In_0,In_2279);
nor U9062 (N_9062,In_3940,In_4629);
and U9063 (N_9063,In_4259,In_20);
xnor U9064 (N_9064,In_825,In_2569);
or U9065 (N_9065,In_3033,In_3334);
and U9066 (N_9066,In_654,In_2812);
xor U9067 (N_9067,In_2574,In_1804);
xor U9068 (N_9068,In_1607,In_4425);
or U9069 (N_9069,In_1638,In_4138);
nand U9070 (N_9070,In_3706,In_1037);
nor U9071 (N_9071,In_211,In_394);
and U9072 (N_9072,In_4066,In_3548);
or U9073 (N_9073,In_3223,In_3559);
nand U9074 (N_9074,In_2440,In_1717);
xnor U9075 (N_9075,In_4584,In_340);
nand U9076 (N_9076,In_2695,In_310);
xnor U9077 (N_9077,In_3559,In_3926);
xnor U9078 (N_9078,In_4991,In_4659);
or U9079 (N_9079,In_17,In_2201);
nand U9080 (N_9080,In_1786,In_3135);
xor U9081 (N_9081,In_797,In_1216);
nand U9082 (N_9082,In_924,In_2929);
and U9083 (N_9083,In_1161,In_1647);
nor U9084 (N_9084,In_4616,In_1004);
or U9085 (N_9085,In_3894,In_4676);
and U9086 (N_9086,In_1859,In_562);
and U9087 (N_9087,In_2757,In_3511);
or U9088 (N_9088,In_1198,In_1178);
xnor U9089 (N_9089,In_3835,In_4528);
nor U9090 (N_9090,In_339,In_585);
or U9091 (N_9091,In_277,In_1194);
nand U9092 (N_9092,In_3671,In_2537);
and U9093 (N_9093,In_3651,In_1235);
xor U9094 (N_9094,In_2411,In_1023);
or U9095 (N_9095,In_274,In_4498);
or U9096 (N_9096,In_4612,In_866);
or U9097 (N_9097,In_3922,In_48);
or U9098 (N_9098,In_549,In_3454);
and U9099 (N_9099,In_3759,In_4880);
xor U9100 (N_9100,In_438,In_592);
nor U9101 (N_9101,In_4284,In_4256);
nor U9102 (N_9102,In_43,In_2145);
or U9103 (N_9103,In_3008,In_3207);
xor U9104 (N_9104,In_4412,In_1583);
nand U9105 (N_9105,In_4053,In_771);
nand U9106 (N_9106,In_2490,In_2298);
xnor U9107 (N_9107,In_627,In_3186);
and U9108 (N_9108,In_2455,In_2301);
and U9109 (N_9109,In_3569,In_1917);
nand U9110 (N_9110,In_3786,In_3219);
xnor U9111 (N_9111,In_2842,In_2693);
nor U9112 (N_9112,In_278,In_970);
and U9113 (N_9113,In_1024,In_3796);
and U9114 (N_9114,In_160,In_3951);
or U9115 (N_9115,In_2771,In_713);
nand U9116 (N_9116,In_736,In_4735);
and U9117 (N_9117,In_3658,In_1015);
or U9118 (N_9118,In_924,In_639);
nor U9119 (N_9119,In_2643,In_4339);
xnor U9120 (N_9120,In_1512,In_3871);
xnor U9121 (N_9121,In_1837,In_2787);
or U9122 (N_9122,In_2969,In_3200);
nand U9123 (N_9123,In_3469,In_1077);
or U9124 (N_9124,In_3476,In_2752);
or U9125 (N_9125,In_474,In_4466);
xor U9126 (N_9126,In_2937,In_3660);
and U9127 (N_9127,In_256,In_2213);
nor U9128 (N_9128,In_1520,In_4532);
nand U9129 (N_9129,In_3843,In_1697);
nor U9130 (N_9130,In_2790,In_2814);
and U9131 (N_9131,In_1969,In_2069);
nor U9132 (N_9132,In_3534,In_3578);
and U9133 (N_9133,In_1580,In_3256);
nor U9134 (N_9134,In_1883,In_3497);
xnor U9135 (N_9135,In_4741,In_3658);
nor U9136 (N_9136,In_3380,In_627);
or U9137 (N_9137,In_4203,In_2497);
nor U9138 (N_9138,In_376,In_383);
xnor U9139 (N_9139,In_4988,In_1011);
and U9140 (N_9140,In_1383,In_403);
and U9141 (N_9141,In_4403,In_3125);
or U9142 (N_9142,In_3075,In_4470);
xnor U9143 (N_9143,In_1937,In_2215);
nor U9144 (N_9144,In_3837,In_529);
nand U9145 (N_9145,In_1647,In_2476);
nor U9146 (N_9146,In_885,In_4917);
and U9147 (N_9147,In_3836,In_3380);
nor U9148 (N_9148,In_4049,In_2096);
nand U9149 (N_9149,In_4831,In_2677);
and U9150 (N_9150,In_607,In_3119);
or U9151 (N_9151,In_1076,In_169);
nand U9152 (N_9152,In_70,In_1132);
and U9153 (N_9153,In_2319,In_1608);
and U9154 (N_9154,In_557,In_1127);
and U9155 (N_9155,In_4220,In_4520);
and U9156 (N_9156,In_4691,In_4734);
xnor U9157 (N_9157,In_4822,In_1727);
xor U9158 (N_9158,In_3340,In_2415);
nor U9159 (N_9159,In_1848,In_2995);
xor U9160 (N_9160,In_2984,In_4041);
xnor U9161 (N_9161,In_3614,In_313);
and U9162 (N_9162,In_2391,In_1850);
nor U9163 (N_9163,In_3250,In_1916);
or U9164 (N_9164,In_2813,In_2701);
nor U9165 (N_9165,In_3732,In_1668);
nor U9166 (N_9166,In_729,In_894);
xnor U9167 (N_9167,In_3563,In_759);
or U9168 (N_9168,In_1984,In_4444);
and U9169 (N_9169,In_1948,In_2342);
and U9170 (N_9170,In_2984,In_391);
nand U9171 (N_9171,In_1398,In_4227);
or U9172 (N_9172,In_2461,In_2377);
nor U9173 (N_9173,In_499,In_3652);
xnor U9174 (N_9174,In_1536,In_3683);
and U9175 (N_9175,In_2683,In_4438);
xor U9176 (N_9176,In_1277,In_3148);
and U9177 (N_9177,In_2893,In_554);
xnor U9178 (N_9178,In_708,In_1433);
nand U9179 (N_9179,In_2618,In_3889);
xor U9180 (N_9180,In_3474,In_2142);
xnor U9181 (N_9181,In_4903,In_3587);
nand U9182 (N_9182,In_2472,In_851);
and U9183 (N_9183,In_1013,In_956);
and U9184 (N_9184,In_254,In_3098);
and U9185 (N_9185,In_631,In_2470);
or U9186 (N_9186,In_891,In_4552);
or U9187 (N_9187,In_1293,In_529);
nand U9188 (N_9188,In_1824,In_4717);
nand U9189 (N_9189,In_723,In_4492);
nand U9190 (N_9190,In_489,In_723);
nor U9191 (N_9191,In_2985,In_813);
or U9192 (N_9192,In_2832,In_2617);
nor U9193 (N_9193,In_4070,In_3498);
or U9194 (N_9194,In_748,In_4955);
nand U9195 (N_9195,In_52,In_3641);
nor U9196 (N_9196,In_4463,In_1510);
nor U9197 (N_9197,In_3583,In_4918);
or U9198 (N_9198,In_3471,In_4282);
nand U9199 (N_9199,In_4220,In_1803);
nand U9200 (N_9200,In_817,In_3763);
nor U9201 (N_9201,In_3682,In_2888);
nor U9202 (N_9202,In_2250,In_3463);
nor U9203 (N_9203,In_2314,In_3308);
xor U9204 (N_9204,In_2322,In_850);
nor U9205 (N_9205,In_257,In_4520);
or U9206 (N_9206,In_4886,In_1542);
nand U9207 (N_9207,In_3141,In_4547);
and U9208 (N_9208,In_2624,In_366);
xor U9209 (N_9209,In_3647,In_1499);
xor U9210 (N_9210,In_1971,In_2718);
xor U9211 (N_9211,In_4469,In_3724);
nor U9212 (N_9212,In_890,In_201);
xnor U9213 (N_9213,In_2838,In_1467);
and U9214 (N_9214,In_3963,In_2376);
nor U9215 (N_9215,In_2302,In_4813);
nand U9216 (N_9216,In_4948,In_3825);
and U9217 (N_9217,In_3952,In_2166);
xor U9218 (N_9218,In_3510,In_2717);
xor U9219 (N_9219,In_2341,In_4639);
or U9220 (N_9220,In_3829,In_3972);
or U9221 (N_9221,In_4620,In_2722);
nor U9222 (N_9222,In_2605,In_323);
and U9223 (N_9223,In_3380,In_1828);
nand U9224 (N_9224,In_19,In_3375);
and U9225 (N_9225,In_3245,In_1535);
and U9226 (N_9226,In_918,In_3479);
nor U9227 (N_9227,In_1914,In_1396);
nor U9228 (N_9228,In_2830,In_1028);
nand U9229 (N_9229,In_3166,In_3048);
nand U9230 (N_9230,In_523,In_2707);
nor U9231 (N_9231,In_329,In_1048);
or U9232 (N_9232,In_3658,In_638);
nand U9233 (N_9233,In_533,In_922);
nand U9234 (N_9234,In_1293,In_1569);
or U9235 (N_9235,In_1328,In_1143);
or U9236 (N_9236,In_2670,In_2250);
xor U9237 (N_9237,In_4076,In_877);
xor U9238 (N_9238,In_884,In_1313);
xor U9239 (N_9239,In_3105,In_4489);
nor U9240 (N_9240,In_4757,In_4948);
nand U9241 (N_9241,In_4448,In_1244);
and U9242 (N_9242,In_3110,In_1046);
nand U9243 (N_9243,In_1262,In_3225);
and U9244 (N_9244,In_2696,In_248);
nor U9245 (N_9245,In_1650,In_543);
or U9246 (N_9246,In_53,In_3781);
or U9247 (N_9247,In_4402,In_4674);
or U9248 (N_9248,In_2779,In_622);
and U9249 (N_9249,In_1964,In_4244);
xnor U9250 (N_9250,In_673,In_460);
nor U9251 (N_9251,In_1580,In_3248);
xnor U9252 (N_9252,In_2678,In_4715);
and U9253 (N_9253,In_4161,In_484);
nor U9254 (N_9254,In_2542,In_1451);
or U9255 (N_9255,In_3174,In_4694);
or U9256 (N_9256,In_3190,In_1096);
nand U9257 (N_9257,In_1856,In_2137);
xnor U9258 (N_9258,In_3222,In_3975);
or U9259 (N_9259,In_368,In_470);
and U9260 (N_9260,In_3540,In_1195);
nand U9261 (N_9261,In_4996,In_3208);
and U9262 (N_9262,In_4000,In_2428);
and U9263 (N_9263,In_264,In_4338);
nor U9264 (N_9264,In_2013,In_2263);
nor U9265 (N_9265,In_2417,In_1254);
nand U9266 (N_9266,In_4385,In_4119);
nor U9267 (N_9267,In_525,In_2531);
nor U9268 (N_9268,In_4011,In_2040);
xor U9269 (N_9269,In_2057,In_769);
nor U9270 (N_9270,In_746,In_1907);
nand U9271 (N_9271,In_3787,In_195);
xor U9272 (N_9272,In_604,In_26);
nor U9273 (N_9273,In_1632,In_3992);
nor U9274 (N_9274,In_1334,In_9);
nand U9275 (N_9275,In_1511,In_1392);
nor U9276 (N_9276,In_3373,In_2303);
xnor U9277 (N_9277,In_2503,In_4232);
nand U9278 (N_9278,In_2463,In_4938);
xnor U9279 (N_9279,In_1426,In_335);
nand U9280 (N_9280,In_3364,In_185);
xnor U9281 (N_9281,In_1064,In_4397);
and U9282 (N_9282,In_258,In_1335);
nand U9283 (N_9283,In_1186,In_357);
nor U9284 (N_9284,In_2675,In_4283);
nor U9285 (N_9285,In_1955,In_513);
and U9286 (N_9286,In_1382,In_4550);
nand U9287 (N_9287,In_4995,In_4361);
nor U9288 (N_9288,In_3696,In_2703);
nand U9289 (N_9289,In_4275,In_6);
xnor U9290 (N_9290,In_1839,In_3525);
nor U9291 (N_9291,In_4455,In_287);
nor U9292 (N_9292,In_4998,In_4598);
and U9293 (N_9293,In_604,In_3469);
or U9294 (N_9294,In_3745,In_1561);
xor U9295 (N_9295,In_4091,In_516);
xnor U9296 (N_9296,In_4836,In_3606);
nor U9297 (N_9297,In_2481,In_3596);
xor U9298 (N_9298,In_951,In_4265);
nor U9299 (N_9299,In_1950,In_911);
nor U9300 (N_9300,In_4963,In_360);
and U9301 (N_9301,In_3805,In_2464);
nor U9302 (N_9302,In_4134,In_3893);
or U9303 (N_9303,In_2323,In_2438);
or U9304 (N_9304,In_152,In_4854);
nor U9305 (N_9305,In_3944,In_3097);
or U9306 (N_9306,In_987,In_3767);
xnor U9307 (N_9307,In_2588,In_2085);
xor U9308 (N_9308,In_4864,In_2745);
nand U9309 (N_9309,In_4343,In_3529);
and U9310 (N_9310,In_4444,In_3982);
or U9311 (N_9311,In_899,In_217);
or U9312 (N_9312,In_579,In_2049);
nand U9313 (N_9313,In_2995,In_1472);
or U9314 (N_9314,In_892,In_4681);
and U9315 (N_9315,In_1181,In_2190);
nor U9316 (N_9316,In_2330,In_1436);
xor U9317 (N_9317,In_2066,In_4038);
or U9318 (N_9318,In_1521,In_3516);
or U9319 (N_9319,In_3947,In_656);
xnor U9320 (N_9320,In_704,In_2374);
xnor U9321 (N_9321,In_1555,In_4182);
xor U9322 (N_9322,In_602,In_597);
nor U9323 (N_9323,In_165,In_3432);
nor U9324 (N_9324,In_4889,In_4000);
or U9325 (N_9325,In_412,In_212);
xnor U9326 (N_9326,In_4873,In_1589);
nor U9327 (N_9327,In_2866,In_4571);
nor U9328 (N_9328,In_4896,In_3562);
xnor U9329 (N_9329,In_4848,In_1847);
nand U9330 (N_9330,In_2551,In_286);
or U9331 (N_9331,In_2344,In_1504);
nor U9332 (N_9332,In_2037,In_456);
or U9333 (N_9333,In_4453,In_3094);
and U9334 (N_9334,In_4164,In_3835);
nand U9335 (N_9335,In_992,In_1645);
nand U9336 (N_9336,In_3252,In_3465);
xnor U9337 (N_9337,In_3936,In_455);
and U9338 (N_9338,In_994,In_803);
nand U9339 (N_9339,In_515,In_2239);
or U9340 (N_9340,In_3856,In_3498);
or U9341 (N_9341,In_1182,In_2830);
nand U9342 (N_9342,In_818,In_4251);
xor U9343 (N_9343,In_1083,In_1737);
nand U9344 (N_9344,In_2774,In_1496);
xnor U9345 (N_9345,In_2640,In_2588);
nand U9346 (N_9346,In_3968,In_1454);
and U9347 (N_9347,In_4810,In_4070);
nor U9348 (N_9348,In_529,In_3109);
and U9349 (N_9349,In_4167,In_1320);
and U9350 (N_9350,In_3139,In_2145);
xnor U9351 (N_9351,In_1921,In_1652);
nand U9352 (N_9352,In_2591,In_3475);
and U9353 (N_9353,In_825,In_460);
or U9354 (N_9354,In_4920,In_2327);
and U9355 (N_9355,In_3521,In_2349);
and U9356 (N_9356,In_3947,In_1878);
and U9357 (N_9357,In_3079,In_3214);
nand U9358 (N_9358,In_1222,In_3573);
and U9359 (N_9359,In_4850,In_478);
and U9360 (N_9360,In_4072,In_913);
or U9361 (N_9361,In_1792,In_83);
xnor U9362 (N_9362,In_3249,In_2574);
xor U9363 (N_9363,In_1809,In_4172);
nand U9364 (N_9364,In_3554,In_2305);
nand U9365 (N_9365,In_4095,In_4781);
xnor U9366 (N_9366,In_2695,In_2640);
or U9367 (N_9367,In_1467,In_2268);
nand U9368 (N_9368,In_1012,In_4673);
nand U9369 (N_9369,In_2488,In_3594);
and U9370 (N_9370,In_3362,In_570);
or U9371 (N_9371,In_3672,In_4911);
and U9372 (N_9372,In_1994,In_3933);
and U9373 (N_9373,In_1206,In_4776);
nor U9374 (N_9374,In_2031,In_1275);
nand U9375 (N_9375,In_3759,In_1412);
or U9376 (N_9376,In_785,In_1606);
nand U9377 (N_9377,In_1991,In_1732);
nand U9378 (N_9378,In_1481,In_4096);
xor U9379 (N_9379,In_4818,In_1214);
xnor U9380 (N_9380,In_705,In_2853);
or U9381 (N_9381,In_346,In_1645);
or U9382 (N_9382,In_3459,In_3587);
nor U9383 (N_9383,In_423,In_377);
xnor U9384 (N_9384,In_535,In_4922);
and U9385 (N_9385,In_1719,In_3108);
or U9386 (N_9386,In_4440,In_1692);
or U9387 (N_9387,In_4459,In_1426);
nand U9388 (N_9388,In_3463,In_1108);
nor U9389 (N_9389,In_376,In_3022);
xnor U9390 (N_9390,In_2652,In_3924);
and U9391 (N_9391,In_2403,In_1861);
or U9392 (N_9392,In_833,In_2792);
nand U9393 (N_9393,In_3825,In_18);
and U9394 (N_9394,In_4450,In_4560);
xnor U9395 (N_9395,In_2154,In_3530);
nor U9396 (N_9396,In_1141,In_441);
nor U9397 (N_9397,In_3118,In_2152);
or U9398 (N_9398,In_4099,In_1739);
xnor U9399 (N_9399,In_4936,In_2793);
and U9400 (N_9400,In_4114,In_535);
xnor U9401 (N_9401,In_1240,In_838);
nand U9402 (N_9402,In_2874,In_2468);
xnor U9403 (N_9403,In_2470,In_1864);
nand U9404 (N_9404,In_2797,In_976);
xnor U9405 (N_9405,In_338,In_2480);
and U9406 (N_9406,In_1935,In_4330);
xor U9407 (N_9407,In_479,In_822);
xor U9408 (N_9408,In_4748,In_4513);
nand U9409 (N_9409,In_1599,In_1494);
and U9410 (N_9410,In_4797,In_4191);
and U9411 (N_9411,In_1173,In_3692);
xnor U9412 (N_9412,In_603,In_3974);
or U9413 (N_9413,In_4846,In_3913);
xnor U9414 (N_9414,In_3860,In_3113);
xnor U9415 (N_9415,In_770,In_1949);
and U9416 (N_9416,In_1305,In_2432);
or U9417 (N_9417,In_4619,In_4679);
nand U9418 (N_9418,In_3650,In_4472);
nor U9419 (N_9419,In_3236,In_1240);
nor U9420 (N_9420,In_766,In_3408);
xor U9421 (N_9421,In_573,In_625);
nand U9422 (N_9422,In_2559,In_1511);
and U9423 (N_9423,In_1598,In_334);
or U9424 (N_9424,In_1791,In_4810);
xnor U9425 (N_9425,In_1198,In_4851);
and U9426 (N_9426,In_558,In_1169);
xnor U9427 (N_9427,In_53,In_623);
nor U9428 (N_9428,In_3790,In_4636);
and U9429 (N_9429,In_4314,In_2665);
nor U9430 (N_9430,In_1388,In_690);
and U9431 (N_9431,In_91,In_2141);
xnor U9432 (N_9432,In_3554,In_4478);
and U9433 (N_9433,In_3903,In_1840);
and U9434 (N_9434,In_2931,In_2665);
or U9435 (N_9435,In_1560,In_2599);
or U9436 (N_9436,In_4306,In_4514);
and U9437 (N_9437,In_3824,In_3732);
and U9438 (N_9438,In_3958,In_1749);
and U9439 (N_9439,In_3461,In_724);
or U9440 (N_9440,In_2173,In_681);
or U9441 (N_9441,In_760,In_3159);
nor U9442 (N_9442,In_2443,In_2566);
and U9443 (N_9443,In_1278,In_3962);
and U9444 (N_9444,In_4375,In_2116);
or U9445 (N_9445,In_4768,In_662);
nor U9446 (N_9446,In_1585,In_2722);
nand U9447 (N_9447,In_511,In_3693);
nand U9448 (N_9448,In_422,In_71);
xnor U9449 (N_9449,In_134,In_2900);
and U9450 (N_9450,In_2818,In_142);
or U9451 (N_9451,In_4970,In_398);
nor U9452 (N_9452,In_1989,In_3378);
and U9453 (N_9453,In_3304,In_3207);
nor U9454 (N_9454,In_265,In_1255);
xnor U9455 (N_9455,In_3696,In_574);
or U9456 (N_9456,In_3046,In_4602);
and U9457 (N_9457,In_1918,In_393);
or U9458 (N_9458,In_1461,In_747);
and U9459 (N_9459,In_2165,In_4212);
xor U9460 (N_9460,In_3645,In_4363);
or U9461 (N_9461,In_1275,In_600);
and U9462 (N_9462,In_1442,In_2533);
nand U9463 (N_9463,In_3094,In_4053);
nand U9464 (N_9464,In_1388,In_1775);
nand U9465 (N_9465,In_4216,In_3322);
nor U9466 (N_9466,In_1286,In_188);
xor U9467 (N_9467,In_1399,In_912);
nand U9468 (N_9468,In_2752,In_4275);
or U9469 (N_9469,In_2926,In_48);
nor U9470 (N_9470,In_1729,In_3471);
and U9471 (N_9471,In_1345,In_3860);
or U9472 (N_9472,In_2221,In_274);
xor U9473 (N_9473,In_1178,In_1732);
or U9474 (N_9474,In_1678,In_926);
and U9475 (N_9475,In_4531,In_804);
nand U9476 (N_9476,In_4405,In_2009);
and U9477 (N_9477,In_2213,In_3946);
nand U9478 (N_9478,In_3294,In_4841);
xor U9479 (N_9479,In_1821,In_1060);
or U9480 (N_9480,In_1335,In_309);
nand U9481 (N_9481,In_3502,In_4920);
and U9482 (N_9482,In_2378,In_2486);
nor U9483 (N_9483,In_3149,In_2961);
or U9484 (N_9484,In_4784,In_2793);
nand U9485 (N_9485,In_4415,In_2075);
nor U9486 (N_9486,In_1740,In_2178);
or U9487 (N_9487,In_2983,In_416);
or U9488 (N_9488,In_409,In_2972);
or U9489 (N_9489,In_753,In_4866);
and U9490 (N_9490,In_1455,In_3524);
nand U9491 (N_9491,In_2549,In_4091);
nand U9492 (N_9492,In_4606,In_3189);
xnor U9493 (N_9493,In_3170,In_2758);
xor U9494 (N_9494,In_3896,In_1089);
nand U9495 (N_9495,In_4912,In_1199);
xor U9496 (N_9496,In_2348,In_1487);
or U9497 (N_9497,In_1520,In_403);
or U9498 (N_9498,In_1372,In_2968);
and U9499 (N_9499,In_3916,In_77);
and U9500 (N_9500,In_1170,In_1985);
xnor U9501 (N_9501,In_4342,In_3846);
nor U9502 (N_9502,In_4788,In_3443);
or U9503 (N_9503,In_4272,In_4877);
nor U9504 (N_9504,In_3895,In_1165);
nor U9505 (N_9505,In_3648,In_1139);
and U9506 (N_9506,In_2524,In_1915);
nand U9507 (N_9507,In_3604,In_4772);
and U9508 (N_9508,In_2900,In_2170);
nand U9509 (N_9509,In_4558,In_1754);
or U9510 (N_9510,In_4859,In_683);
nor U9511 (N_9511,In_2077,In_1554);
nand U9512 (N_9512,In_2815,In_3205);
nand U9513 (N_9513,In_3859,In_4351);
nor U9514 (N_9514,In_3569,In_4854);
nor U9515 (N_9515,In_619,In_486);
and U9516 (N_9516,In_1684,In_4795);
xor U9517 (N_9517,In_1366,In_4767);
nand U9518 (N_9518,In_1297,In_1333);
and U9519 (N_9519,In_1083,In_1027);
xor U9520 (N_9520,In_1488,In_2191);
or U9521 (N_9521,In_1948,In_1265);
nor U9522 (N_9522,In_3013,In_3360);
and U9523 (N_9523,In_1122,In_2245);
or U9524 (N_9524,In_2914,In_219);
nor U9525 (N_9525,In_3653,In_4971);
and U9526 (N_9526,In_4764,In_691);
or U9527 (N_9527,In_3167,In_326);
nand U9528 (N_9528,In_4723,In_474);
or U9529 (N_9529,In_1550,In_444);
or U9530 (N_9530,In_402,In_600);
nand U9531 (N_9531,In_3991,In_3270);
xor U9532 (N_9532,In_3943,In_4144);
or U9533 (N_9533,In_1779,In_1588);
or U9534 (N_9534,In_2423,In_1746);
and U9535 (N_9535,In_3479,In_4844);
nand U9536 (N_9536,In_2603,In_4582);
or U9537 (N_9537,In_4253,In_4602);
xnor U9538 (N_9538,In_2956,In_2586);
nor U9539 (N_9539,In_4425,In_3382);
nor U9540 (N_9540,In_1289,In_596);
xnor U9541 (N_9541,In_4641,In_1960);
and U9542 (N_9542,In_4721,In_990);
or U9543 (N_9543,In_1930,In_2152);
xor U9544 (N_9544,In_2975,In_2100);
xnor U9545 (N_9545,In_749,In_4963);
or U9546 (N_9546,In_3613,In_2490);
nor U9547 (N_9547,In_905,In_45);
and U9548 (N_9548,In_1075,In_1499);
or U9549 (N_9549,In_323,In_2776);
nor U9550 (N_9550,In_4489,In_1823);
and U9551 (N_9551,In_710,In_2319);
nand U9552 (N_9552,In_4190,In_1709);
nand U9553 (N_9553,In_2765,In_1485);
xor U9554 (N_9554,In_241,In_3726);
or U9555 (N_9555,In_1785,In_115);
or U9556 (N_9556,In_1375,In_4809);
nor U9557 (N_9557,In_4443,In_2785);
nor U9558 (N_9558,In_2490,In_4089);
and U9559 (N_9559,In_3611,In_4434);
and U9560 (N_9560,In_3136,In_4391);
xnor U9561 (N_9561,In_4582,In_1868);
xnor U9562 (N_9562,In_172,In_4003);
nand U9563 (N_9563,In_465,In_4193);
nand U9564 (N_9564,In_3114,In_4267);
xor U9565 (N_9565,In_2977,In_313);
nand U9566 (N_9566,In_2349,In_2949);
nand U9567 (N_9567,In_2554,In_3150);
nor U9568 (N_9568,In_3126,In_2287);
or U9569 (N_9569,In_2760,In_2784);
or U9570 (N_9570,In_2201,In_1116);
and U9571 (N_9571,In_4785,In_4506);
or U9572 (N_9572,In_2396,In_2634);
nor U9573 (N_9573,In_2709,In_3217);
nor U9574 (N_9574,In_2295,In_4039);
nor U9575 (N_9575,In_2941,In_3541);
xnor U9576 (N_9576,In_3358,In_3937);
and U9577 (N_9577,In_4186,In_4687);
or U9578 (N_9578,In_196,In_1295);
nor U9579 (N_9579,In_896,In_824);
nand U9580 (N_9580,In_1906,In_891);
nor U9581 (N_9581,In_4777,In_4118);
xnor U9582 (N_9582,In_824,In_1049);
and U9583 (N_9583,In_3546,In_3069);
nand U9584 (N_9584,In_3759,In_4934);
and U9585 (N_9585,In_1075,In_1357);
xor U9586 (N_9586,In_3423,In_2062);
and U9587 (N_9587,In_1598,In_1478);
nor U9588 (N_9588,In_4353,In_229);
or U9589 (N_9589,In_1346,In_1706);
and U9590 (N_9590,In_4731,In_3925);
or U9591 (N_9591,In_673,In_127);
nand U9592 (N_9592,In_1514,In_2052);
and U9593 (N_9593,In_2407,In_3363);
and U9594 (N_9594,In_1161,In_4380);
xor U9595 (N_9595,In_3286,In_4534);
nand U9596 (N_9596,In_1967,In_3721);
nand U9597 (N_9597,In_3826,In_1276);
nor U9598 (N_9598,In_3679,In_4492);
xnor U9599 (N_9599,In_4471,In_3926);
xor U9600 (N_9600,In_3258,In_828);
nand U9601 (N_9601,In_3204,In_1180);
and U9602 (N_9602,In_3418,In_3612);
nand U9603 (N_9603,In_4016,In_1389);
and U9604 (N_9604,In_420,In_3437);
or U9605 (N_9605,In_1178,In_724);
or U9606 (N_9606,In_300,In_186);
xor U9607 (N_9607,In_1685,In_3758);
nor U9608 (N_9608,In_4103,In_1057);
or U9609 (N_9609,In_1547,In_4474);
nand U9610 (N_9610,In_3880,In_2524);
nand U9611 (N_9611,In_3234,In_4986);
nor U9612 (N_9612,In_1209,In_188);
xor U9613 (N_9613,In_4967,In_3099);
nor U9614 (N_9614,In_4308,In_3583);
xor U9615 (N_9615,In_2004,In_1641);
and U9616 (N_9616,In_67,In_4047);
or U9617 (N_9617,In_829,In_1468);
nand U9618 (N_9618,In_3829,In_933);
or U9619 (N_9619,In_96,In_73);
and U9620 (N_9620,In_2341,In_3039);
or U9621 (N_9621,In_199,In_2080);
xnor U9622 (N_9622,In_4713,In_639);
nor U9623 (N_9623,In_3871,In_276);
nand U9624 (N_9624,In_4468,In_2003);
and U9625 (N_9625,In_2160,In_353);
and U9626 (N_9626,In_2174,In_1723);
and U9627 (N_9627,In_4088,In_4219);
nand U9628 (N_9628,In_3617,In_1203);
and U9629 (N_9629,In_3411,In_4667);
nor U9630 (N_9630,In_4435,In_1285);
xnor U9631 (N_9631,In_2566,In_2556);
and U9632 (N_9632,In_3786,In_2715);
xor U9633 (N_9633,In_3173,In_3195);
and U9634 (N_9634,In_2573,In_3940);
nand U9635 (N_9635,In_310,In_1982);
xnor U9636 (N_9636,In_845,In_1025);
xor U9637 (N_9637,In_4664,In_251);
xnor U9638 (N_9638,In_391,In_1349);
or U9639 (N_9639,In_253,In_255);
or U9640 (N_9640,In_4941,In_3053);
nor U9641 (N_9641,In_1964,In_4255);
and U9642 (N_9642,In_4824,In_570);
nand U9643 (N_9643,In_454,In_3245);
nor U9644 (N_9644,In_2653,In_1907);
nand U9645 (N_9645,In_1281,In_942);
xor U9646 (N_9646,In_497,In_3947);
and U9647 (N_9647,In_2589,In_2627);
nand U9648 (N_9648,In_2467,In_1597);
nand U9649 (N_9649,In_2296,In_4048);
or U9650 (N_9650,In_2009,In_4226);
xor U9651 (N_9651,In_101,In_3327);
xnor U9652 (N_9652,In_834,In_1122);
nand U9653 (N_9653,In_4522,In_356);
xor U9654 (N_9654,In_722,In_3824);
nand U9655 (N_9655,In_1169,In_2095);
nand U9656 (N_9656,In_520,In_4169);
and U9657 (N_9657,In_3676,In_2667);
and U9658 (N_9658,In_734,In_909);
nand U9659 (N_9659,In_936,In_2152);
and U9660 (N_9660,In_1076,In_297);
nor U9661 (N_9661,In_47,In_1244);
nand U9662 (N_9662,In_3801,In_1197);
and U9663 (N_9663,In_1056,In_3577);
or U9664 (N_9664,In_2809,In_2837);
xnor U9665 (N_9665,In_632,In_1612);
xnor U9666 (N_9666,In_1612,In_1567);
or U9667 (N_9667,In_13,In_1762);
xnor U9668 (N_9668,In_2338,In_2922);
or U9669 (N_9669,In_2552,In_3815);
or U9670 (N_9670,In_4032,In_3510);
or U9671 (N_9671,In_184,In_2005);
or U9672 (N_9672,In_4442,In_1750);
nor U9673 (N_9673,In_3785,In_1244);
and U9674 (N_9674,In_2267,In_2237);
nor U9675 (N_9675,In_4377,In_1108);
nand U9676 (N_9676,In_1930,In_1885);
and U9677 (N_9677,In_370,In_1190);
xnor U9678 (N_9678,In_754,In_4148);
and U9679 (N_9679,In_881,In_3863);
nand U9680 (N_9680,In_1228,In_4304);
xnor U9681 (N_9681,In_2180,In_1959);
nor U9682 (N_9682,In_4190,In_3504);
and U9683 (N_9683,In_2497,In_3712);
and U9684 (N_9684,In_4861,In_3795);
xor U9685 (N_9685,In_2726,In_3700);
or U9686 (N_9686,In_4931,In_4923);
xor U9687 (N_9687,In_1819,In_1160);
nand U9688 (N_9688,In_4942,In_1535);
or U9689 (N_9689,In_4212,In_152);
nand U9690 (N_9690,In_31,In_2048);
xor U9691 (N_9691,In_556,In_3061);
nand U9692 (N_9692,In_1812,In_4595);
and U9693 (N_9693,In_572,In_1949);
nor U9694 (N_9694,In_4061,In_3778);
or U9695 (N_9695,In_1909,In_2246);
and U9696 (N_9696,In_3865,In_1661);
xnor U9697 (N_9697,In_1952,In_4672);
and U9698 (N_9698,In_2418,In_3495);
nor U9699 (N_9699,In_1878,In_4032);
nand U9700 (N_9700,In_1500,In_123);
nand U9701 (N_9701,In_3022,In_634);
xnor U9702 (N_9702,In_2063,In_3203);
nand U9703 (N_9703,In_3970,In_521);
xnor U9704 (N_9704,In_3077,In_4195);
xor U9705 (N_9705,In_3887,In_223);
xor U9706 (N_9706,In_2648,In_1195);
xor U9707 (N_9707,In_4598,In_3427);
nand U9708 (N_9708,In_1542,In_382);
xnor U9709 (N_9709,In_2372,In_1231);
xor U9710 (N_9710,In_3529,In_4498);
nor U9711 (N_9711,In_4644,In_622);
nand U9712 (N_9712,In_4557,In_3487);
nand U9713 (N_9713,In_4596,In_4813);
and U9714 (N_9714,In_2898,In_1680);
nand U9715 (N_9715,In_3810,In_2686);
xnor U9716 (N_9716,In_1440,In_4176);
nor U9717 (N_9717,In_1876,In_1715);
nand U9718 (N_9718,In_4407,In_285);
nor U9719 (N_9719,In_2142,In_1182);
or U9720 (N_9720,In_246,In_3440);
nor U9721 (N_9721,In_4779,In_4209);
nand U9722 (N_9722,In_2601,In_4164);
xor U9723 (N_9723,In_587,In_2351);
or U9724 (N_9724,In_2109,In_1311);
nand U9725 (N_9725,In_6,In_4373);
and U9726 (N_9726,In_1090,In_3594);
or U9727 (N_9727,In_3339,In_3434);
xor U9728 (N_9728,In_4192,In_1313);
and U9729 (N_9729,In_4637,In_1113);
nand U9730 (N_9730,In_4683,In_4334);
or U9731 (N_9731,In_2842,In_1105);
nand U9732 (N_9732,In_434,In_4304);
nand U9733 (N_9733,In_981,In_319);
nand U9734 (N_9734,In_4018,In_2387);
xnor U9735 (N_9735,In_181,In_112);
and U9736 (N_9736,In_378,In_3840);
nand U9737 (N_9737,In_2758,In_4303);
xor U9738 (N_9738,In_1654,In_1);
or U9739 (N_9739,In_1223,In_4429);
nand U9740 (N_9740,In_2451,In_3850);
nor U9741 (N_9741,In_2097,In_3852);
nor U9742 (N_9742,In_4577,In_3210);
nor U9743 (N_9743,In_4890,In_3488);
xor U9744 (N_9744,In_3038,In_4468);
xnor U9745 (N_9745,In_663,In_1400);
xor U9746 (N_9746,In_3079,In_3898);
or U9747 (N_9747,In_2207,In_3085);
and U9748 (N_9748,In_4848,In_2941);
nand U9749 (N_9749,In_3106,In_1667);
xnor U9750 (N_9750,In_113,In_4669);
or U9751 (N_9751,In_3751,In_4841);
nor U9752 (N_9752,In_3792,In_574);
xor U9753 (N_9753,In_4890,In_3262);
and U9754 (N_9754,In_2312,In_2122);
and U9755 (N_9755,In_2301,In_2483);
nand U9756 (N_9756,In_1591,In_117);
or U9757 (N_9757,In_3266,In_339);
nand U9758 (N_9758,In_4038,In_4520);
xor U9759 (N_9759,In_3282,In_2947);
and U9760 (N_9760,In_3224,In_4229);
nand U9761 (N_9761,In_2007,In_2354);
xnor U9762 (N_9762,In_3324,In_160);
nor U9763 (N_9763,In_2183,In_3635);
nand U9764 (N_9764,In_2654,In_1019);
nor U9765 (N_9765,In_3710,In_3850);
and U9766 (N_9766,In_2111,In_4186);
nor U9767 (N_9767,In_4697,In_4861);
nor U9768 (N_9768,In_1126,In_3719);
and U9769 (N_9769,In_2139,In_2191);
nor U9770 (N_9770,In_1107,In_1788);
nor U9771 (N_9771,In_1808,In_2176);
nor U9772 (N_9772,In_1913,In_3106);
and U9773 (N_9773,In_2167,In_116);
and U9774 (N_9774,In_1316,In_3425);
or U9775 (N_9775,In_4185,In_792);
nor U9776 (N_9776,In_661,In_3146);
and U9777 (N_9777,In_4105,In_3787);
and U9778 (N_9778,In_1604,In_3464);
or U9779 (N_9779,In_4759,In_3790);
or U9780 (N_9780,In_3977,In_1370);
or U9781 (N_9781,In_1323,In_2533);
xnor U9782 (N_9782,In_3719,In_3188);
and U9783 (N_9783,In_1048,In_380);
nand U9784 (N_9784,In_484,In_2161);
xnor U9785 (N_9785,In_1823,In_2040);
or U9786 (N_9786,In_3070,In_3985);
and U9787 (N_9787,In_453,In_3196);
xor U9788 (N_9788,In_4838,In_1928);
and U9789 (N_9789,In_1283,In_3499);
or U9790 (N_9790,In_1077,In_4171);
or U9791 (N_9791,In_2688,In_3086);
nor U9792 (N_9792,In_2871,In_409);
or U9793 (N_9793,In_514,In_4051);
nor U9794 (N_9794,In_4185,In_4048);
nor U9795 (N_9795,In_2883,In_454);
xnor U9796 (N_9796,In_4763,In_1502);
nand U9797 (N_9797,In_692,In_2198);
and U9798 (N_9798,In_4512,In_3545);
or U9799 (N_9799,In_1355,In_1016);
or U9800 (N_9800,In_4550,In_2975);
nand U9801 (N_9801,In_4101,In_4926);
xor U9802 (N_9802,In_387,In_4963);
and U9803 (N_9803,In_4099,In_2390);
or U9804 (N_9804,In_370,In_3339);
and U9805 (N_9805,In_868,In_1841);
or U9806 (N_9806,In_2148,In_3541);
and U9807 (N_9807,In_1079,In_3529);
nor U9808 (N_9808,In_70,In_3187);
or U9809 (N_9809,In_1336,In_2584);
xnor U9810 (N_9810,In_419,In_210);
or U9811 (N_9811,In_568,In_1377);
nand U9812 (N_9812,In_4254,In_1637);
xnor U9813 (N_9813,In_3267,In_4999);
xnor U9814 (N_9814,In_698,In_1380);
xor U9815 (N_9815,In_3111,In_2262);
or U9816 (N_9816,In_2484,In_3388);
nand U9817 (N_9817,In_2661,In_1690);
or U9818 (N_9818,In_2155,In_355);
nand U9819 (N_9819,In_268,In_4942);
and U9820 (N_9820,In_4571,In_1090);
nand U9821 (N_9821,In_3950,In_1843);
nor U9822 (N_9822,In_342,In_4958);
xor U9823 (N_9823,In_513,In_2563);
nor U9824 (N_9824,In_1341,In_1288);
xor U9825 (N_9825,In_1973,In_1647);
xnor U9826 (N_9826,In_417,In_1645);
xor U9827 (N_9827,In_2422,In_1955);
and U9828 (N_9828,In_2883,In_3193);
xor U9829 (N_9829,In_3897,In_4033);
nor U9830 (N_9830,In_3581,In_1076);
nor U9831 (N_9831,In_3114,In_4212);
xor U9832 (N_9832,In_1812,In_798);
or U9833 (N_9833,In_4132,In_4788);
xnor U9834 (N_9834,In_2747,In_1153);
or U9835 (N_9835,In_1974,In_1348);
xnor U9836 (N_9836,In_232,In_1019);
nor U9837 (N_9837,In_34,In_4542);
or U9838 (N_9838,In_4581,In_4504);
and U9839 (N_9839,In_1666,In_590);
nor U9840 (N_9840,In_1932,In_3465);
and U9841 (N_9841,In_2634,In_4576);
and U9842 (N_9842,In_4025,In_2848);
nand U9843 (N_9843,In_1846,In_2001);
or U9844 (N_9844,In_4828,In_3218);
and U9845 (N_9845,In_1573,In_3999);
or U9846 (N_9846,In_3427,In_3522);
nand U9847 (N_9847,In_4352,In_305);
or U9848 (N_9848,In_4083,In_453);
xor U9849 (N_9849,In_3196,In_2914);
nor U9850 (N_9850,In_2682,In_2621);
and U9851 (N_9851,In_4196,In_2838);
nand U9852 (N_9852,In_2118,In_266);
or U9853 (N_9853,In_3280,In_3760);
xor U9854 (N_9854,In_3427,In_1837);
nand U9855 (N_9855,In_4378,In_1375);
or U9856 (N_9856,In_1645,In_4829);
or U9857 (N_9857,In_3708,In_1765);
and U9858 (N_9858,In_9,In_1041);
nor U9859 (N_9859,In_4081,In_312);
nand U9860 (N_9860,In_4942,In_797);
and U9861 (N_9861,In_2467,In_3094);
nand U9862 (N_9862,In_3869,In_3138);
nand U9863 (N_9863,In_1936,In_878);
nand U9864 (N_9864,In_2234,In_80);
nor U9865 (N_9865,In_1935,In_3724);
nand U9866 (N_9866,In_1464,In_638);
nand U9867 (N_9867,In_1653,In_4061);
or U9868 (N_9868,In_640,In_3199);
and U9869 (N_9869,In_731,In_4569);
xnor U9870 (N_9870,In_2005,In_1774);
xor U9871 (N_9871,In_3067,In_1797);
or U9872 (N_9872,In_1808,In_205);
or U9873 (N_9873,In_2043,In_4297);
xor U9874 (N_9874,In_2990,In_4385);
nand U9875 (N_9875,In_3673,In_1450);
and U9876 (N_9876,In_2534,In_775);
nor U9877 (N_9877,In_1867,In_2452);
or U9878 (N_9878,In_2181,In_4584);
or U9879 (N_9879,In_2601,In_1756);
nor U9880 (N_9880,In_4979,In_3960);
and U9881 (N_9881,In_1787,In_723);
or U9882 (N_9882,In_1701,In_642);
nand U9883 (N_9883,In_2947,In_1638);
nor U9884 (N_9884,In_3733,In_1168);
nor U9885 (N_9885,In_4006,In_4736);
nand U9886 (N_9886,In_4499,In_480);
nand U9887 (N_9887,In_2760,In_4476);
xnor U9888 (N_9888,In_3077,In_1226);
nor U9889 (N_9889,In_1578,In_4823);
xor U9890 (N_9890,In_2906,In_3038);
and U9891 (N_9891,In_2095,In_2280);
nor U9892 (N_9892,In_2439,In_3502);
or U9893 (N_9893,In_1538,In_258);
or U9894 (N_9894,In_3903,In_4138);
nand U9895 (N_9895,In_4482,In_3272);
xor U9896 (N_9896,In_1892,In_500);
or U9897 (N_9897,In_4154,In_4772);
nand U9898 (N_9898,In_480,In_3198);
nand U9899 (N_9899,In_1725,In_2231);
nor U9900 (N_9900,In_2854,In_4636);
or U9901 (N_9901,In_4507,In_4244);
and U9902 (N_9902,In_3614,In_3858);
or U9903 (N_9903,In_2350,In_451);
xnor U9904 (N_9904,In_1946,In_1040);
xnor U9905 (N_9905,In_4039,In_1511);
nand U9906 (N_9906,In_192,In_3161);
xnor U9907 (N_9907,In_2599,In_288);
nor U9908 (N_9908,In_1678,In_272);
xnor U9909 (N_9909,In_1611,In_2396);
nor U9910 (N_9910,In_691,In_502);
xnor U9911 (N_9911,In_35,In_4970);
xnor U9912 (N_9912,In_1802,In_1819);
or U9913 (N_9913,In_4491,In_908);
or U9914 (N_9914,In_3270,In_3887);
nor U9915 (N_9915,In_914,In_4791);
and U9916 (N_9916,In_374,In_2136);
or U9917 (N_9917,In_2796,In_3743);
or U9918 (N_9918,In_1745,In_2033);
xnor U9919 (N_9919,In_1814,In_4739);
and U9920 (N_9920,In_1498,In_2804);
nor U9921 (N_9921,In_2204,In_2313);
or U9922 (N_9922,In_4787,In_1989);
or U9923 (N_9923,In_1993,In_4948);
and U9924 (N_9924,In_4885,In_1400);
or U9925 (N_9925,In_4146,In_1092);
nor U9926 (N_9926,In_1059,In_4654);
and U9927 (N_9927,In_2809,In_3155);
and U9928 (N_9928,In_1941,In_1130);
nor U9929 (N_9929,In_1245,In_2835);
or U9930 (N_9930,In_77,In_4796);
xor U9931 (N_9931,In_1701,In_3781);
and U9932 (N_9932,In_2403,In_4992);
nand U9933 (N_9933,In_2019,In_4220);
nand U9934 (N_9934,In_2423,In_3534);
xor U9935 (N_9935,In_2354,In_251);
or U9936 (N_9936,In_4242,In_1086);
nor U9937 (N_9937,In_1211,In_3788);
xor U9938 (N_9938,In_2560,In_2484);
nand U9939 (N_9939,In_1681,In_4893);
nand U9940 (N_9940,In_1794,In_1663);
and U9941 (N_9941,In_3066,In_4052);
nand U9942 (N_9942,In_694,In_527);
and U9943 (N_9943,In_746,In_2906);
nand U9944 (N_9944,In_493,In_3544);
nand U9945 (N_9945,In_917,In_2143);
xnor U9946 (N_9946,In_3551,In_1315);
xor U9947 (N_9947,In_2600,In_504);
or U9948 (N_9948,In_1418,In_3896);
or U9949 (N_9949,In_3630,In_321);
and U9950 (N_9950,In_2213,In_2271);
and U9951 (N_9951,In_538,In_3329);
and U9952 (N_9952,In_2021,In_4522);
xnor U9953 (N_9953,In_4216,In_4325);
or U9954 (N_9954,In_2399,In_141);
nand U9955 (N_9955,In_215,In_2408);
or U9956 (N_9956,In_4462,In_4053);
nor U9957 (N_9957,In_2192,In_308);
nand U9958 (N_9958,In_1295,In_1906);
and U9959 (N_9959,In_4785,In_4845);
xnor U9960 (N_9960,In_2697,In_3601);
and U9961 (N_9961,In_3574,In_2987);
or U9962 (N_9962,In_3350,In_2447);
and U9963 (N_9963,In_3508,In_2562);
and U9964 (N_9964,In_582,In_1779);
and U9965 (N_9965,In_4854,In_1903);
nand U9966 (N_9966,In_2072,In_1610);
nand U9967 (N_9967,In_3522,In_605);
and U9968 (N_9968,In_1810,In_3358);
nand U9969 (N_9969,In_151,In_2154);
and U9970 (N_9970,In_1428,In_2684);
nand U9971 (N_9971,In_1072,In_3543);
and U9972 (N_9972,In_147,In_3217);
xor U9973 (N_9973,In_4270,In_527);
or U9974 (N_9974,In_133,In_3985);
and U9975 (N_9975,In_3599,In_1133);
or U9976 (N_9976,In_3338,In_1669);
or U9977 (N_9977,In_1968,In_4803);
xnor U9978 (N_9978,In_4396,In_1017);
nand U9979 (N_9979,In_107,In_3261);
xnor U9980 (N_9980,In_3714,In_580);
xnor U9981 (N_9981,In_3344,In_3450);
or U9982 (N_9982,In_3185,In_2509);
or U9983 (N_9983,In_4430,In_1973);
xor U9984 (N_9984,In_2222,In_303);
nor U9985 (N_9985,In_545,In_2214);
nor U9986 (N_9986,In_4721,In_370);
xor U9987 (N_9987,In_585,In_4126);
xnor U9988 (N_9988,In_1736,In_4868);
xor U9989 (N_9989,In_2700,In_3055);
and U9990 (N_9990,In_4680,In_4978);
or U9991 (N_9991,In_4565,In_3913);
xor U9992 (N_9992,In_3678,In_1735);
nor U9993 (N_9993,In_859,In_3482);
xnor U9994 (N_9994,In_36,In_2990);
nand U9995 (N_9995,In_3389,In_3233);
xor U9996 (N_9996,In_2212,In_1023);
and U9997 (N_9997,In_2888,In_551);
xor U9998 (N_9998,In_2022,In_1590);
nand U9999 (N_9999,In_3801,In_2509);
xnor U10000 (N_10000,N_590,N_3007);
or U10001 (N_10001,N_4391,N_5715);
nand U10002 (N_10002,N_358,N_1757);
nand U10003 (N_10003,N_2374,N_2948);
or U10004 (N_10004,N_7101,N_5335);
nor U10005 (N_10005,N_5919,N_3023);
nor U10006 (N_10006,N_6307,N_1772);
nand U10007 (N_10007,N_2113,N_4214);
nor U10008 (N_10008,N_9442,N_7660);
or U10009 (N_10009,N_9172,N_7842);
nor U10010 (N_10010,N_3450,N_9917);
or U10011 (N_10011,N_4922,N_2058);
and U10012 (N_10012,N_1175,N_803);
or U10013 (N_10013,N_4616,N_1500);
nand U10014 (N_10014,N_9905,N_6337);
nand U10015 (N_10015,N_3268,N_8122);
nor U10016 (N_10016,N_8287,N_635);
nor U10017 (N_10017,N_5490,N_6936);
nor U10018 (N_10018,N_9072,N_220);
and U10019 (N_10019,N_6122,N_3514);
and U10020 (N_10020,N_4625,N_5977);
xnor U10021 (N_10021,N_5750,N_6059);
and U10022 (N_10022,N_4373,N_9900);
and U10023 (N_10023,N_4550,N_7252);
and U10024 (N_10024,N_7197,N_2737);
nand U10025 (N_10025,N_9750,N_9018);
or U10026 (N_10026,N_537,N_4583);
xor U10027 (N_10027,N_2221,N_4547);
nand U10028 (N_10028,N_1965,N_343);
nor U10029 (N_10029,N_5430,N_957);
xnor U10030 (N_10030,N_2073,N_9711);
xor U10031 (N_10031,N_3530,N_15);
nor U10032 (N_10032,N_6147,N_5610);
and U10033 (N_10033,N_5488,N_6844);
or U10034 (N_10034,N_9594,N_5938);
xor U10035 (N_10035,N_7217,N_389);
nor U10036 (N_10036,N_3112,N_5535);
nand U10037 (N_10037,N_5954,N_7644);
nor U10038 (N_10038,N_3383,N_558);
and U10039 (N_10039,N_3274,N_3878);
nand U10040 (N_10040,N_8754,N_5662);
xnor U10041 (N_10041,N_1813,N_819);
nand U10042 (N_10042,N_2979,N_1047);
nor U10043 (N_10043,N_305,N_4406);
nor U10044 (N_10044,N_3697,N_2734);
nand U10045 (N_10045,N_3305,N_9187);
nor U10046 (N_10046,N_6159,N_1233);
nand U10047 (N_10047,N_9841,N_8386);
or U10048 (N_10048,N_6662,N_4417);
or U10049 (N_10049,N_5766,N_2750);
nor U10050 (N_10050,N_6322,N_3439);
nor U10051 (N_10051,N_118,N_4405);
or U10052 (N_10052,N_6983,N_8948);
nor U10053 (N_10053,N_8016,N_3942);
xor U10054 (N_10054,N_5136,N_5093);
xnor U10055 (N_10055,N_2436,N_1623);
nand U10056 (N_10056,N_6670,N_5146);
or U10057 (N_10057,N_5097,N_9955);
nand U10058 (N_10058,N_514,N_7773);
or U10059 (N_10059,N_1415,N_9358);
or U10060 (N_10060,N_8614,N_9873);
and U10061 (N_10061,N_1519,N_6206);
or U10062 (N_10062,N_9011,N_6016);
nor U10063 (N_10063,N_8739,N_3640);
or U10064 (N_10064,N_2447,N_4939);
nand U10065 (N_10065,N_9333,N_3216);
nor U10066 (N_10066,N_13,N_473);
nand U10067 (N_10067,N_4269,N_6861);
nand U10068 (N_10068,N_7940,N_5310);
xnor U10069 (N_10069,N_6341,N_3438);
and U10070 (N_10070,N_6990,N_7584);
or U10071 (N_10071,N_7485,N_9014);
xnor U10072 (N_10072,N_3582,N_9892);
and U10073 (N_10073,N_5680,N_1786);
nor U10074 (N_10074,N_7903,N_3080);
and U10075 (N_10075,N_4067,N_345);
nor U10076 (N_10076,N_594,N_8362);
nand U10077 (N_10077,N_2187,N_1379);
nand U10078 (N_10078,N_1144,N_2259);
or U10079 (N_10079,N_2205,N_9287);
nor U10080 (N_10080,N_1326,N_9648);
xor U10081 (N_10081,N_5753,N_4513);
xor U10082 (N_10082,N_9296,N_9528);
and U10083 (N_10083,N_4370,N_615);
or U10084 (N_10084,N_7027,N_5953);
xnor U10085 (N_10085,N_7672,N_4367);
or U10086 (N_10086,N_3277,N_3494);
nor U10087 (N_10087,N_6911,N_8758);
nor U10088 (N_10088,N_7016,N_2049);
and U10089 (N_10089,N_2014,N_9311);
or U10090 (N_10090,N_5171,N_5684);
xnor U10091 (N_10091,N_7099,N_1115);
nor U10092 (N_10092,N_6223,N_5131);
nand U10093 (N_10093,N_2983,N_692);
xor U10094 (N_10094,N_3453,N_6812);
xor U10095 (N_10095,N_7415,N_8067);
nor U10096 (N_10096,N_307,N_3498);
and U10097 (N_10097,N_9035,N_5264);
and U10098 (N_10098,N_1560,N_5621);
xnor U10099 (N_10099,N_6103,N_9874);
and U10100 (N_10100,N_8012,N_5914);
nand U10101 (N_10101,N_8908,N_7215);
and U10102 (N_10102,N_1961,N_1774);
nand U10103 (N_10103,N_3072,N_1354);
nand U10104 (N_10104,N_3721,N_2477);
nor U10105 (N_10105,N_7618,N_1896);
nand U10106 (N_10106,N_9719,N_3234);
xnor U10107 (N_10107,N_8609,N_6187);
and U10108 (N_10108,N_297,N_7708);
nand U10109 (N_10109,N_409,N_8606);
nor U10110 (N_10110,N_8280,N_4908);
and U10111 (N_10111,N_7780,N_7130);
nor U10112 (N_10112,N_526,N_7715);
xnor U10113 (N_10113,N_7854,N_5137);
nor U10114 (N_10114,N_9469,N_1974);
and U10115 (N_10115,N_7952,N_1223);
xor U10116 (N_10116,N_9978,N_5786);
nor U10117 (N_10117,N_7668,N_3435);
or U10118 (N_10118,N_6344,N_8451);
and U10119 (N_10119,N_5456,N_1750);
xnor U10120 (N_10120,N_2284,N_8681);
or U10121 (N_10121,N_528,N_3066);
xor U10122 (N_10122,N_7566,N_1240);
nand U10123 (N_10123,N_8987,N_9151);
or U10124 (N_10124,N_9268,N_3114);
xnor U10125 (N_10125,N_6919,N_4027);
nand U10126 (N_10126,N_4945,N_7435);
and U10127 (N_10127,N_9045,N_6826);
and U10128 (N_10128,N_5364,N_5757);
nor U10129 (N_10129,N_6247,N_6849);
xor U10130 (N_10130,N_4867,N_9419);
nand U10131 (N_10131,N_5832,N_458);
and U10132 (N_10132,N_5036,N_3143);
or U10133 (N_10133,N_7491,N_7790);
nor U10134 (N_10134,N_481,N_4895);
or U10135 (N_10135,N_269,N_1893);
nand U10136 (N_10136,N_3533,N_5679);
nor U10137 (N_10137,N_8194,N_1990);
nand U10138 (N_10138,N_3712,N_6809);
or U10139 (N_10139,N_1296,N_9846);
or U10140 (N_10140,N_4471,N_9183);
xor U10141 (N_10141,N_9027,N_4551);
nand U10142 (N_10142,N_6415,N_7983);
or U10143 (N_10143,N_1709,N_2346);
nor U10144 (N_10144,N_8111,N_9694);
xnor U10145 (N_10145,N_9756,N_5507);
xnor U10146 (N_10146,N_9833,N_3454);
nor U10147 (N_10147,N_1833,N_9348);
nand U10148 (N_10148,N_6981,N_2790);
xor U10149 (N_10149,N_3356,N_9844);
or U10150 (N_10150,N_6044,N_4495);
xor U10151 (N_10151,N_3681,N_8811);
and U10152 (N_10152,N_7034,N_5439);
nand U10153 (N_10153,N_3018,N_3748);
nor U10154 (N_10154,N_5319,N_3009);
nor U10155 (N_10155,N_1459,N_240);
and U10156 (N_10156,N_3008,N_3089);
or U10157 (N_10157,N_7817,N_8581);
nor U10158 (N_10158,N_1673,N_9610);
or U10159 (N_10159,N_9328,N_4745);
and U10160 (N_10160,N_4851,N_1465);
or U10161 (N_10161,N_9357,N_49);
or U10162 (N_10162,N_9332,N_69);
xor U10163 (N_10163,N_2548,N_6719);
or U10164 (N_10164,N_1116,N_4138);
or U10165 (N_10165,N_5215,N_5699);
and U10166 (N_10166,N_3281,N_9486);
and U10167 (N_10167,N_7126,N_237);
and U10168 (N_10168,N_7918,N_153);
and U10169 (N_10169,N_1551,N_5024);
and U10170 (N_10170,N_4469,N_6660);
nor U10171 (N_10171,N_893,N_2458);
nor U10172 (N_10172,N_1511,N_644);
nor U10173 (N_10173,N_6342,N_5934);
nor U10174 (N_10174,N_7813,N_785);
nand U10175 (N_10175,N_7797,N_8544);
nand U10176 (N_10176,N_5927,N_8215);
nand U10177 (N_10177,N_1764,N_1302);
or U10178 (N_10178,N_3367,N_7527);
and U10179 (N_10179,N_7581,N_2672);
xor U10180 (N_10180,N_2903,N_3192);
xnor U10181 (N_10181,N_5401,N_6186);
and U10182 (N_10182,N_4000,N_2044);
nor U10183 (N_10183,N_1928,N_6758);
and U10184 (N_10184,N_758,N_3586);
and U10185 (N_10185,N_1298,N_8075);
xnor U10186 (N_10186,N_6182,N_5880);
and U10187 (N_10187,N_5465,N_6293);
nor U10188 (N_10188,N_1315,N_5744);
xnor U10189 (N_10189,N_199,N_6105);
xor U10190 (N_10190,N_2765,N_9150);
nand U10191 (N_10191,N_5170,N_7592);
xor U10192 (N_10192,N_8181,N_2461);
nor U10193 (N_10193,N_1044,N_4688);
nor U10194 (N_10194,N_5645,N_3391);
xnor U10195 (N_10195,N_751,N_1275);
nor U10196 (N_10196,N_1962,N_175);
nand U10197 (N_10197,N_7506,N_7171);
xor U10198 (N_10198,N_1858,N_6237);
and U10199 (N_10199,N_5257,N_3529);
xnor U10200 (N_10200,N_914,N_7320);
and U10201 (N_10201,N_8186,N_7191);
and U10202 (N_10202,N_9670,N_6906);
and U10203 (N_10203,N_283,N_844);
nand U10204 (N_10204,N_715,N_8588);
nand U10205 (N_10205,N_8178,N_5790);
nor U10206 (N_10206,N_3412,N_1052);
or U10207 (N_10207,N_9732,N_3934);
and U10208 (N_10208,N_6638,N_4894);
nand U10209 (N_10209,N_5182,N_7315);
or U10210 (N_10210,N_8636,N_9920);
xnor U10211 (N_10211,N_8116,N_7489);
xor U10212 (N_10212,N_410,N_6822);
nor U10213 (N_10213,N_3132,N_9208);
nor U10214 (N_10214,N_9281,N_4170);
xnor U10215 (N_10215,N_825,N_2176);
or U10216 (N_10216,N_8951,N_7728);
nand U10217 (N_10217,N_5932,N_4629);
and U10218 (N_10218,N_9827,N_3146);
nand U10219 (N_10219,N_399,N_7530);
and U10220 (N_10220,N_2364,N_2762);
or U10221 (N_10221,N_5886,N_1518);
nor U10222 (N_10222,N_545,N_9201);
nand U10223 (N_10223,N_614,N_2587);
nor U10224 (N_10224,N_2572,N_8395);
nor U10225 (N_10225,N_6360,N_3799);
and U10226 (N_10226,N_6878,N_2571);
and U10227 (N_10227,N_9983,N_9205);
or U10228 (N_10228,N_6114,N_9365);
or U10229 (N_10229,N_365,N_8697);
and U10230 (N_10230,N_4504,N_7949);
or U10231 (N_10231,N_1871,N_6284);
nor U10232 (N_10232,N_4549,N_6495);
or U10233 (N_10233,N_1823,N_8808);
nor U10234 (N_10234,N_9310,N_7440);
or U10235 (N_10235,N_7685,N_9293);
or U10236 (N_10236,N_2839,N_7310);
or U10237 (N_10237,N_189,N_4892);
or U10238 (N_10238,N_598,N_1508);
and U10239 (N_10239,N_6586,N_2094);
and U10240 (N_10240,N_717,N_3695);
xnor U10241 (N_10241,N_3816,N_1700);
nand U10242 (N_10242,N_2151,N_1129);
nand U10243 (N_10243,N_1466,N_3403);
and U10244 (N_10244,N_9555,N_649);
nor U10245 (N_10245,N_9468,N_2303);
nand U10246 (N_10246,N_2636,N_16);
nor U10247 (N_10247,N_8110,N_8323);
xnor U10248 (N_10248,N_584,N_2013);
xnor U10249 (N_10249,N_9288,N_1916);
and U10250 (N_10250,N_1314,N_1978);
nand U10251 (N_10251,N_6302,N_6332);
nor U10252 (N_10252,N_7501,N_764);
and U10253 (N_10253,N_2833,N_7718);
nor U10254 (N_10254,N_2862,N_6995);
nand U10255 (N_10255,N_4208,N_6816);
nand U10256 (N_10256,N_9508,N_2615);
and U10257 (N_10257,N_4252,N_2656);
and U10258 (N_10258,N_7233,N_5613);
xnor U10259 (N_10259,N_1093,N_4213);
xnor U10260 (N_10260,N_9093,N_6250);
or U10261 (N_10261,N_2626,N_1413);
and U10262 (N_10262,N_147,N_1731);
nand U10263 (N_10263,N_7412,N_3945);
xor U10264 (N_10264,N_517,N_8664);
xor U10265 (N_10265,N_9678,N_6417);
and U10266 (N_10266,N_9532,N_8611);
xnor U10267 (N_10267,N_723,N_1096);
and U10268 (N_10268,N_8521,N_8649);
xor U10269 (N_10269,N_6007,N_7703);
nor U10270 (N_10270,N_1967,N_7755);
nor U10271 (N_10271,N_3730,N_5411);
xnor U10272 (N_10272,N_8780,N_7284);
nand U10273 (N_10273,N_4730,N_1783);
and U10274 (N_10274,N_7053,N_5126);
nand U10275 (N_10275,N_5628,N_2699);
and U10276 (N_10276,N_166,N_4496);
xnor U10277 (N_10277,N_3488,N_6492);
xor U10278 (N_10278,N_994,N_333);
xnor U10279 (N_10279,N_8904,N_63);
xnor U10280 (N_10280,N_4147,N_2373);
nand U10281 (N_10281,N_898,N_2499);
xnor U10282 (N_10282,N_7505,N_9659);
or U10283 (N_10283,N_9485,N_7097);
xnor U10284 (N_10284,N_7182,N_3421);
xor U10285 (N_10285,N_1311,N_6760);
xor U10286 (N_10286,N_2122,N_2555);
nor U10287 (N_10287,N_3986,N_603);
nand U10288 (N_10288,N_8394,N_6209);
xnor U10289 (N_10289,N_1472,N_1086);
nor U10290 (N_10290,N_8199,N_5225);
or U10291 (N_10291,N_4979,N_7855);
nor U10292 (N_10292,N_7067,N_293);
nor U10293 (N_10293,N_5768,N_8434);
nand U10294 (N_10294,N_7555,N_8410);
nor U10295 (N_10295,N_6508,N_5139);
nand U10296 (N_10296,N_2085,N_9086);
nand U10297 (N_10297,N_9099,N_4489);
nor U10298 (N_10298,N_6072,N_2133);
nor U10299 (N_10299,N_9117,N_1778);
or U10300 (N_10300,N_472,N_9336);
xor U10301 (N_10301,N_4320,N_2334);
nand U10302 (N_10302,N_6125,N_1549);
or U10303 (N_10303,N_7828,N_7492);
xnor U10304 (N_10304,N_314,N_8331);
or U10305 (N_10305,N_727,N_3394);
and U10306 (N_10306,N_7049,N_4742);
nor U10307 (N_10307,N_2383,N_5177);
xor U10308 (N_10308,N_4186,N_7343);
nor U10309 (N_10309,N_3223,N_8349);
nand U10310 (N_10310,N_7932,N_6241);
nand U10311 (N_10311,N_2271,N_4412);
nand U10312 (N_10312,N_5788,N_836);
nand U10313 (N_10313,N_1534,N_7590);
or U10314 (N_10314,N_8034,N_5643);
or U10315 (N_10315,N_6633,N_5890);
and U10316 (N_10316,N_8656,N_120);
or U10317 (N_10317,N_8932,N_7963);
nand U10318 (N_10318,N_5818,N_2584);
and U10319 (N_10319,N_625,N_5062);
or U10320 (N_10320,N_9292,N_601);
nor U10321 (N_10321,N_7168,N_6315);
nor U10322 (N_10322,N_7470,N_3914);
nor U10323 (N_10323,N_2460,N_6974);
nand U10324 (N_10324,N_8982,N_6248);
nand U10325 (N_10325,N_178,N_5326);
nand U10326 (N_10326,N_779,N_3536);
or U10327 (N_10327,N_7086,N_7464);
or U10328 (N_10328,N_4256,N_6326);
nor U10329 (N_10329,N_6409,N_4791);
xor U10330 (N_10330,N_2008,N_9621);
nand U10331 (N_10331,N_3041,N_5227);
xnor U10332 (N_10332,N_9974,N_7852);
and U10333 (N_10333,N_5553,N_1132);
nand U10334 (N_10334,N_7239,N_2649);
nor U10335 (N_10335,N_8081,N_9182);
or U10336 (N_10336,N_4007,N_4578);
nor U10337 (N_10337,N_7712,N_6785);
nor U10338 (N_10338,N_3155,N_8984);
nand U10339 (N_10339,N_4703,N_1167);
nor U10340 (N_10340,N_52,N_3167);
xnor U10341 (N_10341,N_5503,N_2134);
and U10342 (N_10342,N_2479,N_5314);
nand U10343 (N_10343,N_8615,N_9097);
nor U10344 (N_10344,N_5244,N_5362);
and U10345 (N_10345,N_6138,N_7976);
and U10346 (N_10346,N_8840,N_2442);
xnor U10347 (N_10347,N_8393,N_9466);
or U10348 (N_10348,N_8831,N_8930);
nand U10349 (N_10349,N_5591,N_7561);
and U10350 (N_10350,N_1147,N_4961);
or U10351 (N_10351,N_1590,N_2585);
or U10352 (N_10352,N_9590,N_4064);
or U10353 (N_10353,N_5917,N_464);
nor U10354 (N_10354,N_9586,N_8241);
or U10355 (N_10355,N_2145,N_2298);
and U10356 (N_10356,N_4967,N_2998);
nor U10357 (N_10357,N_2405,N_7975);
or U10358 (N_10358,N_8103,N_5506);
nor U10359 (N_10359,N_5254,N_6454);
nand U10360 (N_10360,N_3795,N_8712);
xor U10361 (N_10361,N_3145,N_8715);
and U10362 (N_10362,N_9735,N_9138);
and U10363 (N_10363,N_6972,N_5915);
nand U10364 (N_10364,N_5756,N_684);
xor U10365 (N_10365,N_5212,N_5395);
or U10366 (N_10366,N_8525,N_9580);
nand U10367 (N_10367,N_8628,N_5267);
nor U10368 (N_10368,N_8452,N_3701);
or U10369 (N_10369,N_5423,N_418);
and U10370 (N_10370,N_6874,N_3366);
nand U10371 (N_10371,N_7298,N_9828);
or U10372 (N_10372,N_1140,N_9647);
nor U10373 (N_10373,N_3059,N_1800);
nand U10374 (N_10374,N_2067,N_7871);
nor U10375 (N_10375,N_4805,N_3437);
xnor U10376 (N_10376,N_84,N_8028);
or U10377 (N_10377,N_9990,N_7811);
xor U10378 (N_10378,N_3840,N_8756);
nor U10379 (N_10379,N_2234,N_7178);
nor U10380 (N_10380,N_3344,N_460);
nor U10381 (N_10381,N_1966,N_802);
or U10382 (N_10382,N_6458,N_5622);
and U10383 (N_10383,N_5900,N_9509);
and U10384 (N_10384,N_6452,N_890);
xor U10385 (N_10385,N_209,N_8600);
nor U10386 (N_10386,N_5285,N_1707);
nor U10387 (N_10387,N_7570,N_4997);
xnor U10388 (N_10388,N_6652,N_7895);
or U10389 (N_10389,N_5547,N_9388);
nor U10390 (N_10390,N_4907,N_6355);
xor U10391 (N_10391,N_8257,N_8979);
or U10392 (N_10392,N_2798,N_6519);
or U10393 (N_10393,N_2939,N_8747);
and U10394 (N_10394,N_6957,N_8476);
nor U10395 (N_10395,N_8316,N_933);
xor U10396 (N_10396,N_7972,N_3219);
and U10397 (N_10397,N_1815,N_8926);
and U10398 (N_10398,N_7410,N_4746);
or U10399 (N_10399,N_8850,N_8643);
nand U10400 (N_10400,N_9375,N_619);
nand U10401 (N_10401,N_1826,N_3452);
nand U10402 (N_10402,N_5677,N_7694);
or U10403 (N_10403,N_9574,N_8854);
nor U10404 (N_10404,N_1148,N_8813);
or U10405 (N_10405,N_7833,N_1934);
xnor U10406 (N_10406,N_4649,N_883);
nand U10407 (N_10407,N_5731,N_422);
and U10408 (N_10408,N_3989,N_6202);
or U10409 (N_10409,N_1489,N_2003);
or U10410 (N_10410,N_5425,N_7772);
xnor U10411 (N_10411,N_2770,N_6163);
and U10412 (N_10412,N_4998,N_8722);
nand U10413 (N_10413,N_2116,N_9588);
or U10414 (N_10414,N_6265,N_8304);
and U10415 (N_10415,N_8219,N_813);
nor U10416 (N_10416,N_9726,N_6889);
and U10417 (N_10417,N_1881,N_2789);
and U10418 (N_10418,N_3195,N_7756);
and U10419 (N_10419,N_5438,N_4721);
nand U10420 (N_10420,N_6087,N_3778);
nand U10421 (N_10421,N_3347,N_6065);
nand U10422 (N_10422,N_8013,N_7025);
and U10423 (N_10423,N_3246,N_7229);
and U10424 (N_10424,N_9262,N_5164);
xnor U10425 (N_10425,N_936,N_2716);
xnor U10426 (N_10426,N_2439,N_1758);
xor U10427 (N_10427,N_4592,N_1727);
nor U10428 (N_10428,N_7848,N_6493);
and U10429 (N_10429,N_3897,N_702);
nand U10430 (N_10430,N_9370,N_9767);
nand U10431 (N_10431,N_6353,N_6965);
nor U10432 (N_10432,N_162,N_3233);
xor U10433 (N_10433,N_7427,N_2752);
nor U10434 (N_10434,N_8235,N_9884);
xor U10435 (N_10435,N_6870,N_5966);
nor U10436 (N_10436,N_4807,N_6742);
and U10437 (N_10437,N_8245,N_4457);
nor U10438 (N_10438,N_4679,N_2472);
or U10439 (N_10439,N_6023,N_1292);
or U10440 (N_10440,N_7846,N_9077);
or U10441 (N_10441,N_8557,N_2118);
nand U10442 (N_10442,N_4891,N_9526);
or U10443 (N_10443,N_3621,N_5612);
nand U10444 (N_10444,N_3098,N_4789);
and U10445 (N_10445,N_3263,N_6102);
and U10446 (N_10446,N_1343,N_6388);
or U10447 (N_10447,N_3961,N_1122);
or U10448 (N_10448,N_1887,N_7847);
nand U10449 (N_10449,N_6455,N_91);
xor U10450 (N_10450,N_2412,N_2466);
nand U10451 (N_10451,N_5711,N_732);
xor U10452 (N_10452,N_3829,N_2288);
and U10453 (N_10453,N_8140,N_5572);
nor U10454 (N_10454,N_578,N_7341);
and U10455 (N_10455,N_4983,N_1293);
nand U10456 (N_10456,N_3655,N_8915);
nand U10457 (N_10457,N_1937,N_2285);
nand U10458 (N_10458,N_2257,N_1564);
nand U10459 (N_10459,N_8786,N_9277);
nand U10460 (N_10460,N_9992,N_2146);
xor U10461 (N_10461,N_2300,N_8734);
nand U10462 (N_10462,N_8517,N_9229);
and U10463 (N_10463,N_4350,N_258);
xnor U10464 (N_10464,N_6278,N_4283);
and U10465 (N_10465,N_6430,N_316);
nor U10466 (N_10466,N_7122,N_6160);
or U10467 (N_10467,N_1621,N_7368);
nand U10468 (N_10468,N_6435,N_9209);
nand U10469 (N_10469,N_9657,N_3976);
nor U10470 (N_10470,N_2805,N_6323);
xor U10471 (N_10471,N_4875,N_2247);
or U10472 (N_10472,N_5010,N_907);
nand U10473 (N_10473,N_9455,N_5482);
nand U10474 (N_10474,N_2806,N_3821);
nor U10475 (N_10475,N_6563,N_321);
and U10476 (N_10476,N_9959,N_2821);
xor U10477 (N_10477,N_4317,N_6759);
nand U10478 (N_10478,N_9351,N_882);
or U10479 (N_10479,N_3339,N_737);
nand U10480 (N_10480,N_8274,N_6609);
xnor U10481 (N_10481,N_7682,N_8425);
or U10482 (N_10482,N_2494,N_4397);
nor U10483 (N_10483,N_1171,N_3544);
nor U10484 (N_10484,N_5947,N_77);
or U10485 (N_10485,N_5467,N_5841);
and U10486 (N_10486,N_7657,N_8164);
and U10487 (N_10487,N_9251,N_9169);
or U10488 (N_10488,N_100,N_784);
nand U10489 (N_10489,N_908,N_3979);
and U10490 (N_10490,N_8085,N_3372);
nand U10491 (N_10491,N_5193,N_122);
nand U10492 (N_10492,N_279,N_5123);
and U10493 (N_10493,N_5476,N_4624);
xor U10494 (N_10494,N_2242,N_4254);
nand U10495 (N_10495,N_9289,N_5592);
xnor U10496 (N_10496,N_6646,N_6041);
and U10497 (N_10497,N_561,N_1756);
and U10498 (N_10498,N_1403,N_8101);
or U10499 (N_10499,N_2385,N_2427);
or U10500 (N_10500,N_5210,N_7236);
and U10501 (N_10501,N_6015,N_1127);
and U10502 (N_10502,N_9489,N_5400);
or U10503 (N_10503,N_9671,N_9677);
or U10504 (N_10504,N_6200,N_9108);
and U10505 (N_10505,N_4190,N_5197);
or U10506 (N_10506,N_6530,N_4438);
nor U10507 (N_10507,N_5992,N_7861);
xor U10508 (N_10508,N_3725,N_2504);
and U10509 (N_10509,N_7532,N_8379);
or U10510 (N_10510,N_7212,N_7115);
xor U10511 (N_10511,N_9710,N_1531);
and U10512 (N_10512,N_7992,N_7798);
xnor U10513 (N_10513,N_6650,N_7008);
nand U10514 (N_10514,N_4300,N_8318);
and U10515 (N_10515,N_9459,N_2199);
and U10516 (N_10516,N_1532,N_8743);
and U10517 (N_10517,N_1824,N_7782);
or U10518 (N_10518,N_3430,N_7907);
xor U10519 (N_10519,N_6386,N_9156);
or U10520 (N_10520,N_2888,N_6988);
xnor U10521 (N_10521,N_7373,N_4106);
or U10522 (N_10522,N_4279,N_9561);
nand U10523 (N_10523,N_1514,N_8232);
nor U10524 (N_10524,N_1168,N_3568);
xor U10525 (N_10525,N_3165,N_6941);
or U10526 (N_10526,N_6205,N_2712);
nor U10527 (N_10527,N_9931,N_8853);
nor U10528 (N_10528,N_1570,N_3519);
nor U10529 (N_10529,N_2689,N_5402);
and U10530 (N_10530,N_5047,N_131);
or U10531 (N_10531,N_1036,N_1796);
or U10532 (N_10532,N_6659,N_9786);
nor U10533 (N_10533,N_5811,N_8849);
or U10534 (N_10534,N_1988,N_5039);
nand U10535 (N_10535,N_5153,N_4402);
nor U10536 (N_10536,N_6158,N_565);
or U10537 (N_10537,N_3176,N_8817);
and U10538 (N_10538,N_7075,N_3447);
xor U10539 (N_10539,N_6828,N_2627);
nor U10540 (N_10540,N_46,N_4392);
xnor U10541 (N_10541,N_5236,N_6599);
and U10542 (N_10542,N_2827,N_2224);
nor U10543 (N_10543,N_3938,N_7098);
and U10544 (N_10544,N_6133,N_2529);
or U10545 (N_10545,N_824,N_2139);
nor U10546 (N_10546,N_4611,N_8036);
or U10547 (N_10547,N_4498,N_7020);
and U10548 (N_10548,N_8157,N_397);
nand U10549 (N_10549,N_7981,N_6642);
xnor U10550 (N_10550,N_7249,N_5732);
xor U10551 (N_10551,N_6776,N_4034);
or U10552 (N_10552,N_3658,N_4015);
xnor U10553 (N_10553,N_5183,N_9241);
nand U10554 (N_10554,N_9971,N_2226);
xnor U10555 (N_10555,N_7244,N_6286);
nand U10556 (N_10556,N_407,N_3014);
and U10557 (N_10557,N_3699,N_210);
xor U10558 (N_10558,N_3483,N_7795);
or U10559 (N_10559,N_7863,N_1630);
xor U10560 (N_10560,N_4662,N_1062);
xor U10561 (N_10561,N_2108,N_609);
nand U10562 (N_10562,N_3033,N_434);
nand U10563 (N_10563,N_7185,N_2419);
and U10564 (N_10564,N_4752,N_2976);
nand U10565 (N_10565,N_4607,N_4435);
nand U10566 (N_10566,N_7942,N_3972);
or U10567 (N_10567,N_3370,N_7063);
and U10568 (N_10568,N_695,N_745);
and U10569 (N_10569,N_7328,N_7404);
nor U10570 (N_10570,N_6077,N_7493);
nor U10571 (N_10571,N_750,N_3502);
xor U10572 (N_10572,N_4385,N_1393);
nand U10573 (N_10573,N_3857,N_467);
nor U10574 (N_10574,N_8065,N_4839);
nand U10575 (N_10575,N_2550,N_2832);
and U10576 (N_10576,N_1559,N_7796);
or U10577 (N_10577,N_1153,N_7308);
and U10578 (N_10578,N_776,N_843);
xnor U10579 (N_10579,N_1087,N_3111);
nand U10580 (N_10580,N_330,N_6526);
nand U10581 (N_10581,N_8418,N_1577);
and U10582 (N_10582,N_9912,N_5845);
or U10583 (N_10583,N_5050,N_2476);
nand U10584 (N_10584,N_4445,N_3011);
nand U10585 (N_10585,N_7752,N_797);
and U10586 (N_10586,N_6212,N_721);
xor U10587 (N_10587,N_5971,N_2808);
xnor U10588 (N_10588,N_4856,N_2886);
or U10589 (N_10589,N_477,N_5195);
xnor U10590 (N_10590,N_2793,N_8574);
nor U10591 (N_10591,N_5976,N_5445);
and U10592 (N_10592,N_2055,N_996);
or U10593 (N_10593,N_7413,N_4131);
nand U10594 (N_10594,N_7525,N_197);
nand U10595 (N_10595,N_3707,N_5865);
or U10596 (N_10596,N_9910,N_1976);
xor U10597 (N_10597,N_5325,N_7367);
nor U10598 (N_10598,N_6850,N_9948);
nor U10599 (N_10599,N_7457,N_9755);
and U10600 (N_10600,N_6305,N_4656);
or U10601 (N_10601,N_8233,N_2966);
or U10602 (N_10602,N_6153,N_6291);
xnor U10603 (N_10603,N_3136,N_1189);
and U10604 (N_10604,N_977,N_5330);
nand U10605 (N_10605,N_9502,N_3485);
nand U10606 (N_10606,N_7022,N_5200);
or U10607 (N_10607,N_2202,N_3204);
and U10608 (N_10608,N_2528,N_5031);
and U10609 (N_10609,N_8298,N_538);
nor U10610 (N_10610,N_4073,N_5801);
or U10611 (N_10611,N_2840,N_292);
xor U10612 (N_10612,N_2060,N_6413);
nand U10613 (N_10613,N_6256,N_3302);
and U10614 (N_10614,N_4126,N_9361);
nor U10615 (N_10615,N_5410,N_9359);
nor U10616 (N_10616,N_1899,N_3675);
or U10617 (N_10617,N_4816,N_3814);
nor U10618 (N_10618,N_9123,N_9503);
xor U10619 (N_10619,N_4292,N_8490);
nor U10620 (N_10620,N_8498,N_8935);
and U10621 (N_10621,N_9772,N_1377);
or U10622 (N_10622,N_6523,N_2204);
nor U10623 (N_10623,N_7741,N_7814);
nand U10624 (N_10624,N_2150,N_7356);
and U10625 (N_10625,N_966,N_3160);
and U10626 (N_10626,N_1540,N_3528);
xor U10627 (N_10627,N_4880,N_4570);
nor U10628 (N_10628,N_2953,N_1640);
nand U10629 (N_10629,N_1432,N_5484);
nor U10630 (N_10630,N_653,N_5155);
nand U10631 (N_10631,N_3758,N_6687);
or U10632 (N_10632,N_4904,N_1117);
or U10633 (N_10633,N_642,N_1777);
and U10634 (N_10634,N_1475,N_7611);
xnor U10635 (N_10635,N_5656,N_4796);
or U10636 (N_10636,N_177,N_5304);
nor U10637 (N_10637,N_6000,N_1324);
nor U10638 (N_10638,N_3107,N_8568);
nor U10639 (N_10639,N_4520,N_5946);
xor U10640 (N_10640,N_1694,N_8254);
nand U10641 (N_10641,N_3682,N_56);
or U10642 (N_10642,N_2917,N_9167);
nor U10643 (N_10643,N_4331,N_8259);
nor U10644 (N_10644,N_2648,N_8376);
nand U10645 (N_10645,N_8768,N_3491);
and U10646 (N_10646,N_892,N_8744);
or U10647 (N_10647,N_2153,N_9052);
xor U10648 (N_10648,N_2381,N_7395);
or U10649 (N_10649,N_3270,N_7390);
nor U10650 (N_10650,N_6270,N_9674);
xnor U10651 (N_10651,N_1991,N_4650);
or U10652 (N_10652,N_4817,N_298);
nand U10653 (N_10653,N_3292,N_725);
xor U10654 (N_10654,N_3134,N_8934);
nand U10655 (N_10655,N_9661,N_6274);
and U10656 (N_10656,N_3024,N_9128);
or U10657 (N_10657,N_6335,N_8227);
and U10658 (N_10658,N_2331,N_4051);
nand U10659 (N_10659,N_8303,N_5831);
xnor U10660 (N_10660,N_960,N_432);
xnor U10661 (N_10661,N_999,N_479);
or U10662 (N_10662,N_6180,N_4597);
xnor U10663 (N_10663,N_7749,N_6425);
xor U10664 (N_10664,N_8185,N_6569);
and U10665 (N_10665,N_6804,N_4026);
nand U10666 (N_10666,N_6005,N_5975);
and U10667 (N_10667,N_7962,N_6537);
nor U10668 (N_10668,N_8991,N_2024);
xor U10669 (N_10669,N_1536,N_2090);
or U10670 (N_10670,N_4451,N_6369);
nor U10671 (N_10671,N_2639,N_8570);
xor U10672 (N_10672,N_3660,N_9338);
xnor U10673 (N_10673,N_8753,N_620);
and U10674 (N_10674,N_7524,N_1023);
nand U10675 (N_10675,N_2543,N_4665);
nor U10676 (N_10676,N_7656,N_9320);
or U10677 (N_10677,N_6833,N_4844);
nand U10678 (N_10678,N_6439,N_2913);
or U10679 (N_10679,N_1555,N_7921);
and U10680 (N_10680,N_682,N_3627);
nand U10681 (N_10681,N_5246,N_568);
and U10682 (N_10682,N_2777,N_9222);
or U10683 (N_10683,N_4352,N_4127);
nor U10684 (N_10684,N_1625,N_6310);
and U10685 (N_10685,N_2600,N_8735);
nand U10686 (N_10686,N_4116,N_1769);
xnor U10687 (N_10687,N_9126,N_2465);
nand U10688 (N_10688,N_5279,N_9302);
or U10689 (N_10689,N_9626,N_5663);
xnor U10690 (N_10690,N_6479,N_3873);
and U10691 (N_10691,N_4295,N_2158);
or U10692 (N_10692,N_9460,N_3249);
nor U10693 (N_10693,N_6648,N_72);
and U10694 (N_10694,N_3998,N_6422);
nor U10695 (N_10695,N_2229,N_991);
or U10696 (N_10696,N_1773,N_7118);
nor U10697 (N_10697,N_1521,N_6014);
or U10698 (N_10698,N_3194,N_1571);
or U10699 (N_10699,N_4973,N_5898);
nand U10700 (N_10700,N_8532,N_6451);
xnor U10701 (N_10701,N_2606,N_7735);
and U10702 (N_10702,N_9452,N_8914);
nand U10703 (N_10703,N_1479,N_359);
nand U10704 (N_10704,N_820,N_3404);
nor U10705 (N_10705,N_7339,N_2359);
xnor U10706 (N_10706,N_478,N_9084);
and U10707 (N_10707,N_6703,N_3571);
or U10708 (N_10708,N_3074,N_408);
nand U10709 (N_10709,N_3045,N_962);
nand U10710 (N_10710,N_9991,N_7338);
or U10711 (N_10711,N_6933,N_752);
xnor U10712 (N_10712,N_1619,N_264);
xor U10713 (N_10713,N_4840,N_9422);
or U10714 (N_10714,N_494,N_4809);
xnor U10715 (N_10715,N_7528,N_6379);
and U10716 (N_10716,N_1533,N_2809);
nand U10717 (N_10717,N_287,N_3933);
or U10718 (N_10718,N_1771,N_311);
or U10719 (N_10719,N_6637,N_9865);
nand U10720 (N_10720,N_5113,N_2698);
and U10721 (N_10721,N_6285,N_8839);
xnor U10722 (N_10722,N_2829,N_70);
nor U10723 (N_10723,N_5196,N_1002);
nand U10724 (N_10724,N_8941,N_7956);
xor U10725 (N_10725,N_4778,N_3638);
xor U10726 (N_10726,N_1431,N_2182);
and U10727 (N_10727,N_9542,N_8020);
or U10728 (N_10728,N_944,N_738);
nor U10729 (N_10729,N_4784,N_4680);
xor U10730 (N_10730,N_5986,N_2391);
nor U10731 (N_10731,N_9471,N_847);
xnor U10732 (N_10732,N_9109,N_107);
nand U10733 (N_10733,N_3684,N_2842);
xor U10734 (N_10734,N_9386,N_2490);
and U10735 (N_10735,N_7475,N_792);
or U10736 (N_10736,N_7238,N_9491);
and U10737 (N_10737,N_700,N_78);
and U10738 (N_10738,N_1434,N_3225);
xnor U10739 (N_10739,N_9438,N_1425);
xor U10740 (N_10740,N_8842,N_9953);
xnor U10741 (N_10741,N_846,N_7700);
and U10742 (N_10742,N_7585,N_7727);
or U10743 (N_10743,N_2893,N_276);
nor U10744 (N_10744,N_5119,N_5338);
or U10745 (N_10745,N_236,N_3713);
nand U10746 (N_10746,N_4797,N_5867);
xor U10747 (N_10747,N_3200,N_4847);
nand U10748 (N_10748,N_2254,N_8988);
nor U10749 (N_10749,N_1239,N_1552);
or U10750 (N_10750,N_9023,N_6946);
nor U10751 (N_10751,N_3461,N_4179);
and U10752 (N_10752,N_8052,N_9313);
nand U10753 (N_10753,N_8936,N_9856);
or U10754 (N_10754,N_6068,N_8213);
or U10755 (N_10755,N_8420,N_4461);
nor U10756 (N_10756,N_9548,N_2673);
xor U10757 (N_10757,N_6730,N_5950);
xnor U10758 (N_10758,N_570,N_5633);
and U10759 (N_10759,N_704,N_1950);
nand U10760 (N_10760,N_979,N_2131);
or U10761 (N_10761,N_2323,N_5284);
nor U10762 (N_10762,N_1799,N_8960);
and U10763 (N_10763,N_7393,N_9240);
nand U10764 (N_10764,N_3785,N_8563);
nor U10765 (N_10765,N_5833,N_5765);
xor U10766 (N_10766,N_9003,N_7980);
nand U10767 (N_10767,N_3543,N_6688);
xor U10768 (N_10768,N_3248,N_5256);
xor U10769 (N_10769,N_1244,N_5696);
or U10770 (N_10770,N_1868,N_5798);
and U10771 (N_10771,N_2287,N_9557);
nor U10772 (N_10772,N_8487,N_8702);
and U10773 (N_10773,N_1689,N_8733);
and U10774 (N_10774,N_8086,N_3079);
and U10775 (N_10775,N_8343,N_8283);
nand U10776 (N_10776,N_1603,N_7991);
nand U10777 (N_10777,N_3848,N_8799);
and U10778 (N_10778,N_7288,N_3092);
xnor U10779 (N_10779,N_7031,N_747);
and U10780 (N_10780,N_8260,N_5435);
and U10781 (N_10781,N_2588,N_4658);
and U10782 (N_10782,N_8737,N_57);
nand U10783 (N_10783,N_1723,N_5152);
and U10784 (N_10784,N_290,N_1595);
and U10785 (N_10785,N_6140,N_7629);
or U10786 (N_10786,N_6443,N_3517);
nor U10787 (N_10787,N_8249,N_9571);
xnor U10788 (N_10788,N_1703,N_6741);
xnor U10789 (N_10789,N_679,N_8748);
or U10790 (N_10790,N_9643,N_9831);
nand U10791 (N_10791,N_2305,N_2875);
and U10792 (N_10792,N_4002,N_8321);
nor U10793 (N_10793,N_1502,N_9963);
or U10794 (N_10794,N_4639,N_5211);
nor U10795 (N_10795,N_9071,N_6778);
and U10796 (N_10796,N_1467,N_6621);
xor U10797 (N_10797,N_8123,N_9255);
nor U10798 (N_10798,N_375,N_8230);
nor U10799 (N_10799,N_5657,N_270);
nand U10800 (N_10800,N_7465,N_5923);
nand U10801 (N_10801,N_4492,N_9704);
xnor U10802 (N_10802,N_8704,N_4931);
and U10803 (N_10803,N_6277,N_5180);
or U10804 (N_10804,N_7079,N_58);
or U10805 (N_10805,N_1740,N_3278);
nand U10806 (N_10806,N_1693,N_622);
nand U10807 (N_10807,N_3547,N_1163);
or U10808 (N_10808,N_7114,N_7179);
nor U10809 (N_10809,N_1567,N_567);
nand U10810 (N_10810,N_7117,N_7050);
and U10811 (N_10811,N_8064,N_6192);
and U10812 (N_10812,N_2744,N_6984);
xnor U10813 (N_10813,N_7389,N_5147);
and U10814 (N_10814,N_9285,N_2455);
nor U10815 (N_10815,N_2006,N_5040);
and U10816 (N_10816,N_9120,N_8610);
or U10817 (N_10817,N_9295,N_1157);
nor U10818 (N_10818,N_8506,N_4409);
or U10819 (N_10819,N_6997,N_2591);
and U10820 (N_10820,N_3665,N_8668);
nand U10821 (N_10821,N_9769,N_3924);
xor U10822 (N_10822,N_4355,N_5080);
and U10823 (N_10823,N_9324,N_7737);
and U10824 (N_10824,N_4691,N_9415);
nor U10825 (N_10825,N_4188,N_1016);
xnor U10826 (N_10826,N_9558,N_2791);
xor U10827 (N_10827,N_8821,N_5522);
nand U10828 (N_10828,N_6944,N_6398);
or U10829 (N_10829,N_9581,N_6161);
nor U10830 (N_10830,N_919,N_3809);
nor U10831 (N_10831,N_831,N_7783);
or U10832 (N_10832,N_1105,N_6832);
nand U10833 (N_10833,N_7607,N_7274);
nor U10834 (N_10834,N_3931,N_8);
nand U10835 (N_10835,N_1894,N_9691);
nor U10836 (N_10836,N_7586,N_1411);
nor U10837 (N_10837,N_1269,N_8795);
xor U10838 (N_10838,N_5802,N_4910);
nor U10839 (N_10839,N_9111,N_7048);
nor U10840 (N_10840,N_8029,N_5707);
nor U10841 (N_10841,N_3946,N_9775);
and U10842 (N_10842,N_5721,N_1987);
and U10843 (N_10843,N_1279,N_6666);
and U10844 (N_10844,N_7147,N_3449);
or U10845 (N_10845,N_8617,N_2345);
xor U10846 (N_10846,N_2052,N_8832);
xnor U10847 (N_10847,N_2048,N_746);
nand U10848 (N_10848,N_8177,N_1809);
and U10849 (N_10849,N_3869,N_7466);
or U10850 (N_10850,N_9002,N_6266);
or U10851 (N_10851,N_3957,N_3516);
and U10852 (N_10852,N_23,N_509);
or U10853 (N_10853,N_7624,N_4375);
and U10854 (N_10854,N_867,N_2163);
xor U10855 (N_10855,N_1726,N_9968);
or U10856 (N_10856,N_4403,N_2923);
xnor U10857 (N_10857,N_90,N_8772);
nand U10858 (N_10858,N_1190,N_8158);
or U10859 (N_10859,N_9799,N_7597);
and U10860 (N_10860,N_9115,N_7998);
nor U10861 (N_10861,N_271,N_6185);
and U10862 (N_10862,N_7224,N_381);
nand U10863 (N_10863,N_45,N_7536);
or U10864 (N_10864,N_3419,N_6594);
xor U10865 (N_10865,N_225,N_3800);
nor U10866 (N_10866,N_3317,N_9470);
nand U10867 (N_10867,N_1312,N_7647);
or U10868 (N_10868,N_8363,N_9999);
nand U10869 (N_10869,N_1220,N_6643);
nor U10870 (N_10870,N_2509,N_5859);
or U10871 (N_10871,N_7503,N_6763);
and U10872 (N_10872,N_3731,N_7927);
nand U10873 (N_10873,N_9883,N_7136);
nor U10874 (N_10874,N_1545,N_9740);
xor U10875 (N_10875,N_4265,N_2051);
and U10876 (N_10876,N_9308,N_9136);
and U10877 (N_10877,N_2594,N_7810);
and U10878 (N_10878,N_7865,N_4579);
or U10879 (N_10879,N_6574,N_8706);
nand U10880 (N_10880,N_4747,N_1054);
nand U10881 (N_10881,N_5130,N_6907);
nand U10882 (N_10882,N_9270,N_404);
or U10883 (N_10883,N_5101,N_2884);
and U10884 (N_10884,N_903,N_3279);
nor U10885 (N_10885,N_6431,N_9384);
or U10886 (N_10886,N_8599,N_7643);
nand U10887 (N_10887,N_4923,N_5561);
and U10888 (N_10888,N_3696,N_6359);
xor U10889 (N_10889,N_573,N_7623);
nand U10890 (N_10890,N_3981,N_9664);
or U10891 (N_10891,N_8147,N_8200);
and U10892 (N_10892,N_2993,N_6313);
nor U10893 (N_10893,N_8285,N_3896);
and U10894 (N_10894,N_9430,N_9090);
and U10895 (N_10895,N_6879,N_5542);
and U10896 (N_10896,N_2002,N_1131);
or U10897 (N_10897,N_2015,N_8039);
xor U10898 (N_10898,N_5052,N_6045);
nand U10899 (N_10899,N_6644,N_5616);
nor U10900 (N_10900,N_7369,N_3996);
or U10901 (N_10901,N_7996,N_8463);
or U10902 (N_10902,N_5884,N_1507);
nor U10903 (N_10903,N_9290,N_504);
or U10904 (N_10904,N_2112,N_976);
and U10905 (N_10905,N_6475,N_1322);
nor U10906 (N_10906,N_9849,N_3511);
and U10907 (N_10907,N_8770,N_8218);
or U10908 (N_10908,N_5640,N_3070);
xnor U10909 (N_10909,N_1170,N_1303);
or U10910 (N_10910,N_475,N_8587);
nor U10911 (N_10911,N_5230,N_1781);
nand U10912 (N_10912,N_8634,N_2686);
xor U10913 (N_10913,N_4927,N_2642);
xor U10914 (N_10914,N_5372,N_2995);
xnor U10915 (N_10915,N_8251,N_459);
or U10916 (N_10916,N_340,N_9076);
nand U10917 (N_10917,N_3674,N_5562);
and U10918 (N_10918,N_8974,N_128);
nand U10919 (N_10919,N_5829,N_888);
and U10920 (N_10920,N_3183,N_1460);
or U10921 (N_10921,N_3564,N_1344);
nor U10922 (N_10922,N_8675,N_6863);
and U10923 (N_10923,N_4092,N_8007);
and U10924 (N_10924,N_2489,N_7997);
xnor U10925 (N_10925,N_3867,N_4953);
or U10926 (N_10926,N_3481,N_187);
nor U10927 (N_10927,N_1845,N_542);
xor U10928 (N_10928,N_8350,N_2082);
nor U10929 (N_10929,N_1042,N_7558);
or U10930 (N_10930,N_3093,N_4985);
and U10931 (N_10931,N_7784,N_2902);
xnor U10932 (N_10932,N_4506,N_4737);
nor U10933 (N_10933,N_6771,N_8872);
and U10934 (N_10934,N_8243,N_9942);
or U10935 (N_10935,N_2240,N_8155);
xor U10936 (N_10936,N_5373,N_2179);
xor U10937 (N_10937,N_9863,N_7336);
nor U10938 (N_10938,N_1468,N_4158);
and U10939 (N_10939,N_3860,N_3604);
nor U10940 (N_10940,N_6927,N_1067);
nand U10941 (N_10941,N_6155,N_2937);
nand U10942 (N_10942,N_336,N_9665);
or U10943 (N_10943,N_2926,N_5499);
and U10944 (N_10944,N_446,N_7480);
nor U10945 (N_10945,N_6472,N_4342);
and U10946 (N_10946,N_8830,N_4857);
and U10947 (N_10947,N_9798,N_4057);
nor U10948 (N_10948,N_1218,N_3057);
or U10949 (N_10949,N_6612,N_2722);
nand U10950 (N_10950,N_132,N_6464);
xnor U10951 (N_10951,N_3068,N_8878);
xnor U10952 (N_10952,N_926,N_9811);
xor U10953 (N_10953,N_6841,N_3900);
and U10954 (N_10954,N_1106,N_5382);
nor U10955 (N_10955,N_102,N_274);
xnor U10956 (N_10956,N_6597,N_427);
and U10957 (N_10957,N_5283,N_7691);
xor U10958 (N_10958,N_4582,N_7385);
or U10959 (N_10959,N_412,N_8149);
nand U10960 (N_10960,N_8431,N_5742);
nand U10961 (N_10961,N_6536,N_3923);
or U10962 (N_10962,N_5970,N_7826);
or U10963 (N_10963,N_2258,N_1186);
xnor U10964 (N_10964,N_2890,N_2402);
nor U10965 (N_10965,N_931,N_8151);
xor U10966 (N_10966,N_3916,N_6798);
xnor U10967 (N_10967,N_9007,N_7091);
nor U10968 (N_10968,N_6521,N_7542);
and U10969 (N_10969,N_5419,N_4824);
and U10970 (N_10970,N_7448,N_1162);
nor U10971 (N_10971,N_7658,N_379);
nand U10972 (N_10972,N_83,N_1213);
nor U10973 (N_10973,N_7891,N_3532);
nand U10974 (N_10974,N_9265,N_8464);
xor U10975 (N_10975,N_3757,N_2037);
nand U10976 (N_10976,N_9872,N_2760);
and U10977 (N_10977,N_1583,N_3351);
nand U10978 (N_10978,N_3508,N_186);
nand U10979 (N_10979,N_1490,N_2774);
nor U10980 (N_10980,N_7273,N_6755);
nor U10981 (N_10981,N_1046,N_2909);
or U10982 (N_10982,N_2231,N_8571);
nand U10983 (N_10983,N_1286,N_7380);
or U10984 (N_10984,N_7150,N_2238);
nor U10985 (N_10985,N_8977,N_9796);
nor U10986 (N_10986,N_6080,N_157);
or U10987 (N_10987,N_3425,N_7676);
nor U10988 (N_10988,N_6722,N_2418);
or U10989 (N_10989,N_5396,N_7850);
nand U10990 (N_10990,N_4760,N_2807);
or U10991 (N_10991,N_7580,N_3850);
nor U10992 (N_10992,N_93,N_2941);
nand U10993 (N_10993,N_1337,N_151);
nand U10994 (N_10994,N_4160,N_9504);
and U10995 (N_10995,N_726,N_2784);
or U10996 (N_10996,N_2445,N_8548);
xnor U10997 (N_10997,N_7541,N_8197);
and U10998 (N_10998,N_315,N_1506);
nor U10999 (N_10999,N_6107,N_2420);
nand U11000 (N_11000,N_6485,N_1546);
or U11001 (N_11001,N_1548,N_94);
nor U11002 (N_11002,N_9048,N_4507);
xor U11003 (N_11003,N_4071,N_496);
nor U11004 (N_11004,N_7764,N_1333);
xor U11005 (N_11005,N_7128,N_871);
xnor U11006 (N_11006,N_3887,N_5609);
or U11007 (N_11007,N_3101,N_3537);
nand U11008 (N_11008,N_4404,N_7093);
and U11009 (N_11009,N_2530,N_4768);
nor U11010 (N_11010,N_9440,N_3987);
or U11011 (N_11011,N_8855,N_7039);
and U11012 (N_11012,N_1025,N_9342);
nand U11013 (N_11013,N_5617,N_1482);
and U11014 (N_11014,N_975,N_6295);
nand U11015 (N_11015,N_965,N_3838);
nor U11016 (N_11016,N_3587,N_9);
nand U11017 (N_11017,N_1427,N_610);
xnor U11018 (N_11018,N_9940,N_34);
and U11019 (N_11019,N_3591,N_8719);
xnor U11020 (N_11020,N_8397,N_3043);
xnor U11021 (N_11021,N_7759,N_232);
nand U11022 (N_11022,N_1289,N_44);
or U11023 (N_11023,N_2197,N_9770);
nor U11024 (N_11024,N_8278,N_7924);
nand U11025 (N_11025,N_6440,N_3877);
or U11026 (N_11026,N_302,N_8509);
nand U11027 (N_11027,N_3196,N_9977);
and U11028 (N_11028,N_7556,N_5608);
xnor U11029 (N_11029,N_5174,N_5602);
nor U11030 (N_11030,N_8577,N_1980);
and U11031 (N_11031,N_3717,N_447);
and U11032 (N_11032,N_1702,N_9142);
xor U11033 (N_11033,N_6934,N_3740);
or U11034 (N_11034,N_2281,N_9947);
or U11035 (N_11035,N_7653,N_337);
xor U11036 (N_11036,N_6112,N_5088);
xor U11037 (N_11037,N_3287,N_9781);
nor U11038 (N_11038,N_6132,N_3975);
and U11039 (N_11039,N_6287,N_7060);
and U11040 (N_11040,N_1626,N_476);
nand U11041 (N_11041,N_650,N_1092);
nor U11042 (N_11042,N_9656,N_378);
and U11043 (N_11043,N_9802,N_6097);
xor U11044 (N_11044,N_2135,N_406);
nor U11045 (N_11045,N_1734,N_3962);
xor U11046 (N_11046,N_9776,N_7857);
nand U11047 (N_11047,N_953,N_9500);
nor U11048 (N_11048,N_8468,N_9601);
nand U11049 (N_11049,N_5259,N_2971);
nand U11050 (N_11050,N_5858,N_8881);
and U11051 (N_11051,N_9985,N_1715);
nor U11052 (N_11052,N_2329,N_534);
nor U11053 (N_11053,N_2035,N_4089);
nor U11054 (N_11054,N_1510,N_5392);
nand U11055 (N_11055,N_2456,N_2604);
or U11056 (N_11056,N_9334,N_3206);
xor U11057 (N_11057,N_3687,N_6069);
xor U11058 (N_11058,N_9381,N_5121);
nor U11059 (N_11059,N_7825,N_6336);
nor U11060 (N_11060,N_3148,N_7129);
or U11061 (N_11061,N_8782,N_8791);
and U11062 (N_11062,N_4884,N_3879);
nand U11063 (N_11063,N_470,N_2674);
xnor U11064 (N_11064,N_7264,N_2718);
or U11065 (N_11065,N_8992,N_5922);
nor U11066 (N_11066,N_1158,N_8640);
or U11067 (N_11067,N_8352,N_1663);
and U11068 (N_11068,N_3105,N_5769);
or U11069 (N_11069,N_152,N_9033);
and U11070 (N_11070,N_9527,N_2089);
nand U11071 (N_11071,N_5860,N_3307);
or U11072 (N_11072,N_5669,N_6561);
and U11073 (N_11073,N_7628,N_4200);
xor U11074 (N_11074,N_2586,N_1779);
and U11075 (N_11075,N_4173,N_6325);
nor U11076 (N_11076,N_5469,N_4574);
and U11077 (N_11077,N_9600,N_6260);
nand U11078 (N_11078,N_8815,N_948);
xnor U11079 (N_11079,N_5887,N_5999);
nand U11080 (N_11080,N_2767,N_8450);
and U11081 (N_11081,N_2032,N_9450);
and U11082 (N_11082,N_6349,N_4081);
nand U11083 (N_11083,N_3965,N_6004);
nor U11084 (N_11084,N_8317,N_7262);
and U11085 (N_11085,N_5074,N_9020);
or U11086 (N_11086,N_1859,N_7951);
and U11087 (N_11087,N_2741,N_4548);
xor U11088 (N_11088,N_1187,N_9127);
nor U11089 (N_11089,N_9929,N_8693);
nand U11090 (N_11090,N_7194,N_7766);
xnor U11091 (N_11091,N_3144,N_5899);
and U11092 (N_11092,N_4533,N_2446);
or U11093 (N_11093,N_2629,N_3926);
and U11094 (N_11094,N_6092,N_9585);
or U11095 (N_11095,N_1435,N_925);
nand U11096 (N_11096,N_9989,N_5717);
nor U11097 (N_11097,N_5064,N_5458);
or U11098 (N_11098,N_5727,N_4099);
nor U11099 (N_11099,N_4423,N_1628);
nand U11100 (N_11100,N_3752,N_8592);
or U11101 (N_11101,N_3807,N_2868);
nand U11102 (N_11102,N_4372,N_6220);
and U11103 (N_11103,N_6620,N_634);
or U11104 (N_11104,N_3913,N_6607);
xor U11105 (N_11105,N_2357,N_3863);
or U11106 (N_11106,N_7361,N_5460);
and U11107 (N_11107,N_5879,N_5087);
nand U11108 (N_11108,N_6786,N_4755);
nor U11109 (N_11109,N_9812,N_2356);
or U11110 (N_11110,N_9521,N_9520);
xnor U11111 (N_11111,N_1211,N_3935);
and U11112 (N_11112,N_2969,N_3230);
and U11113 (N_11113,N_5399,N_7324);
and U11114 (N_11114,N_1448,N_5847);
xor U11115 (N_11115,N_4171,N_7550);
and U11116 (N_11116,N_7801,N_708);
or U11117 (N_11117,N_4659,N_1563);
nand U11118 (N_11118,N_2361,N_5988);
and U11119 (N_11119,N_4719,N_420);
nor U11120 (N_11120,N_1242,N_9875);
nor U11121 (N_11121,N_5713,N_2115);
or U11122 (N_11122,N_2394,N_5450);
and U11123 (N_11123,N_6226,N_2954);
nor U11124 (N_11124,N_9170,N_3797);
xnor U11125 (N_11125,N_7061,N_858);
nor U11126 (N_11126,N_4918,N_2539);
nand U11127 (N_11127,N_722,N_4990);
and U11128 (N_11128,N_2093,N_9261);
nor U11129 (N_11129,N_2742,N_2776);
or U11130 (N_11130,N_1793,N_190);
and U11131 (N_11131,N_6514,N_7335);
and U11132 (N_11132,N_1806,N_1125);
or U11133 (N_11133,N_6476,N_4458);
nor U11134 (N_11134,N_1718,N_7837);
or U11135 (N_11135,N_4514,N_519);
nand U11136 (N_11136,N_453,N_5081);
nor U11137 (N_11137,N_6596,N_376);
nand U11138 (N_11138,N_8484,N_6219);
nand U11139 (N_11139,N_6539,N_2175);
xor U11140 (N_11140,N_9447,N_7579);
and U11141 (N_11141,N_3509,N_3084);
nor U11142 (N_11142,N_1638,N_349);
or U11143 (N_11143,N_9851,N_4340);
or U11144 (N_11144,N_4019,N_2924);
or U11145 (N_11145,N_8383,N_8228);
nand U11146 (N_11146,N_7788,N_364);
nor U11147 (N_11147,N_4614,N_6966);
nor U11148 (N_11148,N_6792,N_1606);
xor U11149 (N_11149,N_3977,N_2788);
nand U11150 (N_11150,N_3052,N_4952);
xor U11151 (N_11151,N_2508,N_7969);
nor U11152 (N_11152,N_6471,N_4631);
or U11153 (N_11153,N_9736,N_8398);
nand U11154 (N_11154,N_7275,N_291);
or U11155 (N_11155,N_4212,N_50);
and U11156 (N_11156,N_5415,N_3496);
xor U11157 (N_11157,N_3232,N_20);
nand U11158 (N_11158,N_7546,N_756);
xnor U11159 (N_11159,N_869,N_351);
xnor U11160 (N_11160,N_8478,N_9927);
or U11161 (N_11161,N_3188,N_6154);
xor U11162 (N_11162,N_2911,N_5129);
nor U11163 (N_11163,N_922,N_8174);
or U11164 (N_11164,N_1004,N_1785);
or U11165 (N_11165,N_9692,N_335);
nand U11166 (N_11166,N_6710,N_1231);
or U11167 (N_11167,N_2388,N_5406);
xor U11168 (N_11168,N_2835,N_4459);
xor U11169 (N_11169,N_7925,N_1486);
nor U11170 (N_11170,N_587,N_181);
nor U11171 (N_11171,N_5764,N_1357);
or U11172 (N_11172,N_9427,N_6576);
nor U11173 (N_11173,N_9829,N_5299);
and U11174 (N_11174,N_1616,N_8042);
and U11175 (N_11175,N_2625,N_9256);
nor U11176 (N_11176,N_6470,N_3459);
nor U11177 (N_11177,N_1109,N_318);
and U11178 (N_11178,N_1059,N_9216);
nand U11179 (N_11179,N_7853,N_8896);
xor U11180 (N_11180,N_1249,N_4628);
and U11181 (N_11181,N_8422,N_2069);
nand U11182 (N_11182,N_1075,N_6211);
or U11183 (N_11183,N_1201,N_7545);
nor U11184 (N_11184,N_7021,N_5035);
nor U11185 (N_11185,N_5595,N_935);
nor U11186 (N_11186,N_1964,N_2302);
and U11187 (N_11187,N_3492,N_6690);
xnor U11188 (N_11188,N_1605,N_4782);
xnor U11189 (N_11189,N_3775,N_2423);
nor U11190 (N_11190,N_4030,N_8441);
nor U11191 (N_11191,N_7082,N_9939);
nand U11192 (N_11192,N_5302,N_4255);
or U11193 (N_11193,N_5082,N_2810);
and U11194 (N_11194,N_2904,N_4668);
or U11195 (N_11195,N_2430,N_874);
and U11196 (N_11196,N_7779,N_6497);
and U11197 (N_11197,N_6756,N_3028);
nor U11198 (N_11198,N_4876,N_5515);
nand U11199 (N_11199,N_3149,N_2493);
xnor U11200 (N_11200,N_7460,N_2831);
nand U11201 (N_11201,N_4638,N_7729);
and U11202 (N_11202,N_140,N_3320);
xor U11203 (N_11203,N_6021,N_3704);
xor U11204 (N_11204,N_5324,N_942);
nor U11205 (N_11205,N_3593,N_1045);
or U11206 (N_11206,N_1070,N_5220);
or U11207 (N_11207,N_3895,N_8417);
or U11208 (N_11208,N_4337,N_9056);
xor U11209 (N_11209,N_1679,N_2511);
xnor U11210 (N_11210,N_6768,N_4733);
and U11211 (N_11211,N_6062,N_2252);
and U11212 (N_11212,N_9632,N_7966);
xnor U11213 (N_11213,N_7775,N_8652);
and U11214 (N_11214,N_1191,N_163);
or U11215 (N_11215,N_3737,N_4959);
and U11216 (N_11216,N_4793,N_1048);
xnor U11217 (N_11217,N_663,N_9637);
or U11218 (N_11218,N_5333,N_4848);
nor U11219 (N_11219,N_8438,N_1753);
or U11220 (N_11220,N_3121,N_7512);
and U11221 (N_11221,N_9956,N_2454);
and U11222 (N_11222,N_6813,N_3692);
and U11223 (N_11223,N_3166,N_4485);
xnor U11224 (N_11224,N_5930,N_2522);
nor U11225 (N_11225,N_312,N_4900);
nor U11226 (N_11226,N_5967,N_9178);
xnor U11227 (N_11227,N_1040,N_5537);
nand U11228 (N_11228,N_3739,N_9496);
nand U11229 (N_11229,N_1541,N_2081);
and U11230 (N_11230,N_6244,N_7250);
xor U11231 (N_11231,N_5583,N_9506);
and U11232 (N_11232,N_5292,N_9805);
and U11233 (N_11233,N_4661,N_9105);
or U11234 (N_11234,N_9995,N_2915);
nand U11235 (N_11235,N_1933,N_8256);
or U11236 (N_11236,N_7549,N_1790);
nor U11237 (N_11237,N_5981,N_2428);
nand U11238 (N_11238,N_8143,N_7218);
and U11239 (N_11239,N_2451,N_4453);
nand U11240 (N_11240,N_1442,N_8226);
and U11241 (N_11241,N_879,N_450);
xnor U11242 (N_11242,N_5501,N_1665);
nand U11243 (N_11243,N_3734,N_4418);
nor U11244 (N_11244,N_7183,N_6538);
xor U11245 (N_11245,N_8367,N_9110);
nand U11246 (N_11246,N_7261,N_1948);
nor U11247 (N_11247,N_9973,N_6992);
and U11248 (N_11248,N_198,N_9028);
nand U11249 (N_11249,N_2070,N_1573);
nor U11250 (N_11250,N_1527,N_8154);
nand U11251 (N_11251,N_9325,N_8823);
nor U11252 (N_11252,N_353,N_6857);
or U11253 (N_11253,N_1026,N_2544);
xor U11254 (N_11254,N_1989,N_5546);
nor U11255 (N_11255,N_681,N_6961);
nand U11256 (N_11256,N_7622,N_3583);
nor U11257 (N_11257,N_4946,N_6605);
or U11258 (N_11258,N_895,N_5496);
or U11259 (N_11259,N_6296,N_317);
xor U11260 (N_11260,N_6969,N_1839);
nand U11261 (N_11261,N_8261,N_4911);
xnor U11262 (N_11262,N_5331,N_7246);
nand U11263 (N_11263,N_3915,N_492);
or U11264 (N_11264,N_3615,N_8138);
and U11265 (N_11265,N_4488,N_8079);
nand U11266 (N_11266,N_2425,N_2662);
and U11267 (N_11267,N_9439,N_5512);
nand U11268 (N_11268,N_9457,N_2392);
and U11269 (N_11269,N_2989,N_5468);
nor U11270 (N_11270,N_9766,N_7679);
or U11271 (N_11271,N_3173,N_4834);
nor U11272 (N_11272,N_3661,N_8961);
nand U11273 (N_11273,N_1953,N_9330);
nor U11274 (N_11274,N_3289,N_6806);
and U11275 (N_11275,N_2990,N_6428);
nor U11276 (N_11276,N_6204,N_4813);
nor U11277 (N_11277,N_9619,N_5589);
and U11278 (N_11278,N_5383,N_9390);
or U11279 (N_11279,N_637,N_4821);
nor U11280 (N_11280,N_205,N_5683);
xor U11281 (N_11281,N_7568,N_8766);
nand U11282 (N_11282,N_4100,N_4144);
nor U11283 (N_11283,N_3619,N_1226);
xor U11284 (N_11284,N_6559,N_3892);
xor U11285 (N_11285,N_3743,N_6917);
xor U11286 (N_11286,N_9057,N_7286);
and U11287 (N_11287,N_2860,N_5951);
and U11288 (N_11288,N_4981,N_4376);
xnor U11289 (N_11289,N_5350,N_4486);
nor U11290 (N_11290,N_546,N_7010);
nand U11291 (N_11291,N_6991,N_8391);
nor U11292 (N_11292,N_2910,N_4686);
nand U11293 (N_11293,N_9857,N_5857);
or U11294 (N_11294,N_6165,N_7726);
or U11295 (N_11295,N_3598,N_368);
xnor U11296 (N_11296,N_1787,N_8901);
and U11297 (N_11297,N_1643,N_5295);
nor U11298 (N_11298,N_9383,N_3291);
and U11299 (N_11299,N_5440,N_9335);
or U11300 (N_11300,N_6289,N_3139);
nand U11301 (N_11301,N_5070,N_8535);
nor U11302 (N_11302,N_5743,N_8236);
and U11303 (N_11303,N_4647,N_5327);
nor U11304 (N_11304,N_9021,N_8802);
nand U11305 (N_11305,N_6649,N_5293);
nand U11306 (N_11306,N_7327,N_6085);
and U11307 (N_11307,N_3688,N_2272);
or U11308 (N_11308,N_8790,N_1864);
nand U11309 (N_11309,N_730,N_9297);
and U11310 (N_11310,N_9878,N_2537);
and U11311 (N_11311,N_429,N_7192);
nor U11312 (N_11312,N_7948,N_5217);
nand U11313 (N_11313,N_3310,N_7402);
xor U11314 (N_11314,N_402,N_9681);
xor U11315 (N_11315,N_4511,N_4420);
nand U11316 (N_11316,N_7862,N_640);
nor U11317 (N_11317,N_1674,N_3796);
or U11318 (N_11318,N_9890,N_8388);
nand U11319 (N_11319,N_7318,N_6376);
nor U11320 (N_11320,N_7518,N_5198);
and U11321 (N_11321,N_7879,N_5730);
nor U11322 (N_11322,N_6855,N_3469);
xor U11323 (N_11323,N_5436,N_9727);
xor U11324 (N_11324,N_6783,N_5869);
nor U11325 (N_11325,N_9171,N_2246);
nand U11326 (N_11326,N_5738,N_7767);
nand U11327 (N_11327,N_3662,N_6772);
xnor U11328 (N_11328,N_7135,N_8752);
or U11329 (N_11329,N_2276,N_8319);
xor U11330 (N_11330,N_1505,N_2265);
nor U11331 (N_11331,N_493,N_6836);
nand U11332 (N_11332,N_4140,N_2441);
xor U11333 (N_11333,N_6176,N_3766);
nand U11334 (N_11334,N_9488,N_4697);
or U11335 (N_11335,N_3240,N_2800);
xnor U11336 (N_11336,N_2660,N_1539);
nand U11337 (N_11337,N_1480,N_3157);
nand U11338 (N_11338,N_3170,N_6484);
and U11339 (N_11339,N_7401,N_628);
xnor U11340 (N_11340,N_8726,N_8237);
or U11341 (N_11341,N_7890,N_1394);
nand U11342 (N_11342,N_8579,N_8905);
nor U11343 (N_11343,N_1134,N_4808);
nand U11344 (N_11344,N_5574,N_1102);
xor U11345 (N_11345,N_9331,N_5386);
and U11346 (N_11346,N_911,N_8078);
xor U11347 (N_11347,N_4787,N_8683);
and U11348 (N_11348,N_8531,N_5263);
nor U11349 (N_11349,N_7446,N_7146);
xnor U11350 (N_11350,N_6190,N_1947);
and U11351 (N_11351,N_4526,N_8594);
nand U11352 (N_11352,N_2483,N_8162);
or U11353 (N_11353,N_877,N_6877);
nor U11354 (N_11354,N_6852,N_3715);
or U11355 (N_11355,N_3429,N_8294);
nor U11356 (N_11356,N_9184,N_6316);
nand U11357 (N_11357,N_4779,N_7112);
and U11358 (N_11358,N_5762,N_1543);
nand U11359 (N_11359,N_6060,N_2679);
and U11360 (N_11360,N_6762,N_6039);
and U11361 (N_11361,N_9143,N_5913);
nand U11362 (N_11362,N_9094,N_8499);
xor U11363 (N_11363,N_1391,N_9283);
or U11364 (N_11364,N_1265,N_9998);
and U11365 (N_11365,N_6144,N_3520);
nor U11366 (N_11366,N_8329,N_6904);
nand U11367 (N_11367,N_7461,N_1985);
and U11368 (N_11368,N_1918,N_260);
or U11369 (N_11369,N_4708,N_11);
and U11370 (N_11370,N_2080,N_9418);
or U11371 (N_11371,N_1457,N_5498);
xnor U11372 (N_11372,N_2,N_7675);
or U11373 (N_11373,N_1612,N_6168);
or U11374 (N_11374,N_188,N_3738);
nand U11375 (N_11375,N_7960,N_3119);
and U11376 (N_11376,N_2043,N_822);
nand U11377 (N_11377,N_6233,N_8045);
xnor U11378 (N_11378,N_8868,N_3476);
nand U11379 (N_11379,N_9923,N_4359);
or U11380 (N_11380,N_9597,N_2880);
or U11381 (N_11381,N_9921,N_3727);
xor U11382 (N_11382,N_4462,N_7270);
nand U11383 (N_11383,N_438,N_3130);
or U11384 (N_11384,N_8596,N_7175);
nand U11385 (N_11385,N_2817,N_8713);
or U11386 (N_11386,N_149,N_6267);
or U11387 (N_11387,N_3632,N_9505);
xor U11388 (N_11388,N_1395,N_5412);
nor U11389 (N_11389,N_3950,N_6675);
or U11390 (N_11390,N_9487,N_4260);
nand U11391 (N_11391,N_8449,N_8871);
and U11392 (N_11392,N_9154,N_1861);
nor U11393 (N_11393,N_3858,N_8663);
nor U11394 (N_11394,N_9551,N_7452);
xnor U11395 (N_11395,N_469,N_6162);
or U11396 (N_11396,N_8847,N_1463);
xnor U11397 (N_11397,N_8760,N_6663);
and U11398 (N_11398,N_8764,N_7301);
or U11399 (N_11399,N_9175,N_5505);
or U11400 (N_11400,N_3830,N_3269);
and U11401 (N_11401,N_1013,N_1126);
xnor U11402 (N_11402,N_6767,N_3880);
and U11403 (N_11403,N_6960,N_8180);
xor U11404 (N_11404,N_9723,N_2792);
xnor U11405 (N_11405,N_9038,N_6383);
nor U11406 (N_11406,N_2208,N_6231);
and U11407 (N_11407,N_5607,N_7411);
nor U11408 (N_11408,N_8322,N_7231);
or U11409 (N_11409,N_3237,N_6130);
nand U11410 (N_11410,N_1041,N_6592);
nor U11411 (N_11411,N_1596,N_1000);
or U11412 (N_11412,N_5579,N_207);
or U11413 (N_11413,N_4543,N_9173);
and U11414 (N_11414,N_363,N_9957);
or U11415 (N_11415,N_6447,N_9981);
or U11416 (N_11416,N_8969,N_4210);
xor U11417 (N_11417,N_8876,N_2925);
xor U11418 (N_11418,N_9967,N_8958);
xor U11419 (N_11419,N_5500,N_5700);
nand U11420 (N_11420,N_7886,N_3329);
nand U11421 (N_11421,N_9385,N_361);
and U11422 (N_11422,N_9360,N_1080);
nor U11423 (N_11423,N_2895,N_1325);
nor U11424 (N_11424,N_4201,N_1885);
nor U11425 (N_11425,N_6234,N_3983);
xnor U11426 (N_11426,N_1012,N_9969);
and U11427 (N_11427,N_4426,N_2952);
or U11428 (N_11428,N_8248,N_95);
and U11429 (N_11429,N_9706,N_9928);
or U11430 (N_11430,N_7994,N_3129);
nor U11431 (N_11431,N_2506,N_9053);
nand U11432 (N_11432,N_7713,N_2172);
nor U11433 (N_11433,N_618,N_2961);
nand U11434 (N_11434,N_605,N_2484);
nand U11435 (N_11435,N_536,N_2421);
and U11436 (N_11436,N_2654,N_5755);
xnor U11437 (N_11437,N_660,N_4455);
and U11438 (N_11438,N_4361,N_984);
and U11439 (N_11439,N_7702,N_2617);
or U11440 (N_11440,N_5073,N_37);
nand U11441 (N_11441,N_7696,N_1652);
or U11442 (N_11442,N_6900,N_6363);
nand U11443 (N_11443,N_3417,N_9765);
nand U11444 (N_11444,N_2190,N_4117);
nand U11445 (N_11445,N_9702,N_9389);
nor U11446 (N_11446,N_5686,N_244);
or U11447 (N_11447,N_6465,N_9362);
or U11448 (N_11448,N_4575,N_5421);
nand U11449 (N_11449,N_7625,N_1088);
or U11450 (N_11450,N_3364,N_9758);
xnor U11451 (N_11451,N_2366,N_7583);
nand U11452 (N_11452,N_7481,N_1021);
and U11453 (N_11453,N_204,N_8826);
and U11454 (N_11454,N_2619,N_821);
or U11455 (N_11455,N_4285,N_4399);
or U11456 (N_11456,N_4076,N_6752);
nor U11457 (N_11457,N_4999,N_5653);
xnor U11458 (N_11458,N_4011,N_3503);
and U11459 (N_11459,N_7388,N_9728);
xnor U11460 (N_11460,N_7517,N_6578);
and U11461 (N_11461,N_1176,N_2413);
xnor U11462 (N_11462,N_3990,N_1421);
nor U11463 (N_11463,N_5104,N_1035);
or U11464 (N_11464,N_1891,N_4177);
nor U11465 (N_11465,N_1951,N_1334);
nor U11466 (N_11466,N_6509,N_1373);
xor U11467 (N_11467,N_295,N_6588);
nand U11468 (N_11468,N_2137,N_5056);
nand U11469 (N_11469,N_4012,N_2403);
or U11470 (N_11470,N_1214,N_621);
xor U11471 (N_11471,N_3639,N_4693);
xnor U11472 (N_11472,N_6947,N_2250);
and U11473 (N_11473,N_1637,N_2754);
nand U11474 (N_11474,N_8875,N_8360);
nand U11475 (N_11475,N_1281,N_110);
and U11476 (N_11476,N_1574,N_4436);
nand U11477 (N_11477,N_9446,N_4456);
and U11478 (N_11478,N_8127,N_4244);
nor U11479 (N_11479,N_774,N_4969);
xnor U11480 (N_11480,N_1923,N_6886);
nand U11481 (N_11481,N_4077,N_2072);
nand U11482 (N_11482,N_5148,N_696);
nand U11483 (N_11483,N_3940,N_2450);
and U11484 (N_11484,N_5751,N_4560);
or U11485 (N_11485,N_6916,N_4653);
and U11486 (N_11486,N_2275,N_9135);
and U11487 (N_11487,N_8307,N_1353);
nand U11488 (N_11488,N_1469,N_9595);
nor U11489 (N_11489,N_7819,N_4242);
nor U11490 (N_11490,N_4281,N_775);
or U11491 (N_11491,N_3891,N_5659);
or U11492 (N_11492,N_5272,N_2869);
and U11493 (N_11493,N_8415,N_2074);
nand U11494 (N_11494,N_5497,N_2852);
nand U11495 (N_11495,N_9673,N_3460);
xnor U11496 (N_11496,N_5577,N_3600);
xor U11497 (N_11497,N_5517,N_6463);
xnor U11498 (N_11498,N_9029,N_8859);
or U11499 (N_11499,N_4181,N_6726);
nand U11500 (N_11500,N_4726,N_3456);
nor U11501 (N_11501,N_136,N_7589);
nand U11502 (N_11502,N_445,N_2524);
and U11503 (N_11503,N_2350,N_7257);
or U11504 (N_11504,N_9499,N_6253);
xor U11505 (N_11505,N_3590,N_5948);
or U11506 (N_11506,N_2759,N_8074);
and U11507 (N_11507,N_5452,N_6392);
nand U11508 (N_11508,N_5199,N_3613);
or U11509 (N_11509,N_6423,N_524);
xnor U11510 (N_11510,N_2071,N_2397);
nor U11511 (N_11511,N_9044,N_1672);
or U11512 (N_11512,N_2194,N_9181);
and U11513 (N_11513,N_1501,N_2097);
nor U11514 (N_11514,N_6749,N_8315);
and U11515 (N_11515,N_4541,N_8040);
nand U11516 (N_11516,N_3286,N_7332);
and U11517 (N_11517,N_6541,N_5008);
or U11518 (N_11518,N_6298,N_4262);
or U11519 (N_11519,N_2216,N_4770);
and U11520 (N_11520,N_7880,N_4970);
nor U11521 (N_11521,N_4394,N_1805);
nor U11522 (N_11522,N_8017,N_8679);
nand U11523 (N_11523,N_8944,N_5235);
xor U11524 (N_11524,N_2424,N_6054);
and U11525 (N_11525,N_4792,N_6245);
or U11526 (N_11526,N_2457,N_9149);
xnor U11527 (N_11527,N_5407,N_2950);
nor U11528 (N_11528,N_9576,N_2865);
nor U11529 (N_11529,N_9559,N_683);
xor U11530 (N_11530,N_3282,N_1139);
xor U11531 (N_11531,N_5390,N_7985);
nor U11532 (N_11532,N_3095,N_5808);
or U11533 (N_11533,N_8691,N_5413);
xor U11534 (N_11534,N_8184,N_3654);
nor U11535 (N_11535,N_1477,N_6922);
nor U11536 (N_11536,N_2932,N_5158);
and U11537 (N_11537,N_845,N_360);
and U11538 (N_11538,N_9049,N_9202);
or U11539 (N_11539,N_1720,N_9264);
and U11540 (N_11540,N_8407,N_6525);
and U11541 (N_11541,N_651,N_5556);
or U11542 (N_11542,N_8076,N_1483);
nor U11543 (N_11543,N_8493,N_5289);
nor U11544 (N_11544,N_7923,N_2437);
nand U11545 (N_11545,N_362,N_6043);
or U11546 (N_11546,N_2670,N_4304);
nor U11547 (N_11547,N_1870,N_4701);
or U11548 (N_11548,N_8130,N_1668);
or U11549 (N_11549,N_9337,N_126);
or U11550 (N_11550,N_3605,N_5718);
nand U11551 (N_11551,N_4236,N_2558);
xnor U11552 (N_11552,N_589,N_4935);
xnor U11553 (N_11553,N_9943,N_3929);
nand U11554 (N_11554,N_3433,N_4622);
xor U11555 (N_11555,N_6729,N_8777);
nand U11556 (N_11556,N_5134,N_2157);
xnor U11557 (N_11557,N_8002,N_6548);
xnor U11558 (N_11558,N_8508,N_3767);
nand U11559 (N_11559,N_4272,N_6028);
and U11560 (N_11560,N_7026,N_497);
and U11561 (N_11561,N_5904,N_4934);
nor U11562 (N_11562,N_5897,N_3539);
and U11563 (N_11563,N_9344,N_7451);
xnor U11564 (N_11564,N_9259,N_1995);
nand U11565 (N_11565,N_2876,N_9572);
and U11566 (N_11566,N_8698,N_442);
nand U11567 (N_11567,N_5754,N_7674);
nand U11568 (N_11568,N_9065,N_3645);
nand U11569 (N_11569,N_7567,N_6696);
nand U11570 (N_11570,N_4648,N_2333);
nor U11571 (N_11571,N_5161,N_2147);
and U11572 (N_11572,N_7569,N_9221);
or U11573 (N_11573,N_4066,N_6111);
nor U11574 (N_11574,N_8286,N_2871);
or U11575 (N_11575,N_1696,N_8623);
and U11576 (N_11576,N_9318,N_6528);
or U11577 (N_11577,N_4233,N_7384);
or U11578 (N_11578,N_4716,N_8520);
and U11579 (N_11579,N_5861,N_5026);
and U11580 (N_11580,N_3825,N_2471);
nand U11581 (N_11581,N_1076,N_7226);
nand U11582 (N_11582,N_9853,N_4306);
or U11583 (N_11583,N_3423,N_9392);
or U11584 (N_11584,N_1686,N_8253);
or U11585 (N_11585,N_7984,N_872);
or U11586 (N_11586,N_1137,N_9666);
nor U11587 (N_11587,N_5068,N_8959);
nand U11588 (N_11588,N_9893,N_5341);
nand U11589 (N_11589,N_7409,N_382);
nor U11590 (N_11590,N_4613,N_6031);
and U11591 (N_11591,N_6312,N_7012);
xor U11592 (N_11592,N_6482,N_771);
and U11593 (N_11593,N_9368,N_5809);
nand U11594 (N_11594,N_7744,N_6110);
xnor U11595 (N_11595,N_9435,N_4556);
nand U11596 (N_11596,N_4115,N_3004);
and U11597 (N_11597,N_2320,N_4274);
xor U11598 (N_11598,N_6395,N_1763);
nor U11599 (N_11599,N_238,N_1494);
nand U11600 (N_11600,N_4415,N_7751);
nor U11601 (N_11601,N_4850,N_5000);
or U11602 (N_11602,N_3995,N_5763);
xor U11603 (N_11603,N_9326,N_71);
xnor U11604 (N_11604,N_5911,N_4532);
and U11605 (N_11605,N_3756,N_261);
xor U11606 (N_11606,N_2616,N_9306);
or U11607 (N_11607,N_9025,N_275);
and U11608 (N_11608,N_4109,N_4763);
or U11609 (N_11609,N_2256,N_4590);
nand U11610 (N_11610,N_3067,N_5172);
or U11611 (N_11611,N_2161,N_5944);
xnor U11612 (N_11612,N_8927,N_5462);
and U11613 (N_11613,N_1580,N_1372);
xnor U11614 (N_11614,N_4509,N_5962);
or U11615 (N_11615,N_4729,N_4529);
nand U11616 (N_11616,N_4005,N_2772);
or U11617 (N_11617,N_8938,N_9552);
nand U11618 (N_11618,N_7750,N_3793);
nand U11619 (N_11619,N_1658,N_7838);
nor U11620 (N_11620,N_8454,N_4666);
nor U11621 (N_11621,N_3290,N_7311);
xor U11622 (N_11622,N_9235,N_3313);
xor U11623 (N_11623,N_6264,N_2878);
and U11624 (N_11624,N_2610,N_556);
and U11625 (N_11625,N_4334,N_2687);
xnor U11626 (N_11626,N_1712,N_5586);
and U11627 (N_11627,N_828,N_8800);
xnor U11628 (N_11628,N_5020,N_2557);
or U11629 (N_11629,N_4604,N_1617);
or U11630 (N_11630,N_2974,N_6945);
or U11631 (N_11631,N_8673,N_4139);
or U11632 (N_11632,N_7007,N_3889);
xor U11633 (N_11633,N_1422,N_829);
nand U11634 (N_11634,N_9085,N_9473);
nor U11635 (N_11635,N_2589,N_1316);
xnor U11636 (N_11636,N_2645,N_8968);
nor U11637 (N_11637,N_9935,N_6810);
nand U11638 (N_11638,N_912,N_3314);
and U11639 (N_11639,N_168,N_2975);
nand U11640 (N_11640,N_9997,N_9596);
nor U11641 (N_11641,N_1404,N_1825);
or U11642 (N_11642,N_4154,N_3884);
nand U11643 (N_11643,N_4564,N_9544);
xor U11644 (N_11644,N_5018,N_1855);
xnor U11645 (N_11645,N_4134,N_2582);
xnor U11646 (N_11646,N_2857,N_9022);
nor U11647 (N_11647,N_6913,N_9790);
and U11648 (N_11648,N_74,N_495);
nand U11649 (N_11649,N_8553,N_6174);
xor U11650 (N_11650,N_3055,N_8714);
and U11651 (N_11651,N_3273,N_2046);
and U11652 (N_11652,N_6308,N_6321);
and U11653 (N_11653,N_2159,N_5844);
xor U11654 (N_11654,N_1924,N_6737);
xnor U11655 (N_11655,N_2184,N_2928);
xor U11656 (N_11656,N_5667,N_5102);
or U11657 (N_11657,N_2059,N_8222);
nor U11658 (N_11658,N_4825,N_9733);
and U11659 (N_11659,N_2416,N_3847);
and U11660 (N_11660,N_3811,N_8135);
nor U11661 (N_11661,N_8308,N_719);
or U11662 (N_11662,N_5638,N_4660);
nor U11663 (N_11663,N_1602,N_2541);
or U11664 (N_11664,N_3595,N_4209);
nand U11665 (N_11665,N_1355,N_8524);
or U11666 (N_11666,N_8150,N_9252);
xnor U11667 (N_11667,N_3845,N_5916);
xor U11668 (N_11668,N_6468,N_3826);
or U11669 (N_11669,N_1118,N_2747);
or U11670 (N_11670,N_6682,N_4351);
nand U11671 (N_11671,N_7906,N_5611);
and U11672 (N_11672,N_4197,N_1128);
nand U11673 (N_11673,N_5367,N_3955);
xnor U11674 (N_11674,N_6681,N_7692);
xor U11675 (N_11675,N_5614,N_7447);
and U11676 (N_11676,N_928,N_503);
and U11677 (N_11677,N_5569,N_2628);
nor U11678 (N_11678,N_7354,N_1676);
or U11679 (N_11679,N_4855,N_6725);
nand U11680 (N_11680,N_6128,N_9307);
xnor U11681 (N_11681,N_1094,N_1204);
and U11682 (N_11682,N_3574,N_3899);
and U11683 (N_11683,N_2731,N_5830);
nor U11684 (N_11684,N_7445,N_856);
nor U11685 (N_11685,N_7355,N_2905);
nand U11686 (N_11686,N_789,N_9433);
nand U11687 (N_11687,N_9714,N_741);
xor U11688 (N_11688,N_8054,N_5173);
nor U11689 (N_11689,N_5792,N_2542);
and U11690 (N_11690,N_1677,N_2443);
nand U11691 (N_11691,N_950,N_9792);
and U11692 (N_11692,N_7047,N_5936);
and U11693 (N_11693,N_18,N_9575);
nand U11694 (N_11694,N_1971,N_5308);
nand U11695 (N_11695,N_2422,N_8725);
xor U11696 (N_11696,N_7602,N_4882);
or U11697 (N_11697,N_8271,N_3876);
or U11698 (N_11698,N_7970,N_2711);
nor U11699 (N_11699,N_8999,N_6429);
or U11700 (N_11700,N_4205,N_4187);
nor U11701 (N_11701,N_2951,N_4045);
nand U11702 (N_11702,N_548,N_8160);
xnor U11703 (N_11703,N_8846,N_8338);
xor U11704 (N_11704,N_8037,N_129);
and U11705 (N_11705,N_1660,N_2025);
xnor U11706 (N_11706,N_5740,N_3673);
nor U11707 (N_11707,N_1804,N_8467);
xor U11708 (N_11708,N_2882,N_6723);
nor U11709 (N_11709,N_539,N_1028);
xnor U11710 (N_11710,N_7351,N_6634);
nand U11711 (N_11711,N_8492,N_243);
nor U11712 (N_11712,N_9591,N_346);
nand U11713 (N_11713,N_6581,N_5560);
and U11714 (N_11714,N_2906,N_1503);
nor U11715 (N_11715,N_8044,N_2580);
nor U11716 (N_11716,N_647,N_7241);
nor U11717 (N_11717,N_1061,N_357);
xor U11718 (N_11718,N_2010,N_5531);
xor U11719 (N_11719,N_9789,N_4467);
nand U11720 (N_11720,N_9687,N_3974);
or U11721 (N_11721,N_9401,N_7263);
and U11722 (N_11722,N_6700,N_6228);
nand U11723 (N_11723,N_5427,N_9019);
nor U11724 (N_11724,N_5188,N_3465);
nand U11725 (N_11725,N_2512,N_1613);
or U11726 (N_11726,N_9966,N_5590);
nor U11727 (N_11727,N_3010,N_8728);
or U11728 (N_11728,N_8687,N_9951);
or U11729 (N_11729,N_6735,N_7294);
xor U11730 (N_11730,N_2185,N_3335);
xor U11731 (N_11731,N_6866,N_8885);
nand U11732 (N_11732,N_4587,N_7621);
nor U11733 (N_11733,N_9826,N_3239);
nor U11734 (N_11734,N_3440,N_3379);
nand U11735 (N_11735,N_4683,N_5079);
and U11736 (N_11736,N_9699,N_7916);
xnor U11737 (N_11737,N_8621,N_3579);
nor U11738 (N_11738,N_3540,N_5746);
nand U11739 (N_11739,N_9535,N_5472);
nor U11740 (N_11740,N_4148,N_1581);
or U11741 (N_11741,N_9824,N_2658);
xnor U11742 (N_11742,N_5606,N_7176);
nand U11743 (N_11743,N_963,N_2843);
or U11744 (N_11744,N_6357,N_6554);
nor U11745 (N_11745,N_3868,N_5925);
or U11746 (N_11746,N_7930,N_9683);
xnor U11747 (N_11747,N_1732,N_1547);
xnor U11748 (N_11748,N_9747,N_5044);
nor U11749 (N_11749,N_7993,N_1537);
and U11750 (N_11750,N_956,N_9145);
nand U11751 (N_11751,N_3813,N_6238);
nor U11752 (N_11752,N_1684,N_9822);
or U11753 (N_11753,N_338,N_3644);
xnor U11754 (N_11754,N_9063,N_480);
nor U11755 (N_11755,N_2045,N_8411);
nand U11756 (N_11756,N_2056,N_689);
nand U11757 (N_11757,N_8678,N_2705);
nor U11758 (N_11758,N_9668,N_4353);
or U11759 (N_11759,N_1225,N_3309);
or U11760 (N_11760,N_2653,N_1282);
or U11761 (N_11761,N_2877,N_3177);
or U11762 (N_11762,N_2621,N_9889);
or U11763 (N_11763,N_4010,N_1745);
nand U11764 (N_11764,N_1418,N_2624);
nor U11765 (N_11765,N_3960,N_7306);
nor U11766 (N_11766,N_3444,N_4416);
and U11767 (N_11767,N_8990,N_3299);
nor U11768 (N_11768,N_36,N_5138);
nand U11769 (N_11769,N_533,N_8561);
nand U11770 (N_11770,N_2751,N_899);
xnor U11771 (N_11771,N_1585,N_2510);
or U11772 (N_11772,N_4083,N_5151);
and U11773 (N_11773,N_6684,N_8112);
xor U11774 (N_11774,N_7230,N_9037);
nand U11775 (N_11775,N_4610,N_9043);
xor U11776 (N_11776,N_7347,N_2062);
xnor U11777 (N_11777,N_9564,N_3328);
nor U11778 (N_11778,N_2523,N_431);
or U11779 (N_11779,N_6281,N_665);
nor U11780 (N_11780,N_1512,N_5345);
xor U11781 (N_11781,N_8041,N_543);
nor U11782 (N_11782,N_861,N_616);
and U11783 (N_11783,N_4795,N_9612);
nor U11784 (N_11784,N_9952,N_1301);
nand U11785 (N_11785,N_840,N_8745);
nand U11786 (N_11786,N_7776,N_2826);
nor U11787 (N_11787,N_2632,N_8193);
or U11788 (N_11788,N_3832,N_3409);
or U11789 (N_11789,N_2569,N_2726);
nand U11790 (N_11790,N_2312,N_125);
and U11791 (N_11791,N_9016,N_32);
and U11792 (N_11792,N_3408,N_9223);
xnor U11793 (N_11793,N_5824,N_1181);
nor U11794 (N_11794,N_1939,N_2130);
xor U11795 (N_11795,N_216,N_9107);
and U11796 (N_11796,N_8738,N_2534);
xor U11797 (N_11797,N_390,N_5115);
and U11798 (N_11798,N_6701,N_9166);
xnor U11799 (N_11799,N_2268,N_826);
and U11800 (N_11800,N_1993,N_9174);
or U11801 (N_11801,N_9982,N_7211);
nor U11802 (N_11802,N_8505,N_2177);
and U11803 (N_11803,N_5685,N_4941);
nor U11804 (N_11804,N_3,N_7014);
nand U11805 (N_11805,N_3617,N_3862);
and U11806 (N_11806,N_9197,N_6604);
and U11807 (N_11807,N_5003,N_5566);
or U11808 (N_11808,N_6542,N_2375);
or U11809 (N_11809,N_4502,N_3355);
nand U11810 (N_11810,N_3495,N_8220);
xnor U11811 (N_11811,N_5528,N_8460);
xor U11812 (N_11812,N_7511,N_709);
nor U11813 (N_11813,N_3259,N_2496);
xor U11814 (N_11814,N_5671,N_7519);
nand U11815 (N_11815,N_791,N_423);
nand U11816 (N_11816,N_1371,N_2592);
xor U11817 (N_11817,N_9377,N_2715);
or U11818 (N_11818,N_334,N_4014);
xor U11819 (N_11819,N_6673,N_3118);
xor U11820 (N_11820,N_5247,N_5232);
nor U11821 (N_11821,N_1273,N_5022);
nand U11822 (N_11822,N_3245,N_6121);
nor U11823 (N_11823,N_2730,N_7134);
or U11824 (N_11824,N_7765,N_2262);
nand U11825 (N_11825,N_4224,N_685);
and U11826 (N_11826,N_9031,N_3570);
or U11827 (N_11827,N_356,N_3802);
nor U11828 (N_11828,N_7725,N_7605);
xnor U11829 (N_11829,N_1742,N_9258);
or U11830 (N_11830,N_1250,N_6513);
xor U11831 (N_11831,N_1270,N_8133);
and U11832 (N_11832,N_1941,N_3267);
or U11833 (N_11833,N_7614,N_4919);
or U11834 (N_11834,N_8244,N_3158);
nand U11835 (N_11835,N_3185,N_9432);
xor U11836 (N_11836,N_2671,N_9685);
xnor U11837 (N_11837,N_8804,N_1915);
nand U11838 (N_11838,N_1589,N_8651);
nor U11839 (N_11839,N_7499,N_2729);
nand U11840 (N_11840,N_9239,N_5509);
or U11841 (N_11841,N_183,N_3783);
xnor U11842 (N_11842,N_7870,N_2028);
nor U11843 (N_11843,N_5260,N_9536);
xor U11844 (N_11844,N_5255,N_9282);
nor U11845 (N_11845,N_4859,N_9801);
and U11846 (N_11846,N_5552,N_3623);
and U11847 (N_11847,N_2568,N_9599);
and U11848 (N_11848,N_9319,N_9842);
nand U11849 (N_11849,N_33,N_6524);
nand U11850 (N_11850,N_5315,N_5794);
nor U11851 (N_11851,N_1340,N_854);
or U11852 (N_11852,N_7575,N_4589);
nand U11853 (N_11853,N_2717,N_222);
nor U11854 (N_11854,N_1935,N_6631);
and U11855 (N_11855,N_2766,N_8775);
nand U11856 (N_11856,N_5719,N_606);
xnor U11857 (N_11857,N_8494,N_1905);
nor U11858 (N_11858,N_3407,N_9494);
or U11859 (N_11859,N_4105,N_5931);
and U11860 (N_11860,N_6175,N_7707);
and U11861 (N_11861,N_8414,N_5214);
xor U11862 (N_11862,N_9417,N_7322);
or U11863 (N_11863,N_9257,N_1999);
nand U11864 (N_11864,N_8266,N_5998);
or U11865 (N_11865,N_2063,N_2414);
or U11866 (N_11866,N_7256,N_835);
or U11867 (N_11867,N_805,N_6527);
nand U11868 (N_11868,N_535,N_380);
nor U11869 (N_11869,N_7899,N_1607);
nand U11870 (N_11870,N_1584,N_2823);
and U11871 (N_11871,N_8749,N_7032);
or U11872 (N_11872,N_8144,N_670);
or U11873 (N_11873,N_4899,N_4600);
nand U11874 (N_11874,N_2664,N_5705);
or U11875 (N_11875,N_386,N_4180);
nor U11876 (N_11876,N_9582,N_4738);
xor U11877 (N_11877,N_6948,N_8198);
xor U11878 (N_11878,N_2536,N_8667);
and U11879 (N_11879,N_2255,N_2438);
nand U11880 (N_11880,N_6843,N_6928);
and U11881 (N_11881,N_5848,N_3854);
or U11882 (N_11882,N_9034,N_2462);
and U11883 (N_11883,N_9782,N_2919);
nor U11884 (N_11884,N_2521,N_515);
xor U11885 (N_11885,N_2680,N_2212);
or U11886 (N_11886,N_1022,N_9795);
nor U11887 (N_11887,N_6667,N_3881);
xor U11888 (N_11888,N_3318,N_1682);
or U11889 (N_11889,N_7076,N_5162);
nand U11890 (N_11890,N_171,N_9180);
nand U11891 (N_11891,N_2814,N_201);
xor U11892 (N_11892,N_857,N_8937);
or U11893 (N_11893,N_1257,N_8920);
or U11894 (N_11894,N_3012,N_3174);
and U11895 (N_11895,N_3614,N_474);
or U11896 (N_11896,N_5694,N_4478);
nor U11897 (N_11897,N_7108,N_8148);
xor U11898 (N_11898,N_7407,N_7778);
and U11899 (N_11899,N_6800,N_8019);
or U11900 (N_11900,N_1497,N_9720);
xor U11901 (N_11901,N_6568,N_4443);
nor U11902 (N_11902,N_8654,N_1388);
xnor U11903 (N_11903,N_1556,N_4984);
nor U11904 (N_11904,N_3780,N_4699);
nand U11905 (N_11905,N_7498,N_1032);
nand U11906 (N_11906,N_9329,N_1535);
nand U11907 (N_11907,N_8137,N_1053);
nor U11908 (N_11908,N_121,N_6146);
nor U11909 (N_11909,N_9976,N_8573);
nand U11910 (N_11910,N_6901,N_3647);
and U11911 (N_11911,N_6669,N_2663);
nor U11912 (N_11912,N_3150,N_4764);
and U11913 (N_11913,N_4108,N_7326);
and U11914 (N_11914,N_5175,N_1848);
or U11915 (N_11915,N_8311,N_4386);
nor U11916 (N_11916,N_932,N_6603);
or U11917 (N_11917,N_2228,N_5288);
nand U11918 (N_11918,N_5624,N_917);
nand U11919 (N_11919,N_6801,N_9895);
xnor U11920 (N_11920,N_6143,N_9010);
or U11921 (N_11921,N_3044,N_5243);
nand U11922 (N_11922,N_2576,N_7290);
xnor U11923 (N_11923,N_8419,N_4827);
nand U11924 (N_11924,N_2620,N_3589);
and U11925 (N_11925,N_4032,N_4831);
and U11926 (N_11926,N_8665,N_6457);
or U11927 (N_11927,N_21,N_5805);
xnor U11928 (N_11928,N_4280,N_1653);
and U11929 (N_11929,N_1001,N_8255);
xnor U11930 (N_11930,N_959,N_6910);
nand U11931 (N_11931,N_2459,N_3051);
nand U11932 (N_11932,N_6704,N_4971);
xnor U11933 (N_11933,N_5903,N_4750);
nor U11934 (N_11934,N_9519,N_3208);
nand U11935 (N_11935,N_4951,N_6481);
or U11936 (N_11936,N_4159,N_3789);
and U11937 (N_11937,N_1832,N_5037);
nand U11938 (N_11938,N_8597,N_7399);
xnor U11939 (N_11939,N_6821,N_3395);
xor U11940 (N_11940,N_8807,N_4696);
xor U11941 (N_11941,N_4301,N_1650);
nand U11942 (N_11942,N_3443,N_6361);
nor U11943 (N_11943,N_7734,N_116);
nor U11944 (N_11944,N_5827,N_4830);
xnor U11945 (N_11945,N_1099,N_9986);
xnor U11946 (N_11946,N_2348,N_387);
or U11947 (N_11947,N_8677,N_9709);
nor U11948 (N_11948,N_834,N_693);
nand U11949 (N_11949,N_7296,N_4704);
or U11950 (N_11950,N_1455,N_985);
and U11951 (N_11951,N_5233,N_7160);
xnor U11952 (N_11952,N_8892,N_8526);
nor U11953 (N_11953,N_5620,N_2299);
nand U11954 (N_11954,N_7045,N_8239);
and U11955 (N_11955,N_9155,N_4207);
and U11956 (N_11956,N_7087,N_1484);
xnor U11957 (N_11957,N_972,N_8047);
or U11958 (N_11958,N_5258,N_2691);
or U11959 (N_11959,N_2488,N_597);
and U11960 (N_11960,N_377,N_6288);
nand U11961 (N_11961,N_6421,N_2007);
nor U11962 (N_11962,N_593,N_7441);
and U11963 (N_11963,N_8191,N_8566);
nand U11964 (N_11964,N_6734,N_8765);
or U11965 (N_11965,N_5058,N_7382);
nor U11966 (N_11966,N_3049,N_6025);
or U11967 (N_11967,N_8789,N_1217);
xnor U11968 (N_11968,N_6770,N_9078);
xor U11969 (N_11969,N_6702,N_7497);
and U11970 (N_11970,N_6272,N_439);
or U11971 (N_11971,N_4534,N_7321);
xor U11972 (N_11972,N_1895,N_4090);
and U11973 (N_11973,N_4263,N_5508);
or U11974 (N_11974,N_4474,N_3603);
and U11975 (N_11975,N_623,N_7138);
nor U11976 (N_11976,N_1256,N_6614);
xor U11977 (N_11977,N_7714,N_4327);
xor U11978 (N_11978,N_1889,N_7449);
and U11979 (N_11979,N_2482,N_267);
xor U11980 (N_11980,N_1697,N_5278);
xnor U11981 (N_11981,N_8637,N_3357);
xor U11982 (N_11982,N_3448,N_4008);
or U11983 (N_11983,N_3576,N_564);
or U11984 (N_11984,N_8495,N_997);
nor U11985 (N_11985,N_5862,N_9353);
nor U11986 (N_11986,N_3843,N_4707);
nor U11987 (N_11987,N_6868,N_1492);
or U11988 (N_11988,N_4539,N_4569);
and U11989 (N_11989,N_5674,N_1819);
nor U11990 (N_11990,N_6846,N_6556);
nand U11991 (N_11991,N_5864,N_6268);
nor U11992 (N_11992,N_2669,N_5649);
nand U11993 (N_11993,N_355,N_1452);
or U11994 (N_11994,N_6898,N_9456);
xnor U11995 (N_11995,N_8684,N_9068);
nand U11996 (N_11996,N_4920,N_1554);
nor U11997 (N_11997,N_4039,N_2992);
or U11998 (N_11998,N_1038,N_9379);
nor U11999 (N_11999,N_9984,N_1822);
nor U12000 (N_12000,N_9490,N_6600);
or U12001 (N_12001,N_2763,N_9922);
xnor U12002 (N_12002,N_4940,N_8891);
xor U12003 (N_12003,N_4641,N_8098);
and U12004 (N_12004,N_6150,N_786);
and U12005 (N_12005,N_7131,N_3386);
or U12006 (N_12006,N_6550,N_7001);
xor U12007 (N_12007,N_1836,N_2444);
or U12008 (N_12008,N_5218,N_3561);
nand U12009 (N_12009,N_655,N_3333);
nor U12010 (N_12010,N_8055,N_3428);
nand U12011 (N_12011,N_4387,N_1538);
xnor U12012 (N_12012,N_2566,N_7822);
nor U12013 (N_12013,N_2009,N_668);
xor U12014 (N_12014,N_2084,N_4278);
and U12015 (N_12015,N_2646,N_3521);
nor U12016 (N_12016,N_1338,N_9954);
xor U12017 (N_12017,N_3663,N_3818);
or U12018 (N_12018,N_8341,N_6938);
nand U12019 (N_12019,N_7019,N_1205);
nand U12020 (N_12020,N_6871,N_1695);
xnor U12021 (N_12021,N_4559,N_5323);
nor U12022 (N_12022,N_8650,N_5516);
nand U12023 (N_12023,N_9274,N_4702);
nand U12024 (N_12024,N_4024,N_9630);
and U12025 (N_12025,N_6893,N_5061);
and U12026 (N_12026,N_7717,N_3597);
or U12027 (N_12027,N_4801,N_3901);
and U12028 (N_12028,N_7601,N_2192);
nand U12029 (N_12029,N_4323,N_5605);
nand U12030 (N_12030,N_4229,N_5826);
xnor U12031 (N_12031,N_2815,N_4166);
or U12032 (N_12032,N_3670,N_9547);
xor U12033 (N_12033,N_5455,N_4448);
or U12034 (N_12034,N_4562,N_838);
nand U12035 (N_12035,N_7271,N_4786);
nand U12036 (N_12036,N_3140,N_4175);
or U12037 (N_12037,N_3471,N_3833);
nor U12038 (N_12038,N_710,N_4176);
or U12039 (N_12039,N_4111,N_3578);
or U12040 (N_12040,N_8462,N_2431);
and U12041 (N_12041,N_7885,N_6891);
and U12042 (N_12042,N_9962,N_5371);
or U12043 (N_12043,N_7965,N_9987);
and U12044 (N_12044,N_4906,N_2365);
or U12045 (N_12045,N_6145,N_7397);
xnor U12046 (N_12046,N_185,N_9220);
nand U12047 (N_12047,N_5487,N_6207);
nand U12048 (N_12048,N_251,N_5356);
nor U12049 (N_12049,N_8204,N_8345);
nand U12050 (N_12050,N_5449,N_257);
and U12051 (N_12051,N_1711,N_6042);
xor U12052 (N_12052,N_1883,N_3991);
xor U12053 (N_12053,N_4943,N_4240);
xnor U12054 (N_12054,N_5828,N_3213);
or U12055 (N_12055,N_5687,N_7535);
nand U12056 (N_12056,N_507,N_7200);
nand U12057 (N_12057,N_6511,N_6297);
nor U12058 (N_12058,N_8229,N_4146);
nor U12059 (N_12059,N_3054,N_6534);
nand U12060 (N_12060,N_4341,N_9793);
nor U12061 (N_12061,N_7688,N_8921);
or U12062 (N_12062,N_6503,N_6636);
xnor U12063 (N_12063,N_7316,N_5360);
nor U12064 (N_12064,N_4145,N_9915);
nor U12065 (N_12065,N_6999,N_8993);
nor U12066 (N_12066,N_6567,N_7043);
nand U12067 (N_12067,N_17,N_3163);
or U12068 (N_12068,N_7198,N_2149);
nand U12069 (N_12069,N_2675,N_2999);
or U12070 (N_12070,N_463,N_4615);
and U12071 (N_12071,N_1768,N_3075);
or U12072 (N_12072,N_3610,N_43);
or U12073 (N_12073,N_9980,N_1588);
and U12074 (N_12074,N_5623,N_4490);
xnor U12075 (N_12075,N_8642,N_9402);
or U12076 (N_12076,N_2283,N_6066);
nor U12077 (N_12077,N_8630,N_4921);
and U12078 (N_12078,N_3345,N_8169);
nand U12079 (N_12079,N_823,N_5567);
nor U12080 (N_12080,N_373,N_1150);
and U12081 (N_12081,N_5475,N_1396);
nor U12082 (N_12082,N_7858,N_483);
and U12083 (N_12083,N_6978,N_7800);
nand U12084 (N_12084,N_111,N_2096);
nor U12085 (N_12085,N_5150,N_955);
nor U12086 (N_12086,N_8551,N_4022);
or U12087 (N_12087,N_5357,N_3175);
xnor U12088 (N_12088,N_4577,N_8100);
and U12089 (N_12089,N_1725,N_415);
nand U12090 (N_12090,N_2997,N_3207);
nand U12091 (N_12091,N_6510,N_9441);
xnor U12092 (N_12092,N_8302,N_7908);
and U12093 (N_12093,N_9584,N_1675);
nand U12094 (N_12094,N_6057,N_7467);
and U12095 (N_12095,N_4276,N_8629);
xnor U12096 (N_12096,N_3526,N_2068);
xnor U12097 (N_12097,N_7582,N_3569);
and U12098 (N_12098,N_4868,N_7282);
or U12099 (N_12099,N_4555,N_6036);
xnor U12100 (N_12100,N_2914,N_8529);
or U12101 (N_12101,N_8161,N_5417);
or U12102 (N_12102,N_4434,N_4464);
and U12103 (N_12103,N_2514,N_5905);
xor U12104 (N_12104,N_8970,N_645);
and U12105 (N_12105,N_6765,N_8762);
nand U12106 (N_12106,N_7878,N_4896);
nand U12107 (N_12107,N_920,N_6393);
nand U12108 (N_12108,N_9453,N_923);
nand U12109 (N_12109,N_3365,N_1347);
or U12110 (N_12110,N_400,N_3346);
and U12111 (N_12111,N_5968,N_5376);
nand U12112 (N_12112,N_3585,N_3026);
and U12113 (N_12113,N_3126,N_2758);
nor U12114 (N_12114,N_5712,N_6501);
xor U12115 (N_12115,N_5665,N_9881);
and U12116 (N_12116,N_4853,N_5133);
nor U12117 (N_12117,N_7523,N_6427);
and U12118 (N_12118,N_9079,N_4500);
nand U12119 (N_12119,N_2982,N_1979);
nor U12120 (N_12120,N_4774,N_8560);
xnor U12121 (N_12121,N_5822,N_7662);
or U12122 (N_12122,N_6506,N_4996);
nor U12123 (N_12123,N_1495,N_2143);
xnor U12124 (N_12124,N_6340,N_7299);
nor U12125 (N_12125,N_7565,N_7593);
nor U12126 (N_12126,N_6279,N_5075);
and U12127 (N_12127,N_4865,N_4221);
or U12128 (N_12128,N_2152,N_8645);
nor U12129 (N_12129,N_2200,N_3822);
and U12130 (N_12130,N_706,N_3982);
nand U12131 (N_12131,N_3413,N_4132);
nand U12132 (N_12132,N_9836,N_2315);
nor U12133 (N_12133,N_5557,N_4088);
and U12134 (N_12134,N_9204,N_8694);
nor U12135 (N_12135,N_3742,N_5057);
nand U12136 (N_12136,N_1618,N_3749);
and U12137 (N_12137,N_790,N_1635);
and U12138 (N_12138,N_8797,N_5374);
nor U12139 (N_12139,N_8546,N_6853);
nor U12140 (N_12140,N_4761,N_3769);
nor U12141 (N_12141,N_9909,N_7187);
xor U12142 (N_12142,N_3455,N_8136);
and U12143 (N_12143,N_3358,N_8409);
nor U12144 (N_12144,N_1049,N_9818);
xnor U12145 (N_12145,N_1370,N_5142);
xnor U12146 (N_12146,N_2123,N_9238);
nand U12147 (N_12147,N_4085,N_8189);
nand U12148 (N_12148,N_5297,N_7739);
nand U12149 (N_12149,N_4192,N_7245);
nor U12150 (N_12150,N_3479,N_7873);
nor U12151 (N_12151,N_40,N_2050);
nor U12152 (N_12152,N_3100,N_3828);
and U12153 (N_12153,N_9894,N_2721);
and U12154 (N_12154,N_5837,N_4246);
xor U12155 (N_12155,N_9877,N_213);
xor U12156 (N_12156,N_5159,N_7379);
and U12157 (N_12157,N_303,N_5874);
nand U12158 (N_12158,N_1295,N_1717);
xor U12159 (N_12159,N_4298,N_1641);
or U12160 (N_12160,N_6164,N_7552);
nand U12161 (N_12161,N_8485,N_7058);
nand U12162 (N_12162,N_6580,N_3501);
xor U12163 (N_12163,N_1798,N_9236);
nor U12164 (N_12164,N_6019,N_4058);
nor U12165 (N_12165,N_3909,N_3556);
and U12166 (N_12166,N_4079,N_3039);
xor U12167 (N_12167,N_5815,N_6591);
xnor U12168 (N_12168,N_2166,N_1615);
xnor U12169 (N_12169,N_8201,N_3276);
xor U12170 (N_12170,N_4362,N_4568);
nand U12171 (N_12171,N_82,N_4466);
nand U12172 (N_12172,N_2107,N_7375);
nand U12173 (N_12173,N_8210,N_6714);
nand U12174 (N_12174,N_6827,N_5739);
or U12175 (N_12175,N_7689,N_1149);
or U12176 (N_12176,N_3091,N_5585);
or U12177 (N_12177,N_4799,N_970);
nor U12178 (N_12178,N_9267,N_4358);
and U12179 (N_12179,N_973,N_4947);
xnor U12180 (N_12180,N_1491,N_8502);
nor U12181 (N_12181,N_5889,N_4886);
and U12182 (N_12182,N_4863,N_841);
and U12183 (N_12183,N_9653,N_5166);
nand U12184 (N_12184,N_9949,N_109);
or U12185 (N_12185,N_6499,N_4989);
and U12186 (N_12186,N_8332,N_5346);
nor U12187 (N_12187,N_7594,N_8680);
nor U12188 (N_12188,N_2735,N_7793);
xnor U12189 (N_12189,N_3135,N_3871);
and U12190 (N_12190,N_2517,N_8129);
xor U12191 (N_12191,N_8894,N_3558);
or U12192 (N_12192,N_7978,N_8554);
xnor U12193 (N_12193,N_1867,N_5641);
and U12194 (N_12194,N_9669,N_9463);
nand U12195 (N_12195,N_1212,N_7823);
or U12196 (N_12196,N_266,N_3303);
nor U12197 (N_12197,N_1721,N_2327);
nor U12198 (N_12198,N_604,N_1678);
or U12199 (N_12199,N_6851,N_8769);
and U12200 (N_12200,N_6803,N_4390);
and U12201 (N_12201,N_9393,N_9880);
xnor U12202 (N_12202,N_5587,N_3231);
nor U12203 (N_12203,N_6009,N_5194);
and U12204 (N_12204,N_7304,N_6747);
xnor U12205 (N_12205,N_3133,N_4150);
and U12206 (N_12206,N_7914,N_8326);
and U12207 (N_12207,N_7300,N_4314);
and U12208 (N_12208,N_1470,N_241);
nor U12209 (N_12209,N_3765,N_6680);
nor U12210 (N_12210,N_1683,N_6167);
and U12211 (N_12211,N_7297,N_9778);
and U12212 (N_12212,N_5192,N_8093);
or U12213 (N_12213,N_4937,N_2183);
nor U12214 (N_12214,N_6419,N_4881);
and U12215 (N_12215,N_3451,N_6123);
and U12216 (N_12216,N_4053,N_5433);
nor U12217 (N_12217,N_4717,N_9907);
nor U12218 (N_12218,N_3189,N_8528);
xnor U12219 (N_12219,N_8655,N_2685);
nand U12220 (N_12220,N_754,N_9374);
nand U12221 (N_12221,N_7155,N_6101);
xor U12222 (N_12222,N_765,N_2395);
or U12223 (N_12223,N_6629,N_596);
and U12224 (N_12224,N_6090,N_9887);
and U12225 (N_12225,N_1890,N_7405);
nand U12226 (N_12226,N_9309,N_506);
xor U12227 (N_12227,N_4130,N_7901);
or U12228 (N_12228,N_4470,N_294);
nor U12229 (N_12229,N_4585,N_4772);
nand U12230 (N_12230,N_1901,N_6210);
xnor U12231 (N_12231,N_5576,N_484);
xnor U12232 (N_12232,N_8496,N_4047);
nand U12233 (N_12233,N_9304,N_3735);
nand U12234 (N_12234,N_3473,N_9914);
nor U12235 (N_12235,N_3716,N_176);
xor U12236 (N_12236,N_3193,N_1362);
nand U12237 (N_12237,N_6436,N_778);
and U12238 (N_12238,N_7543,N_416);
or U12239 (N_12239,N_1030,N_5493);
and U12240 (N_12240,N_8862,N_9191);
nor U12241 (N_12241,N_9745,N_990);
and U12242 (N_12242,N_4606,N_174);
nand U12243 (N_12243,N_9160,N_4087);
or U12244 (N_12244,N_5252,N_4936);
nand U12245 (N_12245,N_7904,N_5593);
and U12246 (N_12246,N_1285,N_7159);
and U12247 (N_12247,N_878,N_5084);
xor U12248 (N_12248,N_8724,N_941);
or U12249 (N_12249,N_8783,N_8608);
nor U12250 (N_12250,N_9534,N_4335);
or U12251 (N_12251,N_3515,N_6977);
and U12252 (N_12252,N_1910,N_3546);
xor U12253 (N_12253,N_7432,N_6236);
or U12254 (N_12254,N_1736,N_1688);
or U12255 (N_12255,N_7073,N_4195);
xor U12256 (N_12256,N_5676,N_9106);
nor U12257 (N_12257,N_673,N_4297);
nor U12258 (N_12258,N_2170,N_1927);
nor U12259 (N_12259,N_4371,N_1636);
xnor U12260 (N_12260,N_4396,N_3861);
or U12261 (N_12261,N_8297,N_8583);
nor U12262 (N_12262,N_7259,N_3761);
or U12263 (N_12263,N_9317,N_1722);
nor U12264 (N_12264,N_4241,N_5107);
nand U12265 (N_12265,N_643,N_7571);
or U12266 (N_12266,N_6931,N_6545);
xnor U12267 (N_12267,N_1027,N_9082);
nand U12268 (N_12268,N_641,N_1610);
or U12269 (N_12269,N_1356,N_5736);
or U12270 (N_12270,N_3322,N_6179);
nand U12271 (N_12271,N_8835,N_4640);
nand U12272 (N_12272,N_7695,N_1866);
and U12273 (N_12273,N_633,N_8176);
nand U12274 (N_12274,N_6235,N_6402);
or U12275 (N_12275,N_2088,N_1994);
xor U12276 (N_12276,N_4601,N_7170);
nand U12277 (N_12277,N_6372,N_8361);
nor U12278 (N_12278,N_2812,N_7000);
nand U12279 (N_12279,N_9902,N_3470);
and U12280 (N_12280,N_1738,N_6456);
nor U12281 (N_12281,N_7033,N_2874);
xor U12282 (N_12282,N_5420,N_5536);
and U12283 (N_12283,N_7762,N_711);
and U12284 (N_12284,N_4565,N_4382);
nor U12285 (N_12285,N_6364,N_5454);
nand U12286 (N_12286,N_6873,N_6037);
nand U12287 (N_12287,N_4125,N_342);
xor U12288 (N_12288,N_2803,N_638);
or U12289 (N_12289,N_4968,N_5103);
nand U12290 (N_12290,N_5807,N_8732);
xnor U12291 (N_12291,N_1386,N_7900);
nor U12292 (N_12292,N_2850,N_1136);
nand U12293 (N_12293,N_9217,N_8669);
xor U12294 (N_12294,N_1352,N_5144);
nand U12295 (N_12295,N_1194,N_4107);
and U12296 (N_12296,N_5334,N_3202);
xor U12297 (N_12297,N_4226,N_8845);
xor U12298 (N_12298,N_6775,N_4419);
nor U12299 (N_12299,N_5997,N_5681);
nand U12300 (N_12300,N_7205,N_8082);
xnor U12301 (N_12301,N_2955,N_4449);
and U12302 (N_12302,N_4705,N_8018);
nor U12303 (N_12303,N_7302,N_7818);
xnor U12304 (N_12304,N_7851,N_8690);
nor U12305 (N_12305,N_160,N_6529);
nor U12306 (N_12306,N_9141,N_4667);
or U12307 (N_12307,N_7055,N_9554);
nand U12308 (N_12308,N_92,N_6540);
nand U12309 (N_12309,N_148,N_9567);
or U12310 (N_12310,N_7123,N_7634);
and U12311 (N_12311,N_1977,N_1409);
nor U12312 (N_12312,N_6830,N_6230);
or U12313 (N_12313,N_680,N_4096);
or U12314 (N_12314,N_4437,N_1110);
or U12315 (N_12315,N_4068,N_9616);
nor U12316 (N_12316,N_2978,N_5709);
xor U12317 (N_12317,N_172,N_1444);
nor U12318 (N_12318,N_1165,N_426);
and U12319 (N_12319,N_8396,N_4633);
nor U12320 (N_12320,N_8547,N_5239);
and U12321 (N_12321,N_3363,N_6399);
nor U12322 (N_12322,N_4913,N_370);
xor U12323 (N_12323,N_1561,N_7799);
or U12324 (N_12324,N_3762,N_1929);
or U12325 (N_12325,N_4168,N_7889);
nor U12326 (N_12326,N_3680,N_7830);
xor U12327 (N_12327,N_7083,N_9682);
and U12328 (N_12328,N_9247,N_5474);
and U12329 (N_12329,N_7563,N_6089);
xnor U12330 (N_12330,N_4669,N_6099);
nand U12331 (N_12331,N_5099,N_5511);
or U12332 (N_12332,N_7348,N_9087);
nand U12333 (N_12333,N_8899,N_881);
nand U12334 (N_12334,N_6555,N_6854);
nor U12335 (N_12335,N_4183,N_7610);
xor U12336 (N_12336,N_4781,N_7366);
or U12337 (N_12337,N_164,N_3741);
nor U12338 (N_12338,N_6815,N_86);
xnor U12339 (N_12339,N_2985,N_9618);
or U12340 (N_12340,N_3336,N_7721);
or U12341 (N_12341,N_5481,N_9114);
nor U12342 (N_12342,N_6964,N_8771);
xnor U12343 (N_12343,N_5806,N_5464);
and U12344 (N_12344,N_5540,N_8685);
or U12345 (N_12345,N_9605,N_1193);
nor U12346 (N_12346,N_4566,N_5910);
nand U12347 (N_12347,N_1005,N_5494);
nor U12348 (N_12348,N_6136,N_2191);
nand U12349 (N_12349,N_3251,N_6490);
nand U12350 (N_12350,N_9215,N_6718);
nand U12351 (N_12351,N_1305,N_2091);
or U12352 (N_12352,N_2797,N_2562);
xnor U12353 (N_12353,N_9858,N_2464);
xor U12354 (N_12354,N_2273,N_8601);
and U12355 (N_12355,N_12,N_1389);
nor U12356 (N_12356,N_3700,N_1816);
nand U12357 (N_12357,N_60,N_6839);
nand U12358 (N_12358,N_3396,N_1182);
nor U12359 (N_12359,N_6925,N_915);
nor U12360 (N_12360,N_8225,N_1445);
xor U12361 (N_12361,N_51,N_322);
xor U12362 (N_12362,N_5351,N_4519);
and U12363 (N_12363,N_8857,N_6450);
nand U12364 (N_12364,N_5298,N_1104);
nor U12365 (N_12365,N_3350,N_6390);
nand U12366 (N_12366,N_5710,N_4994);
or U12367 (N_12367,N_3159,N_8096);
and U12368 (N_12368,N_8120,N_228);
nand U12369 (N_12369,N_9925,N_5814);
or U12370 (N_12370,N_5025,N_2241);
xor U12371 (N_12371,N_1234,N_9363);
nor U12372 (N_12372,N_5344,N_815);
and U12373 (N_12373,N_2171,N_1998);
xor U12374 (N_12374,N_9437,N_1575);
nand U12375 (N_12375,N_273,N_9729);
xnor U12376 (N_12376,N_2565,N_3253);
nor U12377 (N_12377,N_3389,N_6396);
nor U12378 (N_12378,N_1810,N_9157);
or U12379 (N_12379,N_4491,N_4228);
xor U12380 (N_12380,N_490,N_2830);
xnor U12381 (N_12381,N_3064,N_229);
and U12382 (N_12382,N_4956,N_4344);
and U12383 (N_12383,N_8061,N_4157);
and U12384 (N_12384,N_7065,N_113);
or U12385 (N_12385,N_2560,N_4245);
and U12386 (N_12386,N_2169,N_2690);
or U12387 (N_12387,N_6115,N_6869);
xor U12388 (N_12388,N_520,N_5186);
or U12389 (N_12389,N_724,N_9609);
and U12390 (N_12390,N_2322,N_9481);
and U12391 (N_12391,N_9834,N_5795);
nor U12392 (N_12392,N_7057,N_2641);
nand U12393 (N_12393,N_7704,N_3787);
nand U12394 (N_12394,N_2981,N_223);
or U12395 (N_12395,N_2195,N_1073);
nor U12396 (N_12396,N_1060,N_3782);
or U12397 (N_12397,N_5432,N_1851);
and U12398 (N_12398,N_3947,N_1849);
or U12399 (N_12399,N_4378,N_5529);
nor U12400 (N_12400,N_6985,N_2538);
nand U12401 (N_12401,N_7426,N_4901);
xnor U12402 (N_12402,N_3110,N_5163);
xor U12403 (N_12403,N_8773,N_4974);
and U12404 (N_12404,N_9611,N_5090);
nand U12405 (N_12405,N_2533,N_5092);
or U12406 (N_12406,N_949,N_9051);
nand U12407 (N_12407,N_2367,N_2870);
or U12408 (N_12408,N_3152,N_5870);
and U12409 (N_12409,N_3908,N_4441);
and U12410 (N_12410,N_5135,N_3178);
nand U12411 (N_12411,N_2841,N_7849);
nor U12412 (N_12412,N_8913,N_1058);
xnor U12413 (N_12413,N_1342,N_2291);
nand U12414 (N_12414,N_99,N_4189);
or U12415 (N_12415,N_4059,N_6544);
or U12416 (N_12416,N_3951,N_8423);
nand U12417 (N_12417,N_4975,N_4800);
xor U12418 (N_12418,N_61,N_5964);
and U12419 (N_12419,N_8015,N_8217);
or U12420 (N_12420,N_9870,N_3921);
nor U12421 (N_12421,N_6790,N_5752);
or U12422 (N_12422,N_8435,N_8809);
xor U12423 (N_12423,N_1499,N_9994);
xor U12424 (N_12424,N_6049,N_3750);
or U12425 (N_12425,N_7929,N_4271);
nor U12426 (N_12426,N_3375,N_3754);
and U12427 (N_12427,N_1056,N_4731);
nand U12428 (N_12428,N_2155,N_6354);
or U12429 (N_12429,N_4191,N_8384);
xnor U12430 (N_12430,N_6796,N_4374);
nor U12431 (N_12431,N_2020,N_3197);
or U12432 (N_12432,N_75,N_5492);
nand U12433 (N_12433,N_1114,N_5912);
nand U12434 (N_12434,N_5873,N_9314);
or U12435 (N_12435,N_8192,N_5631);
and U12436 (N_12436,N_7378,N_7896);
nand U12437 (N_12437,N_4754,N_1307);
xnor U12438 (N_12438,N_7968,N_2881);
and U12439 (N_12439,N_3349,N_3771);
and U12440 (N_12440,N_4135,N_4357);
xnor U12441 (N_12441,N_6169,N_3839);
or U12442 (N_12442,N_6943,N_6350);
and U12443 (N_12443,N_6754,N_7578);
nand U12444 (N_12444,N_6820,N_3958);
nor U12445 (N_12445,N_5176,N_2532);
or U12446 (N_12446,N_6912,N_7502);
nand U12447 (N_12447,N_8533,N_1817);
nor U12448 (N_12448,N_1359,N_3393);
and U12449 (N_12449,N_7084,N_2824);
or U12450 (N_12450,N_1066,N_5941);
nand U12451 (N_12451,N_2453,N_527);
nor U12452 (N_12452,N_5437,N_4287);
nand U12453 (N_12453,N_1173,N_6118);
or U12454 (N_12454,N_3410,N_8759);
xnor U12455 (N_12455,N_571,N_9734);
nand U12456 (N_12456,N_7468,N_891);
nor U12457 (N_12457,N_2838,N_73);
nor U12458 (N_12458,N_6222,N_6356);
nor U12459 (N_12459,N_1237,N_5042);
nand U12460 (N_12460,N_1820,N_3323);
nand U12461 (N_12461,N_482,N_3400);
or U12462 (N_12462,N_3888,N_1632);
and U12463 (N_12463,N_5316,N_8412);
and U12464 (N_12464,N_4315,N_5071);
nor U12465 (N_12465,N_5463,N_1339);
nand U12466 (N_12466,N_4421,N_9237);
nor U12467 (N_12467,N_4841,N_1579);
and U12468 (N_12468,N_9642,N_4364);
and U12469 (N_12469,N_7462,N_8480);
nor U12470 (N_12470,N_4036,N_3551);
nand U12471 (N_12471,N_2160,N_807);
nand U12472 (N_12472,N_4869,N_913);
xnor U12473 (N_12473,N_9930,N_4381);
xor U12474 (N_12474,N_7153,N_2677);
and U12475 (N_12475,N_7180,N_6845);
and U12476 (N_12476,N_8333,N_9738);
nand U12477 (N_12477,N_3612,N_5444);
nor U12478 (N_12478,N_5203,N_2054);
or U12479 (N_12479,N_617,N_4955);
or U12480 (N_12480,N_6104,N_4777);
and U12481 (N_12481,N_6781,N_219);
and U12482 (N_12482,N_8084,N_6368);
xor U12483 (N_12483,N_8829,N_9850);
xnor U12484 (N_12484,N_8837,N_8355);
nand U12485 (N_12485,N_7279,N_3804);
xor U12486 (N_12486,N_391,N_7121);
xor U12487 (N_12487,N_8132,N_3784);
and U12488 (N_12488,N_7186,N_2036);
or U12489 (N_12489,N_7216,N_5523);
or U12490 (N_12490,N_5974,N_5872);
nand U12491 (N_12491,N_3168,N_6982);
and U12492 (N_12492,N_8497,N_7654);
xnor U12493 (N_12493,N_5539,N_602);
or U12494 (N_12494,N_1509,N_8030);
and U12495 (N_12495,N_1766,N_4977);
and U12496 (N_12496,N_937,N_6252);
nand U12497 (N_12497,N_6715,N_3652);
or U12498 (N_12498,N_918,N_8646);
and U12499 (N_12499,N_3405,N_2495);
or U12500 (N_12500,N_9835,N_1888);
nor U12501 (N_12501,N_4694,N_9227);
nor U12502 (N_12502,N_3337,N_6055);
xnor U12503 (N_12503,N_5959,N_7163);
nor U12504 (N_12504,N_5127,N_6937);
nand U12505 (N_12505,N_1701,N_4481);
and U12506 (N_12506,N_7471,N_8619);
nor U12507 (N_12507,N_3728,N_1245);
xnor U12508 (N_12508,N_4542,N_6199);
nor U12509 (N_12509,N_7677,N_6329);
and U12510 (N_12510,N_7052,N_4709);
nor U12511 (N_12511,N_2898,N_4042);
nor U12512 (N_12512,N_2004,N_5668);
nand U12513 (N_12513,N_2503,N_510);
or U12514 (N_12514,N_7006,N_7520);
nor U12515 (N_12515,N_4780,N_7392);
and U12516 (N_12516,N_9757,N_9633);
nor U12517 (N_12517,N_4567,N_1930);
nor U12518 (N_12518,N_1179,N_9926);
xor U12519 (N_12519,N_8474,N_7201);
nor U12520 (N_12520,N_6384,N_5906);
nor U12521 (N_12521,N_6166,N_7806);
xor U12522 (N_12522,N_6940,N_5504);
or U12523 (N_12523,N_6654,N_8950);
or U12524 (N_12524,N_9327,N_5630);
or U12525 (N_12525,N_8718,N_707);
nand U12526 (N_12526,N_3436,N_4303);
or U12527 (N_12527,N_1453,N_4164);
xnor U12528 (N_12528,N_4250,N_7248);
nand U12529 (N_12529,N_5013,N_4538);
xnor U12530 (N_12530,N_8985,N_6294);
nor U12531 (N_12531,N_2156,N_5520);
or U12532 (N_12532,N_2837,N_8755);
and U12533 (N_12533,N_2330,N_7330);
or U12534 (N_12534,N_1646,N_6318);
or U12535 (N_12535,N_3210,N_341);
or U12536 (N_12536,N_8620,N_4576);
nand U12537 (N_12537,N_7051,N_607);
and U12538 (N_12538,N_2019,N_8995);
nand U12539 (N_12539,N_4249,N_2280);
nand U12540 (N_12540,N_4889,N_6817);
xor U12541 (N_12541,N_1328,N_6674);
and U12542 (N_12542,N_9578,N_2114);
nor U12543 (N_12543,N_9577,N_2351);
nor U12544 (N_12544,N_3172,N_7418);
xor U12545 (N_12545,N_2209,N_4980);
nand U12546 (N_12546,N_6498,N_986);
nand U12547 (N_12547,N_4499,N_3352);
and U12548 (N_12548,N_1920,N_832);
and U12549 (N_12549,N_1450,N_2783);
nand U12550 (N_12550,N_2733,N_7631);
or U12551 (N_12551,N_2614,N_5532);
xor U12552 (N_12552,N_7719,N_8472);
nand U12553 (N_12553,N_7189,N_1648);
nand U12554 (N_12554,N_3431,N_2401);
xnor U12555 (N_12555,N_1290,N_2041);
nand U12556 (N_12556,N_4843,N_5714);
or U12557 (N_12557,N_4305,N_8545);
nor U12558 (N_12558,N_5871,N_8819);
nand U12559 (N_12559,N_6213,N_773);
xor U12560 (N_12560,N_7663,N_6547);
and U12561 (N_12561,N_5237,N_1458);
and U12562 (N_12562,N_676,N_1874);
nand U12563 (N_12563,N_5695,N_7722);
or U12564 (N_12564,N_4275,N_4206);
nor U12565 (N_12565,N_9639,N_1215);
nand U12566 (N_12566,N_4740,N_1121);
nand U12567 (N_12567,N_5379,N_6317);
nor U12568 (N_12568,N_396,N_2987);
xnor U12569 (N_12569,N_6474,N_9512);
nand U12570 (N_12570,N_868,N_2933);
nor U12571 (N_12571,N_8059,N_339);
and U12572 (N_12572,N_1360,N_8051);
nand U12573 (N_12573,N_2290,N_3625);
or U12574 (N_12574,N_4814,N_4685);
nand U12575 (N_12575,N_6589,N_998);
nand U12576 (N_12576,N_6951,N_7041);
and U12577 (N_12577,N_1208,N_2564);
nor U12578 (N_12578,N_1274,N_4618);
or U12579 (N_12579,N_9654,N_2707);
and U12580 (N_12580,N_7143,N_8470);
and U12581 (N_12581,N_1228,N_8827);
nor U12582 (N_12582,N_4091,N_1111);
nor U12583 (N_12583,N_8866,N_8305);
nor U12584 (N_12584,N_1776,N_586);
or U12585 (N_12585,N_2740,N_4097);
and U12586 (N_12586,N_9472,N_1710);
xnor U12587 (N_12587,N_2125,N_4427);
nand U12588 (N_12588,N_9667,N_7928);
or U12589 (N_12589,N_2239,N_7113);
xor U12590 (N_12590,N_8708,N_1791);
nand U12591 (N_12591,N_749,N_4218);
xnor U12592 (N_12592,N_2970,N_842);
nor U12593 (N_12593,N_6100,N_7514);
nand U12594 (N_12594,N_5642,N_1185);
nor U12595 (N_12595,N_6691,N_4494);
nor U12596 (N_12596,N_8851,N_6518);
or U12597 (N_12597,N_5049,N_1255);
nand U12598 (N_12598,N_4253,N_323);
and U12599 (N_12599,N_9399,N_7095);
or U12600 (N_12600,N_5544,N_8964);
nor U12601 (N_12601,N_3798,N_1426);
xnor U12602 (N_12602,N_3334,N_6405);
or U12603 (N_12603,N_6777,N_3288);
nand U12604 (N_12604,N_7710,N_9830);
nand U12605 (N_12605,N_1178,N_4651);
or U12606 (N_12606,N_3102,N_5534);
or U12607 (N_12607,N_4038,N_781);
xnor U12608 (N_12608,N_2377,N_3029);
nor U12609 (N_12609,N_2215,N_5716);
nand U12610 (N_12610,N_9941,N_4198);
or U12611 (N_12611,N_2203,N_6553);
xor U12612 (N_12612,N_8399,N_191);
and U12613 (N_12613,N_2739,N_2573);
nand U12614 (N_12614,N_6618,N_1266);
nand U12615 (N_12615,N_6141,N_938);
and U12616 (N_12616,N_532,N_9913);
nand U12617 (N_12617,N_8139,N_4635);
nand U12618 (N_12618,N_1461,N_599);
nor U12619 (N_12619,N_6418,N_6324);
nand U12620 (N_12620,N_3147,N_7874);
nand U12621 (N_12621,N_6249,N_1897);
nor U12622 (N_12622,N_3426,N_9501);
nor U12623 (N_12623,N_1216,N_6071);
xor U12624 (N_12624,N_7655,N_2380);
nor U12625 (N_12625,N_1759,N_9416);
xor U12626 (N_12626,N_896,N_4925);
or U12627 (N_12627,N_5122,N_8121);
nand U12628 (N_12628,N_1542,N_1838);
xnor U12629 (N_12629,N_7961,N_1142);
nor U12630 (N_12630,N_3855,N_7424);
or U12631 (N_12631,N_951,N_4991);
nor U12632 (N_12632,N_3131,N_5800);
and U12633 (N_12633,N_1006,N_7482);
or U12634 (N_12634,N_8430,N_4861);
xnor U12635 (N_12635,N_3341,N_3016);
xor U12636 (N_12636,N_8751,N_8559);
and U12637 (N_12637,N_2553,N_2964);
xnor U12638 (N_12638,N_7285,N_5582);
xor U12639 (N_12639,N_6939,N_5111);
and U12640 (N_12640,N_9566,N_7510);
nor U12641 (N_12641,N_67,N_4082);
and U12642 (N_12642,N_6989,N_1330);
xnor U12643 (N_12643,N_3343,N_8910);
nand U12644 (N_12644,N_9777,N_7742);
nand U12645 (N_12645,N_2704,N_761);
xor U12646 (N_12646,N_7812,N_8616);
xnor U12647 (N_12647,N_394,N_5984);
xnor U12648 (N_12648,N_9650,N_1160);
nor U12649 (N_12649,N_8428,N_4329);
nand U12650 (N_12650,N_2935,N_6751);
nor U12651 (N_12651,N_1207,N_8825);
xor U12652 (N_12652,N_7533,N_1246);
nand U12653 (N_12653,N_8442,N_9640);
nand U12654 (N_12654,N_1367,N_1945);
and U12655 (N_12655,N_3633,N_987);
xnor U12656 (N_12656,N_3319,N_8328);
nand U12657 (N_12657,N_4734,N_2396);
or U12658 (N_12658,N_6838,N_2230);
nand U12659 (N_12659,N_4151,N_5120);
nor U12660 (N_12660,N_8268,N_6679);
nand U12661 (N_12661,N_9779,N_4724);
nand U12662 (N_12662,N_9347,N_4771);
or U12663 (N_12663,N_8295,N_4013);
nor U12664 (N_12664,N_252,N_3941);
xor U12665 (N_12665,N_6373,N_9743);
or U12666 (N_12666,N_4294,N_4118);
or U12667 (N_12667,N_3229,N_6083);
nand U12668 (N_12668,N_9478,N_8709);
xor U12669 (N_12669,N_5083,N_5006);
xor U12670 (N_12670,N_1879,N_9860);
and U12671 (N_12671,N_6201,N_9474);
nor U12672 (N_12672,N_2319,N_7771);
nand U12673 (N_12673,N_491,N_6261);
xnor U12674 (N_12674,N_5207,N_3763);
nor U12675 (N_12675,N_5573,N_9213);
nor U12676 (N_12676,N_1197,N_8072);
or U12677 (N_12677,N_85,N_7883);
and U12678 (N_12678,N_6794,N_8108);
nand U12679 (N_12679,N_1361,N_8527);
nor U12680 (N_12680,N_7037,N_7490);
nand U12681 (N_12681,N_455,N_5580);
nand U12682 (N_12682,N_6448,N_2164);
nor U12683 (N_12683,N_7173,N_7944);
xnor U12684 (N_12684,N_993,N_1661);
and U12685 (N_12685,N_553,N_4289);
xnor U12686 (N_12686,N_2761,N_6695);
xor U12687 (N_12687,N_8647,N_5883);
or U12688 (N_12688,N_6584,N_5322);
nand U12689 (N_12689,N_1687,N_3373);
nand U12690 (N_12690,N_2574,N_3398);
or U12691 (N_12691,N_930,N_1782);
xor U12692 (N_12692,N_3013,N_6434);
xnor U12693 (N_12693,N_8152,N_9312);
nand U12694 (N_12694,N_5836,N_9741);
or U12695 (N_12695,N_6632,N_5027);
or U12696 (N_12696,N_2764,N_8696);
xor U12697 (N_12697,N_8912,N_1345);
nand U12698 (N_12698,N_1566,N_5128);
nor U12699 (N_12699,N_698,N_3293);
and U12700 (N_12700,N_6602,N_1936);
nor U12701 (N_12701,N_7665,N_4480);
nor U12702 (N_12702,N_4238,N_5342);
or U12703 (N_12703,N_2371,N_7151);
xnor U12704 (N_12704,N_5276,N_1200);
xnor U12705 (N_12705,N_4887,N_7394);
and U12706 (N_12706,N_7363,N_5778);
xnor U12707 (N_12707,N_1671,N_7760);
nor U12708 (N_12708,N_2105,N_3588);
xnor U12709 (N_12709,N_6860,N_8269);
xnor U12710 (N_12710,N_7056,N_4517);
nand U12711 (N_12711,N_8590,N_1180);
xor U12712 (N_12712,N_9760,N_254);
xor U12713 (N_12713,N_4395,N_2409);
nor U12714 (N_12714,N_3050,N_3199);
xnor U12715 (N_12715,N_8264,N_626);
xnor U12716 (N_12716,N_2920,N_1957);
nand U12717 (N_12717,N_5558,N_6477);
xnor U12718 (N_12718,N_3808,N_203);
nand U12719 (N_12719,N_7905,N_4021);
and U12720 (N_12720,N_3065,N_2787);
nor U12721 (N_12721,N_8512,N_5208);
and U12722 (N_12722,N_7829,N_8195);
nand U12723 (N_12723,N_6640,N_8032);
xnor U12724 (N_12724,N_8994,N_4930);
nor U12725 (N_12725,N_3841,N_2100);
nor U12726 (N_12726,N_9579,N_5471);
nor U12727 (N_12727,N_5952,N_9190);
and U12728 (N_12728,N_3953,N_2138);
or U12729 (N_12729,N_8156,N_7716);
and U12730 (N_12730,N_4001,N_1808);
xnor U12731 (N_12731,N_2650,N_9186);
and U12732 (N_12732,N_7616,N_9672);
or U12733 (N_12733,N_5525,N_3554);
and U12734 (N_12734,N_3864,N_4512);
nand U12735 (N_12735,N_3624,N_8843);
nor U12736 (N_12736,N_8069,N_1729);
nand U12737 (N_12737,N_1713,N_8903);
nand U12738 (N_12738,N_7941,N_4225);
nor U12739 (N_12739,N_8240,N_3510);
nand U12740 (N_12740,N_6971,N_7222);
nor U12741 (N_12741,N_7172,N_5048);
and U12742 (N_12742,N_3584,N_2263);
and U12743 (N_12743,N_9195,N_9346);
or U12744 (N_12744,N_5581,N_48);
nand U12745 (N_12745,N_425,N_8864);
xnor U12746 (N_12746,N_2991,N_9946);
nand U12747 (N_12747,N_1063,N_133);
nor U12748 (N_12748,N_7289,N_6979);
or U12749 (N_12749,N_6949,N_4929);
and U12750 (N_12750,N_5154,N_8071);
xnor U12751 (N_12751,N_5791,N_2994);
and U12752 (N_12752,N_1609,N_2181);
nor U12753 (N_12753,N_8605,N_2526);
xor U12754 (N_12754,N_8115,N_3542);
nand U12755 (N_12755,N_5877,N_7832);
nand U12756 (N_12756,N_8262,N_7454);
and U12757 (N_12757,N_4322,N_8514);
nor U12758 (N_12758,N_4156,N_104);
and U12759 (N_12759,N_7898,N_3886);
or U12760 (N_12760,N_5673,N_3747);
or U12761 (N_12761,N_4762,N_6126);
xnor U12762 (N_12762,N_2104,N_8347);
or U12763 (N_12763,N_2836,N_7709);
or U12764 (N_12764,N_1765,N_7453);
or U12765 (N_12765,N_1384,N_1419);
nand U12766 (N_12766,N_4308,N_4450);
nand U12767 (N_12767,N_2984,N_8272);
and U12768 (N_12768,N_8598,N_6705);
nand U12769 (N_12769,N_6738,N_2332);
nor U12770 (N_12770,N_2647,N_7442);
or U12771 (N_12771,N_6713,N_5140);
nor U12772 (N_12772,N_8962,N_674);
nor U12773 (N_12773,N_2554,N_6377);
or U12774 (N_12774,N_2218,N_4826);
or U12775 (N_12775,N_6280,N_794);
xor U12776 (N_12776,N_6026,N_4093);
nand U12777 (N_12777,N_173,N_530);
nor U12778 (N_12778,N_9722,N_5575);
xor U12779 (N_12779,N_6818,N_6292);
nor U12780 (N_12780,N_7260,N_5328);
and U12781 (N_12781,N_165,N_686);
or U12782 (N_12782,N_5038,N_5850);
nand U12783 (N_12783,N_8172,N_1195);
nor U12784 (N_12784,N_4433,N_4266);
and U12785 (N_12785,N_8124,N_8005);
or U12786 (N_12786,N_3959,N_5366);
and U12787 (N_12787,N_5397,N_8456);
nor U12788 (N_12788,N_5767,N_5545);
and U12789 (N_12789,N_1260,N_1471);
xnor U12790 (N_12790,N_3019,N_235);
or U12791 (N_12791,N_9696,N_2738);
xor U12792 (N_12792,N_6094,N_4028);
xor U12793 (N_12793,N_1113,N_4122);
or U12794 (N_12794,N_9762,N_3385);
xnor U12795 (N_12795,N_4219,N_8335);
xnor U12796 (N_12796,N_8676,N_3061);
nor U12797 (N_12797,N_5321,N_4609);
nand U12798 (N_12798,N_7110,N_810);
nand U12799 (N_12799,N_864,N_1942);
or U12800 (N_12800,N_248,N_3090);
nand U12801 (N_12801,N_9273,N_9194);
xor U12802 (N_12802,N_6598,N_4803);
or U12803 (N_12803,N_313,N_4483);
nor U12804 (N_12804,N_7977,N_2942);
and U12805 (N_12805,N_139,N_3401);
and U12806 (N_12806,N_661,N_2106);
xor U12807 (N_12807,N_452,N_5016);
xnor U12808 (N_12808,N_7723,N_8427);
and U12809 (N_12809,N_2270,N_2408);
or U12810 (N_12810,N_3257,N_1900);
nand U12811 (N_12811,N_7364,N_3653);
xor U12812 (N_12812,N_4025,N_9635);
xor U12813 (N_12813,N_9026,N_7745);
nor U12814 (N_12814,N_557,N_3214);
and U12815 (N_12815,N_7438,N_5294);
and U12816 (N_12816,N_5184,N_8443);
or U12817 (N_12817,N_6086,N_9412);
xnor U12818 (N_12818,N_6254,N_4123);
xnor U12819 (N_12819,N_6311,N_2570);
or U12820 (N_12820,N_9378,N_5893);
or U12821 (N_12821,N_6459,N_9543);
nor U12822 (N_12822,N_1029,N_167);
and U12823 (N_12823,N_2775,N_2119);
xnor U12824 (N_12824,N_8275,N_865);
nand U12825 (N_12825,N_2474,N_6352);
and U12826 (N_12826,N_5340,N_5261);
and U12827 (N_12827,N_4528,N_3852);
xor U12828 (N_12828,N_3036,N_8203);
nor U12829 (N_12829,N_161,N_9206);
nor U12830 (N_12830,N_7630,N_7472);
xor U12831 (N_12831,N_3636,N_6677);
nand U12832 (N_12832,N_2899,N_5489);
nor U12833 (N_12833,N_2144,N_5179);
nand U12834 (N_12834,N_2501,N_7615);
or U12835 (N_12835,N_5329,N_5124);
or U12836 (N_12836,N_8863,N_1381);
xor U12837 (N_12837,N_4060,N_9475);
and U12838 (N_12838,N_3746,N_4769);
xnor U12839 (N_12839,N_3922,N_9945);
nand U12840 (N_12840,N_566,N_1090);
or U12841 (N_12841,N_2347,N_8503);
xnor U12842 (N_12842,N_2593,N_2651);
nand U12843 (N_12843,N_885,N_9119);
xnor U12844 (N_12844,N_6724,N_9164);
nand U12845 (N_12845,N_7474,N_6303);
nor U12846 (N_12846,N_8277,N_6480);
nor U12847 (N_12847,N_4137,N_6880);
xor U12848 (N_12848,N_7724,N_8918);
or U12849 (N_12849,N_8475,N_8867);
and U12850 (N_12850,N_7680,N_8267);
nand U12851 (N_12851,N_66,N_4120);
or U12852 (N_12852,N_9864,N_2706);
and U12853 (N_12853,N_2613,N_2918);
nand U12854 (N_12854,N_1907,N_8963);
nor U12855 (N_12855,N_4299,N_4811);
nand U12856 (N_12856,N_3801,N_5530);
nor U12857 (N_12857,N_272,N_731);
and U12858 (N_12858,N_7989,N_8793);
nor U12859 (N_12859,N_2266,N_4167);
and U12860 (N_12860,N_2556,N_9005);
nor U12861 (N_12861,N_3890,N_4664);
xnor U12862 (N_12862,N_103,N_8357);
nand U12863 (N_12863,N_1238,N_424);
nor U12864 (N_12864,N_9121,N_8660);
and U12865 (N_12865,N_7346,N_4670);
or U12866 (N_12866,N_5647,N_7999);
nand U12867 (N_12867,N_1869,N_5991);
nand U12868 (N_12868,N_8109,N_8070);
nand U12869 (N_12869,N_8612,N_777);
xnor U12870 (N_12870,N_3217,N_1938);
nand U12871 (N_12871,N_9210,N_4343);
nand U12872 (N_12872,N_7820,N_3262);
nor U12873 (N_12873,N_6746,N_9800);
or U12874 (N_12874,N_1248,N_9649);
nand U12875 (N_12875,N_6404,N_7769);
nand U12876 (N_12876,N_2492,N_669);
or U12877 (N_12877,N_9176,N_5648);
and U12878 (N_12878,N_1704,N_7111);
and U12879 (N_12879,N_2500,N_5041);
or U12880 (N_12880,N_4425,N_8207);
or U12881 (N_12881,N_7070,N_8205);
nor U12882 (N_12882,N_158,N_6897);
xor U12883 (N_12883,N_8153,N_5697);
nand U12884 (N_12884,N_6953,N_7038);
and U12885 (N_12885,N_6819,N_2844);
xnor U12886 (N_12886,N_2771,N_8858);
and U12887 (N_12887,N_2749,N_1143);
nor U12888 (N_12888,N_4290,N_8822);
and U12889 (N_12889,N_540,N_8956);
nand U12890 (N_12890,N_6259,N_9409);
nor U12891 (N_12891,N_6807,N_200);
nand U12892 (N_12892,N_816,N_6784);
nor U12893 (N_12893,N_115,N_6987);
nand U12894 (N_12894,N_529,N_4302);
nand U12895 (N_12895,N_4363,N_96);
or U12896 (N_12896,N_6616,N_1909);
and U12897 (N_12897,N_8022,N_8097);
or U12898 (N_12898,N_4217,N_5726);
nor U12899 (N_12899,N_9083,N_7207);
or U12900 (N_12900,N_4133,N_9233);
or U12901 (N_12901,N_4440,N_9972);
and U12902 (N_12902,N_5245,N_7551);
nand U12903 (N_12903,N_8008,N_964);
xnor U12904 (N_12904,N_5939,N_9382);
and U12905 (N_12905,N_8761,N_4098);
and U12906 (N_12906,N_4468,N_8792);
nand U12907 (N_12907,N_6088,N_3667);
nand U12908 (N_12908,N_9125,N_7881);
xor U12909 (N_12909,N_8884,N_7277);
nor U12910 (N_12910,N_1236,N_7092);
and U12911 (N_12911,N_1846,N_929);
nand U12912 (N_12912,N_3952,N_9598);
xnor U12913 (N_12913,N_8159,N_3894);
xor U12914 (N_12914,N_212,N_6263);
nor U12915 (N_12915,N_630,N_2210);
xnor U12916 (N_12916,N_8674,N_1363);
nor U12917 (N_12917,N_4684,N_7247);
xnor U12918 (N_12918,N_3768,N_2057);
xnor U12919 (N_12919,N_6788,N_6135);
xor U12920 (N_12920,N_79,N_1973);
nor U12921 (N_12921,N_3664,N_4128);
xor U12922 (N_12922,N_850,N_9039);
or U12923 (N_12923,N_6188,N_1719);
or U12924 (N_12924,N_101,N_5825);
and U12925 (N_12925,N_5229,N_5533);
xnor U12926 (N_12926,N_862,N_4874);
or U12927 (N_12927,N_8296,N_7557);
and U12928 (N_12928,N_4521,N_6930);
or U12929 (N_12929,N_4463,N_7537);
and U12930 (N_12930,N_3930,N_1708);
and U12931 (N_12931,N_7743,N_6108);
or U12932 (N_12932,N_5253,N_4259);
nand U12933 (N_12933,N_2237,N_7089);
nor U12934 (N_12934,N_5181,N_8983);
xor U12935 (N_12935,N_137,N_4654);
and U12936 (N_12936,N_8515,N_4933);
xor U12937 (N_12937,N_3374,N_3040);
xnor U12938 (N_12938,N_2938,N_3980);
xor U12939 (N_12939,N_8716,N_5384);
or U12940 (N_12940,N_8356,N_8922);
xnor U12941 (N_12941,N_309,N_7572);
and U12942 (N_12942,N_1827,N_6575);
or U12943 (N_12943,N_559,N_1931);
and U12944 (N_12944,N_8094,N_6958);
xor U12945 (N_12945,N_5908,N_5635);
or U12946 (N_12946,N_550,N_6445);
nor U12947 (N_12947,N_3967,N_4878);
or U12948 (N_12948,N_8009,N_7421);
and U12949 (N_12949,N_4172,N_6709);
and U12950 (N_12950,N_9530,N_6903);
and U12951 (N_12951,N_5604,N_5568);
or U12952 (N_12952,N_4681,N_4756);
xnor U12953 (N_12953,N_4775,N_7144);
nand U12954 (N_12954,N_1199,N_7876);
or U12955 (N_12955,N_6882,N_5698);
and U12956 (N_12956,N_1184,N_2887);
and U12957 (N_12957,N_215,N_8056);
and U12958 (N_12958,N_5882,N_3668);
nor U12959 (N_12959,N_1651,N_8542);
or U12960 (N_12960,N_8033,N_1627);
nor U12961 (N_12961,N_9724,N_8543);
nor U12962 (N_12962,N_3552,N_5201);
or U12963 (N_12963,N_6064,N_1954);
nand U12964 (N_12964,N_5206,N_7132);
xnor U12965 (N_12965,N_3062,N_2487);
nor U12966 (N_12966,N_7872,N_462);
xnor U12967 (N_12967,N_2822,N_4976);
or U12968 (N_12968,N_9794,N_1481);
nor U12969 (N_12969,N_9248,N_1078);
and U12970 (N_12970,N_2220,N_3978);
xor U12971 (N_12971,N_5007,N_3201);
and U12972 (N_12972,N_4389,N_5238);
nor U12973 (N_12973,N_2547,N_7821);
nor U12974 (N_12974,N_1412,N_3153);
nor U12975 (N_12975,N_1159,N_7588);
and U12976 (N_12976,N_1959,N_5804);
and U12977 (N_12977,N_2861,N_5414);
or U12978 (N_12978,N_2342,N_1662);
xor U12979 (N_12979,N_814,N_8168);
and U12980 (N_12980,N_9785,N_6327);
nand U12981 (N_12981,N_2561,N_9395);
and U12982 (N_12982,N_691,N_560);
nand U12983 (N_12983,N_5251,N_2140);
nand U12984 (N_12984,N_9754,N_1599);
nor U12985 (N_12985,N_2000,N_7103);
and U12986 (N_12986,N_7383,N_6076);
nand U12987 (N_12987,N_2213,N_8406);
nand U12988 (N_12988,N_1523,N_8459);
and U12989 (N_12989,N_2847,N_8483);
or U12990 (N_12990,N_7196,N_7317);
or U12991 (N_12991,N_2390,N_7559);
nand U12992 (N_12992,N_4942,N_7255);
nor U12993 (N_12993,N_8658,N_87);
xnor U12994 (N_12994,N_6433,N_6208);
and U12995 (N_12995,N_7638,N_8300);
and U12996 (N_12996,N_5495,N_4424);
nand U12997 (N_12997,N_1196,N_9343);
nor U12998 (N_12998,N_2934,N_2260);
nor U12999 (N_12999,N_2863,N_6780);
xnor U13000 (N_13000,N_2768,N_9212);
nand U13001 (N_13001,N_8955,N_9518);
xnor U13002 (N_13002,N_9752,N_4822);
xnor U13003 (N_13003,N_31,N_2720);
xor U13004 (N_13004,N_5935,N_8519);
and U13005 (N_13005,N_3480,N_2638);
xnor U13006 (N_13006,N_8247,N_1321);
and U13007 (N_13007,N_5978,N_523);
or U13008 (N_13008,N_3806,N_9124);
or U13009 (N_13009,N_5728,N_4537);
and U13010 (N_13010,N_6894,N_1291);
or U13011 (N_13011,N_1955,N_6573);
nor U13012 (N_13012,N_3184,N_4732);
xor U13013 (N_13013,N_3368,N_1251);
or U13014 (N_13014,N_3377,N_1428);
or U13015 (N_13015,N_8721,N_7370);
nand U13016 (N_13016,N_310,N_4031);
nand U13017 (N_13017,N_8940,N_2232);
or U13018 (N_13018,N_6658,N_8522);
or U13019 (N_13019,N_1529,N_1375);
or U13020 (N_13020,N_1065,N_5019);
nand U13021 (N_13021,N_8703,N_154);
nand U13022 (N_13022,N_6401,N_664);
nor U13023 (N_13023,N_5275,N_1288);
xnor U13024 (N_13024,N_4444,N_5265);
and U13025 (N_13025,N_6151,N_3777);
xnor U13026 (N_13026,N_2618,N_7669);
xnor U13027 (N_13027,N_5729,N_7544);
xnor U13028 (N_13028,N_1089,N_8584);
xnor U13029 (N_13029,N_2540,N_555);
nor U13030 (N_13030,N_7386,N_1691);
nor U13031 (N_13031,N_4675,N_2958);
nand U13032 (N_13032,N_2245,N_114);
or U13033 (N_13033,N_6926,N_1762);
nand U13034 (N_13034,N_3954,N_2518);
nand U13035 (N_13035,N_3504,N_753);
nand U13036 (N_13036,N_5627,N_2379);
and U13037 (N_13037,N_1378,N_1365);
xor U13038 (N_13038,N_6172,N_1705);
and U13039 (N_13039,N_4765,N_3971);
and U13040 (N_13040,N_6229,N_6171);
xor U13041 (N_13041,N_3038,N_2282);
nand U13042 (N_13042,N_9075,N_4384);
or U13043 (N_13043,N_9623,N_6920);
or U13044 (N_13044,N_9539,N_6797);
and U13045 (N_13045,N_5069,N_7106);
or U13046 (N_13046,N_8106,N_7681);
nand U13047 (N_13047,N_5055,N_1821);
xnor U13048 (N_13048,N_2794,N_1017);
and U13049 (N_13049,N_25,N_5368);
or U13050 (N_13050,N_3790,N_9054);
xnor U13051 (N_13051,N_7429,N_224);
and U13052 (N_13052,N_9196,N_9628);
nand U13053 (N_13053,N_7670,N_1198);
and U13054 (N_13054,N_6006,N_5190);
or U13055 (N_13055,N_9394,N_4858);
or U13056 (N_13056,N_6717,N_8552);
and U13057 (N_13057,N_5571,N_9116);
or U13058 (N_13058,N_3058,N_3744);
or U13059 (N_13059,N_1374,N_9708);
or U13060 (N_13060,N_8707,N_5816);
xnor U13061 (N_13061,N_6120,N_9906);
nand U13062 (N_13062,N_1366,N_1235);
nand U13063 (N_13063,N_863,N_1405);
and U13064 (N_13064,N_4835,N_9380);
and U13065 (N_13065,N_7419,N_7591);
nor U13066 (N_13066,N_2064,N_8602);
or U13067 (N_13067,N_9316,N_9933);
xnor U13068 (N_13068,N_3326,N_8534);
and U13069 (N_13069,N_9560,N_59);
nor U13070 (N_13070,N_9058,N_6805);
nand U13071 (N_13071,N_3330,N_7495);
or U13072 (N_13072,N_579,N_2040);
nand U13073 (N_13073,N_1318,N_8925);
or U13074 (N_13074,N_8641,N_9636);
and U13075 (N_13075,N_3280,N_8063);
nor U13076 (N_13076,N_6905,N_9651);
or U13077 (N_13077,N_1267,N_3463);
xor U13078 (N_13078,N_8648,N_945);
nand U13079 (N_13079,N_2338,N_2142);
or U13080 (N_13080,N_2652,N_8479);
nor U13081 (N_13081,N_2261,N_6358);
and U13082 (N_13082,N_1659,N_6692);
xnor U13083 (N_13083,N_2481,N_577);
and U13084 (N_13084,N_123,N_940);
and U13085 (N_13085,N_414,N_2676);
or U13086 (N_13086,N_6929,N_2912);
xnor U13087 (N_13087,N_3851,N_562);
nor U13088 (N_13088,N_9725,N_3563);
xnor U13089 (N_13089,N_3906,N_202);
or U13090 (N_13090,N_3315,N_1007);
xnor U13091 (N_13091,N_8212,N_6214);
and U13092 (N_13092,N_7937,N_5787);
xnor U13093 (N_13093,N_8585,N_714);
or U13094 (N_13094,N_7573,N_9081);
xor U13095 (N_13095,N_2622,N_9199);
and U13096 (N_13096,N_9341,N_8949);
xnor U13097 (N_13097,N_1568,N_8796);
xnor U13098 (N_13098,N_5637,N_4530);
and U13099 (N_13099,N_3939,N_3466);
and U13100 (N_13100,N_4049,N_6748);
and U13101 (N_13101,N_8371,N_3853);
nor U13102 (N_13102,N_5358,N_2678);
nand U13103 (N_13103,N_8880,N_5352);
or U13104 (N_13104,N_6585,N_4643);
xor U13105 (N_13105,N_3628,N_8731);
and U13106 (N_13106,N_5958,N_2858);
nand U13107 (N_13107,N_600,N_5221);
or U13108 (N_13108,N_6024,N_1634);
nor U13109 (N_13109,N_9032,N_1264);
or U13110 (N_13110,N_372,N_8073);
and U13111 (N_13111,N_1880,N_9868);
nand U13112 (N_13112,N_7028,N_5086);
nand U13113 (N_13113,N_2463,N_9449);
xnor U13114 (N_13114,N_5032,N_8372);
nor U13115 (N_13115,N_2778,N_2598);
nor U13116 (N_13116,N_6959,N_8784);
or U13117 (N_13117,N_1390,N_106);
nand U13118 (N_13118,N_7124,N_8933);
nor U13119 (N_13119,N_9662,N_4617);
or U13120 (N_13120,N_9397,N_413);
and U13121 (N_13121,N_806,N_7221);
nand U13122 (N_13122,N_1008,N_8146);
nor U13123 (N_13123,N_6290,N_108);
or U13124 (N_13124,N_7377,N_428);
or U13125 (N_13125,N_5937,N_7059);
and U13126 (N_13126,N_995,N_7142);
nand U13127 (N_13127,N_487,N_788);
or U13128 (N_13128,N_8701,N_9614);
and U13129 (N_13129,N_3732,N_6986);
or U13130 (N_13130,N_6753,N_8556);
nand U13131 (N_13131,N_4408,N_5881);
or U13132 (N_13132,N_5046,N_8258);
and U13133 (N_13133,N_1795,N_6795);
or U13134 (N_13134,N_8025,N_894);
xnor U13135 (N_13135,N_6773,N_8284);
nor U13136 (N_13136,N_4476,N_897);
nand U13137 (N_13137,N_6864,N_3710);
nor U13138 (N_13138,N_8779,N_9400);
nand U13139 (N_13139,N_4544,N_7860);
or U13140 (N_13140,N_5110,N_4673);
xnor U13141 (N_13141,N_2885,N_7733);
nor U13142 (N_13142,N_211,N_2980);
or U13143 (N_13143,N_3416,N_8433);
and U13144 (N_13144,N_9993,N_3755);
or U13145 (N_13145,N_580,N_8705);
nor U13146 (N_13146,N_5933,N_1124);
xor U13147 (N_13147,N_6706,N_3324);
xor U13148 (N_13148,N_4588,N_5043);
and U13149 (N_13149,N_5416,N_2683);
nand U13150 (N_13150,N_2047,N_5303);
xor U13151 (N_13151,N_22,N_4017);
nand U13152 (N_13152,N_2076,N_1172);
nand U13153 (N_13153,N_5222,N_9573);
and U13154 (N_13154,N_3180,N_7353);
nor U13155 (N_13155,N_3099,N_631);
nor U13156 (N_13156,N_4184,N_9773);
xnor U13157 (N_13157,N_6113,N_9866);
xnor U13158 (N_13158,N_8104,N_5863);
or U13159 (N_13159,N_6299,N_9200);
nand U13160 (N_13160,N_1926,N_8895);
nor U13161 (N_13161,N_7705,N_3241);
nor U13162 (N_13162,N_6571,N_8473);
nand U13163 (N_13163,N_9146,N_5980);
xnor U13164 (N_13164,N_6512,N_2891);
nand U13165 (N_13165,N_8776,N_7228);
nand U13166 (N_13166,N_5011,N_3902);
and U13167 (N_13167,N_3467,N_8365);
nand U13168 (N_13168,N_4383,N_7982);
xnor U13169 (N_13169,N_4581,N_8613);
or U13170 (N_13170,N_3831,N_348);
or U13171 (N_13171,N_9482,N_1010);
nor U13172 (N_13172,N_3125,N_7754);
and U13173 (N_13173,N_7933,N_4178);
or U13174 (N_13174,N_3774,N_8053);
nor U13175 (N_13175,N_5892,N_9113);
and U13176 (N_13176,N_1600,N_1161);
nand U13177 (N_13177,N_5337,N_1639);
or U13178 (N_13178,N_7893,N_3296);
and U13179 (N_13179,N_9339,N_916);
nand U13180 (N_13180,N_9904,N_7251);
or U13181 (N_13181,N_7633,N_7437);
nand U13182 (N_13182,N_7313,N_5675);
or U13183 (N_13183,N_591,N_7209);
nand U13184 (N_13184,N_849,N_2637);
or U13185 (N_13185,N_3656,N_6834);
nor U13186 (N_13186,N_3304,N_1830);
nand U13187 (N_13187,N_9513,N_5002);
and U13188 (N_13188,N_6119,N_1308);
and U13189 (N_13189,N_9625,N_9008);
nand U13190 (N_13190,N_2755,N_498);
xor U13191 (N_13191,N_1130,N_8090);
or U13192 (N_13192,N_7352,N_6867);
and U13193 (N_13193,N_3097,N_6647);
nand U13194 (N_13194,N_4677,N_4744);
and U13195 (N_13195,N_2779,N_7154);
or U13196 (N_13196,N_2785,N_486);
xor U13197 (N_13197,N_4964,N_8856);
xor U13198 (N_13198,N_4152,N_6993);
or U13199 (N_13199,N_6196,N_5957);
xnor U13200 (N_13200,N_8114,N_4348);
or U13201 (N_13201,N_9224,N_1402);
and U13202 (N_13202,N_8558,N_656);
or U13203 (N_13203,N_8873,N_4063);
or U13204 (N_13204,N_6081,N_7149);
xnor U13205 (N_13205,N_1368,N_3781);
and U13206 (N_13206,N_8750,N_2449);
nand U13207 (N_13207,N_384,N_6432);
or U13208 (N_13208,N_2314,N_6823);
and U13209 (N_13209,N_500,N_9713);
nor U13210 (N_13210,N_666,N_552);
nand U13211 (N_13211,N_2243,N_748);
and U13212 (N_13212,N_4104,N_135);
xor U13213 (N_13213,N_9592,N_2567);
and U13214 (N_13214,N_8686,N_9421);
or U13215 (N_13215,N_8342,N_2306);
nand U13216 (N_13216,N_6802,N_2684);
nor U13217 (N_13217,N_9896,N_3081);
xor U13218 (N_13218,N_8980,N_8242);
nor U13219 (N_13219,N_8695,N_227);
or U13220 (N_13220,N_3534,N_6814);
nor U13221 (N_13221,N_6345,N_5426);
and U13222 (N_13222,N_1770,N_1911);
and U13223 (N_13223,N_9398,N_8424);
nand U13224 (N_13224,N_6408,N_1751);
or U13225 (N_13225,N_7213,N_3513);
or U13226 (N_13226,N_6487,N_5896);
nor U13227 (N_13227,N_6403,N_3581);
or U13228 (N_13228,N_531,N_7522);
xnor U13229 (N_13229,N_3331,N_9260);
xnor U13230 (N_13230,N_787,N_2505);
and U13231 (N_13231,N_8986,N_9908);
nor U13232 (N_13232,N_5309,N_7761);
nand U13233 (N_13233,N_2012,N_3592);
nor U13234 (N_13234,N_6883,N_2668);
nand U13235 (N_13235,N_9823,N_9245);
and U13236 (N_13236,N_6656,N_7009);
xor U13237 (N_13237,N_6375,N_1854);
nor U13238 (N_13238,N_8803,N_2834);
nor U13239 (N_13239,N_860,N_3298);
nand U13240 (N_13240,N_9104,N_2328);
nor U13241 (N_13241,N_9646,N_5405);
nand U13242 (N_13242,N_8023,N_780);
nand U13243 (N_13243,N_5543,N_1424);
or U13244 (N_13244,N_3493,N_833);
nand U13245 (N_13245,N_2577,N_3708);
or U13246 (N_13246,N_145,N_612);
xnor U13247 (N_13247,N_7433,N_3702);
nor U13248 (N_13248,N_3327,N_5418);
nand U13249 (N_13249,N_9272,N_8622);
nor U13250 (N_13250,N_1550,N_2605);
nor U13251 (N_13251,N_6831,N_6996);
and U13252 (N_13252,N_5424,N_2065);
and U13253 (N_13253,N_7548,N_3458);
nand U13254 (N_13254,N_1068,N_4432);
nand U13255 (N_13255,N_8632,N_939);
or U13256 (N_13256,N_2769,N_9148);
and U13257 (N_13257,N_7986,N_3770);
nor U13258 (N_13258,N_5866,N_7223);
nor U13259 (N_13259,N_772,N_3522);
nor U13260 (N_13260,N_8711,N_3943);
nand U13261 (N_13261,N_6420,N_4247);
or U13262 (N_13262,N_1152,N_7529);
and U13263 (N_13263,N_9198,N_1594);
nor U13264 (N_13264,N_7469,N_3035);
xor U13265 (N_13265,N_4605,N_6998);
xnor U13266 (N_13266,N_182,N_502);
nand U13267 (N_13267,N_4112,N_6579);
xnor U13268 (N_13268,N_512,N_2452);
nand U13269 (N_13269,N_8906,N_8375);
and U13270 (N_13270,N_2189,N_142);
nor U13271 (N_13271,N_8886,N_230);
nor U13272 (N_13272,N_2339,N_7203);
and U13273 (N_13273,N_3694,N_7934);
nor U13274 (N_13274,N_2469,N_4965);
nor U13275 (N_13275,N_4227,N_2819);
nor U13276 (N_13276,N_4678,N_3919);
nand U13277 (N_13277,N_6865,N_328);
or U13278 (N_13278,N_4264,N_1876);
nand U13279 (N_13279,N_592,N_9716);
and U13280 (N_13280,N_2497,N_6565);
nand U13281 (N_13281,N_1670,N_1515);
xor U13282 (N_13282,N_8336,N_2136);
nand U13283 (N_13283,N_6890,N_811);
nor U13284 (N_13284,N_521,N_518);
xor U13285 (N_13285,N_8973,N_3497);
or U13286 (N_13286,N_9414,N_3446);
xnor U13287 (N_13287,N_4129,N_7417);
or U13288 (N_13288,N_1578,N_8882);
nand U13289 (N_13289,N_5141,N_5312);
or U13290 (N_13290,N_8402,N_9410);
nand U13291 (N_13291,N_1069,N_6275);
and U13292 (N_13292,N_2579,N_9843);
nor U13293 (N_13293,N_9693,N_3236);
and U13294 (N_13294,N_6494,N_1420);
xnor U13295 (N_13295,N_4422,N_7553);
nand U13296 (N_13296,N_876,N_3087);
nand U13297 (N_13297,N_2310,N_2965);
xnor U13298 (N_13298,N_7042,N_7268);
or U13299 (N_13299,N_6875,N_2111);
xnor U13300 (N_13300,N_6269,N_3984);
nor U13301 (N_13301,N_1784,N_5733);
nand U13302 (N_13302,N_8437,N_301);
and U13303 (N_13303,N_6769,N_9525);
nand U13304 (N_13304,N_8631,N_5843);
nand U13305 (N_13305,N_6385,N_2612);
and U13306 (N_13306,N_9541,N_8978);
nor U13307 (N_13307,N_2141,N_5478);
xnor U13308 (N_13308,N_2211,N_1019);
and U13309 (N_13309,N_2267,N_5632);
or U13310 (N_13310,N_7746,N_7046);
xnor U13311 (N_13311,N_3518,N_4546);
nor U13312 (N_13312,N_9753,N_440);
xor U13313 (N_13313,N_4113,N_6173);
or U13314 (N_13314,N_9000,N_5091);
and U13315 (N_13315,N_9825,N_5598);
nor U13316 (N_13316,N_7479,N_3535);
nor U13317 (N_13317,N_2728,N_4070);
and U13318 (N_13318,N_3630,N_2253);
and U13319 (N_13319,N_3651,N_9066);
or U13320 (N_13320,N_2575,N_7840);
or U13321 (N_13321,N_9744,N_2316);
or U13322 (N_13322,N_8038,N_9686);
xor U13323 (N_13323,N_5672,N_7958);
nand U13324 (N_13324,N_6339,N_9064);
xnor U13325 (N_13325,N_8348,N_5380);
and U13326 (N_13326,N_6757,N_5989);
and U13327 (N_13327,N_8083,N_5009);
or U13328 (N_13328,N_9817,N_5066);
or U13329 (N_13329,N_4518,N_2344);
nand U13330 (N_13330,N_2693,N_569);
or U13331 (N_13331,N_4235,N_905);
xor U13332 (N_13332,N_1752,N_7036);
and U13333 (N_13333,N_639,N_5895);
and U13334 (N_13334,N_2853,N_6557);
or U13335 (N_13335,N_8618,N_8836);
nand U13336 (N_13336,N_8461,N_4748);
and U13337 (N_13337,N_943,N_4339);
nand U13338 (N_13338,N_8369,N_5994);
xnor U13339 (N_13339,N_5408,N_4849);
or U13340 (N_13340,N_889,N_4621);
xor U13341 (N_13341,N_9060,N_8099);
xor U13342 (N_13342,N_9249,N_5354);
xor U13343 (N_13343,N_6333,N_5565);
or U13344 (N_13344,N_2667,N_4715);
xnor U13345 (N_13345,N_7768,N_3478);
nand U13346 (N_13346,N_4898,N_9369);
nor U13347 (N_13347,N_4473,N_6884);
and U13348 (N_13348,N_2021,N_6698);
or U13349 (N_13349,N_5143,N_8946);
or U13350 (N_13350,N_6411,N_8374);
nand U13351 (N_13351,N_3567,N_5381);
or U13352 (N_13352,N_3182,N_8788);
xor U13353 (N_13353,N_7910,N_5810);
nand U13354 (N_13354,N_8364,N_9919);
nand U13355 (N_13355,N_7915,N_6899);
nand U13356 (N_13356,N_4044,N_7845);
and U13357 (N_13357,N_2896,N_6218);
or U13358 (N_13358,N_234,N_5995);
nor U13359 (N_13359,N_7312,N_6001);
or U13360 (N_13360,N_6328,N_8444);
and U13361 (N_13361,N_1416,N_8145);
nor U13362 (N_13362,N_6750,N_1754);
and U13363 (N_13363,N_367,N_4094);
nand U13364 (N_13364,N_4626,N_2376);
and U13365 (N_13365,N_4545,N_9988);
xnor U13366 (N_13366,N_7062,N_7693);
nor U13367 (N_13367,N_924,N_8692);
and U13368 (N_13368,N_1177,N_7165);
nand U13369 (N_13369,N_369,N_7627);
nand U13370 (N_13370,N_3154,N_4169);
or U13371 (N_13371,N_1031,N_2324);
or U13372 (N_13372,N_4864,N_218);
nor U13373 (N_13373,N_3022,N_4065);
or U13374 (N_13374,N_9153,N_4524);
xor U13375 (N_13375,N_4124,N_859);
nand U13376 (N_13376,N_1020,N_7193);
nand U13377 (N_13377,N_9219,N_2415);
and U13378 (N_13378,N_7875,N_3203);
nand U13379 (N_13379,N_5466,N_9070);
or U13380 (N_13380,N_3729,N_4595);
and U13381 (N_13381,N_1313,N_5854);
and U13382 (N_13382,N_7938,N_9936);
xor U13383 (N_13383,N_6764,N_6671);
nand U13384 (N_13384,N_770,N_8900);
or U13385 (N_13385,N_6782,N_6343);
xor U13386 (N_13386,N_7637,N_3911);
and U13387 (N_13387,N_9886,N_7484);
nand U13388 (N_13388,N_2249,N_6848);
nand U13389 (N_13389,N_9137,N_5451);
and U13390 (N_13390,N_2095,N_9891);
and U13391 (N_13391,N_9131,N_7350);
or U13392 (N_13392,N_7841,N_466);
nand U13393 (N_13393,N_9015,N_5491);
xor U13394 (N_13394,N_735,N_1018);
and U13395 (N_13395,N_76,N_7439);
and U13396 (N_13396,N_1642,N_4636);
or U13397 (N_13397,N_5639,N_2325);
and U13398 (N_13398,N_9451,N_9493);
nor U13399 (N_13399,N_3124,N_5644);
xor U13400 (N_13400,N_1792,N_7816);
or U13401 (N_13401,N_4316,N_9784);
xor U13402 (N_13402,N_6406,N_8539);
nand U13403 (N_13403,N_3912,N_4475);
nor U13404 (N_13404,N_5477,N_9163);
nand U13405 (N_13405,N_4296,N_4074);
and U13406 (N_13406,N_1656,N_9739);
xnor U13407 (N_13407,N_7576,N_5600);
nor U13408 (N_13408,N_9225,N_6020);
and U13409 (N_13409,N_1072,N_2264);
xnor U13410 (N_13410,N_2516,N_8183);
nor U13411 (N_13411,N_6048,N_117);
and U13412 (N_13412,N_7701,N_1837);
xor U13413 (N_13413,N_2475,N_3834);
nor U13414 (N_13414,N_4393,N_5149);
nand U13415 (N_13415,N_6370,N_26);
or U13416 (N_13416,N_8889,N_2233);
nand U13417 (N_13417,N_7612,N_8027);
nor U13418 (N_13418,N_9938,N_5250);
or U13419 (N_13419,N_2103,N_1071);
xor U13420 (N_13420,N_9950,N_6635);
or U13421 (N_13421,N_9349,N_2480);
or U13422 (N_13422,N_4557,N_3003);
nor U13423 (N_13423,N_4692,N_4326);
and U13424 (N_13424,N_7827,N_1456);
nand U13425 (N_13425,N_5281,N_7804);
nor U13426 (N_13426,N_5021,N_4862);
and U13427 (N_13427,N_2343,N_7232);
nand U13428 (N_13428,N_5249,N_4237);
nand U13429 (N_13429,N_6469,N_5793);
xor U13430 (N_13430,N_9742,N_1254);
xor U13431 (N_13431,N_4330,N_7909);
nand U13432 (N_13432,N_1407,N_6657);
or U13433 (N_13433,N_3295,N_5702);
and U13434 (N_13434,N_5720,N_6626);
xor U13435 (N_13435,N_5453,N_5248);
nor U13436 (N_13436,N_7266,N_7859);
xnor U13437 (N_13437,N_5780,N_8626);
xor U13438 (N_13438,N_2602,N_8265);
xor U13439 (N_13439,N_6189,N_8377);
xnor U13440 (N_13440,N_1972,N_2018);
nor U13441 (N_13441,N_1112,N_6572);
nor U13442 (N_13442,N_6079,N_6551);
or U13443 (N_13443,N_5821,N_8924);
xnor U13444 (N_13444,N_7003,N_5955);
xnor U13445 (N_13445,N_8504,N_9042);
or U13446 (N_13446,N_5434,N_9903);
nor U13447 (N_13447,N_6073,N_1209);
xor U13448 (N_13448,N_3073,N_4023);
nor U13449 (N_13449,N_8440,N_1141);
or U13450 (N_13450,N_6216,N_5262);
and U13451 (N_13451,N_5691,N_259);
or U13452 (N_13452,N_9695,N_6902);
or U13453 (N_13453,N_2659,N_250);
and U13454 (N_13454,N_1174,N_7486);
xor U13455 (N_13455,N_9356,N_909);
nand U13456 (N_13456,N_3069,N_5690);
nand U13457 (N_13457,N_9516,N_9715);
or U13458 (N_13458,N_2429,N_7023);
nand U13459 (N_13459,N_6914,N_8408);
and U13460 (N_13460,N_7340,N_4960);
nor U13461 (N_13461,N_7253,N_7867);
or U13462 (N_13462,N_9458,N_9538);
or U13463 (N_13463,N_352,N_6084);
nor U13464 (N_13464,N_5722,N_4912);
nand U13465 (N_13465,N_6239,N_4598);
xnor U13466 (N_13466,N_8510,N_3361);
and U13467 (N_13467,N_3733,N_1151);
and U13468 (N_13468,N_4938,N_3999);
nor U13469 (N_13469,N_7090,N_8003);
and U13470 (N_13470,N_7478,N_2206);
and U13471 (N_13471,N_2167,N_2030);
and U13472 (N_13472,N_6382,N_2635);
xnor U13473 (N_13473,N_4223,N_7319);
xor U13474 (N_13474,N_3875,N_7939);
xor U13475 (N_13475,N_3726,N_6181);
or U13476 (N_13476,N_1857,N_2235);
xnor U13477 (N_13477,N_7683,N_9152);
xnor U13478 (N_13478,N_7606,N_3736);
nor U13479 (N_13479,N_8874,N_8607);
or U13480 (N_13480,N_6761,N_8324);
nand U13481 (N_13481,N_8794,N_8089);
and U13482 (N_13482,N_4603,N_4354);
or U13483 (N_13483,N_611,N_3266);
and U13484 (N_13484,N_5502,N_3920);
nor U13485 (N_13485,N_4004,N_8209);
xnor U13486 (N_13486,N_7109,N_9556);
nand U13487 (N_13487,N_3659,N_9305);
nor U13488 (N_13488,N_9746,N_8883);
xnor U13489 (N_13489,N_3629,N_6491);
xnor U13490 (N_13490,N_1253,N_7133);
nand U13491 (N_13491,N_9549,N_7748);
nand U13492 (N_13492,N_1611,N_1399);
nor U13493 (N_13493,N_9965,N_9832);
nor U13494 (N_13494,N_8537,N_8049);
xnor U13495 (N_13495,N_4837,N_3596);
or U13496 (N_13496,N_8582,N_4794);
nor U13497 (N_13497,N_1103,N_1146);
and U13498 (N_13498,N_3997,N_3369);
nor U13499 (N_13499,N_4270,N_9443);
xnor U13500 (N_13500,N_2802,N_4040);
nand U13501 (N_13501,N_3025,N_5741);
or U13502 (N_13502,N_1828,N_1351);
nand U13503 (N_13503,N_4052,N_7459);
xor U13504 (N_13504,N_3106,N_6624);
or U13505 (N_13505,N_7521,N_6050);
xor U13506 (N_13506,N_3944,N_6177);
nor U13507 (N_13507,N_3275,N_3683);
and U13508 (N_13508,N_7278,N_4972);
nor U13509 (N_13509,N_1780,N_6330);
and U13510 (N_13510,N_6858,N_6348);
nand U13511 (N_13511,N_739,N_6460);
or U13512 (N_13512,N_3844,N_4043);
or U13513 (N_13513,N_7988,N_9701);
nor U13514 (N_13514,N_284,N_3117);
and U13515 (N_13515,N_3181,N_2001);
xor U13516 (N_13516,N_5359,N_7494);
xnor U13517 (N_13517,N_193,N_2513);
and U13518 (N_13518,N_705,N_7074);
or U13519 (N_13519,N_7946,N_6486);
nor U13520 (N_13520,N_1852,N_9448);
or U13521 (N_13521,N_7116,N_4706);
nand U13522 (N_13522,N_5878,N_4368);
or U13523 (N_13523,N_3548,N_4194);
or U13524 (N_13524,N_1932,N_263);
nor U13525 (N_13525,N_6271,N_6098);
nand U13526 (N_13526,N_3138,N_3271);
nor U13527 (N_13527,N_4950,N_2743);
or U13528 (N_13528,N_9454,N_8351);
nand U13529 (N_13529,N_9763,N_4311);
nand U13530 (N_13530,N_5761,N_9464);
or U13531 (N_13531,N_3810,N_3805);
or U13532 (N_13532,N_5918,N_2117);
nand U13533 (N_13533,N_6774,N_7066);
or U13534 (N_13534,N_4783,N_6744);
and U13535 (N_13535,N_9803,N_3690);
nand U13536 (N_13536,N_1544,N_5842);
nand U13537 (N_13537,N_9098,N_4525);
and U13538 (N_13538,N_2222,N_659);
nor U13539 (N_13539,N_8482,N_8234);
and U13540 (N_13540,N_3191,N_2527);
nand U13541 (N_13541,N_9434,N_5063);
nand U13542 (N_13542,N_2700,N_1840);
nand U13543 (N_13543,N_5601,N_7314);
or U13544 (N_13544,N_796,N_7922);
nor U13545 (N_13545,N_9593,N_4095);
and U13546 (N_13546,N_296,N_8370);
nand U13547 (N_13547,N_6134,N_3616);
and U13548 (N_13548,N_5851,N_233);
and U13549 (N_13549,N_6516,N_9322);
xnor U13550 (N_13550,N_3937,N_2410);
xnor U13551 (N_13551,N_4982,N_7425);
nand U13552 (N_13552,N_5117,N_2353);
nand U13553 (N_13553,N_9006,N_1423);
xor U13554 (N_13554,N_9269,N_3402);
nor U13555 (N_13555,N_4663,N_1003);
nand U13556 (N_13556,N_2498,N_2515);
nand U13557 (N_13557,N_6243,N_2724);
nand U13558 (N_13558,N_574,N_946);
xor U13559 (N_13559,N_1788,N_1417);
nor U13560 (N_13560,N_4871,N_852);
nand U13561 (N_13561,N_289,N_4736);
nor U13562 (N_13562,N_1914,N_657);
xor U13563 (N_13563,N_9810,N_4751);
nor U13564 (N_13564,N_7156,N_27);
or U13565 (N_13565,N_9629,N_8870);
or U13566 (N_13566,N_1593,N_6608);
and U13567 (N_13567,N_1748,N_1064);
or U13568 (N_13568,N_89,N_9507);
nand U13569 (N_13569,N_3411,N_3071);
nor U13570 (N_13570,N_2387,N_124);
nor U13571 (N_13571,N_98,N_319);
xor U13572 (N_13572,N_7599,N_1299);
nand U13573 (N_13573,N_4758,N_4893);
nand U13574 (N_13574,N_1743,N_4594);
or U13575 (N_13575,N_6622,N_7979);
nor U13576 (N_13576,N_6887,N_3060);
nor U13577 (N_13577,N_1034,N_8447);
nand U13578 (N_13578,N_2378,N_1983);
nor U13579 (N_13579,N_9855,N_2352);
nand U13580 (N_13580,N_1262,N_7035);
and U13581 (N_13581,N_7406,N_5996);
xnor U13582 (N_13582,N_8550,N_3657);
or U13583 (N_13583,N_7888,N_3572);
or U13584 (N_13584,N_5725,N_8489);
and U13585 (N_13585,N_1587,N_6531);
xnor U13586 (N_13586,N_8569,N_5921);
xor U13587 (N_13587,N_9411,N_8401);
xnor U13588 (N_13588,N_1297,N_6507);
xor U13589 (N_13589,N_8088,N_7434);
or U13590 (N_13590,N_6496,N_9234);
nand U13591 (N_13591,N_5443,N_9807);
or U13592 (N_13592,N_2973,N_262);
nand U13593 (N_13593,N_5266,N_3171);
nand U13594 (N_13594,N_5051,N_6888);
xor U13595 (N_13595,N_5385,N_9606);
or U13596 (N_13596,N_3487,N_629);
or U13597 (N_13597,N_7645,N_5945);
or U13598 (N_13598,N_9477,N_8313);
or U13599 (N_13599,N_8292,N_7214);
xnor U13600 (N_13600,N_3477,N_1446);
xnor U13601 (N_13601,N_5339,N_278);
xnor U13602 (N_13602,N_4288,N_8031);
and U13603 (N_13603,N_4672,N_688);
nor U13604 (N_13604,N_5365,N_7483);
xor U13605 (N_13605,N_8381,N_6131);
or U13606 (N_13606,N_1735,N_5459);
nor U13607 (N_13607,N_3378,N_8736);
and U13608 (N_13608,N_5940,N_9979);
xor U13609 (N_13609,N_4309,N_112);
xnor U13610 (N_13610,N_978,N_1569);
or U13611 (N_13611,N_488,N_9788);
or U13612 (N_13612,N_8767,N_226);
nor U13613 (N_13613,N_1487,N_8975);
and U13614 (N_13614,N_7295,N_4720);
nor U13615 (N_13615,N_4637,N_5969);
nor U13616 (N_13616,N_2031,N_2848);
or U13617 (N_13617,N_6362,N_4845);
and U13618 (N_13618,N_6124,N_4379);
and U13619 (N_13619,N_9144,N_1863);
nand U13620 (N_13620,N_1263,N_1860);
nand U13621 (N_13621,N_7732,N_1524);
xor U13622 (N_13622,N_5112,N_5017);
xnor U13623 (N_13623,N_8001,N_9996);
and U13624 (N_13624,N_3618,N_1657);
nand U13625 (N_13625,N_47,N_6453);
nand U13626 (N_13626,N_4962,N_4634);
and U13627 (N_13627,N_6351,N_6095);
xor U13628 (N_13628,N_7309,N_371);
nand U13629 (N_13629,N_3507,N_9861);
nor U13630 (N_13630,N_4293,N_9819);
and U13631 (N_13631,N_1664,N_88);
nand U13632 (N_13632,N_1557,N_624);
xor U13633 (N_13633,N_1107,N_4484);
nor U13634 (N_13634,N_8380,N_697);
nor U13635 (N_13635,N_5268,N_2531);
xnor U13636 (N_13636,N_5030,N_9869);
xor U13637 (N_13637,N_1015,N_5486);
or U13638 (N_13638,N_3968,N_1358);
xnor U13639 (N_13639,N_4759,N_5202);
xor U13640 (N_13640,N_5840,N_6242);
nand U13641 (N_13641,N_9230,N_2719);
nor U13642 (N_13642,N_2017,N_9050);
or U13643 (N_13643,N_736,N_3359);
and U13644 (N_13644,N_3244,N_759);
xnor U13645 (N_13645,N_6954,N_1123);
nor U13646 (N_13646,N_2596,N_7604);
or U13647 (N_13647,N_1077,N_3312);
or U13648 (N_13648,N_2286,N_6378);
or U13649 (N_13649,N_1981,N_6683);
and U13650 (N_13650,N_795,N_9958);
nand U13651 (N_13651,N_3555,N_6570);
nand U13652 (N_13652,N_2608,N_7071);
and U13653 (N_13653,N_9511,N_4061);
xor U13654 (N_13654,N_1441,N_4682);
nor U13655 (N_13655,N_4987,N_7515);
or U13656 (N_13656,N_6314,N_38);
and U13657 (N_13657,N_6106,N_8312);
nand U13658 (N_13658,N_6694,N_4828);
xnor U13659 (N_13659,N_6711,N_4307);
and U13660 (N_13660,N_4365,N_4369);
or U13661 (N_13661,N_3512,N_8263);
and U13662 (N_13662,N_5796,N_2336);
or U13663 (N_13663,N_8672,N_9254);
nand U13664 (N_13664,N_7635,N_7444);
nor U13665 (N_13665,N_2811,N_8801);
and U13666 (N_13666,N_9644,N_7560);
xnor U13667 (N_13667,N_8666,N_1154);
or U13668 (N_13668,N_8860,N_6029);
xor U13669 (N_13669,N_3698,N_8446);
and U13670 (N_13670,N_2075,N_4725);
or U13671 (N_13671,N_6881,N_8288);
or U13672 (N_13672,N_3791,N_6859);
nand U13673 (N_13673,N_827,N_3523);
nor U13674 (N_13674,N_9604,N_2399);
and U13675 (N_13675,N_6093,N_7920);
xor U13676 (N_13676,N_7500,N_6027);
and U13677 (N_13677,N_2400,N_6628);
nand U13678 (N_13678,N_1247,N_6034);
and U13679 (N_13679,N_141,N_5783);
nor U13680 (N_13680,N_249,N_5706);
nor U13681 (N_13681,N_4037,N_6955);
and U13682 (N_13682,N_8540,N_81);
nand U13683 (N_13683,N_7953,N_7805);
nor U13684 (N_13684,N_7254,N_8953);
xor U13685 (N_13685,N_9749,N_4535);
and U13686 (N_13686,N_3622,N_6627);
or U13687 (N_13687,N_1513,N_9546);
and U13688 (N_13688,N_1520,N_8972);
xnor U13689 (N_13689,N_2525,N_9524);
xor U13690 (N_13690,N_7577,N_6665);
xnor U13691 (N_13691,N_1304,N_6549);
or U13692 (N_13692,N_9226,N_6811);
or U13693 (N_13693,N_4103,N_744);
nand U13694 (N_13694,N_8511,N_798);
or U13695 (N_13695,N_159,N_9517);
nor U13696 (N_13696,N_8390,N_4479);
or U13697 (N_13697,N_2165,N_3420);
or U13698 (N_13698,N_6732,N_8844);
and U13699 (N_13699,N_5838,N_2005);
nor U13700 (N_13700,N_8888,N_5204);
xnor U13701 (N_13701,N_7119,N_7358);
nor U13702 (N_13702,N_4714,N_2879);
nor U13703 (N_13703,N_385,N_2694);
nor U13704 (N_13704,N_7868,N_588);
xor U13705 (N_13705,N_3607,N_9690);
nand U13706 (N_13706,N_6835,N_8806);
nor U13707 (N_13707,N_5846,N_1300);
nor U13708 (N_13708,N_572,N_4671);
xor U13709 (N_13709,N_7526,N_5461);
xor U13710 (N_13710,N_4711,N_4619);
xor U13711 (N_13711,N_4411,N_4531);
and U13712 (N_13712,N_8354,N_3096);
or U13713 (N_13713,N_6033,N_3169);
or U13714 (N_13714,N_29,N_398);
xor U13715 (N_13715,N_525,N_8717);
and U13716 (N_13716,N_6500,N_9134);
nand U13717 (N_13717,N_5347,N_9583);
and U13718 (N_13718,N_9276,N_1277);
nor U13719 (N_13719,N_3846,N_6441);
nand U13720 (N_13720,N_8798,N_2936);
xnor U13721 (N_13721,N_1410,N_9340);
nand U13722 (N_13722,N_9162,N_2128);
xor U13723 (N_13723,N_2432,N_7139);
and U13724 (N_13724,N_8657,N_4143);
and U13725 (N_13725,N_6593,N_4790);
or U13726 (N_13726,N_3238,N_8781);
xor U13727 (N_13727,N_5060,N_9497);
nor U13728 (N_13728,N_5774,N_6030);
xnor U13729 (N_13729,N_6655,N_5894);
or U13730 (N_13730,N_8812,N_1037);
nor U13731 (N_13731,N_3557,N_9428);
and U13732 (N_13732,N_6728,N_8126);
or U13733 (N_13733,N_5963,N_6595);
and U13734 (N_13734,N_7902,N_809);
or U13735 (N_13735,N_5820,N_9001);
xor U13736 (N_13736,N_8057,N_1398);
xnor U13737 (N_13737,N_3388,N_2634);
nand U13738 (N_13738,N_4687,N_4866);
or U13739 (N_13739,N_980,N_1898);
or U13740 (N_13740,N_3549,N_4165);
nand U13741 (N_13741,N_2468,N_8358);
and U13742 (N_13742,N_4928,N_7158);
or U13743 (N_13743,N_2960,N_1320);
and U13744 (N_13744,N_7329,N_9263);
and U13745 (N_13745,N_8058,N_7884);
nor U13746 (N_13746,N_8945,N_8000);
and U13747 (N_13747,N_8998,N_417);
and U13748 (N_13748,N_388,N_7420);
xor U13749 (N_13749,N_3472,N_9840);
xnor U13750 (N_13750,N_1230,N_3250);
or U13751 (N_13751,N_4185,N_1892);
and U13752 (N_13752,N_448,N_4630);
nand U13753 (N_13753,N_403,N_5231);
nand U13754 (N_13754,N_3541,N_4220);
or U13755 (N_13755,N_7747,N_9523);
xnor U13756 (N_13756,N_8879,N_9444);
nand U13757 (N_13757,N_608,N_6461);
nand U13758 (N_13758,N_763,N_451);
or U13759 (N_13759,N_3859,N_3316);
and U13760 (N_13760,N_3258,N_7600);
nor U13761 (N_13761,N_5909,N_8898);
or U13762 (N_13762,N_9718,N_2643);
or U13763 (N_13763,N_8202,N_6232);
and U13764 (N_13764,N_8141,N_6653);
xnor U13765 (N_13765,N_9426,N_7720);
nor U13766 (N_13766,N_728,N_6535);
and U13767 (N_13767,N_762,N_8224);
or U13768 (N_13768,N_6522,N_6078);
nor U13769 (N_13769,N_2946,N_3108);
and U13770 (N_13770,N_5779,N_3573);
or U13771 (N_13771,N_2963,N_300);
or U13772 (N_13772,N_9848,N_9193);
or U13773 (N_13773,N_9294,N_1169);
nand U13774 (N_13774,N_441,N_7639);
and U13775 (N_13775,N_2507,N_7337);
and U13776 (N_13776,N_4018,N_8877);
and U13777 (N_13777,N_6942,N_1095);
and U13778 (N_13778,N_3917,N_65);
nor U13779 (N_13779,N_2502,N_4153);
or U13780 (N_13780,N_5223,N_7443);
and U13781 (N_13781,N_742,N_1706);
and U13782 (N_13782,N_4829,N_1730);
nand U13783 (N_13783,N_4773,N_769);
or U13784 (N_13784,N_2296,N_4101);
and U13785 (N_13785,N_8252,N_3127);
or U13786 (N_13786,N_875,N_3686);
nor U13787 (N_13787,N_1329,N_4199);
nand U13788 (N_13788,N_6789,N_7190);
and U13789 (N_13789,N_1739,N_8814);
xor U13790 (N_13790,N_1645,N_3082);
nor U13791 (N_13791,N_5527,N_3254);
nor U13792 (N_13792,N_7697,N_6935);
or U13793 (N_13793,N_1429,N_3083);
or U13794 (N_13794,N_8368,N_554);
nand U13795 (N_13795,N_1401,N_3671);
nor U13796 (N_13796,N_667,N_1350);
and U13797 (N_13797,N_9495,N_6739);
and U13798 (N_13798,N_9101,N_8465);
nor U13799 (N_13799,N_9013,N_1903);
nor U13800 (N_13800,N_242,N_5168);
or U13801 (N_13801,N_9352,N_8670);
xnor U13802 (N_13802,N_1853,N_6437);
xnor U13803 (N_13803,N_1414,N_8530);
nand U13804 (N_13804,N_7974,N_6731);
nand U13805 (N_13805,N_2269,N_7736);
nor U13806 (N_13806,N_1680,N_5369);
or U13807 (N_13807,N_9158,N_5187);
or U13808 (N_13808,N_3414,N_1081);
and U13809 (N_13809,N_1667,N_5856);
or U13810 (N_13810,N_7912,N_5100);
nor U13811 (N_13811,N_4992,N_3812);
nor U13812 (N_13812,N_9899,N_6727);
nand U13813 (N_13813,N_7398,N_239);
nor U13814 (N_13814,N_4142,N_1913);
xnor U13815 (N_13815,N_9088,N_7673);
xor U13816 (N_13816,N_6012,N_3215);
xor U13817 (N_13817,N_1268,N_5564);
nand U13818 (N_13818,N_3441,N_7659);
xnor U13819 (N_13819,N_3836,N_6533);
or U13820 (N_13820,N_1958,N_5734);
nor U13821 (N_13821,N_1164,N_395);
xnor U13822 (N_13822,N_9129,N_430);
nor U13823 (N_13823,N_4593,N_1604);
nor U13824 (N_13824,N_325,N_6053);
nor U13825 (N_13825,N_636,N_9315);
xor U13826 (N_13826,N_5658,N_3198);
or U13827 (N_13827,N_9821,N_3689);
nand U13828 (N_13828,N_8911,N_4136);
or U13829 (N_13829,N_4407,N_9074);
nand U13830 (N_13830,N_4914,N_134);
xor U13831 (N_13831,N_8359,N_3631);
nand U13832 (N_13832,N_4196,N_716);
and U13833 (N_13833,N_8954,N_3760);
or U13834 (N_13834,N_4515,N_4995);
nor U13835 (N_13835,N_2590,N_783);
nand U13836 (N_13836,N_2294,N_1996);
xor U13837 (N_13837,N_5926,N_1944);
nand U13838 (N_13838,N_1271,N_5287);
and U13839 (N_13839,N_3424,N_5014);
xor U13840 (N_13840,N_9480,N_7539);
nor U13841 (N_13841,N_5943,N_3218);
xor U13842 (N_13842,N_2846,N_9280);
or U13843 (N_13843,N_3142,N_9218);
or U13844 (N_13844,N_8967,N_2748);
xnor U13845 (N_13845,N_7334,N_1829);
and U13846 (N_13846,N_1306,N_454);
xor U13847 (N_13847,N_7792,N_3609);
or U13848 (N_13848,N_5749,N_2609);
nor U13849 (N_13849,N_7892,N_5949);
nand U13850 (N_13850,N_1222,N_4749);
and U13851 (N_13851,N_7791,N_873);
and U13852 (N_13852,N_5776,N_5028);
and U13853 (N_13853,N_2129,N_9540);
nor U13854 (N_13854,N_853,N_3242);
and U13855 (N_13855,N_5652,N_4055);
xnor U13856 (N_13856,N_4897,N_9638);
or U13857 (N_13857,N_4273,N_1747);
nand U13858 (N_13858,N_6668,N_7894);
xor U13859 (N_13859,N_4627,N_5023);
and U13860 (N_13860,N_9041,N_7381);
nor U13861 (N_13861,N_2173,N_8087);
xor U13862 (N_13862,N_6743,N_8171);
or U13863 (N_13863,N_7763,N_2398);
xor U13864 (N_13864,N_8834,N_6157);
or U13865 (N_13865,N_1591,N_1397);
and U13866 (N_13866,N_3849,N_9067);
xor U13867 (N_13867,N_5603,N_8330);
nor U13868 (N_13868,N_4230,N_8591);
and U13869 (N_13869,N_6515,N_7141);
nand U13870 (N_13870,N_6197,N_7137);
and U13871 (N_13871,N_1714,N_2467);
and U13872 (N_13872,N_3338,N_9570);
nand U13873 (N_13873,N_326,N_4446);
nand U13874 (N_13874,N_9845,N_9854);
nor U13875 (N_13875,N_1620,N_4447);
nor U13876 (N_13876,N_366,N_7408);
nor U13877 (N_13877,N_8276,N_2225);
xnor U13878 (N_13878,N_2335,N_1629);
or U13879 (N_13879,N_4591,N_4162);
nor U13880 (N_13880,N_4924,N_1633);
xor U13881 (N_13881,N_1101,N_4819);
or U13882 (N_13882,N_4902,N_2595);
nor U13883 (N_13883,N_2411,N_8778);
nand U13884 (N_13884,N_4957,N_1155);
nor U13885 (N_13885,N_1276,N_2340);
or U13886 (N_13886,N_4644,N_5106);
or U13887 (N_13887,N_2278,N_5760);
or U13888 (N_13888,N_9731,N_4282);
xnor U13889 (N_13889,N_9492,N_3601);
nor U13890 (N_13890,N_7477,N_1969);
xnor U13891 (N_13891,N_1439,N_5651);
xor U13892 (N_13892,N_6221,N_7102);
xor U13893 (N_13893,N_9228,N_3381);
or U13894 (N_13894,N_2563,N_7145);
nor U13895 (N_13895,N_4325,N_4388);
nor U13896 (N_13896,N_2727,N_4291);
and U13897 (N_13897,N_9102,N_3382);
xnor U13898 (N_13898,N_8699,N_3047);
or U13899 (N_13899,N_1039,N_9089);
nor U13900 (N_13900,N_9888,N_7237);
nand U13901 (N_13901,N_247,N_8301);
nor U13902 (N_13902,N_8187,N_5524);
and U13903 (N_13903,N_8050,N_5077);
nand U13904 (N_13904,N_2121,N_3406);
nor U13905 (N_13905,N_4284,N_9298);
or U13906 (N_13906,N_9587,N_9820);
or U13907 (N_13907,N_9515,N_4842);
or U13908 (N_13908,N_5550,N_3649);
or U13909 (N_13909,N_3907,N_900);
xor U13910 (N_13910,N_4215,N_1317);
or U13911 (N_13911,N_6040,N_4554);
and U13912 (N_13912,N_7507,N_4324);
nand U13913 (N_13913,N_3538,N_7964);
nand U13914 (N_13914,N_3751,N_8231);
nand U13915 (N_13915,N_2894,N_2311);
nor U13916 (N_13916,N_5317,N_4978);
or U13917 (N_13917,N_9522,N_7204);
xor U13918 (N_13918,N_5901,N_7609);
xor U13919 (N_13919,N_3932,N_766);
nand U13920 (N_13920,N_8290,N_7987);
xnor U13921 (N_13921,N_6257,N_437);
or U13922 (N_13922,N_6096,N_9641);
xnor U13923 (N_13923,N_6319,N_5773);
or U13924 (N_13924,N_4360,N_6449);
or U13925 (N_13925,N_246,N_5688);
nand U13926 (N_13926,N_7210,N_4349);
nand U13927 (N_13927,N_712,N_1192);
and U13928 (N_13928,N_8740,N_1516);
xor U13929 (N_13929,N_9816,N_2666);
or U13930 (N_13930,N_1258,N_1387);
nor U13931 (N_13931,N_7731,N_3006);
nor U13932 (N_13932,N_6707,N_331);
and U13933 (N_13933,N_5770,N_5089);
nor U13934 (N_13934,N_768,N_4713);
nor U13935 (N_13935,N_5655,N_7671);
xnor U13936 (N_13936,N_9046,N_3212);
nand U13937 (N_13937,N_7711,N_6129);
nor U13938 (N_13938,N_9354,N_8216);
and U13939 (N_13939,N_544,N_2384);
or U13940 (N_13940,N_1335,N_2369);
or U13941 (N_13941,N_1649,N_7802);
nand U13942 (N_13942,N_2786,N_8902);
or U13943 (N_13943,N_6924,N_7664);
nand U13944 (N_13944,N_3221,N_7667);
or U13945 (N_13945,N_6956,N_6225);
nand U13946 (N_13946,N_2448,N_8118);
xnor U13947 (N_13947,N_5219,N_9185);
or U13948 (N_13948,N_5004,N_1278);
and U13949 (N_13949,N_7054,N_6467);
nand U13950 (N_13950,N_4727,N_1666);
xor U13951 (N_13951,N_4501,N_7387);
or U13952 (N_13952,N_1576,N_3427);
and U13953 (N_13953,N_9069,N_6994);
nor U13954 (N_13954,N_2078,N_485);
and U13955 (N_13955,N_7652,N_575);
or U13956 (N_13956,N_720,N_4398);
xor U13957 (N_13957,N_1183,N_7242);
nor U13958 (N_13958,N_1100,N_7206);
nor U13959 (N_13959,N_675,N_6583);
nand U13960 (N_13960,N_9299,N_4239);
xor U13961 (N_13961,N_5855,N_8107);
and U13962 (N_13962,N_7824,N_3115);
xor U13963 (N_13963,N_1803,N_6552);
or U13964 (N_13964,N_800,N_5300);
or U13965 (N_13965,N_8320,N_1272);
nor U13966 (N_13966,N_3086,N_8291);
and U13967 (N_13967,N_6195,N_9897);
xnor U13968 (N_13968,N_9698,N_8436);
nor U13969 (N_13969,N_8682,N_6346);
nand U13970 (N_13970,N_1436,N_5078);
and U13971 (N_13971,N_8366,N_9100);
xnor U13972 (N_13972,N_4753,N_3499);
or U13973 (N_13973,N_6193,N_3422);
nand U13974 (N_13974,N_4932,N_6504);
xor U13975 (N_13975,N_3560,N_8852);
nor U13976 (N_13976,N_7431,N_8633);
and U13977 (N_13977,N_2746,N_5597);
xnor U13978 (N_13978,N_1963,N_7487);
or U13979 (N_13979,N_1336,N_7596);
xnor U13980 (N_13980,N_3602,N_4377);
nor U13981 (N_13981,N_3120,N_516);
xnor U13982 (N_13982,N_3885,N_3648);
nor U13983 (N_13983,N_8578,N_2599);
nor U13984 (N_13984,N_880,N_5518);
and U13985 (N_13985,N_1877,N_3227);
xor U13986 (N_13986,N_461,N_1922);
or U13987 (N_13987,N_7396,N_8080);
nor U13988 (N_13988,N_6560,N_8897);
nor U13989 (N_13989,N_6968,N_7777);
or U13990 (N_13990,N_9431,N_9700);
nor U13991 (N_13991,N_3500,N_2773);
and U13992 (N_13992,N_8523,N_8327);
nor U13993 (N_13993,N_2326,N_2665);
nand U13994 (N_13994,N_4993,N_1376);
nand U13995 (N_13995,N_2274,N_799);
and U13996 (N_13996,N_1202,N_9095);
or U13997 (N_13997,N_5629,N_5377);
nand U13998 (N_13998,N_9814,N_9563);
or U13999 (N_13999,N_7181,N_6699);
or U14000 (N_14000,N_2027,N_6224);
or U14001 (N_14001,N_7161,N_3151);
nor U14002 (N_14002,N_2301,N_7843);
and U14003 (N_14003,N_6414,N_1219);
nand U14004 (N_14004,N_7787,N_6178);
xor U14005 (N_14005,N_4110,N_1437);
xor U14006 (N_14006,N_5393,N_4202);
xor U14007 (N_14007,N_817,N_983);
nand U14008 (N_14008,N_2661,N_7877);
xnor U14009 (N_14009,N_9242,N_7856);
xnor U14010 (N_14010,N_5296,N_5888);
nand U14011 (N_14011,N_4080,N_6558);
and U14012 (N_14012,N_5748,N_8805);
xnor U14013 (N_14013,N_6630,N_2098);
or U14014 (N_14014,N_5708,N_3505);
nor U14015 (N_14015,N_8432,N_217);
xor U14016 (N_14016,N_9882,N_2968);
xor U14017 (N_14017,N_8810,N_6791);
or U14018 (N_14018,N_308,N_7834);
or U14019 (N_14019,N_6617,N_4561);
nor U14020 (N_14020,N_3468,N_6017);
nor U14021 (N_14021,N_7815,N_7166);
xor U14022 (N_14022,N_8339,N_1224);
nand U14023 (N_14023,N_7917,N_2360);
xor U14024 (N_14024,N_5876,N_6063);
or U14025 (N_14025,N_3297,N_5241);
nor U14026 (N_14026,N_1327,N_7088);
and U14027 (N_14027,N_8250,N_2293);
nand U14028 (N_14028,N_9901,N_3606);
or U14029 (N_14029,N_206,N_5);
nand U14030 (N_14030,N_3122,N_7220);
nand U14031 (N_14031,N_6676,N_2644);
and U14032 (N_14032,N_6184,N_5389);
or U14033 (N_14033,N_8142,N_8214);
xor U14034 (N_14034,N_6091,N_6847);
or U14035 (N_14035,N_1975,N_6149);
nor U14036 (N_14036,N_119,N_7661);
xnor U14037 (N_14037,N_7698,N_7844);
xnor U14038 (N_14038,N_327,N_7080);
nand U14039 (N_14039,N_6139,N_1408);
nand U14040 (N_14040,N_1522,N_8035);
nor U14041 (N_14041,N_5985,N_2535);
or U14042 (N_14042,N_5875,N_5724);
and U14043 (N_14043,N_7699,N_443);
nand U14044 (N_14044,N_3553,N_5094);
xnor U14045 (N_14045,N_6587,N_8299);
and U14046 (N_14046,N_4472,N_5839);
nand U14047 (N_14047,N_8572,N_3608);
xor U14048 (N_14048,N_2967,N_6693);
or U14049 (N_14049,N_7272,N_221);
and U14050 (N_14050,N_1498,N_8989);
nand U14051 (N_14051,N_1227,N_8373);
and U14052 (N_14052,N_1685,N_1085);
nand U14053 (N_14053,N_4536,N_2702);
and U14054 (N_14054,N_4846,N_1884);
nand U14055 (N_14055,N_7436,N_4493);
nand U14056 (N_14056,N_3723,N_9275);
xnor U14057 (N_14057,N_2921,N_8565);
xor U14058 (N_14058,N_3970,N_6856);
or U14059 (N_14059,N_1943,N_5578);
nor U14060 (N_14060,N_2709,N_7835);
and U14061 (N_14061,N_2695,N_4338);
nor U14062 (N_14062,N_280,N_9301);
nand U14063 (N_14063,N_5034,N_7620);
nand U14064 (N_14064,N_5301,N_8688);
nand U14065 (N_14065,N_1746,N_208);
and U14066 (N_14066,N_6410,N_3088);
or U14067 (N_14067,N_4596,N_5343);
nor U14068 (N_14068,N_9961,N_1082);
xnor U14069 (N_14069,N_662,N_3524);
nor U14070 (N_14070,N_1232,N_9589);
nor U14071 (N_14071,N_4690,N_967);
nor U14072 (N_14072,N_2519,N_9932);
nor U14073 (N_14073,N_8208,N_5987);
nor U14074 (N_14074,N_6842,N_8833);
nor U14075 (N_14075,N_2907,N_672);
xnor U14076 (N_14076,N_9970,N_9133);
and U14077 (N_14077,N_4917,N_4584);
nor U14078 (N_14078,N_4428,N_3792);
nand U14079 (N_14079,N_2549,N_4623);
xor U14080 (N_14080,N_6276,N_5618);
nor U14081 (N_14081,N_8757,N_2825);
nor U14082 (N_14082,N_6562,N_3969);
xor U14083 (N_14083,N_2957,N_1875);
nand U14084 (N_14084,N_6011,N_97);
xor U14085 (N_14085,N_1055,N_6976);
nor U14086 (N_14086,N_9279,N_3186);
nor U14087 (N_14087,N_8309,N_8117);
xor U14088 (N_14088,N_4251,N_1364);
nor U14089 (N_14089,N_2362,N_6564);
xor U14090 (N_14090,N_8516,N_5666);
nand U14091 (N_14091,N_4257,N_1842);
and U14092 (N_14092,N_3634,N_1206);
or U14093 (N_14093,N_9862,N_5781);
nand U14094 (N_14094,N_3966,N_3141);
nand U14095 (N_14095,N_513,N_5242);
xnor U14096 (N_14096,N_4798,N_4050);
or U14097 (N_14097,N_9676,N_1252);
xor U14098 (N_14098,N_5907,N_6610);
nor U14099 (N_14099,N_6282,N_4718);
or U14100 (N_14100,N_9407,N_3820);
nor U14101 (N_14101,N_9177,N_1601);
nand U14102 (N_14102,N_8541,N_9096);
nor U14103 (N_14103,N_6697,N_5703);
nand U14104 (N_14104,N_9266,N_2023);
xnor U14105 (N_14105,N_4695,N_9964);
xor U14106 (N_14106,N_5599,N_7945);
and U14107 (N_14107,N_8011,N_3882);
and U14108 (N_14108,N_5240,N_7770);
and U14109 (N_14109,N_8841,N_7085);
and U14110 (N_14110,N_6708,N_253);
xor U14111 (N_14111,N_8289,N_522);
and U14112 (N_14112,N_6137,N_7807);
nor U14113 (N_14113,N_55,N_6013);
and U14114 (N_14114,N_8929,N_7177);
nor U14115 (N_14115,N_6380,N_9321);
nand U14116 (N_14116,N_8966,N_7646);
and U14117 (N_14117,N_4231,N_3874);
xor U14118 (N_14118,N_6127,N_2986);
nor U14119 (N_14119,N_5157,N_5747);
or U14120 (N_14120,N_701,N_1919);
xnor U14121 (N_14121,N_7227,N_4114);
or U14122 (N_14122,N_39,N_4366);
xnor U14123 (N_14123,N_9721,N_155);
nand U14124 (N_14124,N_3745,N_6950);
nand U14125 (N_14125,N_1079,N_3898);
and U14126 (N_14126,N_547,N_146);
nor U14127 (N_14127,N_5033,N_969);
and U14128 (N_14128,N_2956,N_7738);
or U14129 (N_14129,N_1586,N_5891);
xor U14130 (N_14130,N_7403,N_7803);
nor U14131 (N_14131,N_3380,N_9364);
and U14132 (N_14132,N_7219,N_9712);
nand U14133 (N_14133,N_393,N_7323);
or U14134 (N_14134,N_9073,N_8400);
nand U14135 (N_14135,N_6306,N_179);
nor U14136 (N_14136,N_1009,N_3637);
xnor U14137 (N_14137,N_8448,N_9291);
and U14138 (N_14138,N_5191,N_9847);
or U14139 (N_14139,N_2244,N_9774);
and U14140 (N_14140,N_2295,N_3187);
xnor U14141 (N_14141,N_6400,N_7325);
or U14142 (N_14142,N_5001,N_5588);
xnor U14143 (N_14143,N_3462,N_3893);
or U14144 (N_14144,N_4268,N_7423);
or U14145 (N_14145,N_6331,N_4949);
nor U14146 (N_14146,N_8907,N_468);
nand U14147 (N_14147,N_7473,N_8816);
nor U14148 (N_14148,N_3779,N_1598);
or U14149 (N_14149,N_3550,N_4503);
xnor U14150 (N_14150,N_383,N_6918);
or U14151 (N_14151,N_4854,N_3817);
xor U14152 (N_14152,N_7513,N_4954);
or U14153 (N_14153,N_5549,N_3786);
nand U14154 (N_14154,N_1485,N_4508);
nor U14155 (N_14155,N_2996,N_7786);
or U14156 (N_14156,N_4261,N_3094);
or U14157 (N_14157,N_9232,N_9189);
nor U14158 (N_14158,N_8211,N_9838);
and U14159 (N_14159,N_6394,N_1229);
nor U14160 (N_14160,N_3392,N_901);
nand U14161 (N_14161,N_1166,N_8887);
or U14162 (N_14162,N_8538,N_7690);
xnor U14163 (N_14163,N_6505,N_7148);
nand U14164 (N_14164,N_4572,N_4346);
nor U14165 (N_14165,N_5823,N_9092);
and U14166 (N_14166,N_2959,N_9429);
nor U14167 (N_14167,N_7456,N_2219);
and U14168 (N_14168,N_2279,N_585);
nand U14169 (N_14169,N_9975,N_8942);
nor U14170 (N_14170,N_2703,N_9118);
nor U14171 (N_14171,N_4345,N_2856);
xnor U14172 (N_14172,N_3635,N_8165);
or U14173 (N_14173,N_2201,N_9130);
or U14174 (N_14174,N_6720,N_7706);
nand U14175 (N_14175,N_9809,N_1120);
nand U14176 (N_14176,N_5646,N_9529);
nor U14177 (N_14177,N_3566,N_1631);
nand U14178 (N_14178,N_9004,N_7950);
nand U14179 (N_14179,N_1454,N_5551);
or U14180 (N_14180,N_5387,N_3928);
or U14181 (N_14181,N_1287,N_7044);
nor U14182 (N_14182,N_5054,N_5634);
nand U14183 (N_14183,N_954,N_7018);
nor U14184 (N_14184,N_6625,N_6582);
nand U14185 (N_14185,N_5480,N_1382);
nor U14186 (N_14186,N_9467,N_1582);
or U14187 (N_14187,N_5596,N_1908);
nor U14188 (N_14188,N_8458,N_9425);
nand U14189 (N_14189,N_6462,N_2277);
and U14190 (N_14190,N_7013,N_851);
or U14191 (N_14191,N_8175,N_7574);
nand U14192 (N_14192,N_2630,N_6444);
and U14193 (N_14193,N_2061,N_9806);
nor U14194 (N_14194,N_196,N_4258);
and U14195 (N_14195,N_62,N_5306);
xnor U14196 (N_14196,N_9924,N_1984);
xnor U14197 (N_14197,N_3190,N_6824);
xnor U14198 (N_14198,N_9231,N_6787);
nand U14199 (N_14199,N_9012,N_5442);
xor U14200 (N_14200,N_9391,N_3714);
and U14201 (N_14201,N_4347,N_7152);
or U14202 (N_14202,N_9278,N_1843);
nor U14203 (N_14203,N_299,N_5085);
nor U14204 (N_14204,N_8741,N_7291);
nor U14205 (N_14205,N_1346,N_9689);
and U14206 (N_14206,N_9867,N_9615);
nand U14207 (N_14207,N_6032,N_7774);
or U14208 (N_14208,N_4879,N_4652);
xnor U14209 (N_14209,N_8604,N_4573);
nand U14210 (N_14210,N_7371,N_6963);
and U14211 (N_14211,N_8282,N_3002);
nor U14212 (N_14212,N_374,N_2688);
nand U14213 (N_14213,N_7496,N_5554);
nand U14214 (N_14214,N_3283,N_3856);
and U14215 (N_14215,N_4767,N_4410);
nor U14216 (N_14216,N_8931,N_194);
or U14217 (N_14217,N_7781,N_2781);
xnor U14218 (N_14218,N_3706,N_3973);
nor U14219 (N_14219,N_6018,N_4163);
xnor U14220 (N_14220,N_5735,N_245);
nand U14221 (N_14221,N_1669,N_733);
nand U14222 (N_14222,N_6611,N_1856);
nor U14223 (N_14223,N_541,N_658);
nor U14224 (N_14224,N_1024,N_4852);
nor U14225 (N_14225,N_3103,N_5375);
and U14226 (N_14226,N_3703,N_4723);
nor U14227 (N_14227,N_332,N_4328);
nor U14228 (N_14228,N_1565,N_4442);
nand U14229 (N_14229,N_5307,N_401);
xor U14230 (N_14230,N_2174,N_8943);
and U14231 (N_14231,N_9934,N_9550);
nor U14232 (N_14232,N_4802,N_1440);
and U14233 (N_14233,N_9498,N_7307);
nor U14234 (N_14234,N_7430,N_3077);
nand U14235 (N_14235,N_68,N_5145);
nor U14236 (N_14236,N_2929,N_6142);
nand U14237 (N_14237,N_8340,N_320);
nand U14238 (N_14238,N_3056,N_9684);
or U14239 (N_14239,N_6301,N_9366);
or U14240 (N_14240,N_7450,N_5473);
or U14241 (N_14241,N_2127,N_5682);
nand U14242 (N_14242,N_6685,N_7195);
xor U14243 (N_14243,N_1789,N_8997);
or U14244 (N_14244,N_9284,N_2845);
nor U14245 (N_14245,N_6829,N_8919);
xor U14246 (N_14246,N_3205,N_3042);
and U14247 (N_14247,N_3643,N_3284);
xor U14248 (N_14248,N_2545,N_4602);
nor U14249 (N_14249,N_8746,N_2297);
nand U14250 (N_14250,N_7174,N_6473);
and U14251 (N_14251,N_2804,N_6502);
or U14252 (N_14252,N_7015,N_9631);
and U14253 (N_14253,N_4888,N_3432);
nor U14254 (N_14254,N_4431,N_127);
or U14255 (N_14255,N_8102,N_8466);
or U14256 (N_14256,N_306,N_3709);
nor U14257 (N_14257,N_8405,N_3247);
nor U14258 (N_14258,N_8223,N_4312);
nand U14259 (N_14259,N_6056,N_465);
xor U14260 (N_14260,N_2124,N_4333);
and U14261 (N_14261,N_7931,N_1057);
nand U14262 (N_14262,N_3489,N_4075);
nand U14263 (N_14263,N_1135,N_9483);
xnor U14264 (N_14264,N_8024,N_5965);
xnor U14265 (N_14265,N_8555,N_7188);
nand U14266 (N_14266,N_324,N_4818);
and U14267 (N_14267,N_4612,N_6606);
or U14268 (N_14268,N_4313,N_2406);
nand U14269 (N_14269,N_7455,N_9510);
nor U14270 (N_14270,N_6736,N_1348);
or U14271 (N_14271,N_4086,N_8471);
nor U14272 (N_14272,N_9139,N_5274);
nand U14273 (N_14273,N_3301,N_1476);
or U14274 (N_14274,N_8486,N_4558);
xnor U14275 (N_14275,N_2872,N_8131);
nand U14276 (N_14276,N_4689,N_6980);
and U14277 (N_14277,N_9562,N_3300);
nor U14278 (N_14278,N_4646,N_3032);
nor U14279 (N_14279,N_505,N_6047);
and U14280 (N_14280,N_5559,N_8182);
and U14281 (N_14281,N_3053,N_8861);
nand U14282 (N_14282,N_1872,N_7292);
xor U14283 (N_14283,N_3599,N_6227);
or U14284 (N_14284,N_952,N_1831);
xnor U14285 (N_14285,N_156,N_8077);
and U14286 (N_14286,N_8060,N_5132);
xor U14287 (N_14287,N_8501,N_282);
and U14288 (N_14288,N_9192,N_9062);
xor U14289 (N_14289,N_6381,N_3679);
xnor U14290 (N_14290,N_8603,N_6651);
xor U14291 (N_14291,N_7789,N_1430);
nor U14292 (N_14292,N_3803,N_1188);
and U14293 (N_14293,N_5692,N_7002);
nand U14294 (N_14294,N_1982,N_6613);
and U14295 (N_14295,N_8593,N_782);
xor U14296 (N_14296,N_2681,N_7913);
nor U14297 (N_14297,N_3104,N_2193);
nand U14298 (N_14298,N_411,N_3525);
nand U14299 (N_14299,N_9484,N_1940);
and U14300 (N_14300,N_1997,N_9207);
nand U14301 (N_14301,N_9445,N_5105);
or U14302 (N_14302,N_7730,N_4599);
or U14303 (N_14303,N_3457,N_80);
nand U14304 (N_14304,N_4016,N_7836);
nor U14305 (N_14305,N_6885,N_7564);
nor U14306 (N_14306,N_2309,N_830);
xor U14307 (N_14307,N_7935,N_5269);
or U14308 (N_14308,N_6876,N_1647);
nor U14309 (N_14309,N_7488,N_2818);
nand U14310 (N_14310,N_3794,N_6661);
and U14311 (N_14311,N_2101,N_3948);
or U14312 (N_14312,N_2337,N_3964);
and U14313 (N_14313,N_3306,N_2962);
and U14314 (N_14314,N_5548,N_7678);
xnor U14315 (N_14315,N_304,N_4211);
nor U14316 (N_14316,N_2120,N_2611);
or U14317 (N_14317,N_6546,N_1654);
nor U14318 (N_14318,N_3642,N_8119);
xor U14319 (N_14319,N_632,N_1882);
nor U14320 (N_14320,N_7234,N_6082);
nor U14321 (N_14321,N_255,N_8477);
nand U14322 (N_14322,N_7199,N_3332);
nand U14323 (N_14323,N_5759,N_9036);
or U14324 (N_14324,N_24,N_2940);
and U14325 (N_14325,N_8221,N_3904);
or U14326 (N_14326,N_839,N_7831);
nand U14327 (N_14327,N_9663,N_4232);
and U14328 (N_14328,N_3985,N_8337);
xor U14329 (N_14329,N_1241,N_6896);
xnor U14330 (N_14330,N_5868,N_5065);
xor U14331 (N_14331,N_2186,N_1474);
xor U14332 (N_14332,N_9179,N_6645);
nand U14333 (N_14333,N_8246,N_5704);
xnor U14334 (N_14334,N_1,N_2889);
nand U14335 (N_14335,N_4815,N_7333);
nor U14336 (N_14336,N_549,N_4676);
nor U14337 (N_14337,N_471,N_2026);
nor U14338 (N_14338,N_2440,N_511);
nor U14339 (N_14339,N_2434,N_3442);
xnor U14340 (N_14340,N_4516,N_2341);
xor U14341 (N_14341,N_9211,N_5514);
or U14342 (N_14342,N_3015,N_2631);
and U14343 (N_14343,N_8865,N_4885);
or U14344 (N_14344,N_2011,N_8928);
xnor U14345 (N_14345,N_2866,N_5165);
or U14346 (N_14346,N_3384,N_8392);
xor U14347 (N_14347,N_8334,N_8439);
nand U14348 (N_14348,N_4380,N_8763);
nor U14349 (N_14349,N_2949,N_9680);
or U14350 (N_14350,N_6601,N_2077);
and U14351 (N_14351,N_9624,N_6577);
nor U14352 (N_14352,N_4527,N_9122);
or U14353 (N_14353,N_5457,N_6489);
nand U14354 (N_14354,N_501,N_9808);
nand U14355 (N_14355,N_9565,N_9911);
nor U14356 (N_14356,N_9918,N_9553);
or U14357 (N_14357,N_5479,N_2435);
nor U14358 (N_14358,N_4553,N_2820);
nand U14359 (N_14359,N_9839,N_9250);
or U14360 (N_14360,N_3482,N_2696);
or U14361 (N_14361,N_9608,N_3325);
nand U14362 (N_14362,N_7641,N_9652);
or U14363 (N_14363,N_4046,N_3531);
nor U14364 (N_14364,N_7613,N_9780);
nand U14365 (N_14365,N_4222,N_7374);
nor U14366 (N_14366,N_1083,N_5282);
nand U14367 (N_14367,N_2308,N_2126);
or U14368 (N_14368,N_1655,N_3264);
nand U14369 (N_14369,N_8564,N_9627);
and U14370 (N_14370,N_8453,N_5403);
nand U14371 (N_14371,N_5320,N_583);
xor U14372 (N_14372,N_6194,N_7547);
xor U14373 (N_14373,N_4182,N_8488);
nor U14374 (N_14374,N_5771,N_5012);
nor U14375 (N_14375,N_8068,N_4916);
nand U14376 (N_14376,N_7068,N_7869);
nor U14377 (N_14377,N_4193,N_9165);
and U14378 (N_14378,N_7534,N_8923);
and U14379 (N_14379,N_8310,N_3371);
nor U14380 (N_14380,N_3988,N_1259);
nand U14381 (N_14381,N_8500,N_4883);
nor U14382 (N_14382,N_8196,N_9759);
nand U14383 (N_14383,N_9537,N_1960);
xnor U14384 (N_14384,N_344,N_9533);
nand U14385 (N_14385,N_3342,N_6203);
and U14386 (N_14386,N_1526,N_6003);
nor U14387 (N_14387,N_2780,N_2178);
nor U14388 (N_14388,N_961,N_8026);
or U14389 (N_14389,N_1098,N_981);
nand U14390 (N_14390,N_8062,N_1462);
and U14391 (N_14391,N_433,N_648);
nand U14392 (N_14392,N_3037,N_285);
or U14393 (N_14393,N_6793,N_2407);
nor U14394 (N_14394,N_5355,N_8314);
xnor U14395 (N_14395,N_757,N_1744);
nand U14396 (N_14396,N_5853,N_6975);
xnor U14397 (N_14397,N_6872,N_5799);
and U14398 (N_14398,N_9730,N_4149);
xnor U14399 (N_14399,N_2864,N_4903);
nand U14400 (N_14400,N_760,N_5929);
and U14401 (N_14401,N_5349,N_3910);
or U14402 (N_14402,N_3722,N_1145);
or U14403 (N_14403,N_8403,N_5615);
nand U14404 (N_14404,N_2640,N_6338);
or U14405 (N_14405,N_8947,N_5885);
nand U14406 (N_14406,N_2710,N_2745);
xor U14407 (N_14407,N_5737,N_6074);
nand U14408 (N_14408,N_6892,N_3340);
nor U14409 (N_14409,N_2132,N_6426);
xnor U14410 (N_14410,N_4735,N_9603);
xnor U14411 (N_14411,N_7619,N_8306);
nand U14412 (N_14412,N_6825,N_2947);
or U14413 (N_14413,N_6251,N_7864);
nand U14414 (N_14414,N_436,N_4510);
xor U14415 (N_14415,N_7162,N_678);
nand U14416 (N_14416,N_7169,N_9771);
nand U14417 (N_14417,N_4741,N_1921);
nand U14418 (N_14418,N_4069,N_8004);
nand U14419 (N_14419,N_1438,N_8971);
xnor U14420 (N_14420,N_4121,N_9602);
and U14421 (N_14421,N_7649,N_7030);
nor U14422 (N_14422,N_2354,N_3128);
xor U14423 (N_14423,N_7785,N_1380);
or U14424 (N_14424,N_3870,N_7357);
xnor U14425 (N_14425,N_2927,N_6365);
or U14426 (N_14426,N_7069,N_8727);
and U14427 (N_14427,N_2196,N_2701);
xnor U14428 (N_14428,N_2714,N_6008);
xor U14429 (N_14429,N_9885,N_64);
xor U14430 (N_14430,N_9436,N_4056);
or U14431 (N_14431,N_3594,N_9655);
and U14432 (N_14432,N_4632,N_8273);
and U14433 (N_14433,N_2248,N_7376);
nand U14434 (N_14434,N_3823,N_7345);
xnor U14435 (N_14435,N_457,N_2404);
and U14436 (N_14436,N_8720,N_392);
and U14437 (N_14437,N_2168,N_4203);
and U14438 (N_14438,N_195,N_4084);
or U14439 (N_14439,N_5942,N_3575);
xor U14440 (N_14440,N_8562,N_7540);
nand U14441 (N_14441,N_489,N_1906);
xor U14442 (N_14442,N_1724,N_3179);
nand U14443 (N_14443,N_3017,N_6109);
nand U14444 (N_14444,N_7666,N_7598);
nand U14445 (N_14445,N_9091,N_4482);
xnor U14446 (N_14446,N_3255,N_8625);
or U14447 (N_14447,N_1968,N_2607);
or U14448 (N_14448,N_6967,N_7617);
nor U14449 (N_14449,N_5745,N_8653);
and U14450 (N_14450,N_6442,N_8021);
nand U14451 (N_14451,N_5961,N_3211);
nand U14452 (N_14452,N_1844,N_3565);
xnor U14453 (N_14453,N_8095,N_2470);
or U14454 (N_14454,N_2551,N_5772);
nor U14455 (N_14455,N_6255,N_3559);
or U14456 (N_14456,N_8043,N_3866);
nor U14457 (N_14457,N_3348,N_3776);
nor U14458 (N_14458,N_7955,N_1043);
nor U14459 (N_14459,N_7642,N_1488);
or U14460 (N_14460,N_9852,N_7959);
xnor U14461 (N_14461,N_6895,N_7995);
and U14462 (N_14462,N_2867,N_740);
nor U14463 (N_14463,N_2092,N_3773);
nand U14464 (N_14464,N_3720,N_904);
nor U14465 (N_14465,N_1992,N_2854);
nor U14466 (N_14466,N_6374,N_7064);
and U14467 (N_14467,N_54,N_5513);
and U14468 (N_14468,N_958,N_4810);
nand U14469 (N_14469,N_1986,N_3226);
xnor U14470 (N_14470,N_8389,N_1902);
or U14471 (N_14471,N_6347,N_1794);
or U14472 (N_14472,N_3474,N_1878);
nor U14473 (N_14473,N_6283,N_6923);
and U14474 (N_14474,N_1406,N_8113);
nor U14475 (N_14475,N_4072,N_265);
or U14476 (N_14476,N_9103,N_7463);
xnor U14477 (N_14477,N_5361,N_2601);
nand U14478 (N_14478,N_2892,N_7240);
and U14479 (N_14479,N_3927,N_8638);
xor U14480 (N_14480,N_5409,N_5428);
nor U14481 (N_14481,N_4988,N_971);
and U14482 (N_14482,N_9017,N_1323);
xnor U14483 (N_14483,N_7276,N_1108);
and U14484 (N_14484,N_5982,N_2908);
and U14485 (N_14485,N_4141,N_4860);
xor U14486 (N_14486,N_2217,N_5819);
nand U14487 (N_14487,N_7422,N_1243);
nor U14488 (N_14488,N_2597,N_3256);
xor U14489 (N_14489,N_7954,N_1525);
nand U14490 (N_14490,N_9705,N_5404);
xor U14491 (N_14491,N_7839,N_5526);
xor U14492 (N_14492,N_9188,N_5228);
or U14493 (N_14493,N_6191,N_3085);
and U14494 (N_14494,N_8589,N_9703);
nand U14495 (N_14495,N_9937,N_9764);
and U14496 (N_14496,N_1449,N_1741);
nand U14497 (N_14497,N_694,N_7258);
and U14498 (N_14498,N_1850,N_8170);
and U14499 (N_14499,N_4788,N_4523);
or U14500 (N_14500,N_1283,N_1592);
nand U14501 (N_14501,N_6300,N_5541);
or U14502 (N_14502,N_449,N_3842);
and U14503 (N_14503,N_7081,N_7360);
and U14504 (N_14504,N_7184,N_9387);
xor U14505 (N_14505,N_2039,N_7078);
xnor U14506 (N_14506,N_1385,N_3883);
nand U14507 (N_14507,N_8996,N_9132);
xnor U14508 (N_14508,N_1841,N_6517);
and U14509 (N_14509,N_8455,N_2633);
nor U14510 (N_14510,N_1775,N_6075);
or U14511 (N_14511,N_2148,N_3399);
or U14512 (N_14512,N_1528,N_8206);
or U14513 (N_14513,N_1349,N_1814);
nand U14514 (N_14514,N_419,N_53);
and U14515 (N_14515,N_2034,N_9203);
or U14516 (N_14516,N_405,N_180);
nor U14517 (N_14517,N_2066,N_646);
xnor U14518 (N_14518,N_5277,N_887);
nor U14519 (N_14519,N_4035,N_2486);
xnor U14520 (N_14520,N_5053,N_5723);
and U14521 (N_14521,N_6840,N_3705);
xnor U14522 (N_14522,N_5563,N_8421);
xor U14523 (N_14523,N_9617,N_42);
xor U14524 (N_14524,N_8344,N_3650);
and U14525 (N_14525,N_2033,N_268);
or U14526 (N_14526,N_9300,N_2883);
nor U14527 (N_14527,N_3000,N_2083);
and U14528 (N_14528,N_9568,N_2363);
and U14529 (N_14529,N_8346,N_2849);
or U14530 (N_14530,N_8671,N_6334);
nor U14531 (N_14531,N_4890,N_910);
and U14532 (N_14532,N_8014,N_1862);
and U14533 (N_14533,N_5835,N_2042);
or U14534 (N_14534,N_7077,N_6623);
xor U14535 (N_14535,N_8662,N_9462);
nor U14536 (N_14536,N_9159,N_6799);
and U14537 (N_14537,N_5510,N_3993);
nand U14538 (N_14538,N_6532,N_4400);
nand U14539 (N_14539,N_9345,N_6148);
and U14540 (N_14540,N_2922,N_9748);
nor U14541 (N_14541,N_8293,N_8469);
and U14542 (N_14542,N_7508,N_9622);
or U14543 (N_14543,N_2321,N_804);
xnor U14544 (N_14544,N_4029,N_4915);
or U14545 (N_14545,N_3123,N_8710);
or U14546 (N_14546,N_1203,N_743);
or U14547 (N_14547,N_2317,N_6915);
nand U14548 (N_14548,N_2368,N_1572);
nor U14549 (N_14549,N_8385,N_1400);
or U14550 (N_14550,N_6641,N_3918);
xor U14551 (N_14551,N_6424,N_5584);
and U14552 (N_14552,N_4248,N_2930);
and U14553 (N_14553,N_8167,N_2988);
nor U14554 (N_14554,N_2382,N_1749);
xnor U14555 (N_14555,N_7362,N_2901);
nor U14556 (N_14556,N_6438,N_9660);
xor U14557 (N_14557,N_3819,N_3415);
nor U14558 (N_14558,N_1294,N_4820);
or U14559 (N_14559,N_8518,N_4234);
nor U14560 (N_14560,N_3611,N_9634);
nor U14561 (N_14561,N_1558,N_9479);
and U14562 (N_14562,N_837,N_3464);
nor U14563 (N_14563,N_3360,N_7554);
or U14564 (N_14564,N_2782,N_5701);
and U14565 (N_14565,N_6035,N_9751);
and U14566 (N_14566,N_5313,N_6152);
nor U14567 (N_14567,N_3620,N_7640);
or U14568 (N_14568,N_1761,N_3235);
nor U14569 (N_14569,N_7973,N_3865);
or U14570 (N_14570,N_8838,N_2692);
nor U14571 (N_14571,N_7107,N_2180);
or U14572 (N_14572,N_2358,N_2916);
nor U14573 (N_14573,N_2713,N_1699);
nand U14574 (N_14574,N_3376,N_3161);
nand U14575 (N_14575,N_3261,N_6478);
xnor U14576 (N_14576,N_9461,N_6952);
nor U14577 (N_14577,N_2900,N_6808);
or U14578 (N_14578,N_1369,N_5332);
or U14579 (N_14579,N_6488,N_1811);
or U14580 (N_14580,N_8580,N_2796);
or U14581 (N_14581,N_6716,N_3764);
nand U14582 (N_14582,N_1383,N_5311);
nor U14583 (N_14583,N_5213,N_7808);
nand U14584 (N_14584,N_2214,N_1760);
or U14585 (N_14585,N_4465,N_8818);
nand U14586 (N_14586,N_4216,N_2355);
nor U14587 (N_14587,N_1716,N_5650);
or U14588 (N_14588,N_5979,N_1138);
nand U14589 (N_14589,N_5398,N_5660);
nand U14590 (N_14590,N_5619,N_4062);
and U14591 (N_14591,N_1133,N_5924);
nor U14592 (N_14592,N_4414,N_4401);
or U14593 (N_14593,N_5777,N_5928);
nand U14594 (N_14594,N_5226,N_1517);
nor U14595 (N_14595,N_5291,N_9405);
xnor U14596 (N_14596,N_6686,N_6712);
or U14597 (N_14597,N_9607,N_1473);
and U14598 (N_14598,N_8325,N_508);
or U14599 (N_14599,N_5990,N_9797);
or U14600 (N_14600,N_6240,N_4700);
or U14601 (N_14601,N_5785,N_7414);
nand U14602 (N_14602,N_105,N_5661);
nor U14603 (N_14603,N_7636,N_1946);
xnor U14604 (N_14604,N_5960,N_4319);
and U14605 (N_14605,N_4804,N_6590);
xnor U14606 (N_14606,N_3676,N_1917);
or U14607 (N_14607,N_5538,N_5160);
xnor U14608 (N_14608,N_906,N_870);
or U14609 (N_14609,N_5973,N_1562);
or U14610 (N_14610,N_3027,N_9413);
xnor U14611 (N_14611,N_5156,N_812);
xnor U14612 (N_14612,N_5108,N_2756);
and U14613 (N_14613,N_718,N_5378);
xnor U14614 (N_14614,N_1812,N_3353);
nand U14615 (N_14615,N_7342,N_5664);
nor U14616 (N_14616,N_5429,N_2603);
nor U14617 (N_14617,N_5318,N_2801);
nor U14618 (N_14618,N_4161,N_3672);
and U14619 (N_14619,N_7269,N_8413);
nor U14620 (N_14620,N_9717,N_6371);
xor U14621 (N_14621,N_8010,N_3001);
nor U14622 (N_14622,N_8387,N_8635);
xor U14623 (N_14623,N_5059,N_7416);
nand U14624 (N_14624,N_4336,N_4452);
and U14625 (N_14625,N_7017,N_7757);
nor U14626 (N_14626,N_2029,N_1341);
xnor U14627 (N_14627,N_801,N_9059);
or U14628 (N_14628,N_5290,N_256);
xor U14629 (N_14629,N_9675,N_2855);
nor U14630 (N_14630,N_5983,N_7011);
nor U14631 (N_14631,N_3562,N_6779);
xnor U14632 (N_14632,N_7428,N_3835);
nor U14633 (N_14633,N_4743,N_2038);
nand U14634 (N_14634,N_2313,N_9403);
and U14635 (N_14635,N_5849,N_144);
or U14636 (N_14636,N_5817,N_3260);
and U14637 (N_14637,N_3759,N_7349);
or U14638 (N_14638,N_8981,N_2227);
and U14639 (N_14639,N_7651,N_5834);
and U14640 (N_14640,N_4698,N_3872);
xor U14641 (N_14641,N_3772,N_9545);
xnor U14642 (N_14642,N_1755,N_6217);
nor U14643 (N_14643,N_6407,N_28);
xnor U14644 (N_14644,N_7936,N_7753);
nand U14645 (N_14645,N_2736,N_5015);
or U14646 (N_14646,N_1097,N_184);
nor U14647 (N_14647,N_3815,N_5519);
and U14648 (N_14648,N_6183,N_7626);
nor U14649 (N_14649,N_1865,N_7024);
and U14650 (N_14650,N_9373,N_1834);
nand U14651 (N_14651,N_6973,N_3224);
or U14652 (N_14652,N_2682,N_6962);
xor U14653 (N_14653,N_1447,N_7140);
nor U14654 (N_14654,N_4674,N_1210);
xor U14655 (N_14655,N_2292,N_8128);
nand U14656 (N_14656,N_4823,N_4009);
nor U14657 (N_14657,N_5813,N_3956);
nand U14658 (N_14658,N_6483,N_6921);
nor U14659 (N_14659,N_6862,N_3021);
or U14660 (N_14660,N_7267,N_2099);
nor U14661 (N_14661,N_4487,N_3484);
nor U14662 (N_14662,N_9024,N_1624);
nor U14663 (N_14663,N_2372,N_7127);
and U14664 (N_14664,N_9047,N_350);
xnor U14665 (N_14665,N_5045,N_6022);
xnor U14666 (N_14666,N_2223,N_9707);
nand U14667 (N_14667,N_7809,N_435);
nor U14668 (N_14668,N_5689,N_581);
nand U14669 (N_14669,N_8624,N_8382);
nand U14670 (N_14670,N_5394,N_6117);
and U14671 (N_14671,N_5273,N_5118);
nor U14672 (N_14672,N_1886,N_7516);
nand U14673 (N_14673,N_4586,N_7957);
xor U14674 (N_14674,N_2725,N_3475);
nor U14675 (N_14675,N_7897,N_4776);
and U14676 (N_14676,N_982,N_7372);
and U14677 (N_14677,N_988,N_9787);
or U14678 (N_14678,N_3490,N_3390);
or U14679 (N_14679,N_4832,N_5678);
nand U14680 (N_14680,N_7926,N_7104);
nand U14681 (N_14681,N_734,N_927);
xor U14682 (N_14682,N_4963,N_8457);
and U14683 (N_14683,N_6246,N_1504);
xor U14684 (N_14684,N_1433,N_5167);
and U14685 (N_14685,N_8976,N_4806);
and U14686 (N_14686,N_1319,N_2873);
xnor U14687 (N_14687,N_2154,N_5286);
or U14688 (N_14688,N_4645,N_1011);
or U14689 (N_14689,N_9514,N_8723);
nand U14690 (N_14690,N_5271,N_3905);
nand U14691 (N_14691,N_6543,N_5920);
nand U14692 (N_14692,N_4006,N_3691);
nand U14693 (N_14693,N_6061,N_7476);
nand U14694 (N_14694,N_2198,N_329);
and U14695 (N_14695,N_8893,N_3046);
or U14696 (N_14696,N_2016,N_855);
nand U14697 (N_14697,N_4497,N_9061);
or U14698 (N_14698,N_3669,N_3992);
and U14699 (N_14699,N_6198,N_1949);
nor U14700 (N_14700,N_9161,N_3925);
and U14701 (N_14701,N_3936,N_8378);
nand U14702 (N_14702,N_7866,N_4877);
nand U14703 (N_14703,N_3162,N_8429);
xor U14704 (N_14704,N_143,N_8567);
nand U14705 (N_14705,N_4429,N_2944);
nor U14706 (N_14706,N_582,N_3252);
and U14707 (N_14707,N_286,N_3308);
nand U14708 (N_14708,N_2307,N_1873);
nor U14709 (N_14709,N_9140,N_5067);
or U14710 (N_14710,N_4966,N_7911);
or U14711 (N_14711,N_8952,N_1221);
nand U14712 (N_14712,N_6566,N_9898);
or U14713 (N_14713,N_5209,N_4620);
and U14714 (N_14714,N_4838,N_9371);
xnor U14715 (N_14715,N_7684,N_2110);
xor U14716 (N_14716,N_1614,N_7990);
nand U14717 (N_14717,N_5270,N_3677);
or U14718 (N_14718,N_3228,N_2813);
xor U14719 (N_14719,N_9916,N_4571);
nor U14720 (N_14720,N_8066,N_7265);
or U14721 (N_14721,N_8586,N_8787);
and U14722 (N_14722,N_1284,N_2583);
or U14723 (N_14723,N_9303,N_902);
or U14724 (N_14724,N_8179,N_5422);
xor U14725 (N_14725,N_8828,N_5956);
xnor U14726 (N_14726,N_3220,N_9697);
nor U14727 (N_14727,N_2816,N_1033);
or U14728 (N_14728,N_2559,N_6678);
nand U14729 (N_14729,N_9286,N_3397);
nor U14730 (N_14730,N_989,N_9465);
and U14731 (N_14731,N_7632,N_2552);
and U14732 (N_14732,N_6366,N_2304);
or U14733 (N_14733,N_4267,N_5803);
or U14734 (N_14734,N_5280,N_1767);
xor U14735 (N_14735,N_4054,N_9804);
or U14736 (N_14736,N_6,N_2795);
and U14737 (N_14737,N_7287,N_7125);
nand U14738 (N_14738,N_703,N_2393);
nor U14739 (N_14739,N_6520,N_5178);
xor U14740 (N_14740,N_5625,N_1970);
nor U14741 (N_14741,N_7919,N_4873);
or U14742 (N_14742,N_1331,N_5305);
nor U14743 (N_14743,N_4926,N_2102);
nand U14744 (N_14744,N_2520,N_4944);
or U14745 (N_14745,N_3434,N_6038);
nand U14746 (N_14746,N_3626,N_4833);
nand U14747 (N_14747,N_921,N_6391);
and U14748 (N_14748,N_7967,N_1728);
nand U14749 (N_14749,N_677,N_5446);
and U14750 (N_14750,N_4505,N_5521);
or U14751 (N_14751,N_9960,N_3903);
nor U14752 (N_14752,N_4812,N_5216);
nor U14753 (N_14753,N_1690,N_5109);
or U14754 (N_14754,N_6215,N_3445);
and U14755 (N_14755,N_6412,N_7029);
nand U14756 (N_14756,N_170,N_8445);
nand U14757 (N_14757,N_2753,N_2708);
nand U14758 (N_14758,N_1681,N_4958);
nand U14759 (N_14759,N_7365,N_6909);
nand U14760 (N_14760,N_5388,N_4655);
nor U14761 (N_14761,N_5125,N_9813);
nand U14762 (N_14762,N_8125,N_6466);
nand U14763 (N_14763,N_8700,N_4020);
and U14764 (N_14764,N_652,N_6070);
nor U14765 (N_14765,N_2349,N_3109);
or U14766 (N_14766,N_9613,N_3724);
xor U14767 (N_14767,N_9679,N_8190);
xor U14768 (N_14768,N_2022,N_5029);
xnor U14769 (N_14769,N_5636,N_3294);
nor U14770 (N_14770,N_4657,N_10);
xnor U14771 (N_14771,N_2732,N_4454);
nor U14772 (N_14772,N_8909,N_8270);
nor U14773 (N_14773,N_5114,N_2799);
nand U14774 (N_14774,N_1074,N_2318);
or U14775 (N_14775,N_192,N_7243);
or U14776 (N_14776,N_6046,N_5076);
xnor U14777 (N_14777,N_6304,N_7072);
nand U14778 (N_14778,N_8536,N_8595);
and U14779 (N_14779,N_1904,N_9658);
xnor U14780 (N_14780,N_6067,N_5902);
and U14781 (N_14781,N_421,N_9055);
and U14782 (N_14782,N_2162,N_5169);
xor U14783 (N_14783,N_6908,N_4540);
nor U14784 (N_14784,N_8644,N_7882);
xnor U14785 (N_14785,N_9367,N_8163);
xor U14786 (N_14786,N_3949,N_848);
or U14787 (N_14787,N_7344,N_1847);
xor U14788 (N_14788,N_7235,N_2386);
nand U14789 (N_14789,N_9244,N_7562);
xnor U14790 (N_14790,N_4836,N_5797);
xnor U14791 (N_14791,N_5626,N_9791);
nor U14792 (N_14792,N_8549,N_7538);
nor U14793 (N_14793,N_9815,N_1051);
xor U14794 (N_14794,N_3222,N_7094);
or U14795 (N_14795,N_7509,N_9476);
and U14796 (N_14796,N_9323,N_7100);
nor U14797 (N_14797,N_7971,N_3718);
xnor U14798 (N_14798,N_2972,N_2053);
nand U14799 (N_14799,N_7096,N_7208);
or U14800 (N_14800,N_6766,N_6837);
xor U14801 (N_14801,N_9871,N_7281);
xor U14802 (N_14802,N_6721,N_1952);
xor U14803 (N_14803,N_992,N_9620);
and U14804 (N_14804,N_5370,N_7105);
and U14805 (N_14805,N_1309,N_4757);
nand U14806 (N_14806,N_563,N_5205);
or U14807 (N_14807,N_8848,N_5072);
xor U14808 (N_14808,N_5185,N_6262);
and U14809 (N_14809,N_5789,N_7331);
nand U14810 (N_14810,N_9406,N_3837);
and U14811 (N_14811,N_974,N_4439);
nand U14812 (N_14812,N_9420,N_7359);
nand U14813 (N_14813,N_1553,N_2851);
or U14814 (N_14814,N_5485,N_3719);
or U14815 (N_14815,N_3788,N_9569);
xor U14816 (N_14816,N_8730,N_8173);
xor U14817 (N_14817,N_5993,N_3113);
nor U14818 (N_14818,N_5353,N_5096);
and U14819 (N_14819,N_5447,N_8917);
nand U14820 (N_14820,N_551,N_4766);
nor U14821 (N_14821,N_4872,N_3063);
or U14822 (N_14822,N_9246,N_9876);
or U14823 (N_14823,N_2485,N_818);
and U14824 (N_14824,N_5441,N_2087);
nand U14825 (N_14825,N_214,N_0);
and U14826 (N_14826,N_5189,N_2236);
nor U14827 (N_14827,N_7303,N_1119);
or U14828 (N_14828,N_2546,N_8916);
nor U14829 (N_14829,N_3666,N_456);
xnor U14830 (N_14830,N_8092,N_1451);
or U14831 (N_14831,N_866,N_2623);
and U14832 (N_14832,N_654,N_9168);
nand U14833 (N_14833,N_4905,N_3693);
nor U14834 (N_14834,N_1698,N_8661);
or U14835 (N_14835,N_9350,N_2086);
or U14836 (N_14836,N_9372,N_5782);
and U14837 (N_14837,N_5116,N_5758);
or U14838 (N_14838,N_5483,N_4739);
and U14839 (N_14839,N_6689,N_4712);
or U14840 (N_14840,N_4722,N_613);
nand U14841 (N_14841,N_4332,N_5775);
nor U14842 (N_14842,N_7603,N_7608);
and U14843 (N_14843,N_3580,N_1912);
or U14844 (N_14844,N_277,N_7202);
xnor U14845 (N_14845,N_6397,N_2757);
and U14846 (N_14846,N_7283,N_8965);
or U14847 (N_14847,N_3418,N_5555);
nand U14848 (N_14848,N_6258,N_1443);
or U14849 (N_14849,N_4909,N_8091);
and U14850 (N_14850,N_4870,N_7400);
nand U14851 (N_14851,N_2370,N_2723);
xor U14852 (N_14852,N_1802,N_288);
nand U14853 (N_14853,N_4078,N_7391);
nor U14854 (N_14854,N_1807,N_3078);
nand U14855 (N_14855,N_3156,N_9944);
and U14856 (N_14856,N_3164,N_19);
xnor U14857 (N_14857,N_130,N_169);
nor U14858 (N_14858,N_6970,N_3994);
xor U14859 (N_14859,N_4310,N_8729);
or U14860 (N_14860,N_2578,N_6309);
xor U14861 (N_14861,N_2207,N_3486);
xor U14862 (N_14862,N_30,N_4552);
xor U14863 (N_14863,N_3116,N_1925);
or U14864 (N_14864,N_5654,N_7887);
nand U14865 (N_14865,N_4430,N_8006);
nand U14866 (N_14866,N_7587,N_8774);
or U14867 (N_14867,N_8576,N_6273);
and U14868 (N_14868,N_5391,N_5224);
nand U14869 (N_14869,N_2251,N_8491);
or U14870 (N_14870,N_7650,N_5336);
xnor U14871 (N_14871,N_8939,N_3243);
and U14872 (N_14872,N_7005,N_1644);
or U14873 (N_14873,N_7758,N_9112);
or U14874 (N_14874,N_1464,N_729);
or U14875 (N_14875,N_4003,N_6615);
xor U14876 (N_14876,N_3048,N_2897);
or U14877 (N_14877,N_6446,N_8105);
nor U14878 (N_14878,N_3005,N_5095);
and U14879 (N_14879,N_3527,N_687);
and U14880 (N_14880,N_1014,N_6639);
nor U14881 (N_14881,N_8575,N_3577);
xnor U14882 (N_14882,N_3265,N_9423);
nor U14883 (N_14883,N_7167,N_9424);
nor U14884 (N_14884,N_2697,N_6740);
nor U14885 (N_14885,N_884,N_2657);
nor U14886 (N_14886,N_2977,N_7531);
xor U14887 (N_14887,N_5448,N_7225);
xor U14888 (N_14888,N_3209,N_4048);
xnor U14889 (N_14889,N_1280,N_6932);
xor U14890 (N_14890,N_6672,N_713);
and U14891 (N_14891,N_2828,N_6051);
nor U14892 (N_14892,N_9404,N_6389);
nor U14893 (N_14893,N_4986,N_4642);
xnor U14894 (N_14894,N_968,N_7040);
and U14895 (N_14895,N_3641,N_5363);
nand U14896 (N_14896,N_2389,N_8046);
nand U14897 (N_14897,N_2931,N_7458);
or U14898 (N_14898,N_3685,N_1496);
and U14899 (N_14899,N_627,N_7004);
nor U14900 (N_14900,N_4318,N_231);
xor U14901 (N_14901,N_2426,N_4356);
nor U14902 (N_14902,N_8824,N_6320);
nand U14903 (N_14903,N_7293,N_3076);
xnor U14904 (N_14904,N_7740,N_14);
nor U14905 (N_14905,N_8659,N_6002);
xor U14906 (N_14906,N_5570,N_7686);
nand U14907 (N_14907,N_6387,N_1835);
xor U14908 (N_14908,N_3963,N_886);
nor U14909 (N_14909,N_8820,N_1261);
nor U14910 (N_14910,N_9376,N_3020);
nor U14911 (N_14911,N_2433,N_4563);
nor U14912 (N_14912,N_4102,N_354);
xnor U14913 (N_14913,N_8048,N_2188);
or U14914 (N_14914,N_1478,N_9737);
xor U14915 (N_14915,N_5784,N_7595);
nand U14916 (N_14916,N_4948,N_3678);
nand U14917 (N_14917,N_2473,N_3646);
xnor U14918 (N_14918,N_7120,N_3311);
or U14919 (N_14919,N_5594,N_6416);
nor U14920 (N_14920,N_1050,N_699);
nor U14921 (N_14921,N_4785,N_6010);
nor U14922 (N_14922,N_4321,N_2109);
nand U14923 (N_14923,N_3030,N_8188);
xor U14924 (N_14924,N_9879,N_3827);
or U14925 (N_14925,N_7,N_8353);
and U14926 (N_14926,N_595,N_3354);
or U14927 (N_14927,N_7943,N_5098);
or U14928 (N_14928,N_9009,N_8689);
nand U14929 (N_14929,N_8742,N_4033);
or U14930 (N_14930,N_793,N_3285);
nor U14931 (N_14931,N_7504,N_1956);
nor U14932 (N_14932,N_1091,N_755);
nand U14933 (N_14933,N_3545,N_9243);
nand U14934 (N_14934,N_8481,N_8785);
or U14935 (N_14935,N_9147,N_4286);
nand U14936 (N_14936,N_444,N_5234);
xor U14937 (N_14937,N_4477,N_9080);
nor U14938 (N_14938,N_6058,N_5005);
nor U14939 (N_14939,N_2945,N_9783);
and U14940 (N_14940,N_1392,N_3753);
xnor U14941 (N_14941,N_8134,N_3034);
nand U14942 (N_14942,N_3031,N_2943);
xnor U14943 (N_14943,N_8416,N_1084);
nor U14944 (N_14944,N_41,N_4608);
nor U14945 (N_14945,N_6619,N_4204);
and U14946 (N_14946,N_4119,N_7947);
nand U14947 (N_14947,N_7648,N_4728);
nand U14948 (N_14948,N_9355,N_9645);
nand U14949 (N_14949,N_3272,N_8238);
nand U14950 (N_14950,N_1156,N_9531);
nand U14951 (N_14951,N_1608,N_4710);
and U14952 (N_14952,N_3711,N_4277);
or U14953 (N_14953,N_3506,N_5670);
nand U14954 (N_14954,N_8957,N_2289);
and U14955 (N_14955,N_690,N_3387);
nand U14956 (N_14956,N_7305,N_8639);
nand U14957 (N_14957,N_1733,N_808);
nand U14958 (N_14958,N_5812,N_8890);
and U14959 (N_14959,N_3362,N_5852);
nor U14960 (N_14960,N_7687,N_2478);
nand U14961 (N_14961,N_4041,N_4460);
nand U14962 (N_14962,N_1332,N_576);
nand U14963 (N_14963,N_2491,N_3824);
or U14964 (N_14964,N_6156,N_150);
nand U14965 (N_14965,N_9408,N_7157);
or U14966 (N_14966,N_7280,N_1797);
xnor U14967 (N_14967,N_5470,N_2417);
nor U14968 (N_14968,N_8426,N_1493);
and U14969 (N_14969,N_1310,N_5431);
xor U14970 (N_14970,N_2581,N_7794);
xor U14971 (N_14971,N_8281,N_281);
or U14972 (N_14972,N_9214,N_347);
nor U14973 (N_14973,N_9253,N_4413);
and U14974 (N_14974,N_6116,N_1801);
and U14975 (N_14975,N_1737,N_1818);
xnor U14976 (N_14976,N_4522,N_5348);
or U14977 (N_14977,N_2859,N_5693);
nand U14978 (N_14978,N_9271,N_3321);
and U14979 (N_14979,N_6733,N_6745);
and U14980 (N_14980,N_6170,N_35);
or U14981 (N_14981,N_2079,N_671);
and U14982 (N_14982,N_9688,N_499);
or U14983 (N_14983,N_9030,N_2655);
nor U14984 (N_14984,N_4580,N_9768);
nand U14985 (N_14985,N_4243,N_7164);
xnor U14986 (N_14986,N_9837,N_1530);
and U14987 (N_14987,N_6664,N_8513);
xor U14988 (N_14988,N_1597,N_4174);
and U14989 (N_14989,N_9040,N_947);
and U14990 (N_14990,N_3137,N_9859);
xor U14991 (N_14991,N_9761,N_934);
nor U14992 (N_14992,N_138,N_5972);
nor U14993 (N_14993,N_8279,N_4155);
nor U14994 (N_14994,N_8627,N_1692);
xnor U14995 (N_14995,N_4,N_8404);
xnor U14996 (N_14996,N_8507,N_1622);
and U14997 (N_14997,N_6052,N_6367);
and U14998 (N_14998,N_8869,N_8166);
or U14999 (N_14999,N_9396,N_767);
or U15000 (N_15000,N_2954,N_1898);
and U15001 (N_15001,N_2920,N_5085);
nand U15002 (N_15002,N_4402,N_77);
or U15003 (N_15003,N_6264,N_6783);
or U15004 (N_15004,N_5219,N_1897);
nand U15005 (N_15005,N_5843,N_4202);
and U15006 (N_15006,N_4590,N_1121);
or U15007 (N_15007,N_1757,N_1085);
nor U15008 (N_15008,N_6433,N_6836);
or U15009 (N_15009,N_5193,N_537);
and U15010 (N_15010,N_8178,N_9051);
xnor U15011 (N_15011,N_2696,N_9536);
nand U15012 (N_15012,N_7799,N_4662);
xor U15013 (N_15013,N_6152,N_8491);
nand U15014 (N_15014,N_5558,N_1455);
xor U15015 (N_15015,N_9597,N_8297);
or U15016 (N_15016,N_2257,N_9791);
xnor U15017 (N_15017,N_1543,N_3628);
nor U15018 (N_15018,N_7498,N_6528);
or U15019 (N_15019,N_8941,N_6223);
or U15020 (N_15020,N_9432,N_7180);
and U15021 (N_15021,N_3309,N_6826);
or U15022 (N_15022,N_7012,N_3418);
nor U15023 (N_15023,N_4277,N_462);
or U15024 (N_15024,N_6740,N_3204);
nor U15025 (N_15025,N_7398,N_8292);
nand U15026 (N_15026,N_9823,N_7627);
xnor U15027 (N_15027,N_3432,N_8659);
nand U15028 (N_15028,N_1815,N_699);
nand U15029 (N_15029,N_1439,N_3173);
or U15030 (N_15030,N_5788,N_7750);
xnor U15031 (N_15031,N_1973,N_8045);
and U15032 (N_15032,N_3876,N_4882);
nand U15033 (N_15033,N_8719,N_9444);
nand U15034 (N_15034,N_2647,N_616);
xnor U15035 (N_15035,N_6757,N_634);
and U15036 (N_15036,N_305,N_2754);
xnor U15037 (N_15037,N_1356,N_675);
nand U15038 (N_15038,N_207,N_2724);
nand U15039 (N_15039,N_264,N_3140);
and U15040 (N_15040,N_4990,N_1842);
nor U15041 (N_15041,N_3771,N_7707);
and U15042 (N_15042,N_6201,N_9333);
xnor U15043 (N_15043,N_42,N_2902);
nand U15044 (N_15044,N_6701,N_6658);
nand U15045 (N_15045,N_3849,N_3625);
nor U15046 (N_15046,N_388,N_5643);
nand U15047 (N_15047,N_1395,N_7344);
nand U15048 (N_15048,N_4403,N_3484);
and U15049 (N_15049,N_3286,N_5011);
and U15050 (N_15050,N_8800,N_849);
and U15051 (N_15051,N_1575,N_5131);
or U15052 (N_15052,N_5959,N_9045);
and U15053 (N_15053,N_3277,N_9445);
and U15054 (N_15054,N_4863,N_5650);
nand U15055 (N_15055,N_9239,N_1014);
nor U15056 (N_15056,N_7700,N_9238);
and U15057 (N_15057,N_3161,N_7267);
or U15058 (N_15058,N_3787,N_3428);
and U15059 (N_15059,N_5584,N_9777);
or U15060 (N_15060,N_562,N_8555);
xor U15061 (N_15061,N_9387,N_6654);
xor U15062 (N_15062,N_3227,N_9010);
xor U15063 (N_15063,N_776,N_7734);
nor U15064 (N_15064,N_1830,N_9551);
nand U15065 (N_15065,N_81,N_2585);
or U15066 (N_15066,N_224,N_4789);
nor U15067 (N_15067,N_1186,N_6746);
or U15068 (N_15068,N_9616,N_7045);
and U15069 (N_15069,N_4360,N_1138);
nand U15070 (N_15070,N_3665,N_5803);
and U15071 (N_15071,N_4127,N_8393);
and U15072 (N_15072,N_6989,N_4328);
and U15073 (N_15073,N_4669,N_5460);
nor U15074 (N_15074,N_9464,N_3391);
nand U15075 (N_15075,N_6977,N_8830);
nor U15076 (N_15076,N_9661,N_3013);
or U15077 (N_15077,N_4513,N_6412);
nand U15078 (N_15078,N_2505,N_2337);
nand U15079 (N_15079,N_4748,N_720);
nor U15080 (N_15080,N_9847,N_2395);
and U15081 (N_15081,N_4111,N_2344);
nor U15082 (N_15082,N_9138,N_206);
nand U15083 (N_15083,N_9610,N_7406);
and U15084 (N_15084,N_1134,N_9100);
nor U15085 (N_15085,N_8797,N_1890);
nor U15086 (N_15086,N_5222,N_6902);
and U15087 (N_15087,N_3649,N_7348);
or U15088 (N_15088,N_2129,N_2562);
xor U15089 (N_15089,N_8389,N_6173);
nand U15090 (N_15090,N_8475,N_1938);
xnor U15091 (N_15091,N_8377,N_4702);
and U15092 (N_15092,N_1022,N_7697);
and U15093 (N_15093,N_1285,N_7133);
and U15094 (N_15094,N_7638,N_6054);
nor U15095 (N_15095,N_9097,N_661);
and U15096 (N_15096,N_6873,N_3602);
xor U15097 (N_15097,N_6781,N_3477);
and U15098 (N_15098,N_1484,N_8153);
xnor U15099 (N_15099,N_774,N_6119);
nand U15100 (N_15100,N_7421,N_7567);
nor U15101 (N_15101,N_7392,N_42);
nand U15102 (N_15102,N_5880,N_9812);
xnor U15103 (N_15103,N_8760,N_7232);
nand U15104 (N_15104,N_9070,N_4451);
or U15105 (N_15105,N_1222,N_7206);
or U15106 (N_15106,N_2795,N_7503);
or U15107 (N_15107,N_4568,N_2119);
nand U15108 (N_15108,N_8459,N_5589);
nand U15109 (N_15109,N_4564,N_7711);
and U15110 (N_15110,N_4001,N_2211);
nand U15111 (N_15111,N_7684,N_4050);
nor U15112 (N_15112,N_9922,N_2006);
and U15113 (N_15113,N_3418,N_1228);
nor U15114 (N_15114,N_2450,N_887);
or U15115 (N_15115,N_3569,N_1927);
xor U15116 (N_15116,N_8273,N_682);
or U15117 (N_15117,N_1095,N_8493);
nor U15118 (N_15118,N_2512,N_4890);
xor U15119 (N_15119,N_2521,N_3609);
nand U15120 (N_15120,N_3814,N_3158);
xor U15121 (N_15121,N_7299,N_3044);
nor U15122 (N_15122,N_8704,N_6919);
or U15123 (N_15123,N_8805,N_8679);
nand U15124 (N_15124,N_3842,N_2712);
and U15125 (N_15125,N_5630,N_6498);
and U15126 (N_15126,N_8049,N_5116);
or U15127 (N_15127,N_6096,N_4505);
xnor U15128 (N_15128,N_9603,N_9345);
xnor U15129 (N_15129,N_3772,N_9041);
xor U15130 (N_15130,N_552,N_902);
nor U15131 (N_15131,N_6763,N_2053);
or U15132 (N_15132,N_1108,N_3785);
nor U15133 (N_15133,N_2646,N_91);
nor U15134 (N_15134,N_733,N_7183);
nand U15135 (N_15135,N_6583,N_1150);
or U15136 (N_15136,N_8461,N_8957);
nand U15137 (N_15137,N_6816,N_5421);
nand U15138 (N_15138,N_810,N_219);
nand U15139 (N_15139,N_6365,N_2473);
and U15140 (N_15140,N_9920,N_2656);
or U15141 (N_15141,N_684,N_9237);
xor U15142 (N_15142,N_7575,N_8794);
nand U15143 (N_15143,N_2253,N_5152);
nand U15144 (N_15144,N_2548,N_3938);
nand U15145 (N_15145,N_9478,N_6196);
nand U15146 (N_15146,N_8439,N_8676);
and U15147 (N_15147,N_6171,N_4988);
or U15148 (N_15148,N_5327,N_7302);
nor U15149 (N_15149,N_4407,N_3234);
and U15150 (N_15150,N_1259,N_1802);
nand U15151 (N_15151,N_5691,N_5720);
nand U15152 (N_15152,N_8744,N_3973);
or U15153 (N_15153,N_6765,N_2063);
nand U15154 (N_15154,N_3891,N_7624);
nor U15155 (N_15155,N_1853,N_8574);
xnor U15156 (N_15156,N_7207,N_7050);
nand U15157 (N_15157,N_3098,N_4486);
nand U15158 (N_15158,N_8656,N_6635);
xor U15159 (N_15159,N_9187,N_4340);
xor U15160 (N_15160,N_5422,N_163);
and U15161 (N_15161,N_7251,N_323);
and U15162 (N_15162,N_6275,N_9125);
and U15163 (N_15163,N_8864,N_2332);
nor U15164 (N_15164,N_8319,N_2894);
or U15165 (N_15165,N_5401,N_2111);
or U15166 (N_15166,N_2561,N_132);
xor U15167 (N_15167,N_2129,N_3918);
xnor U15168 (N_15168,N_8979,N_5634);
and U15169 (N_15169,N_3010,N_1490);
xor U15170 (N_15170,N_9375,N_6025);
nand U15171 (N_15171,N_7442,N_3654);
nand U15172 (N_15172,N_9720,N_8747);
nand U15173 (N_15173,N_8392,N_2939);
xor U15174 (N_15174,N_1557,N_8167);
nor U15175 (N_15175,N_7544,N_1485);
or U15176 (N_15176,N_3215,N_3547);
and U15177 (N_15177,N_6825,N_3733);
and U15178 (N_15178,N_6595,N_4700);
and U15179 (N_15179,N_3316,N_7449);
nor U15180 (N_15180,N_1223,N_6091);
or U15181 (N_15181,N_8193,N_4035);
and U15182 (N_15182,N_5566,N_5435);
nor U15183 (N_15183,N_3538,N_9425);
and U15184 (N_15184,N_7486,N_923);
xnor U15185 (N_15185,N_3822,N_8619);
nand U15186 (N_15186,N_4329,N_3318);
nor U15187 (N_15187,N_4661,N_5113);
nand U15188 (N_15188,N_4874,N_2661);
nor U15189 (N_15189,N_4863,N_3625);
and U15190 (N_15190,N_2365,N_9214);
nor U15191 (N_15191,N_6017,N_6679);
and U15192 (N_15192,N_3078,N_8554);
xnor U15193 (N_15193,N_7117,N_4526);
or U15194 (N_15194,N_4576,N_5550);
nand U15195 (N_15195,N_8427,N_7641);
xnor U15196 (N_15196,N_2419,N_4936);
and U15197 (N_15197,N_4121,N_3558);
and U15198 (N_15198,N_4178,N_7766);
and U15199 (N_15199,N_1257,N_4183);
or U15200 (N_15200,N_590,N_6566);
and U15201 (N_15201,N_8496,N_9642);
and U15202 (N_15202,N_8888,N_5828);
nand U15203 (N_15203,N_7570,N_454);
or U15204 (N_15204,N_7539,N_7374);
xnor U15205 (N_15205,N_7262,N_7650);
nand U15206 (N_15206,N_337,N_4881);
or U15207 (N_15207,N_4950,N_289);
and U15208 (N_15208,N_2622,N_6610);
nor U15209 (N_15209,N_3859,N_633);
nor U15210 (N_15210,N_3982,N_7018);
nand U15211 (N_15211,N_8485,N_1746);
xnor U15212 (N_15212,N_1969,N_786);
nand U15213 (N_15213,N_4680,N_5978);
nor U15214 (N_15214,N_1688,N_1809);
xor U15215 (N_15215,N_4375,N_994);
and U15216 (N_15216,N_3137,N_7409);
nor U15217 (N_15217,N_401,N_7856);
nand U15218 (N_15218,N_6665,N_1122);
or U15219 (N_15219,N_2250,N_8402);
and U15220 (N_15220,N_404,N_221);
nor U15221 (N_15221,N_3404,N_1828);
nand U15222 (N_15222,N_7432,N_1001);
xnor U15223 (N_15223,N_3705,N_2112);
and U15224 (N_15224,N_1866,N_6268);
or U15225 (N_15225,N_7800,N_1424);
xnor U15226 (N_15226,N_9028,N_8174);
and U15227 (N_15227,N_241,N_2214);
xnor U15228 (N_15228,N_8001,N_8305);
and U15229 (N_15229,N_1302,N_5597);
nor U15230 (N_15230,N_1029,N_944);
nor U15231 (N_15231,N_9052,N_8118);
xor U15232 (N_15232,N_9227,N_9256);
or U15233 (N_15233,N_2564,N_1102);
xnor U15234 (N_15234,N_3938,N_8815);
nand U15235 (N_15235,N_8373,N_3242);
nor U15236 (N_15236,N_3202,N_4742);
nor U15237 (N_15237,N_9830,N_4449);
nor U15238 (N_15238,N_1842,N_4447);
or U15239 (N_15239,N_8082,N_9621);
and U15240 (N_15240,N_4867,N_812);
and U15241 (N_15241,N_3604,N_3775);
xnor U15242 (N_15242,N_4052,N_4995);
or U15243 (N_15243,N_62,N_1808);
nand U15244 (N_15244,N_4718,N_7467);
and U15245 (N_15245,N_3880,N_2818);
or U15246 (N_15246,N_8618,N_2670);
nor U15247 (N_15247,N_5552,N_3495);
nor U15248 (N_15248,N_4713,N_8936);
nor U15249 (N_15249,N_3757,N_851);
nor U15250 (N_15250,N_4990,N_3241);
xor U15251 (N_15251,N_2440,N_1742);
xnor U15252 (N_15252,N_5969,N_8547);
and U15253 (N_15253,N_5481,N_5725);
nor U15254 (N_15254,N_5296,N_6743);
and U15255 (N_15255,N_1605,N_1937);
nand U15256 (N_15256,N_4538,N_2908);
nand U15257 (N_15257,N_7193,N_8611);
nor U15258 (N_15258,N_3666,N_3395);
xnor U15259 (N_15259,N_4856,N_7706);
nand U15260 (N_15260,N_7232,N_1160);
and U15261 (N_15261,N_115,N_5514);
nand U15262 (N_15262,N_9159,N_8798);
nor U15263 (N_15263,N_9533,N_9613);
and U15264 (N_15264,N_6427,N_7719);
xor U15265 (N_15265,N_3194,N_3338);
and U15266 (N_15266,N_7938,N_5060);
and U15267 (N_15267,N_8465,N_9120);
nand U15268 (N_15268,N_1918,N_3740);
nor U15269 (N_15269,N_648,N_4769);
nor U15270 (N_15270,N_864,N_3598);
or U15271 (N_15271,N_978,N_2953);
or U15272 (N_15272,N_8200,N_5541);
or U15273 (N_15273,N_2807,N_2697);
nor U15274 (N_15274,N_6064,N_9647);
nand U15275 (N_15275,N_2963,N_3365);
or U15276 (N_15276,N_9366,N_6217);
xor U15277 (N_15277,N_8034,N_7233);
or U15278 (N_15278,N_8215,N_5005);
nand U15279 (N_15279,N_5518,N_4684);
xnor U15280 (N_15280,N_4672,N_9559);
and U15281 (N_15281,N_8198,N_989);
nor U15282 (N_15282,N_1007,N_8096);
nor U15283 (N_15283,N_9672,N_8673);
nor U15284 (N_15284,N_6309,N_5442);
and U15285 (N_15285,N_3714,N_833);
and U15286 (N_15286,N_4877,N_626);
xor U15287 (N_15287,N_2913,N_3700);
nand U15288 (N_15288,N_4509,N_7381);
or U15289 (N_15289,N_3601,N_8434);
nor U15290 (N_15290,N_818,N_3507);
and U15291 (N_15291,N_6139,N_4637);
and U15292 (N_15292,N_6005,N_9384);
nor U15293 (N_15293,N_5530,N_5228);
nand U15294 (N_15294,N_3575,N_3932);
or U15295 (N_15295,N_5526,N_130);
nand U15296 (N_15296,N_1649,N_5550);
or U15297 (N_15297,N_8863,N_2555);
or U15298 (N_15298,N_4875,N_6174);
nand U15299 (N_15299,N_4207,N_9224);
xnor U15300 (N_15300,N_3963,N_2833);
or U15301 (N_15301,N_8772,N_1941);
or U15302 (N_15302,N_8948,N_2633);
nand U15303 (N_15303,N_68,N_4282);
or U15304 (N_15304,N_8234,N_8015);
or U15305 (N_15305,N_7082,N_2028);
nand U15306 (N_15306,N_9576,N_3467);
or U15307 (N_15307,N_5579,N_7512);
xor U15308 (N_15308,N_7588,N_1493);
and U15309 (N_15309,N_5893,N_4494);
nand U15310 (N_15310,N_1436,N_9167);
xnor U15311 (N_15311,N_5615,N_5303);
or U15312 (N_15312,N_1890,N_7682);
or U15313 (N_15313,N_7076,N_4733);
nor U15314 (N_15314,N_2179,N_335);
xnor U15315 (N_15315,N_3725,N_3655);
and U15316 (N_15316,N_293,N_1668);
nor U15317 (N_15317,N_6461,N_4007);
or U15318 (N_15318,N_178,N_8632);
xor U15319 (N_15319,N_4686,N_2746);
and U15320 (N_15320,N_3106,N_8813);
nand U15321 (N_15321,N_244,N_6320);
nand U15322 (N_15322,N_2382,N_6515);
and U15323 (N_15323,N_7164,N_9006);
and U15324 (N_15324,N_2718,N_4764);
and U15325 (N_15325,N_1185,N_3455);
xnor U15326 (N_15326,N_7417,N_9023);
nand U15327 (N_15327,N_4165,N_170);
and U15328 (N_15328,N_9411,N_9515);
or U15329 (N_15329,N_812,N_211);
xor U15330 (N_15330,N_4434,N_7623);
nand U15331 (N_15331,N_3655,N_9615);
and U15332 (N_15332,N_7892,N_1359);
nor U15333 (N_15333,N_675,N_3265);
nor U15334 (N_15334,N_1132,N_827);
or U15335 (N_15335,N_2762,N_3223);
nand U15336 (N_15336,N_5450,N_2329);
and U15337 (N_15337,N_2595,N_3479);
and U15338 (N_15338,N_3899,N_464);
nor U15339 (N_15339,N_3516,N_6454);
nor U15340 (N_15340,N_920,N_6525);
and U15341 (N_15341,N_1736,N_3613);
xnor U15342 (N_15342,N_2074,N_6324);
xor U15343 (N_15343,N_838,N_7532);
and U15344 (N_15344,N_852,N_1103);
nand U15345 (N_15345,N_6277,N_1904);
xor U15346 (N_15346,N_4390,N_8716);
xor U15347 (N_15347,N_1633,N_1365);
nor U15348 (N_15348,N_1239,N_885);
and U15349 (N_15349,N_5335,N_4713);
or U15350 (N_15350,N_5702,N_7727);
xor U15351 (N_15351,N_3921,N_1028);
nor U15352 (N_15352,N_9577,N_3254);
nor U15353 (N_15353,N_9704,N_9115);
nand U15354 (N_15354,N_2926,N_9831);
xor U15355 (N_15355,N_5812,N_2623);
nor U15356 (N_15356,N_5453,N_5772);
xor U15357 (N_15357,N_1656,N_4122);
nor U15358 (N_15358,N_9816,N_3874);
or U15359 (N_15359,N_8824,N_830);
xnor U15360 (N_15360,N_2663,N_3574);
or U15361 (N_15361,N_4222,N_2042);
nor U15362 (N_15362,N_4807,N_2436);
or U15363 (N_15363,N_881,N_3589);
nand U15364 (N_15364,N_8587,N_9095);
or U15365 (N_15365,N_9171,N_732);
and U15366 (N_15366,N_9911,N_4412);
or U15367 (N_15367,N_1419,N_7181);
nand U15368 (N_15368,N_9252,N_3534);
and U15369 (N_15369,N_4558,N_3977);
and U15370 (N_15370,N_9401,N_13);
nor U15371 (N_15371,N_5169,N_6170);
nand U15372 (N_15372,N_8823,N_6887);
and U15373 (N_15373,N_6990,N_2151);
xnor U15374 (N_15374,N_6592,N_1822);
xor U15375 (N_15375,N_2737,N_2878);
nand U15376 (N_15376,N_1527,N_2519);
and U15377 (N_15377,N_5037,N_2724);
nand U15378 (N_15378,N_565,N_3849);
nand U15379 (N_15379,N_8699,N_6419);
xor U15380 (N_15380,N_859,N_3614);
or U15381 (N_15381,N_8892,N_8603);
nor U15382 (N_15382,N_2535,N_2150);
or U15383 (N_15383,N_7769,N_899);
and U15384 (N_15384,N_4330,N_1609);
xor U15385 (N_15385,N_423,N_9585);
nand U15386 (N_15386,N_25,N_3369);
xor U15387 (N_15387,N_9782,N_6108);
and U15388 (N_15388,N_1173,N_3993);
nand U15389 (N_15389,N_2345,N_7122);
and U15390 (N_15390,N_7967,N_8135);
xnor U15391 (N_15391,N_9947,N_7999);
or U15392 (N_15392,N_6884,N_5550);
or U15393 (N_15393,N_3717,N_4033);
nor U15394 (N_15394,N_2203,N_8608);
and U15395 (N_15395,N_7847,N_9084);
nor U15396 (N_15396,N_5979,N_9788);
and U15397 (N_15397,N_3253,N_1328);
nand U15398 (N_15398,N_9548,N_3573);
and U15399 (N_15399,N_4380,N_5483);
or U15400 (N_15400,N_9998,N_9585);
nand U15401 (N_15401,N_9349,N_2643);
nor U15402 (N_15402,N_1902,N_1973);
nor U15403 (N_15403,N_2291,N_1779);
nand U15404 (N_15404,N_1611,N_4138);
nor U15405 (N_15405,N_9847,N_3355);
and U15406 (N_15406,N_2670,N_6758);
and U15407 (N_15407,N_9037,N_3751);
nor U15408 (N_15408,N_5117,N_5174);
or U15409 (N_15409,N_1064,N_9012);
nor U15410 (N_15410,N_3399,N_720);
xor U15411 (N_15411,N_8475,N_4052);
xor U15412 (N_15412,N_4724,N_2161);
nand U15413 (N_15413,N_6202,N_8010);
or U15414 (N_15414,N_545,N_5259);
and U15415 (N_15415,N_4586,N_8054);
and U15416 (N_15416,N_6374,N_1068);
or U15417 (N_15417,N_6092,N_8907);
nor U15418 (N_15418,N_8255,N_2586);
xnor U15419 (N_15419,N_6679,N_4429);
nor U15420 (N_15420,N_6960,N_5583);
nand U15421 (N_15421,N_7695,N_3644);
nor U15422 (N_15422,N_856,N_2603);
or U15423 (N_15423,N_1724,N_8934);
and U15424 (N_15424,N_4543,N_2839);
and U15425 (N_15425,N_6697,N_2217);
nand U15426 (N_15426,N_9669,N_6844);
nor U15427 (N_15427,N_5752,N_8403);
and U15428 (N_15428,N_8195,N_5565);
nand U15429 (N_15429,N_7840,N_9798);
nor U15430 (N_15430,N_838,N_4139);
nor U15431 (N_15431,N_9667,N_5487);
xnor U15432 (N_15432,N_8291,N_2492);
xnor U15433 (N_15433,N_3945,N_3560);
xor U15434 (N_15434,N_5174,N_5229);
nand U15435 (N_15435,N_7140,N_8205);
and U15436 (N_15436,N_8950,N_8093);
nand U15437 (N_15437,N_8164,N_3022);
or U15438 (N_15438,N_9066,N_3229);
nand U15439 (N_15439,N_1459,N_4405);
xor U15440 (N_15440,N_417,N_3263);
xnor U15441 (N_15441,N_1811,N_4525);
nor U15442 (N_15442,N_1521,N_7546);
or U15443 (N_15443,N_459,N_5438);
nor U15444 (N_15444,N_9175,N_8776);
xor U15445 (N_15445,N_8351,N_6716);
xor U15446 (N_15446,N_4504,N_3609);
and U15447 (N_15447,N_663,N_1086);
nand U15448 (N_15448,N_1909,N_1170);
and U15449 (N_15449,N_4153,N_4697);
xor U15450 (N_15450,N_2629,N_1054);
or U15451 (N_15451,N_1990,N_4232);
nor U15452 (N_15452,N_7301,N_1672);
xnor U15453 (N_15453,N_434,N_7643);
nor U15454 (N_15454,N_4450,N_9352);
and U15455 (N_15455,N_6770,N_1186);
or U15456 (N_15456,N_8889,N_8872);
or U15457 (N_15457,N_1878,N_962);
xnor U15458 (N_15458,N_9136,N_3643);
or U15459 (N_15459,N_4868,N_9700);
xnor U15460 (N_15460,N_1466,N_1932);
and U15461 (N_15461,N_707,N_9588);
or U15462 (N_15462,N_5543,N_3080);
xor U15463 (N_15463,N_5426,N_6589);
and U15464 (N_15464,N_594,N_7491);
nand U15465 (N_15465,N_8644,N_6782);
xor U15466 (N_15466,N_6260,N_9777);
or U15467 (N_15467,N_3747,N_3252);
nand U15468 (N_15468,N_1737,N_6775);
nand U15469 (N_15469,N_4470,N_3491);
or U15470 (N_15470,N_4442,N_2890);
and U15471 (N_15471,N_6382,N_7984);
and U15472 (N_15472,N_5979,N_761);
or U15473 (N_15473,N_5044,N_8795);
xor U15474 (N_15474,N_3813,N_4922);
nand U15475 (N_15475,N_9274,N_7473);
nand U15476 (N_15476,N_8268,N_7550);
xnor U15477 (N_15477,N_4058,N_324);
and U15478 (N_15478,N_9410,N_4385);
and U15479 (N_15479,N_2027,N_2644);
nor U15480 (N_15480,N_101,N_2749);
or U15481 (N_15481,N_8210,N_5396);
and U15482 (N_15482,N_1804,N_6307);
nand U15483 (N_15483,N_1133,N_3575);
nor U15484 (N_15484,N_7536,N_233);
nor U15485 (N_15485,N_2134,N_6768);
nand U15486 (N_15486,N_4397,N_1448);
nor U15487 (N_15487,N_6304,N_4342);
and U15488 (N_15488,N_3847,N_8566);
xnor U15489 (N_15489,N_223,N_3927);
xor U15490 (N_15490,N_5043,N_3677);
or U15491 (N_15491,N_8481,N_7874);
nor U15492 (N_15492,N_8951,N_9905);
nor U15493 (N_15493,N_8724,N_3246);
or U15494 (N_15494,N_2055,N_3159);
nand U15495 (N_15495,N_9240,N_9302);
nor U15496 (N_15496,N_9071,N_2896);
nor U15497 (N_15497,N_8704,N_3786);
and U15498 (N_15498,N_9410,N_1355);
nand U15499 (N_15499,N_6270,N_4995);
and U15500 (N_15500,N_2658,N_8491);
nand U15501 (N_15501,N_7371,N_9989);
and U15502 (N_15502,N_6411,N_7708);
and U15503 (N_15503,N_7726,N_801);
and U15504 (N_15504,N_9295,N_9014);
nand U15505 (N_15505,N_1132,N_1412);
nand U15506 (N_15506,N_1068,N_164);
and U15507 (N_15507,N_1233,N_2434);
or U15508 (N_15508,N_8315,N_8853);
and U15509 (N_15509,N_4962,N_4661);
nand U15510 (N_15510,N_2695,N_2994);
nor U15511 (N_15511,N_2059,N_455);
and U15512 (N_15512,N_3137,N_2676);
nand U15513 (N_15513,N_2318,N_9127);
and U15514 (N_15514,N_1150,N_3164);
nor U15515 (N_15515,N_4626,N_4597);
xnor U15516 (N_15516,N_170,N_1767);
xnor U15517 (N_15517,N_5731,N_1999);
nand U15518 (N_15518,N_9948,N_9912);
nand U15519 (N_15519,N_6388,N_9737);
nor U15520 (N_15520,N_9469,N_167);
and U15521 (N_15521,N_4826,N_1376);
and U15522 (N_15522,N_2312,N_4893);
nor U15523 (N_15523,N_356,N_2320);
and U15524 (N_15524,N_8582,N_867);
nor U15525 (N_15525,N_5569,N_3133);
and U15526 (N_15526,N_534,N_9582);
nand U15527 (N_15527,N_7858,N_3960);
or U15528 (N_15528,N_5310,N_5275);
nor U15529 (N_15529,N_9715,N_5555);
nand U15530 (N_15530,N_5551,N_6469);
xor U15531 (N_15531,N_6247,N_755);
or U15532 (N_15532,N_1789,N_730);
and U15533 (N_15533,N_9277,N_5941);
nor U15534 (N_15534,N_2141,N_719);
nand U15535 (N_15535,N_7822,N_3540);
nand U15536 (N_15536,N_7911,N_3865);
and U15537 (N_15537,N_2710,N_8610);
xor U15538 (N_15538,N_9691,N_1925);
xnor U15539 (N_15539,N_74,N_9739);
xor U15540 (N_15540,N_8466,N_3168);
and U15541 (N_15541,N_1417,N_2110);
nand U15542 (N_15542,N_7546,N_3265);
or U15543 (N_15543,N_278,N_3984);
nand U15544 (N_15544,N_2181,N_9156);
xnor U15545 (N_15545,N_8990,N_9496);
nand U15546 (N_15546,N_1332,N_8040);
or U15547 (N_15547,N_8303,N_8782);
nor U15548 (N_15548,N_5191,N_6561);
or U15549 (N_15549,N_6154,N_5062);
xnor U15550 (N_15550,N_3102,N_7479);
xor U15551 (N_15551,N_5671,N_6694);
nor U15552 (N_15552,N_7835,N_6306);
and U15553 (N_15553,N_1202,N_1789);
nor U15554 (N_15554,N_4199,N_3728);
nand U15555 (N_15555,N_8015,N_9964);
or U15556 (N_15556,N_1914,N_4621);
nor U15557 (N_15557,N_5065,N_610);
nand U15558 (N_15558,N_1156,N_1249);
xor U15559 (N_15559,N_139,N_7588);
xnor U15560 (N_15560,N_8337,N_8208);
and U15561 (N_15561,N_539,N_8686);
and U15562 (N_15562,N_7395,N_3022);
nor U15563 (N_15563,N_4409,N_2871);
and U15564 (N_15564,N_210,N_9858);
and U15565 (N_15565,N_860,N_6154);
nand U15566 (N_15566,N_580,N_4712);
xor U15567 (N_15567,N_3522,N_3769);
nand U15568 (N_15568,N_7956,N_1861);
or U15569 (N_15569,N_5700,N_8929);
nand U15570 (N_15570,N_8413,N_6305);
nand U15571 (N_15571,N_2733,N_321);
nor U15572 (N_15572,N_7015,N_6119);
nand U15573 (N_15573,N_5722,N_4689);
and U15574 (N_15574,N_3995,N_6628);
or U15575 (N_15575,N_6901,N_1348);
xnor U15576 (N_15576,N_1362,N_3574);
or U15577 (N_15577,N_4580,N_5670);
xnor U15578 (N_15578,N_5071,N_9347);
nor U15579 (N_15579,N_2825,N_7321);
or U15580 (N_15580,N_2387,N_6067);
and U15581 (N_15581,N_3043,N_2240);
xnor U15582 (N_15582,N_2826,N_857);
xnor U15583 (N_15583,N_2274,N_7252);
or U15584 (N_15584,N_8864,N_6289);
nor U15585 (N_15585,N_5386,N_4557);
and U15586 (N_15586,N_6018,N_654);
nand U15587 (N_15587,N_3249,N_3576);
or U15588 (N_15588,N_8953,N_5735);
nor U15589 (N_15589,N_6542,N_8981);
or U15590 (N_15590,N_4349,N_7361);
nor U15591 (N_15591,N_6109,N_8687);
or U15592 (N_15592,N_1831,N_7754);
nor U15593 (N_15593,N_2964,N_4599);
xnor U15594 (N_15594,N_672,N_4951);
nor U15595 (N_15595,N_4525,N_7300);
nand U15596 (N_15596,N_4157,N_4971);
and U15597 (N_15597,N_2688,N_2278);
or U15598 (N_15598,N_3477,N_9345);
xor U15599 (N_15599,N_737,N_9395);
and U15600 (N_15600,N_1191,N_1707);
nand U15601 (N_15601,N_6740,N_6602);
nand U15602 (N_15602,N_6265,N_9535);
nand U15603 (N_15603,N_5573,N_3397);
or U15604 (N_15604,N_8054,N_7242);
and U15605 (N_15605,N_8095,N_8258);
xnor U15606 (N_15606,N_4111,N_3035);
or U15607 (N_15607,N_6100,N_168);
nor U15608 (N_15608,N_861,N_5081);
and U15609 (N_15609,N_2907,N_8383);
nand U15610 (N_15610,N_7186,N_673);
or U15611 (N_15611,N_394,N_1608);
xor U15612 (N_15612,N_203,N_572);
and U15613 (N_15613,N_7569,N_7077);
and U15614 (N_15614,N_8976,N_7105);
xnor U15615 (N_15615,N_3366,N_5924);
xor U15616 (N_15616,N_3487,N_1272);
or U15617 (N_15617,N_6360,N_130);
nor U15618 (N_15618,N_5510,N_7884);
and U15619 (N_15619,N_7323,N_5222);
nor U15620 (N_15620,N_9755,N_8864);
nand U15621 (N_15621,N_5622,N_3432);
and U15622 (N_15622,N_7044,N_8526);
xnor U15623 (N_15623,N_6738,N_9850);
and U15624 (N_15624,N_2562,N_260);
nand U15625 (N_15625,N_2317,N_9482);
nor U15626 (N_15626,N_8015,N_666);
and U15627 (N_15627,N_8024,N_4705);
and U15628 (N_15628,N_8270,N_6774);
or U15629 (N_15629,N_9512,N_9913);
and U15630 (N_15630,N_2534,N_1091);
nor U15631 (N_15631,N_4442,N_5649);
nand U15632 (N_15632,N_5240,N_2722);
nand U15633 (N_15633,N_6072,N_7532);
nand U15634 (N_15634,N_8521,N_8793);
nor U15635 (N_15635,N_7273,N_6939);
nor U15636 (N_15636,N_7647,N_5909);
and U15637 (N_15637,N_61,N_9855);
nand U15638 (N_15638,N_6301,N_1557);
nand U15639 (N_15639,N_1866,N_9747);
xnor U15640 (N_15640,N_9604,N_1501);
and U15641 (N_15641,N_8165,N_3098);
and U15642 (N_15642,N_8598,N_5260);
nand U15643 (N_15643,N_6149,N_1885);
and U15644 (N_15644,N_6643,N_3249);
or U15645 (N_15645,N_7733,N_7747);
or U15646 (N_15646,N_2773,N_721);
and U15647 (N_15647,N_956,N_5712);
nand U15648 (N_15648,N_8762,N_6024);
xnor U15649 (N_15649,N_1608,N_2416);
nor U15650 (N_15650,N_2187,N_7539);
or U15651 (N_15651,N_2825,N_3083);
nand U15652 (N_15652,N_7818,N_1767);
nor U15653 (N_15653,N_9543,N_7881);
nor U15654 (N_15654,N_3296,N_6347);
nor U15655 (N_15655,N_6480,N_4503);
xor U15656 (N_15656,N_1977,N_2552);
nand U15657 (N_15657,N_3938,N_860);
nand U15658 (N_15658,N_8610,N_7267);
xor U15659 (N_15659,N_6964,N_9736);
or U15660 (N_15660,N_304,N_6861);
and U15661 (N_15661,N_8611,N_458);
xor U15662 (N_15662,N_5159,N_4867);
or U15663 (N_15663,N_5740,N_3151);
xnor U15664 (N_15664,N_269,N_7862);
or U15665 (N_15665,N_6479,N_1599);
xnor U15666 (N_15666,N_4086,N_1269);
and U15667 (N_15667,N_9725,N_5429);
or U15668 (N_15668,N_1393,N_6860);
xnor U15669 (N_15669,N_1542,N_4418);
or U15670 (N_15670,N_5803,N_937);
xnor U15671 (N_15671,N_417,N_8666);
nand U15672 (N_15672,N_5994,N_6504);
nor U15673 (N_15673,N_1491,N_7141);
or U15674 (N_15674,N_9011,N_2726);
and U15675 (N_15675,N_9961,N_641);
nand U15676 (N_15676,N_4547,N_381);
or U15677 (N_15677,N_991,N_9932);
nand U15678 (N_15678,N_6461,N_8669);
and U15679 (N_15679,N_6786,N_5449);
nand U15680 (N_15680,N_8615,N_521);
and U15681 (N_15681,N_9707,N_8971);
xnor U15682 (N_15682,N_5464,N_3555);
nor U15683 (N_15683,N_3402,N_1259);
nand U15684 (N_15684,N_4772,N_4135);
nand U15685 (N_15685,N_2523,N_4934);
or U15686 (N_15686,N_791,N_3932);
nand U15687 (N_15687,N_3303,N_156);
and U15688 (N_15688,N_2337,N_221);
and U15689 (N_15689,N_2023,N_2313);
or U15690 (N_15690,N_4267,N_986);
nor U15691 (N_15691,N_2965,N_2064);
nand U15692 (N_15692,N_4383,N_263);
xnor U15693 (N_15693,N_4921,N_2351);
nor U15694 (N_15694,N_3171,N_9398);
or U15695 (N_15695,N_5545,N_6167);
or U15696 (N_15696,N_3770,N_9684);
xnor U15697 (N_15697,N_8317,N_2092);
xnor U15698 (N_15698,N_5138,N_3503);
nand U15699 (N_15699,N_2317,N_2666);
xnor U15700 (N_15700,N_8808,N_4687);
or U15701 (N_15701,N_4179,N_2044);
and U15702 (N_15702,N_2537,N_2914);
nand U15703 (N_15703,N_8800,N_8398);
and U15704 (N_15704,N_5593,N_5130);
or U15705 (N_15705,N_4935,N_1243);
nor U15706 (N_15706,N_1584,N_3993);
xor U15707 (N_15707,N_1049,N_4342);
nor U15708 (N_15708,N_3272,N_4298);
or U15709 (N_15709,N_9179,N_913);
or U15710 (N_15710,N_4864,N_5467);
and U15711 (N_15711,N_6195,N_1910);
nand U15712 (N_15712,N_5446,N_990);
and U15713 (N_15713,N_1368,N_381);
or U15714 (N_15714,N_5783,N_8470);
nand U15715 (N_15715,N_4420,N_8633);
nor U15716 (N_15716,N_6309,N_1994);
xnor U15717 (N_15717,N_7945,N_1225);
nor U15718 (N_15718,N_2893,N_188);
or U15719 (N_15719,N_9717,N_2208);
or U15720 (N_15720,N_3825,N_6104);
xnor U15721 (N_15721,N_7998,N_1165);
xor U15722 (N_15722,N_6362,N_5725);
nand U15723 (N_15723,N_4236,N_2942);
nand U15724 (N_15724,N_4871,N_4339);
and U15725 (N_15725,N_9516,N_827);
xor U15726 (N_15726,N_2786,N_3662);
xor U15727 (N_15727,N_9481,N_4771);
nor U15728 (N_15728,N_1649,N_5731);
nor U15729 (N_15729,N_3949,N_1711);
xor U15730 (N_15730,N_4825,N_4528);
nor U15731 (N_15731,N_2961,N_8998);
or U15732 (N_15732,N_9628,N_1505);
or U15733 (N_15733,N_9783,N_8518);
nand U15734 (N_15734,N_1756,N_8345);
nand U15735 (N_15735,N_8166,N_1589);
nand U15736 (N_15736,N_5301,N_6950);
nor U15737 (N_15737,N_2676,N_654);
xnor U15738 (N_15738,N_6399,N_850);
and U15739 (N_15739,N_3873,N_8450);
nor U15740 (N_15740,N_55,N_5087);
and U15741 (N_15741,N_7399,N_7181);
and U15742 (N_15742,N_2453,N_86);
nor U15743 (N_15743,N_9438,N_2139);
xnor U15744 (N_15744,N_3048,N_5024);
nand U15745 (N_15745,N_1862,N_9512);
xor U15746 (N_15746,N_2240,N_1674);
nand U15747 (N_15747,N_4753,N_7144);
nor U15748 (N_15748,N_479,N_7055);
and U15749 (N_15749,N_2076,N_8091);
and U15750 (N_15750,N_2614,N_8450);
or U15751 (N_15751,N_9153,N_4182);
or U15752 (N_15752,N_8521,N_2250);
or U15753 (N_15753,N_2944,N_7741);
nand U15754 (N_15754,N_3913,N_893);
nand U15755 (N_15755,N_2695,N_5784);
and U15756 (N_15756,N_6787,N_2035);
or U15757 (N_15757,N_7930,N_701);
xnor U15758 (N_15758,N_9430,N_4931);
nand U15759 (N_15759,N_5057,N_3724);
nand U15760 (N_15760,N_9346,N_2424);
and U15761 (N_15761,N_6566,N_5930);
nand U15762 (N_15762,N_7164,N_6480);
nand U15763 (N_15763,N_5652,N_1796);
and U15764 (N_15764,N_258,N_133);
nand U15765 (N_15765,N_7575,N_9381);
nor U15766 (N_15766,N_8675,N_3923);
or U15767 (N_15767,N_8532,N_5493);
xor U15768 (N_15768,N_3372,N_9538);
or U15769 (N_15769,N_820,N_6559);
and U15770 (N_15770,N_6293,N_8446);
and U15771 (N_15771,N_6637,N_2254);
or U15772 (N_15772,N_4522,N_614);
nor U15773 (N_15773,N_7500,N_1868);
xnor U15774 (N_15774,N_9156,N_8971);
nor U15775 (N_15775,N_2300,N_891);
nand U15776 (N_15776,N_9092,N_9656);
nand U15777 (N_15777,N_4627,N_6007);
and U15778 (N_15778,N_5109,N_2858);
or U15779 (N_15779,N_7178,N_3322);
xnor U15780 (N_15780,N_2609,N_8687);
or U15781 (N_15781,N_4287,N_4073);
nand U15782 (N_15782,N_9888,N_7160);
and U15783 (N_15783,N_712,N_3964);
nand U15784 (N_15784,N_5588,N_4438);
and U15785 (N_15785,N_7198,N_5483);
or U15786 (N_15786,N_4064,N_5104);
and U15787 (N_15787,N_7961,N_1843);
and U15788 (N_15788,N_4143,N_8879);
or U15789 (N_15789,N_4400,N_5586);
xnor U15790 (N_15790,N_3253,N_8636);
xor U15791 (N_15791,N_8973,N_747);
or U15792 (N_15792,N_4240,N_7864);
xnor U15793 (N_15793,N_2752,N_7411);
nand U15794 (N_15794,N_1350,N_5455);
and U15795 (N_15795,N_9605,N_459);
and U15796 (N_15796,N_242,N_5244);
xor U15797 (N_15797,N_2731,N_3454);
or U15798 (N_15798,N_6046,N_9008);
xor U15799 (N_15799,N_2661,N_80);
nand U15800 (N_15800,N_3748,N_8386);
nor U15801 (N_15801,N_8616,N_9016);
xnor U15802 (N_15802,N_1198,N_6204);
xor U15803 (N_15803,N_1848,N_7379);
or U15804 (N_15804,N_7302,N_9357);
nand U15805 (N_15805,N_8042,N_7682);
xor U15806 (N_15806,N_9676,N_1396);
nand U15807 (N_15807,N_4064,N_8656);
xor U15808 (N_15808,N_2823,N_3224);
or U15809 (N_15809,N_4581,N_3256);
and U15810 (N_15810,N_2724,N_3163);
and U15811 (N_15811,N_9205,N_3593);
or U15812 (N_15812,N_4600,N_9849);
or U15813 (N_15813,N_9422,N_8341);
and U15814 (N_15814,N_1225,N_7498);
or U15815 (N_15815,N_1660,N_6445);
nor U15816 (N_15816,N_2335,N_9344);
or U15817 (N_15817,N_1782,N_9232);
nor U15818 (N_15818,N_7970,N_6073);
and U15819 (N_15819,N_2605,N_2676);
or U15820 (N_15820,N_9935,N_8846);
xnor U15821 (N_15821,N_6580,N_2474);
and U15822 (N_15822,N_2917,N_5887);
nor U15823 (N_15823,N_7145,N_5170);
nand U15824 (N_15824,N_2498,N_882);
and U15825 (N_15825,N_2233,N_8564);
or U15826 (N_15826,N_4238,N_3406);
xor U15827 (N_15827,N_4270,N_2466);
and U15828 (N_15828,N_7222,N_3295);
xor U15829 (N_15829,N_1446,N_6866);
nor U15830 (N_15830,N_5469,N_9040);
and U15831 (N_15831,N_8368,N_4016);
nand U15832 (N_15832,N_9224,N_1869);
nand U15833 (N_15833,N_1906,N_9099);
or U15834 (N_15834,N_5270,N_3920);
xor U15835 (N_15835,N_6532,N_7108);
nor U15836 (N_15836,N_3111,N_6624);
nand U15837 (N_15837,N_4669,N_635);
nand U15838 (N_15838,N_3062,N_2557);
or U15839 (N_15839,N_2864,N_348);
xnor U15840 (N_15840,N_9672,N_8771);
and U15841 (N_15841,N_3777,N_7458);
nand U15842 (N_15842,N_2366,N_5935);
and U15843 (N_15843,N_1937,N_31);
nor U15844 (N_15844,N_555,N_1497);
nor U15845 (N_15845,N_3137,N_2123);
nand U15846 (N_15846,N_8229,N_4935);
xor U15847 (N_15847,N_2696,N_4315);
and U15848 (N_15848,N_3187,N_2095);
and U15849 (N_15849,N_9788,N_8335);
and U15850 (N_15850,N_7167,N_5719);
nand U15851 (N_15851,N_8023,N_6007);
nand U15852 (N_15852,N_7544,N_1154);
nor U15853 (N_15853,N_9418,N_5458);
or U15854 (N_15854,N_8691,N_7532);
and U15855 (N_15855,N_5670,N_2186);
and U15856 (N_15856,N_5826,N_8646);
nor U15857 (N_15857,N_5090,N_4528);
and U15858 (N_15858,N_2210,N_1429);
xor U15859 (N_15859,N_3314,N_7173);
nand U15860 (N_15860,N_7618,N_4031);
and U15861 (N_15861,N_3174,N_2553);
xnor U15862 (N_15862,N_5134,N_1135);
nor U15863 (N_15863,N_9203,N_7525);
nand U15864 (N_15864,N_4074,N_9517);
nor U15865 (N_15865,N_5582,N_9350);
nor U15866 (N_15866,N_3743,N_7924);
or U15867 (N_15867,N_9151,N_1290);
nand U15868 (N_15868,N_1241,N_9445);
nor U15869 (N_15869,N_4680,N_1803);
or U15870 (N_15870,N_6438,N_8869);
nor U15871 (N_15871,N_7752,N_9246);
nand U15872 (N_15872,N_5480,N_4738);
nand U15873 (N_15873,N_6835,N_4090);
xor U15874 (N_15874,N_81,N_910);
or U15875 (N_15875,N_557,N_1412);
nand U15876 (N_15876,N_4957,N_2275);
xor U15877 (N_15877,N_9546,N_1110);
nor U15878 (N_15878,N_2433,N_6599);
nand U15879 (N_15879,N_7291,N_9430);
nor U15880 (N_15880,N_1940,N_1836);
xor U15881 (N_15881,N_9519,N_5838);
or U15882 (N_15882,N_9208,N_2714);
and U15883 (N_15883,N_1155,N_7755);
or U15884 (N_15884,N_5216,N_1008);
xor U15885 (N_15885,N_6676,N_5672);
or U15886 (N_15886,N_1607,N_1922);
xnor U15887 (N_15887,N_9037,N_5127);
nand U15888 (N_15888,N_9202,N_3276);
and U15889 (N_15889,N_9313,N_6085);
xor U15890 (N_15890,N_2026,N_1734);
and U15891 (N_15891,N_7126,N_3786);
nor U15892 (N_15892,N_7932,N_9096);
nor U15893 (N_15893,N_576,N_6373);
nor U15894 (N_15894,N_8590,N_9836);
or U15895 (N_15895,N_5990,N_7314);
and U15896 (N_15896,N_7842,N_515);
or U15897 (N_15897,N_8607,N_5554);
and U15898 (N_15898,N_1690,N_5622);
nand U15899 (N_15899,N_1526,N_7455);
or U15900 (N_15900,N_5251,N_854);
and U15901 (N_15901,N_7135,N_5578);
and U15902 (N_15902,N_3777,N_2317);
and U15903 (N_15903,N_32,N_5566);
nor U15904 (N_15904,N_2551,N_1355);
and U15905 (N_15905,N_8552,N_8968);
and U15906 (N_15906,N_9652,N_8533);
nand U15907 (N_15907,N_1075,N_2525);
nand U15908 (N_15908,N_6323,N_1049);
and U15909 (N_15909,N_1024,N_8371);
nor U15910 (N_15910,N_8520,N_6549);
and U15911 (N_15911,N_129,N_1513);
and U15912 (N_15912,N_7556,N_9655);
nor U15913 (N_15913,N_9543,N_6212);
nand U15914 (N_15914,N_6141,N_5010);
and U15915 (N_15915,N_4552,N_1083);
xnor U15916 (N_15916,N_5963,N_894);
nor U15917 (N_15917,N_7171,N_3977);
and U15918 (N_15918,N_5577,N_3900);
or U15919 (N_15919,N_5571,N_9880);
xnor U15920 (N_15920,N_4237,N_4284);
and U15921 (N_15921,N_5147,N_1969);
and U15922 (N_15922,N_9198,N_4400);
and U15923 (N_15923,N_512,N_736);
nand U15924 (N_15924,N_1893,N_3038);
nor U15925 (N_15925,N_6971,N_3396);
nand U15926 (N_15926,N_4753,N_9937);
nand U15927 (N_15927,N_8790,N_1356);
or U15928 (N_15928,N_9279,N_7111);
nor U15929 (N_15929,N_9059,N_6026);
nor U15930 (N_15930,N_4605,N_5314);
and U15931 (N_15931,N_6324,N_5358);
or U15932 (N_15932,N_2543,N_2955);
or U15933 (N_15933,N_791,N_3536);
or U15934 (N_15934,N_1268,N_4732);
or U15935 (N_15935,N_3870,N_7980);
or U15936 (N_15936,N_6976,N_2727);
or U15937 (N_15937,N_7106,N_9714);
and U15938 (N_15938,N_8643,N_4045);
xnor U15939 (N_15939,N_5964,N_7717);
xnor U15940 (N_15940,N_1850,N_5681);
xor U15941 (N_15941,N_8592,N_2542);
or U15942 (N_15942,N_5840,N_9298);
xnor U15943 (N_15943,N_7883,N_1991);
nand U15944 (N_15944,N_331,N_3387);
and U15945 (N_15945,N_3802,N_8191);
xor U15946 (N_15946,N_1506,N_6317);
xnor U15947 (N_15947,N_1213,N_614);
xnor U15948 (N_15948,N_5243,N_2910);
nand U15949 (N_15949,N_4198,N_8311);
or U15950 (N_15950,N_7552,N_9757);
or U15951 (N_15951,N_5347,N_3864);
nor U15952 (N_15952,N_6864,N_8400);
and U15953 (N_15953,N_5749,N_7856);
nor U15954 (N_15954,N_3897,N_4717);
nand U15955 (N_15955,N_8716,N_484);
and U15956 (N_15956,N_1496,N_7470);
xnor U15957 (N_15957,N_8030,N_9469);
nand U15958 (N_15958,N_8449,N_7786);
nor U15959 (N_15959,N_4849,N_2528);
nor U15960 (N_15960,N_1334,N_6729);
xor U15961 (N_15961,N_1596,N_2821);
nor U15962 (N_15962,N_2196,N_8562);
nand U15963 (N_15963,N_6984,N_8736);
nor U15964 (N_15964,N_1666,N_9838);
xnor U15965 (N_15965,N_8687,N_2526);
or U15966 (N_15966,N_5980,N_1639);
nand U15967 (N_15967,N_1665,N_4734);
xor U15968 (N_15968,N_6593,N_282);
nand U15969 (N_15969,N_2271,N_2755);
nand U15970 (N_15970,N_5126,N_7509);
or U15971 (N_15971,N_1560,N_661);
and U15972 (N_15972,N_496,N_4225);
and U15973 (N_15973,N_34,N_3694);
and U15974 (N_15974,N_1581,N_5889);
nor U15975 (N_15975,N_3551,N_5838);
and U15976 (N_15976,N_1465,N_6035);
nand U15977 (N_15977,N_3900,N_6339);
xnor U15978 (N_15978,N_4603,N_7234);
nor U15979 (N_15979,N_1518,N_3988);
nand U15980 (N_15980,N_4277,N_5417);
xor U15981 (N_15981,N_7137,N_8323);
nand U15982 (N_15982,N_1132,N_6394);
and U15983 (N_15983,N_6848,N_1066);
and U15984 (N_15984,N_4625,N_2395);
and U15985 (N_15985,N_4689,N_9090);
nor U15986 (N_15986,N_7232,N_6745);
and U15987 (N_15987,N_2424,N_2302);
or U15988 (N_15988,N_8855,N_2887);
xnor U15989 (N_15989,N_8604,N_8715);
xor U15990 (N_15990,N_2393,N_7251);
nand U15991 (N_15991,N_9103,N_1952);
xnor U15992 (N_15992,N_1135,N_2367);
or U15993 (N_15993,N_1032,N_7545);
xor U15994 (N_15994,N_3945,N_1073);
and U15995 (N_15995,N_6053,N_9529);
nand U15996 (N_15996,N_3671,N_7946);
or U15997 (N_15997,N_7614,N_4940);
xnor U15998 (N_15998,N_4104,N_4471);
nand U15999 (N_15999,N_425,N_1940);
and U16000 (N_16000,N_6587,N_7939);
nor U16001 (N_16001,N_337,N_8856);
and U16002 (N_16002,N_2879,N_7994);
xor U16003 (N_16003,N_2159,N_8398);
nand U16004 (N_16004,N_7877,N_1706);
xnor U16005 (N_16005,N_9333,N_608);
nor U16006 (N_16006,N_5272,N_1805);
nor U16007 (N_16007,N_4734,N_6945);
and U16008 (N_16008,N_1918,N_8471);
nor U16009 (N_16009,N_8720,N_8928);
nor U16010 (N_16010,N_963,N_5617);
nand U16011 (N_16011,N_3397,N_8030);
nand U16012 (N_16012,N_6044,N_4111);
or U16013 (N_16013,N_5581,N_8041);
and U16014 (N_16014,N_9870,N_1330);
or U16015 (N_16015,N_9707,N_5987);
and U16016 (N_16016,N_3908,N_158);
or U16017 (N_16017,N_5297,N_509);
nand U16018 (N_16018,N_8312,N_1297);
or U16019 (N_16019,N_283,N_1957);
xnor U16020 (N_16020,N_4176,N_5226);
and U16021 (N_16021,N_5270,N_4941);
xnor U16022 (N_16022,N_2436,N_4071);
xnor U16023 (N_16023,N_1619,N_2176);
nor U16024 (N_16024,N_8873,N_5659);
nand U16025 (N_16025,N_5513,N_4326);
or U16026 (N_16026,N_5497,N_761);
nand U16027 (N_16027,N_1258,N_5751);
nand U16028 (N_16028,N_4631,N_9301);
and U16029 (N_16029,N_2104,N_8769);
xnor U16030 (N_16030,N_5254,N_6679);
and U16031 (N_16031,N_4498,N_8155);
xnor U16032 (N_16032,N_9357,N_6509);
and U16033 (N_16033,N_5814,N_436);
nor U16034 (N_16034,N_2167,N_372);
xor U16035 (N_16035,N_4979,N_7844);
xnor U16036 (N_16036,N_7137,N_1923);
nand U16037 (N_16037,N_4845,N_6444);
and U16038 (N_16038,N_7718,N_1213);
xnor U16039 (N_16039,N_4459,N_9535);
nor U16040 (N_16040,N_2142,N_8010);
and U16041 (N_16041,N_3574,N_7158);
nor U16042 (N_16042,N_9958,N_8218);
nand U16043 (N_16043,N_8945,N_6483);
nand U16044 (N_16044,N_4115,N_4257);
or U16045 (N_16045,N_8818,N_8794);
nor U16046 (N_16046,N_5484,N_5590);
and U16047 (N_16047,N_2087,N_5661);
xnor U16048 (N_16048,N_5919,N_5140);
and U16049 (N_16049,N_4166,N_674);
and U16050 (N_16050,N_5004,N_9756);
nor U16051 (N_16051,N_8991,N_1965);
xnor U16052 (N_16052,N_1883,N_3812);
nor U16053 (N_16053,N_9292,N_1424);
nand U16054 (N_16054,N_7321,N_5648);
nand U16055 (N_16055,N_8748,N_8805);
or U16056 (N_16056,N_8779,N_1481);
xnor U16057 (N_16057,N_9964,N_1211);
or U16058 (N_16058,N_8485,N_1751);
and U16059 (N_16059,N_6490,N_4801);
nor U16060 (N_16060,N_6426,N_6943);
nand U16061 (N_16061,N_9482,N_3427);
and U16062 (N_16062,N_5164,N_7807);
xor U16063 (N_16063,N_5247,N_6045);
and U16064 (N_16064,N_250,N_7517);
and U16065 (N_16065,N_1062,N_5543);
nand U16066 (N_16066,N_5650,N_8768);
or U16067 (N_16067,N_9568,N_1381);
nand U16068 (N_16068,N_6790,N_8157);
xor U16069 (N_16069,N_5805,N_7893);
nor U16070 (N_16070,N_1408,N_5161);
and U16071 (N_16071,N_6436,N_2505);
nand U16072 (N_16072,N_84,N_4296);
nand U16073 (N_16073,N_7188,N_5725);
nor U16074 (N_16074,N_9866,N_4767);
nand U16075 (N_16075,N_1694,N_6486);
xnor U16076 (N_16076,N_2691,N_8854);
nor U16077 (N_16077,N_7642,N_8909);
and U16078 (N_16078,N_8754,N_4257);
and U16079 (N_16079,N_2430,N_5777);
or U16080 (N_16080,N_7880,N_5957);
and U16081 (N_16081,N_8235,N_4335);
and U16082 (N_16082,N_2417,N_8907);
and U16083 (N_16083,N_8013,N_3464);
nor U16084 (N_16084,N_1136,N_8741);
or U16085 (N_16085,N_6955,N_9224);
nand U16086 (N_16086,N_5699,N_4558);
nand U16087 (N_16087,N_2479,N_9633);
and U16088 (N_16088,N_1473,N_2568);
nor U16089 (N_16089,N_3038,N_8685);
or U16090 (N_16090,N_2848,N_4848);
xor U16091 (N_16091,N_4862,N_1037);
nor U16092 (N_16092,N_3833,N_7363);
or U16093 (N_16093,N_2972,N_7135);
or U16094 (N_16094,N_3502,N_1970);
xnor U16095 (N_16095,N_9492,N_2603);
nor U16096 (N_16096,N_841,N_6082);
nand U16097 (N_16097,N_3879,N_6840);
nand U16098 (N_16098,N_2578,N_1665);
and U16099 (N_16099,N_9688,N_885);
or U16100 (N_16100,N_9504,N_2218);
nor U16101 (N_16101,N_8538,N_5867);
nor U16102 (N_16102,N_5102,N_2783);
nor U16103 (N_16103,N_7744,N_3093);
nand U16104 (N_16104,N_8438,N_6080);
or U16105 (N_16105,N_4338,N_7786);
nand U16106 (N_16106,N_2313,N_34);
or U16107 (N_16107,N_3529,N_7621);
nor U16108 (N_16108,N_4177,N_8877);
nor U16109 (N_16109,N_4092,N_9150);
xor U16110 (N_16110,N_5823,N_7306);
or U16111 (N_16111,N_8520,N_3755);
nand U16112 (N_16112,N_8914,N_1695);
xnor U16113 (N_16113,N_6768,N_2261);
and U16114 (N_16114,N_8076,N_4419);
and U16115 (N_16115,N_168,N_4307);
and U16116 (N_16116,N_6130,N_2464);
and U16117 (N_16117,N_6487,N_1127);
nor U16118 (N_16118,N_6643,N_839);
nand U16119 (N_16119,N_3887,N_7591);
nor U16120 (N_16120,N_3607,N_3821);
and U16121 (N_16121,N_4262,N_1563);
and U16122 (N_16122,N_903,N_2666);
nor U16123 (N_16123,N_8920,N_8112);
or U16124 (N_16124,N_3021,N_7460);
xnor U16125 (N_16125,N_5173,N_9184);
or U16126 (N_16126,N_5445,N_259);
and U16127 (N_16127,N_8957,N_8757);
and U16128 (N_16128,N_4778,N_4754);
nor U16129 (N_16129,N_2575,N_4104);
and U16130 (N_16130,N_9542,N_5412);
nor U16131 (N_16131,N_7514,N_1482);
nand U16132 (N_16132,N_1939,N_192);
or U16133 (N_16133,N_7258,N_987);
xnor U16134 (N_16134,N_5951,N_9273);
nor U16135 (N_16135,N_5769,N_7558);
and U16136 (N_16136,N_6559,N_3488);
xnor U16137 (N_16137,N_4951,N_926);
and U16138 (N_16138,N_1223,N_999);
nand U16139 (N_16139,N_5466,N_465);
xor U16140 (N_16140,N_1856,N_8785);
and U16141 (N_16141,N_7545,N_9597);
nor U16142 (N_16142,N_1002,N_3607);
and U16143 (N_16143,N_680,N_5406);
nand U16144 (N_16144,N_842,N_7216);
nand U16145 (N_16145,N_9962,N_2941);
or U16146 (N_16146,N_8643,N_9177);
and U16147 (N_16147,N_7707,N_5834);
or U16148 (N_16148,N_566,N_1074);
nor U16149 (N_16149,N_4510,N_2576);
nor U16150 (N_16150,N_2166,N_6898);
xor U16151 (N_16151,N_125,N_6630);
and U16152 (N_16152,N_2329,N_7408);
nor U16153 (N_16153,N_7071,N_3975);
nand U16154 (N_16154,N_1052,N_102);
nor U16155 (N_16155,N_6087,N_5494);
nand U16156 (N_16156,N_459,N_6960);
nor U16157 (N_16157,N_9729,N_9099);
or U16158 (N_16158,N_9910,N_424);
nor U16159 (N_16159,N_4340,N_1907);
and U16160 (N_16160,N_9938,N_3206);
and U16161 (N_16161,N_4613,N_1572);
xor U16162 (N_16162,N_1046,N_823);
nor U16163 (N_16163,N_9783,N_5769);
nand U16164 (N_16164,N_4443,N_6108);
xor U16165 (N_16165,N_4560,N_4402);
xor U16166 (N_16166,N_6478,N_2272);
nand U16167 (N_16167,N_2478,N_5939);
or U16168 (N_16168,N_3192,N_6038);
nand U16169 (N_16169,N_8769,N_9439);
xnor U16170 (N_16170,N_9326,N_5654);
nand U16171 (N_16171,N_1972,N_7553);
nor U16172 (N_16172,N_1483,N_5773);
nor U16173 (N_16173,N_4904,N_6323);
nor U16174 (N_16174,N_9017,N_5222);
nand U16175 (N_16175,N_4268,N_383);
xor U16176 (N_16176,N_8499,N_3736);
nand U16177 (N_16177,N_5133,N_3583);
nand U16178 (N_16178,N_2872,N_5134);
nand U16179 (N_16179,N_7268,N_812);
or U16180 (N_16180,N_6559,N_4054);
or U16181 (N_16181,N_4694,N_553);
nand U16182 (N_16182,N_5211,N_4609);
xnor U16183 (N_16183,N_7074,N_3631);
nor U16184 (N_16184,N_7960,N_1144);
nand U16185 (N_16185,N_130,N_4581);
or U16186 (N_16186,N_3094,N_4718);
nor U16187 (N_16187,N_1785,N_7281);
nand U16188 (N_16188,N_6010,N_1097);
nand U16189 (N_16189,N_6491,N_1878);
or U16190 (N_16190,N_1012,N_4607);
or U16191 (N_16191,N_6073,N_7868);
and U16192 (N_16192,N_859,N_2399);
or U16193 (N_16193,N_259,N_9826);
and U16194 (N_16194,N_881,N_5888);
nor U16195 (N_16195,N_6585,N_8831);
or U16196 (N_16196,N_9208,N_6);
and U16197 (N_16197,N_1581,N_2876);
and U16198 (N_16198,N_6767,N_9833);
xnor U16199 (N_16199,N_5730,N_5692);
or U16200 (N_16200,N_6721,N_2527);
nor U16201 (N_16201,N_1203,N_8999);
nand U16202 (N_16202,N_5013,N_7515);
or U16203 (N_16203,N_6632,N_7960);
nand U16204 (N_16204,N_5371,N_3394);
nor U16205 (N_16205,N_3760,N_197);
nor U16206 (N_16206,N_6309,N_5025);
nor U16207 (N_16207,N_8406,N_1522);
and U16208 (N_16208,N_2019,N_4919);
or U16209 (N_16209,N_3790,N_926);
nor U16210 (N_16210,N_201,N_2707);
and U16211 (N_16211,N_1280,N_3499);
nand U16212 (N_16212,N_3530,N_3242);
and U16213 (N_16213,N_1969,N_6496);
or U16214 (N_16214,N_8747,N_1295);
or U16215 (N_16215,N_702,N_2871);
nor U16216 (N_16216,N_8453,N_6161);
nand U16217 (N_16217,N_8401,N_3766);
and U16218 (N_16218,N_8745,N_7421);
xor U16219 (N_16219,N_2650,N_6351);
xnor U16220 (N_16220,N_6106,N_1501);
nand U16221 (N_16221,N_6012,N_7988);
nand U16222 (N_16222,N_3757,N_4446);
xnor U16223 (N_16223,N_6364,N_4107);
or U16224 (N_16224,N_8690,N_7824);
xnor U16225 (N_16225,N_9778,N_3570);
nand U16226 (N_16226,N_8318,N_1876);
and U16227 (N_16227,N_1216,N_254);
nor U16228 (N_16228,N_6354,N_1513);
nor U16229 (N_16229,N_5851,N_6640);
and U16230 (N_16230,N_7092,N_4162);
nand U16231 (N_16231,N_271,N_5814);
or U16232 (N_16232,N_6575,N_1707);
xnor U16233 (N_16233,N_7750,N_6056);
or U16234 (N_16234,N_8007,N_5739);
nor U16235 (N_16235,N_2025,N_3993);
xor U16236 (N_16236,N_8680,N_3504);
xor U16237 (N_16237,N_7032,N_8914);
and U16238 (N_16238,N_6301,N_3008);
nor U16239 (N_16239,N_2486,N_80);
or U16240 (N_16240,N_7291,N_3557);
nor U16241 (N_16241,N_3888,N_4844);
and U16242 (N_16242,N_9789,N_944);
nand U16243 (N_16243,N_5278,N_1940);
nor U16244 (N_16244,N_502,N_2006);
xor U16245 (N_16245,N_424,N_4892);
nand U16246 (N_16246,N_7830,N_4902);
xnor U16247 (N_16247,N_5032,N_7663);
nand U16248 (N_16248,N_6755,N_3547);
nand U16249 (N_16249,N_2170,N_7579);
and U16250 (N_16250,N_2250,N_2517);
or U16251 (N_16251,N_6691,N_7167);
and U16252 (N_16252,N_1343,N_6732);
xnor U16253 (N_16253,N_1011,N_8158);
nor U16254 (N_16254,N_942,N_1692);
nor U16255 (N_16255,N_4232,N_5691);
nor U16256 (N_16256,N_2831,N_9520);
nor U16257 (N_16257,N_9297,N_1877);
xor U16258 (N_16258,N_1131,N_9451);
and U16259 (N_16259,N_957,N_7668);
xor U16260 (N_16260,N_1620,N_8556);
and U16261 (N_16261,N_2300,N_2575);
nand U16262 (N_16262,N_4965,N_6557);
nor U16263 (N_16263,N_1781,N_5315);
and U16264 (N_16264,N_1823,N_6099);
nor U16265 (N_16265,N_5945,N_1082);
nor U16266 (N_16266,N_2583,N_31);
nor U16267 (N_16267,N_792,N_8980);
nand U16268 (N_16268,N_1684,N_2052);
and U16269 (N_16269,N_2001,N_3978);
and U16270 (N_16270,N_7202,N_4063);
or U16271 (N_16271,N_4236,N_233);
and U16272 (N_16272,N_538,N_5000);
xor U16273 (N_16273,N_8639,N_1073);
nor U16274 (N_16274,N_4051,N_3834);
and U16275 (N_16275,N_5740,N_6702);
or U16276 (N_16276,N_1835,N_6501);
or U16277 (N_16277,N_5387,N_3808);
xnor U16278 (N_16278,N_418,N_9960);
nor U16279 (N_16279,N_942,N_2795);
nand U16280 (N_16280,N_6350,N_8294);
xor U16281 (N_16281,N_7876,N_8430);
xor U16282 (N_16282,N_714,N_6930);
xnor U16283 (N_16283,N_3306,N_6617);
and U16284 (N_16284,N_5920,N_3985);
nand U16285 (N_16285,N_1649,N_7042);
and U16286 (N_16286,N_7468,N_1508);
and U16287 (N_16287,N_1684,N_463);
nand U16288 (N_16288,N_8904,N_5699);
nand U16289 (N_16289,N_2176,N_7403);
nand U16290 (N_16290,N_5254,N_8697);
xor U16291 (N_16291,N_19,N_6242);
nand U16292 (N_16292,N_1021,N_597);
and U16293 (N_16293,N_6552,N_195);
xnor U16294 (N_16294,N_2214,N_1419);
nor U16295 (N_16295,N_3521,N_4033);
xor U16296 (N_16296,N_6159,N_4168);
nor U16297 (N_16297,N_3668,N_6315);
and U16298 (N_16298,N_5970,N_2565);
nand U16299 (N_16299,N_5872,N_8803);
nor U16300 (N_16300,N_6105,N_8881);
xnor U16301 (N_16301,N_3846,N_3987);
nor U16302 (N_16302,N_4400,N_997);
nand U16303 (N_16303,N_6019,N_2494);
xnor U16304 (N_16304,N_869,N_7063);
or U16305 (N_16305,N_1144,N_5050);
or U16306 (N_16306,N_6336,N_9713);
or U16307 (N_16307,N_4487,N_7861);
and U16308 (N_16308,N_5685,N_6448);
nand U16309 (N_16309,N_756,N_1003);
nor U16310 (N_16310,N_8026,N_9126);
xor U16311 (N_16311,N_3567,N_2518);
or U16312 (N_16312,N_6614,N_5131);
xnor U16313 (N_16313,N_5361,N_7691);
or U16314 (N_16314,N_1353,N_4195);
xor U16315 (N_16315,N_3493,N_549);
and U16316 (N_16316,N_8391,N_755);
or U16317 (N_16317,N_8993,N_1070);
or U16318 (N_16318,N_4128,N_2137);
xor U16319 (N_16319,N_1174,N_8683);
nand U16320 (N_16320,N_2589,N_410);
or U16321 (N_16321,N_623,N_4605);
xnor U16322 (N_16322,N_8349,N_5655);
or U16323 (N_16323,N_9370,N_1748);
and U16324 (N_16324,N_8661,N_5753);
nand U16325 (N_16325,N_6090,N_5539);
or U16326 (N_16326,N_5106,N_8101);
nor U16327 (N_16327,N_9721,N_1197);
xnor U16328 (N_16328,N_6128,N_2186);
or U16329 (N_16329,N_7827,N_7911);
or U16330 (N_16330,N_3192,N_2795);
and U16331 (N_16331,N_580,N_5642);
xor U16332 (N_16332,N_9011,N_9776);
and U16333 (N_16333,N_1201,N_6558);
nand U16334 (N_16334,N_957,N_9095);
xnor U16335 (N_16335,N_3658,N_9793);
or U16336 (N_16336,N_467,N_4710);
xor U16337 (N_16337,N_5436,N_422);
nand U16338 (N_16338,N_6187,N_5673);
nor U16339 (N_16339,N_9732,N_3874);
and U16340 (N_16340,N_1906,N_2376);
or U16341 (N_16341,N_1731,N_1302);
nor U16342 (N_16342,N_9439,N_9876);
xor U16343 (N_16343,N_3259,N_6341);
or U16344 (N_16344,N_4787,N_4399);
and U16345 (N_16345,N_5849,N_5907);
and U16346 (N_16346,N_829,N_6370);
xor U16347 (N_16347,N_7138,N_5172);
xnor U16348 (N_16348,N_5293,N_9206);
and U16349 (N_16349,N_840,N_5396);
or U16350 (N_16350,N_8784,N_2234);
nor U16351 (N_16351,N_2162,N_7296);
and U16352 (N_16352,N_6975,N_3136);
xor U16353 (N_16353,N_4670,N_930);
xor U16354 (N_16354,N_3296,N_3083);
nand U16355 (N_16355,N_7216,N_7408);
and U16356 (N_16356,N_7939,N_2413);
and U16357 (N_16357,N_9467,N_4634);
and U16358 (N_16358,N_2428,N_6940);
nor U16359 (N_16359,N_657,N_7535);
nand U16360 (N_16360,N_7104,N_5537);
nor U16361 (N_16361,N_5267,N_5490);
or U16362 (N_16362,N_4587,N_764);
and U16363 (N_16363,N_351,N_885);
or U16364 (N_16364,N_8608,N_9609);
and U16365 (N_16365,N_6855,N_9331);
nand U16366 (N_16366,N_2827,N_457);
or U16367 (N_16367,N_7300,N_7065);
nor U16368 (N_16368,N_4097,N_6062);
nor U16369 (N_16369,N_9497,N_2780);
nor U16370 (N_16370,N_7577,N_8918);
xor U16371 (N_16371,N_7903,N_9484);
or U16372 (N_16372,N_1027,N_6155);
nor U16373 (N_16373,N_6879,N_6986);
nor U16374 (N_16374,N_8568,N_4604);
or U16375 (N_16375,N_3896,N_2545);
nor U16376 (N_16376,N_2419,N_7674);
or U16377 (N_16377,N_6437,N_8491);
and U16378 (N_16378,N_4407,N_9113);
and U16379 (N_16379,N_5142,N_5531);
nor U16380 (N_16380,N_9000,N_3157);
and U16381 (N_16381,N_5689,N_1573);
nor U16382 (N_16382,N_4292,N_6225);
nor U16383 (N_16383,N_7140,N_7718);
or U16384 (N_16384,N_4712,N_1653);
or U16385 (N_16385,N_8043,N_9045);
and U16386 (N_16386,N_9641,N_5311);
nand U16387 (N_16387,N_8634,N_8711);
nand U16388 (N_16388,N_61,N_3467);
nor U16389 (N_16389,N_653,N_6440);
and U16390 (N_16390,N_2805,N_8774);
or U16391 (N_16391,N_6819,N_249);
or U16392 (N_16392,N_7,N_899);
and U16393 (N_16393,N_240,N_4403);
nand U16394 (N_16394,N_4776,N_9118);
and U16395 (N_16395,N_8193,N_4675);
xor U16396 (N_16396,N_2303,N_6856);
nand U16397 (N_16397,N_7160,N_9549);
xnor U16398 (N_16398,N_8793,N_7009);
xor U16399 (N_16399,N_4726,N_7526);
or U16400 (N_16400,N_7850,N_3454);
or U16401 (N_16401,N_2791,N_7963);
xnor U16402 (N_16402,N_8368,N_3977);
xor U16403 (N_16403,N_3465,N_1022);
nand U16404 (N_16404,N_5649,N_1252);
xor U16405 (N_16405,N_6310,N_2122);
xnor U16406 (N_16406,N_6643,N_601);
xor U16407 (N_16407,N_5681,N_2018);
xor U16408 (N_16408,N_1461,N_7303);
or U16409 (N_16409,N_7330,N_9187);
nand U16410 (N_16410,N_8664,N_7079);
or U16411 (N_16411,N_1656,N_916);
nor U16412 (N_16412,N_7237,N_9776);
nor U16413 (N_16413,N_9799,N_5538);
and U16414 (N_16414,N_7547,N_9899);
or U16415 (N_16415,N_6046,N_8526);
or U16416 (N_16416,N_3482,N_3526);
nor U16417 (N_16417,N_4614,N_8434);
or U16418 (N_16418,N_5441,N_3366);
nand U16419 (N_16419,N_5952,N_6761);
nor U16420 (N_16420,N_2436,N_9017);
and U16421 (N_16421,N_5436,N_6554);
and U16422 (N_16422,N_4394,N_7327);
or U16423 (N_16423,N_2427,N_3896);
xor U16424 (N_16424,N_389,N_2928);
and U16425 (N_16425,N_4085,N_4498);
or U16426 (N_16426,N_7734,N_9549);
and U16427 (N_16427,N_3832,N_5716);
and U16428 (N_16428,N_1879,N_5153);
and U16429 (N_16429,N_763,N_7464);
nor U16430 (N_16430,N_9040,N_6415);
and U16431 (N_16431,N_9818,N_584);
nor U16432 (N_16432,N_9730,N_254);
nand U16433 (N_16433,N_9602,N_3948);
nand U16434 (N_16434,N_1739,N_2720);
and U16435 (N_16435,N_7920,N_2654);
nor U16436 (N_16436,N_7717,N_5720);
or U16437 (N_16437,N_2082,N_9829);
and U16438 (N_16438,N_4046,N_9513);
or U16439 (N_16439,N_1107,N_600);
and U16440 (N_16440,N_5093,N_342);
xnor U16441 (N_16441,N_1918,N_9801);
nor U16442 (N_16442,N_331,N_4792);
and U16443 (N_16443,N_9338,N_4769);
nand U16444 (N_16444,N_6179,N_221);
and U16445 (N_16445,N_4696,N_9256);
or U16446 (N_16446,N_2605,N_3955);
xor U16447 (N_16447,N_1309,N_5831);
and U16448 (N_16448,N_6746,N_2586);
or U16449 (N_16449,N_9261,N_7691);
xor U16450 (N_16450,N_1044,N_9960);
or U16451 (N_16451,N_5979,N_3112);
nor U16452 (N_16452,N_9259,N_6217);
nand U16453 (N_16453,N_4479,N_8658);
nor U16454 (N_16454,N_5614,N_4939);
xor U16455 (N_16455,N_2859,N_7118);
or U16456 (N_16456,N_374,N_3045);
nor U16457 (N_16457,N_8364,N_9851);
nor U16458 (N_16458,N_3286,N_530);
nor U16459 (N_16459,N_6952,N_641);
nor U16460 (N_16460,N_8116,N_4459);
nor U16461 (N_16461,N_2752,N_8828);
nand U16462 (N_16462,N_3264,N_7222);
or U16463 (N_16463,N_9201,N_6733);
nor U16464 (N_16464,N_5168,N_366);
and U16465 (N_16465,N_1341,N_7907);
xnor U16466 (N_16466,N_9178,N_118);
or U16467 (N_16467,N_1890,N_8501);
xnor U16468 (N_16468,N_1432,N_7345);
nand U16469 (N_16469,N_9239,N_6722);
nand U16470 (N_16470,N_4974,N_9213);
or U16471 (N_16471,N_2406,N_162);
xnor U16472 (N_16472,N_9360,N_2039);
nand U16473 (N_16473,N_1364,N_7494);
or U16474 (N_16474,N_4379,N_1014);
and U16475 (N_16475,N_9126,N_8346);
or U16476 (N_16476,N_4701,N_8459);
nand U16477 (N_16477,N_6488,N_4170);
and U16478 (N_16478,N_4643,N_7883);
nand U16479 (N_16479,N_862,N_4688);
nor U16480 (N_16480,N_3393,N_6707);
nand U16481 (N_16481,N_5356,N_1175);
and U16482 (N_16482,N_8805,N_2392);
nor U16483 (N_16483,N_3779,N_2169);
or U16484 (N_16484,N_3120,N_7568);
xor U16485 (N_16485,N_7627,N_2066);
or U16486 (N_16486,N_7500,N_4766);
and U16487 (N_16487,N_9166,N_2602);
nand U16488 (N_16488,N_2210,N_4496);
and U16489 (N_16489,N_3791,N_6192);
nand U16490 (N_16490,N_2832,N_8260);
nor U16491 (N_16491,N_5540,N_1034);
or U16492 (N_16492,N_9186,N_1098);
and U16493 (N_16493,N_4272,N_9328);
and U16494 (N_16494,N_2659,N_3810);
or U16495 (N_16495,N_6114,N_8950);
and U16496 (N_16496,N_2650,N_8345);
and U16497 (N_16497,N_6557,N_6363);
and U16498 (N_16498,N_5658,N_8313);
and U16499 (N_16499,N_4467,N_3858);
and U16500 (N_16500,N_515,N_534);
nor U16501 (N_16501,N_1767,N_2152);
and U16502 (N_16502,N_5993,N_2607);
or U16503 (N_16503,N_7257,N_397);
nor U16504 (N_16504,N_4540,N_4381);
nor U16505 (N_16505,N_2717,N_4755);
or U16506 (N_16506,N_881,N_601);
or U16507 (N_16507,N_9041,N_6965);
nor U16508 (N_16508,N_3016,N_2620);
or U16509 (N_16509,N_2498,N_5064);
or U16510 (N_16510,N_2630,N_2530);
xnor U16511 (N_16511,N_1799,N_8669);
or U16512 (N_16512,N_297,N_8196);
nor U16513 (N_16513,N_3651,N_1477);
xor U16514 (N_16514,N_5591,N_3506);
nand U16515 (N_16515,N_879,N_4188);
nor U16516 (N_16516,N_5789,N_8615);
or U16517 (N_16517,N_8363,N_4161);
xor U16518 (N_16518,N_5422,N_4927);
and U16519 (N_16519,N_2536,N_8439);
and U16520 (N_16520,N_3845,N_9572);
or U16521 (N_16521,N_8413,N_7462);
or U16522 (N_16522,N_8564,N_8521);
nand U16523 (N_16523,N_8680,N_3657);
and U16524 (N_16524,N_7498,N_1860);
nor U16525 (N_16525,N_998,N_6448);
nor U16526 (N_16526,N_1784,N_5335);
or U16527 (N_16527,N_3962,N_8753);
nand U16528 (N_16528,N_8145,N_8894);
nor U16529 (N_16529,N_7406,N_3354);
xor U16530 (N_16530,N_7269,N_3354);
or U16531 (N_16531,N_5180,N_263);
or U16532 (N_16532,N_9591,N_4232);
nor U16533 (N_16533,N_7708,N_6754);
or U16534 (N_16534,N_449,N_4);
nand U16535 (N_16535,N_4843,N_9780);
nand U16536 (N_16536,N_5630,N_8758);
nor U16537 (N_16537,N_5034,N_7840);
or U16538 (N_16538,N_7663,N_1541);
xor U16539 (N_16539,N_296,N_1057);
or U16540 (N_16540,N_400,N_4745);
or U16541 (N_16541,N_7017,N_3048);
nor U16542 (N_16542,N_6382,N_7113);
nor U16543 (N_16543,N_4146,N_7097);
or U16544 (N_16544,N_4147,N_762);
nand U16545 (N_16545,N_8665,N_2665);
xnor U16546 (N_16546,N_1443,N_6812);
or U16547 (N_16547,N_6108,N_1218);
xor U16548 (N_16548,N_471,N_841);
nand U16549 (N_16549,N_9465,N_3469);
nor U16550 (N_16550,N_4422,N_2166);
nand U16551 (N_16551,N_2098,N_6296);
xnor U16552 (N_16552,N_9647,N_7016);
or U16553 (N_16553,N_7109,N_8243);
nand U16554 (N_16554,N_714,N_4515);
nor U16555 (N_16555,N_6859,N_644);
nor U16556 (N_16556,N_3798,N_3217);
nor U16557 (N_16557,N_7131,N_8621);
nor U16558 (N_16558,N_9364,N_5066);
nand U16559 (N_16559,N_8131,N_6137);
xor U16560 (N_16560,N_6628,N_7202);
xor U16561 (N_16561,N_3389,N_7688);
or U16562 (N_16562,N_2599,N_8009);
nor U16563 (N_16563,N_3716,N_6034);
or U16564 (N_16564,N_5251,N_467);
and U16565 (N_16565,N_976,N_7298);
nor U16566 (N_16566,N_1254,N_5507);
nor U16567 (N_16567,N_8661,N_9613);
and U16568 (N_16568,N_2309,N_4174);
nor U16569 (N_16569,N_5157,N_6348);
and U16570 (N_16570,N_3652,N_1597);
xor U16571 (N_16571,N_146,N_9725);
xor U16572 (N_16572,N_373,N_6402);
nor U16573 (N_16573,N_4976,N_398);
or U16574 (N_16574,N_2255,N_8321);
nand U16575 (N_16575,N_4281,N_8983);
nand U16576 (N_16576,N_1744,N_9463);
xnor U16577 (N_16577,N_174,N_5503);
nand U16578 (N_16578,N_8325,N_1057);
xor U16579 (N_16579,N_5971,N_8521);
nand U16580 (N_16580,N_4293,N_8191);
and U16581 (N_16581,N_4198,N_1425);
and U16582 (N_16582,N_5910,N_7562);
and U16583 (N_16583,N_5315,N_5796);
and U16584 (N_16584,N_16,N_7388);
nand U16585 (N_16585,N_8173,N_5720);
nand U16586 (N_16586,N_5089,N_1322);
nor U16587 (N_16587,N_8210,N_9013);
or U16588 (N_16588,N_537,N_7708);
or U16589 (N_16589,N_347,N_9720);
and U16590 (N_16590,N_4433,N_5689);
nand U16591 (N_16591,N_4933,N_1336);
nor U16592 (N_16592,N_8140,N_407);
xnor U16593 (N_16593,N_7192,N_1646);
and U16594 (N_16594,N_8471,N_646);
nor U16595 (N_16595,N_1061,N_4253);
nand U16596 (N_16596,N_8297,N_8787);
and U16597 (N_16597,N_2930,N_9819);
or U16598 (N_16598,N_5498,N_9854);
xnor U16599 (N_16599,N_4487,N_4703);
xor U16600 (N_16600,N_9503,N_6818);
xnor U16601 (N_16601,N_9716,N_8480);
nor U16602 (N_16602,N_9046,N_4091);
xnor U16603 (N_16603,N_2797,N_3346);
nand U16604 (N_16604,N_9243,N_9485);
or U16605 (N_16605,N_8,N_912);
or U16606 (N_16606,N_8831,N_4647);
nor U16607 (N_16607,N_5627,N_616);
xor U16608 (N_16608,N_7053,N_7069);
and U16609 (N_16609,N_4361,N_9879);
nand U16610 (N_16610,N_2290,N_1421);
nand U16611 (N_16611,N_7453,N_4118);
nand U16612 (N_16612,N_195,N_4294);
and U16613 (N_16613,N_8004,N_1208);
xor U16614 (N_16614,N_6143,N_4984);
xnor U16615 (N_16615,N_3957,N_8406);
or U16616 (N_16616,N_1886,N_1371);
nand U16617 (N_16617,N_9592,N_7018);
nor U16618 (N_16618,N_9372,N_3057);
and U16619 (N_16619,N_676,N_2496);
xor U16620 (N_16620,N_4596,N_2059);
xnor U16621 (N_16621,N_4368,N_109);
nor U16622 (N_16622,N_1775,N_9958);
nor U16623 (N_16623,N_1740,N_5418);
nand U16624 (N_16624,N_356,N_4056);
nand U16625 (N_16625,N_9530,N_9018);
nand U16626 (N_16626,N_8548,N_7322);
nand U16627 (N_16627,N_6836,N_7597);
nor U16628 (N_16628,N_2053,N_1055);
nand U16629 (N_16629,N_1757,N_9711);
or U16630 (N_16630,N_7977,N_8764);
nand U16631 (N_16631,N_3191,N_6465);
and U16632 (N_16632,N_3468,N_2726);
or U16633 (N_16633,N_6595,N_5672);
xor U16634 (N_16634,N_8023,N_7203);
and U16635 (N_16635,N_2506,N_2173);
nor U16636 (N_16636,N_3057,N_9615);
nand U16637 (N_16637,N_28,N_7210);
or U16638 (N_16638,N_9378,N_8206);
xnor U16639 (N_16639,N_2199,N_7856);
xor U16640 (N_16640,N_3368,N_3953);
or U16641 (N_16641,N_5139,N_7661);
nor U16642 (N_16642,N_4093,N_9169);
and U16643 (N_16643,N_296,N_9662);
nor U16644 (N_16644,N_4732,N_4272);
xor U16645 (N_16645,N_6615,N_68);
nand U16646 (N_16646,N_9726,N_9849);
or U16647 (N_16647,N_5955,N_5698);
nor U16648 (N_16648,N_3504,N_2460);
nor U16649 (N_16649,N_7562,N_373);
and U16650 (N_16650,N_9196,N_6384);
nand U16651 (N_16651,N_861,N_3899);
nor U16652 (N_16652,N_669,N_1509);
nand U16653 (N_16653,N_696,N_1173);
nor U16654 (N_16654,N_37,N_9285);
nand U16655 (N_16655,N_458,N_3215);
and U16656 (N_16656,N_9153,N_3769);
nor U16657 (N_16657,N_4282,N_9560);
or U16658 (N_16658,N_1361,N_4526);
or U16659 (N_16659,N_4052,N_7486);
nand U16660 (N_16660,N_210,N_8014);
nor U16661 (N_16661,N_3316,N_7682);
xor U16662 (N_16662,N_3278,N_1347);
nor U16663 (N_16663,N_6389,N_8332);
xor U16664 (N_16664,N_9393,N_8031);
xor U16665 (N_16665,N_9365,N_5241);
nor U16666 (N_16666,N_2275,N_788);
xor U16667 (N_16667,N_6134,N_6896);
nor U16668 (N_16668,N_4749,N_881);
or U16669 (N_16669,N_7729,N_5680);
and U16670 (N_16670,N_5899,N_2000);
xor U16671 (N_16671,N_5554,N_5193);
and U16672 (N_16672,N_9225,N_7352);
nand U16673 (N_16673,N_6184,N_4013);
nand U16674 (N_16674,N_5386,N_6703);
nand U16675 (N_16675,N_1955,N_1515);
xnor U16676 (N_16676,N_5409,N_9853);
nor U16677 (N_16677,N_6230,N_3252);
xnor U16678 (N_16678,N_5039,N_8870);
nor U16679 (N_16679,N_3128,N_5029);
nor U16680 (N_16680,N_3311,N_1714);
xnor U16681 (N_16681,N_5150,N_6042);
or U16682 (N_16682,N_5242,N_7243);
nand U16683 (N_16683,N_8087,N_4679);
nand U16684 (N_16684,N_6216,N_7914);
nor U16685 (N_16685,N_2939,N_9433);
and U16686 (N_16686,N_8644,N_4644);
nor U16687 (N_16687,N_8991,N_9990);
nand U16688 (N_16688,N_8459,N_5392);
or U16689 (N_16689,N_3787,N_6703);
or U16690 (N_16690,N_947,N_5160);
and U16691 (N_16691,N_5474,N_3201);
xnor U16692 (N_16692,N_1335,N_9774);
xor U16693 (N_16693,N_3583,N_6752);
nand U16694 (N_16694,N_8193,N_7736);
or U16695 (N_16695,N_5808,N_9511);
or U16696 (N_16696,N_1938,N_5065);
nor U16697 (N_16697,N_1420,N_2481);
nor U16698 (N_16698,N_8920,N_4356);
xor U16699 (N_16699,N_4514,N_4411);
or U16700 (N_16700,N_3618,N_4220);
nor U16701 (N_16701,N_3729,N_7365);
nor U16702 (N_16702,N_9774,N_1452);
and U16703 (N_16703,N_7309,N_9928);
xnor U16704 (N_16704,N_1696,N_1434);
xor U16705 (N_16705,N_8945,N_6400);
xnor U16706 (N_16706,N_2711,N_7070);
nor U16707 (N_16707,N_9405,N_7319);
xnor U16708 (N_16708,N_8573,N_6127);
or U16709 (N_16709,N_3581,N_4665);
xnor U16710 (N_16710,N_5355,N_8947);
nor U16711 (N_16711,N_1403,N_217);
xnor U16712 (N_16712,N_6773,N_5320);
nor U16713 (N_16713,N_1672,N_4597);
or U16714 (N_16714,N_4174,N_1106);
xnor U16715 (N_16715,N_9187,N_4161);
or U16716 (N_16716,N_6336,N_8266);
or U16717 (N_16717,N_1321,N_3981);
or U16718 (N_16718,N_1552,N_6241);
nand U16719 (N_16719,N_7327,N_7909);
xnor U16720 (N_16720,N_2996,N_2531);
xnor U16721 (N_16721,N_7194,N_559);
nor U16722 (N_16722,N_1218,N_119);
and U16723 (N_16723,N_6811,N_1687);
and U16724 (N_16724,N_9127,N_6299);
and U16725 (N_16725,N_2758,N_9934);
nand U16726 (N_16726,N_4645,N_493);
xnor U16727 (N_16727,N_2475,N_397);
nor U16728 (N_16728,N_2603,N_3443);
nor U16729 (N_16729,N_6811,N_3429);
nand U16730 (N_16730,N_6183,N_7811);
xor U16731 (N_16731,N_9874,N_1596);
or U16732 (N_16732,N_1954,N_4395);
nand U16733 (N_16733,N_9065,N_9051);
xor U16734 (N_16734,N_5856,N_4826);
or U16735 (N_16735,N_2246,N_2536);
or U16736 (N_16736,N_9110,N_1729);
and U16737 (N_16737,N_8087,N_8567);
nand U16738 (N_16738,N_7841,N_1392);
or U16739 (N_16739,N_4807,N_2462);
nand U16740 (N_16740,N_7352,N_7069);
nor U16741 (N_16741,N_2372,N_6180);
xnor U16742 (N_16742,N_645,N_6725);
nor U16743 (N_16743,N_6157,N_7848);
or U16744 (N_16744,N_6676,N_2367);
or U16745 (N_16745,N_5203,N_8907);
nor U16746 (N_16746,N_2593,N_821);
xor U16747 (N_16747,N_5276,N_4194);
xor U16748 (N_16748,N_828,N_8736);
nor U16749 (N_16749,N_7311,N_1795);
xor U16750 (N_16750,N_5610,N_5668);
nor U16751 (N_16751,N_2313,N_168);
nor U16752 (N_16752,N_312,N_7313);
and U16753 (N_16753,N_9543,N_3628);
and U16754 (N_16754,N_6304,N_1249);
or U16755 (N_16755,N_9433,N_9253);
and U16756 (N_16756,N_6972,N_6494);
nor U16757 (N_16757,N_1271,N_8056);
nand U16758 (N_16758,N_2204,N_7573);
nand U16759 (N_16759,N_7825,N_5385);
xnor U16760 (N_16760,N_8964,N_5129);
or U16761 (N_16761,N_334,N_5);
and U16762 (N_16762,N_2213,N_7936);
and U16763 (N_16763,N_4488,N_7474);
nor U16764 (N_16764,N_3382,N_713);
nor U16765 (N_16765,N_638,N_5025);
or U16766 (N_16766,N_4958,N_1753);
nand U16767 (N_16767,N_5275,N_706);
and U16768 (N_16768,N_1363,N_9045);
xor U16769 (N_16769,N_7494,N_3243);
nand U16770 (N_16770,N_7747,N_2420);
nand U16771 (N_16771,N_6374,N_4382);
and U16772 (N_16772,N_6970,N_8988);
xor U16773 (N_16773,N_3460,N_4081);
or U16774 (N_16774,N_7075,N_808);
or U16775 (N_16775,N_6118,N_2029);
and U16776 (N_16776,N_414,N_2937);
and U16777 (N_16777,N_7487,N_2854);
xnor U16778 (N_16778,N_933,N_9617);
nand U16779 (N_16779,N_6207,N_5870);
nor U16780 (N_16780,N_4766,N_669);
or U16781 (N_16781,N_4932,N_4279);
nand U16782 (N_16782,N_2817,N_3858);
and U16783 (N_16783,N_3877,N_2848);
xor U16784 (N_16784,N_9744,N_7203);
nand U16785 (N_16785,N_8674,N_375);
nor U16786 (N_16786,N_8459,N_9416);
and U16787 (N_16787,N_2413,N_9590);
and U16788 (N_16788,N_7736,N_1558);
nor U16789 (N_16789,N_9858,N_8187);
or U16790 (N_16790,N_3169,N_1064);
nand U16791 (N_16791,N_8634,N_6804);
or U16792 (N_16792,N_1809,N_5194);
or U16793 (N_16793,N_9635,N_4399);
and U16794 (N_16794,N_1506,N_9821);
or U16795 (N_16795,N_2865,N_842);
xor U16796 (N_16796,N_9290,N_6178);
nand U16797 (N_16797,N_5168,N_9693);
or U16798 (N_16798,N_8623,N_5640);
xor U16799 (N_16799,N_8214,N_6750);
or U16800 (N_16800,N_4971,N_9476);
nor U16801 (N_16801,N_3716,N_4275);
nor U16802 (N_16802,N_9113,N_4230);
nor U16803 (N_16803,N_9115,N_8733);
xor U16804 (N_16804,N_9413,N_2584);
and U16805 (N_16805,N_8684,N_9649);
or U16806 (N_16806,N_5086,N_3099);
and U16807 (N_16807,N_9061,N_9756);
or U16808 (N_16808,N_4476,N_4941);
nand U16809 (N_16809,N_8732,N_1169);
nand U16810 (N_16810,N_6577,N_7307);
nor U16811 (N_16811,N_1543,N_780);
nand U16812 (N_16812,N_6657,N_4625);
nand U16813 (N_16813,N_7722,N_1206);
xor U16814 (N_16814,N_7660,N_4225);
nor U16815 (N_16815,N_3736,N_8100);
nand U16816 (N_16816,N_3072,N_3739);
xnor U16817 (N_16817,N_3456,N_934);
nor U16818 (N_16818,N_8436,N_686);
nor U16819 (N_16819,N_6384,N_4053);
and U16820 (N_16820,N_3921,N_5896);
or U16821 (N_16821,N_1009,N_6506);
nand U16822 (N_16822,N_3966,N_2645);
and U16823 (N_16823,N_7181,N_304);
nand U16824 (N_16824,N_9993,N_7038);
nand U16825 (N_16825,N_1848,N_4331);
and U16826 (N_16826,N_7178,N_377);
and U16827 (N_16827,N_573,N_7294);
nand U16828 (N_16828,N_1342,N_7865);
nor U16829 (N_16829,N_5385,N_944);
xor U16830 (N_16830,N_362,N_488);
or U16831 (N_16831,N_9454,N_3704);
nand U16832 (N_16832,N_7831,N_8743);
or U16833 (N_16833,N_3244,N_2520);
or U16834 (N_16834,N_8746,N_871);
and U16835 (N_16835,N_2223,N_9657);
nand U16836 (N_16836,N_9598,N_479);
xnor U16837 (N_16837,N_441,N_6161);
nor U16838 (N_16838,N_7820,N_320);
nor U16839 (N_16839,N_1865,N_1166);
nand U16840 (N_16840,N_9950,N_665);
nand U16841 (N_16841,N_3608,N_9662);
and U16842 (N_16842,N_1690,N_4243);
or U16843 (N_16843,N_2470,N_7784);
or U16844 (N_16844,N_6009,N_3973);
nand U16845 (N_16845,N_7053,N_8371);
or U16846 (N_16846,N_2997,N_1143);
nor U16847 (N_16847,N_6294,N_4595);
xnor U16848 (N_16848,N_767,N_848);
nand U16849 (N_16849,N_3776,N_4902);
or U16850 (N_16850,N_2239,N_877);
xor U16851 (N_16851,N_8454,N_2429);
and U16852 (N_16852,N_2477,N_2563);
xor U16853 (N_16853,N_9337,N_5141);
or U16854 (N_16854,N_934,N_1336);
nand U16855 (N_16855,N_1666,N_9592);
nor U16856 (N_16856,N_5834,N_8887);
nand U16857 (N_16857,N_2993,N_5014);
nand U16858 (N_16858,N_4723,N_6081);
xnor U16859 (N_16859,N_2381,N_5889);
xor U16860 (N_16860,N_8065,N_7159);
and U16861 (N_16861,N_7128,N_1575);
or U16862 (N_16862,N_9802,N_2952);
and U16863 (N_16863,N_9206,N_7468);
or U16864 (N_16864,N_1384,N_247);
nand U16865 (N_16865,N_8482,N_3033);
or U16866 (N_16866,N_9308,N_6258);
or U16867 (N_16867,N_3787,N_1113);
and U16868 (N_16868,N_6255,N_7666);
nand U16869 (N_16869,N_3856,N_9661);
nor U16870 (N_16870,N_8490,N_1934);
or U16871 (N_16871,N_2684,N_725);
nand U16872 (N_16872,N_5512,N_3198);
xnor U16873 (N_16873,N_5608,N_6888);
nor U16874 (N_16874,N_8,N_2500);
and U16875 (N_16875,N_9536,N_602);
or U16876 (N_16876,N_9914,N_4963);
xor U16877 (N_16877,N_7146,N_2658);
xnor U16878 (N_16878,N_9455,N_5766);
nor U16879 (N_16879,N_2752,N_5520);
xor U16880 (N_16880,N_6290,N_6910);
and U16881 (N_16881,N_8370,N_3035);
xnor U16882 (N_16882,N_9618,N_4758);
xnor U16883 (N_16883,N_9956,N_6312);
and U16884 (N_16884,N_3491,N_6171);
xnor U16885 (N_16885,N_8915,N_9652);
xor U16886 (N_16886,N_7940,N_6932);
or U16887 (N_16887,N_8111,N_5795);
and U16888 (N_16888,N_7928,N_8998);
nand U16889 (N_16889,N_3269,N_9193);
nor U16890 (N_16890,N_4930,N_1270);
nand U16891 (N_16891,N_6233,N_4756);
xor U16892 (N_16892,N_8402,N_5384);
or U16893 (N_16893,N_6705,N_1463);
and U16894 (N_16894,N_4566,N_7852);
nor U16895 (N_16895,N_9633,N_3596);
or U16896 (N_16896,N_4457,N_200);
or U16897 (N_16897,N_887,N_9198);
and U16898 (N_16898,N_1999,N_6368);
nand U16899 (N_16899,N_4603,N_393);
or U16900 (N_16900,N_5892,N_1415);
xnor U16901 (N_16901,N_2252,N_8241);
or U16902 (N_16902,N_249,N_8819);
or U16903 (N_16903,N_8154,N_9330);
xnor U16904 (N_16904,N_9097,N_1511);
xor U16905 (N_16905,N_1191,N_9831);
nor U16906 (N_16906,N_5529,N_4256);
or U16907 (N_16907,N_7554,N_114);
nor U16908 (N_16908,N_4520,N_8926);
or U16909 (N_16909,N_2779,N_2652);
nand U16910 (N_16910,N_5685,N_7514);
and U16911 (N_16911,N_8155,N_8041);
and U16912 (N_16912,N_7935,N_276);
or U16913 (N_16913,N_6396,N_5778);
or U16914 (N_16914,N_7500,N_2736);
xnor U16915 (N_16915,N_9015,N_9240);
nor U16916 (N_16916,N_5589,N_5163);
xor U16917 (N_16917,N_6915,N_831);
nand U16918 (N_16918,N_213,N_4508);
xor U16919 (N_16919,N_3820,N_7565);
nor U16920 (N_16920,N_3746,N_600);
xnor U16921 (N_16921,N_2924,N_4739);
nand U16922 (N_16922,N_7320,N_3932);
nand U16923 (N_16923,N_930,N_6034);
nor U16924 (N_16924,N_6769,N_961);
nand U16925 (N_16925,N_9457,N_5105);
xor U16926 (N_16926,N_4274,N_9409);
or U16927 (N_16927,N_1104,N_8403);
xnor U16928 (N_16928,N_1377,N_7627);
nor U16929 (N_16929,N_8813,N_7224);
and U16930 (N_16930,N_4906,N_1925);
nand U16931 (N_16931,N_3949,N_7206);
nor U16932 (N_16932,N_384,N_3182);
and U16933 (N_16933,N_2947,N_1773);
nand U16934 (N_16934,N_2092,N_4738);
nand U16935 (N_16935,N_2268,N_6367);
and U16936 (N_16936,N_7895,N_4368);
xor U16937 (N_16937,N_1516,N_9174);
nor U16938 (N_16938,N_8036,N_3401);
nand U16939 (N_16939,N_5372,N_775);
nor U16940 (N_16940,N_4549,N_4931);
xor U16941 (N_16941,N_5396,N_8843);
or U16942 (N_16942,N_2432,N_3015);
or U16943 (N_16943,N_4644,N_4102);
and U16944 (N_16944,N_2442,N_2146);
and U16945 (N_16945,N_3125,N_4838);
and U16946 (N_16946,N_2630,N_6230);
nor U16947 (N_16947,N_673,N_1704);
or U16948 (N_16948,N_4885,N_9177);
and U16949 (N_16949,N_7953,N_8833);
xor U16950 (N_16950,N_3958,N_4596);
or U16951 (N_16951,N_4086,N_9695);
xor U16952 (N_16952,N_8152,N_115);
or U16953 (N_16953,N_4870,N_7853);
or U16954 (N_16954,N_8211,N_8688);
or U16955 (N_16955,N_9428,N_5970);
nor U16956 (N_16956,N_477,N_1527);
nor U16957 (N_16957,N_9507,N_495);
or U16958 (N_16958,N_7845,N_3783);
or U16959 (N_16959,N_4680,N_9453);
nand U16960 (N_16960,N_3261,N_7155);
or U16961 (N_16961,N_339,N_4438);
or U16962 (N_16962,N_4668,N_2570);
and U16963 (N_16963,N_3555,N_8621);
nor U16964 (N_16964,N_3714,N_2912);
and U16965 (N_16965,N_2662,N_2296);
and U16966 (N_16966,N_3453,N_4151);
and U16967 (N_16967,N_430,N_1438);
nor U16968 (N_16968,N_7129,N_6610);
xor U16969 (N_16969,N_4348,N_2652);
nor U16970 (N_16970,N_9560,N_3771);
and U16971 (N_16971,N_6528,N_8721);
xnor U16972 (N_16972,N_6434,N_4595);
or U16973 (N_16973,N_9364,N_2134);
nand U16974 (N_16974,N_3401,N_273);
and U16975 (N_16975,N_7671,N_4646);
or U16976 (N_16976,N_4715,N_7332);
or U16977 (N_16977,N_6102,N_2748);
and U16978 (N_16978,N_1370,N_4560);
and U16979 (N_16979,N_5989,N_34);
xnor U16980 (N_16980,N_8100,N_9535);
and U16981 (N_16981,N_4870,N_5325);
xnor U16982 (N_16982,N_5076,N_4526);
nor U16983 (N_16983,N_8978,N_676);
nand U16984 (N_16984,N_5268,N_2886);
and U16985 (N_16985,N_5250,N_8074);
xor U16986 (N_16986,N_5139,N_9455);
or U16987 (N_16987,N_6896,N_4509);
xnor U16988 (N_16988,N_5243,N_3011);
nand U16989 (N_16989,N_7781,N_1226);
or U16990 (N_16990,N_4422,N_3542);
and U16991 (N_16991,N_7653,N_9502);
and U16992 (N_16992,N_1835,N_1691);
nand U16993 (N_16993,N_9851,N_9551);
xnor U16994 (N_16994,N_4681,N_9847);
or U16995 (N_16995,N_1447,N_4991);
or U16996 (N_16996,N_374,N_9087);
xnor U16997 (N_16997,N_2663,N_8221);
or U16998 (N_16998,N_5917,N_6495);
nand U16999 (N_16999,N_4808,N_5658);
xor U17000 (N_17000,N_8727,N_8927);
nand U17001 (N_17001,N_4065,N_9439);
nor U17002 (N_17002,N_4914,N_8639);
nor U17003 (N_17003,N_5064,N_7118);
xor U17004 (N_17004,N_2281,N_1340);
nand U17005 (N_17005,N_2130,N_2636);
or U17006 (N_17006,N_298,N_8550);
xor U17007 (N_17007,N_4291,N_3063);
nand U17008 (N_17008,N_8442,N_1650);
and U17009 (N_17009,N_9894,N_6635);
or U17010 (N_17010,N_145,N_8583);
and U17011 (N_17011,N_7782,N_6967);
nand U17012 (N_17012,N_1477,N_312);
nand U17013 (N_17013,N_9456,N_7515);
xor U17014 (N_17014,N_5506,N_8203);
nor U17015 (N_17015,N_4875,N_6217);
or U17016 (N_17016,N_1347,N_4282);
and U17017 (N_17017,N_4841,N_6941);
or U17018 (N_17018,N_7271,N_6309);
nand U17019 (N_17019,N_6676,N_435);
nor U17020 (N_17020,N_812,N_6752);
xor U17021 (N_17021,N_1928,N_5770);
xnor U17022 (N_17022,N_8919,N_1448);
or U17023 (N_17023,N_9455,N_8609);
nor U17024 (N_17024,N_3123,N_1345);
or U17025 (N_17025,N_9578,N_9634);
nor U17026 (N_17026,N_8338,N_9259);
nor U17027 (N_17027,N_2442,N_3570);
xor U17028 (N_17028,N_3225,N_6088);
xnor U17029 (N_17029,N_9170,N_460);
xnor U17030 (N_17030,N_1884,N_5358);
nor U17031 (N_17031,N_2695,N_489);
or U17032 (N_17032,N_6499,N_8711);
or U17033 (N_17033,N_9326,N_1273);
or U17034 (N_17034,N_4523,N_3217);
or U17035 (N_17035,N_3831,N_9560);
and U17036 (N_17036,N_1802,N_606);
nand U17037 (N_17037,N_5893,N_8232);
nand U17038 (N_17038,N_8484,N_3815);
nor U17039 (N_17039,N_892,N_9671);
nand U17040 (N_17040,N_5303,N_6475);
and U17041 (N_17041,N_7406,N_298);
xor U17042 (N_17042,N_9881,N_5072);
nor U17043 (N_17043,N_9465,N_1258);
or U17044 (N_17044,N_2791,N_945);
nor U17045 (N_17045,N_1710,N_4824);
xor U17046 (N_17046,N_9155,N_4036);
or U17047 (N_17047,N_8053,N_1374);
or U17048 (N_17048,N_7336,N_9256);
nor U17049 (N_17049,N_138,N_3296);
nand U17050 (N_17050,N_6641,N_2337);
nor U17051 (N_17051,N_9161,N_1497);
xor U17052 (N_17052,N_8131,N_2027);
and U17053 (N_17053,N_6398,N_1262);
xor U17054 (N_17054,N_6627,N_7266);
or U17055 (N_17055,N_5481,N_1015);
or U17056 (N_17056,N_435,N_7076);
and U17057 (N_17057,N_7651,N_6390);
and U17058 (N_17058,N_8284,N_1252);
and U17059 (N_17059,N_6711,N_6966);
xor U17060 (N_17060,N_5658,N_8784);
and U17061 (N_17061,N_585,N_7980);
xnor U17062 (N_17062,N_2926,N_9337);
nand U17063 (N_17063,N_7430,N_5932);
nand U17064 (N_17064,N_1647,N_2203);
and U17065 (N_17065,N_9954,N_4764);
and U17066 (N_17066,N_6345,N_3196);
or U17067 (N_17067,N_5146,N_7498);
nand U17068 (N_17068,N_6305,N_4328);
and U17069 (N_17069,N_8489,N_8512);
xnor U17070 (N_17070,N_8589,N_3750);
nor U17071 (N_17071,N_425,N_6818);
and U17072 (N_17072,N_4311,N_2371);
and U17073 (N_17073,N_3317,N_2597);
and U17074 (N_17074,N_6088,N_6336);
and U17075 (N_17075,N_783,N_9070);
and U17076 (N_17076,N_9852,N_9491);
nand U17077 (N_17077,N_5594,N_2524);
nor U17078 (N_17078,N_5134,N_1210);
or U17079 (N_17079,N_9913,N_4696);
xor U17080 (N_17080,N_2032,N_7590);
xnor U17081 (N_17081,N_2177,N_1071);
and U17082 (N_17082,N_1406,N_5115);
and U17083 (N_17083,N_5470,N_1619);
nand U17084 (N_17084,N_4371,N_8659);
nand U17085 (N_17085,N_6506,N_7574);
nand U17086 (N_17086,N_1323,N_540);
or U17087 (N_17087,N_5033,N_9279);
xnor U17088 (N_17088,N_3301,N_6551);
nand U17089 (N_17089,N_4761,N_7230);
xnor U17090 (N_17090,N_2457,N_3209);
xnor U17091 (N_17091,N_3378,N_6243);
xnor U17092 (N_17092,N_7344,N_2896);
or U17093 (N_17093,N_3120,N_7939);
and U17094 (N_17094,N_6373,N_4866);
and U17095 (N_17095,N_8035,N_2304);
nand U17096 (N_17096,N_8577,N_5237);
xor U17097 (N_17097,N_4393,N_9588);
xor U17098 (N_17098,N_3898,N_4757);
nor U17099 (N_17099,N_3517,N_9408);
xnor U17100 (N_17100,N_1886,N_5881);
or U17101 (N_17101,N_3235,N_405);
xnor U17102 (N_17102,N_8739,N_4259);
or U17103 (N_17103,N_1198,N_8455);
nor U17104 (N_17104,N_3462,N_7690);
and U17105 (N_17105,N_9171,N_7522);
xor U17106 (N_17106,N_5966,N_1043);
and U17107 (N_17107,N_7197,N_1431);
xor U17108 (N_17108,N_1289,N_1302);
and U17109 (N_17109,N_2410,N_7735);
nor U17110 (N_17110,N_1104,N_5214);
nor U17111 (N_17111,N_1806,N_6735);
and U17112 (N_17112,N_8801,N_8598);
or U17113 (N_17113,N_6450,N_9458);
and U17114 (N_17114,N_9762,N_3344);
nand U17115 (N_17115,N_1998,N_1038);
or U17116 (N_17116,N_7694,N_1280);
nand U17117 (N_17117,N_9189,N_4234);
or U17118 (N_17118,N_24,N_9338);
and U17119 (N_17119,N_5713,N_1598);
and U17120 (N_17120,N_5749,N_512);
nor U17121 (N_17121,N_387,N_6295);
xnor U17122 (N_17122,N_582,N_2410);
nand U17123 (N_17123,N_4479,N_1653);
nor U17124 (N_17124,N_2668,N_5014);
nor U17125 (N_17125,N_4230,N_6666);
and U17126 (N_17126,N_6103,N_9882);
or U17127 (N_17127,N_9226,N_5517);
xnor U17128 (N_17128,N_8441,N_7574);
xor U17129 (N_17129,N_5596,N_5439);
nand U17130 (N_17130,N_1095,N_5999);
nor U17131 (N_17131,N_8849,N_9168);
xnor U17132 (N_17132,N_6786,N_5087);
nor U17133 (N_17133,N_3117,N_9074);
nand U17134 (N_17134,N_5753,N_817);
nor U17135 (N_17135,N_6636,N_7511);
xnor U17136 (N_17136,N_4634,N_8333);
nand U17137 (N_17137,N_3611,N_7403);
and U17138 (N_17138,N_6927,N_1918);
nor U17139 (N_17139,N_9041,N_4739);
and U17140 (N_17140,N_6020,N_3107);
nand U17141 (N_17141,N_6729,N_4870);
or U17142 (N_17142,N_9016,N_8942);
or U17143 (N_17143,N_790,N_7972);
nor U17144 (N_17144,N_3047,N_3681);
nor U17145 (N_17145,N_7669,N_1965);
nand U17146 (N_17146,N_6050,N_1242);
nor U17147 (N_17147,N_1000,N_4947);
and U17148 (N_17148,N_2678,N_6690);
and U17149 (N_17149,N_2259,N_2339);
nand U17150 (N_17150,N_2218,N_6707);
and U17151 (N_17151,N_5546,N_313);
or U17152 (N_17152,N_3209,N_7316);
xnor U17153 (N_17153,N_8734,N_2050);
and U17154 (N_17154,N_435,N_1507);
nand U17155 (N_17155,N_4860,N_7696);
nand U17156 (N_17156,N_3427,N_9700);
nor U17157 (N_17157,N_1173,N_8463);
and U17158 (N_17158,N_590,N_1854);
nor U17159 (N_17159,N_5400,N_3733);
xnor U17160 (N_17160,N_5046,N_5422);
or U17161 (N_17161,N_4468,N_5597);
nor U17162 (N_17162,N_437,N_9373);
nor U17163 (N_17163,N_537,N_1431);
or U17164 (N_17164,N_9577,N_7397);
or U17165 (N_17165,N_4826,N_9405);
xor U17166 (N_17166,N_7910,N_5614);
or U17167 (N_17167,N_8755,N_4987);
nand U17168 (N_17168,N_9163,N_4208);
nor U17169 (N_17169,N_4570,N_5955);
xor U17170 (N_17170,N_5035,N_6908);
xor U17171 (N_17171,N_5883,N_3058);
xor U17172 (N_17172,N_4151,N_8325);
nand U17173 (N_17173,N_8848,N_9595);
xor U17174 (N_17174,N_7179,N_1642);
and U17175 (N_17175,N_8660,N_7493);
xnor U17176 (N_17176,N_2020,N_3833);
nor U17177 (N_17177,N_7753,N_4655);
xnor U17178 (N_17178,N_924,N_455);
nand U17179 (N_17179,N_4532,N_5796);
nor U17180 (N_17180,N_692,N_1391);
nor U17181 (N_17181,N_5902,N_608);
nand U17182 (N_17182,N_5345,N_6335);
nor U17183 (N_17183,N_1478,N_8987);
nor U17184 (N_17184,N_6161,N_2836);
or U17185 (N_17185,N_1013,N_8726);
or U17186 (N_17186,N_8166,N_5504);
xor U17187 (N_17187,N_9218,N_9150);
nor U17188 (N_17188,N_6063,N_1768);
nand U17189 (N_17189,N_540,N_8004);
or U17190 (N_17190,N_607,N_6864);
nand U17191 (N_17191,N_551,N_5325);
xnor U17192 (N_17192,N_8950,N_7403);
or U17193 (N_17193,N_7430,N_5061);
and U17194 (N_17194,N_8599,N_1979);
and U17195 (N_17195,N_3910,N_2927);
xor U17196 (N_17196,N_9741,N_3961);
xnor U17197 (N_17197,N_8004,N_2892);
nand U17198 (N_17198,N_8199,N_6257);
or U17199 (N_17199,N_5615,N_6491);
nand U17200 (N_17200,N_6878,N_5843);
nand U17201 (N_17201,N_9828,N_2387);
nor U17202 (N_17202,N_1934,N_7108);
and U17203 (N_17203,N_7487,N_4936);
nand U17204 (N_17204,N_4546,N_3456);
nor U17205 (N_17205,N_9338,N_7691);
nand U17206 (N_17206,N_7451,N_6581);
nor U17207 (N_17207,N_9875,N_6879);
xor U17208 (N_17208,N_2826,N_1815);
xor U17209 (N_17209,N_4326,N_9977);
nand U17210 (N_17210,N_9071,N_6044);
nor U17211 (N_17211,N_3618,N_6594);
nor U17212 (N_17212,N_2114,N_6319);
xnor U17213 (N_17213,N_9762,N_4245);
and U17214 (N_17214,N_5302,N_6704);
xnor U17215 (N_17215,N_728,N_8096);
and U17216 (N_17216,N_9714,N_885);
nor U17217 (N_17217,N_3261,N_7843);
and U17218 (N_17218,N_1411,N_9588);
nor U17219 (N_17219,N_3949,N_1424);
xnor U17220 (N_17220,N_7413,N_309);
and U17221 (N_17221,N_4430,N_5574);
or U17222 (N_17222,N_6207,N_79);
xor U17223 (N_17223,N_4538,N_2063);
or U17224 (N_17224,N_4719,N_1760);
nand U17225 (N_17225,N_6037,N_4898);
xnor U17226 (N_17226,N_2091,N_9467);
xor U17227 (N_17227,N_7926,N_677);
nor U17228 (N_17228,N_6841,N_8492);
xor U17229 (N_17229,N_8480,N_2092);
nand U17230 (N_17230,N_1192,N_2428);
nor U17231 (N_17231,N_4037,N_6029);
nand U17232 (N_17232,N_7001,N_4994);
nor U17233 (N_17233,N_6004,N_4346);
nand U17234 (N_17234,N_6912,N_6877);
xor U17235 (N_17235,N_2637,N_6761);
xor U17236 (N_17236,N_55,N_930);
xor U17237 (N_17237,N_7017,N_2788);
and U17238 (N_17238,N_5525,N_9570);
nor U17239 (N_17239,N_1365,N_3317);
nand U17240 (N_17240,N_2753,N_100);
and U17241 (N_17241,N_3575,N_1836);
nand U17242 (N_17242,N_306,N_885);
and U17243 (N_17243,N_3332,N_968);
nand U17244 (N_17244,N_6379,N_986);
or U17245 (N_17245,N_5514,N_4073);
nand U17246 (N_17246,N_7765,N_6779);
nor U17247 (N_17247,N_6203,N_3320);
nand U17248 (N_17248,N_7629,N_3928);
nor U17249 (N_17249,N_3668,N_7754);
xnor U17250 (N_17250,N_1778,N_7977);
nand U17251 (N_17251,N_5760,N_5946);
and U17252 (N_17252,N_5302,N_7048);
and U17253 (N_17253,N_3787,N_6470);
xnor U17254 (N_17254,N_2817,N_5355);
nand U17255 (N_17255,N_5925,N_4179);
and U17256 (N_17256,N_9665,N_5281);
or U17257 (N_17257,N_7466,N_2576);
or U17258 (N_17258,N_8539,N_4726);
xor U17259 (N_17259,N_5022,N_2047);
nand U17260 (N_17260,N_3298,N_8685);
xor U17261 (N_17261,N_6442,N_6145);
or U17262 (N_17262,N_1963,N_5382);
nand U17263 (N_17263,N_9290,N_2137);
xor U17264 (N_17264,N_8035,N_4597);
nor U17265 (N_17265,N_2137,N_6984);
nor U17266 (N_17266,N_6696,N_3862);
or U17267 (N_17267,N_3691,N_3072);
and U17268 (N_17268,N_1456,N_4131);
nand U17269 (N_17269,N_1529,N_2303);
or U17270 (N_17270,N_2931,N_8015);
or U17271 (N_17271,N_1838,N_8311);
nor U17272 (N_17272,N_1704,N_7316);
or U17273 (N_17273,N_3478,N_3156);
or U17274 (N_17274,N_9885,N_3408);
nand U17275 (N_17275,N_1444,N_4983);
nand U17276 (N_17276,N_821,N_7177);
or U17277 (N_17277,N_2324,N_6059);
or U17278 (N_17278,N_4888,N_5248);
nand U17279 (N_17279,N_8530,N_1426);
nor U17280 (N_17280,N_8683,N_5620);
nor U17281 (N_17281,N_3107,N_938);
nand U17282 (N_17282,N_48,N_2116);
nor U17283 (N_17283,N_3837,N_2065);
and U17284 (N_17284,N_3126,N_2770);
xnor U17285 (N_17285,N_1452,N_639);
nand U17286 (N_17286,N_5,N_4571);
nor U17287 (N_17287,N_3383,N_7251);
xnor U17288 (N_17288,N_5836,N_8508);
xnor U17289 (N_17289,N_8056,N_9256);
nand U17290 (N_17290,N_2639,N_6216);
or U17291 (N_17291,N_718,N_4706);
or U17292 (N_17292,N_9020,N_4544);
nand U17293 (N_17293,N_2140,N_1074);
nor U17294 (N_17294,N_1615,N_3450);
xor U17295 (N_17295,N_6722,N_5280);
xnor U17296 (N_17296,N_9664,N_1236);
xnor U17297 (N_17297,N_6336,N_1554);
or U17298 (N_17298,N_3126,N_5638);
xor U17299 (N_17299,N_4792,N_5201);
nor U17300 (N_17300,N_4041,N_9873);
nand U17301 (N_17301,N_455,N_5358);
nand U17302 (N_17302,N_3512,N_9329);
xnor U17303 (N_17303,N_1402,N_565);
or U17304 (N_17304,N_9991,N_7910);
or U17305 (N_17305,N_9795,N_8194);
and U17306 (N_17306,N_2804,N_6118);
nor U17307 (N_17307,N_7095,N_1754);
and U17308 (N_17308,N_9689,N_4569);
nand U17309 (N_17309,N_2187,N_8319);
xor U17310 (N_17310,N_2518,N_2086);
and U17311 (N_17311,N_3148,N_1988);
or U17312 (N_17312,N_8112,N_4889);
nand U17313 (N_17313,N_6376,N_3434);
nor U17314 (N_17314,N_1694,N_4690);
nand U17315 (N_17315,N_786,N_9904);
or U17316 (N_17316,N_6722,N_7875);
and U17317 (N_17317,N_2380,N_2047);
xnor U17318 (N_17318,N_9857,N_1538);
and U17319 (N_17319,N_7928,N_5647);
and U17320 (N_17320,N_7384,N_6137);
and U17321 (N_17321,N_9483,N_1215);
nor U17322 (N_17322,N_2211,N_5702);
or U17323 (N_17323,N_9391,N_3478);
nand U17324 (N_17324,N_9261,N_9804);
and U17325 (N_17325,N_8686,N_6171);
or U17326 (N_17326,N_1864,N_418);
or U17327 (N_17327,N_6868,N_3086);
nand U17328 (N_17328,N_5181,N_5286);
nand U17329 (N_17329,N_2501,N_7461);
and U17330 (N_17330,N_6715,N_4614);
nor U17331 (N_17331,N_1379,N_2274);
or U17332 (N_17332,N_9660,N_8529);
nor U17333 (N_17333,N_5629,N_3571);
xor U17334 (N_17334,N_4476,N_37);
and U17335 (N_17335,N_1164,N_5908);
and U17336 (N_17336,N_2852,N_1142);
nor U17337 (N_17337,N_7493,N_4562);
and U17338 (N_17338,N_74,N_2941);
nand U17339 (N_17339,N_4928,N_1609);
nor U17340 (N_17340,N_7805,N_8114);
nand U17341 (N_17341,N_6414,N_5171);
xnor U17342 (N_17342,N_3915,N_5098);
nor U17343 (N_17343,N_1389,N_8179);
and U17344 (N_17344,N_42,N_9905);
or U17345 (N_17345,N_788,N_659);
nor U17346 (N_17346,N_6018,N_1178);
nor U17347 (N_17347,N_970,N_5764);
xor U17348 (N_17348,N_508,N_3184);
nand U17349 (N_17349,N_2096,N_1644);
nand U17350 (N_17350,N_8864,N_7977);
xor U17351 (N_17351,N_1487,N_8734);
xor U17352 (N_17352,N_5799,N_2715);
nand U17353 (N_17353,N_2326,N_7454);
xor U17354 (N_17354,N_3958,N_5934);
nand U17355 (N_17355,N_3922,N_5794);
xor U17356 (N_17356,N_1958,N_6840);
or U17357 (N_17357,N_1456,N_2019);
and U17358 (N_17358,N_301,N_5495);
or U17359 (N_17359,N_1087,N_6855);
xor U17360 (N_17360,N_4812,N_604);
or U17361 (N_17361,N_7849,N_9856);
xnor U17362 (N_17362,N_6872,N_6875);
nor U17363 (N_17363,N_1153,N_7310);
nand U17364 (N_17364,N_7605,N_1530);
xnor U17365 (N_17365,N_6192,N_5843);
xnor U17366 (N_17366,N_1086,N_8721);
nor U17367 (N_17367,N_555,N_5524);
or U17368 (N_17368,N_9804,N_749);
xor U17369 (N_17369,N_1970,N_800);
nor U17370 (N_17370,N_9863,N_895);
or U17371 (N_17371,N_7219,N_308);
xnor U17372 (N_17372,N_385,N_9834);
nand U17373 (N_17373,N_8888,N_7479);
nor U17374 (N_17374,N_1328,N_8183);
nor U17375 (N_17375,N_172,N_9388);
nand U17376 (N_17376,N_1107,N_9032);
and U17377 (N_17377,N_2754,N_3158);
nor U17378 (N_17378,N_9621,N_9671);
xor U17379 (N_17379,N_4156,N_517);
and U17380 (N_17380,N_3515,N_9303);
xnor U17381 (N_17381,N_2035,N_7541);
xor U17382 (N_17382,N_2308,N_216);
or U17383 (N_17383,N_3531,N_4841);
nor U17384 (N_17384,N_976,N_3574);
or U17385 (N_17385,N_9705,N_3954);
and U17386 (N_17386,N_1850,N_8285);
nor U17387 (N_17387,N_2941,N_740);
nor U17388 (N_17388,N_6545,N_9957);
or U17389 (N_17389,N_7411,N_1524);
and U17390 (N_17390,N_4306,N_3838);
nand U17391 (N_17391,N_6583,N_2584);
xor U17392 (N_17392,N_3372,N_442);
and U17393 (N_17393,N_4071,N_655);
or U17394 (N_17394,N_7133,N_2166);
nand U17395 (N_17395,N_5776,N_2322);
nand U17396 (N_17396,N_4423,N_7679);
xor U17397 (N_17397,N_8565,N_930);
and U17398 (N_17398,N_9039,N_5201);
nand U17399 (N_17399,N_3927,N_729);
and U17400 (N_17400,N_3659,N_9354);
or U17401 (N_17401,N_379,N_9850);
or U17402 (N_17402,N_2367,N_142);
xor U17403 (N_17403,N_1427,N_3026);
nor U17404 (N_17404,N_1415,N_8145);
xnor U17405 (N_17405,N_4997,N_3294);
or U17406 (N_17406,N_5172,N_6131);
nor U17407 (N_17407,N_7416,N_65);
nor U17408 (N_17408,N_6210,N_7917);
nor U17409 (N_17409,N_2492,N_3949);
and U17410 (N_17410,N_5157,N_7172);
nor U17411 (N_17411,N_8162,N_1782);
nand U17412 (N_17412,N_2223,N_2564);
or U17413 (N_17413,N_7798,N_1506);
and U17414 (N_17414,N_3593,N_7823);
and U17415 (N_17415,N_343,N_8933);
xnor U17416 (N_17416,N_2415,N_4350);
xor U17417 (N_17417,N_8657,N_188);
nand U17418 (N_17418,N_2468,N_5359);
and U17419 (N_17419,N_2626,N_8550);
and U17420 (N_17420,N_2234,N_5450);
and U17421 (N_17421,N_9456,N_2615);
and U17422 (N_17422,N_7636,N_7914);
nand U17423 (N_17423,N_138,N_355);
xor U17424 (N_17424,N_4881,N_299);
xnor U17425 (N_17425,N_5062,N_3311);
xnor U17426 (N_17426,N_6754,N_7382);
and U17427 (N_17427,N_2260,N_4007);
nor U17428 (N_17428,N_7156,N_7443);
and U17429 (N_17429,N_6417,N_1692);
nor U17430 (N_17430,N_6109,N_8397);
xor U17431 (N_17431,N_819,N_6440);
nand U17432 (N_17432,N_4221,N_8399);
xor U17433 (N_17433,N_6891,N_2188);
and U17434 (N_17434,N_8319,N_6561);
nand U17435 (N_17435,N_7467,N_733);
or U17436 (N_17436,N_5992,N_2128);
xor U17437 (N_17437,N_16,N_6014);
and U17438 (N_17438,N_4824,N_5552);
and U17439 (N_17439,N_4980,N_1825);
nor U17440 (N_17440,N_2599,N_5861);
nand U17441 (N_17441,N_1288,N_739);
nor U17442 (N_17442,N_7482,N_5707);
nand U17443 (N_17443,N_6615,N_8834);
or U17444 (N_17444,N_9213,N_5135);
nand U17445 (N_17445,N_7785,N_9049);
or U17446 (N_17446,N_3194,N_5226);
and U17447 (N_17447,N_6276,N_5913);
xnor U17448 (N_17448,N_4060,N_5636);
nor U17449 (N_17449,N_59,N_4881);
or U17450 (N_17450,N_4833,N_1999);
nor U17451 (N_17451,N_4733,N_1496);
nor U17452 (N_17452,N_2994,N_8952);
and U17453 (N_17453,N_3037,N_6925);
nor U17454 (N_17454,N_6622,N_2188);
and U17455 (N_17455,N_374,N_7654);
xor U17456 (N_17456,N_2957,N_1788);
nor U17457 (N_17457,N_5154,N_6332);
xnor U17458 (N_17458,N_4910,N_7256);
xnor U17459 (N_17459,N_2513,N_5851);
nand U17460 (N_17460,N_9983,N_8900);
nand U17461 (N_17461,N_6268,N_9706);
or U17462 (N_17462,N_3410,N_5537);
nand U17463 (N_17463,N_4076,N_1935);
and U17464 (N_17464,N_3207,N_7708);
and U17465 (N_17465,N_8137,N_7553);
nand U17466 (N_17466,N_9917,N_4474);
and U17467 (N_17467,N_7066,N_387);
nor U17468 (N_17468,N_2635,N_7416);
and U17469 (N_17469,N_5730,N_4994);
and U17470 (N_17470,N_6638,N_433);
and U17471 (N_17471,N_8034,N_8447);
or U17472 (N_17472,N_8925,N_8201);
and U17473 (N_17473,N_7466,N_4949);
nor U17474 (N_17474,N_3068,N_7316);
nand U17475 (N_17475,N_7698,N_114);
or U17476 (N_17476,N_813,N_2312);
nand U17477 (N_17477,N_3742,N_8978);
nor U17478 (N_17478,N_2962,N_9197);
xnor U17479 (N_17479,N_1610,N_8615);
nor U17480 (N_17480,N_7184,N_1158);
xor U17481 (N_17481,N_1210,N_4849);
or U17482 (N_17482,N_8231,N_6816);
nor U17483 (N_17483,N_8343,N_5911);
and U17484 (N_17484,N_7448,N_8481);
nor U17485 (N_17485,N_2192,N_4087);
nor U17486 (N_17486,N_3751,N_3413);
nand U17487 (N_17487,N_4145,N_9365);
xnor U17488 (N_17488,N_3198,N_1909);
nor U17489 (N_17489,N_3204,N_6979);
xnor U17490 (N_17490,N_7551,N_9709);
nor U17491 (N_17491,N_523,N_1758);
xnor U17492 (N_17492,N_8117,N_91);
nor U17493 (N_17493,N_6255,N_8553);
nand U17494 (N_17494,N_5303,N_6141);
and U17495 (N_17495,N_7813,N_7540);
and U17496 (N_17496,N_2618,N_5175);
or U17497 (N_17497,N_147,N_755);
and U17498 (N_17498,N_6220,N_4355);
or U17499 (N_17499,N_9788,N_3292);
nand U17500 (N_17500,N_6703,N_8501);
or U17501 (N_17501,N_3086,N_85);
nor U17502 (N_17502,N_8952,N_2511);
nand U17503 (N_17503,N_1756,N_68);
nor U17504 (N_17504,N_4589,N_1195);
and U17505 (N_17505,N_8079,N_7155);
and U17506 (N_17506,N_7708,N_1435);
nand U17507 (N_17507,N_3887,N_383);
and U17508 (N_17508,N_3494,N_3349);
xnor U17509 (N_17509,N_2550,N_1823);
xor U17510 (N_17510,N_5050,N_5633);
nor U17511 (N_17511,N_1480,N_1226);
nand U17512 (N_17512,N_1669,N_5185);
nand U17513 (N_17513,N_4323,N_1977);
nand U17514 (N_17514,N_377,N_8881);
nor U17515 (N_17515,N_3670,N_3463);
nor U17516 (N_17516,N_2278,N_7679);
xor U17517 (N_17517,N_9915,N_3474);
and U17518 (N_17518,N_6613,N_4656);
nand U17519 (N_17519,N_8098,N_4804);
or U17520 (N_17520,N_5588,N_3347);
nand U17521 (N_17521,N_9858,N_5493);
xor U17522 (N_17522,N_5562,N_9888);
and U17523 (N_17523,N_5832,N_988);
xnor U17524 (N_17524,N_5526,N_330);
and U17525 (N_17525,N_7855,N_4653);
xnor U17526 (N_17526,N_3,N_3728);
nor U17527 (N_17527,N_750,N_2457);
or U17528 (N_17528,N_1621,N_3541);
nand U17529 (N_17529,N_8482,N_6394);
and U17530 (N_17530,N_8796,N_301);
nand U17531 (N_17531,N_4271,N_5668);
xnor U17532 (N_17532,N_6255,N_4419);
or U17533 (N_17533,N_7053,N_5419);
xor U17534 (N_17534,N_4268,N_6125);
and U17535 (N_17535,N_8955,N_1175);
or U17536 (N_17536,N_6100,N_7589);
xor U17537 (N_17537,N_2800,N_286);
xor U17538 (N_17538,N_6326,N_4274);
or U17539 (N_17539,N_5005,N_3695);
or U17540 (N_17540,N_8056,N_7712);
and U17541 (N_17541,N_8499,N_6217);
or U17542 (N_17542,N_2764,N_8614);
xor U17543 (N_17543,N_143,N_8809);
xnor U17544 (N_17544,N_9710,N_5420);
or U17545 (N_17545,N_6577,N_3768);
or U17546 (N_17546,N_9688,N_994);
nor U17547 (N_17547,N_6925,N_5043);
and U17548 (N_17548,N_4767,N_9949);
or U17549 (N_17549,N_2314,N_3561);
nor U17550 (N_17550,N_971,N_8998);
or U17551 (N_17551,N_5511,N_2585);
xnor U17552 (N_17552,N_3236,N_3093);
and U17553 (N_17553,N_3192,N_9989);
nand U17554 (N_17554,N_8877,N_6690);
nand U17555 (N_17555,N_3450,N_6436);
xor U17556 (N_17556,N_770,N_728);
or U17557 (N_17557,N_2576,N_4867);
nand U17558 (N_17558,N_946,N_9723);
xor U17559 (N_17559,N_4174,N_2983);
and U17560 (N_17560,N_1638,N_6518);
or U17561 (N_17561,N_594,N_4729);
nand U17562 (N_17562,N_7179,N_9310);
and U17563 (N_17563,N_3734,N_3879);
or U17564 (N_17564,N_7184,N_3154);
nor U17565 (N_17565,N_2722,N_2902);
xnor U17566 (N_17566,N_9581,N_644);
xnor U17567 (N_17567,N_2214,N_9090);
or U17568 (N_17568,N_3363,N_9648);
nand U17569 (N_17569,N_2732,N_8858);
xnor U17570 (N_17570,N_3288,N_5813);
and U17571 (N_17571,N_7516,N_4338);
and U17572 (N_17572,N_1623,N_7622);
nor U17573 (N_17573,N_8356,N_7237);
nor U17574 (N_17574,N_9904,N_9784);
or U17575 (N_17575,N_534,N_6550);
nor U17576 (N_17576,N_1404,N_8589);
and U17577 (N_17577,N_2176,N_1919);
xor U17578 (N_17578,N_9797,N_1720);
nor U17579 (N_17579,N_5116,N_8180);
nand U17580 (N_17580,N_901,N_8600);
nor U17581 (N_17581,N_5619,N_9819);
or U17582 (N_17582,N_3346,N_2434);
nor U17583 (N_17583,N_5138,N_195);
nor U17584 (N_17584,N_5633,N_4651);
nand U17585 (N_17585,N_4632,N_6091);
nor U17586 (N_17586,N_9298,N_6157);
nor U17587 (N_17587,N_8391,N_4972);
xor U17588 (N_17588,N_6035,N_605);
xor U17589 (N_17589,N_6215,N_5241);
nand U17590 (N_17590,N_9443,N_8460);
or U17591 (N_17591,N_2429,N_1638);
xnor U17592 (N_17592,N_6580,N_3481);
and U17593 (N_17593,N_7477,N_9944);
nand U17594 (N_17594,N_7740,N_7585);
nand U17595 (N_17595,N_4585,N_4727);
or U17596 (N_17596,N_4637,N_9890);
xnor U17597 (N_17597,N_7167,N_6184);
nor U17598 (N_17598,N_8656,N_7142);
xnor U17599 (N_17599,N_6615,N_8159);
or U17600 (N_17600,N_3597,N_3851);
nand U17601 (N_17601,N_1056,N_8273);
and U17602 (N_17602,N_3694,N_8976);
nand U17603 (N_17603,N_8139,N_4833);
nand U17604 (N_17604,N_9745,N_9270);
and U17605 (N_17605,N_4903,N_532);
nor U17606 (N_17606,N_6597,N_9836);
and U17607 (N_17607,N_4085,N_5716);
nor U17608 (N_17608,N_6868,N_6599);
xor U17609 (N_17609,N_9549,N_9862);
nor U17610 (N_17610,N_7136,N_4642);
nor U17611 (N_17611,N_6278,N_7630);
or U17612 (N_17612,N_9488,N_8050);
nor U17613 (N_17613,N_1481,N_336);
or U17614 (N_17614,N_29,N_3017);
nand U17615 (N_17615,N_3551,N_9196);
nand U17616 (N_17616,N_4255,N_4437);
nor U17617 (N_17617,N_8932,N_557);
xor U17618 (N_17618,N_1417,N_9258);
nand U17619 (N_17619,N_8849,N_8376);
or U17620 (N_17620,N_9257,N_9864);
and U17621 (N_17621,N_2715,N_8036);
xor U17622 (N_17622,N_1695,N_8883);
nor U17623 (N_17623,N_8970,N_6353);
or U17624 (N_17624,N_3103,N_6705);
and U17625 (N_17625,N_110,N_2734);
nor U17626 (N_17626,N_1005,N_7906);
and U17627 (N_17627,N_328,N_9567);
or U17628 (N_17628,N_2197,N_4135);
nor U17629 (N_17629,N_5516,N_2034);
nand U17630 (N_17630,N_3839,N_3456);
or U17631 (N_17631,N_2971,N_8645);
and U17632 (N_17632,N_8116,N_7887);
and U17633 (N_17633,N_9208,N_7110);
xor U17634 (N_17634,N_2596,N_3684);
or U17635 (N_17635,N_3806,N_7105);
or U17636 (N_17636,N_9256,N_4198);
xor U17637 (N_17637,N_8688,N_7876);
or U17638 (N_17638,N_6558,N_4061);
nor U17639 (N_17639,N_9362,N_3772);
and U17640 (N_17640,N_1378,N_3402);
and U17641 (N_17641,N_8854,N_7338);
xor U17642 (N_17642,N_6708,N_36);
xnor U17643 (N_17643,N_5546,N_629);
nand U17644 (N_17644,N_9805,N_880);
and U17645 (N_17645,N_6370,N_8575);
or U17646 (N_17646,N_7953,N_1079);
or U17647 (N_17647,N_8229,N_7339);
nand U17648 (N_17648,N_4663,N_5402);
nor U17649 (N_17649,N_9046,N_6827);
xnor U17650 (N_17650,N_7633,N_7130);
nor U17651 (N_17651,N_3786,N_5056);
nand U17652 (N_17652,N_3517,N_1807);
nor U17653 (N_17653,N_2259,N_6361);
nor U17654 (N_17654,N_5864,N_6036);
nand U17655 (N_17655,N_8290,N_5477);
xor U17656 (N_17656,N_1023,N_5289);
nand U17657 (N_17657,N_7583,N_3262);
and U17658 (N_17658,N_754,N_7722);
or U17659 (N_17659,N_8702,N_1652);
xnor U17660 (N_17660,N_2730,N_9037);
nor U17661 (N_17661,N_2803,N_4382);
or U17662 (N_17662,N_9798,N_7094);
nand U17663 (N_17663,N_2172,N_661);
nor U17664 (N_17664,N_2329,N_1656);
nand U17665 (N_17665,N_1481,N_2769);
xor U17666 (N_17666,N_8665,N_4226);
nor U17667 (N_17667,N_7362,N_1927);
nand U17668 (N_17668,N_7076,N_7960);
xnor U17669 (N_17669,N_5412,N_7329);
or U17670 (N_17670,N_7676,N_2931);
nor U17671 (N_17671,N_464,N_7031);
nor U17672 (N_17672,N_6100,N_429);
nor U17673 (N_17673,N_5881,N_9381);
xnor U17674 (N_17674,N_1337,N_8577);
nor U17675 (N_17675,N_4384,N_8681);
nor U17676 (N_17676,N_8081,N_9999);
xnor U17677 (N_17677,N_1397,N_9508);
or U17678 (N_17678,N_9043,N_4337);
nand U17679 (N_17679,N_7872,N_5031);
and U17680 (N_17680,N_7693,N_9695);
nor U17681 (N_17681,N_4678,N_295);
xor U17682 (N_17682,N_3988,N_3341);
nand U17683 (N_17683,N_1407,N_3380);
and U17684 (N_17684,N_3306,N_2368);
and U17685 (N_17685,N_46,N_9409);
nand U17686 (N_17686,N_6145,N_913);
or U17687 (N_17687,N_191,N_8683);
or U17688 (N_17688,N_6855,N_7261);
and U17689 (N_17689,N_4836,N_704);
and U17690 (N_17690,N_3665,N_3150);
xor U17691 (N_17691,N_6220,N_8684);
xor U17692 (N_17692,N_4208,N_2943);
nand U17693 (N_17693,N_7036,N_1121);
or U17694 (N_17694,N_901,N_7128);
nor U17695 (N_17695,N_6775,N_5564);
nand U17696 (N_17696,N_6845,N_6986);
nor U17697 (N_17697,N_8708,N_945);
nor U17698 (N_17698,N_4742,N_164);
xnor U17699 (N_17699,N_390,N_3981);
xnor U17700 (N_17700,N_6497,N_6718);
and U17701 (N_17701,N_7285,N_8466);
or U17702 (N_17702,N_8630,N_9036);
or U17703 (N_17703,N_9430,N_4359);
xor U17704 (N_17704,N_5016,N_7806);
nor U17705 (N_17705,N_409,N_8580);
and U17706 (N_17706,N_2527,N_3107);
and U17707 (N_17707,N_9438,N_9234);
xnor U17708 (N_17708,N_6771,N_7421);
xor U17709 (N_17709,N_9646,N_6805);
nor U17710 (N_17710,N_4474,N_4630);
xor U17711 (N_17711,N_5580,N_9065);
nor U17712 (N_17712,N_8652,N_3335);
or U17713 (N_17713,N_3052,N_2585);
and U17714 (N_17714,N_6739,N_7489);
nor U17715 (N_17715,N_4779,N_2394);
xnor U17716 (N_17716,N_5026,N_5876);
xor U17717 (N_17717,N_1809,N_2405);
or U17718 (N_17718,N_3558,N_7681);
nand U17719 (N_17719,N_3382,N_4607);
nand U17720 (N_17720,N_2767,N_6227);
and U17721 (N_17721,N_8222,N_2609);
or U17722 (N_17722,N_1443,N_1449);
xnor U17723 (N_17723,N_968,N_9468);
nor U17724 (N_17724,N_7956,N_4844);
and U17725 (N_17725,N_5453,N_3942);
and U17726 (N_17726,N_8156,N_9387);
xor U17727 (N_17727,N_347,N_1459);
and U17728 (N_17728,N_3396,N_1879);
or U17729 (N_17729,N_3128,N_7360);
xnor U17730 (N_17730,N_2791,N_6929);
or U17731 (N_17731,N_8982,N_7394);
nand U17732 (N_17732,N_3895,N_473);
nor U17733 (N_17733,N_3651,N_1294);
or U17734 (N_17734,N_9708,N_2662);
xor U17735 (N_17735,N_1954,N_778);
xor U17736 (N_17736,N_4004,N_8965);
nor U17737 (N_17737,N_4527,N_9249);
nor U17738 (N_17738,N_884,N_5748);
nand U17739 (N_17739,N_1963,N_8072);
nor U17740 (N_17740,N_8596,N_6948);
and U17741 (N_17741,N_5539,N_1242);
nor U17742 (N_17742,N_6212,N_4925);
or U17743 (N_17743,N_1997,N_4772);
and U17744 (N_17744,N_7357,N_863);
or U17745 (N_17745,N_7182,N_558);
xnor U17746 (N_17746,N_1059,N_2601);
and U17747 (N_17747,N_899,N_8884);
nand U17748 (N_17748,N_3057,N_1542);
xnor U17749 (N_17749,N_1280,N_2243);
nor U17750 (N_17750,N_9182,N_9508);
nand U17751 (N_17751,N_3730,N_4826);
and U17752 (N_17752,N_2995,N_5915);
and U17753 (N_17753,N_4506,N_1640);
xor U17754 (N_17754,N_129,N_4003);
or U17755 (N_17755,N_7034,N_5097);
xor U17756 (N_17756,N_3761,N_1243);
or U17757 (N_17757,N_6895,N_3745);
or U17758 (N_17758,N_8425,N_1368);
nor U17759 (N_17759,N_6569,N_7857);
xnor U17760 (N_17760,N_7508,N_5507);
nand U17761 (N_17761,N_8345,N_2214);
nand U17762 (N_17762,N_399,N_7612);
or U17763 (N_17763,N_9606,N_874);
nor U17764 (N_17764,N_82,N_363);
xor U17765 (N_17765,N_1396,N_6736);
and U17766 (N_17766,N_8567,N_6935);
nor U17767 (N_17767,N_6022,N_3684);
nor U17768 (N_17768,N_7221,N_1443);
and U17769 (N_17769,N_2786,N_8522);
or U17770 (N_17770,N_1391,N_2899);
nor U17771 (N_17771,N_6335,N_2939);
or U17772 (N_17772,N_8695,N_7337);
or U17773 (N_17773,N_8642,N_8119);
or U17774 (N_17774,N_6560,N_5052);
nand U17775 (N_17775,N_1394,N_8461);
and U17776 (N_17776,N_2578,N_8259);
nor U17777 (N_17777,N_9299,N_7498);
and U17778 (N_17778,N_6518,N_5461);
xnor U17779 (N_17779,N_190,N_8189);
or U17780 (N_17780,N_3992,N_1116);
nor U17781 (N_17781,N_6554,N_5508);
nor U17782 (N_17782,N_1730,N_3039);
nor U17783 (N_17783,N_3037,N_9727);
or U17784 (N_17784,N_7188,N_6811);
and U17785 (N_17785,N_5330,N_601);
nand U17786 (N_17786,N_4602,N_8437);
and U17787 (N_17787,N_699,N_5489);
nor U17788 (N_17788,N_198,N_6142);
nand U17789 (N_17789,N_4839,N_9061);
and U17790 (N_17790,N_8870,N_1218);
nor U17791 (N_17791,N_8956,N_7960);
xor U17792 (N_17792,N_2123,N_9613);
or U17793 (N_17793,N_3223,N_8023);
xnor U17794 (N_17794,N_4341,N_5910);
xor U17795 (N_17795,N_1240,N_713);
and U17796 (N_17796,N_6548,N_808);
and U17797 (N_17797,N_2417,N_8948);
xnor U17798 (N_17798,N_7226,N_9390);
xor U17799 (N_17799,N_4593,N_2244);
or U17800 (N_17800,N_633,N_8965);
nand U17801 (N_17801,N_7211,N_8952);
nor U17802 (N_17802,N_2289,N_6931);
xnor U17803 (N_17803,N_4981,N_4881);
nand U17804 (N_17804,N_8553,N_7577);
and U17805 (N_17805,N_9735,N_11);
nor U17806 (N_17806,N_249,N_2037);
and U17807 (N_17807,N_2976,N_3280);
nand U17808 (N_17808,N_7436,N_371);
xnor U17809 (N_17809,N_2705,N_7308);
nand U17810 (N_17810,N_8621,N_3054);
nor U17811 (N_17811,N_6752,N_1411);
nor U17812 (N_17812,N_7602,N_6717);
and U17813 (N_17813,N_1775,N_6731);
nor U17814 (N_17814,N_3095,N_6642);
nor U17815 (N_17815,N_8854,N_6247);
nand U17816 (N_17816,N_4470,N_5830);
nand U17817 (N_17817,N_4422,N_5744);
xor U17818 (N_17818,N_7521,N_4072);
and U17819 (N_17819,N_6016,N_1966);
nand U17820 (N_17820,N_4514,N_6443);
nand U17821 (N_17821,N_5709,N_4076);
nand U17822 (N_17822,N_1809,N_9543);
and U17823 (N_17823,N_4116,N_9442);
or U17824 (N_17824,N_1284,N_6512);
and U17825 (N_17825,N_1789,N_2677);
xnor U17826 (N_17826,N_9957,N_1322);
nand U17827 (N_17827,N_5311,N_158);
xor U17828 (N_17828,N_934,N_287);
xnor U17829 (N_17829,N_6861,N_4258);
or U17830 (N_17830,N_4530,N_5123);
and U17831 (N_17831,N_1871,N_1379);
and U17832 (N_17832,N_3714,N_8642);
nor U17833 (N_17833,N_4671,N_8063);
nor U17834 (N_17834,N_7170,N_6901);
and U17835 (N_17835,N_2421,N_6172);
and U17836 (N_17836,N_9514,N_769);
xor U17837 (N_17837,N_7993,N_4371);
and U17838 (N_17838,N_4417,N_1610);
and U17839 (N_17839,N_7221,N_1021);
or U17840 (N_17840,N_1363,N_4302);
nand U17841 (N_17841,N_3766,N_9953);
and U17842 (N_17842,N_2348,N_2135);
or U17843 (N_17843,N_1952,N_1417);
xor U17844 (N_17844,N_6847,N_3801);
xor U17845 (N_17845,N_6405,N_2775);
xnor U17846 (N_17846,N_6865,N_6429);
xnor U17847 (N_17847,N_3311,N_4593);
nor U17848 (N_17848,N_9294,N_5717);
or U17849 (N_17849,N_7564,N_1623);
or U17850 (N_17850,N_2160,N_7206);
nand U17851 (N_17851,N_4343,N_3848);
xnor U17852 (N_17852,N_5604,N_1876);
nor U17853 (N_17853,N_5474,N_3739);
and U17854 (N_17854,N_4270,N_6962);
and U17855 (N_17855,N_3966,N_3803);
nand U17856 (N_17856,N_5146,N_2309);
xor U17857 (N_17857,N_7407,N_1861);
xnor U17858 (N_17858,N_1193,N_894);
and U17859 (N_17859,N_1468,N_2404);
or U17860 (N_17860,N_9916,N_1759);
nor U17861 (N_17861,N_4302,N_3576);
and U17862 (N_17862,N_6677,N_5534);
xor U17863 (N_17863,N_9869,N_6924);
xor U17864 (N_17864,N_3273,N_3709);
nand U17865 (N_17865,N_1316,N_1427);
nor U17866 (N_17866,N_3797,N_5252);
xor U17867 (N_17867,N_2692,N_1951);
nand U17868 (N_17868,N_8368,N_5517);
and U17869 (N_17869,N_8770,N_645);
xnor U17870 (N_17870,N_2207,N_1821);
or U17871 (N_17871,N_9428,N_8905);
or U17872 (N_17872,N_9928,N_1665);
or U17873 (N_17873,N_1630,N_9040);
nand U17874 (N_17874,N_5302,N_5515);
and U17875 (N_17875,N_8799,N_9215);
xor U17876 (N_17876,N_8723,N_1499);
nand U17877 (N_17877,N_4375,N_3981);
or U17878 (N_17878,N_9076,N_9045);
or U17879 (N_17879,N_1573,N_2497);
nand U17880 (N_17880,N_837,N_726);
xor U17881 (N_17881,N_6026,N_5827);
nand U17882 (N_17882,N_6560,N_488);
or U17883 (N_17883,N_7234,N_6154);
nor U17884 (N_17884,N_954,N_1664);
nor U17885 (N_17885,N_4060,N_5067);
nor U17886 (N_17886,N_5272,N_4921);
and U17887 (N_17887,N_1704,N_6854);
nor U17888 (N_17888,N_7118,N_8282);
xor U17889 (N_17889,N_1936,N_4760);
nand U17890 (N_17890,N_6147,N_4955);
nand U17891 (N_17891,N_7478,N_2750);
xnor U17892 (N_17892,N_9093,N_5326);
or U17893 (N_17893,N_4180,N_4623);
xnor U17894 (N_17894,N_3620,N_9784);
nor U17895 (N_17895,N_5175,N_4072);
nand U17896 (N_17896,N_7494,N_2022);
nor U17897 (N_17897,N_6128,N_9862);
nor U17898 (N_17898,N_3185,N_8030);
nand U17899 (N_17899,N_5914,N_1657);
or U17900 (N_17900,N_7931,N_9483);
or U17901 (N_17901,N_6371,N_2331);
nor U17902 (N_17902,N_1817,N_5526);
and U17903 (N_17903,N_8354,N_4985);
nand U17904 (N_17904,N_2055,N_639);
nor U17905 (N_17905,N_7289,N_9180);
xnor U17906 (N_17906,N_6025,N_6183);
and U17907 (N_17907,N_5471,N_9295);
xnor U17908 (N_17908,N_1744,N_1812);
and U17909 (N_17909,N_2027,N_4338);
and U17910 (N_17910,N_7357,N_1224);
and U17911 (N_17911,N_8635,N_9717);
nor U17912 (N_17912,N_3513,N_2029);
nor U17913 (N_17913,N_2337,N_2940);
nand U17914 (N_17914,N_8806,N_2502);
or U17915 (N_17915,N_2016,N_3801);
nand U17916 (N_17916,N_5280,N_4882);
nand U17917 (N_17917,N_7057,N_5332);
nor U17918 (N_17918,N_8433,N_7839);
xor U17919 (N_17919,N_4939,N_606);
nor U17920 (N_17920,N_5973,N_1066);
and U17921 (N_17921,N_5708,N_5199);
and U17922 (N_17922,N_3496,N_1788);
xnor U17923 (N_17923,N_6899,N_9903);
or U17924 (N_17924,N_8435,N_217);
or U17925 (N_17925,N_1596,N_4402);
nand U17926 (N_17926,N_1780,N_7145);
nand U17927 (N_17927,N_1845,N_4480);
and U17928 (N_17928,N_1456,N_5095);
xor U17929 (N_17929,N_1929,N_3524);
or U17930 (N_17930,N_5617,N_1354);
or U17931 (N_17931,N_3385,N_1665);
nand U17932 (N_17932,N_2411,N_1419);
nand U17933 (N_17933,N_3468,N_7505);
or U17934 (N_17934,N_1062,N_7339);
or U17935 (N_17935,N_9697,N_3465);
or U17936 (N_17936,N_9199,N_5315);
nor U17937 (N_17937,N_6419,N_3627);
xor U17938 (N_17938,N_465,N_5392);
xnor U17939 (N_17939,N_9558,N_4846);
xnor U17940 (N_17940,N_5341,N_7306);
xor U17941 (N_17941,N_5022,N_6006);
nand U17942 (N_17942,N_7975,N_1980);
and U17943 (N_17943,N_3003,N_4697);
and U17944 (N_17944,N_4948,N_2966);
xnor U17945 (N_17945,N_7828,N_8461);
or U17946 (N_17946,N_5928,N_5185);
nand U17947 (N_17947,N_1101,N_1841);
nor U17948 (N_17948,N_849,N_5112);
and U17949 (N_17949,N_9332,N_9086);
nand U17950 (N_17950,N_8902,N_8756);
nor U17951 (N_17951,N_2037,N_8287);
nor U17952 (N_17952,N_8964,N_1684);
nor U17953 (N_17953,N_1247,N_9718);
or U17954 (N_17954,N_8673,N_1949);
nand U17955 (N_17955,N_1549,N_4236);
and U17956 (N_17956,N_985,N_4599);
nor U17957 (N_17957,N_817,N_3313);
xnor U17958 (N_17958,N_6401,N_1105);
or U17959 (N_17959,N_4864,N_6314);
nor U17960 (N_17960,N_4675,N_8600);
and U17961 (N_17961,N_5137,N_3834);
nand U17962 (N_17962,N_9083,N_6448);
nand U17963 (N_17963,N_3280,N_7718);
xor U17964 (N_17964,N_571,N_8966);
xor U17965 (N_17965,N_2208,N_7087);
xor U17966 (N_17966,N_4453,N_6498);
nor U17967 (N_17967,N_5851,N_7657);
xor U17968 (N_17968,N_9050,N_3041);
xor U17969 (N_17969,N_7145,N_8955);
and U17970 (N_17970,N_9607,N_6557);
or U17971 (N_17971,N_2051,N_916);
or U17972 (N_17972,N_1174,N_6213);
xnor U17973 (N_17973,N_2735,N_3783);
and U17974 (N_17974,N_3916,N_8060);
nor U17975 (N_17975,N_6064,N_478);
nand U17976 (N_17976,N_5301,N_9730);
nor U17977 (N_17977,N_623,N_5608);
nor U17978 (N_17978,N_6754,N_8244);
nand U17979 (N_17979,N_3148,N_975);
xnor U17980 (N_17980,N_6769,N_3165);
or U17981 (N_17981,N_598,N_3673);
xnor U17982 (N_17982,N_2063,N_3765);
xnor U17983 (N_17983,N_9235,N_2504);
or U17984 (N_17984,N_9108,N_5222);
nor U17985 (N_17985,N_9635,N_9216);
nand U17986 (N_17986,N_405,N_327);
and U17987 (N_17987,N_5060,N_6017);
or U17988 (N_17988,N_9938,N_1419);
xor U17989 (N_17989,N_1067,N_3502);
and U17990 (N_17990,N_5633,N_2488);
nand U17991 (N_17991,N_8485,N_9547);
nor U17992 (N_17992,N_5424,N_9419);
and U17993 (N_17993,N_8820,N_9999);
nand U17994 (N_17994,N_2792,N_8366);
and U17995 (N_17995,N_8612,N_7654);
or U17996 (N_17996,N_8995,N_4654);
xnor U17997 (N_17997,N_5681,N_7836);
and U17998 (N_17998,N_4350,N_683);
and U17999 (N_17999,N_7073,N_7219);
nor U18000 (N_18000,N_6870,N_3676);
or U18001 (N_18001,N_14,N_4209);
or U18002 (N_18002,N_4658,N_7172);
and U18003 (N_18003,N_4232,N_3348);
nor U18004 (N_18004,N_6397,N_8182);
xor U18005 (N_18005,N_8272,N_3712);
or U18006 (N_18006,N_9548,N_3730);
xnor U18007 (N_18007,N_2485,N_4843);
nand U18008 (N_18008,N_2522,N_173);
nor U18009 (N_18009,N_1716,N_4506);
or U18010 (N_18010,N_6810,N_8584);
nor U18011 (N_18011,N_9441,N_5063);
nor U18012 (N_18012,N_1502,N_4772);
or U18013 (N_18013,N_8943,N_207);
nor U18014 (N_18014,N_2228,N_8025);
xor U18015 (N_18015,N_7137,N_4555);
and U18016 (N_18016,N_5385,N_2425);
and U18017 (N_18017,N_550,N_2270);
nor U18018 (N_18018,N_3393,N_1607);
nand U18019 (N_18019,N_6495,N_5216);
nand U18020 (N_18020,N_3956,N_7193);
xnor U18021 (N_18021,N_1434,N_9740);
or U18022 (N_18022,N_4044,N_2416);
xnor U18023 (N_18023,N_2872,N_8680);
xnor U18024 (N_18024,N_8376,N_800);
and U18025 (N_18025,N_3343,N_4478);
xor U18026 (N_18026,N_359,N_7413);
nand U18027 (N_18027,N_2539,N_4660);
nand U18028 (N_18028,N_2114,N_3845);
xnor U18029 (N_18029,N_8681,N_1345);
or U18030 (N_18030,N_6334,N_6195);
nand U18031 (N_18031,N_4978,N_4969);
or U18032 (N_18032,N_6971,N_1815);
nor U18033 (N_18033,N_8274,N_9758);
and U18034 (N_18034,N_6736,N_5995);
or U18035 (N_18035,N_2883,N_7556);
or U18036 (N_18036,N_2800,N_9301);
xor U18037 (N_18037,N_5754,N_7634);
nand U18038 (N_18038,N_959,N_7090);
nor U18039 (N_18039,N_4483,N_8818);
nand U18040 (N_18040,N_5464,N_6932);
and U18041 (N_18041,N_4629,N_6190);
and U18042 (N_18042,N_4286,N_2311);
nand U18043 (N_18043,N_8725,N_2690);
nand U18044 (N_18044,N_4995,N_821);
and U18045 (N_18045,N_383,N_8057);
and U18046 (N_18046,N_2556,N_3781);
nor U18047 (N_18047,N_3321,N_9863);
xnor U18048 (N_18048,N_7033,N_1634);
nor U18049 (N_18049,N_2527,N_6641);
nor U18050 (N_18050,N_4557,N_6742);
xnor U18051 (N_18051,N_4368,N_6301);
nor U18052 (N_18052,N_7454,N_9326);
or U18053 (N_18053,N_4675,N_7061);
or U18054 (N_18054,N_4075,N_439);
nand U18055 (N_18055,N_5356,N_4212);
xnor U18056 (N_18056,N_4829,N_4793);
and U18057 (N_18057,N_6330,N_7483);
or U18058 (N_18058,N_5599,N_9393);
and U18059 (N_18059,N_2340,N_6520);
and U18060 (N_18060,N_4776,N_6541);
xor U18061 (N_18061,N_2465,N_6354);
nand U18062 (N_18062,N_887,N_7093);
or U18063 (N_18063,N_5479,N_9736);
or U18064 (N_18064,N_8749,N_2305);
nor U18065 (N_18065,N_7446,N_417);
xor U18066 (N_18066,N_4456,N_7654);
nor U18067 (N_18067,N_1108,N_8218);
and U18068 (N_18068,N_7397,N_1323);
nand U18069 (N_18069,N_811,N_7928);
or U18070 (N_18070,N_1473,N_7180);
nor U18071 (N_18071,N_692,N_7685);
xor U18072 (N_18072,N_6443,N_115);
and U18073 (N_18073,N_9146,N_9928);
or U18074 (N_18074,N_1317,N_8717);
xnor U18075 (N_18075,N_6904,N_199);
nand U18076 (N_18076,N_5824,N_5289);
xor U18077 (N_18077,N_2454,N_2891);
and U18078 (N_18078,N_2404,N_1679);
xnor U18079 (N_18079,N_9673,N_9007);
nand U18080 (N_18080,N_3911,N_9420);
nor U18081 (N_18081,N_9631,N_6078);
nand U18082 (N_18082,N_5675,N_573);
and U18083 (N_18083,N_7565,N_7551);
nor U18084 (N_18084,N_3448,N_3921);
nand U18085 (N_18085,N_6942,N_6722);
and U18086 (N_18086,N_3352,N_2813);
nor U18087 (N_18087,N_4235,N_4749);
xor U18088 (N_18088,N_2903,N_4596);
nor U18089 (N_18089,N_5148,N_8340);
nand U18090 (N_18090,N_9478,N_3238);
xor U18091 (N_18091,N_1934,N_6886);
nand U18092 (N_18092,N_3490,N_7362);
xnor U18093 (N_18093,N_8874,N_1290);
and U18094 (N_18094,N_7578,N_9955);
nor U18095 (N_18095,N_7564,N_8989);
nor U18096 (N_18096,N_8083,N_1232);
nand U18097 (N_18097,N_8024,N_656);
nand U18098 (N_18098,N_1444,N_5304);
xnor U18099 (N_18099,N_1644,N_2631);
xnor U18100 (N_18100,N_5528,N_2172);
xor U18101 (N_18101,N_9284,N_1044);
and U18102 (N_18102,N_7839,N_2679);
or U18103 (N_18103,N_6404,N_6824);
or U18104 (N_18104,N_4475,N_8898);
xor U18105 (N_18105,N_1195,N_6870);
xnor U18106 (N_18106,N_9823,N_8957);
nand U18107 (N_18107,N_2036,N_9634);
nand U18108 (N_18108,N_7592,N_4190);
or U18109 (N_18109,N_7387,N_7806);
nand U18110 (N_18110,N_439,N_9354);
nand U18111 (N_18111,N_3900,N_7321);
xnor U18112 (N_18112,N_3394,N_4330);
nor U18113 (N_18113,N_1464,N_3302);
or U18114 (N_18114,N_3,N_4032);
or U18115 (N_18115,N_6684,N_6038);
or U18116 (N_18116,N_1542,N_3517);
and U18117 (N_18117,N_2058,N_6752);
nand U18118 (N_18118,N_1875,N_6470);
and U18119 (N_18119,N_5765,N_3198);
xnor U18120 (N_18120,N_6703,N_6390);
nor U18121 (N_18121,N_764,N_3222);
and U18122 (N_18122,N_9919,N_3175);
or U18123 (N_18123,N_1605,N_9443);
xor U18124 (N_18124,N_6353,N_8723);
nand U18125 (N_18125,N_3660,N_6691);
and U18126 (N_18126,N_2521,N_6509);
or U18127 (N_18127,N_1792,N_4400);
nand U18128 (N_18128,N_8414,N_3272);
nor U18129 (N_18129,N_9041,N_6397);
xor U18130 (N_18130,N_1947,N_4454);
and U18131 (N_18131,N_491,N_8466);
or U18132 (N_18132,N_152,N_3906);
and U18133 (N_18133,N_2582,N_1263);
nand U18134 (N_18134,N_8341,N_220);
and U18135 (N_18135,N_9966,N_4321);
or U18136 (N_18136,N_6360,N_7150);
xnor U18137 (N_18137,N_3602,N_4042);
xor U18138 (N_18138,N_8135,N_8769);
nand U18139 (N_18139,N_1422,N_6653);
and U18140 (N_18140,N_6675,N_3870);
nor U18141 (N_18141,N_7700,N_9229);
nand U18142 (N_18142,N_199,N_2431);
nor U18143 (N_18143,N_5367,N_6214);
nor U18144 (N_18144,N_8150,N_9589);
or U18145 (N_18145,N_4968,N_7568);
or U18146 (N_18146,N_607,N_4993);
and U18147 (N_18147,N_9095,N_5602);
and U18148 (N_18148,N_8218,N_5422);
nand U18149 (N_18149,N_316,N_6498);
nor U18150 (N_18150,N_6222,N_6912);
nor U18151 (N_18151,N_886,N_7310);
nand U18152 (N_18152,N_371,N_6277);
and U18153 (N_18153,N_4112,N_4887);
or U18154 (N_18154,N_2701,N_6792);
or U18155 (N_18155,N_75,N_5804);
nor U18156 (N_18156,N_5708,N_5385);
xor U18157 (N_18157,N_6910,N_7891);
nor U18158 (N_18158,N_4579,N_5811);
nand U18159 (N_18159,N_2439,N_3166);
xnor U18160 (N_18160,N_1190,N_5685);
or U18161 (N_18161,N_3830,N_2316);
or U18162 (N_18162,N_4234,N_7062);
xnor U18163 (N_18163,N_6799,N_5617);
nand U18164 (N_18164,N_1474,N_7235);
nor U18165 (N_18165,N_3152,N_4282);
xnor U18166 (N_18166,N_4158,N_7684);
and U18167 (N_18167,N_6335,N_1554);
or U18168 (N_18168,N_1498,N_8458);
and U18169 (N_18169,N_7228,N_8550);
xnor U18170 (N_18170,N_4678,N_1150);
xor U18171 (N_18171,N_3396,N_9982);
nand U18172 (N_18172,N_8833,N_4794);
and U18173 (N_18173,N_1762,N_918);
or U18174 (N_18174,N_8431,N_459);
or U18175 (N_18175,N_7635,N_168);
nand U18176 (N_18176,N_4413,N_1810);
or U18177 (N_18177,N_907,N_435);
and U18178 (N_18178,N_6645,N_9835);
nor U18179 (N_18179,N_3502,N_7053);
or U18180 (N_18180,N_5617,N_9081);
or U18181 (N_18181,N_7840,N_4263);
nor U18182 (N_18182,N_5269,N_4618);
nand U18183 (N_18183,N_848,N_994);
nand U18184 (N_18184,N_9750,N_7243);
nor U18185 (N_18185,N_3506,N_4892);
or U18186 (N_18186,N_1730,N_1916);
and U18187 (N_18187,N_5584,N_7719);
xnor U18188 (N_18188,N_2450,N_5936);
nand U18189 (N_18189,N_3868,N_9778);
nor U18190 (N_18190,N_7151,N_9200);
nand U18191 (N_18191,N_6978,N_3352);
or U18192 (N_18192,N_5702,N_8022);
xnor U18193 (N_18193,N_7712,N_243);
or U18194 (N_18194,N_9395,N_5180);
xor U18195 (N_18195,N_7799,N_8484);
and U18196 (N_18196,N_6829,N_9490);
nand U18197 (N_18197,N_6720,N_8589);
nand U18198 (N_18198,N_3192,N_9621);
nor U18199 (N_18199,N_5119,N_9396);
or U18200 (N_18200,N_9692,N_9507);
nand U18201 (N_18201,N_1493,N_956);
or U18202 (N_18202,N_2796,N_8251);
nor U18203 (N_18203,N_1170,N_4106);
nor U18204 (N_18204,N_1829,N_5912);
xnor U18205 (N_18205,N_5591,N_2604);
or U18206 (N_18206,N_3507,N_2444);
nand U18207 (N_18207,N_4031,N_2309);
or U18208 (N_18208,N_5483,N_7475);
xnor U18209 (N_18209,N_1677,N_4307);
nand U18210 (N_18210,N_9345,N_2093);
nand U18211 (N_18211,N_3716,N_6931);
or U18212 (N_18212,N_188,N_8102);
nor U18213 (N_18213,N_4668,N_2774);
nand U18214 (N_18214,N_7146,N_6659);
and U18215 (N_18215,N_7370,N_3414);
or U18216 (N_18216,N_9476,N_5339);
or U18217 (N_18217,N_7979,N_5552);
nand U18218 (N_18218,N_9309,N_9001);
or U18219 (N_18219,N_2840,N_5883);
nor U18220 (N_18220,N_9402,N_1803);
xnor U18221 (N_18221,N_3438,N_5494);
or U18222 (N_18222,N_8508,N_5245);
or U18223 (N_18223,N_5098,N_28);
and U18224 (N_18224,N_692,N_8873);
or U18225 (N_18225,N_8770,N_8691);
nand U18226 (N_18226,N_8190,N_2124);
nand U18227 (N_18227,N_3310,N_968);
nand U18228 (N_18228,N_1886,N_7917);
and U18229 (N_18229,N_5918,N_2936);
xnor U18230 (N_18230,N_8633,N_4836);
nor U18231 (N_18231,N_5817,N_9779);
nor U18232 (N_18232,N_7484,N_3226);
xnor U18233 (N_18233,N_5074,N_8203);
and U18234 (N_18234,N_748,N_4560);
nor U18235 (N_18235,N_4654,N_4594);
xor U18236 (N_18236,N_7603,N_7094);
nand U18237 (N_18237,N_3063,N_819);
or U18238 (N_18238,N_7827,N_4323);
or U18239 (N_18239,N_6929,N_7496);
nor U18240 (N_18240,N_690,N_5520);
xnor U18241 (N_18241,N_7458,N_7313);
and U18242 (N_18242,N_1322,N_3559);
and U18243 (N_18243,N_4272,N_2690);
nand U18244 (N_18244,N_3949,N_7468);
nand U18245 (N_18245,N_6256,N_3500);
nor U18246 (N_18246,N_4092,N_6800);
nand U18247 (N_18247,N_2262,N_2949);
xor U18248 (N_18248,N_9847,N_2085);
or U18249 (N_18249,N_5267,N_1060);
and U18250 (N_18250,N_9760,N_8327);
and U18251 (N_18251,N_975,N_1097);
nor U18252 (N_18252,N_8325,N_6378);
or U18253 (N_18253,N_6910,N_9893);
xor U18254 (N_18254,N_4880,N_549);
and U18255 (N_18255,N_4053,N_8461);
and U18256 (N_18256,N_1593,N_8647);
xnor U18257 (N_18257,N_6839,N_3103);
or U18258 (N_18258,N_3978,N_5501);
or U18259 (N_18259,N_4078,N_8182);
nand U18260 (N_18260,N_3094,N_5130);
nand U18261 (N_18261,N_114,N_139);
nand U18262 (N_18262,N_1592,N_406);
nand U18263 (N_18263,N_8033,N_4488);
xor U18264 (N_18264,N_7590,N_160);
or U18265 (N_18265,N_157,N_2678);
and U18266 (N_18266,N_7825,N_1132);
nor U18267 (N_18267,N_8618,N_495);
nand U18268 (N_18268,N_3819,N_440);
nand U18269 (N_18269,N_7030,N_5775);
nand U18270 (N_18270,N_4950,N_8193);
nor U18271 (N_18271,N_8785,N_6199);
or U18272 (N_18272,N_5049,N_6304);
and U18273 (N_18273,N_7335,N_794);
nand U18274 (N_18274,N_9447,N_732);
or U18275 (N_18275,N_4052,N_2810);
nor U18276 (N_18276,N_1414,N_3217);
xor U18277 (N_18277,N_3880,N_6988);
xnor U18278 (N_18278,N_271,N_5002);
or U18279 (N_18279,N_1556,N_6264);
xnor U18280 (N_18280,N_7083,N_1895);
and U18281 (N_18281,N_6365,N_132);
or U18282 (N_18282,N_3859,N_599);
nand U18283 (N_18283,N_243,N_4223);
or U18284 (N_18284,N_7125,N_2422);
and U18285 (N_18285,N_2913,N_2581);
xor U18286 (N_18286,N_6029,N_5059);
or U18287 (N_18287,N_2214,N_7892);
or U18288 (N_18288,N_9277,N_921);
nand U18289 (N_18289,N_891,N_7459);
xnor U18290 (N_18290,N_9630,N_916);
xnor U18291 (N_18291,N_3753,N_6210);
nor U18292 (N_18292,N_3556,N_3896);
xnor U18293 (N_18293,N_4417,N_6338);
and U18294 (N_18294,N_6144,N_9699);
xnor U18295 (N_18295,N_1513,N_629);
nand U18296 (N_18296,N_1735,N_4994);
xor U18297 (N_18297,N_2122,N_680);
nand U18298 (N_18298,N_5994,N_9970);
nor U18299 (N_18299,N_1616,N_7589);
nand U18300 (N_18300,N_5691,N_8923);
or U18301 (N_18301,N_745,N_570);
nand U18302 (N_18302,N_6093,N_4291);
nor U18303 (N_18303,N_9548,N_1597);
nand U18304 (N_18304,N_6392,N_4932);
nand U18305 (N_18305,N_3261,N_7743);
nand U18306 (N_18306,N_604,N_1079);
and U18307 (N_18307,N_323,N_3536);
xor U18308 (N_18308,N_2179,N_4838);
or U18309 (N_18309,N_4548,N_1172);
nand U18310 (N_18310,N_9407,N_9420);
nand U18311 (N_18311,N_9411,N_1678);
nor U18312 (N_18312,N_6339,N_9587);
xnor U18313 (N_18313,N_1273,N_5575);
nor U18314 (N_18314,N_4079,N_840);
nor U18315 (N_18315,N_8361,N_2283);
or U18316 (N_18316,N_4012,N_6638);
nor U18317 (N_18317,N_7412,N_3726);
and U18318 (N_18318,N_5829,N_3661);
nand U18319 (N_18319,N_6946,N_7877);
and U18320 (N_18320,N_8723,N_4846);
or U18321 (N_18321,N_4536,N_4518);
and U18322 (N_18322,N_8578,N_4227);
and U18323 (N_18323,N_5023,N_7800);
or U18324 (N_18324,N_3739,N_5085);
nor U18325 (N_18325,N_9604,N_2061);
xnor U18326 (N_18326,N_3802,N_4593);
or U18327 (N_18327,N_7586,N_52);
nor U18328 (N_18328,N_4657,N_8652);
nor U18329 (N_18329,N_3649,N_4323);
xnor U18330 (N_18330,N_3388,N_240);
nor U18331 (N_18331,N_8161,N_6110);
and U18332 (N_18332,N_2053,N_3506);
xor U18333 (N_18333,N_4905,N_7234);
and U18334 (N_18334,N_6387,N_6123);
nand U18335 (N_18335,N_8604,N_9519);
nor U18336 (N_18336,N_8985,N_6093);
and U18337 (N_18337,N_7502,N_9623);
xnor U18338 (N_18338,N_7447,N_4989);
or U18339 (N_18339,N_817,N_2546);
xnor U18340 (N_18340,N_8217,N_7054);
and U18341 (N_18341,N_5429,N_5902);
nand U18342 (N_18342,N_8043,N_6912);
nor U18343 (N_18343,N_5870,N_8356);
and U18344 (N_18344,N_7975,N_2071);
nor U18345 (N_18345,N_180,N_5598);
and U18346 (N_18346,N_1236,N_8640);
nor U18347 (N_18347,N_5045,N_710);
and U18348 (N_18348,N_9810,N_3902);
nor U18349 (N_18349,N_7059,N_7760);
nor U18350 (N_18350,N_6886,N_1396);
or U18351 (N_18351,N_6702,N_2621);
xor U18352 (N_18352,N_8349,N_6469);
xor U18353 (N_18353,N_5087,N_7863);
nor U18354 (N_18354,N_3527,N_4474);
nand U18355 (N_18355,N_5757,N_9701);
and U18356 (N_18356,N_4282,N_5790);
or U18357 (N_18357,N_3809,N_131);
xnor U18358 (N_18358,N_5051,N_4528);
xor U18359 (N_18359,N_184,N_9572);
nor U18360 (N_18360,N_7526,N_7223);
xnor U18361 (N_18361,N_6106,N_6419);
and U18362 (N_18362,N_2802,N_7215);
and U18363 (N_18363,N_2410,N_415);
and U18364 (N_18364,N_2302,N_3731);
or U18365 (N_18365,N_5583,N_2241);
nand U18366 (N_18366,N_9411,N_3213);
nand U18367 (N_18367,N_5472,N_7301);
nand U18368 (N_18368,N_3348,N_8447);
nor U18369 (N_18369,N_7316,N_5342);
or U18370 (N_18370,N_6411,N_9741);
xnor U18371 (N_18371,N_4797,N_9330);
nand U18372 (N_18372,N_3677,N_1053);
nor U18373 (N_18373,N_4744,N_7007);
nand U18374 (N_18374,N_1953,N_4557);
or U18375 (N_18375,N_6432,N_1419);
nor U18376 (N_18376,N_6880,N_4004);
nand U18377 (N_18377,N_2987,N_3138);
and U18378 (N_18378,N_9927,N_3989);
or U18379 (N_18379,N_7491,N_4294);
nand U18380 (N_18380,N_7295,N_8664);
and U18381 (N_18381,N_5375,N_8772);
nor U18382 (N_18382,N_9319,N_121);
xnor U18383 (N_18383,N_6139,N_4762);
xor U18384 (N_18384,N_8406,N_5081);
xor U18385 (N_18385,N_1247,N_7033);
xor U18386 (N_18386,N_462,N_4953);
and U18387 (N_18387,N_1085,N_2409);
and U18388 (N_18388,N_1457,N_3210);
nor U18389 (N_18389,N_2078,N_5254);
and U18390 (N_18390,N_1214,N_3771);
nor U18391 (N_18391,N_8507,N_1111);
and U18392 (N_18392,N_4105,N_3544);
nor U18393 (N_18393,N_2438,N_1601);
nand U18394 (N_18394,N_9799,N_1532);
nand U18395 (N_18395,N_2821,N_9644);
nor U18396 (N_18396,N_1738,N_2145);
nor U18397 (N_18397,N_2272,N_3287);
nor U18398 (N_18398,N_7727,N_4574);
xnor U18399 (N_18399,N_6934,N_1509);
nor U18400 (N_18400,N_920,N_6180);
nor U18401 (N_18401,N_2791,N_691);
and U18402 (N_18402,N_6823,N_65);
xnor U18403 (N_18403,N_3295,N_9492);
or U18404 (N_18404,N_9015,N_3466);
or U18405 (N_18405,N_8536,N_9849);
and U18406 (N_18406,N_8034,N_5725);
nand U18407 (N_18407,N_5097,N_7801);
nor U18408 (N_18408,N_5804,N_7925);
nand U18409 (N_18409,N_4137,N_4071);
nand U18410 (N_18410,N_7987,N_9582);
or U18411 (N_18411,N_3208,N_8218);
nand U18412 (N_18412,N_5225,N_2488);
xnor U18413 (N_18413,N_7092,N_4525);
xor U18414 (N_18414,N_1873,N_8833);
or U18415 (N_18415,N_1631,N_9437);
xnor U18416 (N_18416,N_4651,N_4594);
nand U18417 (N_18417,N_2793,N_385);
xnor U18418 (N_18418,N_5821,N_5199);
xnor U18419 (N_18419,N_1058,N_202);
and U18420 (N_18420,N_2279,N_6324);
or U18421 (N_18421,N_8462,N_1648);
and U18422 (N_18422,N_3412,N_3493);
and U18423 (N_18423,N_5078,N_2968);
nor U18424 (N_18424,N_7025,N_2737);
and U18425 (N_18425,N_2204,N_5084);
nor U18426 (N_18426,N_4635,N_4498);
or U18427 (N_18427,N_4891,N_2829);
nand U18428 (N_18428,N_8621,N_755);
or U18429 (N_18429,N_2005,N_4557);
and U18430 (N_18430,N_8082,N_28);
xnor U18431 (N_18431,N_3148,N_4242);
or U18432 (N_18432,N_6989,N_28);
and U18433 (N_18433,N_130,N_2187);
xor U18434 (N_18434,N_9546,N_5732);
xnor U18435 (N_18435,N_5612,N_5557);
nand U18436 (N_18436,N_7129,N_6812);
xor U18437 (N_18437,N_8266,N_1092);
nand U18438 (N_18438,N_7747,N_5801);
nand U18439 (N_18439,N_5707,N_2970);
and U18440 (N_18440,N_5789,N_3045);
xor U18441 (N_18441,N_5551,N_1858);
or U18442 (N_18442,N_9434,N_5184);
or U18443 (N_18443,N_1221,N_6926);
xnor U18444 (N_18444,N_6695,N_5857);
xnor U18445 (N_18445,N_4589,N_3172);
nand U18446 (N_18446,N_90,N_4156);
or U18447 (N_18447,N_6323,N_9986);
and U18448 (N_18448,N_3311,N_7011);
xnor U18449 (N_18449,N_153,N_2599);
nand U18450 (N_18450,N_7527,N_2925);
or U18451 (N_18451,N_1833,N_6638);
xor U18452 (N_18452,N_9947,N_4125);
and U18453 (N_18453,N_2484,N_1284);
nor U18454 (N_18454,N_4015,N_8005);
nand U18455 (N_18455,N_318,N_800);
nor U18456 (N_18456,N_7583,N_106);
xor U18457 (N_18457,N_8824,N_9514);
nor U18458 (N_18458,N_5756,N_614);
nor U18459 (N_18459,N_5022,N_8707);
and U18460 (N_18460,N_7144,N_2559);
and U18461 (N_18461,N_8363,N_3929);
nand U18462 (N_18462,N_1700,N_6267);
and U18463 (N_18463,N_7989,N_6300);
nand U18464 (N_18464,N_302,N_165);
nand U18465 (N_18465,N_7804,N_1825);
or U18466 (N_18466,N_9330,N_3653);
and U18467 (N_18467,N_5450,N_873);
nand U18468 (N_18468,N_471,N_338);
nor U18469 (N_18469,N_3940,N_1826);
and U18470 (N_18470,N_849,N_6069);
nand U18471 (N_18471,N_6803,N_519);
nand U18472 (N_18472,N_4018,N_9655);
nor U18473 (N_18473,N_2432,N_8723);
and U18474 (N_18474,N_7155,N_5062);
nor U18475 (N_18475,N_9240,N_3088);
nor U18476 (N_18476,N_4780,N_3703);
nor U18477 (N_18477,N_777,N_2586);
or U18478 (N_18478,N_2050,N_6384);
nor U18479 (N_18479,N_8365,N_9756);
nor U18480 (N_18480,N_7666,N_7082);
or U18481 (N_18481,N_319,N_8495);
nor U18482 (N_18482,N_1818,N_5721);
nor U18483 (N_18483,N_8046,N_4288);
nor U18484 (N_18484,N_2023,N_2696);
nor U18485 (N_18485,N_1077,N_2423);
and U18486 (N_18486,N_1215,N_8046);
and U18487 (N_18487,N_549,N_2920);
nor U18488 (N_18488,N_7605,N_1407);
or U18489 (N_18489,N_9682,N_8260);
xnor U18490 (N_18490,N_1718,N_4236);
and U18491 (N_18491,N_5928,N_7781);
nand U18492 (N_18492,N_2270,N_9052);
or U18493 (N_18493,N_4711,N_8725);
xnor U18494 (N_18494,N_5344,N_6251);
or U18495 (N_18495,N_8741,N_6677);
nand U18496 (N_18496,N_3714,N_1254);
and U18497 (N_18497,N_2681,N_5605);
or U18498 (N_18498,N_1559,N_3919);
xnor U18499 (N_18499,N_5726,N_4370);
or U18500 (N_18500,N_6348,N_403);
nor U18501 (N_18501,N_2125,N_5557);
or U18502 (N_18502,N_838,N_1363);
xnor U18503 (N_18503,N_4808,N_9105);
nand U18504 (N_18504,N_9522,N_3392);
and U18505 (N_18505,N_4081,N_9714);
and U18506 (N_18506,N_422,N_1389);
or U18507 (N_18507,N_4612,N_9865);
or U18508 (N_18508,N_6692,N_9569);
or U18509 (N_18509,N_6067,N_7365);
or U18510 (N_18510,N_6473,N_9042);
and U18511 (N_18511,N_1086,N_3185);
nand U18512 (N_18512,N_2574,N_629);
nand U18513 (N_18513,N_522,N_5901);
and U18514 (N_18514,N_4335,N_141);
nand U18515 (N_18515,N_4498,N_2924);
or U18516 (N_18516,N_4950,N_8511);
xor U18517 (N_18517,N_3999,N_6979);
xor U18518 (N_18518,N_5633,N_5545);
or U18519 (N_18519,N_7308,N_9090);
and U18520 (N_18520,N_4941,N_463);
and U18521 (N_18521,N_2092,N_7004);
and U18522 (N_18522,N_3130,N_8831);
nand U18523 (N_18523,N_693,N_6020);
and U18524 (N_18524,N_8749,N_8997);
xnor U18525 (N_18525,N_7051,N_6002);
nor U18526 (N_18526,N_2160,N_1091);
and U18527 (N_18527,N_6583,N_749);
or U18528 (N_18528,N_3969,N_3042);
or U18529 (N_18529,N_163,N_4489);
nand U18530 (N_18530,N_4682,N_7444);
nor U18531 (N_18531,N_4761,N_1952);
xor U18532 (N_18532,N_694,N_7736);
or U18533 (N_18533,N_6943,N_5108);
nand U18534 (N_18534,N_6024,N_5435);
xnor U18535 (N_18535,N_4197,N_6321);
xnor U18536 (N_18536,N_1233,N_6147);
nor U18537 (N_18537,N_8062,N_7843);
or U18538 (N_18538,N_5026,N_2360);
nand U18539 (N_18539,N_7745,N_1879);
nor U18540 (N_18540,N_1585,N_5698);
xor U18541 (N_18541,N_1648,N_4803);
nor U18542 (N_18542,N_8661,N_3735);
or U18543 (N_18543,N_9878,N_1486);
nand U18544 (N_18544,N_6837,N_8726);
and U18545 (N_18545,N_7717,N_7712);
and U18546 (N_18546,N_3587,N_9385);
nor U18547 (N_18547,N_6581,N_79);
xnor U18548 (N_18548,N_5422,N_2504);
nand U18549 (N_18549,N_9460,N_2441);
xor U18550 (N_18550,N_8956,N_1789);
and U18551 (N_18551,N_1670,N_6768);
nand U18552 (N_18552,N_8956,N_8676);
xnor U18553 (N_18553,N_3461,N_1190);
and U18554 (N_18554,N_1318,N_2060);
xnor U18555 (N_18555,N_7809,N_4815);
and U18556 (N_18556,N_9575,N_6761);
nor U18557 (N_18557,N_1453,N_8996);
or U18558 (N_18558,N_3877,N_33);
nand U18559 (N_18559,N_1135,N_5550);
xnor U18560 (N_18560,N_5709,N_2738);
and U18561 (N_18561,N_4371,N_9452);
nand U18562 (N_18562,N_2659,N_4256);
xor U18563 (N_18563,N_9765,N_4132);
and U18564 (N_18564,N_6044,N_6684);
xor U18565 (N_18565,N_9036,N_8124);
xor U18566 (N_18566,N_7130,N_5105);
or U18567 (N_18567,N_6245,N_9986);
xnor U18568 (N_18568,N_604,N_2505);
nand U18569 (N_18569,N_233,N_3157);
or U18570 (N_18570,N_3865,N_7360);
and U18571 (N_18571,N_5174,N_8687);
xor U18572 (N_18572,N_8901,N_6779);
or U18573 (N_18573,N_1513,N_4506);
nand U18574 (N_18574,N_2395,N_1012);
or U18575 (N_18575,N_7027,N_1568);
nor U18576 (N_18576,N_5445,N_1996);
or U18577 (N_18577,N_2091,N_1118);
or U18578 (N_18578,N_7118,N_9621);
or U18579 (N_18579,N_3922,N_2221);
and U18580 (N_18580,N_9093,N_497);
and U18581 (N_18581,N_5296,N_692);
nand U18582 (N_18582,N_5765,N_5490);
nor U18583 (N_18583,N_7239,N_9467);
nand U18584 (N_18584,N_9779,N_3859);
nor U18585 (N_18585,N_5241,N_3832);
nand U18586 (N_18586,N_7846,N_330);
and U18587 (N_18587,N_7595,N_6822);
xnor U18588 (N_18588,N_1729,N_2526);
nand U18589 (N_18589,N_3371,N_9073);
xor U18590 (N_18590,N_2917,N_4240);
nand U18591 (N_18591,N_92,N_5143);
and U18592 (N_18592,N_9849,N_7781);
nand U18593 (N_18593,N_5553,N_3634);
and U18594 (N_18594,N_9651,N_9189);
and U18595 (N_18595,N_8212,N_2544);
and U18596 (N_18596,N_6397,N_8114);
nor U18597 (N_18597,N_9287,N_4360);
nand U18598 (N_18598,N_9998,N_2639);
and U18599 (N_18599,N_1569,N_2266);
or U18600 (N_18600,N_3970,N_7573);
nor U18601 (N_18601,N_5074,N_8174);
nor U18602 (N_18602,N_1334,N_8136);
or U18603 (N_18603,N_1991,N_9283);
xor U18604 (N_18604,N_912,N_3540);
nor U18605 (N_18605,N_4949,N_402);
xnor U18606 (N_18606,N_7623,N_5720);
or U18607 (N_18607,N_2039,N_2256);
and U18608 (N_18608,N_7848,N_8529);
and U18609 (N_18609,N_5621,N_2642);
nor U18610 (N_18610,N_9635,N_2452);
nand U18611 (N_18611,N_8901,N_5516);
nor U18612 (N_18612,N_9537,N_957);
or U18613 (N_18613,N_2587,N_6565);
nor U18614 (N_18614,N_9781,N_4060);
nand U18615 (N_18615,N_1010,N_4129);
and U18616 (N_18616,N_6109,N_8100);
nor U18617 (N_18617,N_3264,N_9939);
xnor U18618 (N_18618,N_7132,N_6815);
and U18619 (N_18619,N_2905,N_9413);
or U18620 (N_18620,N_9929,N_2323);
nor U18621 (N_18621,N_3391,N_2270);
xnor U18622 (N_18622,N_3040,N_5276);
nor U18623 (N_18623,N_9236,N_1130);
nor U18624 (N_18624,N_8780,N_7451);
nand U18625 (N_18625,N_2239,N_1133);
nand U18626 (N_18626,N_9747,N_7351);
xor U18627 (N_18627,N_3288,N_712);
or U18628 (N_18628,N_2507,N_6856);
or U18629 (N_18629,N_3520,N_3154);
and U18630 (N_18630,N_902,N_9746);
xnor U18631 (N_18631,N_8695,N_386);
nand U18632 (N_18632,N_7044,N_9928);
nand U18633 (N_18633,N_3158,N_4232);
nand U18634 (N_18634,N_2567,N_8326);
and U18635 (N_18635,N_1456,N_2612);
nor U18636 (N_18636,N_8939,N_3532);
nor U18637 (N_18637,N_4077,N_2597);
and U18638 (N_18638,N_2584,N_3254);
nand U18639 (N_18639,N_7959,N_6344);
or U18640 (N_18640,N_1139,N_6583);
or U18641 (N_18641,N_4745,N_7676);
xor U18642 (N_18642,N_5642,N_5711);
and U18643 (N_18643,N_1634,N_3154);
and U18644 (N_18644,N_6816,N_4260);
and U18645 (N_18645,N_1968,N_2355);
and U18646 (N_18646,N_3645,N_7333);
and U18647 (N_18647,N_5233,N_6022);
nand U18648 (N_18648,N_8133,N_3591);
nand U18649 (N_18649,N_7671,N_4811);
and U18650 (N_18650,N_3524,N_9928);
or U18651 (N_18651,N_9801,N_5756);
or U18652 (N_18652,N_8759,N_7826);
and U18653 (N_18653,N_478,N_6658);
nor U18654 (N_18654,N_311,N_7627);
and U18655 (N_18655,N_1165,N_8036);
xnor U18656 (N_18656,N_4678,N_6715);
nand U18657 (N_18657,N_8804,N_4839);
nor U18658 (N_18658,N_3827,N_617);
and U18659 (N_18659,N_6052,N_828);
nand U18660 (N_18660,N_6257,N_8432);
nand U18661 (N_18661,N_924,N_8377);
nand U18662 (N_18662,N_394,N_9663);
or U18663 (N_18663,N_1122,N_6741);
nand U18664 (N_18664,N_7828,N_9332);
nor U18665 (N_18665,N_7709,N_2021);
nor U18666 (N_18666,N_9855,N_3322);
nand U18667 (N_18667,N_3885,N_6547);
nor U18668 (N_18668,N_7142,N_9189);
and U18669 (N_18669,N_9791,N_3125);
nor U18670 (N_18670,N_9181,N_5450);
nand U18671 (N_18671,N_5105,N_4348);
nor U18672 (N_18672,N_2169,N_6645);
or U18673 (N_18673,N_8032,N_1869);
nand U18674 (N_18674,N_5482,N_7627);
nor U18675 (N_18675,N_4496,N_3596);
nor U18676 (N_18676,N_6121,N_5807);
nand U18677 (N_18677,N_4464,N_8618);
xnor U18678 (N_18678,N_7801,N_7587);
and U18679 (N_18679,N_6201,N_8189);
nand U18680 (N_18680,N_5997,N_5074);
or U18681 (N_18681,N_9755,N_962);
and U18682 (N_18682,N_3221,N_3654);
and U18683 (N_18683,N_8375,N_2462);
nor U18684 (N_18684,N_3334,N_3596);
and U18685 (N_18685,N_3923,N_8);
and U18686 (N_18686,N_4580,N_5472);
nand U18687 (N_18687,N_5694,N_2258);
nand U18688 (N_18688,N_8828,N_7583);
and U18689 (N_18689,N_115,N_6737);
xnor U18690 (N_18690,N_6265,N_3964);
nand U18691 (N_18691,N_918,N_4969);
nand U18692 (N_18692,N_7426,N_4193);
xor U18693 (N_18693,N_20,N_4734);
or U18694 (N_18694,N_8380,N_9632);
and U18695 (N_18695,N_7002,N_8246);
and U18696 (N_18696,N_6601,N_6558);
nand U18697 (N_18697,N_5624,N_994);
xor U18698 (N_18698,N_8924,N_3143);
and U18699 (N_18699,N_2746,N_9689);
and U18700 (N_18700,N_8699,N_7403);
nor U18701 (N_18701,N_3541,N_187);
xor U18702 (N_18702,N_5620,N_8013);
xnor U18703 (N_18703,N_9835,N_6999);
xor U18704 (N_18704,N_5756,N_5581);
xor U18705 (N_18705,N_7529,N_4329);
xnor U18706 (N_18706,N_1121,N_3019);
or U18707 (N_18707,N_3041,N_349);
nor U18708 (N_18708,N_7992,N_6121);
and U18709 (N_18709,N_3847,N_2739);
or U18710 (N_18710,N_81,N_540);
nor U18711 (N_18711,N_3201,N_724);
or U18712 (N_18712,N_7176,N_9418);
nor U18713 (N_18713,N_8368,N_4132);
xor U18714 (N_18714,N_6619,N_9115);
xnor U18715 (N_18715,N_1966,N_9466);
and U18716 (N_18716,N_88,N_6806);
nand U18717 (N_18717,N_9994,N_7771);
nand U18718 (N_18718,N_3288,N_1519);
xnor U18719 (N_18719,N_8875,N_8571);
xnor U18720 (N_18720,N_9607,N_1093);
xor U18721 (N_18721,N_7381,N_2001);
and U18722 (N_18722,N_2438,N_6241);
nand U18723 (N_18723,N_3117,N_6220);
and U18724 (N_18724,N_8751,N_6433);
xor U18725 (N_18725,N_5170,N_9880);
or U18726 (N_18726,N_9115,N_1673);
and U18727 (N_18727,N_5766,N_2938);
and U18728 (N_18728,N_4333,N_1309);
or U18729 (N_18729,N_9316,N_4578);
and U18730 (N_18730,N_2628,N_695);
nor U18731 (N_18731,N_580,N_5295);
and U18732 (N_18732,N_4500,N_8112);
nand U18733 (N_18733,N_5614,N_7013);
nor U18734 (N_18734,N_564,N_9558);
or U18735 (N_18735,N_5301,N_8477);
or U18736 (N_18736,N_1341,N_8008);
xor U18737 (N_18737,N_6545,N_3727);
xor U18738 (N_18738,N_3949,N_4067);
nand U18739 (N_18739,N_931,N_5992);
nand U18740 (N_18740,N_5781,N_9865);
and U18741 (N_18741,N_2356,N_187);
xnor U18742 (N_18742,N_2171,N_9660);
nand U18743 (N_18743,N_6941,N_900);
nor U18744 (N_18744,N_8757,N_6855);
or U18745 (N_18745,N_2259,N_5187);
or U18746 (N_18746,N_2216,N_8241);
xor U18747 (N_18747,N_5019,N_5390);
or U18748 (N_18748,N_5683,N_2646);
xnor U18749 (N_18749,N_5883,N_5195);
and U18750 (N_18750,N_2788,N_7404);
nor U18751 (N_18751,N_3227,N_496);
nand U18752 (N_18752,N_5630,N_8158);
xnor U18753 (N_18753,N_916,N_8776);
xor U18754 (N_18754,N_3158,N_6909);
or U18755 (N_18755,N_7630,N_5288);
xnor U18756 (N_18756,N_1158,N_6321);
nand U18757 (N_18757,N_6646,N_5264);
xnor U18758 (N_18758,N_3328,N_809);
and U18759 (N_18759,N_1107,N_7548);
and U18760 (N_18760,N_2277,N_7699);
nor U18761 (N_18761,N_2295,N_8133);
or U18762 (N_18762,N_1023,N_8303);
and U18763 (N_18763,N_4375,N_533);
xnor U18764 (N_18764,N_5370,N_3651);
nand U18765 (N_18765,N_5760,N_9469);
nand U18766 (N_18766,N_1934,N_4597);
or U18767 (N_18767,N_5826,N_82);
and U18768 (N_18768,N_3547,N_466);
xnor U18769 (N_18769,N_6647,N_5398);
nand U18770 (N_18770,N_7388,N_1068);
or U18771 (N_18771,N_3550,N_8637);
xor U18772 (N_18772,N_7367,N_4682);
and U18773 (N_18773,N_4265,N_5302);
and U18774 (N_18774,N_1112,N_1259);
or U18775 (N_18775,N_98,N_2501);
and U18776 (N_18776,N_1678,N_2333);
xor U18777 (N_18777,N_7746,N_7788);
nor U18778 (N_18778,N_2380,N_8701);
or U18779 (N_18779,N_8714,N_2316);
and U18780 (N_18780,N_3947,N_4861);
nand U18781 (N_18781,N_6755,N_3642);
xor U18782 (N_18782,N_102,N_5428);
nor U18783 (N_18783,N_1225,N_9876);
nand U18784 (N_18784,N_4000,N_1839);
nand U18785 (N_18785,N_7346,N_6933);
nor U18786 (N_18786,N_6942,N_7633);
nand U18787 (N_18787,N_5900,N_243);
and U18788 (N_18788,N_7184,N_7132);
nand U18789 (N_18789,N_9468,N_6307);
or U18790 (N_18790,N_6927,N_102);
and U18791 (N_18791,N_8056,N_9652);
and U18792 (N_18792,N_6781,N_1567);
nand U18793 (N_18793,N_2216,N_285);
nor U18794 (N_18794,N_6711,N_3954);
xnor U18795 (N_18795,N_2928,N_8786);
nor U18796 (N_18796,N_9572,N_7159);
or U18797 (N_18797,N_9861,N_2338);
or U18798 (N_18798,N_5418,N_1747);
nand U18799 (N_18799,N_7403,N_8446);
xor U18800 (N_18800,N_1951,N_3900);
or U18801 (N_18801,N_8537,N_8737);
xnor U18802 (N_18802,N_9614,N_111);
or U18803 (N_18803,N_6398,N_4577);
and U18804 (N_18804,N_5250,N_8178);
nand U18805 (N_18805,N_3892,N_3074);
nand U18806 (N_18806,N_4559,N_6445);
xor U18807 (N_18807,N_3396,N_6140);
nand U18808 (N_18808,N_8843,N_3041);
nor U18809 (N_18809,N_2083,N_7174);
and U18810 (N_18810,N_5377,N_6791);
nor U18811 (N_18811,N_4884,N_8833);
and U18812 (N_18812,N_1846,N_5478);
nand U18813 (N_18813,N_5967,N_8547);
nand U18814 (N_18814,N_2701,N_9798);
nor U18815 (N_18815,N_1033,N_8942);
nor U18816 (N_18816,N_5943,N_6054);
xnor U18817 (N_18817,N_6018,N_8624);
or U18818 (N_18818,N_9118,N_7815);
nor U18819 (N_18819,N_8648,N_7781);
nor U18820 (N_18820,N_3671,N_4385);
and U18821 (N_18821,N_8038,N_165);
nor U18822 (N_18822,N_4228,N_6853);
nand U18823 (N_18823,N_1969,N_809);
and U18824 (N_18824,N_3166,N_9345);
nand U18825 (N_18825,N_2835,N_6219);
nand U18826 (N_18826,N_9722,N_1252);
nor U18827 (N_18827,N_2335,N_5352);
xor U18828 (N_18828,N_3543,N_6938);
nor U18829 (N_18829,N_5832,N_3617);
or U18830 (N_18830,N_9544,N_3339);
nor U18831 (N_18831,N_128,N_9750);
or U18832 (N_18832,N_2080,N_2539);
nand U18833 (N_18833,N_3915,N_5711);
and U18834 (N_18834,N_6947,N_4802);
nand U18835 (N_18835,N_8452,N_5342);
or U18836 (N_18836,N_4978,N_790);
nand U18837 (N_18837,N_2483,N_663);
nor U18838 (N_18838,N_2547,N_9890);
nor U18839 (N_18839,N_2880,N_7767);
nor U18840 (N_18840,N_8135,N_6157);
and U18841 (N_18841,N_6636,N_1661);
and U18842 (N_18842,N_1454,N_606);
nand U18843 (N_18843,N_2013,N_1062);
and U18844 (N_18844,N_6406,N_2922);
xor U18845 (N_18845,N_530,N_4433);
nor U18846 (N_18846,N_8498,N_6157);
nand U18847 (N_18847,N_6822,N_9635);
nor U18848 (N_18848,N_7921,N_4097);
nand U18849 (N_18849,N_5282,N_8737);
nor U18850 (N_18850,N_8960,N_7845);
and U18851 (N_18851,N_7027,N_3322);
and U18852 (N_18852,N_5892,N_1490);
xnor U18853 (N_18853,N_4316,N_3203);
and U18854 (N_18854,N_5622,N_4746);
nand U18855 (N_18855,N_7891,N_5961);
or U18856 (N_18856,N_9655,N_5682);
nand U18857 (N_18857,N_5517,N_1675);
nand U18858 (N_18858,N_3101,N_3120);
or U18859 (N_18859,N_7006,N_1603);
and U18860 (N_18860,N_4990,N_1883);
and U18861 (N_18861,N_1282,N_7475);
xor U18862 (N_18862,N_5164,N_4417);
or U18863 (N_18863,N_8979,N_7528);
nand U18864 (N_18864,N_296,N_4307);
nand U18865 (N_18865,N_1219,N_4686);
nand U18866 (N_18866,N_1815,N_8397);
nor U18867 (N_18867,N_2487,N_7720);
or U18868 (N_18868,N_770,N_6673);
or U18869 (N_18869,N_4234,N_7578);
xnor U18870 (N_18870,N_8560,N_227);
nor U18871 (N_18871,N_4453,N_5691);
nor U18872 (N_18872,N_7659,N_3992);
nor U18873 (N_18873,N_9746,N_4406);
and U18874 (N_18874,N_2179,N_2653);
or U18875 (N_18875,N_1881,N_2007);
xor U18876 (N_18876,N_4168,N_4544);
nand U18877 (N_18877,N_5672,N_6807);
and U18878 (N_18878,N_6479,N_8831);
nand U18879 (N_18879,N_5248,N_2316);
xor U18880 (N_18880,N_2655,N_6548);
xor U18881 (N_18881,N_6696,N_1216);
nor U18882 (N_18882,N_5045,N_5087);
and U18883 (N_18883,N_5473,N_1540);
nand U18884 (N_18884,N_6457,N_5734);
or U18885 (N_18885,N_9446,N_3467);
nor U18886 (N_18886,N_8303,N_1167);
nor U18887 (N_18887,N_2138,N_6249);
nand U18888 (N_18888,N_7989,N_8974);
nand U18889 (N_18889,N_6688,N_2649);
and U18890 (N_18890,N_2388,N_4159);
nor U18891 (N_18891,N_2290,N_5739);
xor U18892 (N_18892,N_4336,N_380);
xnor U18893 (N_18893,N_9801,N_2322);
nor U18894 (N_18894,N_1431,N_6563);
nor U18895 (N_18895,N_5049,N_5675);
xor U18896 (N_18896,N_5386,N_9926);
and U18897 (N_18897,N_8783,N_1047);
xor U18898 (N_18898,N_7149,N_8257);
nand U18899 (N_18899,N_8423,N_7493);
nand U18900 (N_18900,N_4153,N_54);
or U18901 (N_18901,N_9183,N_9891);
nand U18902 (N_18902,N_6269,N_9872);
and U18903 (N_18903,N_2451,N_7826);
nand U18904 (N_18904,N_7163,N_6858);
or U18905 (N_18905,N_8880,N_1691);
or U18906 (N_18906,N_5541,N_142);
nand U18907 (N_18907,N_9373,N_1867);
nand U18908 (N_18908,N_9579,N_8192);
nor U18909 (N_18909,N_740,N_1632);
or U18910 (N_18910,N_3991,N_4981);
xor U18911 (N_18911,N_3930,N_4436);
or U18912 (N_18912,N_7268,N_405);
xnor U18913 (N_18913,N_250,N_1325);
nand U18914 (N_18914,N_6966,N_344);
nor U18915 (N_18915,N_2545,N_8841);
or U18916 (N_18916,N_1134,N_4520);
nor U18917 (N_18917,N_6842,N_8810);
and U18918 (N_18918,N_750,N_5392);
nand U18919 (N_18919,N_3090,N_6563);
and U18920 (N_18920,N_9478,N_8168);
nor U18921 (N_18921,N_7598,N_1870);
or U18922 (N_18922,N_8260,N_5006);
nand U18923 (N_18923,N_6166,N_9823);
and U18924 (N_18924,N_3079,N_9694);
or U18925 (N_18925,N_8801,N_7520);
nand U18926 (N_18926,N_5874,N_8850);
nand U18927 (N_18927,N_2743,N_2067);
xnor U18928 (N_18928,N_4798,N_7115);
nor U18929 (N_18929,N_1768,N_7794);
xnor U18930 (N_18930,N_1396,N_6844);
or U18931 (N_18931,N_3689,N_4658);
nand U18932 (N_18932,N_1922,N_6772);
nor U18933 (N_18933,N_1649,N_1329);
nand U18934 (N_18934,N_1933,N_7799);
nor U18935 (N_18935,N_1236,N_3844);
nor U18936 (N_18936,N_9962,N_1908);
nand U18937 (N_18937,N_1188,N_3193);
xor U18938 (N_18938,N_5399,N_5659);
or U18939 (N_18939,N_4684,N_5921);
nand U18940 (N_18940,N_334,N_8339);
nor U18941 (N_18941,N_6588,N_1565);
and U18942 (N_18942,N_4031,N_5556);
and U18943 (N_18943,N_2815,N_8632);
or U18944 (N_18944,N_472,N_703);
and U18945 (N_18945,N_3861,N_3955);
nand U18946 (N_18946,N_2179,N_4070);
and U18947 (N_18947,N_1395,N_3046);
and U18948 (N_18948,N_7362,N_9100);
nand U18949 (N_18949,N_6282,N_2716);
xnor U18950 (N_18950,N_7005,N_1973);
nor U18951 (N_18951,N_3433,N_7941);
xnor U18952 (N_18952,N_4648,N_3311);
nor U18953 (N_18953,N_2959,N_4629);
xor U18954 (N_18954,N_5203,N_3103);
xor U18955 (N_18955,N_8693,N_6015);
and U18956 (N_18956,N_1911,N_7843);
nand U18957 (N_18957,N_2945,N_1245);
xnor U18958 (N_18958,N_5675,N_5969);
and U18959 (N_18959,N_6745,N_6661);
or U18960 (N_18960,N_1587,N_7762);
or U18961 (N_18961,N_8397,N_8183);
or U18962 (N_18962,N_6462,N_6737);
nand U18963 (N_18963,N_1932,N_2172);
nor U18964 (N_18964,N_1289,N_990);
xnor U18965 (N_18965,N_6192,N_2990);
xnor U18966 (N_18966,N_5293,N_6977);
and U18967 (N_18967,N_4847,N_1086);
and U18968 (N_18968,N_3898,N_5085);
xnor U18969 (N_18969,N_1966,N_7305);
xnor U18970 (N_18970,N_38,N_1165);
nor U18971 (N_18971,N_7566,N_7376);
nor U18972 (N_18972,N_1128,N_7289);
nand U18973 (N_18973,N_3945,N_2247);
nand U18974 (N_18974,N_1669,N_740);
nor U18975 (N_18975,N_9274,N_2756);
xnor U18976 (N_18976,N_9275,N_2932);
and U18977 (N_18977,N_4153,N_2094);
nand U18978 (N_18978,N_6414,N_1055);
nand U18979 (N_18979,N_5279,N_8924);
nand U18980 (N_18980,N_5689,N_6703);
xor U18981 (N_18981,N_8961,N_2578);
or U18982 (N_18982,N_2469,N_7718);
or U18983 (N_18983,N_9914,N_2972);
and U18984 (N_18984,N_7440,N_4833);
or U18985 (N_18985,N_4460,N_6293);
and U18986 (N_18986,N_8594,N_9973);
nand U18987 (N_18987,N_7950,N_3228);
nand U18988 (N_18988,N_9802,N_8934);
xor U18989 (N_18989,N_6771,N_6659);
or U18990 (N_18990,N_6852,N_9495);
xnor U18991 (N_18991,N_7388,N_1194);
and U18992 (N_18992,N_7004,N_9115);
xnor U18993 (N_18993,N_6038,N_7523);
or U18994 (N_18994,N_5483,N_1793);
or U18995 (N_18995,N_5660,N_6391);
nor U18996 (N_18996,N_7443,N_6883);
nor U18997 (N_18997,N_4740,N_7333);
nand U18998 (N_18998,N_4630,N_3507);
and U18999 (N_18999,N_7210,N_8583);
or U19000 (N_19000,N_3401,N_9152);
nand U19001 (N_19001,N_6425,N_5683);
or U19002 (N_19002,N_635,N_9039);
nor U19003 (N_19003,N_8632,N_5471);
nor U19004 (N_19004,N_9603,N_7417);
nor U19005 (N_19005,N_9570,N_3977);
and U19006 (N_19006,N_9583,N_4348);
nor U19007 (N_19007,N_6510,N_9902);
and U19008 (N_19008,N_9075,N_8495);
nand U19009 (N_19009,N_9930,N_6969);
and U19010 (N_19010,N_1479,N_8557);
or U19011 (N_19011,N_6215,N_8253);
nand U19012 (N_19012,N_5992,N_7249);
nand U19013 (N_19013,N_585,N_3859);
xor U19014 (N_19014,N_1079,N_6128);
nand U19015 (N_19015,N_6375,N_3461);
nor U19016 (N_19016,N_4596,N_8773);
xor U19017 (N_19017,N_292,N_8365);
xnor U19018 (N_19018,N_6125,N_2050);
or U19019 (N_19019,N_382,N_3626);
nor U19020 (N_19020,N_7002,N_9687);
and U19021 (N_19021,N_7921,N_328);
nand U19022 (N_19022,N_2911,N_2679);
nand U19023 (N_19023,N_8134,N_1513);
nand U19024 (N_19024,N_9497,N_619);
nand U19025 (N_19025,N_2022,N_7925);
and U19026 (N_19026,N_393,N_9980);
nor U19027 (N_19027,N_2905,N_7035);
nor U19028 (N_19028,N_7644,N_7733);
xnor U19029 (N_19029,N_6074,N_7797);
nor U19030 (N_19030,N_8652,N_4109);
nand U19031 (N_19031,N_1083,N_9895);
and U19032 (N_19032,N_9840,N_767);
and U19033 (N_19033,N_5191,N_7737);
and U19034 (N_19034,N_7157,N_84);
or U19035 (N_19035,N_8982,N_9876);
and U19036 (N_19036,N_9190,N_2463);
or U19037 (N_19037,N_277,N_9437);
or U19038 (N_19038,N_2032,N_739);
and U19039 (N_19039,N_4123,N_2670);
nor U19040 (N_19040,N_7928,N_5241);
and U19041 (N_19041,N_312,N_9935);
xor U19042 (N_19042,N_4832,N_573);
xor U19043 (N_19043,N_2206,N_2589);
nand U19044 (N_19044,N_2357,N_9562);
or U19045 (N_19045,N_5025,N_9913);
and U19046 (N_19046,N_2505,N_3660);
or U19047 (N_19047,N_5467,N_7786);
xnor U19048 (N_19048,N_4018,N_7846);
and U19049 (N_19049,N_6161,N_8257);
or U19050 (N_19050,N_7245,N_4224);
or U19051 (N_19051,N_4027,N_2027);
xnor U19052 (N_19052,N_6574,N_5775);
nand U19053 (N_19053,N_1695,N_5094);
nand U19054 (N_19054,N_6234,N_2430);
xor U19055 (N_19055,N_29,N_3174);
xor U19056 (N_19056,N_5455,N_9933);
and U19057 (N_19057,N_807,N_2188);
or U19058 (N_19058,N_1515,N_2605);
nor U19059 (N_19059,N_714,N_4315);
nand U19060 (N_19060,N_618,N_7595);
nor U19061 (N_19061,N_7592,N_3346);
and U19062 (N_19062,N_6783,N_6327);
and U19063 (N_19063,N_2593,N_2675);
or U19064 (N_19064,N_9892,N_2090);
or U19065 (N_19065,N_4285,N_7877);
xnor U19066 (N_19066,N_3525,N_333);
or U19067 (N_19067,N_1973,N_1507);
nand U19068 (N_19068,N_7447,N_1416);
xnor U19069 (N_19069,N_7174,N_3995);
or U19070 (N_19070,N_9564,N_581);
nor U19071 (N_19071,N_8049,N_2011);
nand U19072 (N_19072,N_4372,N_8179);
or U19073 (N_19073,N_3067,N_3763);
and U19074 (N_19074,N_3923,N_4600);
nor U19075 (N_19075,N_4367,N_960);
nor U19076 (N_19076,N_4024,N_302);
xnor U19077 (N_19077,N_4939,N_1904);
nand U19078 (N_19078,N_1995,N_7526);
and U19079 (N_19079,N_275,N_2367);
nand U19080 (N_19080,N_3729,N_1632);
nor U19081 (N_19081,N_8252,N_8270);
nand U19082 (N_19082,N_3578,N_3702);
or U19083 (N_19083,N_9604,N_4823);
or U19084 (N_19084,N_5939,N_7860);
or U19085 (N_19085,N_9130,N_5568);
nor U19086 (N_19086,N_539,N_5616);
nor U19087 (N_19087,N_4693,N_8826);
or U19088 (N_19088,N_2734,N_1022);
and U19089 (N_19089,N_362,N_3038);
xor U19090 (N_19090,N_2464,N_8020);
xnor U19091 (N_19091,N_1793,N_8041);
or U19092 (N_19092,N_8887,N_6750);
xor U19093 (N_19093,N_595,N_7779);
or U19094 (N_19094,N_1038,N_5241);
and U19095 (N_19095,N_3373,N_6369);
xor U19096 (N_19096,N_2436,N_9721);
xor U19097 (N_19097,N_7084,N_8575);
nor U19098 (N_19098,N_7449,N_8568);
and U19099 (N_19099,N_983,N_7356);
nor U19100 (N_19100,N_9245,N_2995);
and U19101 (N_19101,N_8166,N_3342);
or U19102 (N_19102,N_9379,N_9789);
and U19103 (N_19103,N_7427,N_4517);
and U19104 (N_19104,N_7928,N_6038);
and U19105 (N_19105,N_5395,N_7318);
or U19106 (N_19106,N_4992,N_7096);
nand U19107 (N_19107,N_5269,N_5939);
nor U19108 (N_19108,N_7419,N_3536);
and U19109 (N_19109,N_8642,N_4746);
xor U19110 (N_19110,N_5685,N_3158);
nand U19111 (N_19111,N_3491,N_5111);
and U19112 (N_19112,N_7555,N_1824);
xor U19113 (N_19113,N_6425,N_3689);
or U19114 (N_19114,N_9307,N_7455);
and U19115 (N_19115,N_3997,N_7382);
nand U19116 (N_19116,N_4836,N_3112);
or U19117 (N_19117,N_6775,N_9085);
xor U19118 (N_19118,N_4764,N_6986);
nor U19119 (N_19119,N_1192,N_3114);
xor U19120 (N_19120,N_3699,N_1439);
and U19121 (N_19121,N_2991,N_8404);
xor U19122 (N_19122,N_4689,N_4072);
xnor U19123 (N_19123,N_7021,N_8092);
and U19124 (N_19124,N_3905,N_6782);
and U19125 (N_19125,N_7027,N_9880);
nand U19126 (N_19126,N_1850,N_1108);
nor U19127 (N_19127,N_3127,N_9692);
xor U19128 (N_19128,N_6277,N_465);
xnor U19129 (N_19129,N_4144,N_2281);
xor U19130 (N_19130,N_3357,N_8634);
or U19131 (N_19131,N_999,N_8297);
and U19132 (N_19132,N_3795,N_6686);
nor U19133 (N_19133,N_2924,N_8740);
nor U19134 (N_19134,N_1643,N_4749);
nand U19135 (N_19135,N_9806,N_9012);
and U19136 (N_19136,N_1969,N_5066);
and U19137 (N_19137,N_8077,N_1114);
nand U19138 (N_19138,N_6153,N_939);
or U19139 (N_19139,N_3678,N_2648);
and U19140 (N_19140,N_7047,N_843);
nand U19141 (N_19141,N_1562,N_9334);
nand U19142 (N_19142,N_8762,N_351);
nand U19143 (N_19143,N_6963,N_9204);
or U19144 (N_19144,N_2385,N_1582);
and U19145 (N_19145,N_9541,N_8514);
xor U19146 (N_19146,N_5218,N_7651);
or U19147 (N_19147,N_8407,N_1609);
nand U19148 (N_19148,N_8981,N_1271);
nand U19149 (N_19149,N_7450,N_1837);
nor U19150 (N_19150,N_6704,N_4898);
and U19151 (N_19151,N_8764,N_2062);
and U19152 (N_19152,N_2522,N_8813);
xnor U19153 (N_19153,N_8912,N_9003);
or U19154 (N_19154,N_6590,N_8170);
nor U19155 (N_19155,N_7657,N_1806);
and U19156 (N_19156,N_986,N_3267);
and U19157 (N_19157,N_258,N_5749);
nand U19158 (N_19158,N_4668,N_1439);
xnor U19159 (N_19159,N_8676,N_8465);
nand U19160 (N_19160,N_6808,N_4241);
and U19161 (N_19161,N_7295,N_4189);
or U19162 (N_19162,N_3849,N_1802);
nand U19163 (N_19163,N_7007,N_9284);
or U19164 (N_19164,N_6544,N_6899);
or U19165 (N_19165,N_9473,N_3899);
nand U19166 (N_19166,N_9546,N_4796);
or U19167 (N_19167,N_8893,N_7752);
nor U19168 (N_19168,N_6058,N_3465);
xor U19169 (N_19169,N_87,N_4422);
nor U19170 (N_19170,N_7917,N_7959);
and U19171 (N_19171,N_1727,N_6355);
or U19172 (N_19172,N_8131,N_9040);
nand U19173 (N_19173,N_4219,N_2430);
nor U19174 (N_19174,N_1125,N_8377);
xor U19175 (N_19175,N_9270,N_1774);
and U19176 (N_19176,N_8345,N_777);
nor U19177 (N_19177,N_7278,N_1154);
nand U19178 (N_19178,N_5294,N_4917);
or U19179 (N_19179,N_8764,N_1908);
xnor U19180 (N_19180,N_5593,N_1870);
nand U19181 (N_19181,N_7202,N_2807);
or U19182 (N_19182,N_9630,N_179);
nand U19183 (N_19183,N_1309,N_5774);
xnor U19184 (N_19184,N_3883,N_9278);
nor U19185 (N_19185,N_1200,N_4583);
or U19186 (N_19186,N_8809,N_5613);
or U19187 (N_19187,N_5133,N_2500);
xnor U19188 (N_19188,N_2664,N_5606);
nor U19189 (N_19189,N_4243,N_7069);
and U19190 (N_19190,N_3608,N_4773);
or U19191 (N_19191,N_8021,N_5356);
nor U19192 (N_19192,N_6939,N_535);
and U19193 (N_19193,N_1673,N_2018);
and U19194 (N_19194,N_2930,N_7184);
or U19195 (N_19195,N_4734,N_8967);
nor U19196 (N_19196,N_5392,N_2411);
nand U19197 (N_19197,N_3233,N_5703);
nor U19198 (N_19198,N_4162,N_9505);
nand U19199 (N_19199,N_620,N_3088);
and U19200 (N_19200,N_6967,N_4527);
and U19201 (N_19201,N_3259,N_62);
xnor U19202 (N_19202,N_94,N_2816);
and U19203 (N_19203,N_4751,N_4428);
nand U19204 (N_19204,N_6914,N_3278);
xnor U19205 (N_19205,N_9194,N_2102);
nor U19206 (N_19206,N_2918,N_5745);
nor U19207 (N_19207,N_3370,N_8844);
xor U19208 (N_19208,N_8890,N_4635);
xor U19209 (N_19209,N_4743,N_5061);
nor U19210 (N_19210,N_5492,N_8954);
xnor U19211 (N_19211,N_9414,N_4819);
or U19212 (N_19212,N_9577,N_9039);
xnor U19213 (N_19213,N_3924,N_9823);
nor U19214 (N_19214,N_8352,N_9824);
nor U19215 (N_19215,N_2093,N_8749);
and U19216 (N_19216,N_5663,N_2140);
and U19217 (N_19217,N_3343,N_4266);
nor U19218 (N_19218,N_8635,N_6237);
nor U19219 (N_19219,N_2703,N_569);
xnor U19220 (N_19220,N_6442,N_8320);
or U19221 (N_19221,N_5778,N_8595);
or U19222 (N_19222,N_8710,N_9410);
nor U19223 (N_19223,N_4842,N_3605);
or U19224 (N_19224,N_4436,N_8135);
and U19225 (N_19225,N_3016,N_1118);
or U19226 (N_19226,N_7584,N_6983);
xor U19227 (N_19227,N_6831,N_3319);
or U19228 (N_19228,N_6502,N_5781);
nor U19229 (N_19229,N_8823,N_1203);
and U19230 (N_19230,N_539,N_2560);
nor U19231 (N_19231,N_1468,N_9794);
or U19232 (N_19232,N_4219,N_9560);
nor U19233 (N_19233,N_2326,N_221);
or U19234 (N_19234,N_7285,N_7949);
nor U19235 (N_19235,N_23,N_9722);
nand U19236 (N_19236,N_3956,N_5471);
or U19237 (N_19237,N_1975,N_261);
xnor U19238 (N_19238,N_4846,N_9580);
or U19239 (N_19239,N_5971,N_4080);
or U19240 (N_19240,N_3996,N_9216);
or U19241 (N_19241,N_8956,N_2268);
nor U19242 (N_19242,N_5473,N_4071);
nand U19243 (N_19243,N_78,N_588);
or U19244 (N_19244,N_831,N_987);
nand U19245 (N_19245,N_9718,N_3004);
nand U19246 (N_19246,N_800,N_8237);
nor U19247 (N_19247,N_9738,N_8);
nor U19248 (N_19248,N_4495,N_4166);
nor U19249 (N_19249,N_2679,N_8414);
nor U19250 (N_19250,N_6966,N_4944);
nand U19251 (N_19251,N_2994,N_4302);
or U19252 (N_19252,N_9427,N_8209);
or U19253 (N_19253,N_553,N_6463);
or U19254 (N_19254,N_7546,N_8008);
xor U19255 (N_19255,N_9668,N_5632);
xnor U19256 (N_19256,N_2218,N_2036);
or U19257 (N_19257,N_7831,N_5296);
nor U19258 (N_19258,N_2303,N_3402);
nand U19259 (N_19259,N_4187,N_3446);
xor U19260 (N_19260,N_2800,N_7308);
xnor U19261 (N_19261,N_137,N_169);
nand U19262 (N_19262,N_857,N_8012);
xnor U19263 (N_19263,N_1941,N_5118);
nand U19264 (N_19264,N_2624,N_2708);
and U19265 (N_19265,N_3623,N_8943);
nor U19266 (N_19266,N_7118,N_9769);
or U19267 (N_19267,N_4157,N_5085);
and U19268 (N_19268,N_9348,N_3347);
and U19269 (N_19269,N_7117,N_4713);
nand U19270 (N_19270,N_5807,N_7298);
xor U19271 (N_19271,N_653,N_1862);
and U19272 (N_19272,N_2034,N_6819);
and U19273 (N_19273,N_7535,N_409);
nand U19274 (N_19274,N_3105,N_50);
xor U19275 (N_19275,N_1417,N_4366);
and U19276 (N_19276,N_5779,N_4479);
or U19277 (N_19277,N_9339,N_6238);
xnor U19278 (N_19278,N_5602,N_1651);
nand U19279 (N_19279,N_2581,N_7892);
or U19280 (N_19280,N_2417,N_633);
nor U19281 (N_19281,N_345,N_335);
nand U19282 (N_19282,N_7725,N_4366);
nor U19283 (N_19283,N_9221,N_7167);
xnor U19284 (N_19284,N_4019,N_1237);
nor U19285 (N_19285,N_5678,N_3422);
nand U19286 (N_19286,N_8477,N_3307);
or U19287 (N_19287,N_7603,N_9685);
xor U19288 (N_19288,N_4728,N_6662);
or U19289 (N_19289,N_7430,N_8454);
xor U19290 (N_19290,N_1093,N_3267);
xor U19291 (N_19291,N_7343,N_5144);
or U19292 (N_19292,N_9710,N_8361);
xor U19293 (N_19293,N_3116,N_4337);
and U19294 (N_19294,N_8526,N_8926);
and U19295 (N_19295,N_7053,N_5957);
or U19296 (N_19296,N_4202,N_8550);
and U19297 (N_19297,N_913,N_918);
nor U19298 (N_19298,N_7971,N_9376);
or U19299 (N_19299,N_4597,N_2658);
nand U19300 (N_19300,N_6306,N_6750);
and U19301 (N_19301,N_2093,N_8645);
nor U19302 (N_19302,N_3175,N_7529);
or U19303 (N_19303,N_1288,N_2285);
or U19304 (N_19304,N_4633,N_4577);
xor U19305 (N_19305,N_6545,N_5137);
nand U19306 (N_19306,N_6356,N_9128);
nor U19307 (N_19307,N_1578,N_5274);
nor U19308 (N_19308,N_9504,N_208);
nor U19309 (N_19309,N_60,N_8480);
and U19310 (N_19310,N_5830,N_1386);
nor U19311 (N_19311,N_2548,N_2912);
or U19312 (N_19312,N_4257,N_6757);
or U19313 (N_19313,N_7089,N_8618);
and U19314 (N_19314,N_7936,N_2630);
xor U19315 (N_19315,N_563,N_3493);
xnor U19316 (N_19316,N_6091,N_1229);
or U19317 (N_19317,N_6713,N_5592);
nand U19318 (N_19318,N_2802,N_2951);
nand U19319 (N_19319,N_2077,N_2956);
nand U19320 (N_19320,N_4007,N_832);
nor U19321 (N_19321,N_4534,N_3946);
nor U19322 (N_19322,N_6540,N_3122);
xnor U19323 (N_19323,N_2197,N_5757);
or U19324 (N_19324,N_2332,N_6362);
xnor U19325 (N_19325,N_4203,N_1548);
xnor U19326 (N_19326,N_1032,N_1581);
nor U19327 (N_19327,N_3243,N_3093);
nor U19328 (N_19328,N_963,N_3176);
or U19329 (N_19329,N_3035,N_8759);
xnor U19330 (N_19330,N_5730,N_2660);
and U19331 (N_19331,N_1206,N_5194);
nand U19332 (N_19332,N_6049,N_1420);
nor U19333 (N_19333,N_6180,N_3095);
nand U19334 (N_19334,N_4861,N_1964);
nand U19335 (N_19335,N_5104,N_9431);
nor U19336 (N_19336,N_3622,N_6788);
nand U19337 (N_19337,N_7678,N_3284);
or U19338 (N_19338,N_7198,N_6388);
nand U19339 (N_19339,N_8896,N_800);
or U19340 (N_19340,N_9566,N_3648);
nand U19341 (N_19341,N_8669,N_8746);
nor U19342 (N_19342,N_5996,N_3959);
xnor U19343 (N_19343,N_237,N_811);
nor U19344 (N_19344,N_8321,N_9839);
xor U19345 (N_19345,N_6206,N_1028);
or U19346 (N_19346,N_3944,N_7468);
nand U19347 (N_19347,N_5552,N_9659);
nand U19348 (N_19348,N_8320,N_5085);
nand U19349 (N_19349,N_1240,N_882);
xnor U19350 (N_19350,N_123,N_4861);
xnor U19351 (N_19351,N_6587,N_8331);
nor U19352 (N_19352,N_8874,N_5639);
nor U19353 (N_19353,N_5916,N_6575);
or U19354 (N_19354,N_666,N_5317);
xor U19355 (N_19355,N_7687,N_5450);
xnor U19356 (N_19356,N_4495,N_9044);
nand U19357 (N_19357,N_7503,N_6899);
or U19358 (N_19358,N_6306,N_32);
and U19359 (N_19359,N_3880,N_8748);
or U19360 (N_19360,N_5201,N_1155);
and U19361 (N_19361,N_9814,N_4880);
nand U19362 (N_19362,N_8820,N_7672);
nand U19363 (N_19363,N_5842,N_6004);
nor U19364 (N_19364,N_4673,N_8175);
xnor U19365 (N_19365,N_43,N_2369);
nor U19366 (N_19366,N_411,N_8773);
and U19367 (N_19367,N_493,N_2651);
or U19368 (N_19368,N_8093,N_520);
and U19369 (N_19369,N_6285,N_5112);
nor U19370 (N_19370,N_7664,N_3735);
or U19371 (N_19371,N_2163,N_7130);
nand U19372 (N_19372,N_427,N_5797);
nand U19373 (N_19373,N_9309,N_7066);
xor U19374 (N_19374,N_1262,N_1048);
nand U19375 (N_19375,N_2936,N_4241);
nor U19376 (N_19376,N_3678,N_1689);
nand U19377 (N_19377,N_4299,N_6739);
and U19378 (N_19378,N_7355,N_442);
or U19379 (N_19379,N_8306,N_9198);
nor U19380 (N_19380,N_2837,N_3995);
or U19381 (N_19381,N_7148,N_3608);
nor U19382 (N_19382,N_4895,N_7228);
and U19383 (N_19383,N_1520,N_4952);
xor U19384 (N_19384,N_299,N_7814);
nor U19385 (N_19385,N_6896,N_7798);
or U19386 (N_19386,N_7462,N_2462);
nand U19387 (N_19387,N_6156,N_8164);
xor U19388 (N_19388,N_7002,N_3432);
or U19389 (N_19389,N_9538,N_8242);
or U19390 (N_19390,N_1034,N_4443);
nor U19391 (N_19391,N_1852,N_3368);
nor U19392 (N_19392,N_8346,N_6943);
and U19393 (N_19393,N_7166,N_5774);
or U19394 (N_19394,N_1744,N_271);
or U19395 (N_19395,N_4703,N_2760);
nand U19396 (N_19396,N_1531,N_9365);
or U19397 (N_19397,N_2834,N_3070);
or U19398 (N_19398,N_3866,N_3294);
or U19399 (N_19399,N_9620,N_8442);
or U19400 (N_19400,N_3913,N_1915);
nand U19401 (N_19401,N_5566,N_2230);
nor U19402 (N_19402,N_2610,N_160);
nor U19403 (N_19403,N_2368,N_4741);
and U19404 (N_19404,N_8226,N_8986);
nand U19405 (N_19405,N_7297,N_7239);
nand U19406 (N_19406,N_8288,N_9751);
nand U19407 (N_19407,N_4969,N_419);
nand U19408 (N_19408,N_8347,N_7143);
or U19409 (N_19409,N_4846,N_5287);
nand U19410 (N_19410,N_4379,N_5492);
xnor U19411 (N_19411,N_8388,N_7561);
or U19412 (N_19412,N_2726,N_7019);
and U19413 (N_19413,N_3,N_8776);
xnor U19414 (N_19414,N_1324,N_3636);
nor U19415 (N_19415,N_1562,N_990);
or U19416 (N_19416,N_4720,N_4333);
and U19417 (N_19417,N_645,N_9449);
and U19418 (N_19418,N_4088,N_6081);
or U19419 (N_19419,N_8534,N_9847);
xor U19420 (N_19420,N_7221,N_3022);
nand U19421 (N_19421,N_2059,N_2152);
nor U19422 (N_19422,N_900,N_3864);
xnor U19423 (N_19423,N_5481,N_7991);
nand U19424 (N_19424,N_2013,N_8469);
nor U19425 (N_19425,N_1953,N_1187);
and U19426 (N_19426,N_8918,N_8160);
or U19427 (N_19427,N_1684,N_11);
xnor U19428 (N_19428,N_2228,N_4959);
xnor U19429 (N_19429,N_9715,N_854);
nand U19430 (N_19430,N_7644,N_6815);
nor U19431 (N_19431,N_8362,N_7383);
or U19432 (N_19432,N_3116,N_4482);
or U19433 (N_19433,N_2441,N_1248);
and U19434 (N_19434,N_8679,N_7642);
and U19435 (N_19435,N_1969,N_607);
nand U19436 (N_19436,N_5221,N_2961);
xnor U19437 (N_19437,N_6861,N_1232);
nor U19438 (N_19438,N_6669,N_5036);
and U19439 (N_19439,N_3216,N_2877);
and U19440 (N_19440,N_6751,N_5397);
nor U19441 (N_19441,N_523,N_6709);
nor U19442 (N_19442,N_6822,N_5630);
and U19443 (N_19443,N_1542,N_4321);
and U19444 (N_19444,N_3862,N_3809);
nand U19445 (N_19445,N_8696,N_8526);
xnor U19446 (N_19446,N_6874,N_4441);
and U19447 (N_19447,N_426,N_862);
or U19448 (N_19448,N_6549,N_1630);
or U19449 (N_19449,N_2630,N_5491);
xnor U19450 (N_19450,N_843,N_3027);
nand U19451 (N_19451,N_876,N_7441);
nor U19452 (N_19452,N_3980,N_5392);
or U19453 (N_19453,N_756,N_819);
nand U19454 (N_19454,N_3397,N_2972);
nor U19455 (N_19455,N_7455,N_6574);
and U19456 (N_19456,N_1635,N_1835);
xor U19457 (N_19457,N_7736,N_8568);
or U19458 (N_19458,N_4584,N_9767);
and U19459 (N_19459,N_6516,N_6054);
nor U19460 (N_19460,N_4170,N_3622);
nor U19461 (N_19461,N_3092,N_2177);
or U19462 (N_19462,N_1880,N_6167);
or U19463 (N_19463,N_7746,N_6310);
or U19464 (N_19464,N_9451,N_317);
and U19465 (N_19465,N_4492,N_3571);
nor U19466 (N_19466,N_4978,N_5203);
xor U19467 (N_19467,N_3905,N_6505);
nor U19468 (N_19468,N_6206,N_2018);
and U19469 (N_19469,N_6394,N_4675);
xnor U19470 (N_19470,N_7316,N_2717);
and U19471 (N_19471,N_2493,N_8310);
nand U19472 (N_19472,N_5250,N_9887);
and U19473 (N_19473,N_7019,N_2587);
xnor U19474 (N_19474,N_114,N_8141);
or U19475 (N_19475,N_3137,N_5488);
nand U19476 (N_19476,N_8483,N_7139);
xor U19477 (N_19477,N_6986,N_1497);
or U19478 (N_19478,N_2660,N_3130);
xnor U19479 (N_19479,N_1182,N_8604);
and U19480 (N_19480,N_4924,N_2984);
or U19481 (N_19481,N_3907,N_6840);
or U19482 (N_19482,N_8253,N_4985);
nand U19483 (N_19483,N_7724,N_8862);
or U19484 (N_19484,N_6762,N_7000);
and U19485 (N_19485,N_1884,N_7518);
nor U19486 (N_19486,N_9070,N_9781);
and U19487 (N_19487,N_1540,N_5353);
nand U19488 (N_19488,N_6726,N_9444);
or U19489 (N_19489,N_9714,N_3890);
xor U19490 (N_19490,N_3924,N_5164);
nor U19491 (N_19491,N_3238,N_3078);
nand U19492 (N_19492,N_3772,N_3934);
or U19493 (N_19493,N_7037,N_1515);
nor U19494 (N_19494,N_4643,N_2058);
or U19495 (N_19495,N_1563,N_5014);
nor U19496 (N_19496,N_5654,N_7150);
or U19497 (N_19497,N_7327,N_3477);
nor U19498 (N_19498,N_8261,N_1364);
nand U19499 (N_19499,N_5546,N_7326);
or U19500 (N_19500,N_6202,N_892);
nor U19501 (N_19501,N_6006,N_7265);
and U19502 (N_19502,N_7420,N_3632);
nor U19503 (N_19503,N_4483,N_4666);
nor U19504 (N_19504,N_236,N_259);
nand U19505 (N_19505,N_2085,N_8132);
or U19506 (N_19506,N_9164,N_9925);
nand U19507 (N_19507,N_3921,N_8256);
and U19508 (N_19508,N_4580,N_1506);
nand U19509 (N_19509,N_1733,N_674);
xor U19510 (N_19510,N_8394,N_5755);
nor U19511 (N_19511,N_8257,N_8244);
xor U19512 (N_19512,N_9570,N_7983);
nor U19513 (N_19513,N_4864,N_7505);
nor U19514 (N_19514,N_79,N_4110);
nor U19515 (N_19515,N_7068,N_7377);
or U19516 (N_19516,N_5503,N_6870);
or U19517 (N_19517,N_8878,N_2181);
nor U19518 (N_19518,N_2692,N_9644);
nor U19519 (N_19519,N_5178,N_1996);
nand U19520 (N_19520,N_3119,N_3722);
xnor U19521 (N_19521,N_9823,N_2607);
nor U19522 (N_19522,N_3493,N_4285);
xor U19523 (N_19523,N_7401,N_7469);
or U19524 (N_19524,N_2857,N_6315);
xor U19525 (N_19525,N_1858,N_481);
and U19526 (N_19526,N_380,N_7285);
and U19527 (N_19527,N_3844,N_5995);
nor U19528 (N_19528,N_8821,N_9486);
and U19529 (N_19529,N_4821,N_5854);
and U19530 (N_19530,N_1123,N_6944);
and U19531 (N_19531,N_3026,N_674);
xor U19532 (N_19532,N_7151,N_6570);
xnor U19533 (N_19533,N_889,N_8945);
and U19534 (N_19534,N_955,N_8015);
nand U19535 (N_19535,N_2030,N_7873);
nor U19536 (N_19536,N_8549,N_1122);
nor U19537 (N_19537,N_8400,N_899);
nor U19538 (N_19538,N_1258,N_9792);
xnor U19539 (N_19539,N_7792,N_6894);
nor U19540 (N_19540,N_3002,N_9745);
nand U19541 (N_19541,N_8867,N_1159);
nand U19542 (N_19542,N_7357,N_287);
xor U19543 (N_19543,N_3672,N_330);
xnor U19544 (N_19544,N_6212,N_4696);
nand U19545 (N_19545,N_9958,N_1864);
nand U19546 (N_19546,N_4333,N_6913);
and U19547 (N_19547,N_5907,N_1297);
or U19548 (N_19548,N_5006,N_7486);
or U19549 (N_19549,N_8781,N_7553);
or U19550 (N_19550,N_1861,N_9215);
or U19551 (N_19551,N_9115,N_2458);
nor U19552 (N_19552,N_607,N_172);
or U19553 (N_19553,N_6538,N_3659);
and U19554 (N_19554,N_4172,N_5459);
xor U19555 (N_19555,N_6215,N_6021);
xor U19556 (N_19556,N_6886,N_2485);
nor U19557 (N_19557,N_486,N_708);
and U19558 (N_19558,N_6112,N_4329);
xor U19559 (N_19559,N_4762,N_3054);
nand U19560 (N_19560,N_6260,N_9108);
nand U19561 (N_19561,N_1987,N_7232);
xor U19562 (N_19562,N_342,N_9311);
nor U19563 (N_19563,N_9097,N_4192);
or U19564 (N_19564,N_6995,N_4599);
xor U19565 (N_19565,N_2344,N_626);
nand U19566 (N_19566,N_2428,N_6727);
xnor U19567 (N_19567,N_7146,N_7987);
xor U19568 (N_19568,N_7207,N_4143);
and U19569 (N_19569,N_4954,N_3507);
xor U19570 (N_19570,N_1237,N_9079);
and U19571 (N_19571,N_9291,N_2180);
xnor U19572 (N_19572,N_3049,N_7457);
or U19573 (N_19573,N_6324,N_6424);
nor U19574 (N_19574,N_2749,N_9390);
nand U19575 (N_19575,N_5516,N_6219);
nand U19576 (N_19576,N_2232,N_3548);
and U19577 (N_19577,N_571,N_8222);
and U19578 (N_19578,N_1592,N_7682);
xnor U19579 (N_19579,N_3121,N_4003);
nand U19580 (N_19580,N_1916,N_5546);
and U19581 (N_19581,N_3717,N_174);
xnor U19582 (N_19582,N_6312,N_7641);
and U19583 (N_19583,N_8059,N_1684);
xnor U19584 (N_19584,N_3356,N_3203);
nor U19585 (N_19585,N_6534,N_9635);
nor U19586 (N_19586,N_8510,N_7908);
and U19587 (N_19587,N_9522,N_2718);
and U19588 (N_19588,N_9240,N_2115);
nor U19589 (N_19589,N_663,N_3139);
and U19590 (N_19590,N_4447,N_4016);
xnor U19591 (N_19591,N_6036,N_6348);
and U19592 (N_19592,N_304,N_8629);
and U19593 (N_19593,N_9637,N_9042);
nor U19594 (N_19594,N_1033,N_6254);
nand U19595 (N_19595,N_7547,N_8759);
nand U19596 (N_19596,N_8088,N_3861);
nor U19597 (N_19597,N_278,N_2443);
or U19598 (N_19598,N_8337,N_1632);
nor U19599 (N_19599,N_1052,N_7969);
nand U19600 (N_19600,N_9562,N_3490);
nand U19601 (N_19601,N_2182,N_5578);
and U19602 (N_19602,N_7460,N_6946);
and U19603 (N_19603,N_3047,N_8901);
nand U19604 (N_19604,N_6002,N_2883);
or U19605 (N_19605,N_4906,N_7978);
nand U19606 (N_19606,N_5393,N_7684);
and U19607 (N_19607,N_8795,N_2152);
xnor U19608 (N_19608,N_973,N_4519);
nor U19609 (N_19609,N_5213,N_9246);
or U19610 (N_19610,N_3042,N_313);
and U19611 (N_19611,N_7242,N_8931);
nor U19612 (N_19612,N_356,N_4985);
or U19613 (N_19613,N_3507,N_897);
and U19614 (N_19614,N_6627,N_9663);
nor U19615 (N_19615,N_4692,N_2650);
nand U19616 (N_19616,N_7055,N_6143);
and U19617 (N_19617,N_8604,N_1012);
nand U19618 (N_19618,N_2758,N_4121);
nor U19619 (N_19619,N_40,N_6640);
nor U19620 (N_19620,N_5644,N_2741);
nor U19621 (N_19621,N_9147,N_8336);
and U19622 (N_19622,N_5294,N_1500);
or U19623 (N_19623,N_98,N_4287);
and U19624 (N_19624,N_5880,N_6110);
nand U19625 (N_19625,N_5898,N_2992);
nor U19626 (N_19626,N_6081,N_5435);
or U19627 (N_19627,N_8908,N_964);
xor U19628 (N_19628,N_7739,N_4842);
nand U19629 (N_19629,N_4550,N_1598);
nor U19630 (N_19630,N_1994,N_4797);
and U19631 (N_19631,N_421,N_3715);
nor U19632 (N_19632,N_438,N_6838);
or U19633 (N_19633,N_1751,N_4328);
xnor U19634 (N_19634,N_4017,N_2747);
nand U19635 (N_19635,N_8576,N_254);
and U19636 (N_19636,N_1782,N_8609);
nand U19637 (N_19637,N_3444,N_3206);
xnor U19638 (N_19638,N_5401,N_2358);
xor U19639 (N_19639,N_7652,N_4842);
nand U19640 (N_19640,N_7922,N_9290);
or U19641 (N_19641,N_5243,N_4829);
or U19642 (N_19642,N_6254,N_1996);
xnor U19643 (N_19643,N_9616,N_2640);
nand U19644 (N_19644,N_9854,N_6624);
or U19645 (N_19645,N_5364,N_4085);
nor U19646 (N_19646,N_2157,N_2612);
xnor U19647 (N_19647,N_8998,N_3291);
nand U19648 (N_19648,N_2099,N_1272);
nor U19649 (N_19649,N_5832,N_204);
xnor U19650 (N_19650,N_8958,N_5765);
or U19651 (N_19651,N_7775,N_1315);
and U19652 (N_19652,N_3957,N_4027);
and U19653 (N_19653,N_5565,N_1062);
nor U19654 (N_19654,N_8240,N_7205);
or U19655 (N_19655,N_6415,N_3456);
nor U19656 (N_19656,N_7648,N_5735);
or U19657 (N_19657,N_1594,N_3530);
nand U19658 (N_19658,N_7009,N_8532);
xnor U19659 (N_19659,N_8807,N_5265);
nor U19660 (N_19660,N_6198,N_4854);
and U19661 (N_19661,N_1528,N_6470);
nand U19662 (N_19662,N_6580,N_4416);
xor U19663 (N_19663,N_3943,N_9586);
nor U19664 (N_19664,N_8791,N_8686);
nor U19665 (N_19665,N_3351,N_8472);
nor U19666 (N_19666,N_4129,N_5900);
or U19667 (N_19667,N_1824,N_9976);
xor U19668 (N_19668,N_778,N_5474);
or U19669 (N_19669,N_2884,N_1302);
xnor U19670 (N_19670,N_3825,N_2079);
or U19671 (N_19671,N_3155,N_2855);
nand U19672 (N_19672,N_3771,N_3136);
and U19673 (N_19673,N_7682,N_7192);
nand U19674 (N_19674,N_4351,N_2502);
xnor U19675 (N_19675,N_8158,N_9857);
nand U19676 (N_19676,N_3357,N_7);
and U19677 (N_19677,N_4780,N_1768);
and U19678 (N_19678,N_7244,N_4446);
and U19679 (N_19679,N_477,N_1463);
or U19680 (N_19680,N_9754,N_103);
xnor U19681 (N_19681,N_1518,N_5573);
or U19682 (N_19682,N_3888,N_4504);
nor U19683 (N_19683,N_6849,N_2332);
nor U19684 (N_19684,N_4953,N_5231);
and U19685 (N_19685,N_1257,N_8594);
xor U19686 (N_19686,N_7222,N_245);
nand U19687 (N_19687,N_2880,N_1830);
or U19688 (N_19688,N_4165,N_6808);
or U19689 (N_19689,N_7146,N_9508);
xnor U19690 (N_19690,N_7855,N_1025);
nand U19691 (N_19691,N_9642,N_7123);
nor U19692 (N_19692,N_4602,N_9184);
nand U19693 (N_19693,N_7567,N_5864);
nand U19694 (N_19694,N_3444,N_7932);
nor U19695 (N_19695,N_578,N_3585);
and U19696 (N_19696,N_2379,N_6999);
or U19697 (N_19697,N_1596,N_2413);
nor U19698 (N_19698,N_1472,N_3219);
or U19699 (N_19699,N_2682,N_6030);
or U19700 (N_19700,N_5473,N_9466);
nor U19701 (N_19701,N_3348,N_8996);
and U19702 (N_19702,N_3540,N_133);
nand U19703 (N_19703,N_7955,N_2044);
nor U19704 (N_19704,N_4400,N_8400);
nor U19705 (N_19705,N_6668,N_1695);
nand U19706 (N_19706,N_7079,N_2726);
or U19707 (N_19707,N_2477,N_6797);
or U19708 (N_19708,N_2114,N_5252);
nor U19709 (N_19709,N_7704,N_6648);
and U19710 (N_19710,N_3972,N_403);
or U19711 (N_19711,N_9240,N_934);
nand U19712 (N_19712,N_4157,N_5743);
xor U19713 (N_19713,N_7861,N_805);
nand U19714 (N_19714,N_7190,N_3035);
xor U19715 (N_19715,N_9414,N_2769);
or U19716 (N_19716,N_7673,N_4330);
or U19717 (N_19717,N_7581,N_5573);
nor U19718 (N_19718,N_5490,N_3387);
nor U19719 (N_19719,N_7389,N_3447);
and U19720 (N_19720,N_2124,N_887);
xnor U19721 (N_19721,N_7693,N_9164);
and U19722 (N_19722,N_7979,N_6498);
or U19723 (N_19723,N_3306,N_9686);
nand U19724 (N_19724,N_1682,N_4578);
xnor U19725 (N_19725,N_3329,N_5422);
nand U19726 (N_19726,N_1778,N_6806);
and U19727 (N_19727,N_578,N_8248);
nor U19728 (N_19728,N_1134,N_377);
nand U19729 (N_19729,N_3354,N_4360);
nor U19730 (N_19730,N_8716,N_3363);
xnor U19731 (N_19731,N_6397,N_2779);
nand U19732 (N_19732,N_8635,N_7993);
nand U19733 (N_19733,N_569,N_6875);
and U19734 (N_19734,N_8894,N_4061);
nand U19735 (N_19735,N_8528,N_8857);
nor U19736 (N_19736,N_2255,N_8561);
nor U19737 (N_19737,N_7712,N_207);
and U19738 (N_19738,N_1923,N_3736);
and U19739 (N_19739,N_2155,N_4603);
xor U19740 (N_19740,N_5684,N_9529);
or U19741 (N_19741,N_920,N_3559);
nand U19742 (N_19742,N_5862,N_4696);
xnor U19743 (N_19743,N_6538,N_2986);
or U19744 (N_19744,N_1132,N_5181);
xnor U19745 (N_19745,N_9442,N_4044);
nor U19746 (N_19746,N_2004,N_3367);
and U19747 (N_19747,N_4252,N_1115);
and U19748 (N_19748,N_7640,N_2047);
and U19749 (N_19749,N_8015,N_9890);
xnor U19750 (N_19750,N_3392,N_6482);
and U19751 (N_19751,N_1182,N_3283);
and U19752 (N_19752,N_1644,N_2603);
and U19753 (N_19753,N_8788,N_8757);
nor U19754 (N_19754,N_4096,N_1850);
or U19755 (N_19755,N_655,N_3234);
or U19756 (N_19756,N_2802,N_6455);
or U19757 (N_19757,N_8063,N_9668);
nor U19758 (N_19758,N_983,N_309);
and U19759 (N_19759,N_2789,N_2529);
nand U19760 (N_19760,N_3303,N_2512);
and U19761 (N_19761,N_8094,N_3073);
nand U19762 (N_19762,N_4347,N_8549);
xor U19763 (N_19763,N_4119,N_2485);
xor U19764 (N_19764,N_8431,N_152);
nor U19765 (N_19765,N_7375,N_5572);
xor U19766 (N_19766,N_8803,N_3147);
nand U19767 (N_19767,N_5218,N_3159);
nor U19768 (N_19768,N_6507,N_7782);
nor U19769 (N_19769,N_6325,N_4961);
and U19770 (N_19770,N_1496,N_9404);
and U19771 (N_19771,N_7700,N_8114);
or U19772 (N_19772,N_2054,N_6089);
or U19773 (N_19773,N_7692,N_8601);
nor U19774 (N_19774,N_5682,N_567);
nand U19775 (N_19775,N_8151,N_3696);
and U19776 (N_19776,N_8179,N_4596);
and U19777 (N_19777,N_2058,N_1460);
nor U19778 (N_19778,N_6170,N_774);
nand U19779 (N_19779,N_8051,N_2196);
nand U19780 (N_19780,N_2616,N_1036);
and U19781 (N_19781,N_1318,N_8845);
nor U19782 (N_19782,N_4253,N_4928);
or U19783 (N_19783,N_5272,N_6796);
xnor U19784 (N_19784,N_4458,N_4676);
and U19785 (N_19785,N_9974,N_7382);
xor U19786 (N_19786,N_1078,N_3829);
nor U19787 (N_19787,N_5242,N_2161);
nand U19788 (N_19788,N_7839,N_3984);
nor U19789 (N_19789,N_4966,N_9806);
nor U19790 (N_19790,N_7384,N_4845);
nand U19791 (N_19791,N_9761,N_7517);
xnor U19792 (N_19792,N_7295,N_9303);
nand U19793 (N_19793,N_4140,N_6255);
xor U19794 (N_19794,N_7567,N_531);
nand U19795 (N_19795,N_3964,N_8157);
or U19796 (N_19796,N_4193,N_8461);
and U19797 (N_19797,N_4411,N_1265);
and U19798 (N_19798,N_5473,N_9599);
nor U19799 (N_19799,N_9839,N_5905);
and U19800 (N_19800,N_1178,N_9815);
and U19801 (N_19801,N_7261,N_9228);
and U19802 (N_19802,N_6749,N_2964);
or U19803 (N_19803,N_6310,N_3496);
or U19804 (N_19804,N_3878,N_7109);
xor U19805 (N_19805,N_8945,N_2913);
or U19806 (N_19806,N_3410,N_9216);
and U19807 (N_19807,N_4187,N_3222);
nor U19808 (N_19808,N_261,N_256);
and U19809 (N_19809,N_6232,N_2181);
xnor U19810 (N_19810,N_8905,N_6261);
xnor U19811 (N_19811,N_2808,N_8388);
or U19812 (N_19812,N_6008,N_8636);
and U19813 (N_19813,N_9585,N_3226);
nand U19814 (N_19814,N_4288,N_6886);
nor U19815 (N_19815,N_1266,N_6961);
nand U19816 (N_19816,N_7913,N_369);
nand U19817 (N_19817,N_2045,N_1084);
xnor U19818 (N_19818,N_4970,N_3134);
and U19819 (N_19819,N_4132,N_8370);
nor U19820 (N_19820,N_2767,N_3218);
nor U19821 (N_19821,N_1757,N_1906);
and U19822 (N_19822,N_1686,N_6080);
xnor U19823 (N_19823,N_1624,N_4920);
and U19824 (N_19824,N_1140,N_6624);
or U19825 (N_19825,N_1101,N_1402);
and U19826 (N_19826,N_7203,N_6232);
or U19827 (N_19827,N_1012,N_8209);
nand U19828 (N_19828,N_3551,N_3840);
or U19829 (N_19829,N_2761,N_2520);
nand U19830 (N_19830,N_3388,N_2354);
nor U19831 (N_19831,N_8814,N_4643);
or U19832 (N_19832,N_6129,N_8578);
xor U19833 (N_19833,N_5442,N_4449);
nor U19834 (N_19834,N_4049,N_4188);
nor U19835 (N_19835,N_150,N_1792);
nor U19836 (N_19836,N_7168,N_1221);
nor U19837 (N_19837,N_9692,N_9340);
nand U19838 (N_19838,N_8810,N_7779);
xor U19839 (N_19839,N_7817,N_758);
nor U19840 (N_19840,N_7956,N_5157);
and U19841 (N_19841,N_6659,N_4057);
nand U19842 (N_19842,N_4059,N_8637);
and U19843 (N_19843,N_3335,N_4572);
or U19844 (N_19844,N_1426,N_1806);
nor U19845 (N_19845,N_765,N_9133);
nand U19846 (N_19846,N_8983,N_5968);
or U19847 (N_19847,N_2574,N_686);
xor U19848 (N_19848,N_982,N_3864);
nor U19849 (N_19849,N_4302,N_3235);
and U19850 (N_19850,N_8596,N_8924);
nor U19851 (N_19851,N_383,N_577);
nor U19852 (N_19852,N_6894,N_7601);
xnor U19853 (N_19853,N_1144,N_9136);
or U19854 (N_19854,N_9481,N_8060);
nand U19855 (N_19855,N_8514,N_9688);
xor U19856 (N_19856,N_4326,N_1865);
nand U19857 (N_19857,N_14,N_4584);
xor U19858 (N_19858,N_5174,N_3944);
nor U19859 (N_19859,N_5282,N_1525);
xor U19860 (N_19860,N_2639,N_2878);
or U19861 (N_19861,N_4433,N_1038);
nor U19862 (N_19862,N_2466,N_6264);
nor U19863 (N_19863,N_7791,N_9011);
nor U19864 (N_19864,N_7787,N_2199);
nor U19865 (N_19865,N_8199,N_213);
nand U19866 (N_19866,N_9669,N_2262);
nand U19867 (N_19867,N_267,N_6503);
nand U19868 (N_19868,N_1390,N_4276);
and U19869 (N_19869,N_9081,N_6086);
nand U19870 (N_19870,N_1932,N_3780);
nand U19871 (N_19871,N_7613,N_1819);
nand U19872 (N_19872,N_2004,N_2984);
or U19873 (N_19873,N_1498,N_647);
and U19874 (N_19874,N_4231,N_4253);
xor U19875 (N_19875,N_8966,N_3104);
nor U19876 (N_19876,N_1139,N_1171);
nor U19877 (N_19877,N_9187,N_7919);
nand U19878 (N_19878,N_4191,N_4550);
nor U19879 (N_19879,N_5498,N_4561);
xnor U19880 (N_19880,N_3056,N_5593);
nor U19881 (N_19881,N_7260,N_1385);
nor U19882 (N_19882,N_1475,N_5449);
or U19883 (N_19883,N_8150,N_221);
and U19884 (N_19884,N_3335,N_4757);
xor U19885 (N_19885,N_8630,N_1646);
xnor U19886 (N_19886,N_1915,N_1933);
and U19887 (N_19887,N_8660,N_10);
and U19888 (N_19888,N_6463,N_4699);
and U19889 (N_19889,N_3821,N_4894);
xnor U19890 (N_19890,N_9135,N_9892);
xnor U19891 (N_19891,N_470,N_5967);
and U19892 (N_19892,N_6928,N_3025);
nor U19893 (N_19893,N_5000,N_5099);
or U19894 (N_19894,N_3003,N_6407);
and U19895 (N_19895,N_4114,N_8595);
nor U19896 (N_19896,N_2282,N_3132);
or U19897 (N_19897,N_5322,N_4010);
and U19898 (N_19898,N_921,N_7255);
nor U19899 (N_19899,N_2875,N_7513);
nand U19900 (N_19900,N_9347,N_470);
or U19901 (N_19901,N_296,N_523);
nor U19902 (N_19902,N_5978,N_9303);
or U19903 (N_19903,N_1353,N_3662);
or U19904 (N_19904,N_8982,N_5093);
nand U19905 (N_19905,N_929,N_1163);
nand U19906 (N_19906,N_6875,N_4683);
and U19907 (N_19907,N_1842,N_8953);
xnor U19908 (N_19908,N_4617,N_4877);
nor U19909 (N_19909,N_1707,N_5349);
nand U19910 (N_19910,N_7380,N_4114);
nor U19911 (N_19911,N_3989,N_3416);
xnor U19912 (N_19912,N_3364,N_8114);
or U19913 (N_19913,N_2410,N_7626);
xnor U19914 (N_19914,N_6209,N_8915);
or U19915 (N_19915,N_3608,N_3547);
nand U19916 (N_19916,N_6236,N_6144);
xnor U19917 (N_19917,N_3516,N_7434);
xnor U19918 (N_19918,N_5270,N_111);
or U19919 (N_19919,N_9553,N_4133);
and U19920 (N_19920,N_459,N_2624);
nand U19921 (N_19921,N_8970,N_4471);
and U19922 (N_19922,N_9607,N_2799);
nor U19923 (N_19923,N_6330,N_968);
and U19924 (N_19924,N_6672,N_4517);
or U19925 (N_19925,N_7404,N_7152);
xor U19926 (N_19926,N_1827,N_1133);
nor U19927 (N_19927,N_4283,N_5908);
or U19928 (N_19928,N_8079,N_7342);
xnor U19929 (N_19929,N_7136,N_9030);
and U19930 (N_19930,N_9786,N_2744);
and U19931 (N_19931,N_981,N_7305);
nand U19932 (N_19932,N_9303,N_7066);
nor U19933 (N_19933,N_2042,N_9614);
nor U19934 (N_19934,N_400,N_6831);
and U19935 (N_19935,N_5101,N_6921);
xnor U19936 (N_19936,N_115,N_7885);
nor U19937 (N_19937,N_8529,N_3898);
or U19938 (N_19938,N_2937,N_3003);
xnor U19939 (N_19939,N_8625,N_7339);
and U19940 (N_19940,N_991,N_5422);
or U19941 (N_19941,N_5734,N_6834);
or U19942 (N_19942,N_8027,N_9657);
or U19943 (N_19943,N_7288,N_9834);
or U19944 (N_19944,N_7101,N_4952);
nand U19945 (N_19945,N_3484,N_2023);
or U19946 (N_19946,N_3751,N_7439);
nand U19947 (N_19947,N_197,N_8110);
or U19948 (N_19948,N_3214,N_3741);
xor U19949 (N_19949,N_7192,N_4281);
and U19950 (N_19950,N_4168,N_4838);
nor U19951 (N_19951,N_9312,N_390);
nor U19952 (N_19952,N_7199,N_3823);
or U19953 (N_19953,N_9525,N_913);
and U19954 (N_19954,N_5663,N_101);
xor U19955 (N_19955,N_1272,N_4844);
nand U19956 (N_19956,N_2340,N_5316);
or U19957 (N_19957,N_5371,N_4052);
or U19958 (N_19958,N_6849,N_9862);
and U19959 (N_19959,N_1100,N_664);
nor U19960 (N_19960,N_7696,N_4338);
xor U19961 (N_19961,N_668,N_8020);
nand U19962 (N_19962,N_3193,N_3550);
or U19963 (N_19963,N_3607,N_248);
xor U19964 (N_19964,N_7878,N_3146);
or U19965 (N_19965,N_8304,N_8360);
and U19966 (N_19966,N_5157,N_5844);
nor U19967 (N_19967,N_1366,N_1064);
or U19968 (N_19968,N_1189,N_4559);
and U19969 (N_19969,N_3112,N_9644);
nor U19970 (N_19970,N_8149,N_8184);
xor U19971 (N_19971,N_2945,N_2529);
nand U19972 (N_19972,N_2365,N_2075);
or U19973 (N_19973,N_8703,N_5907);
xnor U19974 (N_19974,N_9821,N_1794);
and U19975 (N_19975,N_947,N_7530);
nand U19976 (N_19976,N_1754,N_9302);
or U19977 (N_19977,N_499,N_2131);
nor U19978 (N_19978,N_1300,N_2678);
nand U19979 (N_19979,N_1579,N_6422);
nand U19980 (N_19980,N_2768,N_658);
nor U19981 (N_19981,N_3253,N_6708);
nand U19982 (N_19982,N_7355,N_6165);
xor U19983 (N_19983,N_4636,N_580);
nor U19984 (N_19984,N_6786,N_7859);
and U19985 (N_19985,N_1912,N_6789);
nor U19986 (N_19986,N_4055,N_4097);
nor U19987 (N_19987,N_2402,N_6663);
and U19988 (N_19988,N_5148,N_1075);
xnor U19989 (N_19989,N_8028,N_8849);
nand U19990 (N_19990,N_5177,N_9985);
nor U19991 (N_19991,N_1007,N_826);
xor U19992 (N_19992,N_3730,N_3342);
nor U19993 (N_19993,N_2759,N_8746);
and U19994 (N_19994,N_1090,N_4312);
nand U19995 (N_19995,N_6339,N_9579);
xnor U19996 (N_19996,N_8299,N_3147);
xnor U19997 (N_19997,N_2682,N_808);
xnor U19998 (N_19998,N_6443,N_3701);
xnor U19999 (N_19999,N_8219,N_1207);
nor U20000 (N_20000,N_12912,N_19103);
nand U20001 (N_20001,N_12863,N_17641);
nand U20002 (N_20002,N_15321,N_10572);
xnor U20003 (N_20003,N_14517,N_18540);
or U20004 (N_20004,N_12768,N_17744);
nor U20005 (N_20005,N_17704,N_19953);
and U20006 (N_20006,N_12356,N_11772);
nand U20007 (N_20007,N_14461,N_18528);
and U20008 (N_20008,N_13997,N_17855);
xor U20009 (N_20009,N_17954,N_16998);
xor U20010 (N_20010,N_12093,N_17723);
xor U20011 (N_20011,N_17837,N_19063);
or U20012 (N_20012,N_13597,N_12224);
and U20013 (N_20013,N_14082,N_16178);
or U20014 (N_20014,N_19044,N_14122);
nand U20015 (N_20015,N_12850,N_18767);
nand U20016 (N_20016,N_10600,N_18958);
nor U20017 (N_20017,N_16177,N_10459);
nor U20018 (N_20018,N_13319,N_17212);
xnor U20019 (N_20019,N_17351,N_12019);
xor U20020 (N_20020,N_13940,N_10068);
or U20021 (N_20021,N_17294,N_17273);
nor U20022 (N_20022,N_17213,N_16215);
xnor U20023 (N_20023,N_18274,N_13698);
nand U20024 (N_20024,N_18246,N_12115);
and U20025 (N_20025,N_18896,N_17722);
nand U20026 (N_20026,N_19586,N_18974);
or U20027 (N_20027,N_14588,N_13638);
nor U20028 (N_20028,N_10039,N_13274);
nor U20029 (N_20029,N_13607,N_13441);
xnor U20030 (N_20030,N_18521,N_15017);
nand U20031 (N_20031,N_16159,N_17946);
and U20032 (N_20032,N_14397,N_17112);
or U20033 (N_20033,N_12540,N_19424);
nand U20034 (N_20034,N_12967,N_16446);
xor U20035 (N_20035,N_11408,N_19880);
and U20036 (N_20036,N_11714,N_16133);
xor U20037 (N_20037,N_19995,N_15804);
nor U20038 (N_20038,N_16008,N_15090);
or U20039 (N_20039,N_14556,N_16200);
nor U20040 (N_20040,N_16412,N_13081);
xor U20041 (N_20041,N_15224,N_18456);
xor U20042 (N_20042,N_13007,N_15218);
xnor U20043 (N_20043,N_17842,N_14733);
or U20044 (N_20044,N_16598,N_10843);
nand U20045 (N_20045,N_14958,N_18082);
and U20046 (N_20046,N_10938,N_10974);
or U20047 (N_20047,N_18720,N_19136);
and U20048 (N_20048,N_17795,N_18865);
or U20049 (N_20049,N_13505,N_10747);
and U20050 (N_20050,N_18480,N_10520);
and U20051 (N_20051,N_12926,N_16898);
or U20052 (N_20052,N_13006,N_12068);
nor U20053 (N_20053,N_11810,N_17793);
nand U20054 (N_20054,N_13067,N_16881);
or U20055 (N_20055,N_10597,N_14329);
nor U20056 (N_20056,N_12997,N_19121);
nand U20057 (N_20057,N_10013,N_15523);
xnor U20058 (N_20058,N_12092,N_10909);
and U20059 (N_20059,N_12897,N_17084);
nand U20060 (N_20060,N_12188,N_18931);
or U20061 (N_20061,N_11948,N_13381);
nand U20062 (N_20062,N_17824,N_14219);
or U20063 (N_20063,N_11271,N_14090);
xor U20064 (N_20064,N_16643,N_19758);
nor U20065 (N_20065,N_16730,N_17968);
nand U20066 (N_20066,N_19976,N_19876);
nand U20067 (N_20067,N_17166,N_10614);
nor U20068 (N_20068,N_12659,N_12719);
or U20069 (N_20069,N_11041,N_13909);
nand U20070 (N_20070,N_15262,N_10246);
and U20071 (N_20071,N_16115,N_10823);
nor U20072 (N_20072,N_15293,N_19352);
and U20073 (N_20073,N_13825,N_13741);
xor U20074 (N_20074,N_13804,N_18384);
nor U20075 (N_20075,N_13429,N_12037);
xnor U20076 (N_20076,N_13697,N_19440);
xnor U20077 (N_20077,N_11795,N_13922);
nor U20078 (N_20078,N_11124,N_15171);
nand U20079 (N_20079,N_13417,N_15306);
nor U20080 (N_20080,N_14632,N_18415);
nand U20081 (N_20081,N_17511,N_14077);
xnor U20082 (N_20082,N_16719,N_15598);
xnor U20083 (N_20083,N_11823,N_11179);
xnor U20084 (N_20084,N_15436,N_15081);
nand U20085 (N_20085,N_12461,N_18696);
nand U20086 (N_20086,N_18833,N_12463);
nor U20087 (N_20087,N_13608,N_10899);
xor U20088 (N_20088,N_13211,N_10643);
nor U20089 (N_20089,N_16246,N_16423);
xor U20090 (N_20090,N_19992,N_13742);
or U20091 (N_20091,N_13084,N_14466);
or U20092 (N_20092,N_14773,N_13595);
nand U20093 (N_20093,N_18190,N_19579);
xnor U20094 (N_20094,N_18580,N_14023);
xor U20095 (N_20095,N_16531,N_11218);
nand U20096 (N_20096,N_16541,N_11157);
nand U20097 (N_20097,N_18038,N_10963);
xnor U20098 (N_20098,N_19004,N_15391);
nor U20099 (N_20099,N_18033,N_19200);
nand U20100 (N_20100,N_16289,N_17204);
xnor U20101 (N_20101,N_15876,N_16092);
and U20102 (N_20102,N_16997,N_19653);
or U20103 (N_20103,N_14797,N_17733);
or U20104 (N_20104,N_19080,N_10168);
nor U20105 (N_20105,N_19765,N_14749);
and U20106 (N_20106,N_18137,N_12210);
nor U20107 (N_20107,N_16324,N_13075);
or U20108 (N_20108,N_17767,N_16720);
and U20109 (N_20109,N_10390,N_16611);
and U20110 (N_20110,N_17901,N_19670);
nand U20111 (N_20111,N_11668,N_15476);
and U20112 (N_20112,N_13883,N_17669);
nand U20113 (N_20113,N_14861,N_12052);
nor U20114 (N_20114,N_10344,N_11690);
nor U20115 (N_20115,N_17414,N_19710);
and U20116 (N_20116,N_19861,N_17642);
and U20117 (N_20117,N_13944,N_10975);
xor U20118 (N_20118,N_10099,N_10546);
nor U20119 (N_20119,N_15921,N_14249);
and U20120 (N_20120,N_19607,N_10169);
or U20121 (N_20121,N_17525,N_16050);
and U20122 (N_20122,N_18810,N_14266);
or U20123 (N_20123,N_13532,N_18264);
nor U20124 (N_20124,N_11974,N_10635);
or U20125 (N_20125,N_16606,N_17109);
xnor U20126 (N_20126,N_12699,N_18770);
xor U20127 (N_20127,N_10337,N_19571);
nor U20128 (N_20128,N_13119,N_13017);
and U20129 (N_20129,N_10124,N_16360);
xor U20130 (N_20130,N_12742,N_16853);
nor U20131 (N_20131,N_13030,N_17560);
and U20132 (N_20132,N_11190,N_18866);
or U20133 (N_20133,N_18168,N_13307);
or U20134 (N_20134,N_10134,N_16283);
or U20135 (N_20135,N_13708,N_14086);
xnor U20136 (N_20136,N_14327,N_17776);
nor U20137 (N_20137,N_10454,N_13892);
nor U20138 (N_20138,N_17430,N_18413);
and U20139 (N_20139,N_14566,N_14904);
and U20140 (N_20140,N_10729,N_10019);
nand U20141 (N_20141,N_11490,N_19628);
and U20142 (N_20142,N_11866,N_13513);
or U20143 (N_20143,N_19996,N_14375);
nand U20144 (N_20144,N_17180,N_12415);
nand U20145 (N_20145,N_14172,N_10357);
or U20146 (N_20146,N_16736,N_14347);
nand U20147 (N_20147,N_13263,N_10378);
xnor U20148 (N_20148,N_17222,N_12824);
and U20149 (N_20149,N_19734,N_12515);
nand U20150 (N_20150,N_12158,N_18360);
xnor U20151 (N_20151,N_13982,N_14525);
or U20152 (N_20152,N_19652,N_15108);
or U20153 (N_20153,N_11288,N_19459);
nor U20154 (N_20154,N_12334,N_14010);
nand U20155 (N_20155,N_18562,N_10559);
and U20156 (N_20156,N_11425,N_16439);
and U20157 (N_20157,N_16754,N_14328);
xnor U20158 (N_20158,N_12248,N_11770);
nand U20159 (N_20159,N_17701,N_17115);
xnor U20160 (N_20160,N_17427,N_13252);
xnor U20161 (N_20161,N_18559,N_13719);
nor U20162 (N_20162,N_17546,N_14902);
nand U20163 (N_20163,N_14820,N_15567);
and U20164 (N_20164,N_11878,N_11909);
nand U20165 (N_20165,N_18476,N_10863);
or U20166 (N_20166,N_14317,N_18645);
or U20167 (N_20167,N_19248,N_18475);
nand U20168 (N_20168,N_13853,N_12887);
and U20169 (N_20169,N_18128,N_10319);
or U20170 (N_20170,N_11217,N_11918);
or U20171 (N_20171,N_10308,N_17593);
nand U20172 (N_20172,N_14193,N_19917);
nand U20173 (N_20173,N_18199,N_11361);
and U20174 (N_20174,N_11851,N_12318);
nand U20175 (N_20175,N_16405,N_14918);
xnor U20176 (N_20176,N_13581,N_16681);
xnor U20177 (N_20177,N_11275,N_14721);
nand U20178 (N_20178,N_13079,N_11749);
and U20179 (N_20179,N_14955,N_13677);
nor U20180 (N_20180,N_10623,N_16431);
xnor U20181 (N_20181,N_16395,N_14093);
nand U20182 (N_20182,N_17377,N_18129);
or U20183 (N_20183,N_13822,N_12430);
and U20184 (N_20184,N_13955,N_16271);
and U20185 (N_20185,N_16517,N_19252);
or U20186 (N_20186,N_15770,N_15652);
nor U20187 (N_20187,N_17909,N_10112);
nor U20188 (N_20188,N_10092,N_10640);
and U20189 (N_20189,N_14363,N_12631);
nor U20190 (N_20190,N_16511,N_11906);
nand U20191 (N_20191,N_14159,N_12179);
and U20192 (N_20192,N_14261,N_13561);
nor U20193 (N_20193,N_12593,N_12957);
xor U20194 (N_20194,N_10716,N_11301);
or U20195 (N_20195,N_12447,N_12510);
and U20196 (N_20196,N_17295,N_13460);
and U20197 (N_20197,N_14880,N_19141);
and U20198 (N_20198,N_15382,N_11071);
nand U20199 (N_20199,N_18406,N_18534);
or U20200 (N_20200,N_13947,N_18053);
xnor U20201 (N_20201,N_12520,N_16607);
or U20202 (N_20202,N_16635,N_14735);
nor U20203 (N_20203,N_12145,N_13244);
nand U20204 (N_20204,N_17150,N_18222);
nand U20205 (N_20205,N_12138,N_12012);
xnor U20206 (N_20206,N_10098,N_19193);
and U20207 (N_20207,N_11747,N_14752);
and U20208 (N_20208,N_19598,N_14030);
xor U20209 (N_20209,N_15252,N_12310);
nand U20210 (N_20210,N_14972,N_13515);
nor U20211 (N_20211,N_12893,N_19388);
xnor U20212 (N_20212,N_13098,N_17646);
and U20213 (N_20213,N_16584,N_17743);
nor U20214 (N_20214,N_16655,N_12126);
nand U20215 (N_20215,N_12133,N_10626);
or U20216 (N_20216,N_18189,N_15893);
xor U20217 (N_20217,N_16928,N_17058);
and U20218 (N_20218,N_16729,N_11469);
and U20219 (N_20219,N_14817,N_18817);
and U20220 (N_20220,N_10386,N_19323);
nor U20221 (N_20221,N_17055,N_17029);
nor U20222 (N_20222,N_18322,N_10177);
nor U20223 (N_20223,N_13755,N_13200);
or U20224 (N_20224,N_15905,N_19943);
nand U20225 (N_20225,N_14376,N_12241);
nand U20226 (N_20226,N_18380,N_13525);
and U20227 (N_20227,N_15915,N_12464);
or U20228 (N_20228,N_18683,N_18785);
and U20229 (N_20229,N_14356,N_15590);
nor U20230 (N_20230,N_10430,N_12668);
xnor U20231 (N_20231,N_12419,N_10987);
nand U20232 (N_20232,N_19639,N_14070);
xor U20233 (N_20233,N_17108,N_19254);
nand U20234 (N_20234,N_11415,N_13529);
or U20235 (N_20235,N_14934,N_18088);
xor U20236 (N_20236,N_16612,N_10654);
xnor U20237 (N_20237,N_12835,N_18734);
nand U20238 (N_20238,N_19655,N_17962);
or U20239 (N_20239,N_19946,N_10742);
and U20240 (N_20240,N_10433,N_17667);
xor U20241 (N_20241,N_19854,N_13649);
nand U20242 (N_20242,N_11806,N_11776);
or U20243 (N_20243,N_16514,N_12507);
nand U20244 (N_20244,N_13285,N_14176);
and U20245 (N_20245,N_14806,N_18956);
xnor U20246 (N_20246,N_18546,N_17303);
nor U20247 (N_20247,N_11059,N_14539);
nor U20248 (N_20248,N_14352,N_15377);
and U20249 (N_20249,N_13146,N_10889);
and U20250 (N_20250,N_10170,N_18601);
and U20251 (N_20251,N_17557,N_10836);
xnor U20252 (N_20252,N_17320,N_16544);
nand U20253 (N_20253,N_13855,N_17566);
or U20254 (N_20254,N_14884,N_16308);
nor U20255 (N_20255,N_10289,N_10898);
nor U20256 (N_20256,N_12313,N_19503);
or U20257 (N_20257,N_18486,N_15862);
xnor U20258 (N_20258,N_12658,N_10267);
nand U20259 (N_20259,N_13670,N_11169);
or U20260 (N_20260,N_17556,N_18936);
nand U20261 (N_20261,N_15214,N_15671);
nand U20262 (N_20262,N_11307,N_11409);
nand U20263 (N_20263,N_18541,N_17170);
nand U20264 (N_20264,N_11493,N_14758);
nand U20265 (N_20265,N_16104,N_12116);
or U20266 (N_20266,N_17153,N_10897);
and U20267 (N_20267,N_15107,N_14034);
xnor U20268 (N_20268,N_19206,N_11122);
or U20269 (N_20269,N_10399,N_18115);
nor U20270 (N_20270,N_13207,N_12345);
or U20271 (N_20271,N_13680,N_15731);
nand U20272 (N_20272,N_15228,N_19023);
or U20273 (N_20273,N_11984,N_16817);
nand U20274 (N_20274,N_15756,N_13536);
nand U20275 (N_20275,N_17503,N_14960);
nand U20276 (N_20276,N_19460,N_14672);
nand U20277 (N_20277,N_14544,N_13340);
and U20278 (N_20278,N_19951,N_17355);
nor U20279 (N_20279,N_16233,N_12482);
and U20280 (N_20280,N_15023,N_12605);
nand U20281 (N_20281,N_13629,N_19530);
nor U20282 (N_20282,N_17741,N_14149);
nand U20283 (N_20283,N_12557,N_14547);
nor U20284 (N_20284,N_19894,N_16839);
xnor U20285 (N_20285,N_15376,N_11193);
xnor U20286 (N_20286,N_15557,N_11608);
and U20287 (N_20287,N_18050,N_10095);
or U20288 (N_20288,N_17230,N_13267);
xnor U20289 (N_20289,N_18520,N_15439);
or U20290 (N_20290,N_14342,N_17478);
nor U20291 (N_20291,N_18832,N_17007);
and U20292 (N_20292,N_18165,N_18211);
or U20293 (N_20293,N_17436,N_15982);
or U20294 (N_20294,N_12214,N_10947);
and U20295 (N_20295,N_11802,N_16313);
nand U20296 (N_20296,N_10647,N_17220);
or U20297 (N_20297,N_14741,N_12247);
nor U20298 (N_20298,N_15481,N_19093);
nor U20299 (N_20299,N_15609,N_14118);
nor U20300 (N_20300,N_17886,N_11221);
nand U20301 (N_20301,N_14433,N_10783);
xor U20302 (N_20302,N_12531,N_10787);
xnor U20303 (N_20303,N_19508,N_11173);
and U20304 (N_20304,N_18943,N_18048);
xnor U20305 (N_20305,N_17532,N_11870);
xor U20306 (N_20306,N_16500,N_13647);
nand U20307 (N_20307,N_17528,N_18909);
and U20308 (N_20308,N_13701,N_10165);
nand U20309 (N_20309,N_18789,N_14102);
and U20310 (N_20310,N_16018,N_11534);
xor U20311 (N_20311,N_13627,N_12743);
xor U20312 (N_20312,N_10193,N_17844);
nor U20313 (N_20313,N_16987,N_11834);
xnor U20314 (N_20314,N_18019,N_18252);
or U20315 (N_20315,N_19017,N_19648);
nor U20316 (N_20316,N_18243,N_17944);
nor U20317 (N_20317,N_15020,N_11072);
and U20318 (N_20318,N_15858,N_11981);
and U20319 (N_20319,N_11101,N_17512);
and U20320 (N_20320,N_14739,N_14924);
or U20321 (N_20321,N_18828,N_16145);
or U20322 (N_20322,N_19569,N_14607);
xor U20323 (N_20323,N_15009,N_14892);
or U20324 (N_20324,N_18568,N_18704);
and U20325 (N_20325,N_19957,N_18642);
xnor U20326 (N_20326,N_18272,N_15486);
nand U20327 (N_20327,N_13448,N_16477);
xnor U20328 (N_20328,N_18530,N_15510);
xnor U20329 (N_20329,N_18763,N_12089);
and U20330 (N_20330,N_14475,N_18056);
and U20331 (N_20331,N_12434,N_12074);
and U20332 (N_20332,N_15012,N_15786);
or U20333 (N_20333,N_10715,N_15478);
xor U20334 (N_20334,N_17671,N_17361);
nand U20335 (N_20335,N_18621,N_15895);
xnor U20336 (N_20336,N_18441,N_17534);
nand U20337 (N_20337,N_10813,N_12911);
xor U20338 (N_20338,N_15698,N_18790);
nor U20339 (N_20339,N_12990,N_15570);
xnor U20340 (N_20340,N_15713,N_16440);
and U20341 (N_20341,N_15519,N_14882);
xnor U20342 (N_20342,N_18339,N_14681);
nand U20343 (N_20343,N_13409,N_18085);
xor U20344 (N_20344,N_12069,N_17548);
xor U20345 (N_20345,N_19721,N_11254);
nor U20346 (N_20346,N_13082,N_15592);
nor U20347 (N_20347,N_13848,N_18013);
nand U20348 (N_20348,N_14899,N_15873);
and U20349 (N_20349,N_14346,N_17043);
or U20350 (N_20350,N_17062,N_11499);
nor U20351 (N_20351,N_14450,N_13398);
xnor U20352 (N_20352,N_12284,N_17165);
nor U20353 (N_20353,N_18145,N_10438);
or U20354 (N_20354,N_14241,N_14473);
or U20355 (N_20355,N_12793,N_15029);
or U20356 (N_20356,N_18836,N_17174);
nor U20357 (N_20357,N_18118,N_18868);
xor U20358 (N_20358,N_19126,N_10324);
nand U20359 (N_20359,N_18849,N_16799);
nand U20360 (N_20360,N_12873,N_19296);
nor U20361 (N_20361,N_19194,N_13384);
and U20362 (N_20362,N_19788,N_16242);
and U20363 (N_20363,N_11967,N_10610);
or U20364 (N_20364,N_12387,N_17782);
nand U20365 (N_20365,N_19757,N_11144);
and U20366 (N_20366,N_15619,N_18965);
or U20367 (N_20367,N_19640,N_10435);
or U20368 (N_20368,N_11300,N_12099);
and U20369 (N_20369,N_11335,N_15465);
or U20370 (N_20370,N_11927,N_16379);
and U20371 (N_20371,N_10833,N_15960);
or U20372 (N_20372,N_13569,N_15419);
nor U20373 (N_20373,N_13273,N_18175);
or U20374 (N_20374,N_13476,N_19983);
nor U20375 (N_20375,N_14152,N_12888);
and U20376 (N_20376,N_14848,N_12101);
nand U20377 (N_20377,N_17138,N_15189);
nor U20378 (N_20378,N_15312,N_16015);
nor U20379 (N_20379,N_18648,N_16421);
or U20380 (N_20380,N_12866,N_19134);
or U20381 (N_20381,N_13353,N_16205);
and U20382 (N_20382,N_10114,N_12333);
or U20383 (N_20383,N_10026,N_13364);
and U20384 (N_20384,N_17890,N_16521);
nand U20385 (N_20385,N_17473,N_10927);
xor U20386 (N_20386,N_17602,N_12468);
and U20387 (N_20387,N_12806,N_13758);
nor U20388 (N_20388,N_18182,N_17707);
or U20389 (N_20389,N_18316,N_15359);
or U20390 (N_20390,N_14710,N_18049);
xnor U20391 (N_20391,N_12193,N_11936);
nor U20392 (N_20392,N_10029,N_12038);
or U20393 (N_20393,N_13115,N_12685);
nor U20394 (N_20394,N_19318,N_13113);
or U20395 (N_20395,N_17329,N_18309);
or U20396 (N_20396,N_14609,N_18196);
xor U20397 (N_20397,N_17087,N_10856);
xnor U20398 (N_20398,N_10969,N_19947);
and U20399 (N_20399,N_12181,N_11379);
or U20400 (N_20400,N_15339,N_18698);
and U20401 (N_20401,N_13522,N_10340);
and U20402 (N_20402,N_11842,N_19591);
xor U20403 (N_20403,N_17461,N_14906);
xnor U20404 (N_20404,N_18951,N_11571);
nand U20405 (N_20405,N_11090,N_10639);
nor U20406 (N_20406,N_14558,N_11624);
nand U20407 (N_20407,N_18814,N_18929);
and U20408 (N_20408,N_18939,N_15146);
nand U20409 (N_20409,N_13373,N_15130);
and U20410 (N_20410,N_12112,N_10213);
nor U20411 (N_20411,N_19094,N_17880);
nand U20412 (N_20412,N_10450,N_17307);
or U20413 (N_20413,N_15539,N_10629);
nand U20414 (N_20414,N_10443,N_16630);
or U20415 (N_20415,N_16880,N_18314);
xor U20416 (N_20416,N_10458,N_10283);
and U20417 (N_20417,N_19851,N_13432);
or U20418 (N_20418,N_17650,N_17735);
nor U20419 (N_20419,N_11761,N_11491);
nand U20420 (N_20420,N_16221,N_19709);
nand U20421 (N_20421,N_18214,N_16462);
nor U20422 (N_20422,N_19970,N_11051);
nor U20423 (N_20423,N_14876,N_12088);
nand U20424 (N_20424,N_15665,N_15565);
nor U20425 (N_20425,N_12243,N_14463);
nor U20426 (N_20426,N_17616,N_13864);
or U20427 (N_20427,N_10416,N_17093);
or U20428 (N_20428,N_15961,N_14316);
or U20429 (N_20429,N_11045,N_11865);
xor U20430 (N_20430,N_11604,N_14792);
or U20431 (N_20431,N_13814,N_12682);
or U20432 (N_20432,N_18897,N_14519);
nor U20433 (N_20433,N_11556,N_18617);
nand U20434 (N_20434,N_17364,N_16737);
nand U20435 (N_20435,N_16144,N_18543);
xnor U20436 (N_20436,N_18410,N_13458);
nor U20437 (N_20437,N_10375,N_14750);
and U20438 (N_20438,N_14297,N_19267);
and U20439 (N_20439,N_11078,N_12984);
xor U20440 (N_20440,N_17839,N_10085);
nand U20441 (N_20441,N_19576,N_13901);
or U20442 (N_20442,N_14791,N_17270);
and U20443 (N_20443,N_16239,N_10770);
or U20444 (N_20444,N_10736,N_13240);
or U20445 (N_20445,N_11012,N_17468);
or U20446 (N_20446,N_12229,N_17455);
nor U20447 (N_20447,N_12569,N_19186);
xor U20448 (N_20448,N_14011,N_17181);
xnor U20449 (N_20449,N_12006,N_10196);
and U20450 (N_20450,N_18483,N_16025);
and U20451 (N_20451,N_14973,N_19621);
nor U20452 (N_20452,N_10769,N_19552);
nand U20453 (N_20453,N_19708,N_15937);
nor U20454 (N_20454,N_15997,N_16922);
or U20455 (N_20455,N_18982,N_16333);
and U20456 (N_20456,N_14515,N_11476);
nor U20457 (N_20457,N_11165,N_10703);
nor U20458 (N_20458,N_14962,N_17977);
nand U20459 (N_20459,N_11990,N_13555);
or U20460 (N_20460,N_19556,N_14283);
nor U20461 (N_20461,N_16345,N_17136);
nand U20462 (N_20462,N_19188,N_10870);
nor U20463 (N_20463,N_10908,N_11928);
nor U20464 (N_20464,N_17787,N_14803);
nand U20465 (N_20465,N_16358,N_13331);
xnor U20466 (N_20466,N_17344,N_15347);
xor U20467 (N_20467,N_15261,N_12031);
or U20468 (N_20468,N_17484,N_13787);
and U20469 (N_20469,N_18647,N_13457);
nand U20470 (N_20470,N_15370,N_13914);
nand U20471 (N_20471,N_12759,N_18529);
or U20472 (N_20472,N_11889,N_19426);
or U20473 (N_20473,N_19059,N_15636);
nor U20474 (N_20474,N_16011,N_19784);
nand U20475 (N_20475,N_13727,N_19735);
nand U20476 (N_20476,N_11189,N_16091);
and U20477 (N_20477,N_18666,N_14412);
or U20478 (N_20478,N_15734,N_12657);
or U20479 (N_20479,N_19354,N_14895);
nand U20480 (N_20480,N_17737,N_14891);
nor U20481 (N_20481,N_17482,N_16969);
nand U20482 (N_20482,N_16292,N_15718);
nor U20483 (N_20483,N_15892,N_15536);
or U20484 (N_20484,N_18151,N_15288);
xnor U20485 (N_20485,N_13272,N_16934);
or U20486 (N_20486,N_10978,N_19182);
xnor U20487 (N_20487,N_17821,N_15007);
xnor U20488 (N_20488,N_16495,N_18723);
nor U20489 (N_20489,N_12003,N_15479);
nor U20490 (N_20490,N_10391,N_11514);
nand U20491 (N_20491,N_15607,N_10007);
and U20492 (N_20492,N_18589,N_11778);
nor U20493 (N_20493,N_19771,N_18077);
nor U20494 (N_20494,N_14267,N_10310);
xnor U20495 (N_20495,N_18598,N_10009);
and U20496 (N_20496,N_10875,N_16890);
nor U20497 (N_20497,N_13949,N_17146);
and U20498 (N_20498,N_19446,N_15942);
or U20499 (N_20499,N_12071,N_19929);
and U20500 (N_20500,N_14165,N_18492);
or U20501 (N_20501,N_12979,N_17216);
xor U20502 (N_20502,N_19107,N_14754);
or U20503 (N_20503,N_10207,N_17072);
xor U20504 (N_20504,N_15057,N_16910);
nor U20505 (N_20505,N_15569,N_14453);
nand U20506 (N_20506,N_19344,N_13847);
and U20507 (N_20507,N_11393,N_17006);
nand U20508 (N_20508,N_12535,N_16705);
and U20509 (N_20509,N_19219,N_11518);
xor U20510 (N_20510,N_12869,N_17208);
nand U20511 (N_20511,N_19163,N_10535);
nand U20512 (N_20512,N_11565,N_11174);
nand U20513 (N_20513,N_19148,N_11930);
or U20514 (N_20514,N_14119,N_17506);
xnor U20515 (N_20515,N_17801,N_13641);
or U20516 (N_20516,N_12620,N_15043);
or U20517 (N_20517,N_13176,N_18537);
nand U20518 (N_20518,N_10232,N_16148);
or U20519 (N_20519,N_12304,N_19369);
nand U20520 (N_20520,N_18653,N_10877);
nand U20521 (N_20521,N_10505,N_11077);
xnor U20522 (N_20522,N_12885,N_12493);
nor U20523 (N_20523,N_13140,N_19425);
nand U20524 (N_20524,N_14292,N_12586);
or U20525 (N_20525,N_14832,N_10918);
nand U20526 (N_20526,N_19356,N_16813);
and U20527 (N_20527,N_17766,N_16647);
or U20528 (N_20528,N_10936,N_10690);
or U20529 (N_20529,N_12273,N_13474);
xor U20530 (N_20530,N_15250,N_17715);
nor U20531 (N_20531,N_13461,N_17591);
nor U20532 (N_20532,N_15508,N_13877);
and U20533 (N_20533,N_11261,N_11240);
xor U20534 (N_20534,N_10352,N_11332);
or U20535 (N_20535,N_14315,N_15837);
nor U20536 (N_20536,N_19737,N_17149);
or U20537 (N_20537,N_14781,N_19443);
nand U20538 (N_20538,N_11175,N_13372);
nor U20539 (N_20539,N_17878,N_17129);
or U20540 (N_20540,N_18991,N_14427);
nand U20541 (N_20541,N_15572,N_13805);
nand U20542 (N_20542,N_15814,N_14563);
or U20543 (N_20543,N_13105,N_18139);
and U20544 (N_20544,N_19448,N_12774);
or U20545 (N_20545,N_14105,N_17982);
or U20546 (N_20546,N_10942,N_17127);
nor U20547 (N_20547,N_15316,N_13585);
nor U20548 (N_20548,N_11170,N_19283);
nor U20549 (N_20549,N_13796,N_18426);
and U20550 (N_20550,N_17394,N_11095);
nand U20551 (N_20551,N_15237,N_12746);
and U20552 (N_20552,N_10538,N_19828);
xor U20553 (N_20553,N_10268,N_16433);
nand U20554 (N_20554,N_18514,N_10636);
nand U20555 (N_20555,N_18697,N_17033);
and U20556 (N_20556,N_19101,N_10140);
and U20557 (N_20557,N_14929,N_18403);
xor U20558 (N_20558,N_18296,N_12914);
and U20559 (N_20559,N_12820,N_14135);
and U20560 (N_20560,N_18694,N_18787);
nand U20561 (N_20561,N_15583,N_14314);
xnor U20562 (N_20562,N_13134,N_11552);
nand U20563 (N_20563,N_15634,N_17561);
xnor U20564 (N_20564,N_12305,N_10105);
or U20565 (N_20565,N_18321,N_14479);
nor U20566 (N_20566,N_10314,N_15320);
or U20567 (N_20567,N_19945,N_19554);
or U20568 (N_20568,N_19756,N_13812);
nand U20569 (N_20569,N_14970,N_11306);
xnor U20570 (N_20570,N_11322,N_17983);
and U20571 (N_20571,N_13655,N_11248);
or U20572 (N_20572,N_19062,N_15241);
xor U20573 (N_20573,N_19513,N_11805);
nand U20574 (N_20574,N_14012,N_15111);
and U20575 (N_20575,N_16415,N_10494);
nand U20576 (N_20576,N_15736,N_10194);
and U20577 (N_20577,N_12592,N_15074);
and U20578 (N_20578,N_10217,N_15101);
nor U20579 (N_20579,N_12242,N_16551);
xor U20580 (N_20580,N_14560,N_16140);
nand U20581 (N_20581,N_16866,N_13188);
xnor U20582 (N_20582,N_18146,N_19135);
and U20583 (N_20583,N_16161,N_10592);
and U20584 (N_20584,N_13009,N_15402);
xnor U20585 (N_20585,N_11659,N_18421);
and U20586 (N_20586,N_11327,N_11762);
nand U20587 (N_20587,N_15041,N_10149);
or U20588 (N_20588,N_19133,N_17352);
xor U20589 (N_20589,N_10668,N_19674);
and U20590 (N_20590,N_11410,N_15690);
xor U20591 (N_20591,N_18977,N_17951);
nor U20592 (N_20592,N_14628,N_14746);
nand U20593 (N_20593,N_13136,N_13220);
or U20594 (N_20594,N_15063,N_16094);
nor U20595 (N_20595,N_10501,N_13603);
nand U20596 (N_20596,N_17345,N_18488);
or U20597 (N_20597,N_13507,N_19244);
and U20598 (N_20598,N_18891,N_18613);
nor U20599 (N_20599,N_13374,N_10916);
and U20600 (N_20600,N_10052,N_18457);
or U20601 (N_20601,N_17132,N_14348);
or U20602 (N_20602,N_11094,N_14495);
xor U20603 (N_20603,N_12815,N_17337);
nand U20604 (N_20604,N_10141,N_16952);
nand U20605 (N_20605,N_14850,N_11905);
nor U20606 (N_20606,N_14531,N_11914);
nand U20607 (N_20607,N_13270,N_10717);
nor U20608 (N_20608,N_16568,N_12729);
nor U20609 (N_20609,N_17724,N_16834);
nor U20610 (N_20610,N_19139,N_15882);
nand U20611 (N_20611,N_10247,N_19321);
and U20612 (N_20612,N_16121,N_17608);
nor U20613 (N_20613,N_14488,N_15503);
or U20614 (N_20614,N_12162,N_19394);
and U20615 (N_20615,N_17116,N_14636);
nor U20616 (N_20616,N_16776,N_12619);
nor U20617 (N_20617,N_15387,N_12691);
nor U20618 (N_20618,N_15748,N_17665);
nor U20619 (N_20619,N_12915,N_16777);
xor U20620 (N_20620,N_10064,N_14033);
nand U20621 (N_20621,N_15813,N_12120);
nand U20622 (N_20622,N_12960,N_13044);
nor U20623 (N_20623,N_19221,N_12349);
and U20624 (N_20624,N_15825,N_12170);
nand U20625 (N_20625,N_15724,N_18072);
nand U20626 (N_20626,N_16359,N_15187);
nand U20627 (N_20627,N_11607,N_11511);
nor U20628 (N_20628,N_14483,N_12472);
or U20629 (N_20629,N_10849,N_15447);
nor U20630 (N_20630,N_14364,N_10277);
nor U20631 (N_20631,N_13683,N_11989);
nand U20632 (N_20632,N_16768,N_14505);
xor U20633 (N_20633,N_11462,N_13090);
or U20634 (N_20634,N_10713,N_14903);
and U20635 (N_20635,N_12432,N_14440);
or U20636 (N_20636,N_19034,N_15308);
xor U20637 (N_20637,N_14551,N_18886);
and U20638 (N_20638,N_13792,N_14227);
or U20639 (N_20639,N_19463,N_19716);
nand U20640 (N_20640,N_13828,N_16849);
xnor U20641 (N_20641,N_14732,N_18772);
nor U20642 (N_20642,N_12458,N_16175);
nand U20643 (N_20643,N_13418,N_15933);
nand U20644 (N_20644,N_14808,N_17014);
and U20645 (N_20645,N_12673,N_18602);
xnor U20646 (N_20646,N_18761,N_15488);
nor U20647 (N_20647,N_12417,N_12896);
nand U20648 (N_20648,N_14524,N_14582);
nor U20649 (N_20649,N_17135,N_16282);
or U20650 (N_20650,N_11775,N_14325);
nand U20651 (N_20651,N_15532,N_17633);
or U20652 (N_20652,N_18811,N_11040);
nor U20653 (N_20653,N_17318,N_15371);
and U20654 (N_20654,N_11320,N_13336);
and U20655 (N_20655,N_12646,N_14038);
nand U20656 (N_20656,N_13547,N_12606);
or U20657 (N_20657,N_10236,N_16889);
xor U20658 (N_20658,N_18926,N_19881);
or U20659 (N_20659,N_12176,N_13132);
nor U20660 (N_20660,N_13236,N_16422);
or U20661 (N_20661,N_14839,N_15126);
nand U20662 (N_20662,N_12103,N_14615);
nand U20663 (N_20663,N_19511,N_14799);
xnor U20664 (N_20664,N_10650,N_10509);
xnor U20665 (N_20665,N_17171,N_18523);
nand U20666 (N_20666,N_11232,N_11086);
or U20667 (N_20667,N_11372,N_10402);
nor U20668 (N_20668,N_13181,N_19889);
or U20669 (N_20669,N_13681,N_18906);
nor U20670 (N_20670,N_12225,N_10651);
nor U20671 (N_20671,N_13646,N_13225);
nor U20672 (N_20672,N_11529,N_13135);
xnor U20673 (N_20673,N_10240,N_18831);
nor U20674 (N_20674,N_13283,N_18743);
and U20675 (N_20675,N_18315,N_19972);
nand U20676 (N_20676,N_10851,N_14415);
and U20677 (N_20677,N_15600,N_15502);
nor U20678 (N_20678,N_14468,N_16715);
nand U20679 (N_20679,N_10226,N_18673);
nor U20680 (N_20680,N_18109,N_18851);
xor U20681 (N_20681,N_19137,N_12204);
nand U20682 (N_20682,N_19297,N_12546);
nand U20683 (N_20683,N_15277,N_17514);
and U20684 (N_20684,N_14192,N_16741);
or U20685 (N_20685,N_18821,N_11250);
nand U20686 (N_20686,N_12141,N_16786);
nor U20687 (N_20687,N_12744,N_14940);
and U20688 (N_20688,N_18783,N_12218);
or U20689 (N_20689,N_12783,N_19830);
and U20690 (N_20690,N_13589,N_11023);
and U20691 (N_20691,N_19273,N_10686);
and U20692 (N_20692,N_10465,N_18160);
nand U20693 (N_20693,N_19764,N_14840);
and U20694 (N_20694,N_13204,N_11698);
nand U20695 (N_20695,N_15264,N_12568);
nand U20696 (N_20696,N_14703,N_13304);
nand U20697 (N_20697,N_12063,N_12836);
xor U20698 (N_20698,N_12675,N_13129);
nand U20699 (N_20699,N_19761,N_18313);
xnor U20700 (N_20700,N_10730,N_10985);
nor U20701 (N_20701,N_18644,N_11395);
nor U20702 (N_20702,N_14018,N_14860);
xnor U20703 (N_20703,N_12009,N_15575);
or U20704 (N_20704,N_14296,N_15405);
or U20705 (N_20705,N_13194,N_18803);
nand U20706 (N_20706,N_15824,N_17090);
and U20707 (N_20707,N_19719,N_19191);
nor U20708 (N_20708,N_16020,N_10808);
and U20709 (N_20709,N_16173,N_11871);
nor U20710 (N_20710,N_11558,N_15066);
and U20711 (N_20711,N_10531,N_18247);
and U20712 (N_20712,N_11387,N_19543);
xor U20713 (N_20713,N_16231,N_19377);
xnor U20714 (N_20714,N_19821,N_16562);
nor U20715 (N_20715,N_17015,N_16056);
xnor U20716 (N_20716,N_16417,N_11439);
and U20717 (N_20717,N_12151,N_18347);
xnor U20718 (N_20718,N_15275,N_11859);
or U20719 (N_20719,N_18438,N_15418);
nor U20720 (N_20720,N_10408,N_17305);
xnor U20721 (N_20721,N_18289,N_17034);
nand U20722 (N_20722,N_12097,N_13310);
nand U20723 (N_20723,N_17077,N_17107);
or U20724 (N_20724,N_16993,N_12710);
nand U20725 (N_20725,N_12764,N_10492);
xnor U20726 (N_20726,N_16414,N_13577);
and U20727 (N_20727,N_14079,N_12402);
nor U20728 (N_20728,N_10086,N_15484);
and U20729 (N_20729,N_16424,N_16552);
xor U20730 (N_20730,N_12280,N_17476);
nand U20731 (N_20731,N_15313,N_19575);
xor U20732 (N_20732,N_15980,N_14649);
nor U20733 (N_20733,N_11746,N_10162);
and U20734 (N_20734,N_12978,N_17727);
xor U20735 (N_20735,N_17752,N_10081);
xnor U20736 (N_20736,N_19100,N_15427);
nor U20737 (N_20737,N_18287,N_16848);
nand U20738 (N_20738,N_14907,N_15184);
nand U20739 (N_20739,N_13562,N_16836);
xor U20740 (N_20740,N_10763,N_11830);
or U20741 (N_20741,N_17679,N_17655);
and U20742 (N_20742,N_12062,N_19122);
nor U20743 (N_20743,N_10311,N_10163);
nand U20744 (N_20744,N_10235,N_19019);
nor U20745 (N_20745,N_17255,N_18953);
xnor U20746 (N_20746,N_10725,N_10121);
or U20747 (N_20747,N_19959,N_14693);
or U20748 (N_20748,N_19679,N_17647);
xnor U20749 (N_20749,N_11728,N_13192);
or U20750 (N_20750,N_13971,N_13493);
nand U20751 (N_20751,N_13473,N_16767);
and U20752 (N_20752,N_19966,N_10224);
and U20753 (N_20753,N_16646,N_10360);
nand U20754 (N_20754,N_19732,N_13300);
xor U20755 (N_20755,N_12590,N_16526);
nand U20756 (N_20756,N_17717,N_18327);
xnor U20757 (N_20757,N_10700,N_11826);
xnor U20758 (N_20758,N_16806,N_15972);
nand U20759 (N_20759,N_14177,N_18714);
xnor U20760 (N_20760,N_11593,N_17343);
nor U20761 (N_20761,N_10683,N_14308);
or U20762 (N_20762,N_11832,N_13772);
or U20763 (N_20763,N_10934,N_12697);
nand U20764 (N_20764,N_18658,N_13421);
or U20765 (N_20765,N_10981,N_19800);
xnor U20766 (N_20766,N_11184,N_14378);
nor U20767 (N_20767,N_19847,N_19507);
xor U20768 (N_20768,N_19453,N_12585);
and U20769 (N_20769,N_14251,N_11950);
or U20770 (N_20770,N_16740,N_18419);
or U20771 (N_20771,N_19216,N_12228);
or U20772 (N_20772,N_16846,N_11873);
nor U20773 (N_20773,N_16310,N_14944);
or U20774 (N_20774,N_15167,N_11680);
nand U20775 (N_20775,N_11067,N_16734);
nor U20776 (N_20776,N_14581,N_18856);
and U20777 (N_20777,N_17002,N_19436);
xor U20778 (N_20778,N_10073,N_11792);
or U20779 (N_20779,N_16977,N_18364);
and U20780 (N_20780,N_16533,N_15771);
nand U20781 (N_20781,N_16026,N_19694);
nand U20782 (N_20782,N_13053,N_19964);
xor U20783 (N_20783,N_16504,N_10972);
nor U20784 (N_20784,N_12756,N_12974);
and U20785 (N_20785,N_17617,N_12317);
or U20786 (N_20786,N_15341,N_16549);
and U20787 (N_20787,N_16287,N_13572);
and U20788 (N_20788,N_12771,N_13296);
and U20789 (N_20789,N_16083,N_17224);
or U20790 (N_20790,N_10005,N_11768);
or U20791 (N_20791,N_18838,N_19304);
nor U20792 (N_20792,N_12504,N_13995);
xor U20793 (N_20793,N_12414,N_16318);
nor U20794 (N_20794,N_17162,N_12054);
nor U20795 (N_20795,N_16543,N_18005);
and U20796 (N_20796,N_17438,N_18937);
nor U20797 (N_20797,N_15742,N_15676);
and U20798 (N_20798,N_15979,N_14849);
and U20799 (N_20799,N_15263,N_10772);
nor U20800 (N_20800,N_14120,N_13498);
and U20801 (N_20801,N_18362,N_16676);
nor U20802 (N_20802,N_16209,N_12350);
and U20803 (N_20803,N_16400,N_18253);
nand U20804 (N_20804,N_19239,N_17110);
nand U20805 (N_20805,N_16637,N_15670);
nand U20806 (N_20806,N_10895,N_15714);
nor U20807 (N_20807,N_14925,N_19488);
nor U20808 (N_20808,N_12539,N_10518);
or U20809 (N_20809,N_16645,N_10298);
or U20810 (N_20810,N_16795,N_10802);
xor U20811 (N_20811,N_19170,N_13801);
or U20812 (N_20812,N_12598,N_15225);
or U20813 (N_20813,N_17718,N_14063);
xnor U20814 (N_20814,N_10525,N_16463);
and U20815 (N_20815,N_13351,N_18599);
and U20816 (N_20816,N_10275,N_16873);
xor U20817 (N_20817,N_11153,N_14728);
and U20818 (N_20818,N_19226,N_16631);
or U20819 (N_20819,N_18961,N_14989);
and U20820 (N_20820,N_13962,N_15028);
and U20821 (N_20821,N_18954,N_19444);
xor U20822 (N_20822,N_11801,N_13259);
and U20823 (N_20823,N_13916,N_14931);
or U20824 (N_20824,N_10431,N_11540);
and U20825 (N_20825,N_14245,N_12516);
nor U20826 (N_20826,N_18437,N_10880);
and U20827 (N_20827,N_11637,N_17682);
nand U20828 (N_20828,N_14562,N_19641);
and U20829 (N_20829,N_10554,N_12758);
and U20830 (N_20830,N_18998,N_15068);
and U20831 (N_20831,N_15681,N_12524);
and U20832 (N_20832,N_15603,N_10692);
nand U20833 (N_20833,N_13008,N_16404);
xor U20834 (N_20834,N_11504,N_13639);
xor U20835 (N_20835,N_11616,N_10562);
nor U20836 (N_20836,N_12757,N_19489);
and U20837 (N_20837,N_13318,N_14218);
or U20838 (N_20838,N_12879,N_15208);
nor U20839 (N_20839,N_19097,N_19333);
nor U20840 (N_20840,N_16195,N_15954);
and U20841 (N_20841,N_11679,N_15504);
nand U20842 (N_20842,N_13592,N_18203);
xnor U20843 (N_20843,N_11695,N_17811);
nor U20844 (N_20844,N_11586,N_16198);
or U20845 (N_20845,N_13798,N_13654);
and U20846 (N_20846,N_11648,N_16621);
xor U20847 (N_20847,N_17407,N_13110);
nor U20848 (N_20848,N_16679,N_18588);
or U20849 (N_20849,N_14620,N_13746);
nand U20850 (N_20850,N_17598,N_10251);
xor U20851 (N_20851,N_11020,N_10527);
xor U20852 (N_20852,N_14390,N_16689);
or U20853 (N_20853,N_15437,N_18167);
or U20854 (N_20854,N_11622,N_19346);
xor U20855 (N_20855,N_13693,N_13606);
nor U20856 (N_20856,N_15896,N_12169);
nand U20857 (N_20857,N_13175,N_16479);
or U20858 (N_20858,N_14284,N_13975);
xnor U20859 (N_20859,N_18227,N_19330);
nand U20860 (N_20860,N_10313,N_16443);
nor U20861 (N_20861,N_19688,N_19922);
or U20862 (N_20862,N_11670,N_14129);
nor U20863 (N_20863,N_12603,N_11241);
nor U20864 (N_20864,N_17973,N_10405);
or U20865 (N_20865,N_12856,N_11205);
nand U20866 (N_20866,N_18731,N_18600);
and U20867 (N_20867,N_14722,N_14999);
nor U20868 (N_20868,N_12810,N_15901);
or U20869 (N_20869,N_15955,N_19749);
nor U20870 (N_20870,N_12636,N_16380);
or U20871 (N_20871,N_12148,N_12931);
nand U20872 (N_20872,N_12013,N_10829);
xor U20873 (N_20873,N_14387,N_11539);
and U20874 (N_20874,N_13928,N_18009);
nor U20875 (N_20875,N_15953,N_11769);
or U20876 (N_20876,N_17847,N_15330);
nor U20877 (N_20877,N_11457,N_17296);
or U20878 (N_20878,N_19524,N_16906);
xor U20879 (N_20879,N_16954,N_12987);
or U20880 (N_20880,N_11206,N_15538);
or U20881 (N_20881,N_15211,N_19845);
and U20882 (N_20882,N_15723,N_19668);
nor U20883 (N_20883,N_18519,N_10089);
xor U20884 (N_20884,N_10923,N_15751);
or U20885 (N_20885,N_14819,N_14783);
xnor U20886 (N_20886,N_18218,N_16764);
and U20887 (N_20887,N_13102,N_13666);
xnor U20888 (N_20888,N_18975,N_15408);
xor U20889 (N_20889,N_13481,N_10295);
xnor U20890 (N_20890,N_10989,N_13667);
xnor U20891 (N_20891,N_14645,N_10603);
nor U20892 (N_20892,N_19549,N_10145);
xnor U20893 (N_20893,N_17232,N_17833);
and U20894 (N_20894,N_16325,N_12043);
or U20895 (N_20895,N_15487,N_18407);
nand U20896 (N_20896,N_15076,N_16917);
or U20897 (N_20897,N_12327,N_14124);
xor U20898 (N_20898,N_16574,N_13430);
and U20899 (N_20899,N_13829,N_13920);
nor U20900 (N_20900,N_17923,N_16772);
or U20901 (N_20901,N_13957,N_17967);
nor U20902 (N_20902,N_17022,N_18716);
and U20903 (N_20903,N_16134,N_19918);
nor U20904 (N_20904,N_18111,N_11330);
nand U20905 (N_20905,N_19900,N_17448);
and U20906 (N_20906,N_19458,N_16747);
xor U20907 (N_20907,N_14941,N_10785);
or U20908 (N_20908,N_10739,N_11107);
nor U20909 (N_20909,N_18895,N_16371);
nor U20910 (N_20910,N_18014,N_17542);
or U20911 (N_20911,N_10859,N_11893);
or U20912 (N_20912,N_11285,N_14443);
xor U20913 (N_20913,N_18893,N_12381);
or U20914 (N_20914,N_12738,N_18154);
xor U20915 (N_20915,N_11391,N_13747);
nand U20916 (N_20916,N_10374,N_18619);
and U20917 (N_20917,N_12843,N_18756);
and U20918 (N_20918,N_14015,N_16731);
or U20919 (N_20919,N_13037,N_19050);
nand U20920 (N_20920,N_19082,N_12881);
nor U20921 (N_20921,N_12293,N_19203);
and U20922 (N_20922,N_13161,N_12467);
xor U20923 (N_20923,N_13087,N_18740);
and U20924 (N_20924,N_10387,N_14210);
and U20925 (N_20925,N_17283,N_19562);
xor U20926 (N_20926,N_18298,N_10045);
nor U20927 (N_20927,N_10342,N_10680);
xnor U20928 (N_20928,N_17466,N_15560);
nor U20929 (N_20929,N_13403,N_17362);
xnor U20930 (N_20930,N_13887,N_16509);
or U20931 (N_20931,N_18311,N_15719);
xor U20932 (N_20932,N_17258,N_19869);
nand U20933 (N_20933,N_19516,N_12202);
xor U20934 (N_20934,N_10924,N_10348);
xor U20935 (N_20935,N_10627,N_18193);
nor U20936 (N_20936,N_14277,N_17957);
xor U20937 (N_20937,N_11443,N_17994);
nor U20938 (N_20938,N_15757,N_19605);
or U20939 (N_20939,N_17554,N_11960);
xor U20940 (N_20940,N_13556,N_19347);
or U20941 (N_20941,N_17253,N_10886);
xor U20942 (N_20942,N_11507,N_15699);
or U20943 (N_20943,N_13416,N_13154);
and U20944 (N_20944,N_19836,N_19651);
and U20945 (N_20945,N_13586,N_12137);
nand U20946 (N_20946,N_17914,N_14191);
or U20947 (N_20947,N_12294,N_11452);
or U20948 (N_20948,N_12165,N_11786);
or U20949 (N_20949,N_16832,N_14180);
nand U20950 (N_20950,N_12129,N_16608);
xnor U20951 (N_20951,N_11582,N_15552);
and U20952 (N_20952,N_15096,N_19860);
or U20953 (N_20953,N_14996,N_11223);
nor U20954 (N_20954,N_14019,N_11545);
or U20955 (N_20955,N_10185,N_13206);
nor U20956 (N_20956,N_14557,N_11942);
xor U20957 (N_20957,N_13531,N_19981);
nand U20958 (N_20958,N_17798,N_10237);
and U20959 (N_20959,N_12076,N_12973);
or U20960 (N_20960,N_14674,N_13355);
xor U20961 (N_20961,N_17175,N_13672);
and U20962 (N_20962,N_13243,N_17836);
or U20963 (N_20963,N_13454,N_13890);
or U20964 (N_20964,N_13503,N_16603);
xnor U20965 (N_20965,N_18920,N_15033);
nand U20966 (N_20966,N_12470,N_17178);
and U20967 (N_20967,N_18479,N_15372);
nor U20968 (N_20968,N_16078,N_10638);
nand U20969 (N_20969,N_10968,N_19684);
and U20970 (N_20970,N_14605,N_12367);
nor U20971 (N_20971,N_19355,N_19392);
or U20972 (N_20972,N_16920,N_17443);
nand U20973 (N_20973,N_13615,N_10613);
nand U20974 (N_20974,N_12972,N_16070);
or U20975 (N_20975,N_19247,N_17958);
or U20976 (N_20976,N_13938,N_16694);
nand U20977 (N_20977,N_15231,N_15412);
and U20978 (N_20978,N_16807,N_18066);
nand U20979 (N_20979,N_10309,N_16068);
or U20980 (N_20980,N_16702,N_14254);
xnor U20981 (N_20981,N_15367,N_14694);
nor U20982 (N_20982,N_14985,N_18370);
or U20983 (N_20983,N_11931,N_12704);
and U20984 (N_20984,N_11134,N_11703);
nor U20985 (N_20985,N_11743,N_14299);
xnor U20986 (N_20986,N_15244,N_10591);
nor U20987 (N_20987,N_12245,N_11389);
nand U20988 (N_20988,N_18778,N_14391);
nor U20989 (N_20989,N_19573,N_17301);
and U20990 (N_20990,N_15947,N_18796);
and U20991 (N_20991,N_11220,N_13089);
nor U20992 (N_20992,N_13055,N_19197);
and U20993 (N_20993,N_15091,N_10970);
nor U20994 (N_20994,N_12628,N_11968);
nand U20995 (N_20995,N_15245,N_18678);
xnor U20996 (N_20996,N_17064,N_13485);
xnor U20997 (N_20997,N_15094,N_15314);
nand U20998 (N_20998,N_13844,N_18930);
nor U20999 (N_20999,N_10761,N_13214);
or U21000 (N_21000,N_13854,N_19233);
xnor U21001 (N_21001,N_13884,N_18494);
and U21002 (N_21002,N_15201,N_13856);
nand U21003 (N_21003,N_11952,N_17265);
and U21004 (N_21004,N_16739,N_16203);
nor U21005 (N_21005,N_10210,N_14309);
or U21006 (N_21006,N_16662,N_12015);
nor U21007 (N_21007,N_17986,N_14130);
nor U21008 (N_21008,N_11543,N_14589);
nor U21009 (N_21009,N_14623,N_11486);
xor U21010 (N_21010,N_15049,N_13660);
xor U21011 (N_21011,N_18346,N_16589);
nor U21012 (N_21012,N_17024,N_12448);
or U21013 (N_21013,N_10954,N_12563);
or U21014 (N_21014,N_17703,N_10129);
nor U21015 (N_21015,N_16897,N_15852);
or U21016 (N_21016,N_16212,N_14401);
nand U21017 (N_21017,N_12542,N_10496);
xor U21018 (N_21018,N_12451,N_15904);
and U21019 (N_21019,N_13347,N_10202);
nand U21020 (N_21020,N_14874,N_15301);
xor U21021 (N_21021,N_14305,N_13218);
and U21022 (N_21022,N_13150,N_19731);
nor U21023 (N_21023,N_19506,N_17803);
xor U21024 (N_21024,N_17991,N_13325);
xor U21025 (N_21025,N_18052,N_18616);
nand U21026 (N_21026,N_10893,N_19998);
nand U21027 (N_21027,N_10551,N_17788);
or U21028 (N_21028,N_16409,N_17207);
xor U21029 (N_21029,N_17774,N_14590);
or U21030 (N_21030,N_17249,N_13744);
nand U21031 (N_21031,N_14057,N_17037);
xnor U21032 (N_21032,N_10944,N_16941);
xnor U21033 (N_21033,N_16678,N_12837);
or U21034 (N_21034,N_12289,N_15936);
nor U21035 (N_21035,N_11363,N_11860);
nand U21036 (N_21036,N_12544,N_13297);
nand U21037 (N_21037,N_17056,N_17051);
or U21038 (N_21038,N_15496,N_17907);
and U21039 (N_21039,N_12244,N_14789);
nor U21040 (N_21040,N_16788,N_12860);
or U21041 (N_21041,N_12953,N_19664);
xor U21042 (N_21042,N_14720,N_14622);
nor U21043 (N_21043,N_16071,N_19158);
and U21044 (N_21044,N_12992,N_10172);
or U21045 (N_21045,N_17122,N_10914);
nand U21046 (N_21046,N_16916,N_10550);
nand U21047 (N_21047,N_17985,N_18574);
or U21048 (N_21048,N_14388,N_14617);
nand U21049 (N_21049,N_15077,N_18245);
and U21050 (N_21050,N_14911,N_16956);
and U21051 (N_21051,N_17694,N_15270);
and U21052 (N_21052,N_16218,N_16223);
or U21053 (N_21053,N_18045,N_14482);
nor U21054 (N_21054,N_11048,N_17520);
nand U21055 (N_21055,N_14270,N_13527);
nand U21056 (N_21056,N_13534,N_15349);
nor U21057 (N_21057,N_14252,N_15449);
xnor U21058 (N_21058,N_18509,N_11696);
nand U21059 (N_21059,N_11784,N_11430);
nand U21060 (N_21060,N_11678,N_19466);
and U21061 (N_21061,N_18655,N_12517);
xnor U21062 (N_21062,N_10949,N_18394);
and U21063 (N_21063,N_14975,N_18000);
or U21064 (N_21064,N_11505,N_17399);
xnor U21065 (N_21065,N_15417,N_13554);
nand U21066 (N_21066,N_13072,N_15794);
nand U21067 (N_21067,N_13774,N_13610);
nand U21068 (N_21068,N_15119,N_13591);
and U21069 (N_21069,N_12121,N_11238);
and U21070 (N_21070,N_14647,N_15949);
nand U21071 (N_21071,N_15545,N_17759);
or U21072 (N_21072,N_19905,N_13891);
nor U21073 (N_21073,N_15739,N_18163);
xor U21074 (N_21074,N_17375,N_12297);
nor U21075 (N_21075,N_18660,N_14392);
xnor U21076 (N_21076,N_13291,N_12709);
xor U21077 (N_21077,N_12478,N_12270);
nand U21078 (N_21078,N_17293,N_15460);
and U21079 (N_21079,N_18454,N_14413);
xnor U21080 (N_21080,N_19102,N_15880);
nand U21081 (N_21081,N_12454,N_13643);
and U21082 (N_21082,N_15279,N_17552);
or U21083 (N_21083,N_12300,N_17915);
or U21084 (N_21084,N_14619,N_12724);
nor U21085 (N_21085,N_10254,N_17712);
nand U21086 (N_21086,N_15113,N_12683);
nor U21087 (N_21087,N_16507,N_16305);
nor U21088 (N_21088,N_10957,N_19974);
nand U21089 (N_21089,N_19230,N_10257);
and U21090 (N_21090,N_10976,N_12435);
nor U21091 (N_21091,N_11015,N_15444);
or U21092 (N_21092,N_14008,N_15973);
nor U21093 (N_21093,N_11874,N_15989);
nor U21094 (N_21094,N_15403,N_14571);
nand U21095 (N_21095,N_13984,N_15144);
nand U21096 (N_21096,N_11627,N_13311);
nand U21097 (N_21097,N_14930,N_19676);
nand U21098 (N_21098,N_18732,N_16582);
xnor U21099 (N_21099,N_14405,N_10905);
xor U21100 (N_21100,N_19393,N_15162);
nor U21101 (N_21101,N_10135,N_10688);
nor U21102 (N_21102,N_14913,N_13497);
or U21103 (N_21103,N_18657,N_14631);
nor U21104 (N_21104,N_16642,N_15192);
nor U21105 (N_21105,N_10845,N_10058);
nor U21106 (N_21106,N_16202,N_17500);
and U21107 (N_21107,N_12928,N_14005);
or U21108 (N_21108,N_13933,N_12988);
nand U21109 (N_21109,N_10660,N_13768);
or U21110 (N_21110,N_18558,N_19906);
xor U21111 (N_21111,N_14591,N_18065);
nor U21112 (N_21112,N_11621,N_18332);
xnor U21113 (N_21113,N_14586,N_13769);
nor U21114 (N_21114,N_10218,N_14640);
or U21115 (N_21115,N_18060,N_15458);
nor U21116 (N_21116,N_18449,N_15599);
nand U21117 (N_21117,N_19879,N_18352);
and U21118 (N_21118,N_19537,N_17474);
or U21119 (N_21119,N_16277,N_10995);
or U21120 (N_21120,N_15202,N_16847);
nor U21121 (N_21121,N_11231,N_13099);
nor U21122 (N_21122,N_11338,N_14242);
and U21123 (N_21123,N_14434,N_15707);
or U21124 (N_21124,N_19213,N_19769);
and U21125 (N_21125,N_19332,N_15188);
nand U21126 (N_21126,N_14896,N_18430);
and U21127 (N_21127,N_12090,N_19123);
xor U21128 (N_21128,N_12828,N_10493);
xor U21129 (N_21129,N_17285,N_14170);
and U21130 (N_21130,N_17302,N_11716);
and U21131 (N_21131,N_13932,N_19144);
nor U21132 (N_21132,N_10383,N_15325);
and U21133 (N_21133,N_14411,N_10204);
and U21134 (N_21134,N_17882,N_14696);
nand U21135 (N_21135,N_11708,N_13704);
or U21136 (N_21136,N_10634,N_19568);
nor U21137 (N_21137,N_19770,N_18651);
nor U21138 (N_21138,N_12608,N_16456);
xor U21139 (N_21139,N_17054,N_10116);
nand U21140 (N_21140,N_11304,N_12483);
and U21141 (N_21141,N_11964,N_11313);
xnor U21142 (N_21142,N_15498,N_18987);
nor U21143 (N_21143,N_15345,N_16995);
and U21144 (N_21144,N_16634,N_11891);
nor U21145 (N_21145,N_14060,N_16006);
xor U21146 (N_21146,N_10179,N_18912);
nand U21147 (N_21147,N_11245,N_10756);
or U21148 (N_21148,N_19151,N_15755);
or U21149 (N_21149,N_17632,N_13795);
or U21150 (N_21150,N_12580,N_12177);
nand U21151 (N_21151,N_12167,N_10180);
and U21152 (N_21152,N_10563,N_16410);
or U21153 (N_21153,N_18668,N_14410);
nor U21154 (N_21154,N_14257,N_12865);
or U21155 (N_21155,N_16671,N_12252);
and U21156 (N_21156,N_15530,N_10062);
nand U21157 (N_21157,N_18609,N_13130);
and U21158 (N_21158,N_16476,N_16879);
and U21159 (N_21159,N_15448,N_19574);
nor U21160 (N_21160,N_17196,N_10751);
xnor U21161 (N_21161,N_18834,N_11062);
nor U21162 (N_21162,N_13155,N_12848);
xnor U21163 (N_21163,N_17956,N_19696);
or U21164 (N_21164,N_18093,N_16044);
nand U21165 (N_21165,N_12465,N_19667);
xor U21166 (N_21166,N_17999,N_15137);
nor U21167 (N_21167,N_15697,N_11813);
and U21168 (N_21168,N_10080,N_19327);
or U21169 (N_21169,N_10806,N_19211);
xor U21170 (N_21170,N_18824,N_12662);
nand U21171 (N_21171,N_14719,N_17828);
and U21172 (N_21172,N_14705,N_14204);
or U21173 (N_21173,N_16591,N_18465);
nor U21174 (N_21174,N_15150,N_16735);
or U21175 (N_21175,N_18548,N_18329);
or U21176 (N_21176,N_10609,N_16701);
xnor U21177 (N_21177,N_13077,N_12277);
nand U21178 (N_21178,N_11156,N_16196);
or U21179 (N_21179,N_10524,N_15990);
nor U21180 (N_21180,N_10951,N_12376);
or U21181 (N_21181,N_13576,N_17519);
nand U21182 (N_21182,N_12642,N_18840);
nor U21183 (N_21183,N_14873,N_10940);
xnor U21184 (N_21184,N_17144,N_16047);
nand U21185 (N_21185,N_11849,N_14535);
or U21186 (N_21186,N_11587,N_15841);
xor U21187 (N_21187,N_13323,N_18341);
nor U21188 (N_21188,N_13463,N_18972);
xnor U21189 (N_21189,N_18179,N_11253);
nor U21190 (N_21190,N_12077,N_11139);
or U21191 (N_21191,N_12968,N_11619);
and U21192 (N_21192,N_13043,N_16949);
nand U21193 (N_21193,N_17126,N_15774);
xnor U21194 (N_21194,N_11003,N_14755);
xnor U21195 (N_21195,N_13915,N_14024);
xor U21196 (N_21196,N_15730,N_18098);
and U21197 (N_21197,N_19540,N_13101);
or U21198 (N_21198,N_13303,N_14926);
or U21199 (N_21199,N_14056,N_15145);
nor U21200 (N_21200,N_19087,N_11777);
nand U21201 (N_21201,N_19942,N_15910);
xor U21202 (N_21202,N_14510,N_13526);
and U21203 (N_21203,N_17652,N_18988);
and U21204 (N_21204,N_16858,N_16281);
or U21205 (N_21205,N_11120,N_12971);
xnor U21206 (N_21206,N_13262,N_19021);
nor U21207 (N_21207,N_11630,N_19872);
nand U21208 (N_21208,N_15546,N_16829);
and U21209 (N_21209,N_10115,N_10507);
xnor U21210 (N_21210,N_16628,N_19427);
nand U21211 (N_21211,N_12045,N_18682);
and U21212 (N_21212,N_17605,N_15070);
nor U21213 (N_21213,N_12545,N_11319);
xnor U21214 (N_21214,N_19915,N_10423);
nor U21215 (N_21215,N_18560,N_11915);
nand U21216 (N_21216,N_12195,N_16438);
nor U21217 (N_21217,N_10728,N_18236);
or U21218 (N_21218,N_18545,N_19720);
and U21219 (N_21219,N_19582,N_11553);
nand U21220 (N_21220,N_19276,N_13740);
and U21221 (N_21221,N_16994,N_18948);
nand U21222 (N_21222,N_17504,N_16339);
or U21223 (N_21223,N_12551,N_18889);
or U21224 (N_21224,N_18026,N_14355);
nor U21225 (N_21225,N_17580,N_16672);
nor U21226 (N_21226,N_14646,N_18639);
nor U21227 (N_21227,N_19480,N_18952);
nand U21228 (N_21228,N_17076,N_10910);
nor U21229 (N_21229,N_13733,N_17347);
or U21230 (N_21230,N_19056,N_16237);
nor U21231 (N_21231,N_19288,N_15375);
or U21232 (N_21232,N_10701,N_11435);
and U21233 (N_21233,N_13127,N_13093);
nor U21234 (N_21234,N_14878,N_17298);
nand U21235 (N_21235,N_15451,N_12638);
or U21236 (N_21236,N_11956,N_14731);
xnor U21237 (N_21237,N_12316,N_14263);
xor U21238 (N_21238,N_15878,N_17729);
and U21239 (N_21239,N_14253,N_16084);
nor U21240 (N_21240,N_14922,N_13540);
or U21241 (N_21241,N_14377,N_13943);
and U21242 (N_21242,N_18957,N_12020);
xor U21243 (N_21243,N_17876,N_14234);
xor U21244 (N_21244,N_15149,N_11337);
nor U21245 (N_21245,N_19265,N_11998);
nor U21246 (N_21246,N_14639,N_11044);
nand U21247 (N_21247,N_13164,N_12372);
or U21248 (N_21248,N_10820,N_18411);
and U21249 (N_21249,N_17091,N_12811);
xnor U21250 (N_21250,N_14247,N_13686);
or U21251 (N_21251,N_14460,N_12769);
nor U21252 (N_21252,N_12767,N_12932);
nand U21253 (N_21253,N_13508,N_18999);
nor U21254 (N_21254,N_15838,N_12382);
nor U21255 (N_21255,N_17789,N_18582);
nand U21256 (N_21256,N_10675,N_14306);
xnor U21257 (N_21257,N_12386,N_10956);
and U21258 (N_21258,N_14353,N_10533);
nor U21259 (N_21259,N_10633,N_10449);
nand U21260 (N_21260,N_12523,N_15692);
xnor U21261 (N_21261,N_17627,N_11520);
nand U21262 (N_21262,N_17217,N_10866);
nor U21263 (N_21263,N_18733,N_10544);
xor U21264 (N_21264,N_19518,N_16851);
xnor U21265 (N_21265,N_19108,N_12985);
nor U21266 (N_21266,N_19612,N_14393);
and U21267 (N_21267,N_16649,N_19473);
xor U21268 (N_21268,N_18201,N_19820);
and U21269 (N_21269,N_13464,N_19429);
and U21270 (N_21270,N_11276,N_12025);
nand U21271 (N_21271,N_17756,N_10490);
nand U21272 (N_21272,N_16064,N_19535);
and U21273 (N_21273,N_14738,N_16151);
or U21274 (N_21274,N_17585,N_12982);
nand U21275 (N_21275,N_10440,N_12239);
xnor U21276 (N_21276,N_14821,N_18238);
nand U21277 (N_21277,N_10410,N_16580);
nor U21278 (N_21278,N_12886,N_17215);
xor U21279 (N_21279,N_16668,N_19871);
xor U21280 (N_21280,N_14865,N_12993);
and U21281 (N_21281,N_15243,N_19222);
or U21282 (N_21282,N_16619,N_15078);
xnor U21283 (N_21283,N_19541,N_14217);
nand U21284 (N_21284,N_18538,N_18746);
nor U21285 (N_21285,N_12331,N_15909);
or U21286 (N_21286,N_19767,N_17125);
or U21287 (N_21287,N_10349,N_18377);
and U21288 (N_21288,N_10876,N_14981);
nor U21289 (N_21289,N_18835,N_11697);
or U21290 (N_21290,N_15869,N_11902);
or U21291 (N_21291,N_13258,N_11886);
nor U21292 (N_21292,N_13879,N_10615);
xor U21293 (N_21293,N_12528,N_14822);
nand U21294 (N_21294,N_14201,N_15643);
nand U21295 (N_21295,N_12106,N_14294);
nand U21296 (N_21296,N_17426,N_12664);
or U21297 (N_21297,N_19231,N_10334);
nor U21298 (N_21298,N_19350,N_14870);
or U21299 (N_21299,N_17822,N_16035);
or U21300 (N_21300,N_12945,N_14543);
or U21301 (N_21301,N_19692,N_18795);
nor U21302 (N_21302,N_18667,N_13383);
nor U21303 (N_21303,N_17517,N_15992);
or U21304 (N_21304,N_14713,N_16793);
or U21305 (N_21305,N_19977,N_13852);
nand U21306 (N_21306,N_18099,N_12841);
xor U21307 (N_21307,N_17702,N_13994);
or U21308 (N_21308,N_15664,N_13594);
or U21309 (N_21309,N_17976,N_14145);
nor U21310 (N_21310,N_12498,N_13116);
xnor U21311 (N_21311,N_13054,N_15672);
nand U21312 (N_21312,N_17026,N_13664);
and U21313 (N_21313,N_18691,N_19867);
nor U21314 (N_21314,N_15008,N_12104);
and U21315 (N_21315,N_15766,N_11442);
nand U21316 (N_21316,N_15857,N_19452);
or U21317 (N_21317,N_11087,N_13783);
or U21318 (N_21318,N_10545,N_14501);
nor U21319 (N_21319,N_16442,N_12817);
nor U21320 (N_21320,N_11037,N_16073);
nor U21321 (N_21321,N_15374,N_10248);
and U21322 (N_21322,N_11645,N_17905);
xnor U21323 (N_21323,N_19941,N_12499);
and U21324 (N_21324,N_12883,N_15902);
and U21325 (N_21325,N_12895,N_15865);
and U21326 (N_21326,N_17457,N_10757);
and U21327 (N_21327,N_11212,N_10517);
nor U21328 (N_21328,N_12583,N_19428);
nor U21329 (N_21329,N_19173,N_19295);
and U21330 (N_21330,N_15782,N_17799);
nand U21331 (N_21331,N_13378,N_15253);
nand U21332 (N_21332,N_18791,N_19010);
nand U21333 (N_21333,N_10444,N_13104);
nand U21334 (N_21334,N_17188,N_18661);
nand U21335 (N_21335,N_14533,N_11413);
and U21336 (N_21336,N_10900,N_14269);
and U21337 (N_21337,N_11580,N_15788);
and U21338 (N_21338,N_13734,N_10442);
nand U21339 (N_21339,N_10188,N_19833);
and U21340 (N_21340,N_14298,N_11114);
nor U21341 (N_21341,N_12363,N_10466);
nand U21342 (N_21342,N_13873,N_10646);
xor U21343 (N_21343,N_15861,N_11623);
nand U21344 (N_21344,N_10053,N_18579);
nor U21345 (N_21345,N_11700,N_12698);
nand U21346 (N_21346,N_15075,N_10604);
and U21347 (N_21347,N_11551,N_12556);
or U21348 (N_21348,N_10719,N_15025);
and U21349 (N_21349,N_16235,N_11916);
or U21350 (N_21350,N_13111,N_14514);
xnor U21351 (N_21351,N_10258,N_13908);
nand U21352 (N_21352,N_12007,N_18281);
and U21353 (N_21353,N_12839,N_18279);
and U21354 (N_21354,N_19399,N_11727);
and U21355 (N_21355,N_12189,N_14441);
nand U21356 (N_21356,N_17658,N_11006);
and U21357 (N_21357,N_12460,N_19891);
and U21358 (N_21358,N_17761,N_14451);
or U21359 (N_21359,N_16626,N_13295);
and U21360 (N_21360,N_10003,N_18090);
xnor U21361 (N_21361,N_12107,N_18431);
and U21362 (N_21362,N_19154,N_15829);
nand U21363 (N_21363,N_18700,N_14570);
and U21364 (N_21364,N_15461,N_19689);
nor U21365 (N_21365,N_17700,N_13157);
and U21366 (N_21366,N_17049,N_12438);
and U21367 (N_21367,N_11487,N_13245);
nand U21368 (N_21368,N_12184,N_12368);
nor U21369 (N_21369,N_16428,N_18008);
or U21370 (N_21370,N_17736,N_11305);
xor U21371 (N_21371,N_14565,N_19572);
and U21372 (N_21372,N_17879,N_10612);
nand U21373 (N_21373,N_14538,N_11572);
or U21374 (N_21374,N_10699,N_10858);
or U21375 (N_21375,N_14422,N_17437);
nand U21376 (N_21376,N_14770,N_10021);
nand U21377 (N_21377,N_13924,N_17069);
xor U21378 (N_21378,N_15136,N_12705);
and U21379 (N_21379,N_14321,N_12441);
nor U21380 (N_21380,N_16856,N_13886);
nor U21381 (N_21381,N_12473,N_13748);
and U21382 (N_21382,N_17596,N_13467);
or U21383 (N_21383,N_19914,N_18386);
and U21384 (N_21384,N_14435,N_18822);
nand U21385 (N_21385,N_16778,N_15086);
xor U21386 (N_21386,N_12718,N_19275);
or U21387 (N_21387,N_13983,N_12643);
nand U21388 (N_21388,N_16284,N_18627);
and U21389 (N_21389,N_17941,N_11841);
nor U21390 (N_21390,N_14246,N_13999);
nand U21391 (N_21391,N_13992,N_15934);
nand U21392 (N_21392,N_15156,N_16280);
and U21393 (N_21393,N_19902,N_19620);
nor U21394 (N_21394,N_12161,N_11711);
or U21395 (N_21395,N_10002,N_16377);
or U21396 (N_21396,N_14802,N_19630);
and U21397 (N_21397,N_18385,N_10127);
xor U21398 (N_21398,N_13320,N_15594);
xor U21399 (N_21399,N_10656,N_12632);
nand U21400 (N_21400,N_13375,N_10017);
or U21401 (N_21401,N_14107,N_14178);
and U21402 (N_21402,N_16962,N_18522);
and U21403 (N_21403,N_14845,N_10320);
nand U21404 (N_21404,N_11446,N_19181);
and U21405 (N_21405,N_14359,N_17134);
xor U21406 (N_21406,N_18350,N_13968);
nor U21407 (N_21407,N_14014,N_16572);
nand U21408 (N_21408,N_18813,N_14993);
nor U21409 (N_21409,N_18719,N_12282);
and U21410 (N_21410,N_19092,N_10051);
nor U21411 (N_21411,N_15116,N_10854);
nor U21412 (N_21412,N_10060,N_18280);
nor U21413 (N_21413,N_13537,N_19018);
xnor U21414 (N_21414,N_14950,N_10072);
nand U21415 (N_21415,N_14654,N_13571);
xor U21416 (N_21416,N_11819,N_11030);
and U21417 (N_21417,N_14395,N_19910);
or U21418 (N_21418,N_14477,N_17851);
xnor U21419 (N_21419,N_10471,N_17434);
nor U21420 (N_21420,N_10054,N_16569);
xnor U21421 (N_21421,N_13286,N_18531);
and U21422 (N_21422,N_18478,N_13425);
and U21423 (N_21423,N_19961,N_16158);
or U21424 (N_21424,N_15395,N_14480);
nor U21425 (N_21425,N_17147,N_16659);
nor U21426 (N_21426,N_14780,N_19329);
nand U21427 (N_21427,N_14037,N_16141);
and U21428 (N_21428,N_19138,N_17282);
and U21429 (N_21429,N_17281,N_10118);
nor U21430 (N_21430,N_19469,N_19744);
or U21431 (N_21431,N_13499,N_17075);
xor U21432 (N_21432,N_17396,N_18569);
xor U21433 (N_21433,N_10652,N_16982);
nand U21434 (N_21434,N_13293,N_17714);
xnor U21435 (N_21435,N_19982,N_13614);
xor U21436 (N_21436,N_15941,N_13152);
nand U21437 (N_21437,N_16677,N_16697);
and U21438 (N_21438,N_19832,N_18623);
nand U21439 (N_21439,N_12410,N_10522);
xnor U21440 (N_21440,N_12332,N_13048);
xnor U21441 (N_21441,N_17120,N_19924);
xnor U21442 (N_21442,N_10911,N_16798);
nor U21443 (N_21443,N_15490,N_14585);
nand U21444 (N_21444,N_19848,N_17111);
xor U21445 (N_21445,N_19768,N_17357);
xor U21446 (N_21446,N_19072,N_19593);
and U21447 (N_21447,N_13730,N_15141);
and U21448 (N_21448,N_15816,N_18826);
xnor U21449 (N_21449,N_14344,N_17697);
and U21450 (N_21450,N_18170,N_18503);
nor U21451 (N_21451,N_11083,N_14917);
xnor U21452 (N_21452,N_12395,N_14527);
nand U21453 (N_21453,N_10684,N_17830);
nand U21454 (N_21454,N_16867,N_15310);
xnor U21455 (N_21455,N_13633,N_14171);
and U21456 (N_21456,N_17943,N_17677);
nand U21457 (N_21457,N_15287,N_13039);
or U21458 (N_21458,N_10358,N_17016);
or U21459 (N_21459,N_17275,N_11341);
and U21460 (N_21460,N_15352,N_19751);
xor U21461 (N_21461,N_13715,N_15767);
nor U21462 (N_21462,N_17059,N_13806);
xor U21463 (N_21463,N_19358,N_17494);
xnor U21464 (N_21464,N_14190,N_17869);
or U21465 (N_21465,N_12164,N_19656);
xor U21466 (N_21466,N_19927,N_11800);
and U21467 (N_21467,N_14040,N_19269);
nand U21468 (N_21468,N_16216,N_15855);
nor U21469 (N_21469,N_18323,N_13343);
nand U21470 (N_21470,N_11116,N_17575);
or U21471 (N_21471,N_18414,N_13834);
and U21472 (N_21472,N_10239,N_14173);
nand U21473 (N_21473,N_18793,N_19009);
nor U21474 (N_21474,N_19322,N_16699);
and U21475 (N_21475,N_15531,N_12455);
and U21476 (N_21476,N_13523,N_19567);
nor U21477 (N_21477,N_11069,N_18985);
nand U21478 (N_21478,N_14162,N_15872);
and U21479 (N_21479,N_13601,N_19706);
xnor U21480 (N_21480,N_17011,N_16136);
or U21481 (N_21481,N_18830,N_16029);
and U21482 (N_21482,N_14980,N_14642);
or U21483 (N_21483,N_15662,N_19622);
or U21484 (N_21484,N_18859,N_14659);
xnor U21485 (N_21485,N_15140,N_12532);
or U21486 (N_21486,N_19439,N_14465);
or U21487 (N_21487,N_16131,N_15178);
xor U21488 (N_21488,N_14583,N_13766);
or U21489 (N_21489,N_17050,N_14223);
or U21490 (N_21490,N_19225,N_14179);
and U21491 (N_21491,N_16706,N_11653);
or U21492 (N_21492,N_15300,N_18144);
nor U21493 (N_21493,N_14016,N_17872);
xnor U21494 (N_21494,N_13382,N_11729);
xnor U21495 (N_21495,N_19263,N_16774);
and U21496 (N_21496,N_19303,N_14111);
nand U21497 (N_21497,N_17452,N_16529);
nand U21498 (N_21498,N_10345,N_11935);
nand U21499 (N_21499,N_13538,N_19465);
xor U21500 (N_21500,N_11879,N_17479);
nor U21501 (N_21501,N_14357,N_17376);
and U21502 (N_21502,N_12269,N_18398);
or U21503 (N_21503,N_11076,N_11940);
or U21504 (N_21504,N_19699,N_14209);
xnor U21505 (N_21505,N_14887,N_10056);
or U21506 (N_21506,N_15647,N_12396);
nand U21507 (N_21507,N_12064,N_11689);
or U21508 (N_21508,N_13222,N_18680);
nand U21509 (N_21509,N_10720,N_19792);
and U21510 (N_21510,N_17415,N_19223);
and U21511 (N_21511,N_12475,N_10511);
nor U21512 (N_21512,N_11222,N_10429);
nor U21513 (N_21513,N_13145,N_16320);
nand U21514 (N_21514,N_13750,N_17955);
or U21515 (N_21515,N_17381,N_13000);
xnor U21516 (N_21516,N_18288,N_10305);
nand U21517 (N_21517,N_13045,N_11291);
or U21518 (N_21518,N_11715,N_12371);
or U21519 (N_21519,N_13862,N_15669);
nor U21520 (N_21520,N_17268,N_15615);
or U21521 (N_21521,N_17562,N_11488);
xor U21522 (N_21522,N_10994,N_17903);
nor U21523 (N_21523,N_19179,N_16501);
xor U21524 (N_21524,N_10107,N_12083);
nand U21525 (N_21525,N_10175,N_12809);
xnor U21526 (N_21526,N_11364,N_18468);
or U21527 (N_21527,N_14532,N_16512);
nor U21528 (N_21528,N_18054,N_13903);
nor U21529 (N_21529,N_17266,N_15305);
or U21530 (N_21530,N_11748,N_13395);
xnor U21531 (N_21531,N_19637,N_19752);
xor U21532 (N_21532,N_15605,N_10817);
or U21533 (N_21533,N_13679,N_14187);
xor U21534 (N_21534,N_19890,N_12383);
and U21535 (N_21535,N_18703,N_17859);
xor U21536 (N_21536,N_13363,N_15800);
and U21537 (N_21537,N_12521,N_15525);
xor U21538 (N_21538,N_18903,N_16787);
or U21539 (N_21539,N_14366,N_10367);
nand U21540 (N_21540,N_18303,N_16278);
and U21541 (N_21541,N_10125,N_18269);
or U21542 (N_21542,N_12369,N_18328);
or U21543 (N_21543,N_11537,N_10514);
nor U21544 (N_21544,N_12822,N_12733);
or U21545 (N_21545,N_15871,N_10762);
xnor U21546 (N_21546,N_10786,N_13438);
and U21547 (N_21547,N_16342,N_15996);
nor U21548 (N_21548,N_12039,N_19971);
xnor U21549 (N_21549,N_11378,N_10682);
nand U21550 (N_21550,N_19532,N_15299);
nand U21551 (N_21551,N_10826,N_17527);
nand U21552 (N_21552,N_19948,N_11303);
nor U21553 (N_21553,N_10573,N_10255);
xnor U21554 (N_21554,N_16911,N_14920);
nor U21555 (N_21555,N_15913,N_16640);
nor U21556 (N_21556,N_18340,N_12130);
nor U21557 (N_21557,N_11882,N_10946);
xor U21558 (N_21558,N_14601,N_19153);
nand U21559 (N_21559,N_19210,N_11402);
xnor U21560 (N_21560,N_12929,N_11722);
nand U21561 (N_21561,N_18960,N_18104);
or U21562 (N_21562,N_19587,N_11268);
xnor U21563 (N_21563,N_11740,N_15631);
and U21564 (N_21564,N_10307,N_14785);
nand U21565 (N_21565,N_10892,N_10032);
or U21566 (N_21566,N_17619,N_16948);
or U21567 (N_21567,N_10537,N_16234);
nor U21568 (N_21568,N_15036,N_13756);
nand U21569 (N_21569,N_12609,N_10595);
nand U21570 (N_21570,N_19381,N_10710);
and U21571 (N_21571,N_10306,N_19416);
or U21572 (N_21572,N_10231,N_13360);
nand U21573 (N_21573,N_19099,N_11497);
and U21574 (N_21574,N_10552,N_19937);
nand U21575 (N_21575,N_17597,N_11453);
nand U21576 (N_21576,N_11343,N_13990);
or U21577 (N_21577,N_14226,N_18517);
or U21578 (N_21578,N_13446,N_16298);
nand U21579 (N_21579,N_11171,N_13831);
nor U21580 (N_21580,N_10891,N_18875);
or U21581 (N_21581,N_18749,N_11646);
or U21582 (N_21582,N_19035,N_17963);
xnor U21583 (N_21583,N_12389,N_13337);
and U21584 (N_21584,N_10336,N_10396);
xnor U21585 (N_21585,N_12173,N_14711);
nor U21586 (N_21586,N_13985,N_10148);
nor U21587 (N_21587,N_18757,N_11463);
nor U21588 (N_21588,N_18334,N_18671);
xnor U21589 (N_21589,N_15232,N_18404);
xor U21590 (N_21590,N_12600,N_15452);
xnor U21591 (N_21591,N_14574,N_18447);
nor U21592 (N_21592,N_18184,N_11145);
or U21593 (N_21593,N_14214,N_16601);
nand U21594 (N_21594,N_13570,N_11281);
nand U21595 (N_21595,N_18786,N_12075);
nand U21596 (N_21596,N_11135,N_11635);
or U21597 (N_21597,N_16566,N_19299);
or U21598 (N_21598,N_17906,N_11032);
xnor U21599 (N_21599,N_15169,N_11691);
nor U21600 (N_21600,N_13590,N_14350);
xnor U21601 (N_21601,N_10512,N_15463);
or U21602 (N_21602,N_15642,N_18818);
nor U21603 (N_21603,N_12838,N_19795);
or U21604 (N_21604,N_16054,N_12315);
and U21605 (N_21605,N_10871,N_18108);
xor U21606 (N_21606,N_15397,N_18461);
and U21607 (N_21607,N_13506,N_12720);
nand U21608 (N_21608,N_18986,N_12398);
nor U21609 (N_21609,N_12122,N_13120);
nand U21610 (N_21610,N_15073,N_19468);
nor U21611 (N_21611,N_19671,N_16919);
nor U21612 (N_21612,N_10568,N_11501);
xnor U21613 (N_21613,N_13250,N_16096);
and U21614 (N_21614,N_12989,N_15080);
or U21615 (N_21615,N_16302,N_17817);
xnor U21616 (N_21616,N_10166,N_17354);
or U21617 (N_21617,N_10288,N_10670);
nand U21618 (N_21618,N_12623,N_11975);
and U21619 (N_21619,N_18373,N_15761);
nand U21620 (N_21620,N_14511,N_18178);
and U21621 (N_21621,N_17621,N_12859);
xor U21622 (N_21622,N_16958,N_10560);
xnor U21623 (N_21623,N_16332,N_12840);
nor U21624 (N_21624,N_15928,N_18429);
xor U21625 (N_21625,N_19794,N_13764);
and U21626 (N_21626,N_19636,N_12736);
xnor U21627 (N_21627,N_18142,N_12046);
nand U21628 (N_21628,N_12250,N_17751);
nor U21629 (N_21629,N_19781,N_13234);
nor U21630 (N_21630,N_17425,N_15133);
nor U21631 (N_21631,N_13282,N_11742);
xnor U21632 (N_21632,N_11191,N_18918);
nand U21633 (N_21633,N_18843,N_16811);
and U21634 (N_21634,N_17353,N_17505);
nor U21635 (N_21635,N_13095,N_12529);
xor U21636 (N_21636,N_19547,N_15168);
or U21637 (N_21637,N_16505,N_15191);
or U21638 (N_21638,N_18549,N_13046);
nand U21639 (N_21639,N_16515,N_17331);
nor U21640 (N_21640,N_11894,N_17563);
nand U21641 (N_21641,N_12261,N_17130);
nand U21642 (N_21642,N_17565,N_11339);
nor U21643 (N_21643,N_13720,N_19912);
xnor U21644 (N_21644,N_18711,N_17080);
and U21645 (N_21645,N_12073,N_16658);
nand U21646 (N_21646,N_10996,N_16017);
nor U21647 (N_21647,N_19049,N_10662);
and U21648 (N_21648,N_10825,N_11933);
or U21649 (N_21649,N_13197,N_11358);
and U21650 (N_21650,N_17040,N_16565);
xnor U21651 (N_21651,N_16334,N_11138);
nor U21652 (N_21652,N_14648,N_16226);
xnor U21653 (N_21653,N_19690,N_18177);
or U21654 (N_21654,N_18662,N_11065);
nand U21655 (N_21655,N_12326,N_15789);
and U21656 (N_21656,N_12601,N_18873);
or U21657 (N_21657,N_12274,N_15117);
nor U21658 (N_21658,N_19660,N_12923);
and U21659 (N_21659,N_19403,N_17323);
or U21660 (N_21660,N_12678,N_10427);
or U21661 (N_21661,N_10579,N_16624);
or U21662 (N_21662,N_18883,N_12901);
nor U21663 (N_21663,N_13710,N_12426);
xor U21664 (N_21664,N_15810,N_17198);
and U21665 (N_21665,N_14286,N_13391);
nand U21666 (N_21666,N_19088,N_16785);
nand U21667 (N_21667,N_13036,N_17731);
and U21668 (N_21668,N_13963,N_15060);
or U21669 (N_21669,N_11658,N_13032);
or U21670 (N_21670,N_12681,N_18030);
and U21671 (N_21671,N_13842,N_18782);
xor U21672 (N_21672,N_10698,N_11085);
nand U21673 (N_21673,N_10993,N_15951);
or U21674 (N_21674,N_13703,N_16491);
nor U21675 (N_21675,N_14692,N_10365);
nand U21676 (N_21676,N_17338,N_12180);
nand U21677 (N_21677,N_10187,N_19810);
and U21678 (N_21678,N_16021,N_11845);
and U21679 (N_21679,N_15416,N_12732);
nor U21680 (N_21680,N_10711,N_16656);
nor U21681 (N_21681,N_10200,N_11384);
nand U21682 (N_21682,N_18205,N_11269);
and U21683 (N_21683,N_15884,N_12748);
nor U21684 (N_21684,N_19264,N_18636);
nor U21685 (N_21685,N_12597,N_10857);
or U21686 (N_21686,N_19533,N_16219);
nor U21687 (N_21687,N_12579,N_12936);
or U21688 (N_21688,N_14536,N_11208);
or U21689 (N_21689,N_19435,N_17662);
nor U21690 (N_21690,N_18872,N_11955);
and U21691 (N_21691,N_15535,N_10616);
nand U21692 (N_21692,N_18135,N_15752);
and U21693 (N_21693,N_19680,N_15912);
nor U21694 (N_21694,N_15435,N_19391);
xnor U21695 (N_21695,N_13574,N_12801);
nand U21696 (N_21696,N_11579,N_14074);
nand U21697 (N_21697,N_10263,N_12663);
xor U21698 (N_21698,N_12995,N_14737);
nor U21699 (N_21699,N_17140,N_16330);
or U21700 (N_21700,N_14753,N_11555);
nand U21701 (N_21701,N_11166,N_13173);
nand U21702 (N_21702,N_19796,N_10061);
nand U21703 (N_21703,N_14523,N_17334);
or U21704 (N_21704,N_13863,N_16519);
and U21705 (N_21705,N_11944,N_17245);
nand U21706 (N_21706,N_11458,N_13835);
nand U21707 (N_21707,N_19016,N_11544);
and U21708 (N_21708,N_18825,N_11260);
and U21709 (N_21709,N_12621,N_17402);
and U21710 (N_21710,N_16232,N_14809);
or U21711 (N_21711,N_18366,N_14083);
xnor U21712 (N_21712,N_19417,N_19813);
nor U21713 (N_21713,N_11612,N_18759);
nor U21714 (N_21714,N_14365,N_10695);
nand U21715 (N_21715,N_16295,N_15338);
and U21716 (N_21716,N_12227,N_16312);
nor U21717 (N_21717,N_14110,N_15888);
nor U21718 (N_21718,N_15354,N_11684);
nand U21719 (N_21719,N_14168,N_14933);
nand U21720 (N_21720,N_11996,N_14235);
or U21721 (N_21721,N_18378,N_11235);
or U21722 (N_21722,N_19858,N_13128);
nand U21723 (N_21723,N_12374,N_11838);
nor U21724 (N_21724,N_19631,N_10948);
nor U21725 (N_21725,N_19588,N_10323);
nor U21726 (N_21726,N_19411,N_17411);
or U21727 (N_21727,N_11994,N_16718);
and U21728 (N_21728,N_14786,N_18855);
xnor U21729 (N_21729,N_13109,N_15995);
nor U21730 (N_21730,N_12343,N_19520);
nor U21731 (N_21731,N_14414,N_18969);
xnor U21732 (N_21732,N_19643,N_19550);
or U21733 (N_21733,N_16074,N_19826);
xnor U21734 (N_21734,N_10406,N_16220);
nand U21735 (N_21735,N_13478,N_13653);
xnor U21736 (N_21736,N_16416,N_11155);
xnor U21737 (N_21737,N_16636,N_13573);
and U21738 (N_21738,N_12110,N_15203);
nand U21739 (N_21739,N_16150,N_14324);
and U21740 (N_21740,N_12134,N_14163);
and U21741 (N_21741,N_19199,N_13359);
nand U21742 (N_21742,N_11279,N_19545);
or U21743 (N_21743,N_11904,N_17063);
nand U21744 (N_21744,N_13568,N_14189);
xnor U21745 (N_21745,N_18919,N_19956);
xor U21746 (N_21746,N_14048,N_12786);
or U21747 (N_21747,N_10020,N_14684);
xnor U21748 (N_21748,N_14700,N_19973);
and U21749 (N_21749,N_11121,N_15929);
nor U21750 (N_21750,N_13634,N_17071);
nand U21751 (N_21751,N_18096,N_12554);
nor U21752 (N_21752,N_14094,N_16728);
and U21753 (N_21753,N_13392,N_11075);
nor U21754 (N_21754,N_12194,N_16367);
nand U21755 (N_21755,N_17252,N_16929);
nand U21756 (N_21756,N_18829,N_19279);
nor U21757 (N_21757,N_15969,N_11283);
nor U21758 (N_21758,N_16387,N_19849);
and U21759 (N_21759,N_14472,N_18506);
xor U21760 (N_21760,N_10274,N_16043);
and U21761 (N_21761,N_13287,N_17284);
nor U21762 (N_21762,N_16943,N_16499);
nand U21763 (N_21763,N_14871,N_17172);
and U21764 (N_21764,N_18204,N_13777);
and U21765 (N_21765,N_17309,N_17940);
nor U21766 (N_21766,N_16065,N_12514);
nor U21767 (N_21767,N_19728,N_11009);
and U21768 (N_21768,N_11733,N_16055);
nor U21769 (N_21769,N_12335,N_14456);
and U21770 (N_21770,N_13662,N_13802);
xor U21771 (N_21771,N_17540,N_10885);
nand U21772 (N_21772,N_11404,N_15834);
or U21773 (N_21773,N_16627,N_11875);
nand U21774 (N_21774,N_11345,N_14381);
and U21775 (N_21775,N_17300,N_11710);
nand U21776 (N_21776,N_10574,N_12433);
nor U21777 (N_21777,N_18301,N_16354);
and U21778 (N_21778,N_17432,N_19089);
xor U21779 (N_21779,N_11958,N_15926);
and U21780 (N_21780,N_11954,N_13880);
and U21781 (N_21781,N_15195,N_13663);
or U21782 (N_21782,N_12852,N_14442);
nor U21783 (N_21783,N_16391,N_16264);
xnor U21784 (N_21784,N_18337,N_12902);
xnor U21785 (N_21785,N_13315,N_14621);
and U21786 (N_21786,N_17607,N_12028);
nand U21787 (N_21787,N_11013,N_18148);
or U21788 (N_21788,N_19462,N_19147);
xnor U21789 (N_21789,N_15738,N_17768);
and U21790 (N_21790,N_16251,N_14881);
nand U21791 (N_21791,N_17781,N_10658);
nor U21792 (N_21792,N_18634,N_18489);
or U21793 (N_21793,N_14281,N_18707);
or U21794 (N_21794,N_10838,N_14182);
nor U21795 (N_21795,N_19178,N_19505);
nand U21796 (N_21796,N_15064,N_16886);
xor U21797 (N_21797,N_13935,N_19913);
nand U21798 (N_21798,N_13542,N_14610);
and U21799 (N_21799,N_13023,N_16383);
or U21800 (N_21800,N_14199,N_16703);
nor U21801 (N_21801,N_13770,N_11031);
and U21802 (N_21802,N_14596,N_19115);
nor U21803 (N_21803,N_10667,N_18739);
nor U21804 (N_21804,N_13791,N_15938);
xor U21805 (N_21805,N_18412,N_19525);
and U21806 (N_21806,N_13960,N_11481);
nor U21807 (N_21807,N_18921,N_13106);
and U21808 (N_21808,N_15475,N_18213);
and U21809 (N_21809,N_13335,N_16951);
and U21810 (N_21810,N_16835,N_10350);
nor U21811 (N_21811,N_10663,N_14416);
nor U21812 (N_21812,N_19068,N_16478);
nand U21813 (N_21813,N_13038,N_11811);
xnor U21814 (N_21814,N_18392,N_12474);
nor U21815 (N_21815,N_14987,N_19936);
nand U21816 (N_21816,N_11111,N_11583);
and U21817 (N_21817,N_11239,N_18143);
nand U21818 (N_21818,N_18103,N_18342);
nand U21819 (N_21819,N_16214,N_17555);
xnor U21820 (N_21820,N_18755,N_12798);
or U21821 (N_21821,N_16468,N_15083);
nor U21822 (N_21822,N_16693,N_11472);
and U21823 (N_21823,N_10664,N_14224);
nand U21824 (N_21824,N_16558,N_16670);
nor U21825 (N_21825,N_13275,N_14039);
or U21826 (N_21826,N_14036,N_19727);
nand U21827 (N_21827,N_17997,N_18593);
and U21828 (N_21828,N_15018,N_16258);
nor U21829 (N_21829,N_19501,N_12307);
xor U21830 (N_21830,N_18862,N_16469);
and U21831 (N_21831,N_15404,N_11249);
and U21832 (N_21832,N_14326,N_13688);
xor U21833 (N_21833,N_15415,N_18776);
xnor U21834 (N_21834,N_16833,N_10848);
and U21835 (N_21835,N_16132,N_14213);
and U21836 (N_21836,N_14154,N_17400);
nor U21837 (N_21837,N_17009,N_14061);
or U21838 (N_21838,N_10587,N_10528);
or U21839 (N_21839,N_12629,N_17653);
or U21840 (N_21840,N_13449,N_17711);
or U21841 (N_21841,N_10928,N_10265);
xor U21842 (N_21842,N_18870,N_17891);
and U21843 (N_21843,N_11863,N_12795);
nand U21844 (N_21844,N_13182,N_10625);
nor U21845 (N_21845,N_17288,N_15991);
nor U21846 (N_21846,N_19400,N_14447);
nor U21847 (N_21847,N_16779,N_10830);
and U21848 (N_21848,N_16009,N_17930);
xor U21849 (N_21849,N_15220,N_15267);
and U21850 (N_21850,N_11202,N_16651);
nor U21851 (N_21851,N_18032,N_14723);
or U21852 (N_21852,N_13284,N_16769);
xnor U21853 (N_21853,N_16160,N_11049);
xnor U21854 (N_21854,N_13588,N_19843);
and U21855 (N_21855,N_18880,N_12385);
nor U21856 (N_21856,N_16427,N_19564);
xor U21857 (N_21857,N_12669,N_18374);
xor U21858 (N_21858,N_14988,N_12183);
xnor U21859 (N_21859,N_17472,N_14961);
nor U21860 (N_21860,N_19526,N_19842);
and U21861 (N_21861,N_14729,N_11159);
nor U21862 (N_21862,N_18632,N_18076);
nand U21863 (N_21863,N_14229,N_16041);
nand U21864 (N_21864,N_13651,N_13867);
or U21865 (N_21865,N_11959,N_15038);
or U21866 (N_21866,N_13349,N_18180);
and U21867 (N_21867,N_11027,N_19494);
or U21868 (N_21868,N_16164,N_13737);
nor U21869 (N_21869,N_19747,N_12375);
and U21870 (N_21870,N_19865,N_17948);
nor U21871 (N_21871,N_19045,N_17392);
xor U21872 (N_21872,N_16411,N_14701);
nand U21873 (N_21873,N_13549,N_14579);
xor U21874 (N_21874,N_13413,N_16276);
nand U21875 (N_21875,N_13016,N_18262);
or U21876 (N_21876,N_13122,N_10215);
nor U21877 (N_21877,N_16537,N_10945);
nand U21878 (N_21878,N_10906,N_10143);
nand U21879 (N_21879,N_10589,N_11329);
nand U21880 (N_21880,N_12150,N_13495);
nand U21881 (N_21881,N_17874,N_15930);
xnor U21882 (N_21882,N_19470,N_17551);
nand U21883 (N_21883,N_15249,N_19278);
and U21884 (N_21884,N_18556,N_12644);
xor U21885 (N_21885,N_19335,N_19806);
nand U21886 (N_21886,N_19512,N_10329);
nor U21887 (N_21887,N_15425,N_15179);
and U21888 (N_21888,N_13133,N_16490);
or U21889 (N_21889,N_17783,N_16100);
or U21890 (N_21890,N_18239,N_17881);
nand U21891 (N_21891,N_10561,N_18913);
and U21892 (N_21892,N_13431,N_11603);
nand U21893 (N_21893,N_14113,N_13003);
and U21894 (N_21894,N_15394,N_19725);
nor U21895 (N_21895,N_10316,N_15260);
and U21896 (N_21896,N_14689,N_19949);
nand U21897 (N_21897,N_15099,N_12741);
or U21898 (N_21898,N_18620,N_10059);
or U21899 (N_21899,N_12808,N_11617);
nor U21900 (N_21900,N_19553,N_14469);
or U21901 (N_21901,N_17469,N_12513);
and U21902 (N_21902,N_10428,N_19483);
xor U21903 (N_21903,N_12622,N_15164);
nor U21904 (N_21904,N_10558,N_14943);
or U21905 (N_21905,N_11595,N_12459);
and U21906 (N_21906,N_12469,N_10201);
nand U21907 (N_21907,N_19619,N_13512);
xnor U21908 (N_21908,N_15828,N_14763);
xnor U21909 (N_21909,N_16530,N_18605);
nand U21910 (N_21910,N_14320,N_13299);
or U21911 (N_21911,N_15152,N_19580);
and U21912 (N_21912,N_16472,N_17813);
or U21913 (N_21913,N_13575,N_19015);
xnor U21914 (N_21914,N_16169,N_16146);
nor U21915 (N_21915,N_14801,N_17902);
or U21916 (N_21916,N_16327,N_12342);
or U21917 (N_21917,N_17691,N_18234);
xnor U21918 (N_21918,N_17066,N_19529);
or U21919 (N_21919,N_15916,N_13423);
or U21920 (N_21920,N_19175,N_18713);
or U21921 (N_21921,N_12715,N_10279);
nand U21922 (N_21922,N_16748,N_15110);
or U21923 (N_21923,N_15721,N_11973);
and U21924 (N_21924,N_10726,N_19939);
or U21925 (N_21925,N_16386,N_16481);
nand U21926 (N_21926,N_14937,N_16710);
or U21927 (N_21927,N_18036,N_10959);
nor U21928 (N_21928,N_10292,N_16540);
and U21929 (N_21929,N_11336,N_18215);
and U21930 (N_21930,N_15453,N_12185);
nor U21931 (N_21931,N_12191,N_17577);
xor U21932 (N_21932,N_14653,N_12476);
and U21933 (N_21933,N_14633,N_10694);
or U21934 (N_21934,N_13168,N_13501);
nand U21935 (N_21935,N_14936,N_11142);
nor U21936 (N_21936,N_17373,N_11099);
and U21937 (N_21937,N_17492,N_18445);
or U21938 (N_21938,N_10376,N_14486);
nand U21939 (N_21939,N_15659,N_12536);
nor U21940 (N_21940,N_14140,N_16942);
or U21941 (N_21941,N_13771,N_13479);
nor U21942 (N_21942,N_15795,N_11466);
or U21943 (N_21943,N_13648,N_10463);
xnor U21944 (N_21944,N_11562,N_18800);
and U21945 (N_21945,N_14051,N_14503);
or U21946 (N_21946,N_10120,N_11310);
nor U21947 (N_21947,N_18397,N_14939);
or U21948 (N_21948,N_14143,N_14084);
or U21949 (N_21949,N_18266,N_12952);
nand U21950 (N_21950,N_13948,N_13712);
nor U21951 (N_21951,N_19661,N_18917);
xor U21952 (N_21952,N_14455,N_19373);
nand U21953 (N_21953,N_15506,N_16824);
xnor U21954 (N_21954,N_16425,N_11647);
and U21955 (N_21955,N_11730,N_19378);
or U21956 (N_21956,N_15867,N_14407);
nor U21957 (N_21957,N_18907,N_19217);
nor U21958 (N_21958,N_11106,N_11132);
xnor U21959 (N_21959,N_12408,N_19398);
and U21960 (N_21960,N_17028,N_18717);
nor U21961 (N_21961,N_11126,N_12924);
or U21962 (N_21962,N_18155,N_15596);
xnor U21963 (N_21963,N_15514,N_10997);
or U21964 (N_21964,N_15269,N_13073);
nand U21965 (N_21965,N_10101,N_13896);
nor U21966 (N_21966,N_10036,N_13827);
nand U21967 (N_21967,N_18820,N_18935);
xor U21968 (N_21968,N_10846,N_12750);
xnor U21969 (N_21969,N_18123,N_17142);
and U21970 (N_21970,N_18084,N_13442);
or U21971 (N_21971,N_16964,N_11897);
nor U21972 (N_21972,N_11876,N_19120);
or U21973 (N_21973,N_17849,N_14031);
and U21974 (N_21974,N_16837,N_15754);
or U21975 (N_21975,N_18344,N_10816);
xor U21976 (N_21976,N_18210,N_11926);
nand U21977 (N_21977,N_12393,N_15777);
or U21978 (N_21978,N_17734,N_18635);
xnor U21979 (N_21979,N_19157,N_12552);
nor U21980 (N_21980,N_15335,N_11311);
nand U21981 (N_21981,N_15780,N_11187);
nor U21982 (N_21982,N_14150,N_19048);
nand U21983 (N_21983,N_14345,N_15694);
and U21984 (N_21984,N_11331,N_17131);
or U21985 (N_21985,N_11498,N_16901);
nor U21986 (N_21986,N_10132,N_12021);
and U21987 (N_21987,N_10819,N_13623);
and U21988 (N_21988,N_15406,N_12357);
and U21989 (N_21989,N_11180,N_17574);
xnor U21990 (N_21990,N_13096,N_18799);
xnor U21991 (N_21991,N_13658,N_13494);
and U21992 (N_21992,N_18640,N_12639);
nor U21993 (N_21993,N_15576,N_14921);
nor U21994 (N_21994,N_10543,N_14438);
nor U21995 (N_21995,N_12008,N_19349);
nor U21996 (N_21996,N_10138,N_15703);
or U21997 (N_21997,N_11663,N_15860);
nor U21998 (N_21998,N_15823,N_13160);
nand U21999 (N_21999,N_17998,N_16663);
nor U22000 (N_22000,N_18427,N_15875);
nand U22001 (N_22001,N_13228,N_17251);
xnor U22002 (N_22002,N_14658,N_18932);
nand U22003 (N_22003,N_17502,N_19364);
nand U22004 (N_22004,N_15792,N_17366);
nand U22005 (N_22005,N_11626,N_11251);
nor U22006 (N_22006,N_15908,N_13114);
nor U22007 (N_22007,N_18576,N_18712);
or U22008 (N_22008,N_15473,N_14194);
nor U22009 (N_22009,N_12147,N_11354);
nor U22010 (N_22010,N_14360,N_15364);
nor U22011 (N_22011,N_12796,N_11554);
nand U22012 (N_22012,N_16475,N_12618);
and U22013 (N_22013,N_12233,N_12785);
or U22014 (N_22014,N_13544,N_15256);
nand U22015 (N_22015,N_10473,N_12001);
nand U22016 (N_22016,N_10205,N_11941);
nor U22017 (N_22017,N_13158,N_17001);
and U22018 (N_22018,N_14007,N_12172);
nor U22019 (N_22019,N_15827,N_11686);
xor U22020 (N_22020,N_12559,N_14537);
nand U22021 (N_22021,N_15366,N_11298);
or U22022 (N_22022,N_16965,N_13490);
xor U22023 (N_22023,N_11835,N_18074);
nor U22024 (N_22024,N_10828,N_16003);
nand U22025 (N_22025,N_18147,N_12760);
nand U22026 (N_22026,N_16238,N_16484);
nor U22027 (N_22027,N_13729,N_19759);
nand U22028 (N_22028,N_12907,N_15015);
and U22029 (N_22029,N_17939,N_12301);
nand U22030 (N_22030,N_11479,N_15037);
xnor U22031 (N_22031,N_17965,N_16309);
xnor U22032 (N_22032,N_16760,N_13702);
nand U22033 (N_22033,N_15999,N_16652);
nor U22034 (N_22034,N_13839,N_15695);
nand U22035 (N_22035,N_16027,N_15346);
xnor U22036 (N_22036,N_13187,N_11152);
or U22037 (N_22037,N_13869,N_11883);
xnor U22038 (N_22038,N_14666,N_12654);
or U22039 (N_22039,N_11673,N_13941);
xor U22040 (N_22040,N_19804,N_12391);
nor U22041 (N_22041,N_14595,N_12564);
nand U22042 (N_22042,N_18777,N_13714);
nand U22043 (N_22043,N_12418,N_13410);
nor U22044 (N_22044,N_10780,N_13235);
nand U22045 (N_22045,N_12677,N_13502);
xnor U22046 (N_22046,N_14153,N_13203);
xor U22047 (N_22047,N_10050,N_12899);
or U22048 (N_22048,N_13123,N_16254);
nand U22049 (N_22049,N_10487,N_18970);
nor U22050 (N_22050,N_10083,N_16695);
nand U22051 (N_22051,N_13041,N_16045);
or U22052 (N_22052,N_12399,N_11570);
or U22053 (N_22053,N_16506,N_18130);
nor U22054 (N_22054,N_18027,N_12423);
xnor U22055 (N_22055,N_14956,N_19212);
and U22056 (N_22056,N_14664,N_14768);
nor U22057 (N_22057,N_17681,N_15822);
or U22058 (N_22058,N_13314,N_17816);
xnor U22059 (N_22059,N_16445,N_14963);
nand U22060 (N_22060,N_13612,N_10624);
xnor U22061 (N_22061,N_18860,N_18705);
nor U22062 (N_22062,N_18979,N_10672);
and U22063 (N_22063,N_17456,N_13821);
and U22064 (N_22064,N_11949,N_19285);
or U22065 (N_22065,N_11512,N_15638);
and U22066 (N_22066,N_10016,N_13800);
and U22067 (N_22067,N_13063,N_19384);
or U22068 (N_22068,N_15255,N_12949);
nor U22069 (N_22069,N_17947,N_17807);
nand U22070 (N_22070,N_14612,N_14103);
or U22071 (N_22071,N_18140,N_18892);
xor U22072 (N_22072,N_10419,N_17272);
xnor U22073 (N_22073,N_17834,N_14707);
nor U22074 (N_22074,N_11541,N_14829);
xnor U22075 (N_22075,N_14812,N_10142);
nor U22076 (N_22076,N_13815,N_10687);
or U22077 (N_22077,N_16872,N_13426);
nand U22078 (N_22078,N_10590,N_18185);
nor U22079 (N_22079,N_11429,N_14493);
or U22080 (N_22080,N_19864,N_16542);
nor U22081 (N_22081,N_12518,N_17192);
xor U22082 (N_22082,N_18710,N_18284);
nor U22083 (N_22083,N_18042,N_16974);
or U22084 (N_22084,N_15618,N_13237);
nand U22085 (N_22085,N_12905,N_18781);
and U22086 (N_22086,N_10327,N_11233);
or U22087 (N_22087,N_12782,N_16532);
xnor U22088 (N_22088,N_15207,N_15010);
xnor U22089 (N_22089,N_14373,N_16002);
nand U22090 (N_22090,N_15268,N_16900);
nor U22091 (N_22091,N_11774,N_11988);
and U22092 (N_22092,N_19220,N_11137);
xor U22093 (N_22093,N_16966,N_15645);
nand U22094 (N_22094,N_15863,N_16184);
xor U22095 (N_22095,N_16857,N_19076);
xor U22096 (N_22096,N_14361,N_17683);
or U22097 (N_22097,N_10864,N_10596);
nand U22098 (N_22098,N_13543,N_10282);
xnor U22099 (N_22099,N_19999,N_17235);
xnor U22100 (N_22100,N_14507,N_19228);
nor U22101 (N_22101,N_13582,N_13817);
nor U22102 (N_22102,N_17193,N_16525);
nand U22103 (N_22103,N_12205,N_19878);
xnor U22104 (N_22104,N_19491,N_19785);
xor U22105 (N_22105,N_15242,N_11350);
nor U22106 (N_22106,N_13665,N_18775);
nand U22107 (N_22107,N_15396,N_19257);
nand U22108 (N_22108,N_18212,N_13973);
xor U22109 (N_22109,N_12149,N_18257);
and U22110 (N_22110,N_16801,N_18612);
xor U22111 (N_22111,N_11203,N_15131);
or U22112 (N_22112,N_14584,N_12602);
nor U22113 (N_22113,N_17247,N_12267);
nor U22114 (N_22114,N_14843,N_11426);
nand U22115 (N_22115,N_11386,N_13389);
xor U22116 (N_22116,N_15361,N_19449);
xnor U22117 (N_22117,N_14859,N_16382);
or U22118 (N_22118,N_13788,N_10529);
nand U22119 (N_22119,N_12050,N_12696);
or U22120 (N_22120,N_14476,N_15656);
nor U22121 (N_22121,N_16172,N_15874);
xnor U22122 (N_22122,N_17635,N_10012);
nor U22123 (N_22123,N_11353,N_11592);
xor U22124 (N_22124,N_16691,N_17027);
nand U22125 (N_22125,N_12249,N_12511);
nor U22126 (N_22126,N_10608,N_11403);
nor U22127 (N_22127,N_10208,N_18493);
xnor U22128 (N_22128,N_14091,N_11061);
and U22129 (N_22129,N_18752,N_19084);
xnor U22130 (N_22130,N_10965,N_18729);
xor U22131 (N_22131,N_11278,N_10474);
nor U22132 (N_22132,N_16875,N_10038);
xor U22133 (N_22133,N_13640,N_19310);
nor U22134 (N_22134,N_16850,N_19042);
or U22135 (N_22135,N_18984,N_11225);
nor U22136 (N_22136,N_10749,N_10346);
or U22137 (N_22137,N_11736,N_17367);
nand U22138 (N_22138,N_13332,N_10707);
or U22139 (N_22139,N_15159,N_17547);
nand U22140 (N_22140,N_11850,N_17609);
and U22141 (N_22141,N_14706,N_19320);
nor U22142 (N_22142,N_19114,N_18788);
nor U22143 (N_22143,N_11127,N_18277);
and U22144 (N_22144,N_13966,N_14757);
or U22145 (N_22145,N_18585,N_19065);
xor U22146 (N_22146,N_10436,N_18001);
xnor U22147 (N_22147,N_14260,N_11782);
nor U22148 (N_22148,N_16586,N_18202);
xnor U22149 (N_22149,N_14787,N_18539);
nor U22150 (N_22150,N_18922,N_18354);
nand U22151 (N_22151,N_10420,N_19691);
nand U22152 (N_22152,N_18230,N_15410);
nor U22153 (N_22153,N_12543,N_17595);
xor U22154 (N_22154,N_11109,N_19782);
or U22155 (N_22155,N_19693,N_12361);
and U22156 (N_22156,N_12577,N_15281);
nand U22157 (N_22157,N_18183,N_11471);
and U22158 (N_22158,N_19159,N_18216);
nor U22159 (N_22159,N_15628,N_18388);
and U22160 (N_22160,N_11444,N_16197);
nand U22161 (N_22161,N_16457,N_13637);
or U22162 (N_22162,N_14593,N_12452);
or U22163 (N_22163,N_10779,N_11987);
and U22164 (N_22164,N_11797,N_11970);
and U22165 (N_22165,N_18292,N_19698);
and U22166 (N_22166,N_14765,N_19965);
nor U22167 (N_22167,N_16864,N_17488);
or U22168 (N_22168,N_16753,N_17097);
nand U22169 (N_22169,N_15579,N_19389);
xor U22170 (N_22170,N_15812,N_12132);
xnor U22171 (N_22171,N_10113,N_17920);
nand U22172 (N_22172,N_11734,N_12596);
and U22173 (N_22173,N_16353,N_10453);
nand U22174 (N_22174,N_13002,N_13024);
and U22175 (N_22175,N_12481,N_15474);
nor U22176 (N_22176,N_11804,N_11296);
nor U22177 (N_22177,N_17238,N_17036);
nor U22178 (N_22178,N_15687,N_18335);
xor U22179 (N_22179,N_19189,N_11229);
or U22180 (N_22180,N_11937,N_19315);
or U22181 (N_22181,N_17578,N_19898);
xnor U22182 (N_22182,N_10822,N_13361);
xnor U22183 (N_22183,N_19128,N_10793);
or U22184 (N_22184,N_18815,N_11667);
or U22185 (N_22185,N_17820,N_10855);
or U22186 (N_22186,N_16539,N_10330);
or U22187 (N_22187,N_10705,N_19380);
or U22188 (N_22188,N_18220,N_19790);
or U22189 (N_22189,N_17418,N_19882);
nor U22190 (N_22190,N_19447,N_17899);
nor U22191 (N_22191,N_16229,N_15894);
xor U22192 (N_22192,N_12847,N_17470);
and U22193 (N_22193,N_18448,N_15215);
xor U22194 (N_22194,N_19780,N_13736);
and U22195 (N_22195,N_16385,N_18244);
xnor U22196 (N_22196,N_11584,N_17806);
nand U22197 (N_22197,N_13678,N_12290);
xnor U22198 (N_22198,N_19859,N_10077);
xor U22199 (N_22199,N_19055,N_13749);
or U22200 (N_22200,N_12799,N_17279);
nand U22201 (N_22201,N_19307,N_12047);
and U22202 (N_22202,N_14112,N_17221);
xor U22203 (N_22203,N_18044,N_18679);
and U22204 (N_22204,N_10929,N_16174);
or U22205 (N_22205,N_13587,N_18638);
and U22206 (N_22206,N_14431,N_18845);
nand U22207 (N_22207,N_12086,N_12450);
and U22208 (N_22208,N_18007,N_18587);
or U22209 (N_22209,N_13489,N_11196);
and U22210 (N_22210,N_16869,N_14782);
xnor U22211 (N_22211,N_12114,N_10915);
and U22212 (N_22212,N_14774,N_16362);
or U22213 (N_22213,N_14597,N_10222);
xor U22214 (N_22214,N_15793,N_19886);
and U22215 (N_22215,N_16470,N_15657);
or U22216 (N_22216,N_14437,N_18968);
nor U22217 (N_22217,N_12281,N_17926);
nand U22218 (N_22218,N_12775,N_14158);
and U22219 (N_22219,N_19195,N_18472);
nor U22220 (N_22220,N_14499,N_19164);
or U22221 (N_22221,N_11817,N_12067);
xor U22222 (N_22222,N_11385,N_15606);
or U22223 (N_22223,N_10395,N_18442);
or U22224 (N_22224,N_18079,N_18158);
xor U22225 (N_22225,N_11632,N_17168);
or U22226 (N_22226,N_16437,N_10133);
or U22227 (N_22227,N_19515,N_11966);
and U22228 (N_22228,N_11019,N_14050);
or U22229 (N_22229,N_15274,N_15198);
xnor U22230 (N_22230,N_14464,N_11158);
nor U22231 (N_22231,N_19437,N_11536);
and U22232 (N_22232,N_12694,N_11451);
and U22233 (N_22233,N_10834,N_14484);
nor U22234 (N_22234,N_14877,N_16455);
nor U22235 (N_22235,N_17483,N_14496);
nand U22236 (N_22236,N_13434,N_14385);
xnor U22237 (N_22237,N_18643,N_16390);
and U22238 (N_22238,N_13302,N_15981);
xor U22239 (N_22239,N_19603,N_17297);
and U22240 (N_22240,N_10665,N_17250);
nand U22241 (N_22241,N_16036,N_14371);
xnor U22242 (N_22242,N_18933,N_13794);
nand U22243 (N_22243,N_14805,N_12578);
nor U22244 (N_22244,N_11266,N_16750);
nand U22245 (N_22245,N_19940,N_16376);
and U22246 (N_22246,N_19474,N_18941);
and U22247 (N_22247,N_10523,N_17073);
xnor U22248 (N_22248,N_10299,N_17379);
or U22249 (N_22249,N_13691,N_12255);
and U22250 (N_22250,N_18533,N_12872);
xnor U22251 (N_22251,N_15289,N_10841);
nand U22252 (N_22252,N_17770,N_18015);
nor U22253 (N_22253,N_16882,N_16797);
nand U22254 (N_22254,N_12222,N_15353);
nand U22255 (N_22255,N_10455,N_13057);
xor U22256 (N_22256,N_13213,N_16124);
xor U22257 (N_22257,N_13753,N_10256);
or U22258 (N_22258,N_10702,N_12870);
xnor U22259 (N_22259,N_13954,N_14035);
and U22260 (N_22260,N_11178,N_10199);
nor U22261 (N_22261,N_10606,N_16171);
and U22262 (N_22262,N_14838,N_11618);
xnor U22263 (N_22263,N_10078,N_11943);
nand U22264 (N_22264,N_14487,N_12891);
and U22265 (N_22265,N_18737,N_17124);
xor U22266 (N_22266,N_12462,N_13428);
nand U22267 (N_22267,N_14618,N_17440);
nand U22268 (N_22268,N_14256,N_14823);
xnor U22269 (N_22269,N_12365,N_11780);
nand U22270 (N_22270,N_17070,N_14215);
or U22271 (N_22271,N_12541,N_15165);
nand U22272 (N_22272,N_17576,N_19033);
xnor U22273 (N_22273,N_11289,N_16033);
xnor U22274 (N_22274,N_11997,N_16536);
or U22275 (N_22275,N_10815,N_11485);
xor U22276 (N_22276,N_17308,N_16155);
or U22277 (N_22277,N_15661,N_13186);
nand U22278 (N_22278,N_12208,N_11324);
and U22279 (N_22279,N_10303,N_17990);
or U22280 (N_22280,N_10035,N_12648);
nor U22281 (N_22281,N_10788,N_15492);
xnor U22282 (N_22282,N_14139,N_12299);
and U22283 (N_22283,N_18563,N_18659);
or U22284 (N_22284,N_16397,N_10722);
and U22285 (N_22285,N_10797,N_19061);
nor U22286 (N_22286,N_14964,N_18689);
or U22287 (N_22287,N_18744,N_11631);
or U22288 (N_22288,N_14549,N_11084);
nand U22289 (N_22289,N_13061,N_10191);
nand U22290 (N_22290,N_18779,N_13521);
nor U22291 (N_22291,N_12802,N_18507);
nand U22292 (N_22292,N_10495,N_19521);
or U22293 (N_22293,N_11262,N_10025);
nand U22294 (N_22294,N_11455,N_12980);
nor U22295 (N_22295,N_16363,N_11026);
nand U22296 (N_22296,N_17074,N_13580);
or U22297 (N_22297,N_19920,N_14938);
nor U22298 (N_22298,N_15235,N_10238);
nor U22299 (N_22299,N_11625,N_13626);
xnor U22300 (N_22300,N_18715,N_18439);
and U22301 (N_22301,N_12379,N_14834);
and U22302 (N_22302,N_19187,N_19242);
and U22303 (N_22303,N_14274,N_13692);
xor U22304 (N_22304,N_13094,N_19184);
nor U22305 (N_22305,N_14662,N_14290);
or U22306 (N_22306,N_11564,N_16059);
nor U22307 (N_22307,N_17785,N_14080);
nor U22308 (N_22308,N_13552,N_14285);
or U22309 (N_22309,N_14634,N_15957);
nand U22310 (N_22310,N_12739,N_18250);
xnor U22311 (N_22311,N_19868,N_18206);
xnor U22312 (N_22312,N_15541,N_12776);
nand U22313 (N_22313,N_15505,N_15975);
nor U22314 (N_22314,N_17387,N_18754);
xor U22315 (N_22315,N_19980,N_12216);
nand U22316 (N_22316,N_15383,N_19566);
nor U22317 (N_22317,N_14276,N_12745);
xnor U22318 (N_22318,N_11100,N_11001);
xnor U22319 (N_22319,N_18962,N_16502);
or U22320 (N_22320,N_16346,N_17676);
xor U22321 (N_22321,N_18887,N_19251);
xor U22322 (N_22322,N_12846,N_13162);
xnor U22323 (N_22323,N_11209,N_14196);
xor U22324 (N_22324,N_12143,N_17536);
or U22325 (N_22325,N_19925,N_17543);
xor U22326 (N_22326,N_16575,N_18209);
or U22327 (N_22327,N_14423,N_19596);
nor U22328 (N_22328,N_18016,N_18367);
xor U22329 (N_22329,N_12508,N_18132);
and U22330 (N_22330,N_12449,N_12962);
nor U22331 (N_22331,N_12737,N_16486);
xor U22332 (N_22332,N_13131,N_15940);
nand U22333 (N_22333,N_13516,N_17838);
xnor U22334 (N_22334,N_12909,N_17645);
or U22335 (N_22335,N_16927,N_11947);
or U22336 (N_22336,N_15561,N_11812);
or U22337 (N_22337,N_15959,N_12527);
and U22338 (N_22338,N_17356,N_13988);
xor U22339 (N_22339,N_13348,N_11033);
xnor U22340 (N_22340,N_16014,N_19455);
nand U22341 (N_22341,N_14436,N_18727);
or U22342 (N_22342,N_15072,N_10082);
xnor U22343 (N_22343,N_17974,N_15629);
or U22344 (N_22344,N_17092,N_19409);
nand U22345 (N_22345,N_18423,N_19819);
and U22346 (N_22346,N_11392,N_19145);
nor U22347 (N_22347,N_19687,N_18592);
nand U22348 (N_22348,N_19420,N_15578);
or U22349 (N_22349,N_14971,N_15329);
or U22350 (N_22350,N_14408,N_17179);
or U22351 (N_22351,N_16633,N_10249);
xnor U22352 (N_22352,N_18263,N_11683);
nand U22353 (N_22353,N_15835,N_18485);
or U22354 (N_22354,N_19831,N_19007);
or U22355 (N_22355,N_16560,N_13705);
and U22356 (N_22356,N_10599,N_19711);
nand U22357 (N_22357,N_14540,N_12405);
nor U22358 (N_22358,N_11422,N_19372);
xnor U22359 (N_22359,N_19156,N_15380);
and U22360 (N_22360,N_12166,N_11414);
and U22361 (N_22361,N_16010,N_10803);
and U22362 (N_22362,N_11377,N_19246);
nor U22363 (N_22363,N_19726,N_12712);
and U22364 (N_22364,N_12340,N_19504);
xor U22365 (N_22365,N_17276,N_18500);
and U22366 (N_22366,N_17925,N_12324);
nand U22367 (N_22367,N_11702,N_10475);
nand U22368 (N_22368,N_16426,N_17151);
or U22369 (N_22369,N_13921,N_12084);
nor U22370 (N_22370,N_10556,N_11211);
and U22371 (N_22371,N_12930,N_19292);
nand U22372 (N_22372,N_17600,N_13065);
and U22373 (N_22373,N_12235,N_13346);
nor U22374 (N_22374,N_12384,N_15595);
nor U22375 (N_22375,N_10176,N_13424);
nor U22376 (N_22376,N_16610,N_10567);
and U22377 (N_22377,N_12752,N_12238);
or U22378 (N_22378,N_16912,N_11025);
xor U22379 (N_22379,N_12266,N_11294);
or U22380 (N_22380,N_14335,N_19559);
nand U22381 (N_22381,N_14974,N_10679);
nand U22382 (N_22382,N_15123,N_16075);
nor U22383 (N_22383,N_17004,N_19760);
nor U22384 (N_22384,N_10479,N_14228);
and U22385 (N_22385,N_14028,N_17829);
xnor U22386 (N_22386,N_17792,N_16789);
xor U22387 (N_22387,N_14362,N_16053);
nor U22388 (N_22388,N_10832,N_12818);
nand U22389 (N_22389,N_18524,N_16688);
nor U22390 (N_22390,N_13033,N_11525);
and U22391 (N_22391,N_16860,N_14280);
nor U22392 (N_22392,N_19783,N_15291);
xor U22393 (N_22393,N_18925,N_16110);
nor U22394 (N_22394,N_12958,N_19129);
nand U22395 (N_22395,N_11867,N_15781);
nand U22396 (N_22396,N_19232,N_10718);
or U22397 (N_22397,N_19152,N_17114);
xnor U22398 (N_22398,N_11226,N_19578);
nor U22399 (N_22399,N_16650,N_17227);
nor U22400 (N_22400,N_13628,N_15646);
or U22401 (N_22401,N_12604,N_17226);
and U22402 (N_22402,N_17156,N_14698);
nor U22403 (N_22403,N_10070,N_13830);
xnor U22404 (N_22404,N_19201,N_10878);
xnor U22405 (N_22405,N_17061,N_12002);
xor U22406 (N_22406,N_12717,N_11814);
xor U22407 (N_22407,N_17857,N_14682);
and U22408 (N_22408,N_13471,N_10432);
xor U22409 (N_22409,N_18338,N_17912);
nor U22410 (N_22410,N_19786,N_17710);
nand U22411 (N_22411,N_15298,N_12366);
and U22412 (N_22412,N_10184,N_16143);
or U22413 (N_22413,N_18010,N_19962);
and U22414 (N_22414,N_13912,N_10366);
or U22415 (N_22415,N_15732,N_14714);
and U22416 (N_22416,N_11502,N_19073);
and U22417 (N_22417,N_15462,N_15309);
nor U22418 (N_22418,N_17570,N_19916);
nand U22419 (N_22419,N_12480,N_11808);
xnor U22420 (N_22420,N_12098,N_19570);
xor U22421 (N_22421,N_14462,N_11640);
or U22422 (N_22422,N_18477,N_18966);
or U22423 (N_22423,N_10043,N_14399);
nor U22424 (N_22424,N_15768,N_10706);
or U22425 (N_22425,N_18051,N_14207);
and U22426 (N_22426,N_17496,N_10456);
nor U22427 (N_22427,N_12898,N_11681);
or U22428 (N_22428,N_17210,N_16497);
xor U22429 (N_22429,N_14044,N_18631);
nand U22430 (N_22430,N_15411,N_11323);
xnor U22431 (N_22431,N_19884,N_19117);
or U22432 (N_22432,N_12942,N_13177);
and U22433 (N_22433,N_16204,N_14983);
xnor U22434 (N_22434,N_19775,N_19091);
nand U22435 (N_22435,N_17961,N_11982);
nand U22436 (N_22436,N_16841,N_12650);
and U22437 (N_22437,N_11136,N_19301);
or U22438 (N_22438,N_13420,N_12700);
nor U22439 (N_22439,N_13700,N_16335);
xor U22440 (N_22440,N_11039,N_12781);
xor U22441 (N_22441,N_18934,N_18669);
nor U22442 (N_22442,N_14318,N_19807);
or U22443 (N_22443,N_15625,N_19789);
nand U22444 (N_22444,N_12196,N_12753);
xor U22445 (N_22445,N_16802,N_17698);
nand U22446 (N_22446,N_17410,N_13171);
or U22447 (N_22447,N_15745,N_10293);
or U22448 (N_22448,N_14302,N_15551);
or U22449 (N_22449,N_19379,N_16819);
nand U22450 (N_22450,N_18874,N_11542);
and U22451 (N_22451,N_16467,N_15558);
xnor U22452 (N_22452,N_19528,N_12918);
nor U22453 (N_22453,N_11383,N_16698);
nand U22454 (N_22454,N_12955,N_19931);
and U22455 (N_22455,N_14065,N_19441);
nand U22456 (N_22456,N_19339,N_15183);
nand U22457 (N_22457,N_14552,N_13761);
nor U22458 (N_22458,N_10759,N_16034);
and U22459 (N_22459,N_17981,N_17706);
nor U22460 (N_22460,N_17959,N_10418);
or U22461 (N_22461,N_13280,N_17326);
xor U22462 (N_22462,N_16098,N_11924);
or U22463 (N_22463,N_14104,N_16378);
nor U22464 (N_22464,N_15337,N_11474);
nand U22465 (N_22465,N_19818,N_13066);
and U22466 (N_22466,N_10153,N_18496);
nor U22467 (N_22467,N_12049,N_14815);
nor U22468 (N_22468,N_13593,N_14857);
nor U22469 (N_22469,N_13974,N_10776);
nand U22470 (N_22470,N_14386,N_19240);
or U22471 (N_22471,N_19904,N_10372);
or U22472 (N_22472,N_10287,N_17348);
nand U22473 (N_22473,N_16991,N_15373);
and U22474 (N_22474,N_19454,N_14220);
nor U22475 (N_22475,N_17919,N_19495);
nor U22476 (N_22476,N_11043,N_18625);
nand U22477 (N_22477,N_11237,N_17047);
and U22478 (N_22478,N_15385,N_12456);
xor U22479 (N_22479,N_18512,N_18443);
xnor U22480 (N_22480,N_14561,N_18765);
nand U22481 (N_22481,N_16493,N_14155);
nor U22482 (N_22482,N_15006,N_14311);
and U22483 (N_22483,N_16644,N_18994);
and U22484 (N_22484,N_19697,N_19754);
and U22485 (N_22485,N_18444,N_12471);
nand U22486 (N_22486,N_19325,N_19386);
and U22487 (N_22487,N_13936,N_18959);
and U22488 (N_22488,N_10887,N_14846);
nand U22489 (N_22489,N_16272,N_11433);
or U22490 (N_22490,N_14500,N_16461);
and U22491 (N_22491,N_19289,N_17518);
or U22492 (N_22492,N_18629,N_19430);
nand U22493 (N_22493,N_17841,N_18368);
xor U22494 (N_22494,N_12538,N_17161);
xor U22495 (N_22495,N_19739,N_13624);
nor U22496 (N_22496,N_17649,N_19885);
nand U22497 (N_22497,N_14184,N_15134);
nor U22498 (N_22498,N_15351,N_18516);
or U22499 (N_22499,N_16821,N_17648);
nor U22500 (N_22500,N_15886,N_16915);
or U22501 (N_22501,N_14338,N_17424);
and U22502 (N_22502,N_12823,N_18955);
nand U22503 (N_22503,N_18550,N_16859);
nor U22504 (N_22504,N_13107,N_17242);
nor U22505 (N_22505,N_10197,N_14778);
or U22506 (N_22506,N_15051,N_16680);
or U22507 (N_22507,N_17408,N_17539);
xnor U22508 (N_22508,N_13147,N_15088);
or U22509 (N_22509,N_19683,N_16996);
or U22510 (N_22510,N_12070,N_12400);
nor U22511 (N_22511,N_15059,N_12157);
and U22512 (N_22512,N_10621,N_13989);
xnor U22513 (N_22513,N_17843,N_18572);
nor U22514 (N_22514,N_13031,N_18726);
nor U22515 (N_22515,N_18358,N_11371);
nor U22516 (N_22516,N_15421,N_13551);
nand U22517 (N_22517,N_17383,N_10489);
nor U22518 (N_22518,N_10765,N_14991);
nor U22519 (N_22519,N_13050,N_13630);
xor U22520 (N_22520,N_13064,N_19856);
and U22521 (N_22521,N_13256,N_11781);
xor U22522 (N_22522,N_18237,N_18578);
nor U22523 (N_22523,N_12437,N_10181);
nor U22524 (N_22524,N_15381,N_10860);
or U22525 (N_22525,N_13993,N_14616);
xnor U22526 (N_22526,N_18976,N_16665);
or U22527 (N_22527,N_17412,N_15696);
nor U22528 (N_22528,N_12882,N_13560);
nand U22529 (N_22529,N_10351,N_11494);
and U22530 (N_22530,N_10673,N_15702);
and U22531 (N_22531,N_17195,N_12555);
nor U22532 (N_22532,N_12854,N_17815);
nor U22533 (N_22533,N_19502,N_18229);
nand U22534 (N_22534,N_14206,N_17846);
or U22535 (N_22535,N_13433,N_13530);
xor U22536 (N_22536,N_16228,N_17363);
nand U22537 (N_22537,N_13584,N_16449);
nor U22538 (N_22538,N_16759,N_18071);
or U22539 (N_22539,N_14115,N_17417);
nand U22540 (N_22540,N_10582,N_16947);
nor U22541 (N_22541,N_17852,N_17716);
and U22542 (N_22542,N_14986,N_15819);
and U22543 (N_22543,N_14567,N_19646);
and U22544 (N_22544,N_13836,N_10644);
nor U22545 (N_22545,N_10010,N_18003);
nor U22546 (N_22546,N_15340,N_15749);
and U22547 (N_22547,N_12265,N_17018);
nor U22548 (N_22548,N_12765,N_12105);
or U22549 (N_22549,N_18127,N_19835);
nor U22550 (N_22550,N_18232,N_13047);
nor U22551 (N_22551,N_15853,N_15221);
xnor U22552 (N_22552,N_17611,N_15278);
xnor U22553 (N_22553,N_15002,N_10379);
or U22554 (N_22554,N_14663,N_16260);
and U22555 (N_22555,N_15624,N_16028);
and U22556 (N_22556,N_12728,N_13183);
nor U22557 (N_22557,N_13897,N_19777);
and U22558 (N_22558,N_13400,N_17860);
nand U22559 (N_22559,N_19738,N_16012);
and U22560 (N_22560,N_16285,N_14282);
nor U22561 (N_22561,N_17261,N_13979);
nand U22562 (N_22562,N_11639,N_16149);
nand U22563 (N_22563,N_16042,N_19081);
and U22564 (N_22564,N_10642,N_13684);
or U22565 (N_22565,N_15747,N_12095);
nand U22566 (N_22566,N_14810,N_17964);
nand U22567 (N_22567,N_11264,N_14053);
and U22568 (N_22568,N_17521,N_14067);
nand U22569 (N_22569,N_14811,N_16348);
or U22570 (N_22570,N_18276,N_15328);
and U22571 (N_22571,N_19032,N_16185);
nand U22572 (N_22572,N_12142,N_10049);
nand U22573 (N_22573,N_15365,N_11028);
nand U22574 (N_22574,N_11833,N_15173);
or U22575 (N_22575,N_14498,N_11149);
nor U22576 (N_22576,N_11172,N_16452);
and U22577 (N_22577,N_12963,N_11228);
xor U22578 (N_22578,N_14635,N_16316);
nor U22579 (N_22579,N_18762,N_16245);
nor U22580 (N_22580,N_13706,N_16587);
or U22581 (N_22581,N_10074,N_19142);
and U22582 (N_22582,N_19589,N_12944);
nand U22583 (N_22583,N_16217,N_13991);
and U22584 (N_22584,N_15428,N_15471);
xor U22585 (N_22585,N_14026,N_16413);
nor U22586 (N_22586,N_11263,N_11199);
nor U22587 (N_22587,N_14132,N_11753);
nor U22588 (N_22588,N_11656,N_16874);
and U22589 (N_22589,N_17299,N_11412);
nand U22590 (N_22590,N_13216,N_12695);
nor U22591 (N_22591,N_14900,N_15024);
and U22592 (N_22592,N_18467,N_18450);
xor U22593 (N_22593,N_11601,N_12950);
nor U22594 (N_22594,N_17013,N_12867);
and U22595 (N_22595,N_12791,N_19410);
and U22596 (N_22596,N_10764,N_13149);
nor U22597 (N_22597,N_17380,N_13923);
xor U22598 (N_22598,N_12484,N_15485);
nor U22599 (N_22599,N_16564,N_10800);
or U22600 (N_22600,N_15651,N_19098);
xor U22601 (N_22601,N_11119,N_10521);
or U22602 (N_22602,N_13605,N_14001);
nor U22603 (N_22603,N_19298,N_12723);
xor U22604 (N_22604,N_19053,N_16123);
xnor U22605 (N_22605,N_10657,N_12485);
nand U22606 (N_22606,N_16761,N_11309);
and U22607 (N_22607,N_19617,N_18324);
nor U22608 (N_22608,N_14898,N_17393);
or U22609 (N_22609,N_18453,N_17910);
nor U22610 (N_22610,N_10326,N_11388);
nand U22611 (N_22611,N_11448,N_18197);
and U22612 (N_22612,N_16147,N_19923);
nor U22613 (N_22613,N_11857,N_12014);
and U22614 (N_22614,N_14875,N_19047);
xor U22615 (N_22615,N_17244,N_16666);
or U22616 (N_22616,N_15622,N_13659);
xnor U22617 (N_22617,N_14831,N_15887);
nand U22618 (N_22618,N_10641,N_11791);
nor U22619 (N_22619,N_11492,N_13466);
nand U22620 (N_22620,N_11789,N_13778);
or U22621 (N_22621,N_11370,N_12684);
nand U22622 (N_22622,N_17950,N_15013);
and U22623 (N_22623,N_16944,N_16749);
or U22624 (N_22624,N_12734,N_19196);
nand U22625 (N_22625,N_18469,N_16372);
or U22626 (N_22626,N_12322,N_15186);
nor U22627 (N_22627,N_11357,N_19260);
nand U22628 (N_22628,N_12144,N_14058);
and U22629 (N_22629,N_13539,N_14747);
nand U22630 (N_22630,N_16279,N_15234);
and U22631 (N_22631,N_15678,N_18086);
nor U22632 (N_22632,N_17464,N_13153);
nand U22633 (N_22633,N_18305,N_12594);
xor U22634 (N_22634,N_19366,N_19801);
xnor U22635 (N_22635,N_19799,N_15533);
and U22636 (N_22636,N_18940,N_13151);
nand U22637 (N_22637,N_13019,N_15683);
or U22638 (N_22638,N_12981,N_17726);
and U22639 (N_22639,N_16266,N_13163);
nand U22640 (N_22640,N_19509,N_11204);
xor U22641 (N_22641,N_16583,N_13524);
nand U22642 (N_22642,N_13765,N_18353);
xnor U22643 (N_22643,N_16554,N_11256);
or U22644 (N_22644,N_10979,N_13785);
or U22645 (N_22645,N_16060,N_11611);
xnor U22646 (N_22646,N_17760,N_13028);
nor U22647 (N_22647,N_14092,N_15593);
xnor U22648 (N_22648,N_11590,N_15469);
nand U22649 (N_22649,N_17403,N_13546);
nand U22650 (N_22650,N_16435,N_10689);
or U22651 (N_22651,N_12964,N_12751);
or U22652 (N_22652,N_12966,N_17480);
and U22653 (N_22653,N_15039,N_18650);
and U22654 (N_22654,N_15821,N_19165);
nand U22655 (N_22655,N_12032,N_11089);
xor U22656 (N_22656,N_16117,N_14054);
or U22657 (N_22657,N_11662,N_18194);
nand U22658 (N_22658,N_10926,N_14271);
or U22659 (N_22659,N_18275,N_14766);
nand U22660 (N_22660,N_16600,N_18495);
or U22661 (N_22661,N_17674,N_16299);
and U22662 (N_22662,N_17182,N_16408);
and U22663 (N_22663,N_15085,N_16105);
and U22664 (N_22664,N_14978,N_19227);
nand U22665 (N_22665,N_13913,N_18885);
and U22666 (N_22666,N_15785,N_12209);
and U22667 (N_22667,N_14332,N_19866);
or U22668 (N_22668,N_13738,N_16757);
nand U22669 (N_22669,N_15971,N_17922);
and U22670 (N_22670,N_17755,N_18023);
nor U22671 (N_22671,N_13622,N_15128);
nand U22672 (N_22672,N_17239,N_19978);
nand U22673 (N_22673,N_13268,N_15087);
and U22674 (N_22674,N_12288,N_11181);
nor U22675 (N_22675,N_18867,N_14577);
nor U22676 (N_22676,N_18097,N_11060);
nand U22677 (N_22677,N_13052,N_13803);
nor U22678 (N_22678,N_11756,N_16561);
nand U22679 (N_22679,N_17720,N_16399);
and U22680 (N_22680,N_14869,N_10264);
xor U22681 (N_22681,N_17668,N_10084);
and U22682 (N_22682,N_16973,N_13910);
nand U22683 (N_22683,N_18114,N_19041);
nand U22684 (N_22684,N_12617,N_16261);
or U22685 (N_22685,N_11999,N_15870);
or U22686 (N_22686,N_16384,N_16812);
and U22687 (N_22687,N_14966,N_11707);
xor U22688 (N_22688,N_17794,N_15649);
and U22689 (N_22689,N_19713,N_10445);
nor U22690 (N_22690,N_11258,N_17730);
or U22691 (N_22691,N_10932,N_11798);
xor U22692 (N_22692,N_19657,N_17133);
xor U22693 (N_22693,N_17202,N_13668);
nand U22694 (N_22694,N_13013,N_10842);
and U22695 (N_22695,N_12303,N_18387);
or U22696 (N_22696,N_19438,N_19286);
nand U22697 (N_22697,N_16403,N_14935);
nor U22698 (N_22698,N_10343,N_12948);
xnor U22699 (N_22699,N_13779,N_18764);
nor U22700 (N_22700,N_13279,N_17117);
nor U22701 (N_22701,N_15900,N_13281);
and U22702 (N_22702,N_17223,N_14606);
nor U22703 (N_22703,N_10584,N_19584);
xnor U22704 (N_22704,N_14064,N_12935);
xnor U22705 (N_22705,N_17615,N_18784);
and U22706 (N_22706,N_18646,N_12048);
and U22707 (N_22707,N_10198,N_16632);
or U22708 (N_22708,N_14867,N_10566);
or U22709 (N_22709,N_13040,N_16808);
nor U22710 (N_22710,N_17895,N_16669);
and U22711 (N_22711,N_11366,N_18989);
xor U22712 (N_22712,N_15708,N_16961);
xor U22713 (N_22713,N_10206,N_19707);
or U22714 (N_22714,N_10219,N_16179);
nand U22715 (N_22715,N_19901,N_19040);
and U22716 (N_22716,N_11862,N_10983);
xnor U22717 (N_22717,N_16616,N_10291);
and U22718 (N_22718,N_11855,N_18188);
and U22719 (N_22719,N_17254,N_12722);
or U22720 (N_22720,N_13477,N_18002);
nor U22721 (N_22721,N_19406,N_12813);
and U22722 (N_22722,N_10411,N_11369);
nand U22723 (N_22723,N_11068,N_11600);
and U22724 (N_22724,N_15046,N_11576);
and U22725 (N_22725,N_10212,N_16622);
xnor U22726 (N_22726,N_17992,N_13486);
xor U22727 (N_22727,N_10394,N_10631);
nand U22728 (N_22728,N_13967,N_15438);
or U22729 (N_22729,N_10441,N_11219);
nor U22730 (N_22730,N_12526,N_12323);
nand U22731 (N_22731,N_10304,N_17529);
nor U22732 (N_22732,N_10565,N_18525);
xnor U22733 (N_22733,N_16985,N_18173);
xor U22734 (N_22734,N_13945,N_15881);
nor U22735 (N_22735,N_18482,N_13711);
xor U22736 (N_22736,N_17850,N_16892);
nor U22737 (N_22737,N_13851,N_17644);
nor U22738 (N_22738,N_15806,N_15859);
nand U22739 (N_22739,N_12509,N_11969);
nor U22740 (N_22740,N_17229,N_16714);
or U22741 (N_22741,N_19497,N_17031);
nor U22742 (N_22742,N_12740,N_12679);
nand U22743 (N_22743,N_18304,N_10485);
nor U22744 (N_22744,N_14146,N_17205);
and U22745 (N_22745,N_10321,N_16599);
xnor U22746 (N_22746,N_19729,N_16227);
or U22747 (N_22747,N_17601,N_11483);
or U22748 (N_22748,N_18125,N_16559);
nand U22749 (N_22749,N_16109,N_16153);
xor U22750 (N_22750,N_17372,N_15127);
xor U22751 (N_22751,N_13210,N_14798);
nand U22752 (N_22752,N_14426,N_18853);
xor U22753 (N_22753,N_18591,N_15666);
nor U22754 (N_22754,N_14421,N_10476);
nand U22755 (N_22755,N_14494,N_17929);
or U22756 (N_22756,N_19336,N_12727);
nor U22757 (N_22757,N_14331,N_11467);
xor U22758 (N_22758,N_15818,N_15414);
nand U22759 (N_22759,N_16366,N_18149);
nor U22760 (N_22760,N_15480,N_11480);
and U22761 (N_22761,N_12111,N_17928);
nand U22762 (N_22762,N_11460,N_10385);
or U22763 (N_22763,N_10245,N_16494);
or U22764 (N_22764,N_13617,N_17877);
and U22765 (N_22765,N_15537,N_11478);
or U22766 (N_22766,N_19484,N_15746);
nand U22767 (N_22767,N_13600,N_14278);
nor U22768 (N_22768,N_17501,N_16247);
and U22769 (N_22769,N_11080,N_11374);
xnor U22770 (N_22770,N_19718,N_11720);
nand U22771 (N_22771,N_18376,N_15499);
or U22772 (N_22772,N_18993,N_17442);
nor U22773 (N_22773,N_12337,N_17048);
and U22774 (N_22774,N_10156,N_17236);
nor U22775 (N_22775,N_19300,N_14818);
or U22776 (N_22776,N_15958,N_13956);
xor U22777 (N_22777,N_14656,N_11888);
and U22778 (N_22778,N_14021,N_11368);
and U22779 (N_22779,N_17447,N_12125);
or U22780 (N_22780,N_18552,N_15554);
nand U22781 (N_22781,N_17853,N_12023);
nor U22782 (N_22782,N_15630,N_17738);
and U22783 (N_22783,N_15826,N_19348);
xor U22784 (N_22784,N_19544,N_16639);
nand U22785 (N_22785,N_16782,N_11449);
nor U22786 (N_22786,N_14075,N_16240);
xor U22787 (N_22787,N_16609,N_13312);
nand U22788 (N_22788,N_12000,N_17590);
xor U22789 (N_22789,N_13086,N_13138);
nand U22790 (N_22790,N_17445,N_17867);
or U22791 (N_22791,N_19979,N_19935);
xor U22792 (N_22792,N_10158,N_12687);
or U22793 (N_22793,N_17219,N_13469);
or U22794 (N_22794,N_17243,N_15014);
nand U22795 (N_22795,N_15701,N_11284);
nand U22796 (N_22796,N_15843,N_12272);
nand U22797 (N_22797,N_16048,N_14027);
xnor U22798 (N_22798,N_10943,N_14097);
and U22799 (N_22799,N_19014,N_15100);
or U22800 (N_22800,N_14969,N_10919);
and U22801 (N_22801,N_11351,N_15513);
or U22802 (N_22802,N_19029,N_11688);
and U22803 (N_22803,N_17699,N_11581);
and U22804 (N_22804,N_16114,N_19618);
or U22805 (N_22805,N_12217,N_15885);
and U22806 (N_22806,N_15342,N_10840);
nor U22807 (N_22807,N_18081,N_18308);
xnor U22808 (N_22808,N_17808,N_12494);
and U22809 (N_22809,N_10810,N_10901);
nand U22810 (N_22810,N_10273,N_15158);
xor U22811 (N_22811,N_15393,N_13723);
nand U22812 (N_22812,N_17936,N_10355);
nand U22813 (N_22813,N_17541,N_15401);
nor U22814 (N_22814,N_15626,N_13180);
and U22815 (N_22815,N_16314,N_16818);
xor U22816 (N_22816,N_11421,N_12634);
nand U22817 (N_22817,N_16419,N_17980);
and U22818 (N_22818,N_17713,N_11055);
nand U22819 (N_22819,N_10302,N_14459);
xor U22820 (N_22820,N_12814,N_15065);
or U22821 (N_22821,N_18881,N_10100);
and U22822 (N_22822,N_14029,N_19311);
or U22823 (N_22823,N_18356,N_13619);
nand U22824 (N_22824,N_15334,N_16550);
nand U22825 (N_22825,N_11900,N_16052);
xnor U22826 (N_22826,N_16972,N_18124);
or U22827 (N_22827,N_17020,N_16585);
or U22828 (N_22828,N_11669,N_11655);
nand U22829 (N_22829,N_19183,N_13265);
xnor U22830 (N_22830,N_16407,N_19150);
nand U22831 (N_22831,N_14238,N_14559);
and U22832 (N_22832,N_11192,N_16441);
or U22833 (N_22833,N_11431,N_12440);
xor U22834 (N_22834,N_16077,N_12275);
nor U22835 (N_22835,N_18219,N_16840);
or U22836 (N_22836,N_14169,N_11010);
and U22837 (N_22837,N_13058,N_10669);
xnor U22838 (N_22838,N_12321,N_10896);
nor U22839 (N_22839,N_16535,N_17019);
nand U22840 (N_22840,N_15799,N_11515);
nand U22841 (N_22841,N_10057,N_14293);
xnor U22842 (N_22842,N_12291,N_12257);
nor U22843 (N_22843,N_17693,N_14279);
xnor U22844 (N_22844,N_11550,N_19006);
xor U22845 (N_22845,N_19478,N_12645);
and U22846 (N_22846,N_19337,N_13124);
nor U22847 (N_22847,N_17406,N_14106);
or U22848 (N_22848,N_15726,N_14602);
and U22849 (N_22849,N_14942,N_13685);
and U22850 (N_22850,N_11424,N_16165);
nor U22851 (N_22851,N_16099,N_11517);
or U22852 (N_22852,N_14474,N_14088);
or U22853 (N_22853,N_18331,N_10741);
nand U22854 (N_22854,N_14125,N_18876);
xnor U22855 (N_22855,N_15199,N_15986);
xor U22856 (N_22856,N_15691,N_17160);
nand U22857 (N_22857,N_18091,N_15333);
nand U22858 (N_22858,N_17571,N_10109);
and U22859 (N_22859,N_17487,N_19000);
xor U22860 (N_22860,N_16135,N_14471);
or U22861 (N_22861,N_16762,N_11308);
nand U22862 (N_22862,N_18978,N_18747);
or U22863 (N_22863,N_14085,N_16615);
and U22864 (N_22864,N_14512,N_16888);
nor U22865 (N_22865,N_17257,N_18850);
and U22866 (N_22866,N_14947,N_15230);
or U22867 (N_22867,N_14389,N_10865);
nand U22868 (N_22868,N_18995,N_19249);
nand U22869 (N_22869,N_18527,N_18207);
nor U22870 (N_22870,N_13875,N_19131);
or U22871 (N_22871,N_19070,N_18395);
and U22872 (N_22872,N_14677,N_19451);
nor U22873 (N_22873,N_10161,N_13294);
and U22874 (N_22874,N_11705,N_14310);
and U22875 (N_22875,N_13014,N_17088);
xor U22876 (N_22876,N_10044,N_10128);
xnor U22877 (N_22877,N_12947,N_13166);
xnor U22878 (N_22878,N_14630,N_17328);
or U22879 (N_22879,N_11513,N_10500);
nor U22880 (N_22880,N_19852,N_16528);
xnor U22881 (N_22881,N_18268,N_10980);
or U22882 (N_22882,N_17897,N_16683);
nand U22883 (N_22883,N_19887,N_12730);
and U22884 (N_22884,N_13500,N_11755);
and U22885 (N_22885,N_11723,N_15994);
nor U22886 (N_22886,N_14990,N_12190);
or U22887 (N_22887,N_12409,N_15611);
xnor U22888 (N_22888,N_12937,N_17696);
and U22889 (N_22889,N_12215,N_18508);
or U22890 (N_22890,N_15776,N_17666);
and U22891 (N_22891,N_11230,N_17391);
nand U22892 (N_22892,N_10004,N_10102);
nor U22893 (N_22893,N_18094,N_13472);
or U22894 (N_22894,N_19306,N_10913);
nor U22895 (N_22895,N_10022,N_18317);
or U22896 (N_22896,N_14095,N_15363);
or U22897 (N_22897,N_11524,N_14202);
xnor U22898 (N_22898,N_10461,N_16485);
or U22899 (N_22899,N_10617,N_10031);
or U22900 (N_22900,N_17463,N_14745);
nor U22901 (N_22901,N_19106,N_15222);
or U22902 (N_22902,N_14716,N_14641);
or U22903 (N_22903,N_17831,N_12755);
nand U22904 (N_22904,N_13675,N_15103);
or U22905 (N_22905,N_13143,N_17927);
nor U22906 (N_22906,N_12100,N_17467);
nand U22907 (N_22907,N_15931,N_16842);
nand U22908 (N_22908,N_17218,N_16629);
nor U22909 (N_22909,N_12655,N_18101);
or U22910 (N_22910,N_14835,N_13751);
or U22911 (N_22911,N_13368,N_14131);
nand U22912 (N_22912,N_14727,N_12292);
nand U22913 (N_22913,N_16061,N_18688);
and U22914 (N_22914,N_11741,N_14599);
nor U22915 (N_22915,N_15526,N_12022);
nor U22916 (N_22916,N_13271,N_19498);
and U22917 (N_22917,N_14208,N_10413);
and U22918 (N_22918,N_13226,N_17572);
xnor U22919 (N_22919,N_16970,N_18677);
and U22920 (N_22920,N_16520,N_18325);
and U22921 (N_22921,N_15194,N_19359);
xor U22922 (N_22922,N_16257,N_15620);
and U22923 (N_22923,N_13841,N_12614);
nand U22924 (N_22924,N_14341,N_12153);
or U22925 (N_22925,N_19857,N_14680);
and U22926 (N_22926,N_17336,N_15276);
nor U22927 (N_22927,N_14506,N_11796);
and U22928 (N_22928,N_17610,N_12894);
xnor U22929 (N_22929,N_15143,N_12237);
nor U22930 (N_22930,N_10065,N_15454);
nor U22931 (N_22931,N_15798,N_13906);
or U22932 (N_22932,N_19025,N_13868);
nor U22933 (N_22933,N_19119,N_18117);
and U22934 (N_22934,N_17159,N_14886);
nand U22935 (N_22935,N_10447,N_10920);
xor U22936 (N_22936,N_19611,N_11991);
xor U22937 (N_22937,N_14833,N_18186);
and U22938 (N_22938,N_11599,N_11633);
xor U22939 (N_22939,N_19984,N_19825);
and U22940 (N_22940,N_16256,N_13450);
xor U22941 (N_22941,N_19500,N_13998);
xnor U22942 (N_22942,N_18542,N_11844);
xnor U22943 (N_22943,N_18293,N_16863);
nor U22944 (N_22944,N_12640,N_13232);
and U22945 (N_22945,N_10173,N_16527);
and U22946 (N_22946,N_10884,N_11141);
xor U22947 (N_22947,N_11210,N_14047);
nand U22948 (N_22948,N_18017,N_13952);
nor U22949 (N_22949,N_18300,N_13722);
or U22950 (N_22950,N_18564,N_19563);
or U22951 (N_22951,N_19418,N_10037);
or U22952 (N_22952,N_11938,N_19124);
nor U22953 (N_22953,N_13326,N_10174);
nor U22954 (N_22954,N_15851,N_18024);
nor U22955 (N_22955,N_16004,N_14069);
nand U22956 (N_22956,N_14403,N_14657);
and U22957 (N_22957,N_16087,N_19907);
and U22958 (N_22958,N_18474,N_12805);
xor U22959 (N_22959,N_16895,N_11925);
and U22960 (N_22960,N_10723,N_16674);
and U22961 (N_22961,N_11277,N_16620);
or U22962 (N_22962,N_17522,N_11008);
nor U22963 (N_22963,N_18797,N_15970);
or U22964 (N_22964,N_17454,N_17508);
nor U22965 (N_22965,N_19577,N_19370);
nand U22966 (N_22966,N_18905,N_18470);
nor U22967 (N_22967,N_16613,N_12091);
nor U22968 (N_22968,N_12790,N_10950);
or U22969 (N_22969,N_16304,N_10618);
nor U22970 (N_22970,N_16262,N_17164);
and U22971 (N_22971,N_15935,N_13393);
nor U22972 (N_22972,N_14691,N_11356);
xor U22973 (N_22973,N_13784,N_19198);
or U22974 (N_22974,N_14830,N_18320);
nand U22975 (N_22975,N_12908,N_14175);
nand U22976 (N_22976,N_10464,N_13377);
nor U22977 (N_22977,N_19054,N_17599);
nand U22978 (N_22978,N_14534,N_13657);
and U22979 (N_22979,N_13871,N_13322);
and U22980 (N_22980,N_12354,N_10576);
and U22981 (N_22981,N_13376,N_12330);
nor U22982 (N_22982,N_10252,N_16465);
xor U22983 (N_22983,N_16984,N_17622);
xnor U22984 (N_22984,N_11344,N_19433);
or U22985 (N_22985,N_19051,N_10195);
or U22986 (N_22986,N_15660,N_15614);
or U22987 (N_22987,N_19290,N_10748);
and U22988 (N_22988,N_18967,N_15357);
nor U22989 (N_22989,N_13354,N_10088);
or U22990 (N_22990,N_17613,N_15758);
nor U22991 (N_22991,N_15542,N_12550);
nor U22992 (N_22992,N_19457,N_15517);
and U22993 (N_22993,N_15543,N_16758);
or U22994 (N_22994,N_19645,N_11197);
and U22995 (N_22995,N_13026,N_15784);
and U22996 (N_22996,N_14052,N_12714);
xor U22997 (N_22997,N_13435,N_10462);
nor U22998 (N_22998,N_11567,N_19892);
and U22999 (N_22999,N_17594,N_11847);
xor U23000 (N_23000,N_15705,N_14650);
xnor U23001 (N_23001,N_18997,N_14259);
and U23002 (N_23002,N_13069,N_12152);
or U23003 (N_23003,N_16097,N_15491);
and U23004 (N_23004,N_13965,N_10241);
xnor U23005 (N_23005,N_17365,N_18544);
nor U23006 (N_23006,N_10481,N_12401);
or U23007 (N_23007,N_15762,N_18626);
or U23008 (N_23008,N_18399,N_14982);
and U23009 (N_23009,N_12939,N_17067);
nand U23010 (N_23010,N_15477,N_19650);
xor U23011 (N_23011,N_18603,N_15604);
and U23012 (N_23012,N_11477,N_18852);
or U23013 (N_23013,N_16037,N_15079);
nor U23014 (N_23014,N_12421,N_16844);
xor U23015 (N_23015,N_10894,N_13918);
nor U23016 (N_23016,N_15967,N_11744);
and U23017 (N_23017,N_11666,N_13254);
nand U23018 (N_23018,N_17728,N_10353);
and U23019 (N_23019,N_13793,N_19763);
and U23020 (N_23020,N_12487,N_17624);
xnor U23021 (N_23021,N_14676,N_16675);
and U23022 (N_23022,N_16129,N_13565);
or U23023 (N_23023,N_19477,N_18614);
and U23024 (N_23024,N_13306,N_17952);
nor U23025 (N_23025,N_12219,N_19085);
nand U23026 (N_23026,N_11177,N_11359);
nor U23027 (N_23027,N_12610,N_14858);
and U23028 (N_23028,N_16394,N_18823);
nor U23029 (N_23029,N_15050,N_17531);
nor U23030 (N_23030,N_18286,N_15019);
or U23031 (N_23031,N_11495,N_12490);
nand U23032 (N_23032,N_18963,N_18326);
nor U23033 (N_23033,N_16168,N_13316);
and U23034 (N_23034,N_19695,N_16516);
or U23035 (N_23035,N_15177,N_10510);
nor U23036 (N_23036,N_14078,N_11868);
nand U23037 (N_23037,N_12567,N_14491);
nor U23038 (N_23038,N_15053,N_15787);
xor U23039 (N_23039,N_17385,N_12500);
nor U23040 (N_23040,N_13776,N_10571);
or U23041 (N_23041,N_13453,N_10693);
xnor U23042 (N_23042,N_12829,N_19492);
nor U23043 (N_23043,N_10186,N_17749);
and U23044 (N_23044,N_15147,N_13062);
xor U23045 (N_23045,N_12254,N_15968);
or U23046 (N_23046,N_11591,N_14323);
and U23047 (N_23047,N_16120,N_12877);
or U23048 (N_23048,N_19963,N_13514);
nand U23049 (N_23049,N_19968,N_17673);
nor U23050 (N_23050,N_14866,N_16432);
xnor U23051 (N_23051,N_17420,N_11057);
nand U23052 (N_23052,N_17499,N_15093);
or U23053 (N_23053,N_16523,N_17384);
nand U23054 (N_23054,N_17025,N_13004);
nor U23055 (N_23055,N_14138,N_15520);
or U23056 (N_23056,N_17935,N_16007);
nor U23057 (N_23057,N_19548,N_16090);
and U23058 (N_23058,N_16430,N_18348);
xnor U23059 (N_23059,N_10502,N_16727);
or U23060 (N_23060,N_11234,N_11432);
or U23061 (N_23061,N_19594,N_11757);
xnor U23062 (N_23062,N_16444,N_13840);
nor U23063 (N_23063,N_14655,N_17664);
and U23064 (N_23064,N_19116,N_16820);
and U23065 (N_23065,N_10738,N_17446);
and U23066 (N_23066,N_19510,N_16167);
nand U23067 (N_23067,N_16594,N_16206);
or U23068 (N_23068,N_17515,N_11216);
nand U23069 (N_23069,N_17634,N_12735);
or U23070 (N_23070,N_18083,N_11783);
nand U23071 (N_23071,N_19934,N_16038);
and U23072 (N_23072,N_11638,N_15577);
and U23073 (N_23073,N_12411,N_17390);
xor U23074 (N_23074,N_14569,N_11123);
nor U23075 (N_23075,N_13650,N_11977);
nand U23076 (N_23076,N_16369,N_18233);
nand U23077 (N_23077,N_12136,N_16459);
nor U23078 (N_23078,N_10123,N_13362);
or U23079 (N_23079,N_18283,N_11128);
nand U23080 (N_23080,N_18039,N_12976);
and U23081 (N_23081,N_17848,N_18581);
xor U23082 (N_23082,N_16162,N_16349);
nor U23083 (N_23083,N_16563,N_11807);
or U23084 (N_23084,N_16978,N_11577);
nor U23085 (N_23085,N_11035,N_11316);
nor U23086 (N_23086,N_11598,N_18724);
nor U23087 (N_23087,N_17475,N_13488);
xnor U23088 (N_23088,N_14826,N_17550);
nor U23089 (N_23089,N_13414,N_15589);
xor U23090 (N_23090,N_10171,N_16301);
xnor U23091 (N_23091,N_18235,N_19766);
or U23092 (N_23092,N_19043,N_15056);
nor U23093 (N_23093,N_14548,N_19791);
nand U23094 (N_23094,N_13344,N_18708);
xor U23095 (N_23095,N_18878,N_17158);
and U23096 (N_23096,N_13011,N_13567);
xnor U23097 (N_23097,N_15509,N_15483);
xor U23098 (N_23098,N_16790,N_10588);
xnor U23099 (N_23099,N_13388,N_13934);
nor U23100 (N_23100,N_16783,N_12442);
or U23101 (N_23101,N_16770,N_16297);
nand U23102 (N_23102,N_13773,N_19933);
and U23103 (N_23103,N_10632,N_14096);
or U23104 (N_23104,N_13251,N_18981);
nand U23105 (N_23105,N_15163,N_19602);
or U23106 (N_23106,N_18122,N_19293);
xnor U23107 (N_23107,N_13029,N_17017);
xor U23108 (N_23108,N_11665,N_19991);
and U23109 (N_23109,N_19127,N_15432);
nor U23110 (N_23110,N_19067,N_11200);
and U23111 (N_23111,N_16323,N_15709);
and U23112 (N_23112,N_17582,N_11259);
and U23113 (N_23113,N_17335,N_16940);
nand U23114 (N_23114,N_14712,N_11295);
xnor U23115 (N_23115,N_11641,N_13861);
nor U23116 (N_23116,N_10988,N_13385);
nor U23117 (N_23117,N_19632,N_13327);
nand U23118 (N_23118,N_16230,N_16250);
nor U23119 (N_23119,N_18087,N_11881);
xnor U23120 (N_23120,N_19730,N_10284);
nand U23121 (N_23121,N_11052,N_14516);
nand U23122 (N_23122,N_13278,N_11831);
nor U23123 (N_23123,N_18728,N_14794);
nand U23124 (N_23124,N_17322,N_14668);
nor U23125 (N_23125,N_11103,N_15966);
and U23126 (N_23126,N_10371,N_10370);
nor U23127 (N_23127,N_12986,N_11092);
xnor U23128 (N_23128,N_11983,N_11489);
or U23129 (N_23129,N_11605,N_10564);
nand U23130 (N_23130,N_19167,N_18615);
nand U23131 (N_23131,N_14186,N_10964);
or U23132 (N_23132,N_13231,N_19243);
nor U23133 (N_23133,N_15114,N_19268);
or U23134 (N_23134,N_12168,N_18260);
nor U23135 (N_23135,N_18561,N_17444);
and U23136 (N_23136,N_10460,N_16303);
or U23137 (N_23137,N_14824,N_19658);
nor U23138 (N_23138,N_13767,N_10382);
and U23139 (N_23139,N_13148,N_10108);
and U23140 (N_23140,N_11643,N_18624);
xor U23141 (N_23141,N_12199,N_17637);
or U23142 (N_23142,N_15602,N_18171);
xor U23143 (N_23143,N_12424,N_11535);
nand U23144 (N_23144,N_19258,N_14932);
and U23145 (N_23145,N_17584,N_12197);
nor U23146 (N_23146,N_18882,N_18435);
or U23147 (N_23147,N_10157,N_10167);
nand U23148 (N_23148,N_19517,N_15296);
or U23149 (N_23149,N_17311,N_13027);
and U23150 (N_23150,N_19077,N_19343);
nor U23151 (N_23151,N_17191,N_18025);
and U23152 (N_23152,N_12816,N_11022);
or U23153 (N_23153,N_11416,N_13981);
or U23154 (N_23154,N_13205,N_13911);
or U23155 (N_23155,N_19561,N_17631);
nor U23156 (N_23156,N_18063,N_10041);
and U23157 (N_23157,N_19654,N_13241);
and U23158 (N_23158,N_12530,N_19328);
xor U23159 (N_23159,N_14979,N_14945);
nand U23160 (N_23160,N_16296,N_15945);
nor U23161 (N_23161,N_18806,N_11706);
xnor U23162 (N_23162,N_18273,N_18869);
or U23163 (N_23163,N_16682,N_17772);
xnor U23164 (N_23164,N_15809,N_13172);
nor U23165 (N_23165,N_17612,N_14660);
and U23166 (N_23166,N_17687,N_18649);
xnor U23167 (N_23167,N_10253,N_16103);
or U23168 (N_23168,N_10941,N_15155);
and U23169 (N_23169,N_15254,N_19958);
xor U23170 (N_23170,N_18381,N_14055);
nor U23171 (N_23171,N_13165,N_11381);
or U23172 (N_23172,N_16925,N_15389);
nand U23173 (N_23173,N_13859,N_12954);
or U23174 (N_23174,N_15362,N_18555);
and U23175 (N_23175,N_10388,N_12436);
and U23176 (N_23176,N_17039,N_15616);
nor U23177 (N_23177,N_12058,N_15466);
xor U23178 (N_23178,N_13820,N_13370);
nor U23179 (N_23179,N_17845,N_11561);
xnor U23180 (N_23180,N_10912,N_13487);
xnor U23181 (N_23181,N_11788,N_14156);
nand U23182 (N_23182,N_17732,N_10250);
and U23183 (N_23183,N_11903,N_17894);
and U23184 (N_23184,N_15175,N_14225);
xnor U23185 (N_23185,N_17805,N_18156);
nor U23186 (N_23186,N_19614,N_18223);
nor U23187 (N_23187,N_12686,N_11654);
or U23188 (N_23188,N_17898,N_14372);
or U23189 (N_23189,N_15946,N_17764);
nand U23190 (N_23190,N_14688,N_17280);
and U23191 (N_23191,N_11382,N_15257);
or U23192 (N_23192,N_11861,N_14855);
nor U23193 (N_23193,N_16031,N_12503);
or U23194 (N_23194,N_15527,N_11161);
xor U23195 (N_23195,N_15555,N_18390);
nand U23196 (N_23196,N_16224,N_17184);
xnor U23197 (N_23197,N_10380,N_13491);
or U23198 (N_23198,N_14992,N_12857);
or U23199 (N_23199,N_13390,N_17913);
nor U23200 (N_23200,N_16336,N_11839);
nand U23201 (N_23201,N_15803,N_10622);
nand U23202 (N_23202,N_19326,N_12667);
and U23203 (N_23203,N_12416,N_12588);
nand U23204 (N_23204,N_14759,N_16189);
and U23205 (N_23205,N_10674,N_11682);
or U23206 (N_23206,N_17900,N_15318);
nor U23207 (N_23207,N_11752,N_19952);
xor U23208 (N_23208,N_10301,N_17008);
nor U23209 (N_23209,N_11016,N_13345);
nand U23210 (N_23210,N_14406,N_13444);
nand U23211 (N_23211,N_19367,N_14248);
nand U23212 (N_23212,N_19415,N_17419);
nor U23213 (N_23213,N_17663,N_11280);
and U23214 (N_23214,N_17688,N_10867);
and U23215 (N_23215,N_10178,N_19262);
xnor U23216 (N_23216,N_17152,N_10137);
or U23217 (N_23217,N_12260,N_19149);
nand U23218 (N_23218,N_18502,N_17592);
and U23219 (N_23219,N_12230,N_11674);
and U23220 (N_23220,N_11946,N_12940);
and U23221 (N_23221,N_17690,N_17778);
or U23222 (N_23222,N_19736,N_13980);
or U23223 (N_23223,N_17937,N_13159);
nor U23224 (N_23224,N_11962,N_12065);
and U23225 (N_23225,N_16809,N_19740);
or U23226 (N_23226,N_19342,N_12353);
or U23227 (N_23227,N_10882,N_11098);
nand U23228 (N_23228,N_18901,N_10655);
nor U23229 (N_23229,N_13482,N_19130);
nor U23230 (N_23230,N_11427,N_19024);
and U23231 (N_23231,N_15216,N_19362);
nor U23232 (N_23232,N_13387,N_16375);
nand U23233 (N_23233,N_10549,N_12855);
and U23234 (N_23234,N_10671,N_19724);
nand U23235 (N_23235,N_14382,N_15482);
nor U23236 (N_23236,N_19066,N_11441);
xor U23237 (N_23237,N_13889,N_16791);
or U23238 (N_23238,N_11213,N_14273);
nand U23239 (N_23239,N_18511,N_15529);
nor U23240 (N_23240,N_18914,N_17490);
nand U23241 (N_23241,N_15138,N_18557);
nand U23242 (N_23242,N_15210,N_12488);
nor U23243 (N_23243,N_12630,N_19363);
and U23244 (N_23244,N_19988,N_11929);
xnor U23245 (N_23245,N_18176,N_15668);
or U23246 (N_23246,N_11508,N_18436);
or U23247 (N_23247,N_10925,N_15446);
and U23248 (N_23248,N_18349,N_11528);
xor U23249 (N_23249,N_17312,N_10755);
and U23250 (N_23250,N_13970,N_17186);
nand U23251 (N_23251,N_11247,N_11809);
nor U23252 (N_23252,N_17246,N_19606);
and U23253 (N_23253,N_18928,N_13669);
nor U23254 (N_23254,N_10746,N_11093);
and U23255 (N_23255,N_12373,N_13876);
and U23256 (N_23256,N_14002,N_14400);
and U23257 (N_23257,N_19282,N_19395);
nand U23258 (N_23258,N_18043,N_19644);
xor U23259 (N_23259,N_14751,N_13613);
or U23260 (N_23260,N_16717,N_17934);
nand U23261 (N_23261,N_13012,N_10712);
and U23262 (N_23262,N_13059,N_19928);
and U23263 (N_23263,N_19967,N_14446);
nor U23264 (N_23264,N_14264,N_18224);
or U23265 (N_23265,N_13860,N_16340);
nand U23266 (N_23266,N_16023,N_11794);
nand U23267 (N_23267,N_14772,N_19753);
nand U23268 (N_23268,N_15441,N_16181);
nand U23269 (N_23269,N_19678,N_15000);
or U23270 (N_23270,N_11195,N_13674);
or U23271 (N_23271,N_15854,N_19534);
xnor U23272 (N_23272,N_10151,N_12889);
or U23273 (N_23273,N_19776,N_12466);
and U23274 (N_23274,N_14686,N_11799);
and U23275 (N_23275,N_15185,N_13927);
xor U23276 (N_23276,N_15348,N_10790);
and U23277 (N_23277,N_10853,N_13843);
nor U23278 (N_23278,N_16355,N_10209);
nand U23279 (N_23279,N_12011,N_15728);
xnor U23280 (N_23280,N_15166,N_14374);
and U23281 (N_23281,N_13352,N_18745);
and U23282 (N_23282,N_15765,N_17241);
xnor U23283 (N_23283,N_10139,N_17966);
xor U23284 (N_23284,N_18980,N_14072);
or U23285 (N_23285,N_13518,N_13642);
or U23286 (N_23286,N_16118,N_18343);
and U23287 (N_23287,N_13885,N_16473);
nor U23288 (N_23288,N_16660,N_17640);
or U23289 (N_23289,N_16066,N_13823);
nand U23290 (N_23290,N_11779,N_16945);
or U23291 (N_23291,N_13242,N_18466);
and U23292 (N_23292,N_17654,N_17819);
nand U23293 (N_23293,N_17256,N_18473);
xnor U23294 (N_23294,N_19456,N_13483);
xor U23295 (N_23295,N_14025,N_12703);
nand U23296 (N_23296,N_14258,N_12392);
xor U23297 (N_23297,N_11038,N_11297);
xor U23298 (N_23298,N_13558,N_16932);
xnor U23299 (N_23299,N_13217,N_13797);
or U23300 (N_23300,N_14550,N_13167);
nor U23301 (N_23301,N_16328,N_18827);
or U23302 (N_23302,N_12035,N_18526);
nand U23303 (N_23303,N_10530,N_12788);
nand U23304 (N_23304,N_16347,N_12319);
nor U23305 (N_23305,N_10183,N_11367);
or U23306 (N_23306,N_14490,N_12211);
xnor U23307 (N_23307,N_10744,N_18047);
nor U23308 (N_23308,N_15846,N_18798);
or U23309 (N_23309,N_15906,N_17530);
xor U23310 (N_23310,N_11503,N_19870);
or U23311 (N_23311,N_12010,N_16885);
nand U23312 (N_23312,N_16152,N_17933);
and U23313 (N_23313,N_12792,N_11274);
or U23314 (N_23314,N_14726,N_16294);
and U23315 (N_23315,N_13510,N_19592);
nand U23316 (N_23316,N_13564,N_10347);
and U23317 (N_23317,N_16365,N_12884);
nand U23318 (N_23318,N_17862,N_16126);
nor U23319 (N_23319,N_15847,N_13139);
xnor U23320 (N_23320,N_10234,N_15922);
nand U23321 (N_23321,N_17989,N_16815);
nand U23322 (N_23322,N_19673,N_15154);
nand U23323 (N_23323,N_14402,N_16288);
xnor U23324 (N_23324,N_17773,N_12900);
or U23325 (N_23325,N_15573,N_13621);
nor U23326 (N_23326,N_17148,N_13492);
xnor U23327 (N_23327,N_15849,N_11614);
nor U23328 (N_23328,N_10973,N_16364);
xnor U23329 (N_23329,N_14708,N_10904);
or U23330 (N_23330,N_14998,N_10922);
and U23331 (N_23331,N_11606,N_13635);
and U23332 (N_23332,N_14807,N_15102);
and U23333 (N_23333,N_19627,N_15635);
nand U23334 (N_23334,N_19797,N_10297);
nand U23335 (N_23335,N_14862,N_18363);
or U23336 (N_23336,N_17809,N_16567);
xnor U23337 (N_23337,N_14957,N_17523);
nand U23338 (N_23338,N_16709,N_15574);
xnor U23339 (N_23339,N_19542,N_10804);
nand U23340 (N_23340,N_11527,N_17549);
xnor U23341 (N_23341,N_12268,N_11004);
xnor U23342 (N_23342,N_18157,N_16089);
or U23343 (N_23343,N_15219,N_15914);
xnor U23344 (N_23344,N_16810,N_10605);
and U23345 (N_23345,N_15047,N_12082);
or U23346 (N_23346,N_19284,N_16823);
xor U23347 (N_23347,N_11671,N_14049);
and U23348 (N_23348,N_11852,N_10766);
nand U23349 (N_23349,N_18490,N_11411);
nor U23350 (N_23350,N_18590,N_14003);
nor U23351 (N_23351,N_17360,N_19078);
or U23352 (N_23352,N_16950,N_15246);
or U23353 (N_23353,N_15457,N_14542);
nand U23354 (N_23354,N_10539,N_11182);
or U23355 (N_23355,N_12042,N_12163);
nand U23356 (N_23356,N_10278,N_18200);
or U23357 (N_23357,N_16986,N_12329);
and U23358 (N_23358,N_15055,N_14897);
or U23359 (N_23359,N_15763,N_12880);
nor U23360 (N_23360,N_10071,N_18152);
xor U23361 (N_23361,N_15061,N_11373);
or U23362 (N_23362,N_10513,N_11186);
xnor U23363 (N_23363,N_15808,N_11651);
and U23364 (N_23364,N_17740,N_10028);
nor U23365 (N_23365,N_11843,N_14847);
xor U23366 (N_23366,N_18095,N_13504);
and U23367 (N_23367,N_15407,N_12394);
xor U23368 (N_23368,N_16573,N_12422);
nand U23369 (N_23369,N_10704,N_13652);
or U23370 (N_23370,N_15544,N_17214);
nand U23371 (N_23371,N_16938,N_10403);
or U23372 (N_23372,N_10743,N_17780);
nor U23373 (N_23373,N_17286,N_18706);
nand U23374 (N_23374,N_15125,N_15897);
xnor U23375 (N_23375,N_18594,N_15105);
and U23376 (N_23376,N_16352,N_14123);
and U23377 (N_23377,N_15717,N_16597);
nor U23378 (N_23378,N_18586,N_14528);
nor U23379 (N_23379,N_17497,N_14779);
xor U23380 (N_23380,N_11021,N_14157);
xnor U23381 (N_23381,N_19095,N_16255);
and U23382 (N_23382,N_12525,N_12670);
nor U23383 (N_23383,N_14518,N_19816);
and U23384 (N_23384,N_15985,N_14287);
nor U23385 (N_23385,N_13202,N_15390);
xnor U23386 (N_23386,N_19340,N_12665);
or U23387 (N_23387,N_17005,N_12226);
nand U23388 (N_23388,N_11428,N_14454);
or U23389 (N_23389,N_16307,N_17489);
nor U23390 (N_23390,N_14369,N_16557);
xor U23391 (N_23391,N_19712,N_18290);
nand U23392 (N_23392,N_13404,N_19875);
xnor U23393 (N_23393,N_15297,N_17863);
nand U23394 (N_23394,N_15917,N_16374);
nor U23395 (N_23395,N_15655,N_12160);
nand U23396 (N_23396,N_12917,N_10434);
nor U23397 (N_23397,N_12348,N_11718);
and U23398 (N_23398,N_16686,N_11923);
xor U23399 (N_23399,N_11825,N_12128);
and U23400 (N_23400,N_14232,N_19274);
and U23401 (N_23401,N_12056,N_17240);
and U23402 (N_23402,N_16396,N_14977);
nand U23403 (N_23403,N_12807,N_16845);
xor U23404 (N_23404,N_14000,N_19638);
or U23405 (N_23405,N_10446,N_11147);
xor U23406 (N_23406,N_18858,N_14800);
or U23407 (N_23407,N_15633,N_12875);
xor U23408 (N_23408,N_16931,N_13253);
xnor U23409 (N_23409,N_13950,N_11828);
nand U23410 (N_23410,N_14181,N_11763);
or U23411 (N_23411,N_19111,N_13334);
xnor U23412 (N_23412,N_17949,N_17535);
and U23413 (N_23413,N_17330,N_11129);
xor U23414 (N_23414,N_12072,N_12044);
nor U23415 (N_23415,N_14167,N_15919);
xnor U23416 (N_23416,N_16273,N_10091);
or U23417 (N_23417,N_19174,N_12139);
nand U23418 (N_23418,N_11053,N_12271);
and U23419 (N_23419,N_15139,N_15112);
nor U23420 (N_23420,N_14022,N_11360);
xor U23421 (N_23421,N_18846,N_10318);
and U23422 (N_23422,N_13578,N_15588);
or U23423 (N_23423,N_19615,N_15956);
or U23424 (N_23424,N_15977,N_19475);
or U23425 (N_23425,N_11884,N_10962);
or U23426 (N_23426,N_15295,N_13484);
and U23427 (N_23427,N_14669,N_16854);
xor U23428 (N_23428,N_15965,N_12187);
xor U23429 (N_23429,N_17441,N_10601);
xnor U23430 (N_23430,N_16988,N_19625);
nor U23431 (N_23431,N_15500,N_15332);
xor U23432 (N_23432,N_14709,N_13707);
nand U23433 (N_23433,N_13407,N_10271);
or U23434 (N_23434,N_16538,N_16483);
nand U23435 (N_23435,N_19234,N_19038);
nand U23436 (N_23436,N_16588,N_12298);
nand U23437 (N_23437,N_16664,N_18675);
and U23438 (N_23438,N_19595,N_15384);
and U23439 (N_23439,N_10412,N_11596);
nand U23440 (N_23440,N_19496,N_16213);
and U23441 (N_23441,N_17757,N_10782);
nor U23442 (N_23442,N_11418,N_11719);
or U23443 (N_23443,N_17769,N_19132);
xnor U23444 (N_23444,N_18162,N_19313);
xnor U23445 (N_23445,N_18884,N_10214);
xnor U23446 (N_23446,N_12637,N_17485);
nor U23447 (N_23447,N_14334,N_14117);
nand U23448 (N_23448,N_12085,N_17545);
and U23449 (N_23449,N_14071,N_14661);
or U23450 (N_23450,N_16190,N_19863);
nor U23451 (N_23451,N_11864,N_19467);
nand U23452 (N_23452,N_13141,N_16967);
nand U23453 (N_23453,N_15034,N_10280);
or U23454 (N_23454,N_11445,N_19702);
xor U23455 (N_23455,N_16976,N_19294);
xnor U23456 (N_23456,N_13520,N_12502);
nand U23457 (N_23457,N_16183,N_12998);
nor U23458 (N_23458,N_16398,N_12671);
nand U23459 (N_23459,N_17121,N_18267);
xnor U23460 (N_23460,N_11465,N_19805);
xor U23461 (N_23461,N_15003,N_10300);
or U23462 (N_23462,N_13808,N_19031);
nand U23463 (N_23463,N_16290,N_17098);
or U23464 (N_23464,N_12582,N_17932);
and U23465 (N_23465,N_15434,N_18402);
nor U23466 (N_23466,N_14076,N_14183);
or U23467 (N_23467,N_13739,N_14643);
xor U23468 (N_23468,N_13191,N_11610);
and U23469 (N_23469,N_19527,N_16201);
or U23470 (N_23470,N_11214,N_17082);
or U23471 (N_23471,N_10122,N_13602);
nor U23472 (N_23472,N_12589,N_16838);
xnor U23473 (N_23473,N_12302,N_11081);
nor U23474 (N_23474,N_11901,N_16315);
and U23475 (N_23475,N_11456,N_17618);
nor U23476 (N_23476,N_15658,N_10414);
xor U23477 (N_23477,N_19487,N_14062);
nand U23478 (N_23478,N_13599,N_19162);
and U23479 (N_23479,N_19873,N_19105);
or U23480 (N_23480,N_18459,N_18393);
and U23481 (N_23481,N_12959,N_12081);
or U23482 (N_23482,N_17053,N_12479);
and U23483 (N_23483,N_17000,N_14358);
and U23484 (N_23484,N_10096,N_13185);
or U23485 (N_23485,N_16001,N_18567);
nand U23486 (N_23486,N_18819,N_11566);
nand U23487 (N_23487,N_15470,N_13339);
or U23488 (N_23488,N_10540,N_15040);
xnor U23489 (N_23489,N_12278,N_19208);
xor U23490 (N_23490,N_16137,N_19383);
or U23491 (N_23491,N_15157,N_10130);
nor U23492 (N_23492,N_13452,N_19822);
and U23493 (N_23493,N_15400,N_18596);
and U23494 (N_23494,N_13964,N_19155);
or U23495 (N_23495,N_18020,N_12913);
nand U23496 (N_23496,N_15368,N_13366);
xnor U23497 (N_23497,N_15564,N_13930);
nor U23498 (N_23498,N_19485,N_12773);
or U23499 (N_23499,N_12192,N_10575);
nor U23500 (N_23500,N_19969,N_16700);
nor U23501 (N_23501,N_12279,N_11070);
or U23502 (N_23502,N_17625,N_12584);
xor U23503 (N_23503,N_15950,N_15706);
xor U23504 (N_23504,N_19844,N_19371);
and U23505 (N_23505,N_19027,N_14748);
xor U23506 (N_23506,N_16244,N_19214);
nand U23507 (N_23507,N_19701,N_13731);
and U23508 (N_23508,N_13976,N_16828);
or U23509 (N_23509,N_17060,N_10784);
xor U23510 (N_23510,N_11164,N_13125);
or U23511 (N_23511,N_11765,N_13881);
and U23512 (N_23512,N_10754,N_18487);
xor U23513 (N_23513,N_17339,N_12996);
nor U23514 (N_23514,N_13790,N_10508);
nand U23515 (N_23515,N_18628,N_10534);
or U23516 (N_23516,N_10767,N_19207);
or U23517 (N_23517,N_16406,N_14073);
xnor U23518 (N_23518,N_16081,N_18805);
or U23519 (N_23519,N_19950,N_12777);
and U23520 (N_23520,N_18070,N_10677);
nand U23521 (N_23521,N_11286,N_15378);
nor U23522 (N_23522,N_10103,N_13550);
nor U23523 (N_23523,N_16116,N_13846);
nand U23524 (N_23524,N_19113,N_17587);
nor U23525 (N_23525,N_18161,N_13212);
or U23526 (N_23526,N_14687,N_14418);
nand U23527 (N_23527,N_11644,N_16373);
xor U23528 (N_23528,N_18771,N_17206);
and U23529 (N_23529,N_17588,N_14762);
nor U23530 (N_23530,N_11436,N_12616);
and U23531 (N_23531,N_17068,N_15097);
nor U23532 (N_23532,N_18774,N_15750);
xnor U23533 (N_23533,N_16905,N_18249);
or U23534 (N_23534,N_16249,N_14042);
and U23535 (N_23535,N_11917,N_13673);
nor U23536 (N_23536,N_19205,N_12109);
and U23537 (N_23537,N_19546,N_13694);
and U23538 (N_23538,N_10106,N_12702);
nor U23539 (N_23539,N_14637,N_11827);
nand U23540 (N_23540,N_17052,N_12198);
or U23541 (N_23541,N_16926,N_17885);
and U23542 (N_23542,N_18075,N_10868);
and U23543 (N_23543,N_15431,N_14888);
nor U23544 (N_23544,N_15336,N_14905);
and U23545 (N_23545,N_13833,N_19090);
and U23546 (N_23546,N_17786,N_16482);
nor U23547 (N_23547,N_11693,N_12943);
nor U23548 (N_23548,N_12797,N_18228);
nand U23549 (N_23549,N_17321,N_10917);
nand U23550 (N_23550,N_12570,N_17996);
or U23551 (N_23551,N_12154,N_15379);
or U23552 (N_23552,N_14679,N_17614);
nand U23553 (N_23553,N_18187,N_16503);
and U23554 (N_23554,N_17553,N_16291);
nand U23555 (N_23555,N_10425,N_18721);
nor U23556 (N_23556,N_15725,N_19476);
and U23557 (N_23557,N_17010,N_19374);
nand U23558 (N_23558,N_17358,N_11064);
xnor U23559 (N_23559,N_18241,N_16548);
or U23560 (N_23560,N_11750,N_10404);
nor U23561 (N_23561,N_17790,N_17911);
or U23562 (N_23562,N_12571,N_14908);
nand U23563 (N_23563,N_10659,N_13021);
and U23564 (N_23564,N_17342,N_16825);
nand U23565 (N_23565,N_18618,N_12725);
nand U23566 (N_23566,N_13636,N_14949);
nand U23567 (N_23567,N_18801,N_10798);
or U23568 (N_23568,N_18333,N_12558);
nor U23569 (N_23569,N_17103,N_11568);
nand U23570 (N_23570,N_17113,N_12827);
and U23571 (N_23571,N_15206,N_11677);
nand U23572 (N_23572,N_19954,N_11634);
xnor U23573 (N_23573,N_10182,N_19471);
nand U23574 (N_23574,N_11333,N_18595);
nor U23575 (N_23575,N_16211,N_11029);
or U23576 (N_23576,N_18481,N_16046);
nor U23577 (N_23577,N_10397,N_17564);
nand U23578 (N_23578,N_16370,N_17858);
or U23579 (N_23579,N_14638,N_11985);
xnor U23580 (N_23580,N_19557,N_19287);
and U23581 (N_23581,N_12761,N_12347);
nor U23582 (N_23582,N_14478,N_15286);
nand U23583 (N_23583,N_13156,N_18804);
xor U23584 (N_23584,N_13324,N_18231);
or U23585 (N_23585,N_13865,N_18633);
nor U23586 (N_23586,N_17758,N_12553);
nor U23587 (N_23587,N_18848,N_14793);
nor U23588 (N_23588,N_18105,N_10472);
nor U23589 (N_23589,N_15840,N_11148);
xnor U23590 (N_23590,N_16918,N_17639);
xnor U23591 (N_23591,N_10266,N_15534);
or U23592 (N_23592,N_14380,N_13308);
and U23593 (N_23593,N_16128,N_16182);
nor U23594 (N_23594,N_11574,N_17096);
xnor U23595 (N_23595,N_11549,N_19634);
and U23596 (N_23596,N_12378,N_15743);
nand U23597 (N_23597,N_13276,N_17804);
and U23598 (N_23598,N_13080,N_11687);
nor U23599 (N_23599,N_17745,N_10499);
or U23600 (N_23600,N_11709,N_15121);
nor U23601 (N_23601,N_11105,N_16049);
xnor U23602 (N_23602,N_10630,N_16555);
or U23603 (N_23603,N_15559,N_15132);
nor U23604 (N_23604,N_19204,N_10104);
or U23605 (N_23605,N_16831,N_12561);
nor U23606 (N_23606,N_14349,N_15890);
nor U23607 (N_23607,N_17189,N_18915);
nor U23608 (N_23608,N_17678,N_19075);
xor U23609 (N_23609,N_11976,N_11390);
and U23610 (N_23610,N_10811,N_12140);
nor U23611 (N_23611,N_11829,N_18681);
nor U23612 (N_23612,N_19681,N_14504);
nor U23613 (N_23613,N_11014,N_10164);
nor U23614 (N_23614,N_18359,N_10515);
xnor U23615 (N_23615,N_14222,N_15963);
nand U23616 (N_23616,N_15648,N_17825);
nand U23617 (N_23617,N_19834,N_19376);
and U23618 (N_23618,N_11589,N_19169);
xor U23619 (N_23619,N_10335,N_12358);
or U23620 (N_23620,N_15688,N_16107);
or U23621 (N_23621,N_17510,N_18271);
or U23622 (N_23622,N_17507,N_17038);
nor U23623 (N_23623,N_14587,N_11417);
xnor U23624 (N_23624,N_16963,N_12607);
xnor U23625 (N_23625,N_18136,N_13695);
or U23626 (N_23626,N_18110,N_10696);
or U23627 (N_23627,N_14396,N_13782);
xnor U23628 (N_23628,N_13961,N_18365);
and U23629 (N_23629,N_16955,N_14600);
and U23630 (N_23630,N_10154,N_13321);
or U23631 (N_23631,N_19705,N_15582);
xor U23632 (N_23632,N_17083,N_11569);
and U23633 (N_23633,N_17672,N_12999);
or U23634 (N_23634,N_11005,N_14233);
or U23635 (N_23635,N_17747,N_15455);
or U23636 (N_23636,N_10795,N_15549);
and U23637 (N_23637,N_19663,N_16341);
nor U23638 (N_23638,N_18409,N_13309);
or U23639 (N_23639,N_19703,N_19514);
or U23640 (N_23640,N_19897,N_19610);
xor U23641 (N_23641,N_11420,N_12251);
nor U23642 (N_23642,N_19919,N_17626);
or U23643 (N_23643,N_16577,N_12005);
xor U23644 (N_23644,N_11745,N_15521);
and U23645 (N_23645,N_18425,N_19176);
xor U23646 (N_23646,N_15778,N_11821);
nor U23647 (N_23647,N_13097,N_11957);
and U23648 (N_23648,N_12633,N_16236);
nor U23649 (N_23649,N_14288,N_11215);
nand U23650 (N_23650,N_11000,N_15161);
and U23651 (N_23651,N_16673,N_16592);
nor U23652 (N_23652,N_14203,N_12308);
nand U23653 (N_23653,N_18923,N_19808);
nor U23654 (N_23654,N_13969,N_19161);
nor U23655 (N_23655,N_19814,N_15944);
nand U23656 (N_23656,N_16259,N_10498);
nand U23657 (N_23657,N_11042,N_17823);
nor U23658 (N_23658,N_13953,N_17750);
or U23659 (N_23659,N_17784,N_17211);
nand U23660 (N_23660,N_16980,N_13718);
and U23661 (N_23661,N_16989,N_14121);
nand U23662 (N_23662,N_17854,N_10398);
or U23663 (N_23663,N_10883,N_16112);
nand U23664 (N_23664,N_11160,N_16578);
and U23665 (N_23665,N_14188,N_12287);
nand U23666 (N_23666,N_14265,N_11292);
nand U23667 (N_23667,N_13977,N_14520);
and U23668 (N_23668,N_18577,N_12830);
and U23669 (N_23669,N_14351,N_13958);
or U23670 (N_23670,N_13757,N_14521);
and U23671 (N_23671,N_19112,N_11063);
nor U23672 (N_23672,N_10477,N_18899);
and U23673 (N_23673,N_15355,N_10620);
nand U23674 (N_23674,N_13342,N_15623);
or U23675 (N_23675,N_13645,N_10119);
nor U23676 (N_23676,N_14915,N_12537);
xor U23677 (N_23677,N_11657,N_15802);
nand U23678 (N_23678,N_17685,N_12692);
and U23679 (N_23679,N_14851,N_16923);
and U23680 (N_23680,N_11399,N_16924);
nand U23681 (N_23681,N_18491,N_10006);
xor U23682 (N_23682,N_17661,N_11104);
and U23683 (N_23683,N_19778,N_18191);
nor U23684 (N_23684,N_19422,N_13103);
nand U23685 (N_23685,N_11091,N_14087);
nor U23686 (N_23686,N_10159,N_18251);
nand U23687 (N_23687,N_10364,N_11751);
xnor U23688 (N_23688,N_19874,N_11398);
nor U23689 (N_23689,N_15511,N_12061);
xnor U23690 (N_23690,N_12341,N_15729);
nor U23691 (N_23691,N_13440,N_15204);
xor U23692 (N_23692,N_18401,N_14760);
xnor U23693 (N_23693,N_11185,N_17274);
nor U23694 (N_23694,N_16990,N_12186);
xor U23695 (N_23695,N_15920,N_14529);
nor U23696 (N_23696,N_12346,N_14009);
and U23697 (N_23697,N_11007,N_11704);
or U23698 (N_23698,N_15409,N_14910);
nand U23699 (N_23699,N_13317,N_10548);
nor U23700 (N_23700,N_10325,N_16024);
nand U23701 (N_23701,N_17003,N_14160);
nor U23702 (N_23702,N_12970,N_16855);
or U23703 (N_23703,N_16508,N_10272);
or U23704 (N_23704,N_18654,N_16553);
and U23705 (N_23705,N_10581,N_15693);
xnor U23706 (N_23706,N_10160,N_12904);
nor U23707 (N_23707,N_18879,N_11151);
nor U23708 (N_23708,N_15553,N_18174);
xnor U23709 (N_23709,N_15240,N_11547);
nor U23710 (N_23710,N_14670,N_18861);
or U23711 (N_23711,N_12707,N_13618);
nand U23712 (N_23712,N_14239,N_11672);
xnor U23713 (N_23713,N_14045,N_11407);
nor U23714 (N_23714,N_12306,N_13838);
nor U23715 (N_23715,N_18584,N_17695);
nor U23716 (N_23716,N_17248,N_13190);
or U23717 (N_23717,N_12844,N_17259);
nand U23718 (N_23718,N_15568,N_11721);
nand U23719 (N_23719,N_17802,N_19039);
nand U23720 (N_23720,N_18067,N_13025);
and U23721 (N_23721,N_12263,N_13049);
nor U23722 (N_23722,N_17586,N_10424);
xor U23723 (N_23723,N_16337,N_13786);
nor U23724 (N_23724,N_10902,N_16579);
nand U23725 (N_23725,N_11500,N_10971);
xor U23726 (N_23726,N_10982,N_16547);
and U23727 (N_23727,N_12407,N_19472);
and U23728 (N_23728,N_16093,N_15001);
xnor U23729 (N_23729,N_17771,N_16080);
xor U23730 (N_23730,N_14718,N_12096);
or U23731 (N_23731,N_15331,N_10553);
nand U23732 (N_23732,N_11963,N_11921);
and U23733 (N_23733,N_12119,N_17579);
and U23734 (N_23734,N_19338,N_18664);
or U23735 (N_23735,N_10602,N_12842);
and U23736 (N_23736,N_19717,N_17078);
nand U23737 (N_23737,N_19431,N_18990);
and U23738 (N_23738,N_17871,N_17325);
and U23739 (N_23739,N_12519,N_10024);
nand U23740 (N_23740,N_17371,N_18012);
nand U23741 (N_23741,N_14467,N_13196);
or U23742 (N_23742,N_19253,N_12876);
or U23743 (N_23743,N_19046,N_19990);
or U23744 (N_23744,N_19028,N_15098);
or U23745 (N_23745,N_12762,N_11326);
or U23746 (N_23746,N_15848,N_18924);
nand U23747 (N_23747,N_13866,N_19052);
nor U23748 (N_23748,N_16641,N_10930);
and U23749 (N_23749,N_17537,N_16861);
and U23750 (N_23750,N_18396,N_10030);
nor U23751 (N_23751,N_13553,N_16275);
or U23752 (N_23752,N_15952,N_12611);
or U23753 (N_23753,N_18055,N_11246);
and U23754 (N_23754,N_15292,N_12207);
xnor U23755 (N_23755,N_14032,N_18751);
nand U23756 (N_23756,N_12956,N_10998);
and U23757 (N_23757,N_12206,N_14553);
and U23758 (N_23758,N_13583,N_17526);
or U23759 (N_23759,N_15430,N_14100);
or U23760 (N_23760,N_14513,N_17708);
or U23761 (N_23761,N_16451,N_13874);
nor U23762 (N_23762,N_10734,N_18248);
or U23763 (N_23763,N_17892,N_19519);
nand U23764 (N_23764,N_10373,N_11685);
nor U23765 (N_23765,N_13394,N_16830);
nor U23766 (N_23766,N_16771,N_18750);
or U23767 (N_23767,N_11818,N_12951);
or U23768 (N_23768,N_13010,N_13269);
or U23769 (N_23769,N_17118,N_19096);
or U23770 (N_23770,N_13535,N_11877);
xor U23771 (N_23771,N_12576,N_14136);
or U23772 (N_23772,N_15601,N_14502);
xor U23773 (N_23773,N_14573,N_17481);
nand U23774 (N_23774,N_11953,N_15319);
nor U23775 (N_23775,N_17314,N_19302);
or U23776 (N_23776,N_10377,N_15236);
and U23777 (N_23777,N_14613,N_16614);
nand U23778 (N_23778,N_18258,N_12652);
or U23779 (N_23779,N_17021,N_13917);
nor U23780 (N_23780,N_10421,N_19989);
and U23781 (N_23781,N_11050,N_10583);
xor U23782 (N_23782,N_11676,N_12574);
nor U23783 (N_23783,N_11058,N_19837);
xor U23784 (N_23784,N_19877,N_14724);
or U23785 (N_23785,N_19334,N_10317);
or U23786 (N_23786,N_10467,N_11766);
and U23787 (N_23787,N_16321,N_15423);
or U23788 (N_23788,N_19259,N_10362);
nor U23789 (N_23789,N_13717,N_10331);
nor U23790 (N_23790,N_17477,N_10666);
nor U23791 (N_23791,N_18100,N_14625);
nor U23792 (N_23792,N_17884,N_19802);
nor U23793 (N_23793,N_16293,N_15686);
or U23794 (N_23794,N_11362,N_13439);
nand U23795 (N_23795,N_11885,N_17094);
nand U23796 (N_23796,N_15667,N_14134);
and U23797 (N_23797,N_15516,N_16058);
and U23798 (N_23798,N_19600,N_17435);
or U23799 (N_23799,N_10607,N_14114);
nor U23800 (N_23800,N_10136,N_16653);
and U23801 (N_23801,N_11396,N_11510);
nor U23802 (N_23802,N_13978,N_11074);
or U23803 (N_23803,N_12946,N_19314);
xnor U23804 (N_23804,N_10400,N_19280);
xnor U23805 (N_23805,N_16248,N_15923);
nor U23806 (N_23806,N_17200,N_11365);
xnor U23807 (N_23807,N_15258,N_17421);
xor U23808 (N_23808,N_19748,N_12845);
and U23809 (N_23809,N_17453,N_12572);
and U23810 (N_23810,N_12155,N_15727);
or U23811 (N_23811,N_19390,N_18006);
xor U23812 (N_23812,N_15811,N_17439);
nand U23813 (N_23813,N_10709,N_15223);
xnor U23814 (N_23814,N_10578,N_17449);
nor U23815 (N_23815,N_10774,N_16775);
nor U23816 (N_23816,N_11840,N_14604);
or U23817 (N_23817,N_13436,N_16746);
xnor U23818 (N_23818,N_18863,N_19143);
or U23819 (N_23819,N_11110,N_10881);
nor U23820 (N_23820,N_13882,N_15229);
and U23821 (N_23821,N_17709,N_19986);
or U23822 (N_23822,N_12789,N_16187);
or U23823 (N_23823,N_19277,N_14546);
or U23824 (N_23824,N_19715,N_17889);
nor U23825 (N_23825,N_18040,N_13942);
nand U23826 (N_23826,N_14715,N_14864);
nor U23827 (N_23827,N_10069,N_15879);
nor U23828 (N_23828,N_17187,N_15135);
and U23829 (N_23829,N_14231,N_15205);
or U23830 (N_23830,N_19312,N_17988);
nand U23831 (N_23831,N_13690,N_16480);
nand U23832 (N_23832,N_13699,N_13781);
and U23833 (N_23833,N_14458,N_14767);
nor U23834 (N_23834,N_15759,N_16418);
nand U23835 (N_23835,N_12595,N_15898);
or U23836 (N_23836,N_15181,N_13907);
xor U23837 (N_23837,N_16545,N_15190);
nand U23838 (N_23838,N_17317,N_13178);
and U23839 (N_23839,N_18389,N_14439);
nor U23840 (N_23840,N_19997,N_12066);
and U23841 (N_23841,N_11154,N_15654);
nand U23842 (N_23842,N_18518,N_10903);
or U23843 (N_23843,N_16704,N_13239);
nand U23844 (N_23844,N_15722,N_14244);
nor U23845 (N_23845,N_14041,N_16755);
and U23846 (N_23846,N_10837,N_11869);
nor U23847 (N_23847,N_11822,N_10801);
xnor U23848 (N_23848,N_16086,N_14522);
and U23849 (N_23849,N_17814,N_10407);
xnor U23850 (N_23850,N_17684,N_11002);
nand U23851 (N_23851,N_15180,N_10821);
xnor U23852 (N_23852,N_12123,N_15442);
and U23853 (N_23853,N_10281,N_10457);
nand U23854 (N_23854,N_18164,N_15005);
xor U23855 (N_23855,N_13925,N_14592);
nand U23856 (N_23856,N_18973,N_18484);
xnor U23857 (N_23857,N_14099,N_18440);
nor U23858 (N_23858,N_15581,N_16930);
or U23859 (N_23859,N_11509,N_18221);
xnor U23860 (N_23860,N_13411,N_10861);
or U23861 (N_23861,N_19255,N_17209);
and U23862 (N_23862,N_15042,N_11447);
nor U23863 (N_23863,N_10478,N_16154);
nor U23864 (N_23864,N_13289,N_10960);
or U23865 (N_23865,N_15467,N_13926);
or U23866 (N_23866,N_15443,N_19733);
nor U23867 (N_23867,N_10519,N_12203);
or U23868 (N_23868,N_10753,N_12370);
and U23869 (N_23869,N_14764,N_15422);
and U23870 (N_23870,N_18181,N_14221);
xnor U23871 (N_23871,N_13333,N_12812);
nand U23872 (N_23872,N_16402,N_10076);
or U23873 (N_23873,N_15663,N_18685);
xor U23874 (N_23874,N_13443,N_11945);
or U23875 (N_23875,N_19261,N_17203);
and U23876 (N_23876,N_13034,N_14530);
nand U23877 (N_23877,N_17945,N_14126);
and U23878 (N_23878,N_17100,N_17332);
nor U23879 (N_23879,N_17603,N_19633);
or U23880 (N_23880,N_12491,N_10033);
nand U23881 (N_23881,N_12647,N_11434);
nor U23882 (N_23882,N_16971,N_13661);
nand U23883 (N_23883,N_14444,N_12397);
or U23884 (N_23884,N_15839,N_18226);
xnor U23885 (N_23885,N_18291,N_11024);
nand U23886 (N_23886,N_12240,N_12359);
nand U23887 (N_23887,N_15445,N_17413);
nor U23888 (N_23888,N_18983,N_17154);
nor U23889 (N_23889,N_19993,N_17993);
nor U23890 (N_23890,N_17044,N_17101);
nor U23891 (N_23891,N_13533,N_16447);
nor U23892 (N_23892,N_17346,N_14841);
or U23893 (N_23893,N_16263,N_15978);
or U23894 (N_23894,N_12506,N_13209);
xnor U23895 (N_23895,N_16732,N_15899);
and U23896 (N_23896,N_17763,N_17228);
xor U23897 (N_23897,N_17893,N_10451);
nand U23898 (N_23898,N_18138,N_10637);
xnor U23899 (N_23899,N_17875,N_18571);
nand U23900 (N_23900,N_17041,N_19723);
xor U23901 (N_23901,N_10593,N_19827);
nor U23902 (N_23902,N_18676,N_16163);
nand U23903 (N_23903,N_10417,N_17818);
and U23904 (N_23904,N_13929,N_12906);
xnor U23905 (N_23905,N_17079,N_10047);
xnor U23906 (N_23906,N_16979,N_11895);
or U23907 (N_23907,N_18169,N_19202);
xor U23908 (N_23908,N_13169,N_19291);
or U23909 (N_23909,N_12826,N_10486);
or U23910 (N_23910,N_10409,N_18256);
and U23911 (N_23911,N_16546,N_16322);
or U23912 (N_23912,N_18068,N_15817);
nand U23913 (N_23913,N_14445,N_17197);
nor U23914 (N_23914,N_16122,N_19083);
nand U23915 (N_23915,N_14161,N_14667);
and U23916 (N_23916,N_10992,N_19160);
xor U23917 (N_23917,N_17486,N_10422);
or U23918 (N_23918,N_12862,N_16022);
and U23919 (N_23919,N_16800,N_12431);
nor U23920 (N_23920,N_12780,N_13406);
nand U23921 (N_23921,N_11846,N_10286);
or U23922 (N_23922,N_10225,N_17388);
xor U23923 (N_23923,N_18996,N_17887);
and U23924 (N_23924,N_19555,N_17746);
and U23925 (N_23925,N_14211,N_16711);
or U23926 (N_23926,N_15176,N_10242);
or U23927 (N_23927,N_19895,N_17231);
and U23928 (N_23928,N_15054,N_12264);
nand U23929 (N_23929,N_11066,N_10470);
xnor U23930 (N_23930,N_18150,N_10580);
nor U23931 (N_23931,N_19172,N_12127);
and U23932 (N_23932,N_14300,N_13972);
nor U23933 (N_23933,N_11243,N_10067);
xor U23934 (N_23934,N_11454,N_18857);
xor U23935 (N_23935,N_15160,N_13462);
nand U23936 (N_23936,N_14319,N_17237);
nor U23937 (N_23937,N_13809,N_14863);
nand U23938 (N_23938,N_10792,N_19960);
xnor U23939 (N_23939,N_14127,N_18888);
or U23940 (N_23940,N_13290,N_16763);
or U23941 (N_23941,N_14272,N_18842);
and U23942 (N_23942,N_11400,N_10491);
nand U23943 (N_23943,N_17316,N_13076);
nand U23944 (N_23944,N_16326,N_18198);
xor U23945 (N_23945,N_13379,N_19357);
or U23946 (N_23946,N_10569,N_12977);
nand U23947 (N_23947,N_19911,N_12213);
nor U23948 (N_23948,N_17046,N_17225);
nor U23949 (N_23949,N_18964,N_16690);
nor U23950 (N_23950,N_10585,N_11194);
nor U23951 (N_23951,N_15227,N_11992);
nor U23952 (N_23952,N_10093,N_13174);
xor U23953 (N_23953,N_14919,N_15627);
or U23954 (N_23954,N_18355,N_17085);
xor U23955 (N_23955,N_12325,N_15842);
nor U23956 (N_23956,N_19629,N_16909);
nor U23957 (N_23957,N_19662,N_13813);
nand U23958 (N_23958,N_17422,N_17233);
xor U23959 (N_23959,N_19921,N_15495);
and U23960 (N_23960,N_12778,N_14425);
or U23961 (N_23961,N_12212,N_14683);
and U23962 (N_23962,N_13996,N_19104);
nor U23963 (N_23963,N_11176,N_17123);
or U23964 (N_23964,N_17032,N_14576);
xnor U23965 (N_23965,N_11464,N_10874);
or U23966 (N_23966,N_13752,N_12221);
xor U23967 (N_23967,N_11340,N_11758);
nor U23968 (N_23968,N_12413,N_19404);
or U23969 (N_23969,N_10221,N_12794);
nor U23970 (N_23970,N_11609,N_16738);
and U23971 (N_23971,N_18242,N_11082);
xor U23972 (N_23972,N_15151,N_13035);
nand U23973 (N_23973,N_15613,N_17987);
nand U23974 (N_23974,N_19375,N_18725);
or U23975 (N_23975,N_13451,N_16933);
nand U23976 (N_23976,N_10835,N_17431);
or U23977 (N_23977,N_19893,N_12004);
or U23978 (N_23978,N_14704,N_11394);
xnor U23979 (N_23979,N_10452,N_19272);
xor U23980 (N_23980,N_16170,N_19669);
and U23981 (N_23981,N_15122,N_19140);
xnor U23982 (N_23982,N_19601,N_18153);
nand U23983 (N_23983,N_11519,N_11858);
nand U23984 (N_23984,N_12403,N_13732);
nor U23985 (N_23985,N_13455,N_13221);
xor U23986 (N_23986,N_11629,N_13447);
or U23987 (N_23987,N_18261,N_13247);
xnor U23988 (N_23988,N_10192,N_15326);
nand U23989 (N_23989,N_15764,N_16960);
nor U23990 (N_23990,N_17173,N_10547);
xnor U23991 (N_23991,N_17409,N_13939);
nand U23992 (N_23992,N_14470,N_10090);
nand U23993 (N_23993,N_10290,N_18652);
and U23994 (N_23994,N_15653,N_16692);
nor U23995 (N_23995,N_15170,N_15637);
or U23996 (N_23996,N_12961,N_14307);
and U23997 (N_23997,N_13358,N_16180);
nor U23998 (N_23998,N_18141,N_18945);
or U23999 (N_23999,N_16796,N_14043);
nand U24000 (N_24000,N_10733,N_15344);
nor U24001 (N_24001,N_17979,N_11112);
xnor U24002 (N_24002,N_17369,N_15883);
xor U24003 (N_24003,N_12851,N_16878);
nand U24004 (N_24004,N_11348,N_14148);
nor U24005 (N_24005,N_15494,N_14303);
nand U24006 (N_24006,N_15271,N_14736);
nor U24007 (N_24007,N_15783,N_19030);
nand U24008 (N_24008,N_17141,N_17971);
or U24009 (N_24009,N_16887,N_19011);
nor U24010 (N_24010,N_18854,N_18126);
and U24011 (N_24011,N_11899,N_17931);
nor U24012 (N_24012,N_13616,N_12991);
nor U24013 (N_24013,N_16157,N_16981);
xnor U24014 (N_24014,N_13762,N_12412);
nor U24015 (N_24015,N_10369,N_16936);
or U24016 (N_24016,N_17460,N_12406);
nand U24017 (N_24017,N_10312,N_18741);
nand U24018 (N_24018,N_14611,N_10042);
or U24019 (N_24019,N_11820,N_16039);
and U24020 (N_24020,N_17533,N_14046);
and U24021 (N_24021,N_15641,N_15067);
or U24022 (N_24022,N_16492,N_19585);
xnor U24023 (N_24023,N_15924,N_15343);
nand U24024 (N_24024,N_10055,N_19190);
nor U24025 (N_24025,N_15004,N_18611);
nor U24026 (N_24026,N_10034,N_18133);
and U24027 (N_24027,N_17128,N_13264);
and U24028 (N_24028,N_17491,N_17856);
nand U24029 (N_24029,N_12721,N_17864);
nor U24030 (N_24030,N_15801,N_11375);
and U24031 (N_24031,N_15030,N_18265);
and U24032 (N_24032,N_19215,N_12175);
and U24033 (N_24033,N_15021,N_16723);
or U24034 (N_24034,N_19809,N_15148);
or U24035 (N_24035,N_14367,N_10000);
nor U24036 (N_24036,N_16466,N_12113);
xor U24037 (N_24037,N_19442,N_14951);
or U24038 (N_24038,N_16464,N_12625);
and U24039 (N_24039,N_18464,N_11312);
xnor U24040 (N_24040,N_18497,N_11837);
nor U24041 (N_24041,N_17888,N_18674);
and U24042 (N_24042,N_16351,N_10939);
and U24043 (N_24043,N_18942,N_15998);
or U24044 (N_24044,N_19853,N_14827);
nand U24045 (N_24045,N_19005,N_17657);
or U24046 (N_24046,N_16268,N_12027);
nor U24047 (N_24047,N_12573,N_13341);
nor U24048 (N_24048,N_11701,N_15044);
nand U24049 (N_24049,N_15294,N_14813);
nor U24050 (N_24050,N_14243,N_15964);
and U24051 (N_24051,N_11484,N_19608);
or U24052 (N_24052,N_13559,N_19238);
or U24053 (N_24053,N_15639,N_17689);
and U24054 (N_24054,N_17081,N_13386);
xor U24055 (N_24055,N_17045,N_15515);
or U24056 (N_24056,N_18894,N_19649);
nand U24057 (N_24057,N_11227,N_13085);
xor U24058 (N_24058,N_12512,N_17630);
xor U24059 (N_24059,N_18736,N_13760);
xnor U24060 (N_24060,N_16899,N_15058);
and U24061 (N_24061,N_10805,N_12425);
xnor U24062 (N_24062,N_15679,N_19309);
nand U24063 (N_24063,N_15833,N_17382);
or U24064 (N_24064,N_10526,N_12983);
xor U24065 (N_24065,N_11531,N_14725);
xnor U24066 (N_24066,N_12711,N_14743);
or U24067 (N_24067,N_10536,N_10190);
and U24068 (N_24068,N_11046,N_13858);
or U24069 (N_24069,N_13725,N_17429);
or U24070 (N_24070,N_16822,N_17106);
xnor U24071 (N_24071,N_13422,N_19250);
nand U24072 (N_24072,N_14568,N_17386);
or U24073 (N_24073,N_19762,N_19003);
and U24074 (N_24074,N_19224,N_16357);
and U24075 (N_24075,N_11290,N_18195);
nor U24076 (N_24076,N_16654,N_19001);
or U24077 (N_24077,N_15052,N_12404);
and U24078 (N_24078,N_19316,N_18107);
and U24079 (N_24079,N_18844,N_11034);
nand U24080 (N_24080,N_10046,N_18532);
or U24081 (N_24081,N_17423,N_10778);
nand U24082 (N_24082,N_16522,N_12560);
and U24083 (N_24083,N_19229,N_13811);
or U24084 (N_24084,N_15984,N_15109);
nand U24085 (N_24085,N_18225,N_15983);
or U24086 (N_24086,N_15413,N_18089);
nor U24087 (N_24087,N_11102,N_10230);
nor U24088 (N_24088,N_12626,N_18102);
and U24089 (N_24089,N_18037,N_15071);
nor U24090 (N_24090,N_10260,N_19666);
or U24091 (N_24091,N_11143,N_10586);
nor U24092 (N_24092,N_11440,N_15209);
or U24093 (N_24093,N_10557,N_15584);
or U24094 (N_24094,N_13100,N_19742);
or U24095 (N_24095,N_19642,N_15388);
or U24096 (N_24096,N_16937,N_19118);
xnor U24097 (N_24097,N_19888,N_13108);
nand U24098 (N_24098,N_14788,N_14578);
nand U24099 (N_24099,N_18351,N_13396);
or U24100 (N_24100,N_10542,N_17287);
xnor U24101 (N_24101,N_17313,N_10117);
or U24102 (N_24102,N_10697,N_10807);
and U24103 (N_24103,N_16752,N_13137);
or U24104 (N_24104,N_11526,N_16420);
xor U24105 (N_24105,N_18553,N_12833);
or U24106 (N_24106,N_14954,N_10333);
nand U24107 (N_24107,N_10771,N_18768);
xor U24108 (N_24108,N_12053,N_13713);
or U24109 (N_24109,N_16707,N_15124);
and U24110 (N_24110,N_16593,N_14006);
nor U24111 (N_24111,N_16194,N_17450);
nand U24112 (N_24112,N_19281,N_14301);
nor U24113 (N_24113,N_18504,N_16127);
or U24114 (N_24114,N_14968,N_10315);
nor U24115 (N_24115,N_11602,N_17030);
nor U24116 (N_24116,N_11767,N_11282);
nor U24117 (N_24117,N_11380,N_13397);
nor U24118 (N_24118,N_11036,N_19896);
or U24119 (N_24119,N_19074,N_15200);
nand U24120 (N_24120,N_10216,N_10368);
nand U24121 (N_24121,N_17395,N_16448);
xnor U24122 (N_24122,N_16270,N_10984);
nand U24123 (N_24123,N_11732,N_17035);
nand U24124 (N_24124,N_13001,N_10015);
or U24125 (N_24125,N_14545,N_10653);
and U24126 (N_24126,N_15092,N_10844);
xnor U24127 (N_24127,N_10961,N_15106);
xnor U24128 (N_24128,N_18722,N_10228);
nand U24129 (N_24129,N_10155,N_11328);
nand U24130 (N_24130,N_14690,N_11242);
xor U24131 (N_24131,N_14624,N_18753);
nor U24132 (N_24132,N_13837,N_15507);
and U24133 (N_24133,N_16267,N_15684);
nor U24134 (N_24134,N_18428,N_18312);
nand U24135 (N_24135,N_19811,N_19774);
nor U24136 (N_24136,N_19434,N_11273);
or U24137 (N_24137,N_14068,N_15927);
and U24138 (N_24138,N_15550,N_15429);
nor U24139 (N_24139,N_17606,N_16338);
and U24140 (N_24140,N_17163,N_17397);
and U24141 (N_24141,N_19862,N_10243);
and U24142 (N_24142,N_16300,N_10506);
and U24143 (N_24143,N_12443,N_17167);
or U24144 (N_24144,N_17924,N_14580);
xnor U24145 (N_24145,N_12656,N_19405);
nor U24146 (N_24146,N_14185,N_12613);
and U24147 (N_24147,N_11349,N_15796);
nand U24148 (N_24148,N_15317,N_12339);
and U24149 (N_24149,N_10126,N_10775);
nor U24150 (N_24150,N_14885,N_17670);
and U24151 (N_24151,N_14784,N_18031);
xnor U24152 (N_24152,N_14336,N_11971);
and U24153 (N_24153,N_16902,N_11270);
and U24154 (N_24154,N_15943,N_15674);
and U24155 (N_24155,N_11054,N_15032);
nor U24156 (N_24156,N_15285,N_15399);
nor U24157 (N_24157,N_18041,N_11578);
nor U24158 (N_24158,N_11419,N_14429);
xor U24159 (N_24159,N_15016,N_17404);
xor U24160 (N_24160,N_11724,N_16862);
nand U24161 (N_24161,N_17826,N_11315);
xnor U24162 (N_24162,N_16975,N_10773);
nor U24163 (N_24163,N_14572,N_19538);
or U24164 (N_24164,N_13754,N_15062);
nor U24165 (N_24165,N_16453,N_18345);
xor U24166 (N_24166,N_13620,N_10011);
xnor U24167 (N_24167,N_11521,N_19493);
nor U24168 (N_24168,N_19616,N_15716);
xor U24169 (N_24169,N_10401,N_12975);
and U24170 (N_24170,N_16016,N_10259);
xnor U24171 (N_24171,N_12849,N_15120);
xor U24172 (N_24172,N_16210,N_19414);
and U24173 (N_24173,N_12624,N_10967);
nand U24174 (N_24174,N_17692,N_19385);
nor U24175 (N_24175,N_18330,N_14340);
xnor U24176 (N_24176,N_11401,N_18630);
nand U24177 (N_24177,N_17042,N_17137);
or U24178 (N_24178,N_16392,N_12803);
nand U24179 (N_24179,N_12831,N_14497);
nor U24180 (N_24180,N_16708,N_18035);
nor U24181 (N_24181,N_11162,N_15468);
xor U24182 (N_24182,N_17719,N_12078);
nor U24183 (N_24183,N_14255,N_14777);
nand U24184 (N_24184,N_18391,N_16125);
xnor U24185 (N_24185,N_14965,N_14452);
xor U24186 (N_24186,N_13631,N_17368);
nor U24187 (N_24187,N_14151,N_12731);
or U24188 (N_24188,N_14424,N_18028);
and U24189 (N_24189,N_15027,N_18057);
and U24190 (N_24190,N_12903,N_15045);
nor U24191 (N_24191,N_19926,N_10812);
nand U24192 (N_24192,N_12910,N_16450);
nor U24193 (N_24193,N_17306,N_18092);
or U24194 (N_24194,N_11848,N_12754);
nor U24195 (N_24195,N_15925,N_10075);
and U24196 (N_24196,N_14144,N_13625);
nor U24197 (N_24197,N_12312,N_10144);
nor U24198 (N_24198,N_18565,N_16176);
xor U24199 (N_24199,N_10724,N_11880);
xnor U24200 (N_24200,N_11236,N_18622);
nand U24201 (N_24201,N_16712,N_11636);
or U24202 (N_24202,N_13689,N_13260);
nor U24203 (N_24203,N_18573,N_18735);
nand U24204 (N_24204,N_15832,N_19270);
and U24205 (N_24205,N_14923,N_17370);
xor U24206 (N_24206,N_12102,N_12661);
xnor U24207 (N_24207,N_14098,N_17827);
or U24208 (N_24208,N_10999,N_16852);
or U24209 (N_24209,N_11660,N_18369);
or U24210 (N_24210,N_11573,N_12547);
or U24211 (N_24211,N_14626,N_16253);
or U24212 (N_24212,N_12566,N_13229);
nand U24213 (N_24213,N_18121,N_11993);
xor U24214 (N_24214,N_19675,N_18908);
nand U24215 (N_24215,N_14428,N_12599);
and U24216 (N_24216,N_11824,N_14675);
and U24217 (N_24217,N_19536,N_18022);
nand U24218 (N_24218,N_17327,N_14740);
nor U24219 (N_24219,N_12565,N_12861);
xnor U24220 (N_24220,N_12377,N_17680);
xnor U24221 (N_24221,N_15704,N_19079);
nand U24222 (N_24222,N_18400,N_15540);
nand U24223 (N_24223,N_17199,N_13986);
xor U24224 (N_24224,N_10008,N_12320);
and U24225 (N_24225,N_15948,N_19985);
nor U24226 (N_24226,N_11694,N_12380);
nor U24227 (N_24227,N_19345,N_13427);
and U24228 (N_24228,N_14997,N_13257);
or U24229 (N_24229,N_14004,N_14852);
or U24230 (N_24230,N_17686,N_16156);
or U24231 (N_24231,N_17263,N_12680);
xor U24232 (N_24232,N_19037,N_14564);
xor U24233 (N_24233,N_11726,N_10001);
or U24234 (N_24234,N_18295,N_15640);
or U24235 (N_24235,N_15547,N_16192);
xor U24236 (N_24236,N_13230,N_11597);
or U24237 (N_24237,N_18583,N_18837);
or U24238 (N_24238,N_15610,N_13051);
or U24239 (N_24239,N_17559,N_14013);
nor U24240 (N_24240,N_17659,N_12146);
xor U24241 (N_24241,N_13596,N_16265);
or U24242 (N_24242,N_12234,N_19686);
nor U24243 (N_24243,N_18902,N_11506);
and U24244 (N_24244,N_14526,N_10794);
and U24245 (N_24245,N_14142,N_16716);
nor U24246 (N_24246,N_19341,N_13068);
nand U24247 (N_24247,N_12922,N_15685);
or U24248 (N_24248,N_12676,N_11760);
or U24249 (N_24249,N_16138,N_16051);
nand U24250 (N_24250,N_11965,N_10261);
or U24251 (N_24251,N_16604,N_18656);
nor U24252 (N_24252,N_12496,N_13870);
nand U24253 (N_24253,N_18871,N_11594);
and U24254 (N_24254,N_11907,N_15129);
and U24255 (N_24255,N_13261,N_14678);
and U24256 (N_24256,N_17350,N_19002);
xnor U24257 (N_24257,N_15632,N_14872);
nand U24258 (N_24258,N_17835,N_11560);
xor U24259 (N_24259,N_17918,N_18285);
and U24260 (N_24260,N_10831,N_11739);
nand U24261 (N_24261,N_16570,N_17405);
or U24262 (N_24262,N_18916,N_19479);
nand U24263 (N_24263,N_17105,N_16368);
nand U24264 (N_24264,N_12497,N_16939);
and U24265 (N_24265,N_11346,N_11272);
and U24266 (N_24266,N_17921,N_17984);
xnor U24267 (N_24267,N_10328,N_16487);
and U24268 (N_24268,N_11475,N_19413);
or U24269 (N_24269,N_14894,N_17278);
nor U24270 (N_24270,N_18663,N_12533);
nand U24271 (N_24271,N_19317,N_16780);
and U24272 (N_24272,N_17086,N_14879);
or U24273 (N_24273,N_17433,N_10480);
or U24274 (N_24274,N_19266,N_11652);
nand U24275 (N_24275,N_16602,N_18134);
nor U24276 (N_24276,N_14216,N_11267);
and U24277 (N_24277,N_16032,N_13826);
nor U24278 (N_24278,N_13401,N_13604);
and U24279 (N_24279,N_14946,N_13682);
nand U24280 (N_24280,N_19125,N_15673);
nor U24281 (N_24281,N_19171,N_14702);
nor U24282 (N_24282,N_14699,N_17567);
nand U24283 (N_24283,N_14066,N_10760);
nor U24284 (N_24284,N_13248,N_10341);
nor U24285 (N_24285,N_16687,N_18336);
or U24286 (N_24286,N_10018,N_17324);
or U24287 (N_24287,N_16721,N_12223);
nand U24288 (N_24288,N_14928,N_12825);
and U24289 (N_24289,N_14312,N_11096);
nor U24290 (N_24290,N_14313,N_12726);
and U24291 (N_24291,N_18446,N_10937);
or U24292 (N_24292,N_17513,N_10768);
nand U24293 (N_24293,N_14837,N_13445);
nand U24294 (N_24294,N_16085,N_17978);
xor U24295 (N_24295,N_11713,N_14174);
nor U24296 (N_24296,N_17185,N_10079);
xor U24297 (N_24297,N_14796,N_14842);
nand U24298 (N_24298,N_14059,N_12295);
or U24299 (N_24299,N_19522,N_11079);
or U24300 (N_24300,N_18718,N_18807);
xor U24301 (N_24301,N_13437,N_12581);
xor U24302 (N_24302,N_10040,N_13687);
and U24303 (N_24303,N_18946,N_17416);
or U24304 (N_24304,N_14744,N_12033);
nor U24305 (N_24305,N_13056,N_15866);
or U24306 (N_24306,N_15741,N_10986);
nand U24307 (N_24307,N_18021,N_11423);
nand U24308 (N_24308,N_10150,N_17089);
or U24309 (N_24309,N_18217,N_17271);
nor U24310 (N_24310,N_13246,N_19793);
and U24311 (N_24311,N_16638,N_10818);
xor U24312 (N_24312,N_14814,N_14868);
xor U24313 (N_24313,N_10294,N_11898);
or U24314 (N_24314,N_10977,N_16953);
or U24315 (N_24315,N_19798,N_13118);
and U24316 (N_24316,N_17319,N_14419);
nand U24317 (N_24317,N_12427,N_13020);
and U24318 (N_24318,N_10750,N_13763);
xnor U24319 (N_24319,N_11980,N_16667);
and U24320 (N_24320,N_19755,N_19597);
and U24321 (N_24321,N_14236,N_14304);
nor U24322 (N_24322,N_15889,N_14995);
or U24323 (N_24323,N_12457,N_19824);
xnor U24324 (N_24324,N_16513,N_14541);
xnor U24325 (N_24325,N_11047,N_14197);
nand U24326 (N_24326,N_11224,N_19635);
and U24327 (N_24327,N_10094,N_11188);
xnor U24328 (N_24328,N_16781,N_11890);
xnor U24329 (N_24329,N_16904,N_15556);
nor U24330 (N_24330,N_10483,N_10147);
xnor U24331 (N_24331,N_19069,N_18462);
or U24332 (N_24332,N_10990,N_16751);
nand U24333 (N_24333,N_17289,N_10708);
xnor U24334 (N_24334,N_11118,N_14598);
xor U24335 (N_24335,N_19590,N_11854);
and U24336 (N_24336,N_12445,N_18432);
nor U24337 (N_24337,N_16286,N_14409);
and U24338 (N_24338,N_18606,N_12920);
and U24339 (N_24339,N_13018,N_12135);
nand U24340 (N_24340,N_18208,N_15712);
or U24341 (N_24341,N_19419,N_13005);
or U24342 (N_24342,N_12575,N_13305);
or U24343 (N_24343,N_10269,N_15304);
or U24344 (N_24344,N_14398,N_14836);
and U24345 (N_24345,N_12674,N_16274);
nand U24346 (N_24346,N_18433,N_13818);
or U24347 (N_24347,N_15907,N_13465);
nand U24348 (N_24348,N_10681,N_16696);
xor U24349 (N_24349,N_14695,N_19177);
nor U24350 (N_24350,N_13371,N_18383);
nor U24351 (N_24351,N_12311,N_10577);
xor U24352 (N_24352,N_15153,N_14697);
or U24353 (N_24353,N_10322,N_13895);
or U24354 (N_24354,N_11754,N_16590);
or U24355 (N_24355,N_14485,N_15493);
nand U24356 (N_24356,N_16992,N_12314);
nor U24357 (N_24357,N_11939,N_13888);
nor U24358 (N_24358,N_14914,N_14730);
nand U24359 (N_24359,N_12892,N_13541);
and U24360 (N_24360,N_18971,N_14430);
nand U24361 (N_24361,N_11405,N_12259);
and U24362 (N_24362,N_17972,N_16393);
and U24363 (N_24363,N_19899,N_14828);
and U24364 (N_24364,N_17754,N_12026);
nor U24365 (N_24365,N_11115,N_18938);
nor U24366 (N_24366,N_13249,N_17765);
and U24367 (N_24367,N_14756,N_16999);
and U24368 (N_24368,N_12858,N_18302);
or U24369 (N_24369,N_13365,N_18890);
xnor U24370 (N_24370,N_14651,N_18034);
nor U24371 (N_24371,N_11853,N_10233);
xnor U24372 (N_24372,N_11146,N_18375);
xor U24373 (N_24373,N_13676,N_11986);
or U24374 (N_24374,N_10063,N_13223);
nand U24375 (N_24375,N_18742,N_12834);
or U24376 (N_24376,N_18748,N_19623);
nand U24377 (N_24377,N_13415,N_15710);
nor U24378 (N_24378,N_11979,N_10393);
and U24379 (N_24379,N_17883,N_15501);
or U24380 (N_24380,N_16474,N_13367);
nor U24381 (N_24381,N_18417,N_14575);
and U24382 (N_24382,N_19745,N_18950);
or U24383 (N_24383,N_16957,N_10229);
nand U24384 (N_24384,N_10296,N_12749);
nor U24385 (N_24385,N_10146,N_13611);
nand U24386 (N_24386,N_18458,N_15089);
nor U24387 (N_24387,N_12492,N_13266);
nand U24388 (N_24388,N_13780,N_14959);
xnor U24389 (N_24389,N_18282,N_12296);
nand U24390 (N_24390,N_17832,N_19987);
or U24391 (N_24391,N_17471,N_18064);
nor U24392 (N_24392,N_13015,N_16794);
nor U24393 (N_24393,N_16968,N_12200);
nand U24394 (N_24394,N_14893,N_15518);
nand U24395 (N_24395,N_12495,N_18610);
nor U24396 (N_24396,N_12040,N_12587);
xnor U24397 (N_24397,N_11201,N_17651);
or U24398 (N_24398,N_18078,N_12029);
and U24399 (N_24399,N_12034,N_11961);
nor U24400 (N_24400,N_14769,N_12439);
or U24401 (N_24401,N_11712,N_13328);
nand U24402 (N_24402,N_16166,N_12832);
and U24403 (N_24403,N_12591,N_11257);
or U24404 (N_24404,N_14953,N_15976);
xor U24405 (N_24405,N_16556,N_19305);
and U24406 (N_24406,N_17762,N_16458);
nor U24407 (N_24407,N_19022,N_16661);
nor U24408 (N_24408,N_19944,N_14128);
and U24409 (N_24409,N_11731,N_18877);
nor U24410 (N_24410,N_18769,N_12804);
and U24411 (N_24411,N_13092,N_10211);
xnor U24412 (N_24412,N_16766,N_14492);
or U24413 (N_24413,N_16617,N_16344);
or U24414 (N_24414,N_14614,N_12477);
xnor U24415 (N_24415,N_16225,N_12285);
nand U24416 (N_24416,N_12693,N_17660);
nand U24417 (N_24417,N_16471,N_15586);
and U24418 (N_24418,N_13721,N_17779);
or U24419 (N_24419,N_15580,N_15779);
or U24420 (N_24420,N_15358,N_17012);
nor U24421 (N_24421,N_11908,N_18080);
nand U24422 (N_24422,N_16317,N_15587);
or U24423 (N_24423,N_12853,N_19815);
or U24424 (N_24424,N_18424,N_13656);
nand U24425 (N_24425,N_11650,N_16243);
nor U24426 (N_24426,N_15836,N_10097);
nor U24427 (N_24427,N_16765,N_11664);
xnor U24428 (N_24428,N_18535,N_18059);
nor U24429 (N_24429,N_13946,N_13215);
xnor U24430 (N_24430,N_15456,N_18498);
nor U24431 (N_24431,N_18192,N_10691);
xor U24432 (N_24432,N_11725,N_11438);
and U24433 (N_24433,N_11293,N_16119);
nand U24434 (N_24434,N_16079,N_10497);
and U24435 (N_24435,N_10437,N_18515);
or U24436 (N_24436,N_15528,N_17538);
nor U24437 (N_24437,N_12871,N_15489);
nor U24438 (N_24438,N_19012,N_17145);
or U24439 (N_24439,N_11198,N_18451);
and U24440 (N_24440,N_17260,N_18604);
xor U24441 (N_24441,N_15790,N_16072);
and U24442 (N_24442,N_19387,N_11785);
and U24443 (N_24443,N_14291,N_10111);
nor U24444 (N_24444,N_12344,N_12706);
xnor U24445 (N_24445,N_15911,N_19551);
or U24446 (N_24446,N_19700,N_18992);
nand U24447 (N_24447,N_17201,N_17493);
nor U24448 (N_24448,N_18802,N_15830);
nor U24449 (N_24449,N_17023,N_15733);
and U24450 (N_24450,N_18575,N_18422);
nor U24451 (N_24451,N_10276,N_10594);
or U24452 (N_24452,N_18029,N_13224);
or U24453 (N_24453,N_17942,N_14379);
or U24454 (N_24454,N_12051,N_12787);
or U24455 (N_24455,N_10958,N_15775);
or U24456 (N_24456,N_19382,N_13126);
nor U24457 (N_24457,N_10339,N_12921);
or U24458 (N_24458,N_19245,N_11661);
and U24459 (N_24459,N_15392,N_15744);
nand U24460 (N_24460,N_11995,N_15497);
nor U24461 (N_24461,N_18898,N_10503);
nor U24462 (N_24462,N_12286,N_13405);
or U24463 (N_24463,N_16814,N_12355);
nor U24464 (N_24464,N_19146,N_16605);
and U24465 (N_24465,N_18695,N_15082);
xnor U24466 (N_24466,N_18460,N_18106);
xnor U24467 (N_24467,N_10611,N_19626);
xnor U24468 (N_24468,N_13277,N_13088);
or U24469 (N_24469,N_17569,N_14109);
xnor U24470 (N_24470,N_16496,N_15585);
and U24471 (N_24471,N_18637,N_15011);
or U24472 (N_24472,N_17583,N_15426);
and U24473 (N_24473,N_16742,N_12258);
xnor U24474 (N_24474,N_12390,N_12548);
and U24475 (N_24475,N_18505,N_18113);
and U24476 (N_24476,N_18554,N_10087);
nor U24477 (N_24477,N_10555,N_17359);
or U24478 (N_24478,N_14665,N_16069);
nor U24479 (N_24479,N_11856,N_12174);
or U24480 (N_24480,N_18294,N_12747);
xnor U24481 (N_24481,N_10850,N_10676);
and U24482 (N_24482,N_15868,N_18738);
nor U24483 (N_24483,N_10731,N_11347);
xor U24484 (N_24484,N_13726,N_17057);
or U24485 (N_24485,N_17065,N_10966);
xnor U24486 (N_24486,N_18947,N_15398);
nand U24487 (N_24487,N_10714,N_15084);
xor U24488 (N_24488,N_11836,N_14909);
xnor U24489 (N_24489,N_12024,N_14717);
nand U24490 (N_24490,N_10721,N_11920);
xnor U24491 (N_24491,N_15617,N_17866);
nor U24492 (N_24492,N_12925,N_15650);
nor U24493 (N_24493,N_17748,N_11459);
xor U24494 (N_24494,N_18665,N_17800);
and U24495 (N_24495,N_14734,N_10758);
xnor U24496 (N_24496,N_19481,N_10270);
nor U24497 (N_24497,N_16595,N_11468);
and U24498 (N_24498,N_16434,N_13091);
xnor U24499 (N_24499,N_19560,N_15035);
nand U24500 (N_24500,N_19714,N_15464);
nor U24501 (N_24501,N_11913,N_10799);
nand U24502 (N_24502,N_12784,N_11252);
or U24503 (N_24503,N_18166,N_14268);
and U24504 (N_24504,N_14089,N_16524);
nand U24505 (N_24505,N_14594,N_17705);
nor U24506 (N_24506,N_15524,N_14295);
or U24507 (N_24507,N_16576,N_14825);
nand U24508 (N_24508,N_13402,N_12800);
and U24509 (N_24509,N_13208,N_19360);
xnor U24510 (N_24510,N_16361,N_15048);
nor U24511 (N_24511,N_17870,N_15174);
or U24512 (N_24512,N_16088,N_11325);
xnor U24513 (N_24513,N_17623,N_10839);
and U24514 (N_24514,N_16816,N_14984);
and U24515 (N_24515,N_12079,N_18011);
nand U24516 (N_24516,N_18455,N_17277);
nor U24517 (N_24517,N_12256,N_11887);
or U24518 (N_24518,N_17291,N_14394);
nand U24519 (N_24519,N_12336,N_17451);
and U24520 (N_24520,N_10439,N_12934);
xor U24521 (N_24521,N_19235,N_16713);
xor U24522 (N_24522,N_10285,N_16013);
nor U24523 (N_24523,N_19930,N_16724);
nor U24524 (N_24524,N_12919,N_11073);
and U24525 (N_24525,N_19482,N_15571);
nand U24526 (N_24526,N_18372,N_10921);
and U24527 (N_24527,N_11406,N_13745);
or U24528 (N_24528,N_19331,N_16188);
and U24529 (N_24529,N_11910,N_17604);
nand U24530 (N_24530,N_18816,N_10389);
or U24531 (N_24531,N_13902,N_17104);
and U24532 (N_24532,N_13898,N_11287);
and U24533 (N_24533,N_11108,N_14804);
nand U24534 (N_24534,N_15193,N_16843);
nand U24535 (N_24535,N_13480,N_16871);
and U24536 (N_24536,N_12666,N_14240);
or U24537 (N_24537,N_13709,N_17777);
and U24538 (N_24538,N_12309,N_17340);
xnor U24539 (N_24539,N_19665,N_15711);
and U24540 (N_24540,N_17896,N_19855);
and U24541 (N_24541,N_14994,N_19975);
nand U24542 (N_24542,N_16208,N_16186);
and U24543 (N_24543,N_18547,N_19192);
and U24544 (N_24544,N_16331,N_12055);
nand U24545 (N_24545,N_16534,N_13775);
nand U24546 (N_24546,N_12388,N_18240);
and U24547 (N_24547,N_15284,N_16883);
and U24548 (N_24548,N_13824,N_10598);
nor U24549 (N_24549,N_12649,N_16350);
nand U24550 (N_24550,N_14343,N_14368);
or U24551 (N_24551,N_19407,N_11168);
and U24552 (N_24552,N_12688,N_14742);
nor U24553 (N_24553,N_18434,N_17725);
nand U24554 (N_24554,N_11620,N_18684);
xnor U24555 (N_24555,N_16488,N_13566);
nor U24556 (N_24556,N_15608,N_10648);
and U24557 (N_24557,N_10862,N_16827);
nand U24558 (N_24558,N_12018,N_19613);
xor U24559 (N_24559,N_11355,N_11951);
nor U24560 (N_24560,N_12653,N_18499);
or U24561 (N_24561,N_10777,N_17102);
xor U24562 (N_24562,N_18686,N_19071);
and U24563 (N_24563,N_14976,N_16946);
or U24564 (N_24564,N_16581,N_16067);
nand U24565 (N_24565,N_14404,N_10484);
or U24566 (N_24566,N_19450,N_11302);
nor U24567 (N_24567,N_12819,N_13412);
nor U24568 (N_24568,N_18119,N_14383);
or U24569 (N_24569,N_13743,N_15805);
or U24570 (N_24570,N_13789,N_19932);
nor U24571 (N_24571,N_15612,N_19839);
or U24572 (N_24572,N_14195,N_14775);
and U24573 (N_24573,N_12641,N_19396);
nand U24574 (N_24574,N_18701,N_11532);
and U24575 (N_24575,N_16130,N_18699);
or U24576 (N_24576,N_13816,N_19308);
nand U24577 (N_24577,N_15424,N_12182);
or U24578 (N_24578,N_13850,N_12171);
xnor U24579 (N_24579,N_19397,N_12118);
and U24580 (N_24580,N_18405,N_16207);
nor U24581 (N_24581,N_13380,N_15522);
or U24582 (N_24582,N_13563,N_18310);
or U24583 (N_24583,N_10189,N_11131);
xnor U24584 (N_24584,N_17916,N_13022);
or U24585 (N_24585,N_13313,N_11522);
or U24586 (N_24586,N_11437,N_10220);
and U24587 (N_24587,N_12933,N_16510);
and U24588 (N_24588,N_10649,N_11919);
and U24589 (N_24589,N_13198,N_16102);
nor U24590 (N_24590,N_10789,N_12689);
nor U24591 (N_24591,N_19523,N_12131);
nand U24592 (N_24592,N_19361,N_14108);
nand U24593 (N_24593,N_11516,N_16571);
nand U24594 (N_24594,N_15248,N_15675);
xor U24595 (N_24595,N_18452,N_17462);
and U24596 (N_24596,N_15737,N_15740);
and U24597 (N_24597,N_15715,N_13219);
nand U24598 (N_24598,N_12094,N_19829);
xnor U24599 (N_24599,N_11546,N_13517);
xor U24600 (N_24600,N_18408,N_11352);
nor U24601 (N_24601,N_11133,N_18471);
xor U24602 (N_24602,N_19271,N_12534);
nor U24603 (N_24603,N_11018,N_19408);
or U24604 (N_24604,N_19704,N_13735);
or U24605 (N_24605,N_12489,N_14116);
or U24606 (N_24606,N_13199,N_10359);
xor U24607 (N_24607,N_10935,N_11771);
or U24608 (N_24608,N_13696,N_17656);
or U24609 (N_24609,N_19168,N_12428);
and U24610 (N_24610,N_11207,N_12360);
nand U24611 (N_24611,N_18501,N_13070);
or U24612 (N_24612,N_18510,N_12352);
and U24613 (N_24613,N_15512,N_15591);
nand U24614 (N_24614,N_19256,N_11011);
xnor U24615 (N_24615,N_14017,N_10991);
nor U24616 (N_24616,N_16306,N_14020);
or U24617 (N_24617,N_15433,N_16095);
or U24618 (N_24618,N_10852,N_16596);
nand U24619 (N_24619,N_10338,N_12772);
or U24620 (N_24620,N_15239,N_14844);
nand U24621 (N_24621,N_19624,N_13117);
or U24622 (N_24622,N_15266,N_12444);
nor U24623 (N_24623,N_10354,N_13937);
nor U24624 (N_24624,N_18062,N_13255);
xnor U24625 (N_24625,N_10735,N_18120);
xor U24626 (N_24626,N_19994,N_14673);
nand U24627 (N_24627,N_17861,N_14652);
or U24628 (N_24628,N_11376,N_17904);
or U24629 (N_24629,N_17458,N_17573);
nand U24630 (N_24630,N_19772,N_18841);
and U24631 (N_24631,N_14147,N_13330);
xor U24632 (N_24632,N_19218,N_11397);
xnor U24633 (N_24633,N_17292,N_10745);
nand U24634 (N_24634,N_14337,N_13233);
and U24635 (N_24635,N_10066,N_14555);
xnor U24636 (N_24636,N_18949,N_17970);
xnor U24637 (N_24637,N_12916,N_11932);
and U24638 (N_24638,N_16082,N_15720);
and U24639 (N_24639,N_17812,N_14200);
xnor U24640 (N_24640,N_14275,N_14449);
or U24641 (N_24641,N_10363,N_15182);
xor U24642 (N_24642,N_15877,N_13408);
nor U24643 (N_24643,N_12117,N_19565);
nand U24644 (N_24644,N_13905,N_14554);
xnor U24645 (N_24645,N_17840,N_13301);
and U24646 (N_24646,N_13528,N_11922);
xnor U24647 (N_24647,N_14101,N_10448);
xnor U24648 (N_24648,N_16804,N_11314);
nor U24649 (N_24649,N_12232,N_19401);
and U24650 (N_24650,N_11461,N_17304);
xnor U24651 (N_24651,N_17753,N_12779);
nor U24652 (N_24652,N_15918,N_11482);
xnor U24653 (N_24653,N_10955,N_10048);
nor U24654 (N_24654,N_17315,N_18570);
nand U24655 (N_24655,N_11588,N_16389);
nor U24656 (N_24656,N_17938,N_16241);
xnor U24657 (N_24657,N_18306,N_12420);
xnor U24658 (N_24658,N_15807,N_13338);
and U24659 (N_24659,N_10791,N_14856);
nor U24660 (N_24660,N_13899,N_14166);
nand U24661 (N_24661,N_14901,N_17796);
xor U24662 (N_24662,N_14927,N_13350);
or U24663 (N_24663,N_13724,N_17638);
and U24664 (N_24664,N_15031,N_11150);
or U24665 (N_24665,N_16648,N_14508);
or U24666 (N_24666,N_13475,N_12615);
xnor U24667 (N_24667,N_15307,N_10869);
nand U24668 (N_24668,N_13184,N_15327);
nand U24669 (N_24669,N_14816,N_16057);
nor U24670 (N_24670,N_19236,N_17791);
nand U24671 (N_24671,N_18730,N_10244);
nor U24672 (N_24672,N_11816,N_13894);
nand U24673 (N_24673,N_14883,N_18608);
nor U24674 (N_24674,N_18944,N_16191);
nand U24675 (N_24675,N_10203,N_19412);
or U24676 (N_24676,N_11117,N_11815);
xor U24677 (N_24677,N_17465,N_11793);
xnor U24678 (N_24678,N_19746,N_18687);
nand U24679 (N_24679,N_12283,N_15118);
and U24680 (N_24680,N_19185,N_12505);
nand U24681 (N_24681,N_12486,N_13078);
and U24682 (N_24682,N_14685,N_11163);
nor U24683 (N_24683,N_13579,N_12159);
or U24684 (N_24684,N_10356,N_14629);
nand U24685 (N_24685,N_14420,N_11912);
xnor U24686 (N_24686,N_15769,N_13557);
nand U24687 (N_24687,N_15562,N_18046);
nand U24688 (N_24688,N_11759,N_11056);
or U24689 (N_24689,N_17183,N_17194);
or U24690 (N_24690,N_18259,N_19677);
and U24691 (N_24691,N_16319,N_18371);
nand U24692 (N_24692,N_11548,N_14141);
xor U24693 (N_24693,N_13142,N_13819);
xnor U24694 (N_24694,N_13298,N_14795);
nor U24695 (N_24695,N_10931,N_15864);
xnor U24696 (N_24696,N_17620,N_16907);
xor U24697 (N_24697,N_10737,N_15772);
or U24698 (N_24698,N_16625,N_15115);
and U24699 (N_24699,N_12713,N_11628);
xnor U24700 (N_24700,N_14370,N_11872);
xnor U24701 (N_24701,N_17095,N_17267);
and U24702 (N_24702,N_12262,N_19209);
xor U24703 (N_24703,N_16684,N_16744);
nand U24704 (N_24704,N_16139,N_10384);
nand U24705 (N_24705,N_10532,N_18073);
or U24706 (N_24706,N_17310,N_15290);
xor U24707 (N_24707,N_18299,N_14890);
nand U24708 (N_24708,N_14509,N_18418);
and U24709 (N_24709,N_13329,N_19609);
and U24710 (N_24710,N_17589,N_14448);
or U24711 (N_24711,N_10661,N_13170);
nor U24712 (N_24712,N_19841,N_11299);
and U24713 (N_24713,N_12766,N_15988);
nor U24714 (N_24714,N_19672,N_17721);
nand U24715 (N_24715,N_14644,N_16685);
or U24716 (N_24716,N_19026,N_10482);
nor U24717 (N_24717,N_14133,N_15212);
xnor U24718 (N_24718,N_17775,N_14354);
and U24719 (N_24719,N_17643,N_11787);
or U24720 (N_24720,N_13195,N_18670);
and U24721 (N_24721,N_17234,N_16489);
and U24722 (N_24722,N_19423,N_15356);
xor U24723 (N_24723,N_18693,N_11265);
xor U24724 (N_24724,N_17675,N_16193);
xnor U24725 (N_24725,N_17953,N_12201);
and U24726 (N_24726,N_18773,N_18597);
xor U24727 (N_24727,N_11717,N_17262);
or U24728 (N_24728,N_15302,N_17509);
nor U24729 (N_24729,N_19741,N_18566);
and U24730 (N_24730,N_10426,N_15282);
xnor U24731 (N_24731,N_16784,N_15680);
nand U24732 (N_24732,N_12522,N_17341);
nor U24733 (N_24733,N_18416,N_13083);
or U24734 (N_24734,N_11675,N_13919);
and U24735 (N_24735,N_19583,N_15962);
nor U24736 (N_24736,N_14952,N_16436);
and U24737 (N_24737,N_16252,N_12338);
nand U24738 (N_24738,N_19464,N_11496);
nor U24739 (N_24739,N_14205,N_15644);
and U24740 (N_24740,N_10796,N_14322);
nand U24741 (N_24741,N_11450,N_15974);
xnor U24742 (N_24742,N_12627,N_18900);
xor U24743 (N_24743,N_10516,N_10152);
nand U24744 (N_24744,N_10952,N_19955);
nand U24745 (N_24745,N_14164,N_16745);
nor U24746 (N_24746,N_12864,N_13609);
and U24747 (N_24747,N_15273,N_13872);
xor U24748 (N_24748,N_13459,N_14671);
or U24749 (N_24749,N_19773,N_12364);
xnor U24750 (N_24750,N_10809,N_10872);
nand U24751 (N_24751,N_14137,N_10392);
nor U24752 (N_24752,N_12651,N_16657);
nor U24753 (N_24753,N_14790,N_12016);
or U24754 (N_24754,N_12017,N_14912);
nand U24755 (N_24755,N_18116,N_11699);
or U24756 (N_24756,N_18254,N_16030);
or U24757 (N_24757,N_14854,N_10879);
or U24758 (N_24758,N_16921,N_16756);
or U24759 (N_24759,N_11557,N_19604);
and U24760 (N_24760,N_12080,N_19486);
xor U24761 (N_24761,N_12501,N_19850);
nor U24762 (N_24762,N_13959,N_19368);
or U24763 (N_24763,N_15265,N_19353);
nand U24764 (N_24764,N_13060,N_11113);
xnor U24765 (N_24765,N_19166,N_16460);
xnor U24766 (N_24766,N_13288,N_14853);
nand U24767 (N_24767,N_10027,N_12549);
nor U24768 (N_24768,N_12994,N_17544);
xnor U24769 (N_24769,N_13357,N_11523);
nor U24770 (N_24770,N_19787,N_11764);
and U24771 (N_24771,N_15831,N_12938);
and U24772 (N_24772,N_13419,N_15369);
xor U24773 (N_24773,N_14289,N_18780);
xnor U24774 (N_24774,N_16805,N_15760);
nand U24775 (N_24775,N_13849,N_16959);
and U24776 (N_24776,N_19823,N_12672);
nand U24777 (N_24777,N_18297,N_18709);
xnor U24778 (N_24778,N_19531,N_15797);
nand U24779 (N_24779,N_18159,N_19909);
or U24780 (N_24780,N_18839,N_19903);
or U24781 (N_24781,N_19750,N_13857);
and U24782 (N_24782,N_18318,N_14489);
xor U24783 (N_24783,N_18357,N_14262);
nor U24784 (N_24784,N_12231,N_15026);
nand U24785 (N_24785,N_11097,N_19036);
nand U24786 (N_24786,N_19008,N_12927);
nor U24787 (N_24787,N_15753,N_16983);
nand U24788 (N_24788,N_17378,N_10023);
nor U24789 (N_24789,N_15459,N_14627);
or U24790 (N_24790,N_17865,N_16199);
nor U24791 (N_24791,N_10619,N_12060);
nand U24792 (N_24792,N_19558,N_16101);
nor U24793 (N_24793,N_17524,N_18809);
xor U24794 (N_24794,N_10888,N_10361);
or U24795 (N_24795,N_17374,N_14457);
nor U24796 (N_24796,N_19180,N_18131);
and U24797 (N_24797,N_17636,N_13227);
nand U24798 (N_24798,N_15315,N_17269);
and U24799 (N_24799,N_17157,N_19421);
nand U24800 (N_24800,N_10110,N_18112);
nand U24801 (N_24801,N_12453,N_14481);
or U24802 (N_24802,N_15689,N_14967);
or U24803 (N_24803,N_15735,N_13716);
nand U24804 (N_24804,N_15845,N_12156);
nor U24805 (N_24805,N_19817,N_12708);
nor U24806 (N_24806,N_15196,N_18692);
nand U24807 (N_24807,N_10781,N_19365);
and U24808 (N_24808,N_18794,N_12612);
nor U24809 (N_24809,N_17264,N_14237);
nor U24810 (N_24810,N_12635,N_19324);
or U24811 (N_24811,N_16792,N_17290);
nor U24812 (N_24812,N_19647,N_10953);
xnor U24813 (N_24813,N_14608,N_14432);
nand U24814 (N_24814,N_12874,N_10933);
nor U24815 (N_24815,N_11140,N_18911);
nand U24816 (N_24816,N_12253,N_13042);
and U24817 (N_24817,N_19402,N_14948);
and U24818 (N_24818,N_11563,N_15700);
xnor U24819 (N_24819,N_16311,N_10415);
and U24820 (N_24820,N_15247,N_12701);
or U24821 (N_24821,N_19599,N_16908);
xor U24822 (N_24822,N_17498,N_12690);
and U24823 (N_24823,N_13832,N_16142);
and U24824 (N_24824,N_15142,N_19812);
and U24825 (N_24825,N_10570,N_12108);
and U24826 (N_24826,N_19445,N_15069);
xnor U24827 (N_24827,N_15932,N_15563);
nand U24828 (N_24828,N_13193,N_13900);
nand U24829 (N_24829,N_16062,N_19461);
xor U24830 (N_24830,N_12178,N_19685);
and U24831 (N_24831,N_11559,N_18927);
nand U24832 (N_24832,N_11088,N_16773);
nand U24833 (N_24833,N_13728,N_15548);
and U24834 (N_24834,N_11892,N_13468);
and U24835 (N_24835,N_11533,N_11470);
nor U24836 (N_24836,N_16803,N_15259);
nand U24837 (N_24837,N_17969,N_10131);
xor U24838 (N_24838,N_15815,N_13545);
nand U24839 (N_24839,N_17169,N_15773);
or U24840 (N_24840,N_10873,N_17333);
or U24841 (N_24841,N_15993,N_11183);
or U24842 (N_24842,N_14333,N_15197);
nor U24843 (N_24843,N_19722,N_16000);
nor U24844 (N_24844,N_12821,N_16935);
and U24845 (N_24845,N_13519,N_17908);
xnor U24846 (N_24846,N_12276,N_19490);
or U24847 (N_24847,N_17797,N_16381);
nor U24848 (N_24848,N_16894,N_19351);
nand U24849 (N_24849,N_18361,N_13632);
and U24850 (N_24850,N_18792,N_14339);
and U24851 (N_24851,N_11575,N_17155);
nor U24852 (N_24852,N_17568,N_15820);
nor U24853 (N_24853,N_13238,N_16498);
nor U24854 (N_24854,N_17099,N_18255);
or U24855 (N_24855,N_10678,N_12087);
xor U24856 (N_24856,N_15233,N_12446);
xor U24857 (N_24857,N_15850,N_13179);
and U24858 (N_24858,N_18758,N_19499);
or U24859 (N_24859,N_13356,N_19013);
nand U24860 (N_24860,N_17995,N_15213);
nand U24861 (N_24861,N_11130,N_18812);
nand U24862 (N_24862,N_11911,N_11978);
xnor U24863 (N_24863,N_10332,N_11255);
and U24864 (N_24864,N_11473,N_14384);
nor U24865 (N_24865,N_18463,N_13074);
nor U24866 (N_24866,N_19581,N_11017);
nor U24867 (N_24867,N_15856,N_17739);
nor U24868 (N_24868,N_11972,N_13845);
xor U24869 (N_24869,N_16269,N_11342);
and U24870 (N_24870,N_12057,N_15386);
xnor U24871 (N_24871,N_19020,N_19060);
or U24872 (N_24872,N_15280,N_18513);
nor U24873 (N_24873,N_14916,N_15621);
xnor U24874 (N_24874,N_14417,N_11334);
nor U24875 (N_24875,N_12236,N_17516);
nor U24876 (N_24876,N_15472,N_10847);
xnor U24877 (N_24877,N_19803,N_18420);
and U24878 (N_24878,N_15022,N_13121);
and U24879 (N_24879,N_13456,N_19539);
xor U24880 (N_24880,N_12429,N_19743);
or U24881 (N_24881,N_18760,N_18061);
xnor U24882 (N_24882,N_14889,N_12220);
nor U24883 (N_24883,N_15987,N_18690);
nor U24884 (N_24884,N_19319,N_17810);
xor U24885 (N_24885,N_13189,N_12763);
and U24886 (N_24886,N_15322,N_15844);
or U24887 (N_24887,N_15095,N_13292);
xnor U24888 (N_24888,N_18641,N_12660);
nor U24889 (N_24889,N_11692,N_16343);
and U24890 (N_24890,N_14330,N_16743);
nor U24891 (N_24891,N_15272,N_13807);
nor U24892 (N_24892,N_15323,N_17975);
nand U24893 (N_24893,N_17398,N_11773);
and U24894 (N_24894,N_11530,N_18766);
and U24895 (N_24895,N_17176,N_19109);
nor U24896 (N_24896,N_17349,N_11167);
and U24897 (N_24897,N_19846,N_12890);
xnor U24898 (N_24898,N_17459,N_10468);
nand U24899 (N_24899,N_15311,N_17960);
or U24900 (N_24900,N_10645,N_13509);
xnor U24901 (N_24901,N_14230,N_13144);
nand U24902 (N_24902,N_13598,N_12868);
nor U24903 (N_24903,N_16111,N_13071);
xnor U24904 (N_24904,N_16388,N_17629);
xnor U24905 (N_24905,N_12246,N_16108);
and U24906 (N_24906,N_13369,N_18847);
or U24907 (N_24907,N_18607,N_13931);
nor U24908 (N_24908,N_10488,N_17495);
or U24909 (N_24909,N_13548,N_12351);
nor U24910 (N_24910,N_18172,N_17190);
or U24911 (N_24911,N_16518,N_17428);
nor U24912 (N_24912,N_15172,N_17581);
nand U24913 (N_24913,N_13759,N_17917);
or U24914 (N_24914,N_11649,N_12030);
xor U24915 (N_24915,N_13644,N_11896);
nand U24916 (N_24916,N_13511,N_17389);
or U24917 (N_24917,N_16429,N_14603);
nor U24918 (N_24918,N_10685,N_13799);
nor U24919 (N_24919,N_15104,N_15226);
xor U24920 (N_24920,N_17177,N_15791);
nand U24921 (N_24921,N_19779,N_16063);
nand U24922 (N_24922,N_12878,N_11318);
and U24923 (N_24923,N_17628,N_16884);
xor U24924 (N_24924,N_18058,N_10890);
and U24925 (N_24925,N_17868,N_13893);
nor U24926 (N_24926,N_17119,N_18702);
or U24927 (N_24927,N_16019,N_16454);
or U24928 (N_24928,N_16870,N_18904);
or U24929 (N_24929,N_19057,N_18864);
nor U24930 (N_24930,N_15251,N_16113);
nor U24931 (N_24931,N_12059,N_10014);
nor U24932 (N_24932,N_14250,N_10740);
and U24933 (N_24933,N_19682,N_10727);
or U24934 (N_24934,N_15238,N_10227);
or U24935 (N_24935,N_16106,N_11244);
nand U24936 (N_24936,N_17558,N_18808);
and U24937 (N_24937,N_18672,N_10541);
and U24938 (N_24938,N_13878,N_11737);
and U24939 (N_24939,N_10469,N_14198);
or U24940 (N_24940,N_13112,N_18910);
xor U24941 (N_24941,N_15597,N_19086);
nor U24942 (N_24942,N_16329,N_15217);
nand U24943 (N_24943,N_12036,N_10824);
or U24944 (N_24944,N_16733,N_13810);
or U24945 (N_24945,N_18018,N_10223);
or U24946 (N_24946,N_15420,N_16913);
and U24947 (N_24947,N_16865,N_13987);
xnor U24948 (N_24948,N_10814,N_10732);
xor U24949 (N_24949,N_16876,N_11538);
nand U24950 (N_24950,N_16896,N_13951);
nor U24951 (N_24951,N_12716,N_16076);
or U24952 (N_24952,N_12770,N_18319);
xnor U24953 (N_24953,N_17873,N_18307);
and U24954 (N_24954,N_19241,N_16877);
nor U24955 (N_24955,N_14212,N_11803);
nand U24956 (N_24956,N_15450,N_16726);
nand U24957 (N_24957,N_17139,N_15939);
or U24958 (N_24958,N_19659,N_16891);
xor U24959 (N_24959,N_16903,N_19110);
nand U24960 (N_24960,N_18004,N_15682);
or U24961 (N_24961,N_15303,N_10752);
and U24962 (N_24962,N_17401,N_13496);
or U24963 (N_24963,N_16356,N_15360);
nor U24964 (N_24964,N_12362,N_14761);
and U24965 (N_24965,N_16893,N_19938);
nand U24966 (N_24966,N_19838,N_12941);
nand U24967 (N_24967,N_18379,N_16040);
and U24968 (N_24968,N_11317,N_13904);
nand U24969 (N_24969,N_12562,N_11615);
or U24970 (N_24970,N_19064,N_15891);
nand U24971 (N_24971,N_12969,N_15903);
and U24972 (N_24972,N_10907,N_10628);
xnor U24973 (N_24973,N_11321,N_19883);
or U24974 (N_24974,N_16914,N_11738);
or U24975 (N_24975,N_18270,N_19432);
or U24976 (N_24976,N_18536,N_18551);
nor U24977 (N_24977,N_16222,N_12328);
and U24978 (N_24978,N_16725,N_14081);
and U24979 (N_24979,N_19058,N_11934);
nand U24980 (N_24980,N_18069,N_12124);
xnor U24981 (N_24981,N_15440,N_18382);
or U24982 (N_24982,N_11735,N_16826);
and U24983 (N_24983,N_16005,N_17143);
xor U24984 (N_24984,N_15677,N_13470);
nor U24985 (N_24985,N_15283,N_19237);
nand U24986 (N_24986,N_17742,N_19908);
nand U24987 (N_24987,N_15350,N_10262);
nor U24988 (N_24988,N_11125,N_13671);
xnor U24989 (N_24989,N_11642,N_16623);
nor U24990 (N_24990,N_14771,N_11585);
and U24991 (N_24991,N_16401,N_16618);
and U24992 (N_24992,N_18278,N_11790);
and U24993 (N_24993,N_13399,N_16722);
nor U24994 (N_24994,N_16868,N_10827);
or U24995 (N_24995,N_13201,N_14776);
nor U24996 (N_24996,N_15566,N_15324);
xnor U24997 (N_24997,N_19840,N_10504);
nor U24998 (N_24998,N_12041,N_11613);
or U24999 (N_24999,N_12965,N_10381);
xor U25000 (N_25000,N_15272,N_17105);
xnor U25001 (N_25001,N_15979,N_12419);
and U25002 (N_25002,N_19313,N_13321);
nor U25003 (N_25003,N_16886,N_11784);
or U25004 (N_25004,N_18806,N_17246);
nand U25005 (N_25005,N_17632,N_15459);
nand U25006 (N_25006,N_13991,N_12302);
nor U25007 (N_25007,N_11979,N_19372);
nand U25008 (N_25008,N_18890,N_12855);
nor U25009 (N_25009,N_15653,N_17702);
or U25010 (N_25010,N_12960,N_11160);
nor U25011 (N_25011,N_10855,N_18688);
or U25012 (N_25012,N_11740,N_10394);
xor U25013 (N_25013,N_11810,N_13560);
nand U25014 (N_25014,N_16976,N_17478);
xnor U25015 (N_25015,N_15199,N_10555);
xnor U25016 (N_25016,N_11140,N_15740);
nor U25017 (N_25017,N_19313,N_13943);
or U25018 (N_25018,N_16168,N_12102);
or U25019 (N_25019,N_15178,N_10682);
or U25020 (N_25020,N_13007,N_16795);
or U25021 (N_25021,N_17872,N_18141);
or U25022 (N_25022,N_16228,N_17167);
or U25023 (N_25023,N_12059,N_11543);
xnor U25024 (N_25024,N_19739,N_14611);
xor U25025 (N_25025,N_17530,N_10010);
nand U25026 (N_25026,N_16717,N_13794);
and U25027 (N_25027,N_11465,N_18504);
or U25028 (N_25028,N_19174,N_19606);
nor U25029 (N_25029,N_14487,N_10054);
nor U25030 (N_25030,N_19607,N_11857);
or U25031 (N_25031,N_10679,N_14633);
xor U25032 (N_25032,N_14503,N_18986);
or U25033 (N_25033,N_12004,N_17360);
and U25034 (N_25034,N_14819,N_19859);
and U25035 (N_25035,N_12540,N_15773);
or U25036 (N_25036,N_13194,N_13891);
nand U25037 (N_25037,N_14896,N_11620);
xnor U25038 (N_25038,N_12025,N_14731);
and U25039 (N_25039,N_12473,N_13589);
xnor U25040 (N_25040,N_19485,N_12001);
and U25041 (N_25041,N_19021,N_18109);
nor U25042 (N_25042,N_10903,N_14071);
nor U25043 (N_25043,N_11223,N_10072);
and U25044 (N_25044,N_15114,N_13447);
and U25045 (N_25045,N_12527,N_13066);
and U25046 (N_25046,N_18474,N_12101);
xnor U25047 (N_25047,N_16926,N_14811);
nor U25048 (N_25048,N_14643,N_14542);
xnor U25049 (N_25049,N_13512,N_12584);
nor U25050 (N_25050,N_13182,N_19049);
nand U25051 (N_25051,N_13700,N_18676);
xnor U25052 (N_25052,N_11428,N_17342);
nand U25053 (N_25053,N_18349,N_15172);
nor U25054 (N_25054,N_10246,N_13647);
or U25055 (N_25055,N_13573,N_10458);
nand U25056 (N_25056,N_19558,N_11172);
nand U25057 (N_25057,N_15068,N_11009);
and U25058 (N_25058,N_10136,N_17769);
xor U25059 (N_25059,N_16701,N_13084);
nor U25060 (N_25060,N_17906,N_13779);
nor U25061 (N_25061,N_17296,N_17006);
nor U25062 (N_25062,N_13489,N_15019);
and U25063 (N_25063,N_11889,N_12882);
nor U25064 (N_25064,N_11462,N_11660);
and U25065 (N_25065,N_15083,N_11032);
and U25066 (N_25066,N_12847,N_15058);
or U25067 (N_25067,N_17663,N_12363);
and U25068 (N_25068,N_13954,N_17093);
or U25069 (N_25069,N_10228,N_12853);
nor U25070 (N_25070,N_13664,N_13052);
xnor U25071 (N_25071,N_10415,N_17427);
or U25072 (N_25072,N_15362,N_18882);
or U25073 (N_25073,N_15707,N_17041);
or U25074 (N_25074,N_13742,N_18426);
nor U25075 (N_25075,N_18113,N_10709);
nand U25076 (N_25076,N_17021,N_17357);
or U25077 (N_25077,N_18761,N_16655);
nor U25078 (N_25078,N_14083,N_17882);
and U25079 (N_25079,N_16337,N_13873);
and U25080 (N_25080,N_13439,N_17690);
and U25081 (N_25081,N_17266,N_15293);
nor U25082 (N_25082,N_16980,N_11846);
nand U25083 (N_25083,N_17161,N_19415);
xnor U25084 (N_25084,N_14340,N_14151);
nand U25085 (N_25085,N_16815,N_19289);
nand U25086 (N_25086,N_16035,N_10037);
nor U25087 (N_25087,N_19515,N_15233);
nor U25088 (N_25088,N_13948,N_19583);
nand U25089 (N_25089,N_17025,N_17005);
nor U25090 (N_25090,N_15653,N_16636);
or U25091 (N_25091,N_13734,N_18297);
or U25092 (N_25092,N_13189,N_14103);
nand U25093 (N_25093,N_17287,N_15412);
nand U25094 (N_25094,N_16675,N_10006);
and U25095 (N_25095,N_13542,N_15076);
nand U25096 (N_25096,N_10541,N_16933);
and U25097 (N_25097,N_11774,N_11980);
or U25098 (N_25098,N_13998,N_14165);
nand U25099 (N_25099,N_18599,N_19829);
nand U25100 (N_25100,N_16149,N_17979);
and U25101 (N_25101,N_11707,N_15907);
and U25102 (N_25102,N_16708,N_12061);
nand U25103 (N_25103,N_15368,N_15246);
or U25104 (N_25104,N_10622,N_13041);
nand U25105 (N_25105,N_10822,N_11495);
nand U25106 (N_25106,N_12207,N_11069);
nand U25107 (N_25107,N_13828,N_18056);
xnor U25108 (N_25108,N_14615,N_19291);
and U25109 (N_25109,N_15042,N_18173);
nand U25110 (N_25110,N_15062,N_18543);
xnor U25111 (N_25111,N_11742,N_10731);
or U25112 (N_25112,N_14782,N_13904);
nor U25113 (N_25113,N_17268,N_12135);
xnor U25114 (N_25114,N_10714,N_10300);
nand U25115 (N_25115,N_10060,N_17474);
or U25116 (N_25116,N_11801,N_12639);
and U25117 (N_25117,N_14564,N_15084);
xnor U25118 (N_25118,N_12329,N_16579);
nand U25119 (N_25119,N_10479,N_15434);
xnor U25120 (N_25120,N_19623,N_18042);
nand U25121 (N_25121,N_13029,N_15542);
nor U25122 (N_25122,N_13256,N_11746);
xnor U25123 (N_25123,N_18816,N_12086);
nand U25124 (N_25124,N_11270,N_14096);
xor U25125 (N_25125,N_12254,N_19149);
or U25126 (N_25126,N_13299,N_13121);
or U25127 (N_25127,N_11251,N_10511);
xor U25128 (N_25128,N_12190,N_16752);
nand U25129 (N_25129,N_19330,N_12972);
xnor U25130 (N_25130,N_14877,N_19198);
nor U25131 (N_25131,N_13053,N_12668);
nand U25132 (N_25132,N_10638,N_14971);
nor U25133 (N_25133,N_18364,N_10577);
nand U25134 (N_25134,N_13729,N_16621);
xor U25135 (N_25135,N_15111,N_11573);
nand U25136 (N_25136,N_18430,N_16192);
nor U25137 (N_25137,N_14074,N_17676);
or U25138 (N_25138,N_13441,N_18729);
nand U25139 (N_25139,N_15995,N_16102);
nor U25140 (N_25140,N_12774,N_11044);
nand U25141 (N_25141,N_11266,N_14424);
or U25142 (N_25142,N_17968,N_19833);
xor U25143 (N_25143,N_15997,N_16140);
nor U25144 (N_25144,N_16572,N_14467);
nand U25145 (N_25145,N_18469,N_18823);
or U25146 (N_25146,N_18708,N_19802);
or U25147 (N_25147,N_10575,N_18879);
xor U25148 (N_25148,N_14517,N_13031);
nand U25149 (N_25149,N_14951,N_17449);
xnor U25150 (N_25150,N_13722,N_10655);
xnor U25151 (N_25151,N_10860,N_12717);
xor U25152 (N_25152,N_16360,N_19923);
or U25153 (N_25153,N_17667,N_14402);
and U25154 (N_25154,N_18843,N_10215);
or U25155 (N_25155,N_10433,N_14213);
or U25156 (N_25156,N_13513,N_19558);
xnor U25157 (N_25157,N_16415,N_12656);
nor U25158 (N_25158,N_19905,N_17770);
or U25159 (N_25159,N_14265,N_11896);
or U25160 (N_25160,N_18083,N_17822);
and U25161 (N_25161,N_19177,N_13169);
nor U25162 (N_25162,N_11166,N_15005);
nor U25163 (N_25163,N_18433,N_10560);
nor U25164 (N_25164,N_13232,N_17823);
or U25165 (N_25165,N_10461,N_10504);
and U25166 (N_25166,N_16231,N_12376);
nand U25167 (N_25167,N_17053,N_13377);
xor U25168 (N_25168,N_11280,N_12774);
nor U25169 (N_25169,N_15313,N_12213);
xnor U25170 (N_25170,N_16915,N_12677);
or U25171 (N_25171,N_12668,N_15772);
and U25172 (N_25172,N_10617,N_10412);
and U25173 (N_25173,N_13156,N_16239);
or U25174 (N_25174,N_13942,N_16489);
and U25175 (N_25175,N_17605,N_19577);
nor U25176 (N_25176,N_10741,N_16869);
and U25177 (N_25177,N_18231,N_14004);
nand U25178 (N_25178,N_19722,N_12130);
xor U25179 (N_25179,N_10807,N_19186);
and U25180 (N_25180,N_13249,N_19904);
or U25181 (N_25181,N_16921,N_15516);
or U25182 (N_25182,N_11829,N_10019);
or U25183 (N_25183,N_17030,N_18601);
nand U25184 (N_25184,N_15653,N_11689);
and U25185 (N_25185,N_15217,N_16730);
and U25186 (N_25186,N_17524,N_15224);
and U25187 (N_25187,N_12244,N_14547);
xnor U25188 (N_25188,N_19120,N_19882);
and U25189 (N_25189,N_14064,N_10896);
nor U25190 (N_25190,N_13290,N_15966);
and U25191 (N_25191,N_11826,N_13245);
or U25192 (N_25192,N_15406,N_19441);
xor U25193 (N_25193,N_12266,N_12006);
nor U25194 (N_25194,N_15582,N_14414);
nand U25195 (N_25195,N_11446,N_14214);
nor U25196 (N_25196,N_15889,N_19744);
or U25197 (N_25197,N_14401,N_13449);
nor U25198 (N_25198,N_13359,N_11214);
and U25199 (N_25199,N_16341,N_13832);
nor U25200 (N_25200,N_18394,N_19020);
nor U25201 (N_25201,N_13616,N_18332);
nand U25202 (N_25202,N_13510,N_12072);
or U25203 (N_25203,N_19720,N_11037);
nand U25204 (N_25204,N_14876,N_14655);
nor U25205 (N_25205,N_13878,N_19258);
nor U25206 (N_25206,N_10781,N_17208);
or U25207 (N_25207,N_19688,N_17153);
and U25208 (N_25208,N_16390,N_15054);
nand U25209 (N_25209,N_19570,N_17952);
or U25210 (N_25210,N_13860,N_16792);
nand U25211 (N_25211,N_19645,N_15601);
nor U25212 (N_25212,N_16120,N_17196);
and U25213 (N_25213,N_16588,N_13354);
xor U25214 (N_25214,N_15065,N_10345);
and U25215 (N_25215,N_18098,N_12530);
nand U25216 (N_25216,N_18761,N_11195);
and U25217 (N_25217,N_11794,N_15392);
nor U25218 (N_25218,N_19203,N_18503);
and U25219 (N_25219,N_13269,N_14785);
and U25220 (N_25220,N_13840,N_19050);
nand U25221 (N_25221,N_16192,N_15908);
nor U25222 (N_25222,N_18938,N_13431);
or U25223 (N_25223,N_14620,N_13616);
and U25224 (N_25224,N_12587,N_15121);
or U25225 (N_25225,N_13286,N_13315);
xor U25226 (N_25226,N_18216,N_19387);
and U25227 (N_25227,N_11756,N_17505);
xor U25228 (N_25228,N_15096,N_12189);
or U25229 (N_25229,N_16284,N_10304);
and U25230 (N_25230,N_16159,N_17377);
xor U25231 (N_25231,N_13431,N_13542);
and U25232 (N_25232,N_13662,N_15869);
and U25233 (N_25233,N_11400,N_15608);
xor U25234 (N_25234,N_19134,N_11659);
and U25235 (N_25235,N_10947,N_17221);
nor U25236 (N_25236,N_10407,N_16984);
nor U25237 (N_25237,N_18848,N_18055);
nor U25238 (N_25238,N_10767,N_13542);
xnor U25239 (N_25239,N_14638,N_10655);
nor U25240 (N_25240,N_19699,N_12125);
and U25241 (N_25241,N_15857,N_17087);
or U25242 (N_25242,N_10339,N_12811);
or U25243 (N_25243,N_12767,N_12393);
or U25244 (N_25244,N_13146,N_19601);
and U25245 (N_25245,N_10994,N_11212);
nor U25246 (N_25246,N_15531,N_14133);
nor U25247 (N_25247,N_11718,N_11125);
nor U25248 (N_25248,N_15591,N_13519);
xor U25249 (N_25249,N_10432,N_18489);
nand U25250 (N_25250,N_15779,N_19421);
nor U25251 (N_25251,N_19287,N_18980);
and U25252 (N_25252,N_16758,N_14758);
nand U25253 (N_25253,N_10546,N_19901);
xnor U25254 (N_25254,N_19842,N_16402);
nor U25255 (N_25255,N_14849,N_14299);
or U25256 (N_25256,N_13025,N_17058);
nor U25257 (N_25257,N_12119,N_19053);
xor U25258 (N_25258,N_17373,N_16140);
xnor U25259 (N_25259,N_12047,N_10959);
nand U25260 (N_25260,N_17230,N_12472);
nand U25261 (N_25261,N_13206,N_19489);
nand U25262 (N_25262,N_12785,N_12310);
nand U25263 (N_25263,N_10799,N_17048);
and U25264 (N_25264,N_16243,N_10985);
and U25265 (N_25265,N_10695,N_13719);
nor U25266 (N_25266,N_19594,N_12572);
or U25267 (N_25267,N_11071,N_10482);
xnor U25268 (N_25268,N_11900,N_18101);
or U25269 (N_25269,N_17236,N_12237);
xor U25270 (N_25270,N_10658,N_10776);
nand U25271 (N_25271,N_13093,N_15308);
or U25272 (N_25272,N_10073,N_10737);
xor U25273 (N_25273,N_16419,N_16187);
nand U25274 (N_25274,N_14199,N_13747);
nand U25275 (N_25275,N_13812,N_19109);
xnor U25276 (N_25276,N_11984,N_12657);
or U25277 (N_25277,N_15825,N_13082);
and U25278 (N_25278,N_13342,N_13518);
or U25279 (N_25279,N_17648,N_12870);
nor U25280 (N_25280,N_14571,N_15020);
nor U25281 (N_25281,N_16614,N_11620);
and U25282 (N_25282,N_11710,N_19143);
or U25283 (N_25283,N_18823,N_18433);
nor U25284 (N_25284,N_15449,N_15105);
and U25285 (N_25285,N_10327,N_19772);
or U25286 (N_25286,N_16682,N_13309);
and U25287 (N_25287,N_19237,N_13424);
nand U25288 (N_25288,N_18337,N_16885);
or U25289 (N_25289,N_13701,N_10472);
xor U25290 (N_25290,N_13108,N_19547);
nand U25291 (N_25291,N_12334,N_15719);
xnor U25292 (N_25292,N_12477,N_19895);
nand U25293 (N_25293,N_11678,N_16213);
nor U25294 (N_25294,N_12376,N_18151);
xor U25295 (N_25295,N_10963,N_19392);
nand U25296 (N_25296,N_19746,N_17659);
nand U25297 (N_25297,N_15506,N_15883);
xnor U25298 (N_25298,N_18974,N_12986);
nor U25299 (N_25299,N_10386,N_10837);
xor U25300 (N_25300,N_19600,N_17115);
nor U25301 (N_25301,N_19081,N_10164);
xnor U25302 (N_25302,N_15298,N_18589);
and U25303 (N_25303,N_17259,N_14211);
and U25304 (N_25304,N_10229,N_13092);
nand U25305 (N_25305,N_18738,N_12933);
or U25306 (N_25306,N_11151,N_19004);
nor U25307 (N_25307,N_18012,N_17692);
and U25308 (N_25308,N_15207,N_10888);
or U25309 (N_25309,N_11867,N_13125);
nor U25310 (N_25310,N_15008,N_13690);
nand U25311 (N_25311,N_18983,N_16546);
or U25312 (N_25312,N_16167,N_18938);
nand U25313 (N_25313,N_16930,N_12678);
and U25314 (N_25314,N_19285,N_16961);
nor U25315 (N_25315,N_10726,N_12490);
or U25316 (N_25316,N_18410,N_16034);
nand U25317 (N_25317,N_12707,N_12398);
or U25318 (N_25318,N_16640,N_18852);
and U25319 (N_25319,N_12914,N_17886);
nor U25320 (N_25320,N_14257,N_12058);
nand U25321 (N_25321,N_10533,N_18938);
or U25322 (N_25322,N_17775,N_12324);
and U25323 (N_25323,N_10956,N_13790);
and U25324 (N_25324,N_19598,N_18447);
nor U25325 (N_25325,N_16389,N_18151);
or U25326 (N_25326,N_11503,N_11259);
xor U25327 (N_25327,N_10686,N_12851);
nand U25328 (N_25328,N_17434,N_18353);
nand U25329 (N_25329,N_10224,N_12111);
nor U25330 (N_25330,N_13439,N_11987);
nand U25331 (N_25331,N_19001,N_18025);
nor U25332 (N_25332,N_16734,N_12685);
xnor U25333 (N_25333,N_16335,N_12021);
or U25334 (N_25334,N_19169,N_12933);
nand U25335 (N_25335,N_14609,N_11145);
xor U25336 (N_25336,N_19497,N_12575);
or U25337 (N_25337,N_10448,N_16932);
or U25338 (N_25338,N_17056,N_10245);
or U25339 (N_25339,N_12489,N_11334);
and U25340 (N_25340,N_18953,N_11945);
nand U25341 (N_25341,N_11480,N_16170);
nand U25342 (N_25342,N_17205,N_16621);
nor U25343 (N_25343,N_16076,N_18080);
and U25344 (N_25344,N_13047,N_15152);
and U25345 (N_25345,N_11835,N_12211);
nor U25346 (N_25346,N_16724,N_19510);
or U25347 (N_25347,N_17808,N_15640);
and U25348 (N_25348,N_12117,N_12756);
or U25349 (N_25349,N_16794,N_13886);
nand U25350 (N_25350,N_13506,N_12422);
xor U25351 (N_25351,N_10128,N_14177);
or U25352 (N_25352,N_17340,N_15449);
nor U25353 (N_25353,N_14072,N_19466);
and U25354 (N_25354,N_19456,N_15258);
xnor U25355 (N_25355,N_14879,N_16042);
or U25356 (N_25356,N_13783,N_19175);
and U25357 (N_25357,N_18076,N_10299);
xor U25358 (N_25358,N_10508,N_16903);
xnor U25359 (N_25359,N_12662,N_17262);
nor U25360 (N_25360,N_17668,N_12589);
xor U25361 (N_25361,N_18499,N_11516);
nand U25362 (N_25362,N_15085,N_11884);
xor U25363 (N_25363,N_16616,N_14904);
and U25364 (N_25364,N_15351,N_10071);
or U25365 (N_25365,N_14783,N_18343);
and U25366 (N_25366,N_13646,N_14876);
nand U25367 (N_25367,N_12741,N_17266);
and U25368 (N_25368,N_10107,N_17772);
and U25369 (N_25369,N_17129,N_18616);
nor U25370 (N_25370,N_17611,N_13058);
nor U25371 (N_25371,N_11938,N_19815);
or U25372 (N_25372,N_11490,N_15736);
nand U25373 (N_25373,N_16856,N_13587);
nand U25374 (N_25374,N_17422,N_12544);
nand U25375 (N_25375,N_17622,N_10857);
and U25376 (N_25376,N_18568,N_19133);
xor U25377 (N_25377,N_15808,N_12489);
or U25378 (N_25378,N_12458,N_12309);
xor U25379 (N_25379,N_17971,N_13962);
or U25380 (N_25380,N_19006,N_17634);
nor U25381 (N_25381,N_10112,N_18823);
nor U25382 (N_25382,N_14642,N_13979);
xnor U25383 (N_25383,N_13539,N_16602);
nor U25384 (N_25384,N_13915,N_19964);
xnor U25385 (N_25385,N_19077,N_13901);
or U25386 (N_25386,N_13294,N_13056);
or U25387 (N_25387,N_16932,N_18723);
nor U25388 (N_25388,N_16010,N_11389);
xor U25389 (N_25389,N_17703,N_12811);
xor U25390 (N_25390,N_10924,N_18935);
xor U25391 (N_25391,N_10650,N_11962);
nand U25392 (N_25392,N_18981,N_19189);
xor U25393 (N_25393,N_11629,N_12876);
xnor U25394 (N_25394,N_12949,N_17522);
xnor U25395 (N_25395,N_14441,N_10488);
or U25396 (N_25396,N_10750,N_19572);
or U25397 (N_25397,N_19570,N_15845);
or U25398 (N_25398,N_12857,N_18484);
or U25399 (N_25399,N_11941,N_14564);
nand U25400 (N_25400,N_18979,N_10814);
and U25401 (N_25401,N_13353,N_16686);
xnor U25402 (N_25402,N_13901,N_19472);
nand U25403 (N_25403,N_15624,N_12149);
xnor U25404 (N_25404,N_18168,N_19144);
nand U25405 (N_25405,N_18258,N_16844);
or U25406 (N_25406,N_19706,N_13680);
or U25407 (N_25407,N_12458,N_17343);
or U25408 (N_25408,N_15047,N_14784);
or U25409 (N_25409,N_19358,N_11334);
and U25410 (N_25410,N_12126,N_17085);
and U25411 (N_25411,N_18761,N_11463);
xnor U25412 (N_25412,N_17080,N_17656);
and U25413 (N_25413,N_12414,N_12853);
xor U25414 (N_25414,N_14408,N_14038);
or U25415 (N_25415,N_15681,N_14089);
and U25416 (N_25416,N_14297,N_16693);
nor U25417 (N_25417,N_10780,N_13681);
nor U25418 (N_25418,N_17532,N_11026);
or U25419 (N_25419,N_12126,N_13840);
and U25420 (N_25420,N_11036,N_13967);
or U25421 (N_25421,N_14350,N_14962);
or U25422 (N_25422,N_16956,N_11546);
xnor U25423 (N_25423,N_16475,N_11198);
nor U25424 (N_25424,N_17607,N_17096);
xnor U25425 (N_25425,N_14872,N_12782);
nor U25426 (N_25426,N_15964,N_14571);
nand U25427 (N_25427,N_11160,N_18959);
or U25428 (N_25428,N_15837,N_16255);
or U25429 (N_25429,N_18840,N_10172);
xor U25430 (N_25430,N_15101,N_19724);
nor U25431 (N_25431,N_14520,N_18302);
nand U25432 (N_25432,N_14519,N_18514);
nor U25433 (N_25433,N_15306,N_17030);
nand U25434 (N_25434,N_13470,N_19295);
xnor U25435 (N_25435,N_18603,N_11745);
nand U25436 (N_25436,N_19005,N_16798);
nor U25437 (N_25437,N_16350,N_18093);
or U25438 (N_25438,N_15721,N_14306);
nand U25439 (N_25439,N_14479,N_15345);
nand U25440 (N_25440,N_19241,N_11697);
or U25441 (N_25441,N_15670,N_14836);
nand U25442 (N_25442,N_16323,N_18588);
and U25443 (N_25443,N_13134,N_11971);
nand U25444 (N_25444,N_19981,N_16012);
xor U25445 (N_25445,N_11843,N_19170);
nor U25446 (N_25446,N_10039,N_15627);
xor U25447 (N_25447,N_10207,N_18213);
xnor U25448 (N_25448,N_16476,N_18743);
and U25449 (N_25449,N_14085,N_16776);
and U25450 (N_25450,N_10178,N_16303);
nor U25451 (N_25451,N_19191,N_12224);
nand U25452 (N_25452,N_12341,N_13343);
nor U25453 (N_25453,N_18477,N_11716);
or U25454 (N_25454,N_19340,N_18901);
nand U25455 (N_25455,N_16162,N_19249);
or U25456 (N_25456,N_12448,N_17857);
nand U25457 (N_25457,N_13082,N_14351);
or U25458 (N_25458,N_18478,N_12948);
or U25459 (N_25459,N_16438,N_15805);
xnor U25460 (N_25460,N_13481,N_10027);
xnor U25461 (N_25461,N_17669,N_13576);
xor U25462 (N_25462,N_15324,N_14756);
nand U25463 (N_25463,N_18571,N_10640);
and U25464 (N_25464,N_15811,N_10476);
or U25465 (N_25465,N_15680,N_18150);
and U25466 (N_25466,N_10822,N_13700);
or U25467 (N_25467,N_12880,N_16777);
and U25468 (N_25468,N_16746,N_14177);
xnor U25469 (N_25469,N_15969,N_19914);
xor U25470 (N_25470,N_15658,N_12584);
and U25471 (N_25471,N_16902,N_11252);
and U25472 (N_25472,N_11851,N_17509);
and U25473 (N_25473,N_19012,N_15523);
nand U25474 (N_25474,N_16599,N_16248);
and U25475 (N_25475,N_11050,N_10938);
nor U25476 (N_25476,N_17801,N_13670);
xor U25477 (N_25477,N_11790,N_17504);
xor U25478 (N_25478,N_11595,N_11237);
nor U25479 (N_25479,N_15548,N_19282);
nor U25480 (N_25480,N_17299,N_18534);
xnor U25481 (N_25481,N_19536,N_14751);
or U25482 (N_25482,N_16651,N_14620);
or U25483 (N_25483,N_14440,N_12772);
or U25484 (N_25484,N_18411,N_12082);
nor U25485 (N_25485,N_13904,N_17562);
nand U25486 (N_25486,N_16112,N_19287);
or U25487 (N_25487,N_18520,N_10062);
nand U25488 (N_25488,N_17089,N_18409);
and U25489 (N_25489,N_18620,N_13954);
or U25490 (N_25490,N_11043,N_18331);
nor U25491 (N_25491,N_16871,N_11731);
nand U25492 (N_25492,N_10616,N_12995);
xnor U25493 (N_25493,N_17881,N_15242);
nand U25494 (N_25494,N_17236,N_10966);
or U25495 (N_25495,N_10098,N_13993);
nand U25496 (N_25496,N_14256,N_17205);
nor U25497 (N_25497,N_17799,N_15227);
and U25498 (N_25498,N_12932,N_14572);
and U25499 (N_25499,N_17400,N_13470);
nand U25500 (N_25500,N_15168,N_19223);
and U25501 (N_25501,N_19543,N_16377);
nor U25502 (N_25502,N_16896,N_16519);
nand U25503 (N_25503,N_16375,N_18390);
and U25504 (N_25504,N_16042,N_12442);
xor U25505 (N_25505,N_12021,N_13597);
xnor U25506 (N_25506,N_14262,N_11347);
xnor U25507 (N_25507,N_18486,N_16384);
or U25508 (N_25508,N_11935,N_12478);
nor U25509 (N_25509,N_16471,N_10573);
nand U25510 (N_25510,N_13831,N_17358);
xor U25511 (N_25511,N_15475,N_13413);
or U25512 (N_25512,N_12034,N_14205);
or U25513 (N_25513,N_15720,N_12995);
or U25514 (N_25514,N_16801,N_16359);
and U25515 (N_25515,N_17901,N_14004);
and U25516 (N_25516,N_10826,N_11178);
nor U25517 (N_25517,N_11574,N_16690);
nor U25518 (N_25518,N_19341,N_12802);
or U25519 (N_25519,N_16888,N_18270);
and U25520 (N_25520,N_12201,N_13333);
nand U25521 (N_25521,N_11570,N_16673);
xor U25522 (N_25522,N_10455,N_13139);
xnor U25523 (N_25523,N_19513,N_15722);
nand U25524 (N_25524,N_12748,N_13182);
or U25525 (N_25525,N_14485,N_16630);
nor U25526 (N_25526,N_14753,N_19413);
or U25527 (N_25527,N_19012,N_12419);
nor U25528 (N_25528,N_11559,N_14333);
or U25529 (N_25529,N_15861,N_11049);
or U25530 (N_25530,N_11185,N_18478);
or U25531 (N_25531,N_17000,N_13891);
nor U25532 (N_25532,N_10791,N_13562);
xor U25533 (N_25533,N_17960,N_12765);
nor U25534 (N_25534,N_10402,N_17723);
nor U25535 (N_25535,N_19751,N_12852);
nand U25536 (N_25536,N_11356,N_18713);
nand U25537 (N_25537,N_15172,N_11990);
xnor U25538 (N_25538,N_16611,N_11931);
nand U25539 (N_25539,N_15562,N_17848);
xnor U25540 (N_25540,N_18643,N_11991);
xor U25541 (N_25541,N_17940,N_11947);
or U25542 (N_25542,N_11516,N_19138);
nor U25543 (N_25543,N_17048,N_14061);
nand U25544 (N_25544,N_17345,N_14768);
nand U25545 (N_25545,N_14445,N_10934);
nand U25546 (N_25546,N_17237,N_11173);
nor U25547 (N_25547,N_18587,N_10928);
and U25548 (N_25548,N_14616,N_12727);
nand U25549 (N_25549,N_14046,N_12303);
or U25550 (N_25550,N_17539,N_18209);
xor U25551 (N_25551,N_15043,N_13602);
and U25552 (N_25552,N_16897,N_16859);
or U25553 (N_25553,N_17403,N_15270);
or U25554 (N_25554,N_17303,N_19148);
or U25555 (N_25555,N_12774,N_12668);
and U25556 (N_25556,N_15801,N_17666);
or U25557 (N_25557,N_18474,N_11986);
or U25558 (N_25558,N_13748,N_11253);
nor U25559 (N_25559,N_19181,N_19474);
xnor U25560 (N_25560,N_15775,N_19549);
nor U25561 (N_25561,N_15359,N_13897);
nand U25562 (N_25562,N_11301,N_18668);
nand U25563 (N_25563,N_12688,N_11326);
or U25564 (N_25564,N_13241,N_11719);
nand U25565 (N_25565,N_11511,N_11995);
or U25566 (N_25566,N_11441,N_13515);
xnor U25567 (N_25567,N_10404,N_15026);
and U25568 (N_25568,N_18049,N_10737);
and U25569 (N_25569,N_17505,N_11749);
nor U25570 (N_25570,N_14332,N_11629);
nor U25571 (N_25571,N_11303,N_17287);
nor U25572 (N_25572,N_14083,N_12724);
xnor U25573 (N_25573,N_13295,N_19216);
nand U25574 (N_25574,N_13498,N_11070);
nor U25575 (N_25575,N_12381,N_19224);
or U25576 (N_25576,N_14802,N_11236);
nor U25577 (N_25577,N_12918,N_15090);
xnor U25578 (N_25578,N_18887,N_17373);
xor U25579 (N_25579,N_13814,N_12360);
nor U25580 (N_25580,N_14546,N_11555);
or U25581 (N_25581,N_17416,N_12304);
xor U25582 (N_25582,N_17483,N_13595);
and U25583 (N_25583,N_12274,N_13236);
and U25584 (N_25584,N_10645,N_17479);
nand U25585 (N_25585,N_11425,N_15402);
nand U25586 (N_25586,N_15682,N_14710);
nand U25587 (N_25587,N_17619,N_14074);
xor U25588 (N_25588,N_19167,N_17300);
nor U25589 (N_25589,N_18032,N_15843);
nor U25590 (N_25590,N_11137,N_15550);
nand U25591 (N_25591,N_13786,N_13570);
xnor U25592 (N_25592,N_19977,N_15240);
xnor U25593 (N_25593,N_13160,N_19864);
nor U25594 (N_25594,N_18043,N_10441);
nand U25595 (N_25595,N_10982,N_11110);
nand U25596 (N_25596,N_13765,N_15541);
nand U25597 (N_25597,N_10192,N_16733);
or U25598 (N_25598,N_17844,N_14020);
or U25599 (N_25599,N_15023,N_17367);
xor U25600 (N_25600,N_11791,N_18652);
nor U25601 (N_25601,N_10165,N_18235);
or U25602 (N_25602,N_12112,N_13266);
xnor U25603 (N_25603,N_10105,N_15607);
nor U25604 (N_25604,N_17670,N_16712);
or U25605 (N_25605,N_17377,N_12042);
and U25606 (N_25606,N_13489,N_11467);
nor U25607 (N_25607,N_19954,N_15316);
nand U25608 (N_25608,N_16774,N_18913);
and U25609 (N_25609,N_12251,N_14036);
nor U25610 (N_25610,N_19640,N_13113);
and U25611 (N_25611,N_10997,N_19584);
nand U25612 (N_25612,N_18678,N_13161);
nor U25613 (N_25613,N_16570,N_11640);
nand U25614 (N_25614,N_19444,N_13938);
nand U25615 (N_25615,N_16171,N_18956);
nor U25616 (N_25616,N_11034,N_17016);
xnor U25617 (N_25617,N_18011,N_17558);
xor U25618 (N_25618,N_15462,N_16280);
and U25619 (N_25619,N_19154,N_10670);
nand U25620 (N_25620,N_15681,N_12442);
nor U25621 (N_25621,N_16404,N_13164);
xor U25622 (N_25622,N_16544,N_11730);
nand U25623 (N_25623,N_14420,N_13481);
xor U25624 (N_25624,N_12378,N_17258);
nor U25625 (N_25625,N_13629,N_17623);
nand U25626 (N_25626,N_18577,N_10097);
xor U25627 (N_25627,N_19170,N_13105);
or U25628 (N_25628,N_19071,N_12315);
or U25629 (N_25629,N_19200,N_11246);
xor U25630 (N_25630,N_14611,N_18566);
nand U25631 (N_25631,N_10515,N_12022);
nor U25632 (N_25632,N_13945,N_14854);
or U25633 (N_25633,N_14959,N_11252);
nand U25634 (N_25634,N_18892,N_12927);
xnor U25635 (N_25635,N_19501,N_18593);
xor U25636 (N_25636,N_11837,N_10844);
nor U25637 (N_25637,N_18602,N_10132);
nor U25638 (N_25638,N_16256,N_19637);
xnor U25639 (N_25639,N_19256,N_18421);
nor U25640 (N_25640,N_10518,N_12083);
and U25641 (N_25641,N_15997,N_13549);
and U25642 (N_25642,N_17731,N_19284);
xnor U25643 (N_25643,N_18484,N_16325);
or U25644 (N_25644,N_14062,N_14154);
nand U25645 (N_25645,N_15959,N_16365);
nand U25646 (N_25646,N_14380,N_10860);
nor U25647 (N_25647,N_19720,N_16874);
nor U25648 (N_25648,N_16948,N_18152);
or U25649 (N_25649,N_12617,N_11566);
and U25650 (N_25650,N_15496,N_15387);
or U25651 (N_25651,N_14581,N_13872);
or U25652 (N_25652,N_13743,N_19105);
nor U25653 (N_25653,N_17717,N_10355);
xor U25654 (N_25654,N_12846,N_16774);
nand U25655 (N_25655,N_18133,N_16994);
xnor U25656 (N_25656,N_17006,N_17867);
nor U25657 (N_25657,N_11024,N_16053);
and U25658 (N_25658,N_11661,N_19024);
xnor U25659 (N_25659,N_11950,N_13538);
or U25660 (N_25660,N_12075,N_15828);
xor U25661 (N_25661,N_19549,N_10727);
and U25662 (N_25662,N_16610,N_11816);
nand U25663 (N_25663,N_12079,N_12453);
and U25664 (N_25664,N_13715,N_13074);
or U25665 (N_25665,N_12945,N_14128);
nor U25666 (N_25666,N_17220,N_16771);
nand U25667 (N_25667,N_16858,N_16497);
nor U25668 (N_25668,N_12699,N_15646);
nand U25669 (N_25669,N_15210,N_16815);
and U25670 (N_25670,N_17684,N_18671);
nand U25671 (N_25671,N_14876,N_11708);
and U25672 (N_25672,N_18792,N_15548);
or U25673 (N_25673,N_14598,N_17567);
nor U25674 (N_25674,N_13499,N_17868);
nor U25675 (N_25675,N_10149,N_17931);
and U25676 (N_25676,N_15948,N_16924);
nand U25677 (N_25677,N_12055,N_19704);
nor U25678 (N_25678,N_11853,N_18338);
or U25679 (N_25679,N_14979,N_10113);
and U25680 (N_25680,N_18946,N_16095);
nand U25681 (N_25681,N_14730,N_15926);
nand U25682 (N_25682,N_15367,N_10721);
nor U25683 (N_25683,N_13330,N_16819);
nand U25684 (N_25684,N_16262,N_14435);
xor U25685 (N_25685,N_12410,N_10443);
or U25686 (N_25686,N_11198,N_11813);
nor U25687 (N_25687,N_10926,N_19194);
and U25688 (N_25688,N_17779,N_17292);
nor U25689 (N_25689,N_19764,N_18680);
or U25690 (N_25690,N_12799,N_15709);
nand U25691 (N_25691,N_14669,N_19116);
nor U25692 (N_25692,N_15752,N_17928);
or U25693 (N_25693,N_10188,N_12442);
nand U25694 (N_25694,N_10622,N_15688);
or U25695 (N_25695,N_18496,N_19132);
and U25696 (N_25696,N_16165,N_11902);
and U25697 (N_25697,N_12086,N_11279);
xor U25698 (N_25698,N_16181,N_16504);
nor U25699 (N_25699,N_17494,N_17320);
and U25700 (N_25700,N_15892,N_11865);
nor U25701 (N_25701,N_13452,N_16790);
xnor U25702 (N_25702,N_12863,N_16536);
xor U25703 (N_25703,N_16349,N_18246);
nand U25704 (N_25704,N_18502,N_10781);
nor U25705 (N_25705,N_12015,N_17471);
nand U25706 (N_25706,N_12346,N_11552);
nand U25707 (N_25707,N_14519,N_18919);
nor U25708 (N_25708,N_17826,N_16624);
and U25709 (N_25709,N_14069,N_11766);
and U25710 (N_25710,N_11141,N_11482);
xnor U25711 (N_25711,N_17186,N_13782);
nand U25712 (N_25712,N_10089,N_15592);
nand U25713 (N_25713,N_13609,N_12926);
and U25714 (N_25714,N_17145,N_12534);
nand U25715 (N_25715,N_11274,N_12587);
or U25716 (N_25716,N_16500,N_18530);
xnor U25717 (N_25717,N_17690,N_19508);
nand U25718 (N_25718,N_11185,N_10334);
or U25719 (N_25719,N_18486,N_10292);
or U25720 (N_25720,N_13592,N_16420);
nor U25721 (N_25721,N_16666,N_13389);
nand U25722 (N_25722,N_17383,N_12158);
and U25723 (N_25723,N_17326,N_16561);
and U25724 (N_25724,N_10970,N_16486);
xnor U25725 (N_25725,N_18778,N_15689);
xor U25726 (N_25726,N_15176,N_12839);
and U25727 (N_25727,N_13127,N_10431);
nand U25728 (N_25728,N_11805,N_15154);
xor U25729 (N_25729,N_19634,N_19334);
nand U25730 (N_25730,N_16336,N_15607);
xnor U25731 (N_25731,N_11996,N_13760);
nor U25732 (N_25732,N_10590,N_18967);
nor U25733 (N_25733,N_11272,N_17337);
xnor U25734 (N_25734,N_12239,N_17539);
nand U25735 (N_25735,N_13466,N_14014);
nand U25736 (N_25736,N_11047,N_17074);
xnor U25737 (N_25737,N_14379,N_12503);
nand U25738 (N_25738,N_15508,N_11705);
or U25739 (N_25739,N_16783,N_10452);
nand U25740 (N_25740,N_18784,N_13065);
nor U25741 (N_25741,N_13336,N_11125);
and U25742 (N_25742,N_14360,N_18409);
nand U25743 (N_25743,N_19021,N_15302);
xor U25744 (N_25744,N_13847,N_12709);
xor U25745 (N_25745,N_10237,N_11543);
xnor U25746 (N_25746,N_17421,N_18552);
nand U25747 (N_25747,N_11729,N_14224);
nor U25748 (N_25748,N_18018,N_12648);
xnor U25749 (N_25749,N_18286,N_16574);
nand U25750 (N_25750,N_12739,N_19704);
xor U25751 (N_25751,N_12440,N_18453);
nand U25752 (N_25752,N_15360,N_12595);
or U25753 (N_25753,N_12592,N_18801);
xnor U25754 (N_25754,N_13875,N_14013);
nand U25755 (N_25755,N_10456,N_15162);
nand U25756 (N_25756,N_12113,N_12771);
and U25757 (N_25757,N_13174,N_16075);
and U25758 (N_25758,N_14978,N_16635);
and U25759 (N_25759,N_18758,N_12970);
xor U25760 (N_25760,N_17265,N_15867);
xor U25761 (N_25761,N_19181,N_13736);
xnor U25762 (N_25762,N_18282,N_14127);
nand U25763 (N_25763,N_11478,N_17911);
or U25764 (N_25764,N_18293,N_17535);
or U25765 (N_25765,N_15785,N_10306);
or U25766 (N_25766,N_10581,N_10445);
nor U25767 (N_25767,N_18623,N_14520);
nand U25768 (N_25768,N_19269,N_18153);
or U25769 (N_25769,N_17515,N_14032);
and U25770 (N_25770,N_17389,N_11139);
nor U25771 (N_25771,N_18242,N_18831);
or U25772 (N_25772,N_13684,N_16580);
and U25773 (N_25773,N_17682,N_13128);
nand U25774 (N_25774,N_18315,N_17585);
nand U25775 (N_25775,N_17233,N_12903);
xnor U25776 (N_25776,N_16694,N_11153);
and U25777 (N_25777,N_10239,N_14624);
and U25778 (N_25778,N_17004,N_14608);
xor U25779 (N_25779,N_13245,N_19608);
and U25780 (N_25780,N_15730,N_14483);
and U25781 (N_25781,N_16180,N_14986);
nand U25782 (N_25782,N_11107,N_19421);
xnor U25783 (N_25783,N_10921,N_17543);
and U25784 (N_25784,N_14575,N_16744);
nand U25785 (N_25785,N_15631,N_15865);
and U25786 (N_25786,N_13688,N_14922);
xor U25787 (N_25787,N_17959,N_10000);
and U25788 (N_25788,N_13939,N_12140);
or U25789 (N_25789,N_10911,N_15136);
or U25790 (N_25790,N_17844,N_12693);
xor U25791 (N_25791,N_12003,N_12004);
or U25792 (N_25792,N_13581,N_19921);
xnor U25793 (N_25793,N_16109,N_13162);
nor U25794 (N_25794,N_10659,N_16115);
or U25795 (N_25795,N_11573,N_16627);
xnor U25796 (N_25796,N_10625,N_10003);
and U25797 (N_25797,N_16244,N_16625);
or U25798 (N_25798,N_10091,N_11500);
nor U25799 (N_25799,N_10512,N_17173);
or U25800 (N_25800,N_16395,N_12656);
xnor U25801 (N_25801,N_12664,N_13675);
nor U25802 (N_25802,N_19048,N_12311);
nor U25803 (N_25803,N_19982,N_10793);
or U25804 (N_25804,N_19081,N_14152);
and U25805 (N_25805,N_16291,N_13516);
and U25806 (N_25806,N_14376,N_11503);
nand U25807 (N_25807,N_14744,N_13327);
xor U25808 (N_25808,N_15936,N_18884);
and U25809 (N_25809,N_17059,N_11982);
xnor U25810 (N_25810,N_15632,N_14140);
nor U25811 (N_25811,N_10398,N_10294);
or U25812 (N_25812,N_14436,N_11040);
nor U25813 (N_25813,N_16595,N_10640);
xnor U25814 (N_25814,N_11059,N_15197);
nand U25815 (N_25815,N_18738,N_17499);
or U25816 (N_25816,N_18597,N_15547);
nand U25817 (N_25817,N_10939,N_11789);
and U25818 (N_25818,N_11352,N_16699);
xor U25819 (N_25819,N_16367,N_15912);
nor U25820 (N_25820,N_19754,N_16357);
xnor U25821 (N_25821,N_13477,N_11758);
nor U25822 (N_25822,N_17170,N_11763);
xor U25823 (N_25823,N_18969,N_11926);
xnor U25824 (N_25824,N_10656,N_14238);
or U25825 (N_25825,N_19370,N_15362);
or U25826 (N_25826,N_12249,N_16918);
nor U25827 (N_25827,N_10928,N_16333);
nand U25828 (N_25828,N_12189,N_18191);
nand U25829 (N_25829,N_15383,N_13987);
or U25830 (N_25830,N_12468,N_17542);
or U25831 (N_25831,N_11614,N_16932);
nand U25832 (N_25832,N_17709,N_13118);
nor U25833 (N_25833,N_11640,N_16978);
nor U25834 (N_25834,N_14795,N_12545);
or U25835 (N_25835,N_14320,N_12920);
or U25836 (N_25836,N_10830,N_17320);
xnor U25837 (N_25837,N_12686,N_16133);
or U25838 (N_25838,N_10596,N_13515);
nor U25839 (N_25839,N_10839,N_19697);
and U25840 (N_25840,N_14733,N_19641);
nor U25841 (N_25841,N_17742,N_11682);
and U25842 (N_25842,N_18915,N_15736);
nor U25843 (N_25843,N_17949,N_13648);
nand U25844 (N_25844,N_10183,N_10667);
nand U25845 (N_25845,N_12968,N_13034);
nor U25846 (N_25846,N_11346,N_11654);
or U25847 (N_25847,N_19489,N_13284);
or U25848 (N_25848,N_18140,N_14217);
xnor U25849 (N_25849,N_13840,N_17141);
nand U25850 (N_25850,N_17746,N_16064);
and U25851 (N_25851,N_10085,N_19563);
nand U25852 (N_25852,N_16501,N_12152);
xor U25853 (N_25853,N_17325,N_17513);
nand U25854 (N_25854,N_15105,N_14574);
and U25855 (N_25855,N_13881,N_15616);
and U25856 (N_25856,N_18639,N_13296);
nor U25857 (N_25857,N_16356,N_12032);
xor U25858 (N_25858,N_12070,N_19520);
nand U25859 (N_25859,N_16406,N_15662);
xor U25860 (N_25860,N_13571,N_11574);
xor U25861 (N_25861,N_12121,N_17728);
and U25862 (N_25862,N_15645,N_13451);
nor U25863 (N_25863,N_11287,N_14687);
and U25864 (N_25864,N_17521,N_15662);
and U25865 (N_25865,N_17262,N_16001);
or U25866 (N_25866,N_11951,N_19955);
nor U25867 (N_25867,N_10493,N_19643);
nor U25868 (N_25868,N_12690,N_13406);
and U25869 (N_25869,N_12728,N_12006);
and U25870 (N_25870,N_19511,N_18779);
and U25871 (N_25871,N_17845,N_14969);
nand U25872 (N_25872,N_16667,N_11573);
nor U25873 (N_25873,N_11347,N_13900);
xor U25874 (N_25874,N_13798,N_18566);
xor U25875 (N_25875,N_14909,N_11435);
or U25876 (N_25876,N_11387,N_14629);
and U25877 (N_25877,N_13562,N_13460);
or U25878 (N_25878,N_16275,N_17040);
or U25879 (N_25879,N_10824,N_12980);
or U25880 (N_25880,N_15405,N_16184);
xnor U25881 (N_25881,N_12400,N_13060);
nor U25882 (N_25882,N_18549,N_19072);
or U25883 (N_25883,N_15137,N_14679);
and U25884 (N_25884,N_10799,N_12463);
nand U25885 (N_25885,N_11643,N_12982);
and U25886 (N_25886,N_17274,N_13701);
nor U25887 (N_25887,N_12473,N_14352);
xor U25888 (N_25888,N_12266,N_10376);
nand U25889 (N_25889,N_13971,N_13263);
xnor U25890 (N_25890,N_19404,N_19899);
and U25891 (N_25891,N_18992,N_19938);
nand U25892 (N_25892,N_18986,N_17554);
xnor U25893 (N_25893,N_17865,N_15490);
nand U25894 (N_25894,N_18770,N_11913);
xor U25895 (N_25895,N_13817,N_17164);
or U25896 (N_25896,N_19345,N_15163);
and U25897 (N_25897,N_14208,N_13143);
and U25898 (N_25898,N_11363,N_16417);
nor U25899 (N_25899,N_18265,N_12017);
xor U25900 (N_25900,N_11274,N_11602);
xnor U25901 (N_25901,N_16121,N_19617);
nand U25902 (N_25902,N_16659,N_15005);
nor U25903 (N_25903,N_13454,N_18555);
nor U25904 (N_25904,N_17847,N_19746);
nor U25905 (N_25905,N_19192,N_14752);
and U25906 (N_25906,N_18992,N_13777);
or U25907 (N_25907,N_17024,N_18483);
or U25908 (N_25908,N_11818,N_14041);
and U25909 (N_25909,N_17264,N_18661);
nor U25910 (N_25910,N_13376,N_11058);
or U25911 (N_25911,N_13087,N_18743);
and U25912 (N_25912,N_19900,N_14460);
nor U25913 (N_25913,N_19669,N_18374);
nand U25914 (N_25914,N_11902,N_10097);
nand U25915 (N_25915,N_17544,N_11591);
or U25916 (N_25916,N_13515,N_19445);
xnor U25917 (N_25917,N_16050,N_16513);
or U25918 (N_25918,N_18266,N_15249);
nand U25919 (N_25919,N_15464,N_11942);
xnor U25920 (N_25920,N_17560,N_13671);
nand U25921 (N_25921,N_15855,N_17110);
nand U25922 (N_25922,N_13773,N_16100);
nor U25923 (N_25923,N_16169,N_14639);
nor U25924 (N_25924,N_11007,N_15915);
or U25925 (N_25925,N_14467,N_10340);
nor U25926 (N_25926,N_14784,N_14906);
xor U25927 (N_25927,N_15141,N_19467);
nor U25928 (N_25928,N_12329,N_19958);
xor U25929 (N_25929,N_11190,N_13529);
nand U25930 (N_25930,N_15871,N_18131);
nor U25931 (N_25931,N_11830,N_15276);
nand U25932 (N_25932,N_13434,N_15239);
xor U25933 (N_25933,N_18735,N_11487);
or U25934 (N_25934,N_12683,N_14360);
nand U25935 (N_25935,N_19564,N_17544);
and U25936 (N_25936,N_16150,N_13381);
or U25937 (N_25937,N_17373,N_19822);
nor U25938 (N_25938,N_19652,N_10919);
nor U25939 (N_25939,N_15509,N_13438);
xnor U25940 (N_25940,N_16103,N_13591);
xor U25941 (N_25941,N_13154,N_11997);
xnor U25942 (N_25942,N_16341,N_17785);
and U25943 (N_25943,N_12592,N_16543);
nand U25944 (N_25944,N_16684,N_13821);
nand U25945 (N_25945,N_11663,N_13286);
or U25946 (N_25946,N_18383,N_15260);
nand U25947 (N_25947,N_12352,N_16500);
xor U25948 (N_25948,N_12436,N_16389);
nand U25949 (N_25949,N_15327,N_11022);
nand U25950 (N_25950,N_15825,N_13260);
and U25951 (N_25951,N_14196,N_18672);
and U25952 (N_25952,N_15199,N_11637);
or U25953 (N_25953,N_13861,N_18191);
xor U25954 (N_25954,N_11358,N_13033);
or U25955 (N_25955,N_15726,N_14246);
xor U25956 (N_25956,N_13563,N_12582);
or U25957 (N_25957,N_16790,N_14644);
and U25958 (N_25958,N_11187,N_15451);
nand U25959 (N_25959,N_15641,N_13021);
xor U25960 (N_25960,N_10650,N_19025);
and U25961 (N_25961,N_15129,N_11474);
or U25962 (N_25962,N_18065,N_10990);
xnor U25963 (N_25963,N_18908,N_11315);
or U25964 (N_25964,N_18484,N_13402);
nor U25965 (N_25965,N_19106,N_14958);
nand U25966 (N_25966,N_11948,N_12837);
nor U25967 (N_25967,N_16600,N_11762);
or U25968 (N_25968,N_15681,N_13251);
nand U25969 (N_25969,N_10318,N_15904);
nand U25970 (N_25970,N_15475,N_15705);
nor U25971 (N_25971,N_14826,N_19236);
nand U25972 (N_25972,N_14743,N_14050);
or U25973 (N_25973,N_14767,N_15852);
and U25974 (N_25974,N_19245,N_17890);
or U25975 (N_25975,N_12913,N_10461);
xnor U25976 (N_25976,N_11450,N_11069);
nor U25977 (N_25977,N_19984,N_14801);
xnor U25978 (N_25978,N_12205,N_12894);
nand U25979 (N_25979,N_12053,N_16871);
and U25980 (N_25980,N_15088,N_13980);
xor U25981 (N_25981,N_18640,N_14951);
xor U25982 (N_25982,N_16696,N_17169);
and U25983 (N_25983,N_11655,N_11264);
nor U25984 (N_25984,N_16430,N_11303);
nor U25985 (N_25985,N_14719,N_10656);
nor U25986 (N_25986,N_13777,N_17380);
xnor U25987 (N_25987,N_11871,N_17345);
nand U25988 (N_25988,N_19542,N_13222);
nor U25989 (N_25989,N_17533,N_13797);
xnor U25990 (N_25990,N_12657,N_14922);
xor U25991 (N_25991,N_13469,N_15332);
nor U25992 (N_25992,N_12311,N_17677);
or U25993 (N_25993,N_14352,N_15470);
and U25994 (N_25994,N_14452,N_16223);
nand U25995 (N_25995,N_16827,N_10305);
and U25996 (N_25996,N_18519,N_17614);
nand U25997 (N_25997,N_18750,N_17995);
xor U25998 (N_25998,N_12871,N_14028);
nand U25999 (N_25999,N_14427,N_19020);
nand U26000 (N_26000,N_11038,N_15981);
xor U26001 (N_26001,N_17670,N_11517);
nand U26002 (N_26002,N_15578,N_10706);
or U26003 (N_26003,N_17946,N_12475);
nor U26004 (N_26004,N_15943,N_12147);
xnor U26005 (N_26005,N_18026,N_14649);
or U26006 (N_26006,N_18883,N_17444);
xor U26007 (N_26007,N_14056,N_15889);
and U26008 (N_26008,N_14949,N_17337);
xnor U26009 (N_26009,N_14161,N_16820);
and U26010 (N_26010,N_15076,N_12679);
and U26011 (N_26011,N_10881,N_14367);
xor U26012 (N_26012,N_18029,N_10071);
xor U26013 (N_26013,N_11977,N_16509);
xor U26014 (N_26014,N_14118,N_10922);
xor U26015 (N_26015,N_19858,N_14483);
and U26016 (N_26016,N_15855,N_13929);
xor U26017 (N_26017,N_10608,N_16475);
nand U26018 (N_26018,N_15788,N_14317);
xnor U26019 (N_26019,N_17406,N_12509);
xnor U26020 (N_26020,N_12716,N_11015);
and U26021 (N_26021,N_11697,N_19297);
and U26022 (N_26022,N_15403,N_11898);
xor U26023 (N_26023,N_19357,N_10181);
xnor U26024 (N_26024,N_16156,N_13674);
nand U26025 (N_26025,N_10030,N_12276);
and U26026 (N_26026,N_10192,N_11474);
and U26027 (N_26027,N_19468,N_19192);
or U26028 (N_26028,N_17940,N_17163);
and U26029 (N_26029,N_14578,N_15181);
nor U26030 (N_26030,N_17986,N_15377);
xor U26031 (N_26031,N_19992,N_10478);
nor U26032 (N_26032,N_16405,N_17705);
or U26033 (N_26033,N_17182,N_12146);
xnor U26034 (N_26034,N_14081,N_15716);
xnor U26035 (N_26035,N_15896,N_14299);
nand U26036 (N_26036,N_10254,N_13508);
and U26037 (N_26037,N_17483,N_18066);
and U26038 (N_26038,N_15514,N_12116);
nor U26039 (N_26039,N_10718,N_15892);
nand U26040 (N_26040,N_15929,N_18471);
and U26041 (N_26041,N_13504,N_11528);
or U26042 (N_26042,N_16440,N_10765);
nand U26043 (N_26043,N_12866,N_15320);
or U26044 (N_26044,N_13876,N_17226);
nor U26045 (N_26045,N_17081,N_11645);
nor U26046 (N_26046,N_12817,N_15621);
nand U26047 (N_26047,N_15816,N_11095);
xnor U26048 (N_26048,N_18152,N_10422);
or U26049 (N_26049,N_19552,N_19052);
nand U26050 (N_26050,N_10464,N_10594);
nor U26051 (N_26051,N_15256,N_19315);
nand U26052 (N_26052,N_12498,N_18163);
and U26053 (N_26053,N_19834,N_12103);
or U26054 (N_26054,N_10311,N_11541);
and U26055 (N_26055,N_15999,N_17415);
and U26056 (N_26056,N_10064,N_14020);
nand U26057 (N_26057,N_18483,N_16871);
xnor U26058 (N_26058,N_13613,N_13609);
nor U26059 (N_26059,N_15926,N_17386);
or U26060 (N_26060,N_17474,N_14858);
xor U26061 (N_26061,N_10393,N_11465);
nand U26062 (N_26062,N_18870,N_13016);
and U26063 (N_26063,N_17407,N_19323);
xor U26064 (N_26064,N_12349,N_17882);
nand U26065 (N_26065,N_18552,N_19119);
xnor U26066 (N_26066,N_18960,N_13492);
and U26067 (N_26067,N_18767,N_10402);
nor U26068 (N_26068,N_14655,N_14849);
and U26069 (N_26069,N_14695,N_13899);
xnor U26070 (N_26070,N_10776,N_18687);
xor U26071 (N_26071,N_11514,N_17329);
xnor U26072 (N_26072,N_12291,N_18332);
xor U26073 (N_26073,N_16484,N_13271);
nand U26074 (N_26074,N_17970,N_16066);
nor U26075 (N_26075,N_12465,N_17099);
nor U26076 (N_26076,N_15550,N_19211);
nor U26077 (N_26077,N_15876,N_14197);
nor U26078 (N_26078,N_17227,N_19360);
nand U26079 (N_26079,N_13091,N_10490);
and U26080 (N_26080,N_17282,N_19066);
and U26081 (N_26081,N_16433,N_10732);
or U26082 (N_26082,N_11798,N_14717);
nand U26083 (N_26083,N_16017,N_19326);
xor U26084 (N_26084,N_16572,N_17661);
nand U26085 (N_26085,N_18306,N_15019);
nand U26086 (N_26086,N_12020,N_16388);
nand U26087 (N_26087,N_19190,N_14605);
nor U26088 (N_26088,N_14411,N_11844);
xnor U26089 (N_26089,N_13772,N_11903);
or U26090 (N_26090,N_15674,N_17826);
nor U26091 (N_26091,N_14675,N_16161);
nor U26092 (N_26092,N_14067,N_14339);
and U26093 (N_26093,N_12968,N_15618);
nand U26094 (N_26094,N_10297,N_17480);
or U26095 (N_26095,N_13092,N_16257);
or U26096 (N_26096,N_13836,N_12986);
nand U26097 (N_26097,N_12561,N_11822);
nor U26098 (N_26098,N_19567,N_15016);
nand U26099 (N_26099,N_19020,N_19735);
and U26100 (N_26100,N_19342,N_13600);
nand U26101 (N_26101,N_18614,N_18882);
nand U26102 (N_26102,N_12058,N_14009);
nand U26103 (N_26103,N_13528,N_15723);
or U26104 (N_26104,N_14375,N_18088);
and U26105 (N_26105,N_13134,N_18517);
nand U26106 (N_26106,N_11654,N_10975);
and U26107 (N_26107,N_13530,N_15242);
nand U26108 (N_26108,N_13877,N_13722);
nor U26109 (N_26109,N_17307,N_15365);
and U26110 (N_26110,N_19711,N_12190);
or U26111 (N_26111,N_14983,N_15556);
xor U26112 (N_26112,N_16082,N_11381);
xor U26113 (N_26113,N_10510,N_13909);
nor U26114 (N_26114,N_12216,N_13608);
or U26115 (N_26115,N_10218,N_18234);
nor U26116 (N_26116,N_15278,N_13699);
nor U26117 (N_26117,N_10241,N_11382);
nor U26118 (N_26118,N_12741,N_16768);
xor U26119 (N_26119,N_13089,N_15054);
nand U26120 (N_26120,N_17795,N_18288);
nand U26121 (N_26121,N_15203,N_14636);
and U26122 (N_26122,N_13678,N_16690);
or U26123 (N_26123,N_13495,N_16379);
and U26124 (N_26124,N_13851,N_19791);
nor U26125 (N_26125,N_13288,N_11128);
xnor U26126 (N_26126,N_12152,N_19682);
nand U26127 (N_26127,N_13101,N_16809);
xor U26128 (N_26128,N_19235,N_16171);
or U26129 (N_26129,N_15780,N_16006);
nor U26130 (N_26130,N_11825,N_11516);
nor U26131 (N_26131,N_10341,N_18626);
nor U26132 (N_26132,N_19837,N_10142);
or U26133 (N_26133,N_18119,N_14869);
and U26134 (N_26134,N_15775,N_14244);
or U26135 (N_26135,N_19512,N_10256);
nand U26136 (N_26136,N_13126,N_10423);
or U26137 (N_26137,N_10230,N_11666);
nor U26138 (N_26138,N_10608,N_14400);
or U26139 (N_26139,N_17154,N_19899);
and U26140 (N_26140,N_19102,N_19066);
or U26141 (N_26141,N_10927,N_13429);
nor U26142 (N_26142,N_17583,N_18729);
or U26143 (N_26143,N_15992,N_10655);
nand U26144 (N_26144,N_15744,N_14341);
and U26145 (N_26145,N_18302,N_10919);
nor U26146 (N_26146,N_19159,N_14386);
or U26147 (N_26147,N_19028,N_17622);
or U26148 (N_26148,N_15859,N_10854);
nor U26149 (N_26149,N_17252,N_19567);
nor U26150 (N_26150,N_14119,N_17026);
xor U26151 (N_26151,N_19115,N_12745);
xnor U26152 (N_26152,N_18093,N_19304);
nor U26153 (N_26153,N_13971,N_18274);
xnor U26154 (N_26154,N_10206,N_18728);
nand U26155 (N_26155,N_19270,N_17652);
nand U26156 (N_26156,N_18826,N_11883);
xor U26157 (N_26157,N_19764,N_11736);
nor U26158 (N_26158,N_16096,N_12791);
xor U26159 (N_26159,N_10297,N_19383);
and U26160 (N_26160,N_16199,N_13746);
nor U26161 (N_26161,N_11248,N_13816);
nor U26162 (N_26162,N_19577,N_14354);
and U26163 (N_26163,N_16777,N_13893);
xor U26164 (N_26164,N_14063,N_18325);
xor U26165 (N_26165,N_17028,N_13369);
xnor U26166 (N_26166,N_18862,N_12096);
xnor U26167 (N_26167,N_10588,N_19732);
nand U26168 (N_26168,N_13152,N_17029);
and U26169 (N_26169,N_15470,N_12009);
or U26170 (N_26170,N_12832,N_10786);
xnor U26171 (N_26171,N_17172,N_13812);
and U26172 (N_26172,N_14091,N_14760);
or U26173 (N_26173,N_19401,N_13785);
xnor U26174 (N_26174,N_17516,N_16854);
nor U26175 (N_26175,N_13589,N_17272);
nand U26176 (N_26176,N_11499,N_15083);
or U26177 (N_26177,N_10754,N_14852);
nand U26178 (N_26178,N_15239,N_10679);
nor U26179 (N_26179,N_16159,N_17280);
nand U26180 (N_26180,N_11253,N_11706);
xor U26181 (N_26181,N_13567,N_11210);
or U26182 (N_26182,N_12608,N_15608);
and U26183 (N_26183,N_15060,N_10744);
nand U26184 (N_26184,N_19735,N_19670);
and U26185 (N_26185,N_10561,N_13539);
nor U26186 (N_26186,N_12188,N_18178);
nand U26187 (N_26187,N_18737,N_16859);
xnor U26188 (N_26188,N_16309,N_17130);
nand U26189 (N_26189,N_19189,N_14636);
or U26190 (N_26190,N_13884,N_19334);
and U26191 (N_26191,N_15694,N_14348);
or U26192 (N_26192,N_13717,N_17498);
or U26193 (N_26193,N_14447,N_19118);
xor U26194 (N_26194,N_16592,N_18056);
or U26195 (N_26195,N_10037,N_19656);
xor U26196 (N_26196,N_16165,N_10748);
nand U26197 (N_26197,N_16749,N_11649);
nand U26198 (N_26198,N_11108,N_18003);
nor U26199 (N_26199,N_11117,N_15640);
and U26200 (N_26200,N_13428,N_11774);
nand U26201 (N_26201,N_17425,N_16445);
nand U26202 (N_26202,N_11356,N_19368);
nand U26203 (N_26203,N_18471,N_10338);
nor U26204 (N_26204,N_19120,N_13598);
nand U26205 (N_26205,N_13213,N_16000);
nor U26206 (N_26206,N_18372,N_18468);
nand U26207 (N_26207,N_10759,N_12759);
xnor U26208 (N_26208,N_12898,N_19329);
or U26209 (N_26209,N_12060,N_10428);
or U26210 (N_26210,N_12814,N_18303);
nor U26211 (N_26211,N_10001,N_11384);
and U26212 (N_26212,N_12612,N_12661);
xor U26213 (N_26213,N_13571,N_18342);
nor U26214 (N_26214,N_12645,N_17678);
xor U26215 (N_26215,N_14595,N_10257);
nand U26216 (N_26216,N_10682,N_10774);
or U26217 (N_26217,N_16381,N_17350);
xnor U26218 (N_26218,N_11316,N_16151);
nor U26219 (N_26219,N_10843,N_16395);
and U26220 (N_26220,N_11936,N_16690);
nor U26221 (N_26221,N_10097,N_11010);
or U26222 (N_26222,N_12486,N_13587);
or U26223 (N_26223,N_18137,N_18540);
xor U26224 (N_26224,N_15673,N_14995);
or U26225 (N_26225,N_19605,N_13865);
and U26226 (N_26226,N_11481,N_14079);
or U26227 (N_26227,N_10298,N_12889);
nand U26228 (N_26228,N_13022,N_11563);
or U26229 (N_26229,N_14427,N_18099);
or U26230 (N_26230,N_10599,N_12205);
and U26231 (N_26231,N_13924,N_13283);
nand U26232 (N_26232,N_10356,N_17101);
nand U26233 (N_26233,N_19894,N_10094);
nor U26234 (N_26234,N_13099,N_13435);
nor U26235 (N_26235,N_11351,N_13073);
and U26236 (N_26236,N_17862,N_19297);
nor U26237 (N_26237,N_17474,N_10566);
nand U26238 (N_26238,N_15393,N_11096);
nand U26239 (N_26239,N_10526,N_18248);
xnor U26240 (N_26240,N_10265,N_10671);
and U26241 (N_26241,N_17170,N_19646);
xor U26242 (N_26242,N_11932,N_16687);
nor U26243 (N_26243,N_17035,N_14478);
or U26244 (N_26244,N_12882,N_17794);
nor U26245 (N_26245,N_11312,N_15595);
or U26246 (N_26246,N_14392,N_15455);
nor U26247 (N_26247,N_10376,N_10591);
nand U26248 (N_26248,N_12532,N_13082);
xor U26249 (N_26249,N_12257,N_16928);
or U26250 (N_26250,N_11548,N_10729);
nand U26251 (N_26251,N_16764,N_19660);
nor U26252 (N_26252,N_18651,N_14464);
or U26253 (N_26253,N_19493,N_19455);
xnor U26254 (N_26254,N_19663,N_19505);
xor U26255 (N_26255,N_16222,N_19604);
or U26256 (N_26256,N_17359,N_10956);
nor U26257 (N_26257,N_11580,N_19427);
and U26258 (N_26258,N_18158,N_15547);
nor U26259 (N_26259,N_10886,N_17906);
and U26260 (N_26260,N_10383,N_18827);
nand U26261 (N_26261,N_19523,N_19400);
or U26262 (N_26262,N_14951,N_17569);
or U26263 (N_26263,N_11664,N_16266);
nor U26264 (N_26264,N_18496,N_17776);
and U26265 (N_26265,N_15239,N_16124);
nor U26266 (N_26266,N_11460,N_10409);
xor U26267 (N_26267,N_17754,N_17135);
and U26268 (N_26268,N_19572,N_18530);
nand U26269 (N_26269,N_10788,N_13905);
nor U26270 (N_26270,N_15567,N_18127);
nand U26271 (N_26271,N_17190,N_11284);
nand U26272 (N_26272,N_15289,N_19322);
nor U26273 (N_26273,N_17550,N_11600);
or U26274 (N_26274,N_17296,N_11245);
nor U26275 (N_26275,N_12592,N_12362);
and U26276 (N_26276,N_11349,N_13563);
or U26277 (N_26277,N_10678,N_15138);
nor U26278 (N_26278,N_18477,N_11626);
nand U26279 (N_26279,N_15440,N_16067);
nor U26280 (N_26280,N_16751,N_18066);
or U26281 (N_26281,N_15658,N_19907);
and U26282 (N_26282,N_10234,N_13848);
nor U26283 (N_26283,N_14188,N_15359);
and U26284 (N_26284,N_10311,N_18591);
xnor U26285 (N_26285,N_12266,N_19643);
and U26286 (N_26286,N_13470,N_18016);
and U26287 (N_26287,N_16234,N_11302);
or U26288 (N_26288,N_16213,N_17510);
or U26289 (N_26289,N_18574,N_15342);
xnor U26290 (N_26290,N_17661,N_14952);
and U26291 (N_26291,N_18732,N_12788);
xnor U26292 (N_26292,N_14151,N_11380);
xor U26293 (N_26293,N_19574,N_14045);
nor U26294 (N_26294,N_19650,N_10426);
nor U26295 (N_26295,N_12531,N_18535);
and U26296 (N_26296,N_17602,N_19306);
nor U26297 (N_26297,N_14047,N_10333);
nand U26298 (N_26298,N_11446,N_17894);
nand U26299 (N_26299,N_10387,N_18423);
or U26300 (N_26300,N_18072,N_13579);
or U26301 (N_26301,N_13817,N_11319);
nand U26302 (N_26302,N_16487,N_17854);
xnor U26303 (N_26303,N_12572,N_17351);
xor U26304 (N_26304,N_18838,N_13067);
nor U26305 (N_26305,N_13657,N_10181);
xnor U26306 (N_26306,N_13098,N_12478);
or U26307 (N_26307,N_15248,N_16367);
nor U26308 (N_26308,N_16167,N_16229);
nand U26309 (N_26309,N_17142,N_12938);
xor U26310 (N_26310,N_10090,N_12361);
and U26311 (N_26311,N_15711,N_13679);
nand U26312 (N_26312,N_16696,N_13534);
nand U26313 (N_26313,N_16226,N_13543);
nor U26314 (N_26314,N_17067,N_17395);
or U26315 (N_26315,N_16871,N_11822);
or U26316 (N_26316,N_16162,N_19586);
and U26317 (N_26317,N_19193,N_14298);
or U26318 (N_26318,N_12911,N_14570);
or U26319 (N_26319,N_17736,N_11849);
xor U26320 (N_26320,N_17245,N_14639);
or U26321 (N_26321,N_14466,N_10060);
or U26322 (N_26322,N_19634,N_18286);
and U26323 (N_26323,N_12384,N_19549);
or U26324 (N_26324,N_16015,N_11307);
nor U26325 (N_26325,N_17962,N_19251);
nand U26326 (N_26326,N_15981,N_14497);
nor U26327 (N_26327,N_12243,N_16491);
nor U26328 (N_26328,N_16712,N_16998);
xnor U26329 (N_26329,N_15133,N_12665);
nor U26330 (N_26330,N_18249,N_17913);
or U26331 (N_26331,N_17959,N_13191);
nor U26332 (N_26332,N_10005,N_18044);
xnor U26333 (N_26333,N_12889,N_12141);
and U26334 (N_26334,N_10251,N_11762);
and U26335 (N_26335,N_12608,N_17644);
and U26336 (N_26336,N_16072,N_11117);
nand U26337 (N_26337,N_18509,N_15371);
or U26338 (N_26338,N_17603,N_12204);
nand U26339 (N_26339,N_17809,N_11518);
and U26340 (N_26340,N_13634,N_19805);
nand U26341 (N_26341,N_16064,N_13289);
nor U26342 (N_26342,N_19412,N_18051);
or U26343 (N_26343,N_17589,N_13106);
or U26344 (N_26344,N_14125,N_13452);
xnor U26345 (N_26345,N_16706,N_16383);
nor U26346 (N_26346,N_18911,N_15769);
and U26347 (N_26347,N_18483,N_12328);
or U26348 (N_26348,N_10930,N_19860);
or U26349 (N_26349,N_12388,N_17790);
and U26350 (N_26350,N_16664,N_15816);
nor U26351 (N_26351,N_13588,N_15365);
and U26352 (N_26352,N_14028,N_11116);
and U26353 (N_26353,N_11483,N_19781);
nand U26354 (N_26354,N_14510,N_17172);
nand U26355 (N_26355,N_14328,N_17908);
nand U26356 (N_26356,N_11645,N_15249);
nand U26357 (N_26357,N_10263,N_19293);
nand U26358 (N_26358,N_17469,N_13498);
nor U26359 (N_26359,N_17435,N_12945);
xnor U26360 (N_26360,N_12542,N_10757);
xor U26361 (N_26361,N_13291,N_10692);
xnor U26362 (N_26362,N_14614,N_19220);
or U26363 (N_26363,N_17727,N_19509);
nor U26364 (N_26364,N_11994,N_10646);
xor U26365 (N_26365,N_17575,N_15331);
and U26366 (N_26366,N_14665,N_17579);
nor U26367 (N_26367,N_16292,N_13007);
nor U26368 (N_26368,N_16044,N_10213);
nor U26369 (N_26369,N_11581,N_14067);
nor U26370 (N_26370,N_15020,N_16267);
nand U26371 (N_26371,N_16905,N_12091);
or U26372 (N_26372,N_12386,N_17152);
and U26373 (N_26373,N_17494,N_11944);
and U26374 (N_26374,N_16085,N_12305);
or U26375 (N_26375,N_18773,N_13344);
or U26376 (N_26376,N_17754,N_17789);
nor U26377 (N_26377,N_13343,N_15788);
xnor U26378 (N_26378,N_10571,N_11753);
xnor U26379 (N_26379,N_19899,N_18009);
nand U26380 (N_26380,N_10173,N_18372);
or U26381 (N_26381,N_14535,N_14404);
xnor U26382 (N_26382,N_12030,N_11853);
xnor U26383 (N_26383,N_17749,N_18610);
xor U26384 (N_26384,N_16418,N_17005);
nor U26385 (N_26385,N_12220,N_13263);
or U26386 (N_26386,N_12645,N_12508);
nor U26387 (N_26387,N_10780,N_18585);
nand U26388 (N_26388,N_12870,N_16166);
or U26389 (N_26389,N_11098,N_11017);
nand U26390 (N_26390,N_14204,N_17048);
or U26391 (N_26391,N_12865,N_16939);
nor U26392 (N_26392,N_18174,N_18669);
nand U26393 (N_26393,N_10888,N_12797);
and U26394 (N_26394,N_11881,N_12441);
nand U26395 (N_26395,N_10507,N_12550);
or U26396 (N_26396,N_13510,N_16949);
or U26397 (N_26397,N_13690,N_13534);
nand U26398 (N_26398,N_14946,N_16210);
or U26399 (N_26399,N_10103,N_13362);
and U26400 (N_26400,N_12152,N_10218);
or U26401 (N_26401,N_18708,N_14660);
nand U26402 (N_26402,N_13499,N_16263);
xnor U26403 (N_26403,N_14618,N_18482);
nand U26404 (N_26404,N_12056,N_15852);
nand U26405 (N_26405,N_18118,N_11569);
nor U26406 (N_26406,N_12539,N_18430);
xnor U26407 (N_26407,N_13974,N_18115);
or U26408 (N_26408,N_19607,N_11788);
or U26409 (N_26409,N_18670,N_17677);
or U26410 (N_26410,N_10392,N_18729);
nor U26411 (N_26411,N_10570,N_18609);
nand U26412 (N_26412,N_12579,N_13967);
nor U26413 (N_26413,N_13047,N_17012);
nor U26414 (N_26414,N_18510,N_17757);
nand U26415 (N_26415,N_11111,N_19203);
nand U26416 (N_26416,N_16968,N_15248);
xor U26417 (N_26417,N_15604,N_12762);
and U26418 (N_26418,N_18707,N_11907);
nand U26419 (N_26419,N_18665,N_14108);
nand U26420 (N_26420,N_15315,N_16319);
or U26421 (N_26421,N_18914,N_14934);
nand U26422 (N_26422,N_12837,N_19135);
nor U26423 (N_26423,N_15088,N_15834);
nor U26424 (N_26424,N_18947,N_16094);
xnor U26425 (N_26425,N_16222,N_18645);
and U26426 (N_26426,N_12042,N_14372);
xnor U26427 (N_26427,N_18450,N_14716);
or U26428 (N_26428,N_14396,N_17383);
xor U26429 (N_26429,N_19305,N_19568);
nor U26430 (N_26430,N_13673,N_15413);
nor U26431 (N_26431,N_10542,N_18731);
nor U26432 (N_26432,N_17432,N_16077);
or U26433 (N_26433,N_10377,N_17333);
nand U26434 (N_26434,N_10513,N_19045);
nand U26435 (N_26435,N_16803,N_18964);
or U26436 (N_26436,N_13565,N_19693);
nor U26437 (N_26437,N_16168,N_12908);
nor U26438 (N_26438,N_14557,N_19095);
nor U26439 (N_26439,N_11917,N_12729);
nor U26440 (N_26440,N_12859,N_14200);
xnor U26441 (N_26441,N_15523,N_18397);
nand U26442 (N_26442,N_17370,N_17421);
nor U26443 (N_26443,N_14656,N_16236);
nor U26444 (N_26444,N_12342,N_18855);
xnor U26445 (N_26445,N_15109,N_11853);
nand U26446 (N_26446,N_13812,N_19083);
and U26447 (N_26447,N_13071,N_12624);
nor U26448 (N_26448,N_10585,N_15122);
and U26449 (N_26449,N_11456,N_17763);
xnor U26450 (N_26450,N_12157,N_16498);
xnor U26451 (N_26451,N_13046,N_11556);
and U26452 (N_26452,N_16737,N_13607);
or U26453 (N_26453,N_15047,N_18783);
or U26454 (N_26454,N_18097,N_18103);
nand U26455 (N_26455,N_15503,N_17872);
nand U26456 (N_26456,N_16738,N_16959);
or U26457 (N_26457,N_18827,N_16375);
nand U26458 (N_26458,N_11104,N_16741);
xor U26459 (N_26459,N_13635,N_18957);
nor U26460 (N_26460,N_13871,N_16687);
and U26461 (N_26461,N_18876,N_12526);
nand U26462 (N_26462,N_17989,N_14822);
nand U26463 (N_26463,N_13678,N_19338);
xor U26464 (N_26464,N_17300,N_18377);
or U26465 (N_26465,N_10118,N_17976);
and U26466 (N_26466,N_18878,N_10428);
nor U26467 (N_26467,N_15243,N_12588);
nand U26468 (N_26468,N_10682,N_17289);
xnor U26469 (N_26469,N_15134,N_17265);
xnor U26470 (N_26470,N_10102,N_11056);
or U26471 (N_26471,N_14445,N_14133);
and U26472 (N_26472,N_17832,N_14901);
nand U26473 (N_26473,N_12593,N_13030);
and U26474 (N_26474,N_19728,N_13149);
xor U26475 (N_26475,N_13451,N_16584);
or U26476 (N_26476,N_17045,N_18198);
xor U26477 (N_26477,N_17944,N_13879);
or U26478 (N_26478,N_14457,N_11921);
and U26479 (N_26479,N_13707,N_13426);
or U26480 (N_26480,N_16335,N_13363);
or U26481 (N_26481,N_17586,N_11392);
nand U26482 (N_26482,N_14685,N_13663);
nor U26483 (N_26483,N_16440,N_18928);
nand U26484 (N_26484,N_12802,N_11941);
nand U26485 (N_26485,N_19102,N_11422);
or U26486 (N_26486,N_12106,N_19168);
and U26487 (N_26487,N_17552,N_15749);
xnor U26488 (N_26488,N_18782,N_19035);
or U26489 (N_26489,N_11842,N_18739);
nor U26490 (N_26490,N_14222,N_18207);
xnor U26491 (N_26491,N_19692,N_12721);
and U26492 (N_26492,N_11634,N_15808);
and U26493 (N_26493,N_10272,N_14584);
or U26494 (N_26494,N_12065,N_16154);
xnor U26495 (N_26495,N_14094,N_11009);
or U26496 (N_26496,N_11622,N_15783);
xnor U26497 (N_26497,N_18523,N_19646);
nand U26498 (N_26498,N_14234,N_15356);
or U26499 (N_26499,N_10500,N_10713);
nor U26500 (N_26500,N_13839,N_16383);
nand U26501 (N_26501,N_10389,N_11414);
nand U26502 (N_26502,N_16847,N_11115);
xor U26503 (N_26503,N_14788,N_16822);
nand U26504 (N_26504,N_12923,N_12136);
xnor U26505 (N_26505,N_10901,N_16215);
nand U26506 (N_26506,N_11082,N_12421);
or U26507 (N_26507,N_11570,N_16208);
and U26508 (N_26508,N_17112,N_17817);
xnor U26509 (N_26509,N_14777,N_18747);
nand U26510 (N_26510,N_18879,N_10370);
and U26511 (N_26511,N_17501,N_13048);
xor U26512 (N_26512,N_12099,N_13943);
xnor U26513 (N_26513,N_14320,N_16721);
xor U26514 (N_26514,N_11925,N_19522);
xor U26515 (N_26515,N_14243,N_16433);
xnor U26516 (N_26516,N_18463,N_14230);
and U26517 (N_26517,N_14535,N_10803);
xor U26518 (N_26518,N_11922,N_15585);
xnor U26519 (N_26519,N_11976,N_19290);
and U26520 (N_26520,N_19444,N_19546);
xor U26521 (N_26521,N_10783,N_12330);
and U26522 (N_26522,N_12049,N_11678);
nand U26523 (N_26523,N_15616,N_15503);
nor U26524 (N_26524,N_18567,N_17096);
nand U26525 (N_26525,N_13796,N_12951);
or U26526 (N_26526,N_16513,N_17245);
xor U26527 (N_26527,N_15299,N_12249);
nand U26528 (N_26528,N_11730,N_16071);
or U26529 (N_26529,N_16176,N_16898);
xnor U26530 (N_26530,N_15667,N_14521);
or U26531 (N_26531,N_18155,N_15099);
nand U26532 (N_26532,N_12066,N_14609);
xnor U26533 (N_26533,N_10333,N_10799);
or U26534 (N_26534,N_16528,N_13314);
nand U26535 (N_26535,N_18400,N_14446);
xor U26536 (N_26536,N_15202,N_14771);
and U26537 (N_26537,N_11868,N_17948);
or U26538 (N_26538,N_11915,N_11753);
xnor U26539 (N_26539,N_17578,N_12480);
nand U26540 (N_26540,N_18917,N_17921);
or U26541 (N_26541,N_17943,N_12273);
and U26542 (N_26542,N_14674,N_19815);
or U26543 (N_26543,N_13137,N_11928);
nand U26544 (N_26544,N_16637,N_11992);
nand U26545 (N_26545,N_10824,N_17198);
nand U26546 (N_26546,N_14706,N_18893);
nand U26547 (N_26547,N_15964,N_14102);
nor U26548 (N_26548,N_19890,N_10709);
nor U26549 (N_26549,N_13866,N_12582);
and U26550 (N_26550,N_12207,N_19563);
and U26551 (N_26551,N_13305,N_11978);
or U26552 (N_26552,N_19701,N_15073);
nand U26553 (N_26553,N_15772,N_16593);
and U26554 (N_26554,N_15186,N_16673);
xnor U26555 (N_26555,N_18518,N_13315);
and U26556 (N_26556,N_13896,N_12130);
nor U26557 (N_26557,N_18264,N_12532);
and U26558 (N_26558,N_16975,N_19343);
xnor U26559 (N_26559,N_11447,N_10813);
or U26560 (N_26560,N_18029,N_10458);
and U26561 (N_26561,N_11100,N_15916);
or U26562 (N_26562,N_11853,N_19331);
xnor U26563 (N_26563,N_13269,N_13280);
nand U26564 (N_26564,N_15989,N_12394);
xor U26565 (N_26565,N_12904,N_19526);
and U26566 (N_26566,N_18757,N_14322);
nand U26567 (N_26567,N_16625,N_13418);
or U26568 (N_26568,N_10763,N_13204);
nor U26569 (N_26569,N_17245,N_16542);
and U26570 (N_26570,N_11786,N_10004);
or U26571 (N_26571,N_12055,N_13712);
or U26572 (N_26572,N_12694,N_12114);
nor U26573 (N_26573,N_14077,N_12746);
or U26574 (N_26574,N_15737,N_18263);
nand U26575 (N_26575,N_15509,N_19063);
and U26576 (N_26576,N_19455,N_10691);
nand U26577 (N_26577,N_15791,N_16911);
and U26578 (N_26578,N_14278,N_17855);
nor U26579 (N_26579,N_19981,N_16603);
nor U26580 (N_26580,N_19290,N_18285);
and U26581 (N_26581,N_12442,N_12668);
and U26582 (N_26582,N_18389,N_18776);
nand U26583 (N_26583,N_13979,N_14115);
or U26584 (N_26584,N_14410,N_14705);
xor U26585 (N_26585,N_12127,N_11853);
and U26586 (N_26586,N_13011,N_17510);
or U26587 (N_26587,N_10663,N_16343);
or U26588 (N_26588,N_13531,N_16156);
xor U26589 (N_26589,N_16761,N_16632);
xnor U26590 (N_26590,N_19478,N_12542);
nand U26591 (N_26591,N_11201,N_18671);
nand U26592 (N_26592,N_12336,N_19061);
and U26593 (N_26593,N_10559,N_14756);
and U26594 (N_26594,N_15520,N_16450);
nor U26595 (N_26595,N_15950,N_14637);
xor U26596 (N_26596,N_19603,N_19103);
or U26597 (N_26597,N_19086,N_10396);
nor U26598 (N_26598,N_13366,N_19952);
nand U26599 (N_26599,N_15774,N_14295);
xor U26600 (N_26600,N_19634,N_18193);
xnor U26601 (N_26601,N_10158,N_19166);
and U26602 (N_26602,N_12765,N_19031);
or U26603 (N_26603,N_14241,N_15357);
nor U26604 (N_26604,N_14931,N_11539);
nand U26605 (N_26605,N_13737,N_10004);
xnor U26606 (N_26606,N_12295,N_15582);
xnor U26607 (N_26607,N_15400,N_10597);
xor U26608 (N_26608,N_16215,N_14172);
or U26609 (N_26609,N_17047,N_17632);
or U26610 (N_26610,N_11770,N_11958);
nor U26611 (N_26611,N_16423,N_10677);
and U26612 (N_26612,N_15476,N_15413);
nand U26613 (N_26613,N_10391,N_10518);
and U26614 (N_26614,N_17565,N_18925);
nor U26615 (N_26615,N_19058,N_10501);
nand U26616 (N_26616,N_15485,N_12028);
nor U26617 (N_26617,N_16110,N_19071);
nand U26618 (N_26618,N_11199,N_15507);
xnor U26619 (N_26619,N_16731,N_11795);
and U26620 (N_26620,N_17770,N_14370);
nor U26621 (N_26621,N_18587,N_13929);
xnor U26622 (N_26622,N_18543,N_17949);
nand U26623 (N_26623,N_16834,N_11931);
xor U26624 (N_26624,N_17381,N_14711);
xor U26625 (N_26625,N_19284,N_10924);
xnor U26626 (N_26626,N_10640,N_17108);
and U26627 (N_26627,N_16522,N_17730);
and U26628 (N_26628,N_17694,N_15939);
nand U26629 (N_26629,N_16495,N_18594);
nand U26630 (N_26630,N_16863,N_10125);
xnor U26631 (N_26631,N_17418,N_18839);
nand U26632 (N_26632,N_18319,N_11610);
and U26633 (N_26633,N_10030,N_11546);
nand U26634 (N_26634,N_11460,N_17770);
nor U26635 (N_26635,N_19400,N_15789);
or U26636 (N_26636,N_17587,N_19018);
nor U26637 (N_26637,N_15097,N_16461);
xnor U26638 (N_26638,N_13048,N_15000);
nor U26639 (N_26639,N_10469,N_10803);
or U26640 (N_26640,N_17970,N_16357);
xnor U26641 (N_26641,N_13054,N_19543);
nand U26642 (N_26642,N_11832,N_11054);
and U26643 (N_26643,N_15106,N_18540);
or U26644 (N_26644,N_15501,N_17042);
nand U26645 (N_26645,N_17876,N_14354);
xnor U26646 (N_26646,N_16690,N_15509);
nand U26647 (N_26647,N_16555,N_10884);
or U26648 (N_26648,N_10251,N_17880);
nand U26649 (N_26649,N_19801,N_10391);
nand U26650 (N_26650,N_16195,N_19048);
xor U26651 (N_26651,N_10937,N_11815);
nand U26652 (N_26652,N_15787,N_16401);
xor U26653 (N_26653,N_12371,N_16733);
or U26654 (N_26654,N_15847,N_11613);
nor U26655 (N_26655,N_11191,N_13880);
or U26656 (N_26656,N_19752,N_15026);
nand U26657 (N_26657,N_14020,N_14536);
xor U26658 (N_26658,N_12829,N_16502);
or U26659 (N_26659,N_16108,N_13696);
nor U26660 (N_26660,N_18609,N_16628);
and U26661 (N_26661,N_12218,N_17417);
nand U26662 (N_26662,N_18916,N_12528);
nand U26663 (N_26663,N_17034,N_16669);
nor U26664 (N_26664,N_12742,N_13614);
xor U26665 (N_26665,N_14083,N_13091);
nor U26666 (N_26666,N_19565,N_18566);
xnor U26667 (N_26667,N_14289,N_14436);
or U26668 (N_26668,N_12298,N_13060);
nand U26669 (N_26669,N_17154,N_16847);
nand U26670 (N_26670,N_14867,N_12996);
or U26671 (N_26671,N_10381,N_15256);
or U26672 (N_26672,N_19227,N_10148);
or U26673 (N_26673,N_15278,N_18991);
or U26674 (N_26674,N_10958,N_13741);
or U26675 (N_26675,N_12190,N_15281);
or U26676 (N_26676,N_13610,N_17911);
nor U26677 (N_26677,N_14593,N_10702);
or U26678 (N_26678,N_14336,N_12369);
or U26679 (N_26679,N_16302,N_19371);
nor U26680 (N_26680,N_12340,N_19870);
or U26681 (N_26681,N_18918,N_16127);
and U26682 (N_26682,N_18343,N_16831);
or U26683 (N_26683,N_16270,N_10921);
xnor U26684 (N_26684,N_16018,N_17574);
and U26685 (N_26685,N_12594,N_10978);
or U26686 (N_26686,N_13429,N_14746);
nand U26687 (N_26687,N_11708,N_14585);
nor U26688 (N_26688,N_12903,N_10602);
and U26689 (N_26689,N_17417,N_13735);
nor U26690 (N_26690,N_13282,N_12374);
nor U26691 (N_26691,N_16577,N_12063);
or U26692 (N_26692,N_14309,N_15539);
nor U26693 (N_26693,N_13830,N_13605);
and U26694 (N_26694,N_10688,N_18260);
nor U26695 (N_26695,N_12777,N_10595);
and U26696 (N_26696,N_13571,N_17276);
xnor U26697 (N_26697,N_19324,N_14586);
xnor U26698 (N_26698,N_10403,N_11922);
nand U26699 (N_26699,N_18346,N_14143);
or U26700 (N_26700,N_19690,N_19844);
nor U26701 (N_26701,N_10767,N_17976);
xor U26702 (N_26702,N_11665,N_14207);
xor U26703 (N_26703,N_18399,N_19314);
or U26704 (N_26704,N_11389,N_10371);
and U26705 (N_26705,N_15608,N_13562);
xor U26706 (N_26706,N_13428,N_19847);
and U26707 (N_26707,N_10634,N_12642);
or U26708 (N_26708,N_12786,N_11417);
and U26709 (N_26709,N_19013,N_15079);
and U26710 (N_26710,N_10861,N_16606);
and U26711 (N_26711,N_16371,N_19048);
nand U26712 (N_26712,N_12866,N_12945);
nand U26713 (N_26713,N_10125,N_11819);
xnor U26714 (N_26714,N_18213,N_11506);
xor U26715 (N_26715,N_18142,N_18856);
nand U26716 (N_26716,N_13654,N_19071);
and U26717 (N_26717,N_17603,N_10630);
and U26718 (N_26718,N_17444,N_13598);
nor U26719 (N_26719,N_13284,N_12231);
or U26720 (N_26720,N_19294,N_19540);
xor U26721 (N_26721,N_16591,N_13433);
xnor U26722 (N_26722,N_13703,N_11015);
or U26723 (N_26723,N_11948,N_11935);
nand U26724 (N_26724,N_18686,N_13747);
nor U26725 (N_26725,N_18095,N_11633);
and U26726 (N_26726,N_19044,N_12768);
xor U26727 (N_26727,N_12691,N_13948);
nor U26728 (N_26728,N_11692,N_11643);
xnor U26729 (N_26729,N_12023,N_19549);
nor U26730 (N_26730,N_13974,N_14484);
or U26731 (N_26731,N_13410,N_11528);
nor U26732 (N_26732,N_13366,N_18067);
nor U26733 (N_26733,N_18885,N_13679);
nor U26734 (N_26734,N_11437,N_10900);
xnor U26735 (N_26735,N_12414,N_10400);
xnor U26736 (N_26736,N_16443,N_18859);
and U26737 (N_26737,N_16420,N_16227);
nor U26738 (N_26738,N_13764,N_19582);
xnor U26739 (N_26739,N_19175,N_14166);
and U26740 (N_26740,N_17565,N_13287);
and U26741 (N_26741,N_19379,N_15754);
and U26742 (N_26742,N_18462,N_14975);
or U26743 (N_26743,N_14791,N_17024);
and U26744 (N_26744,N_11972,N_19839);
and U26745 (N_26745,N_19686,N_15214);
and U26746 (N_26746,N_14413,N_14553);
and U26747 (N_26747,N_14562,N_10171);
xor U26748 (N_26748,N_15312,N_16721);
nand U26749 (N_26749,N_17936,N_11442);
xnor U26750 (N_26750,N_14114,N_13871);
nand U26751 (N_26751,N_11945,N_17325);
xor U26752 (N_26752,N_11647,N_17492);
and U26753 (N_26753,N_15379,N_19004);
or U26754 (N_26754,N_12344,N_13328);
or U26755 (N_26755,N_16074,N_15094);
xor U26756 (N_26756,N_19105,N_16356);
or U26757 (N_26757,N_19420,N_19553);
nand U26758 (N_26758,N_18758,N_14121);
nand U26759 (N_26759,N_13000,N_11908);
nand U26760 (N_26760,N_12698,N_14901);
and U26761 (N_26761,N_15492,N_11520);
nand U26762 (N_26762,N_11518,N_18521);
or U26763 (N_26763,N_19100,N_13840);
nand U26764 (N_26764,N_19735,N_19191);
or U26765 (N_26765,N_14845,N_16495);
and U26766 (N_26766,N_17653,N_13838);
nor U26767 (N_26767,N_18251,N_19375);
xor U26768 (N_26768,N_16777,N_18688);
and U26769 (N_26769,N_15369,N_11386);
and U26770 (N_26770,N_15306,N_10205);
or U26771 (N_26771,N_19934,N_19850);
and U26772 (N_26772,N_10530,N_10075);
or U26773 (N_26773,N_16028,N_19772);
nand U26774 (N_26774,N_18961,N_13269);
or U26775 (N_26775,N_11480,N_14873);
nor U26776 (N_26776,N_19963,N_11665);
xor U26777 (N_26777,N_16214,N_12348);
or U26778 (N_26778,N_16162,N_16045);
nor U26779 (N_26779,N_15271,N_13452);
nor U26780 (N_26780,N_11431,N_10662);
or U26781 (N_26781,N_16481,N_14763);
nand U26782 (N_26782,N_11596,N_10668);
or U26783 (N_26783,N_15084,N_14305);
or U26784 (N_26784,N_11484,N_13998);
and U26785 (N_26785,N_11182,N_15882);
nand U26786 (N_26786,N_16844,N_11789);
xor U26787 (N_26787,N_16293,N_16208);
or U26788 (N_26788,N_12374,N_19124);
xnor U26789 (N_26789,N_12085,N_18239);
or U26790 (N_26790,N_16886,N_17629);
and U26791 (N_26791,N_11907,N_11209);
nor U26792 (N_26792,N_11246,N_15522);
nand U26793 (N_26793,N_16039,N_19960);
nor U26794 (N_26794,N_12989,N_10432);
or U26795 (N_26795,N_16657,N_19264);
or U26796 (N_26796,N_15985,N_12736);
xnor U26797 (N_26797,N_18552,N_14727);
nor U26798 (N_26798,N_15998,N_16025);
nor U26799 (N_26799,N_15688,N_15638);
xnor U26800 (N_26800,N_12472,N_15415);
xnor U26801 (N_26801,N_13190,N_12171);
or U26802 (N_26802,N_17748,N_19285);
and U26803 (N_26803,N_18591,N_17074);
nor U26804 (N_26804,N_17723,N_19119);
xor U26805 (N_26805,N_14221,N_19046);
and U26806 (N_26806,N_13876,N_19618);
or U26807 (N_26807,N_19383,N_18505);
xor U26808 (N_26808,N_15649,N_14689);
nand U26809 (N_26809,N_12498,N_17515);
or U26810 (N_26810,N_19839,N_19619);
nand U26811 (N_26811,N_14010,N_16364);
xor U26812 (N_26812,N_10195,N_17026);
xor U26813 (N_26813,N_11360,N_11788);
or U26814 (N_26814,N_13721,N_19704);
and U26815 (N_26815,N_18407,N_17302);
nor U26816 (N_26816,N_11232,N_18553);
or U26817 (N_26817,N_10346,N_14825);
xor U26818 (N_26818,N_15670,N_12660);
xor U26819 (N_26819,N_11076,N_11326);
nand U26820 (N_26820,N_10404,N_18970);
xnor U26821 (N_26821,N_18170,N_15298);
and U26822 (N_26822,N_19944,N_12117);
xnor U26823 (N_26823,N_16618,N_19415);
or U26824 (N_26824,N_16990,N_12735);
or U26825 (N_26825,N_11778,N_14000);
nor U26826 (N_26826,N_15085,N_19653);
and U26827 (N_26827,N_17422,N_15723);
nand U26828 (N_26828,N_17362,N_13601);
xor U26829 (N_26829,N_14767,N_10205);
xor U26830 (N_26830,N_15468,N_19377);
nor U26831 (N_26831,N_19433,N_12655);
nor U26832 (N_26832,N_18692,N_11030);
nand U26833 (N_26833,N_12343,N_10601);
xnor U26834 (N_26834,N_17623,N_15131);
or U26835 (N_26835,N_12695,N_18712);
or U26836 (N_26836,N_14520,N_12827);
nor U26837 (N_26837,N_13185,N_10410);
or U26838 (N_26838,N_15622,N_18059);
xnor U26839 (N_26839,N_10720,N_12679);
xor U26840 (N_26840,N_17329,N_16092);
or U26841 (N_26841,N_11975,N_12047);
xor U26842 (N_26842,N_11996,N_12196);
nand U26843 (N_26843,N_14476,N_11290);
nand U26844 (N_26844,N_14010,N_19612);
nor U26845 (N_26845,N_15685,N_15503);
nor U26846 (N_26846,N_19253,N_18953);
and U26847 (N_26847,N_18774,N_12303);
nand U26848 (N_26848,N_15278,N_17474);
or U26849 (N_26849,N_16965,N_15683);
nor U26850 (N_26850,N_13793,N_13949);
nor U26851 (N_26851,N_13519,N_11260);
or U26852 (N_26852,N_14041,N_15263);
nor U26853 (N_26853,N_13853,N_16297);
xor U26854 (N_26854,N_18841,N_19263);
xor U26855 (N_26855,N_15439,N_19724);
nand U26856 (N_26856,N_13525,N_19465);
nor U26857 (N_26857,N_14430,N_18017);
or U26858 (N_26858,N_13742,N_14597);
and U26859 (N_26859,N_11684,N_19507);
nand U26860 (N_26860,N_13471,N_14239);
nor U26861 (N_26861,N_17545,N_17009);
and U26862 (N_26862,N_16931,N_14026);
xnor U26863 (N_26863,N_13164,N_14628);
nand U26864 (N_26864,N_12422,N_14468);
or U26865 (N_26865,N_12241,N_17306);
or U26866 (N_26866,N_10497,N_16654);
nand U26867 (N_26867,N_18843,N_18015);
nor U26868 (N_26868,N_15404,N_10882);
or U26869 (N_26869,N_16087,N_17141);
nand U26870 (N_26870,N_13384,N_17872);
and U26871 (N_26871,N_18855,N_17911);
or U26872 (N_26872,N_19462,N_12329);
nand U26873 (N_26873,N_13920,N_16953);
nor U26874 (N_26874,N_18240,N_12677);
xnor U26875 (N_26875,N_19645,N_10557);
xnor U26876 (N_26876,N_10093,N_14935);
nor U26877 (N_26877,N_16063,N_17078);
or U26878 (N_26878,N_14605,N_10835);
nand U26879 (N_26879,N_15933,N_18911);
nor U26880 (N_26880,N_19973,N_15589);
and U26881 (N_26881,N_14002,N_12962);
xnor U26882 (N_26882,N_14223,N_15282);
or U26883 (N_26883,N_17082,N_17069);
or U26884 (N_26884,N_13986,N_10793);
and U26885 (N_26885,N_15324,N_16901);
and U26886 (N_26886,N_18188,N_12529);
xor U26887 (N_26887,N_16664,N_14570);
xor U26888 (N_26888,N_12040,N_13524);
nand U26889 (N_26889,N_10585,N_17205);
nor U26890 (N_26890,N_19587,N_15586);
or U26891 (N_26891,N_10199,N_15039);
and U26892 (N_26892,N_12802,N_12173);
and U26893 (N_26893,N_14016,N_18093);
nand U26894 (N_26894,N_12169,N_14272);
nand U26895 (N_26895,N_16394,N_17751);
xor U26896 (N_26896,N_16223,N_18188);
or U26897 (N_26897,N_17237,N_11134);
xor U26898 (N_26898,N_14941,N_13102);
or U26899 (N_26899,N_10046,N_13094);
nand U26900 (N_26900,N_18372,N_18088);
nand U26901 (N_26901,N_17247,N_16126);
xnor U26902 (N_26902,N_10841,N_14094);
and U26903 (N_26903,N_19629,N_10968);
nand U26904 (N_26904,N_11968,N_15688);
nand U26905 (N_26905,N_17388,N_15639);
nor U26906 (N_26906,N_11427,N_11270);
xor U26907 (N_26907,N_10456,N_10453);
xor U26908 (N_26908,N_10476,N_14045);
nand U26909 (N_26909,N_12635,N_11092);
nand U26910 (N_26910,N_15501,N_15410);
nand U26911 (N_26911,N_17672,N_17609);
and U26912 (N_26912,N_12479,N_11564);
nand U26913 (N_26913,N_12230,N_10232);
xnor U26914 (N_26914,N_16343,N_11352);
nor U26915 (N_26915,N_16561,N_12627);
and U26916 (N_26916,N_13993,N_15889);
or U26917 (N_26917,N_13715,N_13854);
and U26918 (N_26918,N_18691,N_18622);
xnor U26919 (N_26919,N_15936,N_10093);
xor U26920 (N_26920,N_12229,N_11264);
nand U26921 (N_26921,N_16138,N_19936);
xor U26922 (N_26922,N_14164,N_18697);
xnor U26923 (N_26923,N_13450,N_18009);
nor U26924 (N_26924,N_16731,N_17855);
nand U26925 (N_26925,N_10317,N_16320);
nand U26926 (N_26926,N_17886,N_10598);
nand U26927 (N_26927,N_14457,N_11487);
and U26928 (N_26928,N_17284,N_19274);
nand U26929 (N_26929,N_18898,N_17508);
and U26930 (N_26930,N_11305,N_13590);
nor U26931 (N_26931,N_15994,N_11295);
nand U26932 (N_26932,N_17184,N_10681);
nand U26933 (N_26933,N_10560,N_16476);
nand U26934 (N_26934,N_12328,N_16680);
or U26935 (N_26935,N_19279,N_16960);
nand U26936 (N_26936,N_17243,N_17946);
or U26937 (N_26937,N_13045,N_19519);
and U26938 (N_26938,N_18107,N_12498);
nand U26939 (N_26939,N_15118,N_13537);
and U26940 (N_26940,N_12304,N_18293);
nand U26941 (N_26941,N_17370,N_18667);
or U26942 (N_26942,N_13410,N_19523);
nand U26943 (N_26943,N_13604,N_14638);
nor U26944 (N_26944,N_18137,N_11292);
xnor U26945 (N_26945,N_16190,N_18651);
or U26946 (N_26946,N_16172,N_11958);
or U26947 (N_26947,N_14097,N_14115);
nand U26948 (N_26948,N_14557,N_13616);
and U26949 (N_26949,N_15230,N_16607);
nand U26950 (N_26950,N_13603,N_19212);
and U26951 (N_26951,N_16761,N_12731);
xnor U26952 (N_26952,N_15208,N_13740);
and U26953 (N_26953,N_19861,N_16421);
xnor U26954 (N_26954,N_17210,N_19400);
xor U26955 (N_26955,N_16499,N_18973);
nand U26956 (N_26956,N_17766,N_15629);
or U26957 (N_26957,N_16074,N_12321);
and U26958 (N_26958,N_18855,N_13545);
and U26959 (N_26959,N_17922,N_10480);
nor U26960 (N_26960,N_12857,N_13690);
xor U26961 (N_26961,N_14080,N_18521);
or U26962 (N_26962,N_18138,N_19200);
nor U26963 (N_26963,N_16627,N_18784);
or U26964 (N_26964,N_14700,N_15480);
xnor U26965 (N_26965,N_19795,N_15008);
or U26966 (N_26966,N_19144,N_10631);
xor U26967 (N_26967,N_12830,N_15269);
and U26968 (N_26968,N_18463,N_13354);
and U26969 (N_26969,N_14362,N_17315);
xor U26970 (N_26970,N_13015,N_14295);
or U26971 (N_26971,N_10535,N_19325);
nand U26972 (N_26972,N_15664,N_14815);
or U26973 (N_26973,N_17551,N_15487);
nor U26974 (N_26974,N_14170,N_15901);
nand U26975 (N_26975,N_19511,N_19293);
nor U26976 (N_26976,N_14948,N_13823);
or U26977 (N_26977,N_12486,N_17622);
or U26978 (N_26978,N_13660,N_11681);
nor U26979 (N_26979,N_13080,N_17486);
and U26980 (N_26980,N_15560,N_10395);
nand U26981 (N_26981,N_14641,N_13182);
xnor U26982 (N_26982,N_15958,N_18001);
xnor U26983 (N_26983,N_11241,N_15139);
or U26984 (N_26984,N_15286,N_19006);
and U26985 (N_26985,N_15212,N_11578);
nand U26986 (N_26986,N_11451,N_11706);
nand U26987 (N_26987,N_16533,N_19186);
nand U26988 (N_26988,N_10635,N_15474);
nand U26989 (N_26989,N_16406,N_18398);
nor U26990 (N_26990,N_18314,N_14982);
nor U26991 (N_26991,N_18789,N_19688);
and U26992 (N_26992,N_15756,N_17310);
nand U26993 (N_26993,N_14833,N_17511);
xnor U26994 (N_26994,N_18865,N_10107);
nor U26995 (N_26995,N_13765,N_18909);
xor U26996 (N_26996,N_19037,N_16345);
nor U26997 (N_26997,N_17477,N_17558);
xor U26998 (N_26998,N_15337,N_12420);
nor U26999 (N_26999,N_18898,N_17723);
nor U27000 (N_27000,N_14925,N_10261);
xnor U27001 (N_27001,N_19903,N_10450);
xnor U27002 (N_27002,N_18182,N_18048);
and U27003 (N_27003,N_14947,N_16757);
nand U27004 (N_27004,N_17862,N_19455);
nor U27005 (N_27005,N_11252,N_13158);
and U27006 (N_27006,N_18469,N_15373);
and U27007 (N_27007,N_18840,N_16151);
xnor U27008 (N_27008,N_10429,N_10781);
and U27009 (N_27009,N_16379,N_15132);
xnor U27010 (N_27010,N_17967,N_12522);
nor U27011 (N_27011,N_11452,N_16704);
xor U27012 (N_27012,N_11663,N_12769);
xor U27013 (N_27013,N_17318,N_14296);
or U27014 (N_27014,N_10047,N_16884);
or U27015 (N_27015,N_10310,N_13638);
nor U27016 (N_27016,N_18127,N_19321);
or U27017 (N_27017,N_13797,N_15157);
xor U27018 (N_27018,N_14863,N_19140);
or U27019 (N_27019,N_10251,N_11524);
or U27020 (N_27020,N_11547,N_16604);
nor U27021 (N_27021,N_17066,N_13807);
or U27022 (N_27022,N_11811,N_16160);
and U27023 (N_27023,N_15710,N_11920);
nor U27024 (N_27024,N_19605,N_14975);
and U27025 (N_27025,N_12930,N_14301);
and U27026 (N_27026,N_11305,N_13800);
xor U27027 (N_27027,N_18399,N_17031);
nor U27028 (N_27028,N_13853,N_16010);
and U27029 (N_27029,N_11499,N_14765);
nand U27030 (N_27030,N_19202,N_19035);
xor U27031 (N_27031,N_16178,N_18773);
and U27032 (N_27032,N_10432,N_16174);
and U27033 (N_27033,N_11476,N_11490);
nand U27034 (N_27034,N_17505,N_12526);
or U27035 (N_27035,N_19235,N_10646);
xnor U27036 (N_27036,N_19357,N_18215);
nand U27037 (N_27037,N_16944,N_14991);
or U27038 (N_27038,N_12263,N_19943);
and U27039 (N_27039,N_13662,N_18440);
nand U27040 (N_27040,N_11174,N_14719);
and U27041 (N_27041,N_14876,N_13276);
and U27042 (N_27042,N_14911,N_14154);
and U27043 (N_27043,N_18388,N_16391);
nor U27044 (N_27044,N_19481,N_19131);
or U27045 (N_27045,N_15535,N_10237);
nand U27046 (N_27046,N_19391,N_14436);
nor U27047 (N_27047,N_10501,N_12712);
and U27048 (N_27048,N_18345,N_13035);
and U27049 (N_27049,N_16226,N_17846);
nand U27050 (N_27050,N_18267,N_13727);
or U27051 (N_27051,N_13247,N_14496);
nor U27052 (N_27052,N_11741,N_12271);
xnor U27053 (N_27053,N_11357,N_14153);
xor U27054 (N_27054,N_14574,N_17053);
and U27055 (N_27055,N_13960,N_11138);
or U27056 (N_27056,N_15849,N_19362);
nor U27057 (N_27057,N_17209,N_13308);
and U27058 (N_27058,N_18574,N_19694);
xnor U27059 (N_27059,N_11101,N_19648);
and U27060 (N_27060,N_13387,N_11330);
nor U27061 (N_27061,N_15352,N_13207);
xor U27062 (N_27062,N_13624,N_19056);
nor U27063 (N_27063,N_19926,N_11466);
or U27064 (N_27064,N_16021,N_10379);
xnor U27065 (N_27065,N_10898,N_17125);
xnor U27066 (N_27066,N_19116,N_15303);
or U27067 (N_27067,N_19255,N_18732);
and U27068 (N_27068,N_18482,N_17707);
xor U27069 (N_27069,N_12712,N_14542);
xor U27070 (N_27070,N_18232,N_15745);
or U27071 (N_27071,N_17750,N_11612);
nand U27072 (N_27072,N_11447,N_15707);
xnor U27073 (N_27073,N_13002,N_13729);
nor U27074 (N_27074,N_16623,N_14147);
and U27075 (N_27075,N_16387,N_11755);
nor U27076 (N_27076,N_16495,N_11868);
nor U27077 (N_27077,N_15216,N_10764);
xnor U27078 (N_27078,N_13593,N_10544);
xnor U27079 (N_27079,N_16374,N_19641);
nor U27080 (N_27080,N_10593,N_18349);
nand U27081 (N_27081,N_13147,N_11838);
or U27082 (N_27082,N_17659,N_15889);
nand U27083 (N_27083,N_13833,N_16116);
and U27084 (N_27084,N_19343,N_14001);
and U27085 (N_27085,N_17222,N_16735);
xor U27086 (N_27086,N_16865,N_14629);
nand U27087 (N_27087,N_15366,N_17761);
and U27088 (N_27088,N_16329,N_14814);
or U27089 (N_27089,N_19851,N_10139);
nand U27090 (N_27090,N_12192,N_13120);
nor U27091 (N_27091,N_17440,N_17787);
nand U27092 (N_27092,N_13842,N_18304);
and U27093 (N_27093,N_15477,N_15693);
and U27094 (N_27094,N_10503,N_15948);
nor U27095 (N_27095,N_16999,N_15046);
or U27096 (N_27096,N_12837,N_15504);
nand U27097 (N_27097,N_14292,N_19774);
or U27098 (N_27098,N_10201,N_13821);
nor U27099 (N_27099,N_13008,N_19185);
and U27100 (N_27100,N_18722,N_19966);
nand U27101 (N_27101,N_13352,N_13112);
or U27102 (N_27102,N_16002,N_19114);
and U27103 (N_27103,N_19554,N_10313);
or U27104 (N_27104,N_17482,N_12009);
nand U27105 (N_27105,N_14576,N_14631);
or U27106 (N_27106,N_18949,N_19293);
xor U27107 (N_27107,N_15647,N_16631);
xor U27108 (N_27108,N_13945,N_19783);
nor U27109 (N_27109,N_17125,N_16099);
or U27110 (N_27110,N_15306,N_11177);
nand U27111 (N_27111,N_10957,N_10999);
nand U27112 (N_27112,N_16166,N_12398);
nand U27113 (N_27113,N_14072,N_14207);
nor U27114 (N_27114,N_18484,N_18684);
nand U27115 (N_27115,N_15103,N_11193);
nand U27116 (N_27116,N_15182,N_17269);
nand U27117 (N_27117,N_15987,N_12312);
and U27118 (N_27118,N_14441,N_16753);
xor U27119 (N_27119,N_16878,N_17165);
or U27120 (N_27120,N_10103,N_17418);
and U27121 (N_27121,N_10197,N_16831);
xor U27122 (N_27122,N_13507,N_17679);
or U27123 (N_27123,N_18401,N_19969);
nor U27124 (N_27124,N_11265,N_13304);
nand U27125 (N_27125,N_10148,N_16451);
nor U27126 (N_27126,N_10741,N_11600);
nand U27127 (N_27127,N_18076,N_12767);
nand U27128 (N_27128,N_10033,N_13929);
nand U27129 (N_27129,N_14221,N_11289);
nor U27130 (N_27130,N_15515,N_10292);
xnor U27131 (N_27131,N_11472,N_10618);
and U27132 (N_27132,N_11004,N_12983);
xor U27133 (N_27133,N_12996,N_17929);
or U27134 (N_27134,N_15401,N_10286);
or U27135 (N_27135,N_10259,N_14552);
xor U27136 (N_27136,N_10763,N_10970);
xnor U27137 (N_27137,N_17409,N_19964);
xnor U27138 (N_27138,N_14069,N_14556);
nand U27139 (N_27139,N_17942,N_15537);
nor U27140 (N_27140,N_16048,N_12496);
xnor U27141 (N_27141,N_11535,N_16141);
and U27142 (N_27142,N_10093,N_10567);
nand U27143 (N_27143,N_13814,N_15089);
xnor U27144 (N_27144,N_14791,N_16447);
and U27145 (N_27145,N_12019,N_11245);
xor U27146 (N_27146,N_13168,N_13956);
and U27147 (N_27147,N_17284,N_13192);
nor U27148 (N_27148,N_19679,N_10348);
xnor U27149 (N_27149,N_18891,N_15312);
nand U27150 (N_27150,N_12545,N_18498);
nor U27151 (N_27151,N_16074,N_13037);
nand U27152 (N_27152,N_10809,N_13650);
or U27153 (N_27153,N_18782,N_10733);
and U27154 (N_27154,N_14137,N_14403);
xor U27155 (N_27155,N_14782,N_15136);
or U27156 (N_27156,N_13392,N_14974);
nand U27157 (N_27157,N_10860,N_14876);
or U27158 (N_27158,N_18640,N_10730);
or U27159 (N_27159,N_13679,N_19550);
and U27160 (N_27160,N_12554,N_17853);
xor U27161 (N_27161,N_13235,N_16394);
nand U27162 (N_27162,N_13358,N_16656);
and U27163 (N_27163,N_13790,N_16855);
and U27164 (N_27164,N_10896,N_11103);
or U27165 (N_27165,N_13611,N_17946);
xnor U27166 (N_27166,N_16408,N_16140);
nand U27167 (N_27167,N_15615,N_19068);
and U27168 (N_27168,N_13869,N_11743);
xor U27169 (N_27169,N_19196,N_14467);
and U27170 (N_27170,N_16415,N_10583);
nor U27171 (N_27171,N_10895,N_16684);
nand U27172 (N_27172,N_10860,N_14105);
nor U27173 (N_27173,N_19420,N_15752);
nor U27174 (N_27174,N_18263,N_12528);
or U27175 (N_27175,N_19272,N_11481);
or U27176 (N_27176,N_11174,N_12160);
or U27177 (N_27177,N_10115,N_11050);
and U27178 (N_27178,N_15522,N_14154);
and U27179 (N_27179,N_15928,N_16661);
nor U27180 (N_27180,N_19556,N_17205);
xor U27181 (N_27181,N_16688,N_18880);
nand U27182 (N_27182,N_19061,N_16066);
xnor U27183 (N_27183,N_11669,N_10070);
nand U27184 (N_27184,N_14673,N_11852);
or U27185 (N_27185,N_17540,N_17756);
nand U27186 (N_27186,N_13977,N_10493);
and U27187 (N_27187,N_18456,N_16567);
nand U27188 (N_27188,N_18873,N_17386);
xnor U27189 (N_27189,N_11811,N_14501);
and U27190 (N_27190,N_12729,N_10345);
or U27191 (N_27191,N_19775,N_14908);
xnor U27192 (N_27192,N_14254,N_17089);
or U27193 (N_27193,N_16739,N_10237);
xor U27194 (N_27194,N_19276,N_16363);
xor U27195 (N_27195,N_17067,N_19290);
and U27196 (N_27196,N_15856,N_10708);
xor U27197 (N_27197,N_11704,N_19634);
xnor U27198 (N_27198,N_15113,N_15448);
nand U27199 (N_27199,N_17986,N_15195);
nand U27200 (N_27200,N_16706,N_13924);
xor U27201 (N_27201,N_15115,N_14026);
nor U27202 (N_27202,N_14767,N_11751);
and U27203 (N_27203,N_11562,N_10408);
and U27204 (N_27204,N_18671,N_19432);
nor U27205 (N_27205,N_16283,N_13452);
and U27206 (N_27206,N_12361,N_10101);
or U27207 (N_27207,N_16163,N_13942);
nand U27208 (N_27208,N_12049,N_10282);
or U27209 (N_27209,N_17441,N_17554);
or U27210 (N_27210,N_12940,N_15911);
nand U27211 (N_27211,N_16465,N_19033);
xor U27212 (N_27212,N_15785,N_19349);
xnor U27213 (N_27213,N_11487,N_16530);
nor U27214 (N_27214,N_10206,N_16203);
nor U27215 (N_27215,N_10243,N_14081);
xor U27216 (N_27216,N_15020,N_13354);
nand U27217 (N_27217,N_11128,N_18903);
and U27218 (N_27218,N_16836,N_12720);
nand U27219 (N_27219,N_11557,N_18506);
and U27220 (N_27220,N_15055,N_13584);
nand U27221 (N_27221,N_12248,N_11989);
or U27222 (N_27222,N_16765,N_13714);
nand U27223 (N_27223,N_10195,N_12154);
or U27224 (N_27224,N_13537,N_10065);
or U27225 (N_27225,N_18306,N_16699);
nor U27226 (N_27226,N_15894,N_12271);
xor U27227 (N_27227,N_17483,N_13073);
and U27228 (N_27228,N_14972,N_17739);
and U27229 (N_27229,N_19846,N_14517);
or U27230 (N_27230,N_11633,N_13718);
or U27231 (N_27231,N_14906,N_13554);
nand U27232 (N_27232,N_10749,N_15096);
nor U27233 (N_27233,N_14521,N_13585);
nor U27234 (N_27234,N_18566,N_17556);
and U27235 (N_27235,N_14073,N_17431);
and U27236 (N_27236,N_18701,N_13083);
nand U27237 (N_27237,N_16652,N_13006);
nor U27238 (N_27238,N_13536,N_11835);
nand U27239 (N_27239,N_10779,N_15603);
nor U27240 (N_27240,N_16779,N_16595);
nand U27241 (N_27241,N_19997,N_10288);
nand U27242 (N_27242,N_11211,N_15854);
nor U27243 (N_27243,N_11212,N_17034);
nand U27244 (N_27244,N_19398,N_18662);
nand U27245 (N_27245,N_13280,N_12481);
nand U27246 (N_27246,N_19465,N_16816);
nand U27247 (N_27247,N_14821,N_18975);
nand U27248 (N_27248,N_10253,N_11924);
or U27249 (N_27249,N_19963,N_13670);
xnor U27250 (N_27250,N_16123,N_10494);
xor U27251 (N_27251,N_11590,N_17017);
xor U27252 (N_27252,N_10950,N_16263);
or U27253 (N_27253,N_14781,N_19460);
nand U27254 (N_27254,N_12631,N_13198);
nand U27255 (N_27255,N_11768,N_14735);
xnor U27256 (N_27256,N_15210,N_17444);
and U27257 (N_27257,N_11633,N_11124);
and U27258 (N_27258,N_16917,N_16508);
and U27259 (N_27259,N_13666,N_16661);
nand U27260 (N_27260,N_10368,N_16295);
nand U27261 (N_27261,N_11873,N_10762);
nand U27262 (N_27262,N_11755,N_18106);
and U27263 (N_27263,N_13852,N_11820);
nand U27264 (N_27264,N_10162,N_10488);
or U27265 (N_27265,N_15974,N_12851);
or U27266 (N_27266,N_19758,N_15162);
nor U27267 (N_27267,N_14002,N_15252);
or U27268 (N_27268,N_10037,N_11712);
nor U27269 (N_27269,N_14750,N_15675);
and U27270 (N_27270,N_15985,N_15143);
xor U27271 (N_27271,N_19420,N_19895);
nor U27272 (N_27272,N_15046,N_19863);
xnor U27273 (N_27273,N_16523,N_17307);
nand U27274 (N_27274,N_15088,N_18719);
or U27275 (N_27275,N_16431,N_15708);
nor U27276 (N_27276,N_15958,N_13342);
or U27277 (N_27277,N_18197,N_10196);
xor U27278 (N_27278,N_12761,N_19109);
nand U27279 (N_27279,N_16943,N_11328);
xnor U27280 (N_27280,N_12206,N_16795);
nand U27281 (N_27281,N_14467,N_10511);
and U27282 (N_27282,N_16087,N_12800);
xor U27283 (N_27283,N_18209,N_11666);
xor U27284 (N_27284,N_11693,N_14459);
and U27285 (N_27285,N_12299,N_17827);
and U27286 (N_27286,N_18261,N_11577);
nand U27287 (N_27287,N_12064,N_14957);
and U27288 (N_27288,N_12740,N_15400);
xor U27289 (N_27289,N_10482,N_13210);
nand U27290 (N_27290,N_11450,N_10425);
xor U27291 (N_27291,N_18145,N_19698);
nand U27292 (N_27292,N_16154,N_18416);
or U27293 (N_27293,N_19278,N_17322);
or U27294 (N_27294,N_18010,N_18872);
xor U27295 (N_27295,N_15829,N_18122);
nor U27296 (N_27296,N_16175,N_10050);
nand U27297 (N_27297,N_19531,N_10892);
and U27298 (N_27298,N_10289,N_19462);
and U27299 (N_27299,N_10469,N_16666);
nor U27300 (N_27300,N_19506,N_11012);
nand U27301 (N_27301,N_18748,N_13184);
nor U27302 (N_27302,N_14583,N_10974);
nand U27303 (N_27303,N_10370,N_18952);
nor U27304 (N_27304,N_10968,N_17769);
xnor U27305 (N_27305,N_12852,N_18340);
or U27306 (N_27306,N_19845,N_11106);
and U27307 (N_27307,N_12294,N_14428);
xor U27308 (N_27308,N_14416,N_14524);
nor U27309 (N_27309,N_14275,N_10945);
nor U27310 (N_27310,N_11085,N_10270);
nand U27311 (N_27311,N_19189,N_12911);
and U27312 (N_27312,N_11973,N_15014);
nand U27313 (N_27313,N_19072,N_10820);
or U27314 (N_27314,N_11986,N_15192);
and U27315 (N_27315,N_14836,N_12606);
or U27316 (N_27316,N_10062,N_14409);
nand U27317 (N_27317,N_10830,N_13670);
nor U27318 (N_27318,N_11696,N_13617);
and U27319 (N_27319,N_13559,N_10427);
and U27320 (N_27320,N_12630,N_16968);
nor U27321 (N_27321,N_15317,N_14122);
and U27322 (N_27322,N_13812,N_11498);
nor U27323 (N_27323,N_18096,N_12072);
nor U27324 (N_27324,N_13182,N_13811);
xor U27325 (N_27325,N_19844,N_18958);
nor U27326 (N_27326,N_16783,N_18102);
nand U27327 (N_27327,N_16212,N_13000);
or U27328 (N_27328,N_15473,N_16964);
nor U27329 (N_27329,N_15822,N_10638);
and U27330 (N_27330,N_15237,N_17738);
or U27331 (N_27331,N_12595,N_12764);
nand U27332 (N_27332,N_13444,N_15350);
xor U27333 (N_27333,N_13703,N_13373);
or U27334 (N_27334,N_10582,N_11833);
nor U27335 (N_27335,N_17137,N_12989);
xor U27336 (N_27336,N_14021,N_13781);
xor U27337 (N_27337,N_18948,N_11152);
and U27338 (N_27338,N_19336,N_15865);
and U27339 (N_27339,N_16496,N_18127);
nand U27340 (N_27340,N_16739,N_10393);
and U27341 (N_27341,N_14005,N_16111);
and U27342 (N_27342,N_16842,N_10109);
nand U27343 (N_27343,N_15119,N_15158);
xor U27344 (N_27344,N_18657,N_15710);
or U27345 (N_27345,N_19008,N_18440);
xor U27346 (N_27346,N_15097,N_14455);
or U27347 (N_27347,N_11467,N_17091);
nand U27348 (N_27348,N_19518,N_13869);
nand U27349 (N_27349,N_16201,N_16618);
or U27350 (N_27350,N_10500,N_18363);
xnor U27351 (N_27351,N_18537,N_11888);
or U27352 (N_27352,N_19441,N_13548);
and U27353 (N_27353,N_14074,N_14065);
or U27354 (N_27354,N_17762,N_15611);
or U27355 (N_27355,N_11360,N_11944);
and U27356 (N_27356,N_16498,N_12688);
and U27357 (N_27357,N_12453,N_15394);
nand U27358 (N_27358,N_11358,N_13821);
nand U27359 (N_27359,N_14475,N_13391);
or U27360 (N_27360,N_16346,N_18501);
nor U27361 (N_27361,N_11495,N_12123);
and U27362 (N_27362,N_11785,N_10261);
or U27363 (N_27363,N_16345,N_11310);
nor U27364 (N_27364,N_18390,N_17871);
and U27365 (N_27365,N_12148,N_16346);
and U27366 (N_27366,N_12535,N_18690);
xnor U27367 (N_27367,N_14149,N_13971);
nor U27368 (N_27368,N_12326,N_19551);
or U27369 (N_27369,N_12274,N_13794);
nor U27370 (N_27370,N_14637,N_16066);
nor U27371 (N_27371,N_10920,N_18715);
and U27372 (N_27372,N_12064,N_12284);
and U27373 (N_27373,N_17857,N_12274);
or U27374 (N_27374,N_15886,N_11938);
or U27375 (N_27375,N_19889,N_13539);
and U27376 (N_27376,N_19971,N_13517);
or U27377 (N_27377,N_10174,N_13290);
nor U27378 (N_27378,N_11978,N_19321);
nand U27379 (N_27379,N_18331,N_18478);
nor U27380 (N_27380,N_16953,N_19931);
nor U27381 (N_27381,N_18759,N_12233);
or U27382 (N_27382,N_13897,N_15733);
and U27383 (N_27383,N_13024,N_13958);
nand U27384 (N_27384,N_10549,N_14999);
nand U27385 (N_27385,N_15534,N_18734);
and U27386 (N_27386,N_11515,N_16662);
nand U27387 (N_27387,N_15707,N_18318);
or U27388 (N_27388,N_17786,N_15349);
xnor U27389 (N_27389,N_15195,N_13148);
or U27390 (N_27390,N_19322,N_11742);
nand U27391 (N_27391,N_15415,N_14741);
nand U27392 (N_27392,N_17170,N_12198);
xnor U27393 (N_27393,N_11380,N_15021);
and U27394 (N_27394,N_15468,N_15072);
and U27395 (N_27395,N_13030,N_12476);
and U27396 (N_27396,N_16718,N_15653);
or U27397 (N_27397,N_12027,N_16498);
nand U27398 (N_27398,N_16301,N_16998);
nand U27399 (N_27399,N_15932,N_17271);
nor U27400 (N_27400,N_10739,N_18037);
nand U27401 (N_27401,N_15844,N_13367);
or U27402 (N_27402,N_19489,N_15514);
or U27403 (N_27403,N_15949,N_13232);
or U27404 (N_27404,N_18570,N_11033);
nor U27405 (N_27405,N_17319,N_19660);
nand U27406 (N_27406,N_10348,N_13906);
or U27407 (N_27407,N_19001,N_15949);
and U27408 (N_27408,N_18450,N_18744);
nor U27409 (N_27409,N_19833,N_18530);
nor U27410 (N_27410,N_10770,N_10308);
and U27411 (N_27411,N_18567,N_10975);
nor U27412 (N_27412,N_11457,N_18642);
xor U27413 (N_27413,N_18988,N_12684);
and U27414 (N_27414,N_11323,N_15291);
nand U27415 (N_27415,N_16049,N_16863);
nand U27416 (N_27416,N_17040,N_13730);
or U27417 (N_27417,N_10892,N_17458);
or U27418 (N_27418,N_10911,N_18801);
nand U27419 (N_27419,N_19421,N_14468);
nor U27420 (N_27420,N_11637,N_10071);
xnor U27421 (N_27421,N_13772,N_15741);
or U27422 (N_27422,N_14189,N_13748);
nor U27423 (N_27423,N_18533,N_13934);
and U27424 (N_27424,N_17126,N_10234);
or U27425 (N_27425,N_15093,N_15224);
nor U27426 (N_27426,N_16537,N_19615);
or U27427 (N_27427,N_16284,N_12741);
xnor U27428 (N_27428,N_11521,N_13857);
nand U27429 (N_27429,N_10796,N_19787);
or U27430 (N_27430,N_16094,N_18452);
nand U27431 (N_27431,N_11429,N_16169);
nand U27432 (N_27432,N_10517,N_15979);
and U27433 (N_27433,N_11099,N_15711);
xnor U27434 (N_27434,N_15588,N_18688);
and U27435 (N_27435,N_18021,N_16697);
nand U27436 (N_27436,N_13938,N_13832);
nand U27437 (N_27437,N_17186,N_18096);
nand U27438 (N_27438,N_17967,N_17685);
or U27439 (N_27439,N_19652,N_12585);
or U27440 (N_27440,N_12520,N_12633);
or U27441 (N_27441,N_11841,N_18478);
or U27442 (N_27442,N_12164,N_13352);
nor U27443 (N_27443,N_19287,N_10785);
or U27444 (N_27444,N_15460,N_16782);
nand U27445 (N_27445,N_12648,N_13289);
or U27446 (N_27446,N_11609,N_19080);
or U27447 (N_27447,N_11255,N_17542);
nor U27448 (N_27448,N_18681,N_16900);
nor U27449 (N_27449,N_17815,N_15974);
nand U27450 (N_27450,N_13183,N_16626);
xor U27451 (N_27451,N_11468,N_11714);
nand U27452 (N_27452,N_16942,N_13176);
nand U27453 (N_27453,N_16635,N_16531);
or U27454 (N_27454,N_19062,N_15769);
xor U27455 (N_27455,N_15835,N_17094);
xnor U27456 (N_27456,N_18134,N_14330);
nand U27457 (N_27457,N_19669,N_19427);
or U27458 (N_27458,N_16388,N_19004);
or U27459 (N_27459,N_14047,N_12778);
or U27460 (N_27460,N_17977,N_12765);
nand U27461 (N_27461,N_12755,N_14817);
nand U27462 (N_27462,N_11954,N_17896);
nand U27463 (N_27463,N_18961,N_11751);
xnor U27464 (N_27464,N_11477,N_12156);
and U27465 (N_27465,N_18463,N_11457);
and U27466 (N_27466,N_10222,N_16010);
nor U27467 (N_27467,N_12614,N_14834);
or U27468 (N_27468,N_19934,N_12408);
nor U27469 (N_27469,N_12127,N_14589);
xnor U27470 (N_27470,N_10612,N_11356);
xnor U27471 (N_27471,N_12073,N_14114);
xor U27472 (N_27472,N_18894,N_12060);
xor U27473 (N_27473,N_18462,N_12476);
nand U27474 (N_27474,N_19851,N_15341);
nor U27475 (N_27475,N_10437,N_18941);
nor U27476 (N_27476,N_14244,N_12916);
nand U27477 (N_27477,N_11974,N_15721);
xor U27478 (N_27478,N_16822,N_17944);
nor U27479 (N_27479,N_12736,N_15499);
nor U27480 (N_27480,N_19141,N_15648);
nor U27481 (N_27481,N_15596,N_17264);
or U27482 (N_27482,N_10190,N_19846);
nand U27483 (N_27483,N_17028,N_13570);
and U27484 (N_27484,N_17994,N_16754);
or U27485 (N_27485,N_12285,N_19666);
xnor U27486 (N_27486,N_11049,N_16906);
xnor U27487 (N_27487,N_15405,N_10931);
nor U27488 (N_27488,N_17219,N_11516);
and U27489 (N_27489,N_11311,N_14407);
and U27490 (N_27490,N_10679,N_19927);
or U27491 (N_27491,N_16333,N_12684);
or U27492 (N_27492,N_13858,N_13777);
or U27493 (N_27493,N_11136,N_12257);
xnor U27494 (N_27494,N_10395,N_11474);
and U27495 (N_27495,N_15794,N_10770);
xnor U27496 (N_27496,N_12537,N_17781);
nor U27497 (N_27497,N_14455,N_10012);
or U27498 (N_27498,N_11027,N_16786);
xor U27499 (N_27499,N_14452,N_14902);
xnor U27500 (N_27500,N_10536,N_12884);
or U27501 (N_27501,N_16756,N_11512);
and U27502 (N_27502,N_11054,N_11695);
xnor U27503 (N_27503,N_17328,N_19125);
and U27504 (N_27504,N_16479,N_12362);
xnor U27505 (N_27505,N_12354,N_13774);
or U27506 (N_27506,N_12800,N_14266);
nor U27507 (N_27507,N_15027,N_11057);
and U27508 (N_27508,N_19465,N_19092);
nor U27509 (N_27509,N_16520,N_10515);
nand U27510 (N_27510,N_19956,N_17230);
nand U27511 (N_27511,N_18463,N_10083);
xor U27512 (N_27512,N_17187,N_11032);
and U27513 (N_27513,N_19319,N_13343);
and U27514 (N_27514,N_13362,N_17454);
nor U27515 (N_27515,N_10287,N_10616);
nor U27516 (N_27516,N_13254,N_19132);
and U27517 (N_27517,N_12572,N_19571);
nand U27518 (N_27518,N_15437,N_18915);
or U27519 (N_27519,N_12591,N_13883);
nand U27520 (N_27520,N_10870,N_13678);
nor U27521 (N_27521,N_18615,N_15403);
nor U27522 (N_27522,N_16058,N_17718);
nand U27523 (N_27523,N_13920,N_18186);
xnor U27524 (N_27524,N_12723,N_13516);
and U27525 (N_27525,N_18439,N_16638);
and U27526 (N_27526,N_13420,N_15616);
nand U27527 (N_27527,N_18940,N_17017);
nor U27528 (N_27528,N_13973,N_16008);
xor U27529 (N_27529,N_14027,N_13794);
and U27530 (N_27530,N_10686,N_12820);
xnor U27531 (N_27531,N_13001,N_16689);
xnor U27532 (N_27532,N_18935,N_12168);
or U27533 (N_27533,N_18861,N_15991);
nand U27534 (N_27534,N_17532,N_14462);
xor U27535 (N_27535,N_13931,N_15862);
nand U27536 (N_27536,N_15369,N_18360);
nand U27537 (N_27537,N_13815,N_15881);
and U27538 (N_27538,N_11669,N_18618);
nand U27539 (N_27539,N_15217,N_10703);
nand U27540 (N_27540,N_12671,N_18726);
nand U27541 (N_27541,N_11880,N_16480);
nand U27542 (N_27542,N_14731,N_16563);
or U27543 (N_27543,N_17200,N_17084);
and U27544 (N_27544,N_16036,N_13480);
and U27545 (N_27545,N_10587,N_10096);
or U27546 (N_27546,N_16533,N_12799);
nor U27547 (N_27547,N_18917,N_14193);
or U27548 (N_27548,N_17443,N_16967);
nand U27549 (N_27549,N_10417,N_11123);
and U27550 (N_27550,N_16820,N_14977);
or U27551 (N_27551,N_12329,N_13658);
or U27552 (N_27552,N_14114,N_15044);
and U27553 (N_27553,N_17551,N_13122);
nor U27554 (N_27554,N_10370,N_10204);
nor U27555 (N_27555,N_10950,N_18081);
nor U27556 (N_27556,N_17451,N_11705);
nor U27557 (N_27557,N_10078,N_11068);
nor U27558 (N_27558,N_18332,N_15829);
nand U27559 (N_27559,N_12450,N_13523);
and U27560 (N_27560,N_18865,N_12707);
or U27561 (N_27561,N_18042,N_14046);
xor U27562 (N_27562,N_12594,N_13373);
and U27563 (N_27563,N_18928,N_14566);
nor U27564 (N_27564,N_13918,N_18760);
nor U27565 (N_27565,N_14998,N_12036);
nand U27566 (N_27566,N_11818,N_19570);
nor U27567 (N_27567,N_18655,N_11879);
or U27568 (N_27568,N_15758,N_15746);
nor U27569 (N_27569,N_13750,N_14843);
xnor U27570 (N_27570,N_19943,N_11810);
and U27571 (N_27571,N_10560,N_12529);
nand U27572 (N_27572,N_16866,N_16226);
and U27573 (N_27573,N_10045,N_13332);
or U27574 (N_27574,N_15729,N_17379);
and U27575 (N_27575,N_16347,N_15429);
or U27576 (N_27576,N_18343,N_10447);
nand U27577 (N_27577,N_10664,N_12638);
nor U27578 (N_27578,N_13506,N_12672);
nand U27579 (N_27579,N_15964,N_16459);
nor U27580 (N_27580,N_19987,N_13319);
xnor U27581 (N_27581,N_12295,N_18734);
xnor U27582 (N_27582,N_14544,N_15665);
nor U27583 (N_27583,N_11825,N_16080);
and U27584 (N_27584,N_14611,N_18155);
xnor U27585 (N_27585,N_15252,N_13586);
or U27586 (N_27586,N_16227,N_11510);
xnor U27587 (N_27587,N_17286,N_19444);
nor U27588 (N_27588,N_10944,N_14989);
or U27589 (N_27589,N_11718,N_17495);
and U27590 (N_27590,N_12134,N_16253);
and U27591 (N_27591,N_11059,N_15495);
nand U27592 (N_27592,N_15635,N_17624);
or U27593 (N_27593,N_16661,N_12646);
nor U27594 (N_27594,N_11179,N_17073);
xnor U27595 (N_27595,N_12680,N_14903);
nand U27596 (N_27596,N_17141,N_10970);
nor U27597 (N_27597,N_16287,N_18520);
xnor U27598 (N_27598,N_10684,N_14645);
or U27599 (N_27599,N_15941,N_12597);
or U27600 (N_27600,N_15849,N_13654);
nor U27601 (N_27601,N_15926,N_14859);
and U27602 (N_27602,N_12267,N_12923);
and U27603 (N_27603,N_17323,N_18258);
xnor U27604 (N_27604,N_16148,N_12398);
nor U27605 (N_27605,N_14074,N_13606);
nand U27606 (N_27606,N_17779,N_13344);
nand U27607 (N_27607,N_11577,N_14819);
or U27608 (N_27608,N_10038,N_12235);
xor U27609 (N_27609,N_14494,N_12203);
and U27610 (N_27610,N_19458,N_10441);
and U27611 (N_27611,N_14518,N_13211);
or U27612 (N_27612,N_12855,N_15490);
nand U27613 (N_27613,N_19177,N_18101);
and U27614 (N_27614,N_14207,N_12159);
and U27615 (N_27615,N_11668,N_13001);
nand U27616 (N_27616,N_13464,N_14831);
nand U27617 (N_27617,N_16145,N_18724);
nand U27618 (N_27618,N_15316,N_16003);
xnor U27619 (N_27619,N_19373,N_16760);
nand U27620 (N_27620,N_12276,N_15861);
xor U27621 (N_27621,N_10295,N_14132);
nand U27622 (N_27622,N_19205,N_13609);
xnor U27623 (N_27623,N_12455,N_17780);
nor U27624 (N_27624,N_10157,N_10850);
or U27625 (N_27625,N_17928,N_13365);
or U27626 (N_27626,N_12192,N_13000);
and U27627 (N_27627,N_15739,N_18078);
and U27628 (N_27628,N_14481,N_12020);
or U27629 (N_27629,N_11852,N_17912);
or U27630 (N_27630,N_17773,N_17901);
nand U27631 (N_27631,N_19905,N_13720);
nor U27632 (N_27632,N_19183,N_14985);
nor U27633 (N_27633,N_18344,N_13520);
nand U27634 (N_27634,N_14034,N_19280);
nand U27635 (N_27635,N_14834,N_19818);
xnor U27636 (N_27636,N_17637,N_11146);
nor U27637 (N_27637,N_11416,N_13632);
nor U27638 (N_27638,N_11661,N_13029);
or U27639 (N_27639,N_16909,N_18437);
xnor U27640 (N_27640,N_19798,N_14339);
nor U27641 (N_27641,N_12565,N_17187);
or U27642 (N_27642,N_17666,N_13191);
and U27643 (N_27643,N_12066,N_14820);
nand U27644 (N_27644,N_13173,N_14719);
nand U27645 (N_27645,N_12194,N_17665);
or U27646 (N_27646,N_15606,N_17565);
or U27647 (N_27647,N_12419,N_11357);
or U27648 (N_27648,N_15960,N_10991);
nor U27649 (N_27649,N_13112,N_16346);
and U27650 (N_27650,N_19502,N_19171);
nand U27651 (N_27651,N_16445,N_14013);
nand U27652 (N_27652,N_16113,N_17132);
xor U27653 (N_27653,N_18050,N_10514);
xor U27654 (N_27654,N_19609,N_10886);
or U27655 (N_27655,N_14233,N_10298);
and U27656 (N_27656,N_14471,N_10042);
or U27657 (N_27657,N_12436,N_18009);
xnor U27658 (N_27658,N_14909,N_11406);
nand U27659 (N_27659,N_19381,N_10087);
or U27660 (N_27660,N_11158,N_16019);
nand U27661 (N_27661,N_12673,N_16050);
xnor U27662 (N_27662,N_14702,N_19493);
nor U27663 (N_27663,N_12909,N_18668);
or U27664 (N_27664,N_19367,N_17380);
xnor U27665 (N_27665,N_10220,N_18341);
nand U27666 (N_27666,N_13184,N_14590);
or U27667 (N_27667,N_12548,N_12417);
or U27668 (N_27668,N_19722,N_18506);
nor U27669 (N_27669,N_11188,N_18100);
and U27670 (N_27670,N_19881,N_12247);
nand U27671 (N_27671,N_19115,N_19001);
nor U27672 (N_27672,N_19064,N_16341);
and U27673 (N_27673,N_11262,N_11496);
nand U27674 (N_27674,N_19981,N_10801);
nand U27675 (N_27675,N_13243,N_17366);
xor U27676 (N_27676,N_19407,N_12550);
nand U27677 (N_27677,N_13376,N_16886);
nor U27678 (N_27678,N_10646,N_10337);
xor U27679 (N_27679,N_16407,N_13273);
nor U27680 (N_27680,N_19708,N_11364);
and U27681 (N_27681,N_16504,N_17005);
nand U27682 (N_27682,N_14746,N_11165);
nor U27683 (N_27683,N_13723,N_18259);
or U27684 (N_27684,N_10425,N_12200);
nor U27685 (N_27685,N_18556,N_12437);
xnor U27686 (N_27686,N_13554,N_12487);
xnor U27687 (N_27687,N_10372,N_19446);
nand U27688 (N_27688,N_17663,N_15661);
xor U27689 (N_27689,N_12681,N_10088);
nor U27690 (N_27690,N_19240,N_19915);
nand U27691 (N_27691,N_11648,N_16363);
nand U27692 (N_27692,N_17202,N_18105);
or U27693 (N_27693,N_11392,N_13576);
or U27694 (N_27694,N_14971,N_19687);
nand U27695 (N_27695,N_10893,N_10778);
xnor U27696 (N_27696,N_10145,N_17614);
nand U27697 (N_27697,N_17762,N_17751);
and U27698 (N_27698,N_19494,N_12267);
nand U27699 (N_27699,N_17185,N_12276);
or U27700 (N_27700,N_15531,N_14519);
xor U27701 (N_27701,N_11969,N_13671);
or U27702 (N_27702,N_16942,N_13027);
and U27703 (N_27703,N_18181,N_14069);
or U27704 (N_27704,N_15244,N_11774);
nand U27705 (N_27705,N_11576,N_12764);
nor U27706 (N_27706,N_18443,N_13609);
or U27707 (N_27707,N_19072,N_18302);
and U27708 (N_27708,N_17902,N_16987);
nand U27709 (N_27709,N_17657,N_16281);
nor U27710 (N_27710,N_15848,N_10036);
or U27711 (N_27711,N_15516,N_19644);
nand U27712 (N_27712,N_10471,N_18351);
or U27713 (N_27713,N_12798,N_17577);
or U27714 (N_27714,N_10070,N_14760);
nand U27715 (N_27715,N_13396,N_15920);
xnor U27716 (N_27716,N_19604,N_17543);
nor U27717 (N_27717,N_16060,N_15775);
nor U27718 (N_27718,N_19778,N_19609);
and U27719 (N_27719,N_13466,N_10650);
nor U27720 (N_27720,N_16495,N_16141);
and U27721 (N_27721,N_11950,N_18613);
nor U27722 (N_27722,N_13059,N_14661);
nand U27723 (N_27723,N_16443,N_19849);
nand U27724 (N_27724,N_18120,N_19651);
nand U27725 (N_27725,N_12673,N_15921);
xnor U27726 (N_27726,N_10892,N_12343);
xnor U27727 (N_27727,N_11713,N_10208);
and U27728 (N_27728,N_12859,N_12270);
nor U27729 (N_27729,N_17900,N_15778);
and U27730 (N_27730,N_12310,N_17727);
or U27731 (N_27731,N_11730,N_19298);
nor U27732 (N_27732,N_17540,N_13512);
nand U27733 (N_27733,N_11090,N_15535);
nand U27734 (N_27734,N_14508,N_19354);
or U27735 (N_27735,N_15659,N_11504);
or U27736 (N_27736,N_15973,N_18104);
xor U27737 (N_27737,N_14067,N_12537);
or U27738 (N_27738,N_10362,N_17166);
and U27739 (N_27739,N_10206,N_17855);
nor U27740 (N_27740,N_12360,N_14661);
and U27741 (N_27741,N_16604,N_14647);
or U27742 (N_27742,N_17612,N_13074);
xor U27743 (N_27743,N_15356,N_17834);
and U27744 (N_27744,N_13314,N_19797);
xor U27745 (N_27745,N_10344,N_15904);
xor U27746 (N_27746,N_11936,N_12502);
nor U27747 (N_27747,N_13724,N_11370);
and U27748 (N_27748,N_10587,N_13979);
xnor U27749 (N_27749,N_18869,N_18223);
and U27750 (N_27750,N_13341,N_18427);
and U27751 (N_27751,N_15517,N_17035);
or U27752 (N_27752,N_19239,N_15202);
nand U27753 (N_27753,N_10553,N_19584);
and U27754 (N_27754,N_16489,N_16420);
nand U27755 (N_27755,N_11046,N_19148);
and U27756 (N_27756,N_17061,N_13414);
or U27757 (N_27757,N_18129,N_16364);
and U27758 (N_27758,N_19485,N_15476);
or U27759 (N_27759,N_17861,N_10430);
nor U27760 (N_27760,N_10986,N_16824);
xnor U27761 (N_27761,N_14910,N_14081);
nand U27762 (N_27762,N_14872,N_12788);
or U27763 (N_27763,N_15288,N_17644);
nor U27764 (N_27764,N_12218,N_17449);
xnor U27765 (N_27765,N_11112,N_18169);
or U27766 (N_27766,N_17954,N_12590);
nand U27767 (N_27767,N_11043,N_13940);
or U27768 (N_27768,N_10819,N_18033);
nor U27769 (N_27769,N_15465,N_12455);
xnor U27770 (N_27770,N_13593,N_19338);
nand U27771 (N_27771,N_16556,N_17369);
nand U27772 (N_27772,N_11067,N_16868);
xnor U27773 (N_27773,N_11929,N_19035);
or U27774 (N_27774,N_17634,N_11853);
nor U27775 (N_27775,N_17583,N_13685);
and U27776 (N_27776,N_15803,N_15142);
nor U27777 (N_27777,N_18927,N_12837);
nor U27778 (N_27778,N_17027,N_11751);
nor U27779 (N_27779,N_11857,N_15323);
or U27780 (N_27780,N_15592,N_19735);
nor U27781 (N_27781,N_13680,N_11671);
or U27782 (N_27782,N_11601,N_10163);
nor U27783 (N_27783,N_15881,N_11674);
nand U27784 (N_27784,N_18050,N_19993);
or U27785 (N_27785,N_15085,N_16383);
nor U27786 (N_27786,N_13584,N_18147);
nor U27787 (N_27787,N_16364,N_13921);
or U27788 (N_27788,N_18080,N_14457);
nor U27789 (N_27789,N_14381,N_16635);
or U27790 (N_27790,N_15728,N_11006);
xor U27791 (N_27791,N_16789,N_16352);
xor U27792 (N_27792,N_18000,N_15678);
nor U27793 (N_27793,N_19884,N_16601);
xnor U27794 (N_27794,N_10308,N_15715);
and U27795 (N_27795,N_13998,N_13462);
xor U27796 (N_27796,N_18105,N_13280);
or U27797 (N_27797,N_18997,N_19642);
xor U27798 (N_27798,N_14055,N_17442);
nand U27799 (N_27799,N_17679,N_14446);
xor U27800 (N_27800,N_13544,N_16885);
xnor U27801 (N_27801,N_11667,N_16394);
nand U27802 (N_27802,N_17455,N_18923);
and U27803 (N_27803,N_19711,N_15453);
nor U27804 (N_27804,N_10247,N_12201);
and U27805 (N_27805,N_15953,N_15637);
nor U27806 (N_27806,N_17061,N_14424);
nand U27807 (N_27807,N_13767,N_16907);
nand U27808 (N_27808,N_18692,N_14572);
xnor U27809 (N_27809,N_12266,N_10004);
and U27810 (N_27810,N_10697,N_10393);
or U27811 (N_27811,N_12927,N_16567);
and U27812 (N_27812,N_17758,N_17263);
and U27813 (N_27813,N_14984,N_14119);
and U27814 (N_27814,N_14411,N_18560);
nor U27815 (N_27815,N_19196,N_15045);
and U27816 (N_27816,N_13716,N_11080);
and U27817 (N_27817,N_18587,N_17410);
xor U27818 (N_27818,N_16234,N_19286);
nor U27819 (N_27819,N_18302,N_17319);
xor U27820 (N_27820,N_19513,N_18964);
xnor U27821 (N_27821,N_15840,N_13800);
nand U27822 (N_27822,N_16636,N_16943);
xor U27823 (N_27823,N_14841,N_10787);
and U27824 (N_27824,N_12233,N_13304);
or U27825 (N_27825,N_15708,N_12410);
or U27826 (N_27826,N_11536,N_16906);
and U27827 (N_27827,N_14452,N_13802);
nor U27828 (N_27828,N_17671,N_19041);
or U27829 (N_27829,N_19079,N_17754);
or U27830 (N_27830,N_13020,N_15290);
xor U27831 (N_27831,N_10437,N_16790);
and U27832 (N_27832,N_14447,N_17613);
and U27833 (N_27833,N_12598,N_13709);
nand U27834 (N_27834,N_12539,N_13060);
nand U27835 (N_27835,N_14254,N_15299);
nand U27836 (N_27836,N_19387,N_13813);
xor U27837 (N_27837,N_11324,N_19298);
and U27838 (N_27838,N_15356,N_17179);
or U27839 (N_27839,N_15005,N_19149);
or U27840 (N_27840,N_13299,N_11764);
nor U27841 (N_27841,N_17884,N_19536);
nand U27842 (N_27842,N_17191,N_10677);
nor U27843 (N_27843,N_13810,N_16519);
and U27844 (N_27844,N_17400,N_17995);
and U27845 (N_27845,N_10072,N_12033);
or U27846 (N_27846,N_14822,N_17178);
or U27847 (N_27847,N_17085,N_19300);
and U27848 (N_27848,N_12569,N_16768);
nand U27849 (N_27849,N_15535,N_15934);
or U27850 (N_27850,N_12739,N_15742);
and U27851 (N_27851,N_17989,N_18713);
nand U27852 (N_27852,N_11385,N_12708);
nand U27853 (N_27853,N_14873,N_11322);
xnor U27854 (N_27854,N_19979,N_13847);
or U27855 (N_27855,N_19236,N_12099);
nand U27856 (N_27856,N_14749,N_10765);
or U27857 (N_27857,N_17772,N_15015);
nand U27858 (N_27858,N_18654,N_15725);
nand U27859 (N_27859,N_17040,N_14639);
or U27860 (N_27860,N_13522,N_14973);
or U27861 (N_27861,N_13620,N_10260);
nand U27862 (N_27862,N_15470,N_13077);
xor U27863 (N_27863,N_16290,N_10571);
nand U27864 (N_27864,N_15832,N_15619);
xor U27865 (N_27865,N_14811,N_16662);
nor U27866 (N_27866,N_13159,N_16560);
or U27867 (N_27867,N_18436,N_15962);
nand U27868 (N_27868,N_17701,N_19123);
nand U27869 (N_27869,N_13490,N_10210);
and U27870 (N_27870,N_11524,N_16543);
nor U27871 (N_27871,N_18295,N_12279);
nor U27872 (N_27872,N_16905,N_16836);
xnor U27873 (N_27873,N_17434,N_11245);
and U27874 (N_27874,N_19384,N_11774);
nor U27875 (N_27875,N_10528,N_19233);
and U27876 (N_27876,N_11578,N_11237);
or U27877 (N_27877,N_17971,N_17531);
nor U27878 (N_27878,N_12847,N_15225);
or U27879 (N_27879,N_16670,N_12800);
nand U27880 (N_27880,N_16545,N_19947);
or U27881 (N_27881,N_18689,N_17197);
nand U27882 (N_27882,N_15570,N_14132);
and U27883 (N_27883,N_18577,N_18535);
or U27884 (N_27884,N_11219,N_13667);
nand U27885 (N_27885,N_13487,N_17480);
xnor U27886 (N_27886,N_17334,N_15009);
and U27887 (N_27887,N_15152,N_16275);
or U27888 (N_27888,N_15571,N_10709);
nand U27889 (N_27889,N_18586,N_12842);
or U27890 (N_27890,N_16198,N_14518);
or U27891 (N_27891,N_14349,N_12732);
xnor U27892 (N_27892,N_14468,N_17755);
or U27893 (N_27893,N_13546,N_17987);
nor U27894 (N_27894,N_15918,N_11483);
and U27895 (N_27895,N_14933,N_16384);
and U27896 (N_27896,N_14770,N_15586);
nor U27897 (N_27897,N_14972,N_18016);
nand U27898 (N_27898,N_15464,N_15465);
and U27899 (N_27899,N_11149,N_17762);
xor U27900 (N_27900,N_13936,N_15490);
nand U27901 (N_27901,N_17595,N_18187);
or U27902 (N_27902,N_11530,N_14104);
nor U27903 (N_27903,N_17327,N_18581);
nor U27904 (N_27904,N_12355,N_11701);
xor U27905 (N_27905,N_15825,N_10276);
nor U27906 (N_27906,N_15203,N_19346);
nor U27907 (N_27907,N_16664,N_16394);
nor U27908 (N_27908,N_12563,N_18132);
xor U27909 (N_27909,N_14676,N_11918);
or U27910 (N_27910,N_17987,N_12522);
xnor U27911 (N_27911,N_14254,N_11371);
and U27912 (N_27912,N_10067,N_18106);
or U27913 (N_27913,N_13519,N_10302);
or U27914 (N_27914,N_14434,N_18363);
nand U27915 (N_27915,N_19986,N_14290);
nand U27916 (N_27916,N_17755,N_13639);
nor U27917 (N_27917,N_11214,N_16556);
and U27918 (N_27918,N_12515,N_10371);
nand U27919 (N_27919,N_18074,N_19052);
or U27920 (N_27920,N_12083,N_11248);
or U27921 (N_27921,N_18616,N_13800);
or U27922 (N_27922,N_17370,N_16810);
nor U27923 (N_27923,N_17194,N_15687);
and U27924 (N_27924,N_12836,N_10218);
nor U27925 (N_27925,N_19957,N_17268);
nand U27926 (N_27926,N_15902,N_15683);
and U27927 (N_27927,N_17144,N_10560);
and U27928 (N_27928,N_12789,N_16577);
nand U27929 (N_27929,N_12322,N_17262);
nand U27930 (N_27930,N_12314,N_14767);
nand U27931 (N_27931,N_18324,N_19195);
nand U27932 (N_27932,N_13833,N_19931);
xor U27933 (N_27933,N_11119,N_19140);
and U27934 (N_27934,N_14638,N_17172);
or U27935 (N_27935,N_10757,N_11254);
nand U27936 (N_27936,N_11121,N_15476);
nand U27937 (N_27937,N_11019,N_17173);
xnor U27938 (N_27938,N_10498,N_18413);
nand U27939 (N_27939,N_19207,N_14333);
nand U27940 (N_27940,N_11710,N_18733);
or U27941 (N_27941,N_18792,N_10378);
and U27942 (N_27942,N_18503,N_14008);
nor U27943 (N_27943,N_15476,N_12717);
nand U27944 (N_27944,N_15810,N_13544);
nand U27945 (N_27945,N_13999,N_16285);
nand U27946 (N_27946,N_12209,N_10080);
and U27947 (N_27947,N_13448,N_19659);
xnor U27948 (N_27948,N_17943,N_13583);
or U27949 (N_27949,N_16122,N_16544);
nor U27950 (N_27950,N_10935,N_18915);
nand U27951 (N_27951,N_12757,N_15575);
xnor U27952 (N_27952,N_17718,N_16338);
and U27953 (N_27953,N_12451,N_18303);
nand U27954 (N_27954,N_17443,N_19864);
or U27955 (N_27955,N_15047,N_17416);
xor U27956 (N_27956,N_16599,N_15872);
nor U27957 (N_27957,N_19691,N_18432);
nor U27958 (N_27958,N_10068,N_19581);
and U27959 (N_27959,N_13334,N_17971);
or U27960 (N_27960,N_15316,N_18784);
nand U27961 (N_27961,N_15553,N_14687);
nand U27962 (N_27962,N_10502,N_13591);
nand U27963 (N_27963,N_13928,N_14426);
nor U27964 (N_27964,N_18880,N_18881);
or U27965 (N_27965,N_12428,N_11111);
nor U27966 (N_27966,N_17812,N_18828);
nor U27967 (N_27967,N_15106,N_17138);
and U27968 (N_27968,N_15291,N_14077);
and U27969 (N_27969,N_11855,N_16221);
xor U27970 (N_27970,N_17026,N_16142);
or U27971 (N_27971,N_12401,N_10579);
nor U27972 (N_27972,N_11350,N_14738);
or U27973 (N_27973,N_14314,N_18798);
or U27974 (N_27974,N_15061,N_17863);
or U27975 (N_27975,N_13719,N_13224);
xnor U27976 (N_27976,N_19090,N_14992);
and U27977 (N_27977,N_16803,N_19607);
nor U27978 (N_27978,N_14608,N_18071);
and U27979 (N_27979,N_16436,N_18994);
or U27980 (N_27980,N_15489,N_14470);
nand U27981 (N_27981,N_18624,N_12966);
nor U27982 (N_27982,N_15782,N_12029);
nand U27983 (N_27983,N_13274,N_17204);
nand U27984 (N_27984,N_15988,N_13907);
xor U27985 (N_27985,N_19815,N_18943);
nor U27986 (N_27986,N_11247,N_13539);
and U27987 (N_27987,N_12730,N_12233);
nor U27988 (N_27988,N_11074,N_11823);
or U27989 (N_27989,N_17298,N_19476);
or U27990 (N_27990,N_15779,N_16159);
nand U27991 (N_27991,N_18733,N_13882);
nor U27992 (N_27992,N_10076,N_11087);
or U27993 (N_27993,N_15299,N_19116);
nor U27994 (N_27994,N_11291,N_10729);
or U27995 (N_27995,N_17907,N_18104);
and U27996 (N_27996,N_13169,N_12023);
or U27997 (N_27997,N_19183,N_14148);
nand U27998 (N_27998,N_18515,N_13270);
nor U27999 (N_27999,N_15139,N_15823);
nor U28000 (N_28000,N_18087,N_18656);
nor U28001 (N_28001,N_19566,N_10986);
or U28002 (N_28002,N_11812,N_10368);
or U28003 (N_28003,N_11123,N_17959);
and U28004 (N_28004,N_11819,N_17324);
nand U28005 (N_28005,N_11882,N_10406);
nand U28006 (N_28006,N_14011,N_10725);
nand U28007 (N_28007,N_17260,N_16195);
xnor U28008 (N_28008,N_14845,N_18793);
or U28009 (N_28009,N_19543,N_12805);
nor U28010 (N_28010,N_18060,N_18428);
or U28011 (N_28011,N_19889,N_16369);
nor U28012 (N_28012,N_16247,N_19129);
nand U28013 (N_28013,N_16375,N_16768);
and U28014 (N_28014,N_15636,N_10193);
nand U28015 (N_28015,N_12110,N_14925);
xnor U28016 (N_28016,N_18866,N_15470);
xnor U28017 (N_28017,N_18630,N_13782);
and U28018 (N_28018,N_14050,N_14095);
and U28019 (N_28019,N_12466,N_18526);
nand U28020 (N_28020,N_10506,N_14168);
or U28021 (N_28021,N_15946,N_16768);
nor U28022 (N_28022,N_15729,N_19346);
nor U28023 (N_28023,N_16708,N_17646);
nand U28024 (N_28024,N_10732,N_10993);
or U28025 (N_28025,N_10749,N_18712);
and U28026 (N_28026,N_17758,N_18724);
xor U28027 (N_28027,N_14011,N_16725);
and U28028 (N_28028,N_19312,N_17891);
nor U28029 (N_28029,N_10535,N_12093);
nor U28030 (N_28030,N_12914,N_15341);
nand U28031 (N_28031,N_12092,N_19708);
or U28032 (N_28032,N_14867,N_13197);
nor U28033 (N_28033,N_16820,N_13211);
xor U28034 (N_28034,N_12567,N_12132);
nor U28035 (N_28035,N_14937,N_16643);
xor U28036 (N_28036,N_14875,N_15775);
xor U28037 (N_28037,N_17771,N_17023);
or U28038 (N_28038,N_18637,N_18422);
nand U28039 (N_28039,N_14173,N_19156);
nor U28040 (N_28040,N_13927,N_15655);
xnor U28041 (N_28041,N_15020,N_15111);
xor U28042 (N_28042,N_10024,N_16710);
nor U28043 (N_28043,N_17706,N_15037);
and U28044 (N_28044,N_18467,N_10029);
or U28045 (N_28045,N_11002,N_13425);
or U28046 (N_28046,N_12714,N_18807);
xnor U28047 (N_28047,N_17405,N_17931);
xor U28048 (N_28048,N_13802,N_10096);
and U28049 (N_28049,N_15124,N_13847);
nor U28050 (N_28050,N_18158,N_14256);
nand U28051 (N_28051,N_12071,N_10743);
nor U28052 (N_28052,N_14481,N_17433);
or U28053 (N_28053,N_15503,N_10727);
nor U28054 (N_28054,N_16156,N_18086);
and U28055 (N_28055,N_19714,N_14351);
and U28056 (N_28056,N_14993,N_11329);
nor U28057 (N_28057,N_17797,N_16608);
nor U28058 (N_28058,N_15904,N_10851);
nand U28059 (N_28059,N_12311,N_14032);
nand U28060 (N_28060,N_14753,N_19571);
nand U28061 (N_28061,N_16470,N_13120);
xnor U28062 (N_28062,N_13085,N_11508);
or U28063 (N_28063,N_10902,N_15048);
nand U28064 (N_28064,N_12083,N_17355);
nor U28065 (N_28065,N_17596,N_10289);
or U28066 (N_28066,N_14457,N_13837);
or U28067 (N_28067,N_14556,N_12346);
and U28068 (N_28068,N_15420,N_16892);
nor U28069 (N_28069,N_13817,N_16075);
nor U28070 (N_28070,N_17446,N_15594);
or U28071 (N_28071,N_14769,N_13897);
nor U28072 (N_28072,N_11676,N_18098);
nand U28073 (N_28073,N_12866,N_18063);
nor U28074 (N_28074,N_11859,N_12861);
nor U28075 (N_28075,N_15736,N_10218);
nor U28076 (N_28076,N_13233,N_13758);
nor U28077 (N_28077,N_13114,N_16036);
nor U28078 (N_28078,N_18797,N_18019);
or U28079 (N_28079,N_10455,N_11802);
nand U28080 (N_28080,N_16896,N_14844);
xnor U28081 (N_28081,N_17201,N_12563);
and U28082 (N_28082,N_10500,N_10171);
or U28083 (N_28083,N_19193,N_17154);
nand U28084 (N_28084,N_13962,N_15278);
nor U28085 (N_28085,N_11154,N_11821);
and U28086 (N_28086,N_11876,N_10288);
nand U28087 (N_28087,N_19594,N_13422);
nor U28088 (N_28088,N_19235,N_11400);
nor U28089 (N_28089,N_13780,N_15361);
nand U28090 (N_28090,N_17629,N_12158);
nand U28091 (N_28091,N_16685,N_11207);
xor U28092 (N_28092,N_12120,N_14286);
nand U28093 (N_28093,N_11902,N_16855);
nor U28094 (N_28094,N_13225,N_16444);
and U28095 (N_28095,N_13390,N_14792);
and U28096 (N_28096,N_19095,N_11332);
or U28097 (N_28097,N_12282,N_13309);
xor U28098 (N_28098,N_11097,N_12430);
nand U28099 (N_28099,N_14325,N_15362);
or U28100 (N_28100,N_18241,N_14060);
or U28101 (N_28101,N_14773,N_15948);
xor U28102 (N_28102,N_14328,N_14743);
nand U28103 (N_28103,N_17691,N_16325);
or U28104 (N_28104,N_16108,N_19850);
nand U28105 (N_28105,N_11020,N_17561);
xnor U28106 (N_28106,N_15321,N_13753);
nand U28107 (N_28107,N_13211,N_18091);
nand U28108 (N_28108,N_17115,N_19287);
nor U28109 (N_28109,N_14008,N_10920);
or U28110 (N_28110,N_13754,N_16554);
and U28111 (N_28111,N_12669,N_19343);
and U28112 (N_28112,N_18684,N_19736);
or U28113 (N_28113,N_10791,N_10089);
xnor U28114 (N_28114,N_18615,N_11933);
or U28115 (N_28115,N_17852,N_19550);
and U28116 (N_28116,N_11609,N_13709);
or U28117 (N_28117,N_14809,N_15656);
and U28118 (N_28118,N_13469,N_15438);
and U28119 (N_28119,N_17888,N_13488);
xnor U28120 (N_28120,N_12278,N_15572);
nand U28121 (N_28121,N_11386,N_19259);
xor U28122 (N_28122,N_18432,N_18668);
and U28123 (N_28123,N_16515,N_18766);
nor U28124 (N_28124,N_10533,N_13680);
nor U28125 (N_28125,N_16111,N_18092);
nor U28126 (N_28126,N_15655,N_18617);
and U28127 (N_28127,N_18305,N_14129);
and U28128 (N_28128,N_10411,N_19785);
nand U28129 (N_28129,N_16666,N_12189);
nand U28130 (N_28130,N_16683,N_17105);
xnor U28131 (N_28131,N_17483,N_13297);
nand U28132 (N_28132,N_16744,N_19393);
nand U28133 (N_28133,N_13715,N_18531);
nor U28134 (N_28134,N_10273,N_15352);
and U28135 (N_28135,N_17069,N_11435);
nor U28136 (N_28136,N_14466,N_11515);
xnor U28137 (N_28137,N_19250,N_18705);
nand U28138 (N_28138,N_19900,N_14838);
nand U28139 (N_28139,N_11630,N_17096);
or U28140 (N_28140,N_16438,N_14169);
nand U28141 (N_28141,N_13265,N_10485);
or U28142 (N_28142,N_13664,N_13006);
nor U28143 (N_28143,N_11342,N_18431);
nand U28144 (N_28144,N_14648,N_19248);
xnor U28145 (N_28145,N_11623,N_13432);
or U28146 (N_28146,N_13996,N_16898);
or U28147 (N_28147,N_18958,N_10433);
nor U28148 (N_28148,N_18835,N_11920);
nor U28149 (N_28149,N_12108,N_16056);
xnor U28150 (N_28150,N_17169,N_19103);
or U28151 (N_28151,N_14563,N_15874);
or U28152 (N_28152,N_12738,N_14389);
nor U28153 (N_28153,N_13499,N_11395);
nor U28154 (N_28154,N_18175,N_18644);
nand U28155 (N_28155,N_19178,N_19360);
nor U28156 (N_28156,N_12330,N_12455);
nor U28157 (N_28157,N_15045,N_10334);
nand U28158 (N_28158,N_14881,N_11471);
nor U28159 (N_28159,N_17294,N_10121);
or U28160 (N_28160,N_16815,N_13568);
and U28161 (N_28161,N_10435,N_17271);
or U28162 (N_28162,N_19068,N_18309);
xnor U28163 (N_28163,N_17817,N_10036);
xor U28164 (N_28164,N_10816,N_18112);
or U28165 (N_28165,N_15178,N_17913);
or U28166 (N_28166,N_11111,N_17759);
xnor U28167 (N_28167,N_11403,N_18176);
or U28168 (N_28168,N_10363,N_17918);
and U28169 (N_28169,N_16357,N_16072);
nand U28170 (N_28170,N_18200,N_15635);
or U28171 (N_28171,N_17032,N_16403);
or U28172 (N_28172,N_11115,N_19264);
and U28173 (N_28173,N_17792,N_17087);
or U28174 (N_28174,N_19730,N_10223);
and U28175 (N_28175,N_10732,N_14988);
or U28176 (N_28176,N_14819,N_15122);
or U28177 (N_28177,N_11593,N_13826);
xor U28178 (N_28178,N_10344,N_12791);
and U28179 (N_28179,N_15163,N_15319);
nor U28180 (N_28180,N_17085,N_17879);
nand U28181 (N_28181,N_10211,N_12749);
and U28182 (N_28182,N_16112,N_12722);
nand U28183 (N_28183,N_16353,N_18428);
and U28184 (N_28184,N_10573,N_16852);
xor U28185 (N_28185,N_14660,N_11295);
and U28186 (N_28186,N_16168,N_13870);
or U28187 (N_28187,N_12322,N_16201);
xor U28188 (N_28188,N_19161,N_17931);
nand U28189 (N_28189,N_18613,N_13366);
or U28190 (N_28190,N_17305,N_17375);
or U28191 (N_28191,N_15842,N_17386);
or U28192 (N_28192,N_12259,N_19047);
xor U28193 (N_28193,N_15104,N_12499);
nand U28194 (N_28194,N_13999,N_18021);
nand U28195 (N_28195,N_19476,N_17230);
nand U28196 (N_28196,N_16530,N_18306);
and U28197 (N_28197,N_19874,N_19270);
nand U28198 (N_28198,N_19360,N_15261);
or U28199 (N_28199,N_10919,N_12017);
and U28200 (N_28200,N_15468,N_19041);
or U28201 (N_28201,N_11578,N_17069);
nor U28202 (N_28202,N_15704,N_10126);
and U28203 (N_28203,N_16352,N_19620);
nand U28204 (N_28204,N_17007,N_17161);
and U28205 (N_28205,N_13439,N_14183);
nor U28206 (N_28206,N_19907,N_12392);
or U28207 (N_28207,N_11971,N_16756);
nand U28208 (N_28208,N_18643,N_18082);
and U28209 (N_28209,N_16745,N_17062);
and U28210 (N_28210,N_11203,N_19291);
nand U28211 (N_28211,N_15783,N_13202);
nand U28212 (N_28212,N_15506,N_15448);
or U28213 (N_28213,N_17418,N_17956);
xnor U28214 (N_28214,N_17490,N_18557);
nor U28215 (N_28215,N_19072,N_19085);
xor U28216 (N_28216,N_18961,N_10442);
xnor U28217 (N_28217,N_16115,N_12470);
xor U28218 (N_28218,N_15845,N_15531);
nor U28219 (N_28219,N_19621,N_10456);
xor U28220 (N_28220,N_17767,N_13495);
nand U28221 (N_28221,N_11873,N_12182);
and U28222 (N_28222,N_16661,N_19349);
and U28223 (N_28223,N_18868,N_17945);
or U28224 (N_28224,N_16823,N_10524);
and U28225 (N_28225,N_10379,N_14544);
xnor U28226 (N_28226,N_10876,N_14870);
nand U28227 (N_28227,N_10130,N_19042);
xnor U28228 (N_28228,N_10558,N_15611);
xor U28229 (N_28229,N_12515,N_14277);
nor U28230 (N_28230,N_12855,N_12064);
nand U28231 (N_28231,N_19684,N_18894);
and U28232 (N_28232,N_11388,N_15655);
xnor U28233 (N_28233,N_14040,N_17111);
and U28234 (N_28234,N_14931,N_17040);
and U28235 (N_28235,N_13787,N_14628);
nand U28236 (N_28236,N_17197,N_10076);
or U28237 (N_28237,N_18633,N_17060);
nor U28238 (N_28238,N_19261,N_19371);
nor U28239 (N_28239,N_15097,N_19429);
nand U28240 (N_28240,N_14072,N_18315);
xor U28241 (N_28241,N_14185,N_15326);
nand U28242 (N_28242,N_17805,N_15957);
nor U28243 (N_28243,N_13020,N_11283);
and U28244 (N_28244,N_11797,N_15671);
and U28245 (N_28245,N_11706,N_13704);
nand U28246 (N_28246,N_15870,N_19075);
nand U28247 (N_28247,N_11615,N_19384);
and U28248 (N_28248,N_13973,N_17965);
or U28249 (N_28249,N_16062,N_15199);
nand U28250 (N_28250,N_11372,N_16169);
nand U28251 (N_28251,N_14660,N_15158);
or U28252 (N_28252,N_11043,N_17261);
and U28253 (N_28253,N_10827,N_11714);
and U28254 (N_28254,N_10209,N_14022);
xnor U28255 (N_28255,N_15247,N_12586);
xnor U28256 (N_28256,N_18800,N_15193);
and U28257 (N_28257,N_19704,N_10475);
nand U28258 (N_28258,N_10523,N_18813);
nand U28259 (N_28259,N_17727,N_16695);
nor U28260 (N_28260,N_13842,N_16498);
or U28261 (N_28261,N_13697,N_13718);
nand U28262 (N_28262,N_18904,N_11227);
nand U28263 (N_28263,N_14521,N_19155);
and U28264 (N_28264,N_14404,N_18213);
nand U28265 (N_28265,N_16585,N_14915);
xnor U28266 (N_28266,N_12466,N_10093);
or U28267 (N_28267,N_18389,N_13895);
nor U28268 (N_28268,N_11264,N_19761);
or U28269 (N_28269,N_13144,N_14170);
nor U28270 (N_28270,N_11947,N_16323);
and U28271 (N_28271,N_18395,N_11112);
or U28272 (N_28272,N_10504,N_13839);
or U28273 (N_28273,N_10148,N_10225);
xor U28274 (N_28274,N_19000,N_12445);
or U28275 (N_28275,N_17370,N_12644);
and U28276 (N_28276,N_19354,N_19486);
xor U28277 (N_28277,N_13660,N_13542);
nand U28278 (N_28278,N_16299,N_11012);
and U28279 (N_28279,N_12010,N_14330);
nor U28280 (N_28280,N_17983,N_17257);
nor U28281 (N_28281,N_13417,N_11209);
nor U28282 (N_28282,N_11446,N_18873);
xnor U28283 (N_28283,N_16544,N_17655);
xnor U28284 (N_28284,N_18681,N_16883);
nor U28285 (N_28285,N_11497,N_19436);
or U28286 (N_28286,N_13436,N_15397);
nand U28287 (N_28287,N_14110,N_16222);
and U28288 (N_28288,N_10019,N_16316);
xor U28289 (N_28289,N_18492,N_16361);
nor U28290 (N_28290,N_11625,N_17578);
and U28291 (N_28291,N_11945,N_19114);
xnor U28292 (N_28292,N_13829,N_10143);
and U28293 (N_28293,N_13924,N_18578);
and U28294 (N_28294,N_14909,N_15535);
or U28295 (N_28295,N_19685,N_18060);
nor U28296 (N_28296,N_13654,N_17563);
nand U28297 (N_28297,N_19550,N_13712);
nor U28298 (N_28298,N_12277,N_17370);
xor U28299 (N_28299,N_19287,N_18381);
nor U28300 (N_28300,N_15919,N_18659);
nand U28301 (N_28301,N_10438,N_13187);
and U28302 (N_28302,N_11428,N_13515);
and U28303 (N_28303,N_15213,N_18540);
xnor U28304 (N_28304,N_12557,N_17064);
nand U28305 (N_28305,N_10323,N_17606);
xnor U28306 (N_28306,N_14022,N_16471);
and U28307 (N_28307,N_14129,N_16594);
and U28308 (N_28308,N_18222,N_14358);
nand U28309 (N_28309,N_10489,N_15894);
nor U28310 (N_28310,N_18965,N_15292);
or U28311 (N_28311,N_10749,N_12212);
nor U28312 (N_28312,N_14221,N_12143);
nor U28313 (N_28313,N_19803,N_11607);
xnor U28314 (N_28314,N_16582,N_10897);
and U28315 (N_28315,N_13086,N_13657);
xor U28316 (N_28316,N_19275,N_19528);
or U28317 (N_28317,N_10408,N_16434);
or U28318 (N_28318,N_12714,N_17414);
nor U28319 (N_28319,N_15690,N_13931);
or U28320 (N_28320,N_16975,N_14537);
xnor U28321 (N_28321,N_17245,N_17093);
and U28322 (N_28322,N_11191,N_17093);
and U28323 (N_28323,N_11069,N_10224);
or U28324 (N_28324,N_11434,N_19399);
nor U28325 (N_28325,N_12531,N_11625);
or U28326 (N_28326,N_15034,N_12415);
or U28327 (N_28327,N_18313,N_12160);
nand U28328 (N_28328,N_10672,N_19810);
and U28329 (N_28329,N_17597,N_12504);
and U28330 (N_28330,N_14131,N_16911);
xnor U28331 (N_28331,N_11487,N_18985);
or U28332 (N_28332,N_12878,N_13825);
nand U28333 (N_28333,N_14879,N_18288);
xor U28334 (N_28334,N_17567,N_12360);
xnor U28335 (N_28335,N_11485,N_14087);
and U28336 (N_28336,N_19886,N_16281);
nand U28337 (N_28337,N_11318,N_18642);
nor U28338 (N_28338,N_16147,N_11778);
and U28339 (N_28339,N_19861,N_17917);
nor U28340 (N_28340,N_15653,N_12532);
nand U28341 (N_28341,N_18718,N_19068);
nand U28342 (N_28342,N_11714,N_13216);
nand U28343 (N_28343,N_12834,N_12301);
nor U28344 (N_28344,N_15470,N_12833);
nor U28345 (N_28345,N_11414,N_19734);
nor U28346 (N_28346,N_15873,N_18393);
xor U28347 (N_28347,N_16973,N_10072);
nand U28348 (N_28348,N_11577,N_12291);
or U28349 (N_28349,N_15068,N_18516);
nand U28350 (N_28350,N_19627,N_13970);
xor U28351 (N_28351,N_18755,N_19333);
nand U28352 (N_28352,N_14559,N_16589);
or U28353 (N_28353,N_16874,N_12427);
nand U28354 (N_28354,N_14244,N_12277);
or U28355 (N_28355,N_15515,N_18628);
nor U28356 (N_28356,N_11409,N_11890);
nor U28357 (N_28357,N_19365,N_10033);
nor U28358 (N_28358,N_13855,N_17720);
or U28359 (N_28359,N_14821,N_12491);
nand U28360 (N_28360,N_19876,N_18180);
or U28361 (N_28361,N_11934,N_12542);
nand U28362 (N_28362,N_14120,N_16163);
nand U28363 (N_28363,N_17024,N_13513);
nand U28364 (N_28364,N_18821,N_12446);
nand U28365 (N_28365,N_16071,N_11814);
and U28366 (N_28366,N_11374,N_15382);
and U28367 (N_28367,N_14759,N_16479);
nor U28368 (N_28368,N_17401,N_17246);
nor U28369 (N_28369,N_15326,N_19391);
nor U28370 (N_28370,N_12528,N_10067);
nand U28371 (N_28371,N_11703,N_16466);
nor U28372 (N_28372,N_10046,N_11745);
or U28373 (N_28373,N_19495,N_19786);
nand U28374 (N_28374,N_15294,N_15018);
or U28375 (N_28375,N_15773,N_13775);
nor U28376 (N_28376,N_15502,N_15160);
xor U28377 (N_28377,N_19187,N_11660);
nand U28378 (N_28378,N_17766,N_14072);
nand U28379 (N_28379,N_12867,N_10266);
xor U28380 (N_28380,N_15223,N_19917);
nor U28381 (N_28381,N_13249,N_12294);
or U28382 (N_28382,N_17039,N_10736);
xnor U28383 (N_28383,N_15535,N_10371);
nor U28384 (N_28384,N_19281,N_14650);
and U28385 (N_28385,N_12734,N_15325);
xnor U28386 (N_28386,N_12206,N_18518);
nand U28387 (N_28387,N_18650,N_17144);
nor U28388 (N_28388,N_11582,N_17278);
nor U28389 (N_28389,N_16873,N_13989);
and U28390 (N_28390,N_12092,N_13971);
or U28391 (N_28391,N_16007,N_19394);
or U28392 (N_28392,N_19954,N_10049);
nor U28393 (N_28393,N_19615,N_16670);
nor U28394 (N_28394,N_16232,N_19272);
and U28395 (N_28395,N_15158,N_17557);
and U28396 (N_28396,N_10457,N_13126);
or U28397 (N_28397,N_19458,N_10743);
and U28398 (N_28398,N_17946,N_14179);
and U28399 (N_28399,N_15402,N_16208);
xnor U28400 (N_28400,N_16829,N_12379);
nand U28401 (N_28401,N_13295,N_16712);
or U28402 (N_28402,N_13539,N_14311);
or U28403 (N_28403,N_14746,N_16262);
or U28404 (N_28404,N_12822,N_16734);
and U28405 (N_28405,N_12651,N_10240);
and U28406 (N_28406,N_17719,N_13943);
or U28407 (N_28407,N_17631,N_15515);
or U28408 (N_28408,N_14465,N_16219);
nand U28409 (N_28409,N_11281,N_15739);
nand U28410 (N_28410,N_13243,N_13523);
or U28411 (N_28411,N_11473,N_15873);
or U28412 (N_28412,N_15673,N_10477);
xor U28413 (N_28413,N_12851,N_18593);
nor U28414 (N_28414,N_17520,N_10408);
nand U28415 (N_28415,N_12110,N_10533);
or U28416 (N_28416,N_12653,N_15322);
or U28417 (N_28417,N_17776,N_15444);
xor U28418 (N_28418,N_12211,N_12050);
nor U28419 (N_28419,N_19278,N_14556);
nand U28420 (N_28420,N_18764,N_11675);
nand U28421 (N_28421,N_11830,N_19973);
nand U28422 (N_28422,N_13598,N_13783);
nor U28423 (N_28423,N_16380,N_11049);
and U28424 (N_28424,N_15655,N_12385);
nand U28425 (N_28425,N_10296,N_17316);
or U28426 (N_28426,N_11765,N_15006);
or U28427 (N_28427,N_11528,N_19374);
xnor U28428 (N_28428,N_18412,N_12110);
or U28429 (N_28429,N_13471,N_16834);
and U28430 (N_28430,N_11886,N_10099);
nor U28431 (N_28431,N_17383,N_14871);
nand U28432 (N_28432,N_12854,N_19062);
nor U28433 (N_28433,N_15266,N_11143);
or U28434 (N_28434,N_15118,N_18357);
or U28435 (N_28435,N_19798,N_15179);
nand U28436 (N_28436,N_17295,N_19465);
nand U28437 (N_28437,N_11138,N_12142);
or U28438 (N_28438,N_18103,N_15546);
nor U28439 (N_28439,N_11938,N_14580);
nor U28440 (N_28440,N_14103,N_11184);
nand U28441 (N_28441,N_16674,N_14149);
and U28442 (N_28442,N_12258,N_10413);
and U28443 (N_28443,N_11860,N_14354);
nand U28444 (N_28444,N_11055,N_16371);
and U28445 (N_28445,N_14921,N_16502);
nand U28446 (N_28446,N_12352,N_12041);
nand U28447 (N_28447,N_10196,N_12370);
or U28448 (N_28448,N_11097,N_17787);
nor U28449 (N_28449,N_13053,N_17787);
or U28450 (N_28450,N_14743,N_14260);
and U28451 (N_28451,N_11391,N_12270);
nor U28452 (N_28452,N_14585,N_10998);
nand U28453 (N_28453,N_19121,N_19963);
or U28454 (N_28454,N_10717,N_16258);
and U28455 (N_28455,N_15881,N_14734);
xnor U28456 (N_28456,N_11281,N_13384);
nand U28457 (N_28457,N_11142,N_14739);
nand U28458 (N_28458,N_18882,N_11437);
and U28459 (N_28459,N_18347,N_18287);
nand U28460 (N_28460,N_15408,N_15351);
nor U28461 (N_28461,N_16307,N_17978);
or U28462 (N_28462,N_19020,N_10760);
xor U28463 (N_28463,N_13186,N_11709);
nand U28464 (N_28464,N_12092,N_10255);
and U28465 (N_28465,N_15015,N_17422);
nand U28466 (N_28466,N_14786,N_18954);
nand U28467 (N_28467,N_16485,N_19974);
and U28468 (N_28468,N_11548,N_13475);
and U28469 (N_28469,N_14184,N_11243);
nand U28470 (N_28470,N_11627,N_16141);
nand U28471 (N_28471,N_12807,N_18911);
or U28472 (N_28472,N_13045,N_16426);
or U28473 (N_28473,N_17155,N_10967);
nor U28474 (N_28474,N_12053,N_12535);
or U28475 (N_28475,N_19064,N_15999);
nand U28476 (N_28476,N_13235,N_17935);
and U28477 (N_28477,N_17222,N_18115);
nor U28478 (N_28478,N_13716,N_15525);
nand U28479 (N_28479,N_11294,N_13846);
nand U28480 (N_28480,N_18096,N_19539);
xnor U28481 (N_28481,N_17587,N_16732);
or U28482 (N_28482,N_18532,N_18343);
nor U28483 (N_28483,N_10741,N_12674);
or U28484 (N_28484,N_17568,N_19566);
xnor U28485 (N_28485,N_17832,N_16894);
nand U28486 (N_28486,N_12149,N_17117);
xor U28487 (N_28487,N_10290,N_11745);
nor U28488 (N_28488,N_18919,N_10858);
nand U28489 (N_28489,N_10164,N_10220);
xor U28490 (N_28490,N_19583,N_10423);
and U28491 (N_28491,N_10668,N_19232);
nor U28492 (N_28492,N_14003,N_11681);
xnor U28493 (N_28493,N_17079,N_11584);
xor U28494 (N_28494,N_18067,N_14291);
xnor U28495 (N_28495,N_17826,N_13241);
nand U28496 (N_28496,N_17474,N_15490);
nor U28497 (N_28497,N_13659,N_16397);
and U28498 (N_28498,N_17936,N_15962);
or U28499 (N_28499,N_18946,N_12256);
and U28500 (N_28500,N_15108,N_12406);
xnor U28501 (N_28501,N_11285,N_12569);
or U28502 (N_28502,N_10042,N_16250);
nand U28503 (N_28503,N_18124,N_19473);
nor U28504 (N_28504,N_18264,N_16128);
nand U28505 (N_28505,N_14886,N_13634);
or U28506 (N_28506,N_13113,N_11227);
or U28507 (N_28507,N_17976,N_18370);
nor U28508 (N_28508,N_12396,N_14013);
or U28509 (N_28509,N_10021,N_15062);
nor U28510 (N_28510,N_15975,N_12053);
nand U28511 (N_28511,N_10338,N_13122);
xor U28512 (N_28512,N_11872,N_14973);
nand U28513 (N_28513,N_18063,N_14861);
nand U28514 (N_28514,N_11434,N_10851);
nor U28515 (N_28515,N_15992,N_15075);
and U28516 (N_28516,N_18798,N_18472);
xnor U28517 (N_28517,N_12397,N_14701);
nor U28518 (N_28518,N_12115,N_18434);
or U28519 (N_28519,N_15657,N_13294);
nand U28520 (N_28520,N_11952,N_17899);
and U28521 (N_28521,N_13230,N_15126);
nor U28522 (N_28522,N_18043,N_17934);
nor U28523 (N_28523,N_18690,N_17560);
or U28524 (N_28524,N_18429,N_15064);
xnor U28525 (N_28525,N_16128,N_17695);
nor U28526 (N_28526,N_10211,N_18730);
nor U28527 (N_28527,N_15309,N_12542);
nand U28528 (N_28528,N_11353,N_15717);
or U28529 (N_28529,N_13884,N_17997);
and U28530 (N_28530,N_15996,N_14034);
or U28531 (N_28531,N_10962,N_13370);
xnor U28532 (N_28532,N_13439,N_11422);
nor U28533 (N_28533,N_17694,N_10180);
and U28534 (N_28534,N_13612,N_17177);
xnor U28535 (N_28535,N_18593,N_10865);
xnor U28536 (N_28536,N_15922,N_14336);
xnor U28537 (N_28537,N_11307,N_19256);
nor U28538 (N_28538,N_11866,N_12926);
xnor U28539 (N_28539,N_18124,N_15344);
or U28540 (N_28540,N_16141,N_14999);
and U28541 (N_28541,N_16547,N_13745);
xor U28542 (N_28542,N_19548,N_17421);
xor U28543 (N_28543,N_13023,N_18284);
xnor U28544 (N_28544,N_11806,N_18680);
nor U28545 (N_28545,N_10969,N_19917);
nand U28546 (N_28546,N_12278,N_19355);
nor U28547 (N_28547,N_12764,N_18073);
and U28548 (N_28548,N_12591,N_10613);
nand U28549 (N_28549,N_19768,N_10341);
nor U28550 (N_28550,N_17190,N_16080);
nand U28551 (N_28551,N_14934,N_16734);
or U28552 (N_28552,N_19084,N_10143);
nand U28553 (N_28553,N_11140,N_13958);
xnor U28554 (N_28554,N_17080,N_19793);
nand U28555 (N_28555,N_12949,N_19766);
nand U28556 (N_28556,N_10049,N_19735);
or U28557 (N_28557,N_12968,N_12413);
nand U28558 (N_28558,N_13321,N_13658);
or U28559 (N_28559,N_12750,N_12192);
and U28560 (N_28560,N_11565,N_11102);
nor U28561 (N_28561,N_15664,N_14514);
and U28562 (N_28562,N_11173,N_14150);
or U28563 (N_28563,N_10552,N_12668);
or U28564 (N_28564,N_12990,N_10058);
xor U28565 (N_28565,N_14052,N_13239);
nor U28566 (N_28566,N_18846,N_10996);
and U28567 (N_28567,N_19971,N_15817);
xnor U28568 (N_28568,N_16744,N_11994);
xor U28569 (N_28569,N_18252,N_19285);
and U28570 (N_28570,N_10576,N_10475);
nand U28571 (N_28571,N_13410,N_10930);
xnor U28572 (N_28572,N_16389,N_16132);
nand U28573 (N_28573,N_16795,N_18827);
nand U28574 (N_28574,N_13702,N_14005);
and U28575 (N_28575,N_10401,N_11414);
and U28576 (N_28576,N_16237,N_19300);
or U28577 (N_28577,N_14306,N_13326);
nand U28578 (N_28578,N_14695,N_15864);
nor U28579 (N_28579,N_10316,N_11175);
nand U28580 (N_28580,N_18503,N_10836);
nor U28581 (N_28581,N_15178,N_10761);
xor U28582 (N_28582,N_10214,N_12694);
and U28583 (N_28583,N_10984,N_14737);
nor U28584 (N_28584,N_11865,N_12810);
or U28585 (N_28585,N_10909,N_18697);
nor U28586 (N_28586,N_11913,N_16623);
nand U28587 (N_28587,N_17937,N_15338);
nor U28588 (N_28588,N_11389,N_19077);
nand U28589 (N_28589,N_17400,N_13151);
nor U28590 (N_28590,N_19539,N_10763);
nor U28591 (N_28591,N_17569,N_14689);
or U28592 (N_28592,N_12108,N_12145);
nand U28593 (N_28593,N_11846,N_17206);
xor U28594 (N_28594,N_16896,N_18667);
xnor U28595 (N_28595,N_15437,N_13822);
nand U28596 (N_28596,N_11135,N_19580);
or U28597 (N_28597,N_13123,N_18559);
or U28598 (N_28598,N_19367,N_10632);
and U28599 (N_28599,N_17476,N_11698);
nand U28600 (N_28600,N_15059,N_14099);
or U28601 (N_28601,N_10506,N_19939);
and U28602 (N_28602,N_15706,N_10915);
and U28603 (N_28603,N_15824,N_12948);
nor U28604 (N_28604,N_19005,N_10472);
xnor U28605 (N_28605,N_13588,N_10619);
nand U28606 (N_28606,N_15013,N_17875);
nor U28607 (N_28607,N_16054,N_14456);
or U28608 (N_28608,N_15890,N_18944);
nor U28609 (N_28609,N_11990,N_15003);
nand U28610 (N_28610,N_13441,N_15036);
nor U28611 (N_28611,N_13065,N_15019);
nand U28612 (N_28612,N_19087,N_11014);
xor U28613 (N_28613,N_17950,N_11002);
nor U28614 (N_28614,N_10051,N_13094);
and U28615 (N_28615,N_14900,N_17719);
xor U28616 (N_28616,N_15760,N_16781);
nand U28617 (N_28617,N_10923,N_13198);
xor U28618 (N_28618,N_15627,N_14621);
nor U28619 (N_28619,N_10320,N_14831);
nor U28620 (N_28620,N_17697,N_16868);
nand U28621 (N_28621,N_15393,N_17782);
nand U28622 (N_28622,N_19028,N_13189);
xnor U28623 (N_28623,N_19272,N_13832);
xor U28624 (N_28624,N_18954,N_11189);
or U28625 (N_28625,N_13292,N_15011);
nor U28626 (N_28626,N_13428,N_16971);
and U28627 (N_28627,N_18800,N_18544);
nand U28628 (N_28628,N_13245,N_16802);
or U28629 (N_28629,N_19109,N_14776);
or U28630 (N_28630,N_12219,N_18011);
or U28631 (N_28631,N_15110,N_18415);
nand U28632 (N_28632,N_12465,N_19789);
nand U28633 (N_28633,N_18611,N_17527);
xnor U28634 (N_28634,N_18427,N_13289);
and U28635 (N_28635,N_14578,N_13808);
and U28636 (N_28636,N_18821,N_11028);
nand U28637 (N_28637,N_18461,N_14882);
xnor U28638 (N_28638,N_19529,N_12344);
and U28639 (N_28639,N_18764,N_16313);
nor U28640 (N_28640,N_11176,N_14172);
xnor U28641 (N_28641,N_18210,N_14588);
nand U28642 (N_28642,N_11801,N_19762);
nand U28643 (N_28643,N_17339,N_15862);
nand U28644 (N_28644,N_14268,N_12465);
and U28645 (N_28645,N_11373,N_15983);
and U28646 (N_28646,N_14966,N_12210);
and U28647 (N_28647,N_16952,N_18086);
or U28648 (N_28648,N_13074,N_11778);
nor U28649 (N_28649,N_14243,N_15291);
nor U28650 (N_28650,N_10771,N_12153);
and U28651 (N_28651,N_14691,N_12694);
and U28652 (N_28652,N_17123,N_11868);
and U28653 (N_28653,N_12791,N_13638);
and U28654 (N_28654,N_10305,N_16748);
xor U28655 (N_28655,N_19950,N_12189);
nand U28656 (N_28656,N_14433,N_14619);
or U28657 (N_28657,N_14360,N_11005);
nand U28658 (N_28658,N_16761,N_11550);
xnor U28659 (N_28659,N_10557,N_19216);
xnor U28660 (N_28660,N_14805,N_15447);
xor U28661 (N_28661,N_15313,N_14276);
nor U28662 (N_28662,N_12452,N_12782);
and U28663 (N_28663,N_12270,N_16218);
nor U28664 (N_28664,N_13001,N_17940);
nand U28665 (N_28665,N_14901,N_10533);
and U28666 (N_28666,N_16860,N_13799);
and U28667 (N_28667,N_11272,N_13727);
nor U28668 (N_28668,N_17586,N_19040);
nor U28669 (N_28669,N_10272,N_18092);
or U28670 (N_28670,N_11417,N_16312);
and U28671 (N_28671,N_11887,N_10194);
and U28672 (N_28672,N_11056,N_11506);
and U28673 (N_28673,N_19539,N_18236);
nor U28674 (N_28674,N_16082,N_12639);
or U28675 (N_28675,N_10920,N_12497);
nand U28676 (N_28676,N_14704,N_15853);
and U28677 (N_28677,N_10068,N_13022);
nand U28678 (N_28678,N_15508,N_19477);
nor U28679 (N_28679,N_10601,N_19285);
xnor U28680 (N_28680,N_18718,N_13860);
nor U28681 (N_28681,N_15136,N_13171);
or U28682 (N_28682,N_14065,N_18511);
xnor U28683 (N_28683,N_19526,N_15528);
and U28684 (N_28684,N_19720,N_12711);
and U28685 (N_28685,N_13858,N_14713);
and U28686 (N_28686,N_10446,N_19080);
nor U28687 (N_28687,N_10074,N_11883);
nand U28688 (N_28688,N_13480,N_14711);
xor U28689 (N_28689,N_18125,N_15687);
and U28690 (N_28690,N_11637,N_13093);
nor U28691 (N_28691,N_19110,N_16166);
nand U28692 (N_28692,N_16390,N_19969);
nand U28693 (N_28693,N_19317,N_12916);
or U28694 (N_28694,N_19271,N_10291);
nor U28695 (N_28695,N_12453,N_19069);
xnor U28696 (N_28696,N_18694,N_17438);
nor U28697 (N_28697,N_15017,N_16659);
nand U28698 (N_28698,N_17606,N_12111);
and U28699 (N_28699,N_18569,N_17407);
or U28700 (N_28700,N_19797,N_19033);
and U28701 (N_28701,N_14114,N_15604);
xnor U28702 (N_28702,N_19596,N_14414);
and U28703 (N_28703,N_15600,N_13107);
xor U28704 (N_28704,N_11057,N_18532);
or U28705 (N_28705,N_12643,N_12329);
nand U28706 (N_28706,N_12490,N_12060);
nand U28707 (N_28707,N_16869,N_15065);
nor U28708 (N_28708,N_18642,N_10435);
nor U28709 (N_28709,N_13017,N_18863);
and U28710 (N_28710,N_19604,N_17759);
nor U28711 (N_28711,N_13193,N_13013);
nand U28712 (N_28712,N_10144,N_14723);
and U28713 (N_28713,N_15954,N_10885);
nand U28714 (N_28714,N_17756,N_13101);
nand U28715 (N_28715,N_15671,N_14117);
and U28716 (N_28716,N_19799,N_16380);
or U28717 (N_28717,N_18090,N_10929);
xnor U28718 (N_28718,N_12782,N_18011);
and U28719 (N_28719,N_15777,N_11229);
and U28720 (N_28720,N_11791,N_14053);
and U28721 (N_28721,N_14500,N_10559);
xor U28722 (N_28722,N_13256,N_16125);
and U28723 (N_28723,N_13352,N_15830);
or U28724 (N_28724,N_18209,N_11220);
nor U28725 (N_28725,N_18038,N_19913);
and U28726 (N_28726,N_17184,N_18282);
and U28727 (N_28727,N_11316,N_19872);
xnor U28728 (N_28728,N_10641,N_15084);
or U28729 (N_28729,N_15430,N_13056);
xnor U28730 (N_28730,N_19238,N_14899);
xor U28731 (N_28731,N_17897,N_15439);
nor U28732 (N_28732,N_14710,N_10766);
xnor U28733 (N_28733,N_11584,N_12139);
nor U28734 (N_28734,N_16797,N_12630);
xnor U28735 (N_28735,N_10798,N_12836);
or U28736 (N_28736,N_13444,N_13640);
xnor U28737 (N_28737,N_19153,N_19517);
and U28738 (N_28738,N_11755,N_11390);
xor U28739 (N_28739,N_10002,N_13490);
nand U28740 (N_28740,N_19804,N_14314);
xnor U28741 (N_28741,N_11291,N_11116);
nand U28742 (N_28742,N_11588,N_15105);
xor U28743 (N_28743,N_15805,N_11672);
xnor U28744 (N_28744,N_13802,N_11526);
nor U28745 (N_28745,N_11734,N_12286);
nor U28746 (N_28746,N_19780,N_19648);
and U28747 (N_28747,N_16061,N_16553);
nand U28748 (N_28748,N_11470,N_18052);
or U28749 (N_28749,N_18801,N_19602);
or U28750 (N_28750,N_15645,N_14611);
nand U28751 (N_28751,N_10819,N_16794);
xnor U28752 (N_28752,N_14341,N_15674);
nor U28753 (N_28753,N_16341,N_16121);
or U28754 (N_28754,N_16699,N_14502);
and U28755 (N_28755,N_17712,N_14894);
nor U28756 (N_28756,N_16455,N_17177);
nand U28757 (N_28757,N_16073,N_17559);
nand U28758 (N_28758,N_15337,N_17323);
xor U28759 (N_28759,N_17821,N_15988);
nor U28760 (N_28760,N_18945,N_13998);
or U28761 (N_28761,N_15431,N_13997);
nor U28762 (N_28762,N_13466,N_19292);
nand U28763 (N_28763,N_11460,N_16695);
and U28764 (N_28764,N_16716,N_17468);
nor U28765 (N_28765,N_18371,N_10110);
nor U28766 (N_28766,N_12537,N_11113);
xnor U28767 (N_28767,N_16786,N_11263);
or U28768 (N_28768,N_18654,N_18533);
xor U28769 (N_28769,N_18529,N_18111);
and U28770 (N_28770,N_14593,N_18857);
and U28771 (N_28771,N_15036,N_16480);
or U28772 (N_28772,N_16721,N_15545);
and U28773 (N_28773,N_18920,N_16150);
and U28774 (N_28774,N_17700,N_10008);
or U28775 (N_28775,N_11162,N_13104);
and U28776 (N_28776,N_17728,N_13521);
or U28777 (N_28777,N_19038,N_13271);
nor U28778 (N_28778,N_19247,N_17847);
xnor U28779 (N_28779,N_18307,N_14025);
nand U28780 (N_28780,N_15946,N_13070);
or U28781 (N_28781,N_10292,N_12047);
xnor U28782 (N_28782,N_10699,N_13763);
nor U28783 (N_28783,N_18779,N_12036);
or U28784 (N_28784,N_12322,N_14176);
or U28785 (N_28785,N_19849,N_14960);
nand U28786 (N_28786,N_15189,N_11495);
xnor U28787 (N_28787,N_19771,N_15990);
nor U28788 (N_28788,N_18686,N_16775);
and U28789 (N_28789,N_19374,N_18628);
nand U28790 (N_28790,N_16149,N_16035);
nand U28791 (N_28791,N_17404,N_10277);
nand U28792 (N_28792,N_14259,N_13667);
or U28793 (N_28793,N_17712,N_19750);
xor U28794 (N_28794,N_15867,N_11797);
and U28795 (N_28795,N_16665,N_12608);
nand U28796 (N_28796,N_11260,N_16419);
nand U28797 (N_28797,N_18306,N_16302);
nand U28798 (N_28798,N_17389,N_10703);
xnor U28799 (N_28799,N_18084,N_11124);
nand U28800 (N_28800,N_15971,N_19700);
and U28801 (N_28801,N_10478,N_18596);
nand U28802 (N_28802,N_18331,N_18985);
or U28803 (N_28803,N_15613,N_13606);
nand U28804 (N_28804,N_10500,N_15156);
xor U28805 (N_28805,N_12527,N_13933);
nand U28806 (N_28806,N_14417,N_15586);
and U28807 (N_28807,N_18320,N_18510);
xor U28808 (N_28808,N_19490,N_16811);
or U28809 (N_28809,N_17827,N_14265);
nor U28810 (N_28810,N_17075,N_15933);
or U28811 (N_28811,N_11375,N_17674);
xor U28812 (N_28812,N_18369,N_13610);
or U28813 (N_28813,N_17090,N_12211);
nand U28814 (N_28814,N_11927,N_18364);
xor U28815 (N_28815,N_16511,N_16745);
xnor U28816 (N_28816,N_12730,N_12100);
xor U28817 (N_28817,N_12691,N_16471);
and U28818 (N_28818,N_10610,N_12178);
nor U28819 (N_28819,N_11835,N_13451);
xnor U28820 (N_28820,N_10196,N_12692);
and U28821 (N_28821,N_18813,N_11055);
nand U28822 (N_28822,N_11919,N_15110);
nor U28823 (N_28823,N_13433,N_18466);
and U28824 (N_28824,N_17171,N_12804);
xor U28825 (N_28825,N_18504,N_14233);
and U28826 (N_28826,N_16612,N_18745);
nand U28827 (N_28827,N_18136,N_18704);
nand U28828 (N_28828,N_16547,N_19862);
nor U28829 (N_28829,N_11383,N_14143);
nor U28830 (N_28830,N_13787,N_12653);
nor U28831 (N_28831,N_15294,N_12690);
xor U28832 (N_28832,N_15345,N_19188);
nand U28833 (N_28833,N_11756,N_16291);
nand U28834 (N_28834,N_13065,N_13842);
nor U28835 (N_28835,N_12387,N_13769);
or U28836 (N_28836,N_19080,N_18225);
nand U28837 (N_28837,N_13984,N_12483);
xnor U28838 (N_28838,N_11615,N_12690);
or U28839 (N_28839,N_19312,N_10329);
and U28840 (N_28840,N_13016,N_12150);
xor U28841 (N_28841,N_18999,N_11796);
or U28842 (N_28842,N_15322,N_10785);
or U28843 (N_28843,N_17323,N_14384);
or U28844 (N_28844,N_19213,N_13664);
nor U28845 (N_28845,N_15407,N_17248);
or U28846 (N_28846,N_14570,N_19509);
and U28847 (N_28847,N_17520,N_11527);
and U28848 (N_28848,N_15871,N_14004);
nor U28849 (N_28849,N_14170,N_10664);
and U28850 (N_28850,N_17004,N_11528);
nand U28851 (N_28851,N_13277,N_15254);
nor U28852 (N_28852,N_15640,N_14768);
xor U28853 (N_28853,N_17678,N_10581);
nand U28854 (N_28854,N_14278,N_17630);
nor U28855 (N_28855,N_16018,N_12773);
or U28856 (N_28856,N_19957,N_11403);
or U28857 (N_28857,N_15410,N_14033);
xor U28858 (N_28858,N_19339,N_19055);
nor U28859 (N_28859,N_10927,N_12720);
and U28860 (N_28860,N_17806,N_11349);
nand U28861 (N_28861,N_10946,N_16253);
or U28862 (N_28862,N_14388,N_11814);
and U28863 (N_28863,N_10820,N_16662);
nor U28864 (N_28864,N_13205,N_13595);
and U28865 (N_28865,N_11254,N_17619);
or U28866 (N_28866,N_17024,N_19504);
nand U28867 (N_28867,N_10188,N_16294);
nor U28868 (N_28868,N_17276,N_16747);
xor U28869 (N_28869,N_16819,N_12298);
or U28870 (N_28870,N_19663,N_10860);
nor U28871 (N_28871,N_18920,N_12302);
nand U28872 (N_28872,N_17253,N_18681);
or U28873 (N_28873,N_16519,N_19599);
xnor U28874 (N_28874,N_11698,N_13236);
or U28875 (N_28875,N_11124,N_11896);
nand U28876 (N_28876,N_15668,N_10926);
nor U28877 (N_28877,N_11010,N_13398);
nor U28878 (N_28878,N_17861,N_18172);
nand U28879 (N_28879,N_12882,N_14764);
or U28880 (N_28880,N_14005,N_17111);
and U28881 (N_28881,N_13789,N_13807);
xor U28882 (N_28882,N_14654,N_12125);
nor U28883 (N_28883,N_17823,N_16815);
nand U28884 (N_28884,N_16354,N_15416);
and U28885 (N_28885,N_10287,N_13169);
nand U28886 (N_28886,N_17477,N_14161);
nand U28887 (N_28887,N_14598,N_19773);
or U28888 (N_28888,N_15564,N_13040);
or U28889 (N_28889,N_10762,N_18725);
nand U28890 (N_28890,N_13139,N_15409);
xor U28891 (N_28891,N_13788,N_15680);
or U28892 (N_28892,N_17927,N_10815);
nand U28893 (N_28893,N_16024,N_12614);
or U28894 (N_28894,N_13490,N_14056);
and U28895 (N_28895,N_17902,N_19022);
xor U28896 (N_28896,N_13623,N_19406);
nand U28897 (N_28897,N_14503,N_11380);
or U28898 (N_28898,N_13859,N_13536);
nand U28899 (N_28899,N_11595,N_19503);
and U28900 (N_28900,N_15583,N_11485);
xor U28901 (N_28901,N_17412,N_17072);
and U28902 (N_28902,N_16476,N_13794);
and U28903 (N_28903,N_14372,N_17593);
nand U28904 (N_28904,N_16519,N_17760);
or U28905 (N_28905,N_16378,N_12094);
xor U28906 (N_28906,N_17502,N_17940);
and U28907 (N_28907,N_11064,N_16870);
nor U28908 (N_28908,N_12278,N_17282);
xor U28909 (N_28909,N_12185,N_17403);
or U28910 (N_28910,N_13683,N_18652);
nand U28911 (N_28911,N_19467,N_16099);
nor U28912 (N_28912,N_17915,N_16161);
or U28913 (N_28913,N_15283,N_18912);
nand U28914 (N_28914,N_14454,N_14318);
nand U28915 (N_28915,N_15306,N_13715);
or U28916 (N_28916,N_16174,N_12439);
nand U28917 (N_28917,N_15258,N_14194);
xor U28918 (N_28918,N_17724,N_14361);
and U28919 (N_28919,N_13989,N_10198);
nor U28920 (N_28920,N_18651,N_10095);
or U28921 (N_28921,N_15837,N_17228);
nor U28922 (N_28922,N_16262,N_17863);
and U28923 (N_28923,N_18180,N_12428);
or U28924 (N_28924,N_15641,N_12703);
nand U28925 (N_28925,N_12772,N_14445);
nand U28926 (N_28926,N_12537,N_15922);
nor U28927 (N_28927,N_16781,N_13654);
and U28928 (N_28928,N_16704,N_18039);
and U28929 (N_28929,N_17705,N_15626);
xnor U28930 (N_28930,N_19821,N_16347);
xor U28931 (N_28931,N_14597,N_19722);
nand U28932 (N_28932,N_19167,N_15862);
nand U28933 (N_28933,N_18384,N_10120);
and U28934 (N_28934,N_15841,N_10266);
nand U28935 (N_28935,N_15162,N_13095);
and U28936 (N_28936,N_10898,N_12131);
nor U28937 (N_28937,N_17031,N_13116);
or U28938 (N_28938,N_17166,N_12988);
nand U28939 (N_28939,N_14731,N_19702);
nor U28940 (N_28940,N_13046,N_19112);
nor U28941 (N_28941,N_12326,N_17821);
or U28942 (N_28942,N_15812,N_13074);
nor U28943 (N_28943,N_16480,N_11624);
xor U28944 (N_28944,N_13097,N_16916);
nor U28945 (N_28945,N_11314,N_16829);
xnor U28946 (N_28946,N_16304,N_11287);
nor U28947 (N_28947,N_14574,N_10954);
or U28948 (N_28948,N_16149,N_18559);
nand U28949 (N_28949,N_13582,N_16883);
and U28950 (N_28950,N_13010,N_12561);
xnor U28951 (N_28951,N_18783,N_12450);
and U28952 (N_28952,N_17173,N_19235);
or U28953 (N_28953,N_10821,N_18378);
nor U28954 (N_28954,N_17181,N_18672);
or U28955 (N_28955,N_18700,N_12243);
xnor U28956 (N_28956,N_15649,N_17162);
nand U28957 (N_28957,N_15542,N_17694);
nor U28958 (N_28958,N_13863,N_12633);
xor U28959 (N_28959,N_18669,N_13379);
or U28960 (N_28960,N_12885,N_14642);
and U28961 (N_28961,N_13841,N_10763);
nor U28962 (N_28962,N_16076,N_16471);
or U28963 (N_28963,N_13872,N_11396);
and U28964 (N_28964,N_18905,N_16009);
xnor U28965 (N_28965,N_19964,N_17007);
or U28966 (N_28966,N_11836,N_13240);
or U28967 (N_28967,N_10137,N_14449);
xor U28968 (N_28968,N_15065,N_12934);
xor U28969 (N_28969,N_11305,N_10355);
and U28970 (N_28970,N_14215,N_17188);
nor U28971 (N_28971,N_13595,N_16671);
xor U28972 (N_28972,N_17999,N_19277);
nand U28973 (N_28973,N_10602,N_12520);
xor U28974 (N_28974,N_16238,N_16995);
and U28975 (N_28975,N_14117,N_11808);
or U28976 (N_28976,N_15641,N_12513);
nor U28977 (N_28977,N_16312,N_14333);
or U28978 (N_28978,N_17632,N_16382);
or U28979 (N_28979,N_11534,N_11555);
nand U28980 (N_28980,N_14979,N_18259);
nand U28981 (N_28981,N_12939,N_11339);
and U28982 (N_28982,N_19068,N_13879);
and U28983 (N_28983,N_13242,N_16571);
nor U28984 (N_28984,N_13023,N_15045);
nor U28985 (N_28985,N_10699,N_16028);
nor U28986 (N_28986,N_17696,N_15152);
or U28987 (N_28987,N_13850,N_15080);
or U28988 (N_28988,N_10519,N_10653);
xor U28989 (N_28989,N_19848,N_12127);
or U28990 (N_28990,N_19483,N_16857);
and U28991 (N_28991,N_12784,N_18298);
xnor U28992 (N_28992,N_18689,N_13905);
nor U28993 (N_28993,N_18282,N_17703);
nor U28994 (N_28994,N_19586,N_13158);
nand U28995 (N_28995,N_13057,N_19641);
and U28996 (N_28996,N_13630,N_12372);
xor U28997 (N_28997,N_11526,N_19861);
and U28998 (N_28998,N_19531,N_10503);
or U28999 (N_28999,N_16154,N_18117);
and U29000 (N_29000,N_10899,N_16434);
or U29001 (N_29001,N_11716,N_15455);
or U29002 (N_29002,N_13109,N_19923);
and U29003 (N_29003,N_10778,N_18464);
nand U29004 (N_29004,N_18633,N_19428);
nor U29005 (N_29005,N_17473,N_17125);
or U29006 (N_29006,N_13371,N_17477);
xor U29007 (N_29007,N_12316,N_12933);
xor U29008 (N_29008,N_10979,N_18574);
and U29009 (N_29009,N_12455,N_16483);
and U29010 (N_29010,N_10421,N_11849);
nor U29011 (N_29011,N_19120,N_13393);
or U29012 (N_29012,N_19145,N_14975);
or U29013 (N_29013,N_19344,N_14745);
or U29014 (N_29014,N_15198,N_14281);
and U29015 (N_29015,N_19994,N_16639);
nor U29016 (N_29016,N_15917,N_11707);
nand U29017 (N_29017,N_15469,N_19670);
xor U29018 (N_29018,N_17722,N_16536);
nor U29019 (N_29019,N_16250,N_18062);
nand U29020 (N_29020,N_11502,N_18643);
or U29021 (N_29021,N_11310,N_13453);
and U29022 (N_29022,N_11225,N_18743);
or U29023 (N_29023,N_18963,N_17714);
nor U29024 (N_29024,N_10520,N_15336);
xnor U29025 (N_29025,N_13226,N_18816);
and U29026 (N_29026,N_13310,N_17741);
xor U29027 (N_29027,N_10754,N_18310);
or U29028 (N_29028,N_15142,N_12856);
nand U29029 (N_29029,N_16355,N_17546);
nor U29030 (N_29030,N_15549,N_10778);
or U29031 (N_29031,N_12993,N_12851);
nand U29032 (N_29032,N_14891,N_17924);
or U29033 (N_29033,N_12325,N_17065);
and U29034 (N_29034,N_18320,N_15917);
and U29035 (N_29035,N_17495,N_11738);
or U29036 (N_29036,N_19672,N_19886);
nor U29037 (N_29037,N_14750,N_14845);
xor U29038 (N_29038,N_15386,N_15049);
and U29039 (N_29039,N_18136,N_11070);
or U29040 (N_29040,N_11418,N_16005);
and U29041 (N_29041,N_15749,N_19319);
nor U29042 (N_29042,N_17459,N_12590);
and U29043 (N_29043,N_19090,N_12164);
nand U29044 (N_29044,N_17799,N_17352);
and U29045 (N_29045,N_17793,N_14223);
nand U29046 (N_29046,N_15775,N_12912);
and U29047 (N_29047,N_11918,N_13050);
and U29048 (N_29048,N_15953,N_12537);
nor U29049 (N_29049,N_16244,N_10564);
and U29050 (N_29050,N_13029,N_12933);
xnor U29051 (N_29051,N_13584,N_17184);
nand U29052 (N_29052,N_11189,N_19302);
xor U29053 (N_29053,N_11555,N_18541);
or U29054 (N_29054,N_17088,N_10048);
xor U29055 (N_29055,N_19337,N_18003);
nand U29056 (N_29056,N_16632,N_10725);
and U29057 (N_29057,N_17582,N_18227);
nand U29058 (N_29058,N_14397,N_12479);
nor U29059 (N_29059,N_10208,N_17427);
nand U29060 (N_29060,N_17049,N_12229);
nand U29061 (N_29061,N_10173,N_15766);
xor U29062 (N_29062,N_12876,N_10951);
nor U29063 (N_29063,N_16712,N_16182);
or U29064 (N_29064,N_19372,N_10180);
nor U29065 (N_29065,N_13078,N_13359);
nor U29066 (N_29066,N_10151,N_13183);
or U29067 (N_29067,N_12370,N_11204);
and U29068 (N_29068,N_19386,N_19344);
xnor U29069 (N_29069,N_18349,N_12745);
and U29070 (N_29070,N_15239,N_13541);
nand U29071 (N_29071,N_19685,N_19713);
nor U29072 (N_29072,N_11696,N_13979);
xor U29073 (N_29073,N_11191,N_11461);
xor U29074 (N_29074,N_17943,N_10373);
nand U29075 (N_29075,N_17690,N_14349);
xor U29076 (N_29076,N_17901,N_14875);
nand U29077 (N_29077,N_15314,N_13432);
nand U29078 (N_29078,N_12106,N_11689);
xnor U29079 (N_29079,N_11903,N_11317);
or U29080 (N_29080,N_11488,N_10624);
nand U29081 (N_29081,N_18504,N_15959);
nor U29082 (N_29082,N_18588,N_10364);
and U29083 (N_29083,N_13678,N_14797);
nor U29084 (N_29084,N_10352,N_18213);
or U29085 (N_29085,N_18216,N_14646);
or U29086 (N_29086,N_10673,N_19481);
nor U29087 (N_29087,N_12987,N_12764);
xor U29088 (N_29088,N_12828,N_11068);
and U29089 (N_29089,N_15129,N_15396);
nand U29090 (N_29090,N_19548,N_13835);
and U29091 (N_29091,N_12263,N_12278);
or U29092 (N_29092,N_13282,N_19842);
xnor U29093 (N_29093,N_17099,N_11528);
nor U29094 (N_29094,N_12729,N_10978);
and U29095 (N_29095,N_12242,N_14891);
and U29096 (N_29096,N_19521,N_10839);
xor U29097 (N_29097,N_19698,N_10707);
xor U29098 (N_29098,N_12170,N_15563);
xor U29099 (N_29099,N_19197,N_16610);
and U29100 (N_29100,N_18998,N_15924);
nand U29101 (N_29101,N_18457,N_16772);
nor U29102 (N_29102,N_14427,N_15397);
or U29103 (N_29103,N_18599,N_15256);
and U29104 (N_29104,N_10193,N_14998);
and U29105 (N_29105,N_13345,N_15660);
nor U29106 (N_29106,N_12292,N_15629);
nand U29107 (N_29107,N_14258,N_12422);
and U29108 (N_29108,N_13474,N_12475);
or U29109 (N_29109,N_16528,N_12791);
nor U29110 (N_29110,N_11315,N_17355);
nor U29111 (N_29111,N_18089,N_16161);
nor U29112 (N_29112,N_12216,N_17275);
or U29113 (N_29113,N_13832,N_10413);
and U29114 (N_29114,N_18002,N_17051);
nand U29115 (N_29115,N_13430,N_15171);
xor U29116 (N_29116,N_10337,N_17676);
nor U29117 (N_29117,N_12786,N_13931);
and U29118 (N_29118,N_16107,N_12489);
nand U29119 (N_29119,N_13474,N_15421);
xnor U29120 (N_29120,N_12890,N_16607);
nand U29121 (N_29121,N_16318,N_18890);
nor U29122 (N_29122,N_18464,N_11283);
and U29123 (N_29123,N_17133,N_15048);
or U29124 (N_29124,N_13495,N_15751);
nor U29125 (N_29125,N_17868,N_17645);
nand U29126 (N_29126,N_13934,N_18792);
nand U29127 (N_29127,N_15907,N_13066);
and U29128 (N_29128,N_17132,N_10098);
and U29129 (N_29129,N_15552,N_14295);
nor U29130 (N_29130,N_18310,N_19963);
nor U29131 (N_29131,N_14487,N_19245);
or U29132 (N_29132,N_19441,N_10266);
and U29133 (N_29133,N_19312,N_16992);
xnor U29134 (N_29134,N_10306,N_19410);
or U29135 (N_29135,N_11176,N_11009);
or U29136 (N_29136,N_17096,N_12030);
nor U29137 (N_29137,N_18596,N_10857);
xnor U29138 (N_29138,N_18146,N_16355);
nor U29139 (N_29139,N_11450,N_10858);
nor U29140 (N_29140,N_10420,N_12972);
or U29141 (N_29141,N_12721,N_12297);
nand U29142 (N_29142,N_14370,N_13154);
xnor U29143 (N_29143,N_12338,N_11804);
or U29144 (N_29144,N_14928,N_19576);
nor U29145 (N_29145,N_11439,N_18340);
nand U29146 (N_29146,N_17225,N_12736);
nor U29147 (N_29147,N_14097,N_10992);
and U29148 (N_29148,N_13747,N_12778);
and U29149 (N_29149,N_16218,N_12677);
nand U29150 (N_29150,N_13326,N_11662);
xnor U29151 (N_29151,N_18580,N_10091);
nand U29152 (N_29152,N_10203,N_17049);
nor U29153 (N_29153,N_19390,N_18938);
nor U29154 (N_29154,N_17658,N_12555);
nor U29155 (N_29155,N_11788,N_12222);
nor U29156 (N_29156,N_17754,N_12239);
nand U29157 (N_29157,N_12094,N_13154);
or U29158 (N_29158,N_16074,N_14067);
nand U29159 (N_29159,N_19384,N_15373);
or U29160 (N_29160,N_11253,N_15433);
nand U29161 (N_29161,N_17470,N_19488);
nand U29162 (N_29162,N_10559,N_19950);
xnor U29163 (N_29163,N_15909,N_12261);
and U29164 (N_29164,N_19093,N_13496);
nand U29165 (N_29165,N_17899,N_11902);
nand U29166 (N_29166,N_12119,N_13955);
xor U29167 (N_29167,N_15485,N_16625);
or U29168 (N_29168,N_11097,N_11563);
nand U29169 (N_29169,N_12008,N_17255);
nand U29170 (N_29170,N_10432,N_15061);
nor U29171 (N_29171,N_13582,N_15862);
nor U29172 (N_29172,N_10342,N_19199);
and U29173 (N_29173,N_19759,N_19174);
or U29174 (N_29174,N_18550,N_17076);
or U29175 (N_29175,N_12360,N_11443);
and U29176 (N_29176,N_19862,N_18407);
or U29177 (N_29177,N_10887,N_14944);
or U29178 (N_29178,N_14926,N_11300);
nand U29179 (N_29179,N_10030,N_15287);
and U29180 (N_29180,N_14785,N_17187);
and U29181 (N_29181,N_17443,N_12950);
nand U29182 (N_29182,N_14256,N_14775);
nand U29183 (N_29183,N_13468,N_14258);
nor U29184 (N_29184,N_18649,N_10928);
nand U29185 (N_29185,N_16600,N_19690);
and U29186 (N_29186,N_13838,N_15121);
nor U29187 (N_29187,N_17287,N_11470);
xor U29188 (N_29188,N_18271,N_11517);
or U29189 (N_29189,N_13267,N_16957);
nor U29190 (N_29190,N_18476,N_13721);
or U29191 (N_29191,N_15249,N_14467);
or U29192 (N_29192,N_13818,N_14000);
nand U29193 (N_29193,N_14009,N_18350);
nand U29194 (N_29194,N_12237,N_12658);
xnor U29195 (N_29195,N_13379,N_11477);
xnor U29196 (N_29196,N_17530,N_18657);
and U29197 (N_29197,N_14216,N_15375);
xor U29198 (N_29198,N_10957,N_13099);
nand U29199 (N_29199,N_16994,N_16921);
and U29200 (N_29200,N_15469,N_15058);
or U29201 (N_29201,N_11229,N_19927);
and U29202 (N_29202,N_19538,N_12739);
xnor U29203 (N_29203,N_15963,N_14471);
or U29204 (N_29204,N_12959,N_18737);
nand U29205 (N_29205,N_16929,N_13723);
xor U29206 (N_29206,N_15333,N_14600);
nor U29207 (N_29207,N_14421,N_18433);
and U29208 (N_29208,N_12779,N_18433);
nor U29209 (N_29209,N_12790,N_13925);
nor U29210 (N_29210,N_15306,N_18718);
or U29211 (N_29211,N_12687,N_18745);
nand U29212 (N_29212,N_11630,N_16773);
or U29213 (N_29213,N_11252,N_12224);
and U29214 (N_29214,N_14292,N_17760);
or U29215 (N_29215,N_14986,N_17429);
xor U29216 (N_29216,N_17461,N_10797);
nor U29217 (N_29217,N_16816,N_15239);
xor U29218 (N_29218,N_17764,N_14979);
nor U29219 (N_29219,N_17295,N_10931);
xnor U29220 (N_29220,N_12826,N_16939);
nand U29221 (N_29221,N_14863,N_13479);
nor U29222 (N_29222,N_11650,N_18793);
and U29223 (N_29223,N_16946,N_10230);
and U29224 (N_29224,N_17866,N_11338);
xnor U29225 (N_29225,N_11803,N_12341);
xor U29226 (N_29226,N_18350,N_14452);
xnor U29227 (N_29227,N_19827,N_15273);
and U29228 (N_29228,N_18613,N_15082);
nand U29229 (N_29229,N_19387,N_10939);
nor U29230 (N_29230,N_14210,N_14705);
nor U29231 (N_29231,N_18936,N_13335);
or U29232 (N_29232,N_11682,N_19285);
nor U29233 (N_29233,N_14768,N_10170);
xor U29234 (N_29234,N_13945,N_15382);
xnor U29235 (N_29235,N_18947,N_17345);
xor U29236 (N_29236,N_11051,N_17620);
or U29237 (N_29237,N_15895,N_18277);
and U29238 (N_29238,N_17941,N_11449);
nand U29239 (N_29239,N_10160,N_12406);
or U29240 (N_29240,N_17551,N_19956);
nand U29241 (N_29241,N_19108,N_11994);
or U29242 (N_29242,N_16779,N_11652);
nor U29243 (N_29243,N_11793,N_17565);
nand U29244 (N_29244,N_10090,N_17882);
and U29245 (N_29245,N_13129,N_17822);
nand U29246 (N_29246,N_12974,N_11478);
and U29247 (N_29247,N_18130,N_15997);
nand U29248 (N_29248,N_17392,N_12258);
or U29249 (N_29249,N_14339,N_13954);
and U29250 (N_29250,N_16478,N_17172);
and U29251 (N_29251,N_17899,N_12264);
nand U29252 (N_29252,N_13109,N_12808);
nor U29253 (N_29253,N_13053,N_16445);
nor U29254 (N_29254,N_19714,N_15949);
xnor U29255 (N_29255,N_13135,N_18964);
xnor U29256 (N_29256,N_16549,N_11491);
and U29257 (N_29257,N_17404,N_16190);
nor U29258 (N_29258,N_14647,N_15717);
or U29259 (N_29259,N_14158,N_15777);
xnor U29260 (N_29260,N_13364,N_19902);
nor U29261 (N_29261,N_18208,N_16937);
and U29262 (N_29262,N_12968,N_11045);
and U29263 (N_29263,N_15832,N_14593);
and U29264 (N_29264,N_12195,N_11699);
nor U29265 (N_29265,N_19063,N_12845);
xor U29266 (N_29266,N_17630,N_13586);
xnor U29267 (N_29267,N_16374,N_11766);
and U29268 (N_29268,N_13692,N_18832);
xor U29269 (N_29269,N_13726,N_13845);
nor U29270 (N_29270,N_18571,N_16410);
nor U29271 (N_29271,N_11001,N_13009);
or U29272 (N_29272,N_17541,N_13389);
xor U29273 (N_29273,N_19870,N_16245);
xnor U29274 (N_29274,N_10548,N_12921);
nand U29275 (N_29275,N_15643,N_19937);
xnor U29276 (N_29276,N_19735,N_19343);
nand U29277 (N_29277,N_13365,N_12061);
nand U29278 (N_29278,N_10901,N_10220);
and U29279 (N_29279,N_13883,N_17776);
and U29280 (N_29280,N_14357,N_10241);
nand U29281 (N_29281,N_11450,N_10822);
nand U29282 (N_29282,N_10995,N_18190);
nor U29283 (N_29283,N_17700,N_12003);
or U29284 (N_29284,N_16716,N_15608);
nor U29285 (N_29285,N_17626,N_13876);
nand U29286 (N_29286,N_14803,N_18698);
or U29287 (N_29287,N_17457,N_11637);
xor U29288 (N_29288,N_15069,N_19894);
nor U29289 (N_29289,N_16005,N_15694);
xor U29290 (N_29290,N_13868,N_17150);
or U29291 (N_29291,N_17807,N_11063);
nor U29292 (N_29292,N_14527,N_16058);
and U29293 (N_29293,N_12140,N_18390);
nand U29294 (N_29294,N_13606,N_14068);
nand U29295 (N_29295,N_16445,N_14424);
nor U29296 (N_29296,N_16318,N_16828);
nor U29297 (N_29297,N_15510,N_15214);
and U29298 (N_29298,N_10195,N_16897);
nor U29299 (N_29299,N_15661,N_10525);
xor U29300 (N_29300,N_15485,N_12426);
nor U29301 (N_29301,N_12895,N_17026);
and U29302 (N_29302,N_18718,N_19129);
and U29303 (N_29303,N_18153,N_19484);
nor U29304 (N_29304,N_17875,N_15031);
or U29305 (N_29305,N_15798,N_16516);
or U29306 (N_29306,N_18095,N_15526);
nand U29307 (N_29307,N_11797,N_14509);
and U29308 (N_29308,N_15857,N_16045);
nand U29309 (N_29309,N_11999,N_11623);
nand U29310 (N_29310,N_14121,N_10452);
nand U29311 (N_29311,N_16038,N_18920);
xnor U29312 (N_29312,N_12644,N_13285);
xor U29313 (N_29313,N_16568,N_16411);
nand U29314 (N_29314,N_11347,N_18273);
xor U29315 (N_29315,N_18197,N_14620);
or U29316 (N_29316,N_11192,N_10636);
and U29317 (N_29317,N_19149,N_17796);
or U29318 (N_29318,N_10287,N_12522);
or U29319 (N_29319,N_18799,N_13293);
and U29320 (N_29320,N_19305,N_18286);
nor U29321 (N_29321,N_14555,N_18815);
and U29322 (N_29322,N_13276,N_13544);
nand U29323 (N_29323,N_13673,N_11019);
and U29324 (N_29324,N_12729,N_10080);
and U29325 (N_29325,N_13160,N_19866);
and U29326 (N_29326,N_19600,N_13424);
and U29327 (N_29327,N_12654,N_13536);
xor U29328 (N_29328,N_18147,N_10769);
xnor U29329 (N_29329,N_11817,N_12428);
nand U29330 (N_29330,N_18703,N_12040);
xor U29331 (N_29331,N_19196,N_18407);
xor U29332 (N_29332,N_17855,N_18118);
and U29333 (N_29333,N_18442,N_17778);
or U29334 (N_29334,N_13839,N_16647);
and U29335 (N_29335,N_12195,N_10798);
xnor U29336 (N_29336,N_19617,N_14199);
nand U29337 (N_29337,N_13153,N_12152);
xnor U29338 (N_29338,N_19649,N_15815);
nor U29339 (N_29339,N_15454,N_19482);
and U29340 (N_29340,N_10593,N_18813);
xor U29341 (N_29341,N_13568,N_14056);
and U29342 (N_29342,N_18812,N_12800);
nor U29343 (N_29343,N_17580,N_12416);
nor U29344 (N_29344,N_14668,N_17412);
and U29345 (N_29345,N_18178,N_17893);
and U29346 (N_29346,N_12574,N_17876);
nand U29347 (N_29347,N_11150,N_16098);
nand U29348 (N_29348,N_14988,N_13953);
nand U29349 (N_29349,N_10865,N_13298);
or U29350 (N_29350,N_12955,N_13021);
nand U29351 (N_29351,N_16188,N_15708);
and U29352 (N_29352,N_12472,N_11662);
and U29353 (N_29353,N_16016,N_17831);
nand U29354 (N_29354,N_19703,N_18495);
or U29355 (N_29355,N_19985,N_13202);
and U29356 (N_29356,N_10887,N_17503);
and U29357 (N_29357,N_11093,N_18991);
or U29358 (N_29358,N_15401,N_19960);
or U29359 (N_29359,N_10455,N_18997);
and U29360 (N_29360,N_11862,N_11634);
and U29361 (N_29361,N_12188,N_19073);
and U29362 (N_29362,N_15618,N_14577);
nand U29363 (N_29363,N_11760,N_18081);
xnor U29364 (N_29364,N_18146,N_12049);
xnor U29365 (N_29365,N_10315,N_11307);
nor U29366 (N_29366,N_15176,N_13065);
xnor U29367 (N_29367,N_11512,N_11035);
nand U29368 (N_29368,N_15075,N_14120);
and U29369 (N_29369,N_19961,N_16578);
xor U29370 (N_29370,N_13670,N_15687);
or U29371 (N_29371,N_13904,N_10825);
nor U29372 (N_29372,N_17758,N_16722);
or U29373 (N_29373,N_10388,N_11435);
or U29374 (N_29374,N_16884,N_13952);
or U29375 (N_29375,N_15023,N_16434);
nor U29376 (N_29376,N_19482,N_12217);
or U29377 (N_29377,N_15140,N_15390);
or U29378 (N_29378,N_13386,N_18518);
nor U29379 (N_29379,N_19831,N_19890);
xor U29380 (N_29380,N_10534,N_12996);
nand U29381 (N_29381,N_14567,N_14283);
nor U29382 (N_29382,N_14181,N_10255);
and U29383 (N_29383,N_19276,N_14333);
xnor U29384 (N_29384,N_10898,N_13896);
nand U29385 (N_29385,N_14168,N_19636);
xor U29386 (N_29386,N_16343,N_11656);
xnor U29387 (N_29387,N_15560,N_19156);
nor U29388 (N_29388,N_19182,N_11095);
or U29389 (N_29389,N_19361,N_19471);
and U29390 (N_29390,N_16835,N_10518);
and U29391 (N_29391,N_17393,N_13710);
nand U29392 (N_29392,N_18799,N_12564);
or U29393 (N_29393,N_10237,N_19686);
nor U29394 (N_29394,N_16141,N_18278);
nor U29395 (N_29395,N_18751,N_19895);
xnor U29396 (N_29396,N_10705,N_19122);
and U29397 (N_29397,N_14003,N_11348);
or U29398 (N_29398,N_14627,N_16851);
nand U29399 (N_29399,N_14156,N_10191);
and U29400 (N_29400,N_13211,N_14685);
xnor U29401 (N_29401,N_15149,N_14253);
or U29402 (N_29402,N_11348,N_12466);
xnor U29403 (N_29403,N_17925,N_19905);
xnor U29404 (N_29404,N_11701,N_12794);
and U29405 (N_29405,N_16941,N_13218);
xor U29406 (N_29406,N_16742,N_14530);
xnor U29407 (N_29407,N_10803,N_15522);
or U29408 (N_29408,N_19628,N_10048);
xnor U29409 (N_29409,N_16161,N_11210);
and U29410 (N_29410,N_17457,N_19081);
nor U29411 (N_29411,N_10844,N_13792);
and U29412 (N_29412,N_17596,N_11909);
nor U29413 (N_29413,N_19840,N_10660);
nor U29414 (N_29414,N_15192,N_18635);
xor U29415 (N_29415,N_13058,N_14198);
xnor U29416 (N_29416,N_13076,N_12045);
nor U29417 (N_29417,N_19129,N_14282);
or U29418 (N_29418,N_12520,N_12741);
nand U29419 (N_29419,N_11983,N_19143);
and U29420 (N_29420,N_14716,N_14547);
xnor U29421 (N_29421,N_13958,N_16869);
and U29422 (N_29422,N_16048,N_17279);
nand U29423 (N_29423,N_17316,N_14629);
xnor U29424 (N_29424,N_12198,N_13261);
or U29425 (N_29425,N_12325,N_10568);
or U29426 (N_29426,N_19044,N_14402);
nor U29427 (N_29427,N_11076,N_19113);
xor U29428 (N_29428,N_15147,N_17888);
or U29429 (N_29429,N_14534,N_11802);
nor U29430 (N_29430,N_14046,N_11919);
xor U29431 (N_29431,N_10018,N_15223);
and U29432 (N_29432,N_10831,N_14126);
or U29433 (N_29433,N_19242,N_16915);
nand U29434 (N_29434,N_11231,N_19507);
and U29435 (N_29435,N_15166,N_18377);
nor U29436 (N_29436,N_11083,N_13491);
nor U29437 (N_29437,N_11711,N_11668);
nand U29438 (N_29438,N_19695,N_13199);
xor U29439 (N_29439,N_17850,N_13158);
and U29440 (N_29440,N_15500,N_19500);
nand U29441 (N_29441,N_11940,N_18517);
nor U29442 (N_29442,N_14763,N_13543);
and U29443 (N_29443,N_17554,N_10114);
nor U29444 (N_29444,N_16315,N_10825);
and U29445 (N_29445,N_10618,N_10368);
nand U29446 (N_29446,N_14480,N_12325);
nand U29447 (N_29447,N_10585,N_10061);
and U29448 (N_29448,N_12085,N_13135);
nand U29449 (N_29449,N_17451,N_18722);
xnor U29450 (N_29450,N_15024,N_14604);
or U29451 (N_29451,N_11115,N_16437);
nor U29452 (N_29452,N_10115,N_12658);
or U29453 (N_29453,N_16719,N_11475);
xnor U29454 (N_29454,N_14713,N_18022);
and U29455 (N_29455,N_19470,N_12405);
xor U29456 (N_29456,N_10439,N_10923);
xnor U29457 (N_29457,N_16958,N_10445);
or U29458 (N_29458,N_15199,N_11029);
and U29459 (N_29459,N_16013,N_12619);
nor U29460 (N_29460,N_13752,N_15049);
nor U29461 (N_29461,N_16315,N_10999);
or U29462 (N_29462,N_14715,N_16944);
nor U29463 (N_29463,N_13363,N_16936);
nand U29464 (N_29464,N_13783,N_18610);
xnor U29465 (N_29465,N_15052,N_11564);
or U29466 (N_29466,N_12311,N_13419);
nor U29467 (N_29467,N_15931,N_17373);
nand U29468 (N_29468,N_11936,N_18123);
and U29469 (N_29469,N_10402,N_19432);
and U29470 (N_29470,N_12803,N_19730);
and U29471 (N_29471,N_14877,N_18951);
nand U29472 (N_29472,N_15870,N_18131);
nor U29473 (N_29473,N_10535,N_13090);
xnor U29474 (N_29474,N_14331,N_19839);
or U29475 (N_29475,N_19720,N_16258);
nand U29476 (N_29476,N_13504,N_19514);
nor U29477 (N_29477,N_12942,N_16094);
and U29478 (N_29478,N_18375,N_10288);
xnor U29479 (N_29479,N_11854,N_19919);
xor U29480 (N_29480,N_13290,N_16604);
xnor U29481 (N_29481,N_17420,N_16709);
or U29482 (N_29482,N_15670,N_18634);
xor U29483 (N_29483,N_10566,N_18818);
nor U29484 (N_29484,N_16823,N_10995);
and U29485 (N_29485,N_17655,N_17980);
nand U29486 (N_29486,N_17437,N_16574);
xor U29487 (N_29487,N_10586,N_18537);
nor U29488 (N_29488,N_11831,N_17866);
nand U29489 (N_29489,N_17531,N_14817);
and U29490 (N_29490,N_19255,N_14421);
xor U29491 (N_29491,N_12174,N_13640);
nand U29492 (N_29492,N_10323,N_14627);
or U29493 (N_29493,N_12081,N_17666);
and U29494 (N_29494,N_15814,N_18636);
or U29495 (N_29495,N_11945,N_15343);
and U29496 (N_29496,N_14759,N_12605);
nor U29497 (N_29497,N_10079,N_10737);
xor U29498 (N_29498,N_14093,N_14652);
and U29499 (N_29499,N_15345,N_15536);
nand U29500 (N_29500,N_14154,N_10993);
xnor U29501 (N_29501,N_12469,N_19344);
and U29502 (N_29502,N_18493,N_13943);
nor U29503 (N_29503,N_15999,N_14977);
nand U29504 (N_29504,N_19880,N_16359);
xor U29505 (N_29505,N_11830,N_19346);
nand U29506 (N_29506,N_15924,N_10042);
nand U29507 (N_29507,N_12401,N_17681);
xor U29508 (N_29508,N_10128,N_16241);
or U29509 (N_29509,N_15635,N_14367);
and U29510 (N_29510,N_14131,N_18145);
or U29511 (N_29511,N_16056,N_16793);
and U29512 (N_29512,N_10037,N_19647);
nand U29513 (N_29513,N_19472,N_12096);
or U29514 (N_29514,N_16193,N_17181);
or U29515 (N_29515,N_13234,N_19163);
xor U29516 (N_29516,N_11636,N_12933);
nand U29517 (N_29517,N_19071,N_11242);
nand U29518 (N_29518,N_18559,N_17225);
and U29519 (N_29519,N_10409,N_17353);
and U29520 (N_29520,N_18642,N_14398);
nor U29521 (N_29521,N_19115,N_15302);
xnor U29522 (N_29522,N_10798,N_19158);
nand U29523 (N_29523,N_10541,N_17125);
or U29524 (N_29524,N_15538,N_16808);
and U29525 (N_29525,N_13664,N_12854);
nor U29526 (N_29526,N_10215,N_18451);
and U29527 (N_29527,N_11060,N_18117);
or U29528 (N_29528,N_17151,N_13483);
xor U29529 (N_29529,N_10375,N_13564);
and U29530 (N_29530,N_10399,N_19977);
nand U29531 (N_29531,N_11967,N_10635);
xor U29532 (N_29532,N_14447,N_19632);
nor U29533 (N_29533,N_13195,N_10078);
nand U29534 (N_29534,N_15862,N_18194);
or U29535 (N_29535,N_19153,N_13135);
and U29536 (N_29536,N_12320,N_12065);
nand U29537 (N_29537,N_16188,N_16759);
or U29538 (N_29538,N_12851,N_14040);
nor U29539 (N_29539,N_12193,N_10413);
nor U29540 (N_29540,N_19253,N_17164);
nand U29541 (N_29541,N_11749,N_17344);
or U29542 (N_29542,N_16645,N_11451);
and U29543 (N_29543,N_13817,N_11770);
xnor U29544 (N_29544,N_16555,N_17297);
nor U29545 (N_29545,N_12399,N_18551);
nand U29546 (N_29546,N_14762,N_16227);
and U29547 (N_29547,N_19923,N_17033);
or U29548 (N_29548,N_19153,N_10680);
xnor U29549 (N_29549,N_12665,N_13553);
and U29550 (N_29550,N_12051,N_14364);
nor U29551 (N_29551,N_16749,N_17028);
or U29552 (N_29552,N_19136,N_19186);
and U29553 (N_29553,N_13699,N_16931);
and U29554 (N_29554,N_10985,N_16075);
nor U29555 (N_29555,N_17123,N_18379);
and U29556 (N_29556,N_18509,N_18838);
nand U29557 (N_29557,N_13810,N_16332);
xor U29558 (N_29558,N_13540,N_14359);
nand U29559 (N_29559,N_15536,N_13331);
nand U29560 (N_29560,N_12119,N_13688);
and U29561 (N_29561,N_16496,N_14658);
nand U29562 (N_29562,N_16763,N_17189);
nor U29563 (N_29563,N_18785,N_17953);
nor U29564 (N_29564,N_10359,N_14258);
nor U29565 (N_29565,N_14980,N_14876);
nor U29566 (N_29566,N_10992,N_19371);
and U29567 (N_29567,N_12819,N_19275);
nor U29568 (N_29568,N_10718,N_15352);
nand U29569 (N_29569,N_15791,N_12448);
or U29570 (N_29570,N_17082,N_17915);
or U29571 (N_29571,N_19485,N_17262);
nand U29572 (N_29572,N_14830,N_14099);
xor U29573 (N_29573,N_16802,N_11015);
xor U29574 (N_29574,N_14106,N_14678);
xnor U29575 (N_29575,N_15469,N_17181);
or U29576 (N_29576,N_14318,N_14223);
or U29577 (N_29577,N_14884,N_15125);
nand U29578 (N_29578,N_10853,N_12493);
or U29579 (N_29579,N_18440,N_16652);
xnor U29580 (N_29580,N_17331,N_19554);
nor U29581 (N_29581,N_15665,N_13604);
and U29582 (N_29582,N_18347,N_19670);
or U29583 (N_29583,N_18231,N_12780);
xnor U29584 (N_29584,N_16722,N_14417);
or U29585 (N_29585,N_15747,N_15315);
xor U29586 (N_29586,N_16679,N_15354);
and U29587 (N_29587,N_17850,N_13055);
nor U29588 (N_29588,N_11640,N_10966);
and U29589 (N_29589,N_15816,N_11658);
nand U29590 (N_29590,N_19109,N_17621);
nor U29591 (N_29591,N_12287,N_14127);
nor U29592 (N_29592,N_15758,N_13890);
and U29593 (N_29593,N_16324,N_16252);
xnor U29594 (N_29594,N_16549,N_14778);
nor U29595 (N_29595,N_11978,N_10386);
nand U29596 (N_29596,N_11705,N_12001);
and U29597 (N_29597,N_14995,N_11497);
xnor U29598 (N_29598,N_14503,N_18631);
xnor U29599 (N_29599,N_18069,N_14737);
nand U29600 (N_29600,N_13360,N_13757);
or U29601 (N_29601,N_15612,N_16940);
and U29602 (N_29602,N_12145,N_12570);
and U29603 (N_29603,N_18957,N_14947);
or U29604 (N_29604,N_14904,N_13802);
nand U29605 (N_29605,N_11679,N_14263);
or U29606 (N_29606,N_12803,N_19506);
or U29607 (N_29607,N_16622,N_12839);
nand U29608 (N_29608,N_17683,N_18185);
or U29609 (N_29609,N_16879,N_12637);
xor U29610 (N_29610,N_13503,N_10015);
nor U29611 (N_29611,N_10062,N_15314);
nor U29612 (N_29612,N_17254,N_11425);
nand U29613 (N_29613,N_11739,N_18001);
xnor U29614 (N_29614,N_19278,N_18327);
xnor U29615 (N_29615,N_12664,N_12907);
xnor U29616 (N_29616,N_10178,N_11194);
and U29617 (N_29617,N_10250,N_15999);
xnor U29618 (N_29618,N_16520,N_16948);
and U29619 (N_29619,N_16713,N_13519);
or U29620 (N_29620,N_15163,N_11371);
nand U29621 (N_29621,N_16010,N_11640);
and U29622 (N_29622,N_19127,N_12903);
nor U29623 (N_29623,N_18318,N_11861);
nor U29624 (N_29624,N_19837,N_15965);
nand U29625 (N_29625,N_16625,N_13021);
xor U29626 (N_29626,N_15363,N_18647);
and U29627 (N_29627,N_15048,N_15761);
nor U29628 (N_29628,N_13875,N_18652);
nand U29629 (N_29629,N_10205,N_16090);
nor U29630 (N_29630,N_12583,N_17048);
xor U29631 (N_29631,N_12699,N_11835);
nand U29632 (N_29632,N_19453,N_12737);
nand U29633 (N_29633,N_19338,N_17457);
nand U29634 (N_29634,N_11144,N_19173);
or U29635 (N_29635,N_19583,N_19693);
or U29636 (N_29636,N_16423,N_19108);
or U29637 (N_29637,N_11341,N_14463);
or U29638 (N_29638,N_15547,N_18539);
or U29639 (N_29639,N_15645,N_11529);
nor U29640 (N_29640,N_19270,N_18074);
and U29641 (N_29641,N_12956,N_14056);
nor U29642 (N_29642,N_17202,N_18688);
nor U29643 (N_29643,N_13275,N_11984);
nand U29644 (N_29644,N_19834,N_15867);
nand U29645 (N_29645,N_14774,N_12287);
or U29646 (N_29646,N_13446,N_14697);
xor U29647 (N_29647,N_15719,N_14745);
xor U29648 (N_29648,N_12907,N_13533);
nand U29649 (N_29649,N_12246,N_10630);
or U29650 (N_29650,N_14282,N_16637);
xor U29651 (N_29651,N_17196,N_19571);
and U29652 (N_29652,N_10853,N_15324);
xnor U29653 (N_29653,N_18288,N_13980);
and U29654 (N_29654,N_14691,N_14520);
or U29655 (N_29655,N_15340,N_14703);
nand U29656 (N_29656,N_13457,N_17635);
nand U29657 (N_29657,N_15693,N_12611);
or U29658 (N_29658,N_12380,N_14733);
and U29659 (N_29659,N_18486,N_11524);
nor U29660 (N_29660,N_11974,N_11902);
and U29661 (N_29661,N_12517,N_10365);
and U29662 (N_29662,N_18471,N_14346);
nand U29663 (N_29663,N_12436,N_18821);
or U29664 (N_29664,N_18392,N_19161);
nor U29665 (N_29665,N_16585,N_17565);
and U29666 (N_29666,N_15824,N_10852);
or U29667 (N_29667,N_10493,N_18704);
nor U29668 (N_29668,N_11666,N_17974);
and U29669 (N_29669,N_19181,N_18425);
and U29670 (N_29670,N_10038,N_10379);
or U29671 (N_29671,N_16767,N_14720);
xor U29672 (N_29672,N_11001,N_10033);
or U29673 (N_29673,N_10810,N_13922);
or U29674 (N_29674,N_15889,N_11675);
or U29675 (N_29675,N_12286,N_12413);
and U29676 (N_29676,N_17647,N_19793);
nand U29677 (N_29677,N_12436,N_13733);
nand U29678 (N_29678,N_19766,N_17314);
nor U29679 (N_29679,N_11465,N_14577);
xnor U29680 (N_29680,N_11349,N_14198);
xnor U29681 (N_29681,N_12363,N_17924);
nand U29682 (N_29682,N_12910,N_18357);
and U29683 (N_29683,N_12906,N_17085);
or U29684 (N_29684,N_17836,N_14622);
nor U29685 (N_29685,N_18665,N_16605);
or U29686 (N_29686,N_15793,N_19941);
or U29687 (N_29687,N_11881,N_12639);
xor U29688 (N_29688,N_19781,N_10508);
nor U29689 (N_29689,N_13220,N_12330);
nand U29690 (N_29690,N_19218,N_11320);
nor U29691 (N_29691,N_13937,N_11705);
nand U29692 (N_29692,N_16422,N_16099);
or U29693 (N_29693,N_16067,N_16604);
nand U29694 (N_29694,N_12882,N_15248);
nand U29695 (N_29695,N_12289,N_15512);
and U29696 (N_29696,N_12047,N_13234);
nor U29697 (N_29697,N_16120,N_12876);
nor U29698 (N_29698,N_19058,N_15864);
or U29699 (N_29699,N_11356,N_16970);
or U29700 (N_29700,N_14890,N_10881);
nor U29701 (N_29701,N_12486,N_10775);
xor U29702 (N_29702,N_10961,N_15494);
nand U29703 (N_29703,N_12574,N_13439);
nor U29704 (N_29704,N_14060,N_18096);
xor U29705 (N_29705,N_15379,N_12638);
and U29706 (N_29706,N_14589,N_14926);
xor U29707 (N_29707,N_19721,N_10874);
and U29708 (N_29708,N_11827,N_10075);
xor U29709 (N_29709,N_16102,N_10985);
nand U29710 (N_29710,N_11256,N_15699);
xnor U29711 (N_29711,N_15921,N_17105);
and U29712 (N_29712,N_15668,N_19684);
nor U29713 (N_29713,N_15026,N_18305);
xnor U29714 (N_29714,N_15650,N_17097);
and U29715 (N_29715,N_10392,N_15944);
nand U29716 (N_29716,N_15245,N_18603);
and U29717 (N_29717,N_16918,N_15319);
or U29718 (N_29718,N_11590,N_10308);
or U29719 (N_29719,N_13077,N_17049);
or U29720 (N_29720,N_19036,N_10262);
xor U29721 (N_29721,N_19179,N_16318);
nand U29722 (N_29722,N_11729,N_10760);
xnor U29723 (N_29723,N_11186,N_18509);
xor U29724 (N_29724,N_19176,N_14532);
nand U29725 (N_29725,N_13121,N_15147);
nand U29726 (N_29726,N_15112,N_14947);
nor U29727 (N_29727,N_15774,N_17674);
nand U29728 (N_29728,N_19707,N_15612);
nor U29729 (N_29729,N_18597,N_14878);
nor U29730 (N_29730,N_11270,N_15921);
nor U29731 (N_29731,N_18862,N_13256);
nand U29732 (N_29732,N_13734,N_15705);
or U29733 (N_29733,N_15451,N_12020);
xnor U29734 (N_29734,N_13341,N_14405);
or U29735 (N_29735,N_17859,N_12816);
and U29736 (N_29736,N_11845,N_17498);
xnor U29737 (N_29737,N_19263,N_19844);
nand U29738 (N_29738,N_12901,N_16004);
or U29739 (N_29739,N_14269,N_17959);
nor U29740 (N_29740,N_18638,N_11437);
or U29741 (N_29741,N_15674,N_17717);
and U29742 (N_29742,N_15778,N_15739);
and U29743 (N_29743,N_13256,N_18937);
and U29744 (N_29744,N_14988,N_18602);
and U29745 (N_29745,N_18153,N_13375);
nor U29746 (N_29746,N_11442,N_12782);
nand U29747 (N_29747,N_17680,N_13599);
nand U29748 (N_29748,N_17878,N_13770);
nor U29749 (N_29749,N_11615,N_13827);
or U29750 (N_29750,N_14058,N_16221);
or U29751 (N_29751,N_16585,N_10165);
nand U29752 (N_29752,N_12563,N_10209);
xnor U29753 (N_29753,N_15453,N_16789);
xnor U29754 (N_29754,N_13456,N_19118);
and U29755 (N_29755,N_16429,N_16411);
nor U29756 (N_29756,N_17118,N_13383);
or U29757 (N_29757,N_17080,N_17799);
nor U29758 (N_29758,N_15040,N_10816);
nor U29759 (N_29759,N_12180,N_16360);
and U29760 (N_29760,N_18416,N_17083);
and U29761 (N_29761,N_12623,N_17786);
xnor U29762 (N_29762,N_18397,N_10051);
nor U29763 (N_29763,N_11218,N_15123);
or U29764 (N_29764,N_13772,N_12212);
xnor U29765 (N_29765,N_14013,N_13622);
nand U29766 (N_29766,N_18368,N_13012);
nor U29767 (N_29767,N_10590,N_19400);
xnor U29768 (N_29768,N_11197,N_19392);
or U29769 (N_29769,N_18304,N_19864);
and U29770 (N_29770,N_10480,N_18937);
or U29771 (N_29771,N_15150,N_11206);
xnor U29772 (N_29772,N_13815,N_19374);
or U29773 (N_29773,N_18253,N_14578);
or U29774 (N_29774,N_19513,N_12253);
xor U29775 (N_29775,N_16826,N_17756);
and U29776 (N_29776,N_17466,N_18125);
and U29777 (N_29777,N_16175,N_13922);
xor U29778 (N_29778,N_18014,N_16963);
and U29779 (N_29779,N_18493,N_11199);
nor U29780 (N_29780,N_14490,N_12296);
nand U29781 (N_29781,N_14681,N_15072);
or U29782 (N_29782,N_11164,N_17474);
nor U29783 (N_29783,N_19597,N_16360);
xor U29784 (N_29784,N_12382,N_13680);
and U29785 (N_29785,N_16170,N_14856);
or U29786 (N_29786,N_16819,N_16723);
and U29787 (N_29787,N_16027,N_15244);
or U29788 (N_29788,N_10205,N_14554);
nand U29789 (N_29789,N_14074,N_13665);
xor U29790 (N_29790,N_14784,N_14316);
nor U29791 (N_29791,N_19913,N_14228);
or U29792 (N_29792,N_16657,N_10647);
nand U29793 (N_29793,N_18849,N_10458);
xnor U29794 (N_29794,N_18005,N_14520);
xor U29795 (N_29795,N_17591,N_11654);
and U29796 (N_29796,N_10233,N_12111);
nand U29797 (N_29797,N_17515,N_19765);
xnor U29798 (N_29798,N_18867,N_14823);
xor U29799 (N_29799,N_18326,N_14669);
or U29800 (N_29800,N_10180,N_12783);
nor U29801 (N_29801,N_14276,N_13331);
xnor U29802 (N_29802,N_11767,N_13564);
and U29803 (N_29803,N_13172,N_16702);
nand U29804 (N_29804,N_15459,N_10678);
or U29805 (N_29805,N_14106,N_17225);
xor U29806 (N_29806,N_15430,N_17857);
xor U29807 (N_29807,N_12569,N_19050);
nand U29808 (N_29808,N_18240,N_16684);
and U29809 (N_29809,N_15180,N_10247);
xnor U29810 (N_29810,N_10872,N_13076);
and U29811 (N_29811,N_14378,N_19879);
nor U29812 (N_29812,N_14600,N_15476);
nor U29813 (N_29813,N_19872,N_17215);
or U29814 (N_29814,N_18742,N_11341);
xnor U29815 (N_29815,N_19615,N_16178);
or U29816 (N_29816,N_19690,N_18167);
or U29817 (N_29817,N_15650,N_18783);
nand U29818 (N_29818,N_14806,N_10377);
xnor U29819 (N_29819,N_12579,N_16434);
xnor U29820 (N_29820,N_14515,N_16766);
nand U29821 (N_29821,N_10071,N_14655);
or U29822 (N_29822,N_10174,N_13149);
xnor U29823 (N_29823,N_16774,N_10934);
nand U29824 (N_29824,N_17384,N_14862);
nand U29825 (N_29825,N_12431,N_13038);
or U29826 (N_29826,N_16709,N_11959);
nand U29827 (N_29827,N_17062,N_15901);
nand U29828 (N_29828,N_19295,N_19339);
or U29829 (N_29829,N_15207,N_10850);
or U29830 (N_29830,N_16413,N_19199);
and U29831 (N_29831,N_19666,N_18470);
nor U29832 (N_29832,N_11159,N_10568);
and U29833 (N_29833,N_12998,N_15761);
xor U29834 (N_29834,N_11261,N_15970);
nand U29835 (N_29835,N_15633,N_13107);
xor U29836 (N_29836,N_11558,N_15750);
nand U29837 (N_29837,N_16032,N_13476);
and U29838 (N_29838,N_16967,N_16487);
xnor U29839 (N_29839,N_16445,N_14461);
and U29840 (N_29840,N_17532,N_15997);
nor U29841 (N_29841,N_12339,N_10612);
or U29842 (N_29842,N_17481,N_13793);
nor U29843 (N_29843,N_11186,N_14417);
and U29844 (N_29844,N_12051,N_15353);
nand U29845 (N_29845,N_15915,N_10680);
xor U29846 (N_29846,N_17842,N_12590);
nand U29847 (N_29847,N_19467,N_15503);
or U29848 (N_29848,N_19721,N_12977);
xor U29849 (N_29849,N_18716,N_15344);
nor U29850 (N_29850,N_15277,N_17952);
or U29851 (N_29851,N_19677,N_16470);
nand U29852 (N_29852,N_12162,N_17386);
xor U29853 (N_29853,N_16176,N_17327);
nand U29854 (N_29854,N_10935,N_10523);
or U29855 (N_29855,N_18669,N_18004);
nand U29856 (N_29856,N_18797,N_13306);
xor U29857 (N_29857,N_17539,N_17458);
and U29858 (N_29858,N_12168,N_16098);
or U29859 (N_29859,N_12233,N_13416);
xor U29860 (N_29860,N_17514,N_13540);
or U29861 (N_29861,N_18948,N_14366);
or U29862 (N_29862,N_17458,N_18687);
nor U29863 (N_29863,N_13331,N_15666);
xnor U29864 (N_29864,N_13528,N_13123);
or U29865 (N_29865,N_19396,N_15528);
xnor U29866 (N_29866,N_12280,N_16120);
or U29867 (N_29867,N_14836,N_19453);
and U29868 (N_29868,N_15823,N_10805);
xor U29869 (N_29869,N_12999,N_10154);
or U29870 (N_29870,N_17358,N_15432);
or U29871 (N_29871,N_15059,N_16960);
xnor U29872 (N_29872,N_13031,N_13788);
xor U29873 (N_29873,N_18882,N_10128);
xor U29874 (N_29874,N_16559,N_14399);
xnor U29875 (N_29875,N_10784,N_14692);
xnor U29876 (N_29876,N_15965,N_15641);
or U29877 (N_29877,N_13237,N_16739);
xor U29878 (N_29878,N_11964,N_12989);
and U29879 (N_29879,N_19627,N_19176);
nand U29880 (N_29880,N_17602,N_19186);
xor U29881 (N_29881,N_17563,N_17485);
xor U29882 (N_29882,N_16036,N_18695);
or U29883 (N_29883,N_13171,N_12367);
or U29884 (N_29884,N_18759,N_18169);
and U29885 (N_29885,N_13614,N_14315);
nor U29886 (N_29886,N_16362,N_11605);
nor U29887 (N_29887,N_18374,N_13318);
and U29888 (N_29888,N_13835,N_13815);
and U29889 (N_29889,N_18212,N_11641);
xor U29890 (N_29890,N_13293,N_18539);
or U29891 (N_29891,N_14191,N_12531);
xnor U29892 (N_29892,N_15572,N_10527);
or U29893 (N_29893,N_13593,N_12403);
or U29894 (N_29894,N_19993,N_10892);
or U29895 (N_29895,N_15302,N_17702);
or U29896 (N_29896,N_18827,N_12412);
nor U29897 (N_29897,N_11240,N_18007);
and U29898 (N_29898,N_11406,N_19425);
and U29899 (N_29899,N_11151,N_15567);
or U29900 (N_29900,N_15447,N_15576);
and U29901 (N_29901,N_10736,N_19685);
and U29902 (N_29902,N_17141,N_14079);
nand U29903 (N_29903,N_11182,N_11604);
or U29904 (N_29904,N_19423,N_13494);
nand U29905 (N_29905,N_12947,N_12895);
xor U29906 (N_29906,N_11180,N_14393);
xor U29907 (N_29907,N_11504,N_12670);
nand U29908 (N_29908,N_10511,N_17589);
or U29909 (N_29909,N_17315,N_16625);
nand U29910 (N_29910,N_11125,N_17540);
or U29911 (N_29911,N_13686,N_15418);
or U29912 (N_29912,N_14922,N_19726);
nand U29913 (N_29913,N_13323,N_10965);
or U29914 (N_29914,N_18123,N_17165);
or U29915 (N_29915,N_19327,N_12621);
and U29916 (N_29916,N_14626,N_17910);
nand U29917 (N_29917,N_15639,N_11066);
and U29918 (N_29918,N_11285,N_16471);
and U29919 (N_29919,N_17652,N_10567);
or U29920 (N_29920,N_11811,N_17383);
nand U29921 (N_29921,N_19843,N_11346);
and U29922 (N_29922,N_12579,N_15287);
nand U29923 (N_29923,N_16564,N_15346);
and U29924 (N_29924,N_14973,N_17322);
nor U29925 (N_29925,N_15705,N_19545);
nor U29926 (N_29926,N_19692,N_12614);
or U29927 (N_29927,N_17507,N_15502);
or U29928 (N_29928,N_18830,N_13141);
and U29929 (N_29929,N_11002,N_11888);
and U29930 (N_29930,N_15965,N_19417);
xnor U29931 (N_29931,N_12010,N_11972);
nand U29932 (N_29932,N_16000,N_17307);
nand U29933 (N_29933,N_18676,N_12255);
xnor U29934 (N_29934,N_12700,N_17271);
xor U29935 (N_29935,N_10337,N_12932);
xnor U29936 (N_29936,N_18840,N_15152);
nor U29937 (N_29937,N_15132,N_19270);
nand U29938 (N_29938,N_13637,N_12782);
and U29939 (N_29939,N_14688,N_13075);
and U29940 (N_29940,N_12707,N_11915);
nor U29941 (N_29941,N_19495,N_12927);
and U29942 (N_29942,N_12442,N_18422);
nor U29943 (N_29943,N_14064,N_17940);
xor U29944 (N_29944,N_10319,N_14227);
xor U29945 (N_29945,N_17577,N_11361);
and U29946 (N_29946,N_11108,N_17289);
nand U29947 (N_29947,N_15934,N_14442);
nand U29948 (N_29948,N_13657,N_18926);
xor U29949 (N_29949,N_18499,N_13224);
nor U29950 (N_29950,N_10552,N_10985);
nor U29951 (N_29951,N_15437,N_16381);
xor U29952 (N_29952,N_14288,N_14605);
nand U29953 (N_29953,N_18330,N_13593);
or U29954 (N_29954,N_17969,N_16001);
nand U29955 (N_29955,N_13423,N_17396);
xnor U29956 (N_29956,N_14612,N_10202);
nor U29957 (N_29957,N_11388,N_19487);
or U29958 (N_29958,N_10899,N_13220);
and U29959 (N_29959,N_17655,N_16064);
or U29960 (N_29960,N_13385,N_14924);
or U29961 (N_29961,N_10611,N_17569);
and U29962 (N_29962,N_16762,N_18325);
nand U29963 (N_29963,N_19446,N_16371);
or U29964 (N_29964,N_17736,N_16665);
xnor U29965 (N_29965,N_13982,N_13907);
and U29966 (N_29966,N_15180,N_13205);
xor U29967 (N_29967,N_11293,N_10004);
nand U29968 (N_29968,N_12074,N_17970);
or U29969 (N_29969,N_18225,N_10856);
xor U29970 (N_29970,N_15297,N_16455);
xor U29971 (N_29971,N_17898,N_15242);
nand U29972 (N_29972,N_18019,N_18120);
nor U29973 (N_29973,N_19893,N_11163);
and U29974 (N_29974,N_13941,N_10472);
nand U29975 (N_29975,N_13071,N_19199);
and U29976 (N_29976,N_18764,N_16355);
nor U29977 (N_29977,N_10814,N_19930);
or U29978 (N_29978,N_19916,N_15260);
and U29979 (N_29979,N_13687,N_10555);
xor U29980 (N_29980,N_11361,N_13751);
nand U29981 (N_29981,N_12789,N_19017);
and U29982 (N_29982,N_10579,N_10627);
xnor U29983 (N_29983,N_10088,N_11238);
xor U29984 (N_29984,N_19847,N_13273);
xnor U29985 (N_29985,N_17007,N_10699);
nor U29986 (N_29986,N_18720,N_14392);
xnor U29987 (N_29987,N_16100,N_17352);
xor U29988 (N_29988,N_13388,N_17765);
or U29989 (N_29989,N_14244,N_16129);
and U29990 (N_29990,N_10948,N_16559);
nand U29991 (N_29991,N_18660,N_18087);
xnor U29992 (N_29992,N_11164,N_16256);
nand U29993 (N_29993,N_17467,N_11554);
or U29994 (N_29994,N_12108,N_14200);
nor U29995 (N_29995,N_12300,N_10568);
xnor U29996 (N_29996,N_18482,N_16904);
nand U29997 (N_29997,N_14771,N_10878);
xnor U29998 (N_29998,N_15808,N_17174);
and U29999 (N_29999,N_15744,N_14783);
xnor U30000 (N_30000,N_27989,N_26821);
xor U30001 (N_30001,N_24321,N_27683);
or U30002 (N_30002,N_22959,N_23494);
xor U30003 (N_30003,N_24369,N_22485);
or U30004 (N_30004,N_20502,N_20588);
or U30005 (N_30005,N_21064,N_20049);
xnor U30006 (N_30006,N_28586,N_27156);
or U30007 (N_30007,N_25813,N_24017);
or U30008 (N_30008,N_29538,N_24592);
or U30009 (N_30009,N_28676,N_24507);
xnor U30010 (N_30010,N_25437,N_28423);
xor U30011 (N_30011,N_23628,N_27170);
and U30012 (N_30012,N_27804,N_22994);
nand U30013 (N_30013,N_24874,N_21047);
nor U30014 (N_30014,N_26349,N_29649);
or U30015 (N_30015,N_23205,N_24548);
and U30016 (N_30016,N_27489,N_28693);
or U30017 (N_30017,N_29263,N_20066);
or U30018 (N_30018,N_24806,N_22021);
and U30019 (N_30019,N_26933,N_28845);
and U30020 (N_30020,N_27135,N_23105);
or U30021 (N_30021,N_25763,N_29793);
and U30022 (N_30022,N_21678,N_26092);
nand U30023 (N_30023,N_24420,N_27221);
nand U30024 (N_30024,N_20669,N_22902);
xnor U30025 (N_30025,N_22808,N_20207);
xor U30026 (N_30026,N_28155,N_25331);
nand U30027 (N_30027,N_24946,N_26827);
xor U30028 (N_30028,N_27967,N_23271);
or U30029 (N_30029,N_23386,N_25844);
nor U30030 (N_30030,N_23533,N_29244);
xnor U30031 (N_30031,N_22505,N_27469);
or U30032 (N_30032,N_29723,N_23107);
or U30033 (N_30033,N_24144,N_27866);
and U30034 (N_30034,N_20677,N_28730);
and U30035 (N_30035,N_20014,N_24208);
and U30036 (N_30036,N_22811,N_20539);
xor U30037 (N_30037,N_27441,N_25637);
or U30038 (N_30038,N_27034,N_29280);
and U30039 (N_30039,N_27837,N_26341);
or U30040 (N_30040,N_28794,N_29343);
xor U30041 (N_30041,N_20815,N_24585);
nor U30042 (N_30042,N_25333,N_24694);
nand U30043 (N_30043,N_20348,N_27716);
nor U30044 (N_30044,N_25747,N_21837);
nand U30045 (N_30045,N_23146,N_22300);
xnor U30046 (N_30046,N_21217,N_29906);
and U30047 (N_30047,N_26331,N_25297);
xnor U30048 (N_30048,N_23503,N_27497);
nand U30049 (N_30049,N_26424,N_24239);
xnor U30050 (N_30050,N_20298,N_25795);
or U30051 (N_30051,N_24226,N_28762);
nor U30052 (N_30052,N_28765,N_22032);
or U30053 (N_30053,N_21629,N_25674);
and U30054 (N_30054,N_23474,N_28516);
and U30055 (N_30055,N_21677,N_28497);
nor U30056 (N_30056,N_26145,N_22879);
nand U30057 (N_30057,N_28561,N_28174);
or U30058 (N_30058,N_24060,N_20172);
and U30059 (N_30059,N_28735,N_29541);
nor U30060 (N_30060,N_23539,N_24608);
or U30061 (N_30061,N_25244,N_25607);
and U30062 (N_30062,N_22154,N_20703);
nor U30063 (N_30063,N_29057,N_27163);
xor U30064 (N_30064,N_29051,N_29743);
nand U30065 (N_30065,N_27485,N_22200);
xor U30066 (N_30066,N_22752,N_20915);
nor U30067 (N_30067,N_21891,N_25682);
or U30068 (N_30068,N_24209,N_28906);
or U30069 (N_30069,N_29121,N_21504);
nor U30070 (N_30070,N_25553,N_21222);
nor U30071 (N_30071,N_29481,N_20320);
xnor U30072 (N_30072,N_26287,N_25838);
xnor U30073 (N_30073,N_29861,N_24791);
or U30074 (N_30074,N_25578,N_21490);
or U30075 (N_30075,N_21089,N_25147);
nor U30076 (N_30076,N_23215,N_22182);
xnor U30077 (N_30077,N_23608,N_27955);
nand U30078 (N_30078,N_27768,N_20384);
nand U30079 (N_30079,N_26540,N_25106);
nor U30080 (N_30080,N_21668,N_20259);
and U30081 (N_30081,N_29809,N_23344);
or U30082 (N_30082,N_24130,N_22593);
nand U30083 (N_30083,N_21675,N_22401);
or U30084 (N_30084,N_22135,N_26284);
xor U30085 (N_30085,N_25231,N_23831);
xor U30086 (N_30086,N_20798,N_25234);
nand U30087 (N_30087,N_21092,N_24377);
nor U30088 (N_30088,N_26398,N_22615);
nand U30089 (N_30089,N_22102,N_23597);
nand U30090 (N_30090,N_25898,N_25424);
nor U30091 (N_30091,N_25748,N_29254);
xor U30092 (N_30092,N_26584,N_29171);
xor U30093 (N_30093,N_26844,N_28124);
nand U30094 (N_30094,N_21660,N_24700);
or U30095 (N_30095,N_22209,N_27902);
or U30096 (N_30096,N_22267,N_25011);
nor U30097 (N_30097,N_29209,N_25506);
nor U30098 (N_30098,N_25537,N_24812);
nor U30099 (N_30099,N_20012,N_22239);
xnor U30100 (N_30100,N_20893,N_24170);
nand U30101 (N_30101,N_24508,N_26296);
nor U30102 (N_30102,N_29318,N_25451);
nand U30103 (N_30103,N_24442,N_25890);
or U30104 (N_30104,N_24906,N_21845);
or U30105 (N_30105,N_24088,N_29880);
nor U30106 (N_30106,N_23411,N_29806);
nand U30107 (N_30107,N_29805,N_20488);
and U30108 (N_30108,N_25115,N_28198);
nand U30109 (N_30109,N_27872,N_21904);
nand U30110 (N_30110,N_29627,N_24461);
xor U30111 (N_30111,N_22490,N_24318);
or U30112 (N_30112,N_27946,N_27400);
and U30113 (N_30113,N_22338,N_25953);
xnor U30114 (N_30114,N_24681,N_23629);
nor U30115 (N_30115,N_22988,N_27301);
xnor U30116 (N_30116,N_21104,N_28040);
nor U30117 (N_30117,N_22329,N_29549);
nand U30118 (N_30118,N_26954,N_24002);
xnor U30119 (N_30119,N_27059,N_21354);
xnor U30120 (N_30120,N_20751,N_23330);
or U30121 (N_30121,N_23854,N_25420);
or U30122 (N_30122,N_29108,N_26358);
and U30123 (N_30123,N_29501,N_27936);
nor U30124 (N_30124,N_26602,N_24549);
nor U30125 (N_30125,N_26258,N_21263);
or U30126 (N_30126,N_20901,N_20850);
nor U30127 (N_30127,N_21010,N_25756);
xor U30128 (N_30128,N_25308,N_25501);
nor U30129 (N_30129,N_21373,N_21695);
nor U30130 (N_30130,N_23864,N_27855);
or U30131 (N_30131,N_22223,N_28227);
or U30132 (N_30132,N_29186,N_25037);
nor U30133 (N_30133,N_25332,N_22174);
nor U30134 (N_30134,N_23856,N_22423);
and U30135 (N_30135,N_24721,N_20907);
nor U30136 (N_30136,N_21808,N_26043);
nand U30137 (N_30137,N_24824,N_22483);
nand U30138 (N_30138,N_25622,N_20081);
or U30139 (N_30139,N_23946,N_29686);
and U30140 (N_30140,N_21709,N_28454);
xnor U30141 (N_30141,N_28038,N_24529);
and U30142 (N_30142,N_28449,N_20745);
and U30143 (N_30143,N_22399,N_27010);
or U30144 (N_30144,N_23471,N_21550);
and U30145 (N_30145,N_23700,N_23941);
and U30146 (N_30146,N_26867,N_20610);
and U30147 (N_30147,N_26712,N_23573);
nor U30148 (N_30148,N_28445,N_20167);
nor U30149 (N_30149,N_26193,N_29768);
nand U30150 (N_30150,N_23113,N_28201);
and U30151 (N_30151,N_25862,N_24573);
nand U30152 (N_30152,N_24543,N_21260);
and U30153 (N_30153,N_27054,N_29359);
xnor U30154 (N_30154,N_20950,N_22346);
or U30155 (N_30155,N_25847,N_25870);
nor U30156 (N_30156,N_24654,N_28129);
nor U30157 (N_30157,N_22552,N_29041);
and U30158 (N_30158,N_23722,N_24828);
and U30159 (N_30159,N_28701,N_22681);
nor U30160 (N_30160,N_29037,N_22510);
xnor U30161 (N_30161,N_21184,N_23377);
nand U30162 (N_30162,N_26757,N_21800);
or U30163 (N_30163,N_26134,N_29350);
nor U30164 (N_30164,N_28492,N_21231);
nand U30165 (N_30165,N_26244,N_24020);
and U30166 (N_30166,N_27682,N_28630);
nand U30167 (N_30167,N_29980,N_26314);
and U30168 (N_30168,N_20109,N_28973);
or U30169 (N_30169,N_22464,N_29533);
and U30170 (N_30170,N_26897,N_20995);
nor U30171 (N_30171,N_29147,N_24082);
nor U30172 (N_30172,N_28439,N_24521);
nand U30173 (N_30173,N_20699,N_25216);
nor U30174 (N_30174,N_21117,N_28432);
xnor U30175 (N_30175,N_22380,N_22074);
nand U30176 (N_30176,N_29513,N_26952);
xnor U30177 (N_30177,N_27066,N_23884);
xnor U30178 (N_30178,N_26870,N_22240);
xnor U30179 (N_30179,N_27950,N_27629);
xnor U30180 (N_30180,N_26750,N_26487);
nor U30181 (N_30181,N_28123,N_25427);
nand U30182 (N_30182,N_29000,N_26783);
or U30183 (N_30183,N_29170,N_27265);
or U30184 (N_30184,N_28313,N_21048);
and U30185 (N_30185,N_21429,N_25034);
nor U30186 (N_30186,N_22217,N_27307);
nand U30187 (N_30187,N_22000,N_28000);
nand U30188 (N_30188,N_20152,N_20465);
nor U30189 (N_30189,N_20038,N_24197);
or U30190 (N_30190,N_21824,N_22437);
xor U30191 (N_30191,N_20986,N_26495);
and U30192 (N_30192,N_22829,N_27891);
or U30193 (N_30193,N_21006,N_28650);
nand U30194 (N_30194,N_26200,N_24313);
and U30195 (N_30195,N_24024,N_28804);
xor U30196 (N_30196,N_22215,N_28099);
xnor U30197 (N_30197,N_27092,N_20494);
xnor U30198 (N_30198,N_23585,N_28779);
and U30199 (N_30199,N_24825,N_28412);
or U30200 (N_30200,N_27518,N_28820);
xor U30201 (N_30201,N_23319,N_26709);
nand U30202 (N_30202,N_23255,N_21026);
xor U30203 (N_30203,N_22616,N_24268);
or U30204 (N_30204,N_21991,N_29183);
nand U30205 (N_30205,N_22018,N_27353);
and U30206 (N_30206,N_24409,N_27127);
and U30207 (N_30207,N_25993,N_22192);
or U30208 (N_30208,N_26049,N_27199);
xnor U30209 (N_30209,N_23899,N_26771);
xnor U30210 (N_30210,N_23536,N_25593);
and U30211 (N_30211,N_21063,N_24818);
or U30212 (N_30212,N_29948,N_23500);
or U30213 (N_30213,N_25527,N_21335);
or U30214 (N_30214,N_21135,N_22066);
nor U30215 (N_30215,N_28008,N_20695);
xor U30216 (N_30216,N_26724,N_20782);
nand U30217 (N_30217,N_24089,N_28297);
or U30218 (N_30218,N_28411,N_29437);
nand U30219 (N_30219,N_24183,N_28728);
or U30220 (N_30220,N_21622,N_22295);
nand U30221 (N_30221,N_25525,N_27897);
nor U30222 (N_30222,N_27520,N_21963);
or U30223 (N_30223,N_20379,N_26065);
nand U30224 (N_30224,N_20036,N_29469);
or U30225 (N_30225,N_25171,N_22160);
nor U30226 (N_30226,N_25943,N_28293);
and U30227 (N_30227,N_23203,N_20486);
and U30228 (N_30228,N_29797,N_21012);
or U30229 (N_30229,N_24108,N_27446);
or U30230 (N_30230,N_20341,N_26434);
and U30231 (N_30231,N_26887,N_25690);
xnor U30232 (N_30232,N_26469,N_21269);
or U30233 (N_30233,N_24191,N_26937);
or U30234 (N_30234,N_29427,N_25928);
nor U30235 (N_30235,N_29008,N_27638);
or U30236 (N_30236,N_24685,N_23996);
nor U30237 (N_30237,N_26411,N_20561);
xor U30238 (N_30238,N_27830,N_29908);
or U30239 (N_30239,N_25602,N_20373);
xnor U30240 (N_30240,N_24388,N_25640);
or U30241 (N_30241,N_28504,N_20437);
xnor U30242 (N_30242,N_28408,N_23914);
and U30243 (N_30243,N_29419,N_22585);
nand U30244 (N_30244,N_25175,N_25086);
nand U30245 (N_30245,N_26249,N_28241);
nand U30246 (N_30246,N_26537,N_22537);
nor U30247 (N_30247,N_28685,N_29589);
and U30248 (N_30248,N_25361,N_28004);
xor U30249 (N_30249,N_24302,N_24842);
and U30250 (N_30250,N_28361,N_26586);
or U30251 (N_30251,N_29591,N_26667);
or U30252 (N_30252,N_22716,N_22546);
or U30253 (N_30253,N_22313,N_27146);
nand U30254 (N_30254,N_26585,N_29467);
xnor U30255 (N_30255,N_27733,N_28874);
nor U30256 (N_30256,N_27125,N_27311);
nor U30257 (N_30257,N_21308,N_24075);
and U30258 (N_30258,N_20820,N_22415);
nor U30259 (N_30259,N_28932,N_28643);
xnor U30260 (N_30260,N_25514,N_28646);
and U30261 (N_30261,N_29613,N_21834);
or U30262 (N_30262,N_22062,N_23744);
xor U30263 (N_30263,N_21817,N_25168);
xnor U30264 (N_30264,N_23976,N_28394);
nor U30265 (N_30265,N_25678,N_20071);
xor U30266 (N_30266,N_21646,N_21149);
nand U30267 (N_30267,N_26310,N_27289);
xnor U30268 (N_30268,N_20719,N_23357);
and U30269 (N_30269,N_24742,N_23785);
nor U30270 (N_30270,N_23784,N_20645);
nor U30271 (N_30271,N_20473,N_26105);
nand U30272 (N_30272,N_27041,N_24703);
or U30273 (N_30273,N_22828,N_24662);
nand U30274 (N_30274,N_20190,N_25035);
xnor U30275 (N_30275,N_21948,N_22059);
xor U30276 (N_30276,N_26531,N_29043);
nand U30277 (N_30277,N_28850,N_25941);
nand U30278 (N_30278,N_27115,N_24695);
or U30279 (N_30279,N_20346,N_22765);
xnor U30280 (N_30280,N_29250,N_21836);
nand U30281 (N_30281,N_22414,N_29891);
nor U30282 (N_30282,N_27206,N_23001);
and U30283 (N_30283,N_22722,N_25974);
and U30284 (N_30284,N_27616,N_21398);
and U30285 (N_30285,N_20142,N_28546);
xor U30286 (N_30286,N_24111,N_21000);
nand U30287 (N_30287,N_20999,N_24093);
nand U30288 (N_30288,N_29347,N_20008);
and U30289 (N_30289,N_28175,N_22461);
xnor U30290 (N_30290,N_21513,N_21103);
and U30291 (N_30291,N_26231,N_24135);
nand U30292 (N_30292,N_28409,N_27542);
nor U30293 (N_30293,N_25612,N_23896);
nor U30294 (N_30294,N_27428,N_28360);
nor U30295 (N_30295,N_27618,N_24346);
or U30296 (N_30296,N_23466,N_23659);
nand U30297 (N_30297,N_26617,N_23118);
and U30298 (N_30298,N_25311,N_26290);
and U30299 (N_30299,N_27286,N_21296);
nand U30300 (N_30300,N_21697,N_23367);
nor U30301 (N_30301,N_20085,N_27828);
xnor U30302 (N_30302,N_20403,N_21057);
and U30303 (N_30303,N_27023,N_20533);
and U30304 (N_30304,N_28415,N_28405);
nor U30305 (N_30305,N_28997,N_21031);
or U30306 (N_30306,N_24952,N_20933);
nor U30307 (N_30307,N_29019,N_28603);
or U30308 (N_30308,N_27306,N_23593);
and U30309 (N_30309,N_26230,N_26519);
xnor U30310 (N_30310,N_25883,N_21291);
and U30311 (N_30311,N_28739,N_22030);
and U30312 (N_30312,N_22194,N_24764);
xor U30313 (N_30313,N_22596,N_26390);
and U30314 (N_30314,N_28625,N_24145);
nand U30315 (N_30315,N_28840,N_27103);
nor U30316 (N_30316,N_29257,N_20587);
nand U30317 (N_30317,N_27153,N_24672);
nor U30318 (N_30318,N_24553,N_22232);
or U30319 (N_30319,N_29114,N_26172);
nor U30320 (N_30320,N_26592,N_27669);
nand U30321 (N_30321,N_23038,N_24217);
nand U30322 (N_30322,N_28799,N_22573);
xor U30323 (N_30323,N_28868,N_27749);
xor U30324 (N_30324,N_22337,N_20443);
or U30325 (N_30325,N_26762,N_29623);
and U30326 (N_30326,N_27220,N_20225);
and U30327 (N_30327,N_23522,N_24206);
and U30328 (N_30328,N_27598,N_28253);
and U30329 (N_30329,N_29372,N_26914);
xor U30330 (N_30330,N_23065,N_21146);
and U30331 (N_30331,N_29682,N_25985);
nor U30332 (N_30332,N_21993,N_25080);
and U30333 (N_30333,N_23160,N_29465);
and U30334 (N_30334,N_24370,N_26634);
or U30335 (N_30335,N_23887,N_20663);
and U30336 (N_30336,N_26706,N_20089);
or U30337 (N_30337,N_29242,N_21692);
nand U30338 (N_30338,N_24886,N_28212);
nor U30339 (N_30339,N_26958,N_27611);
nor U30340 (N_30340,N_25850,N_24050);
xnor U30341 (N_30341,N_24912,N_28232);
and U30342 (N_30342,N_23297,N_20394);
nor U30343 (N_30343,N_25729,N_20770);
nand U30344 (N_30344,N_26361,N_23197);
or U30345 (N_30345,N_25348,N_20434);
or U30346 (N_30346,N_24281,N_21610);
nand U30347 (N_30347,N_25393,N_22119);
or U30348 (N_30348,N_23457,N_21727);
or U30349 (N_30349,N_23705,N_29292);
nand U30350 (N_30350,N_24419,N_24305);
nand U30351 (N_30351,N_26833,N_26294);
and U30352 (N_30352,N_22158,N_23764);
xnor U30353 (N_30353,N_20431,N_26129);
or U30354 (N_30354,N_23400,N_28292);
xnor U30355 (N_30355,N_22562,N_23314);
nand U30356 (N_30356,N_28535,N_21218);
or U30357 (N_30357,N_22650,N_27925);
nand U30358 (N_30358,N_24123,N_25962);
or U30359 (N_30359,N_22384,N_22785);
nand U30360 (N_30360,N_26219,N_28855);
nor U30361 (N_30361,N_27114,N_25920);
and U30362 (N_30362,N_29996,N_25705);
and U30363 (N_30363,N_23625,N_22165);
and U30364 (N_30364,N_26595,N_20381);
nand U30365 (N_30365,N_27329,N_21211);
nand U30366 (N_30366,N_22255,N_26546);
nand U30367 (N_30367,N_21542,N_28944);
nor U30368 (N_30368,N_29593,N_20467);
or U30369 (N_30369,N_24792,N_27434);
xor U30370 (N_30370,N_24137,N_24431);
nor U30371 (N_30371,N_23394,N_23791);
nand U30372 (N_30372,N_29751,N_21798);
nor U30373 (N_30373,N_21999,N_28006);
nor U30374 (N_30374,N_23995,N_28353);
or U30375 (N_30375,N_28748,N_22706);
and U30376 (N_30376,N_21912,N_28980);
xor U30377 (N_30377,N_26682,N_23777);
or U30378 (N_30378,N_20455,N_28427);
nor U30379 (N_30379,N_21890,N_23682);
and U30380 (N_30380,N_23492,N_27349);
or U30381 (N_30381,N_29144,N_27850);
nor U30382 (N_30382,N_29022,N_20478);
xnor U30383 (N_30383,N_23620,N_26809);
nand U30384 (N_30384,N_26940,N_26037);
xor U30385 (N_30385,N_21616,N_24414);
or U30386 (N_30386,N_23423,N_23773);
or U30387 (N_30387,N_25353,N_26416);
nor U30388 (N_30388,N_25210,N_22095);
and U30389 (N_30389,N_28462,N_24869);
and U30390 (N_30390,N_24478,N_26376);
nor U30391 (N_30391,N_24113,N_28900);
nand U30392 (N_30392,N_29960,N_26094);
nor U30393 (N_30393,N_28969,N_29458);
nor U30394 (N_30394,N_27931,N_25782);
or U30395 (N_30395,N_23210,N_25724);
nor U30396 (N_30396,N_26456,N_29138);
and U30397 (N_30397,N_20504,N_27342);
nand U30398 (N_30398,N_27351,N_20653);
xor U30399 (N_30399,N_27612,N_24330);
and U30400 (N_30400,N_21451,N_26525);
nand U30401 (N_30401,N_28143,N_20170);
nand U30402 (N_30402,N_21264,N_29354);
nor U30403 (N_30403,N_22574,N_26322);
and U30404 (N_30404,N_25854,N_21742);
xnor U30405 (N_30405,N_23053,N_25293);
nand U30406 (N_30406,N_22053,N_22726);
nand U30407 (N_30407,N_25542,N_28431);
nand U30408 (N_30408,N_21213,N_27184);
and U30409 (N_30409,N_20644,N_23228);
nand U30410 (N_30410,N_24413,N_27444);
nor U30411 (N_30411,N_21722,N_20256);
or U30412 (N_30412,N_23653,N_27303);
or U30413 (N_30413,N_22936,N_25045);
xor U30414 (N_30414,N_27008,N_28047);
nand U30415 (N_30415,N_28512,N_28696);
nand U30416 (N_30416,N_25468,N_25471);
nand U30417 (N_30417,N_20721,N_29860);
nand U30418 (N_30418,N_28108,N_26074);
xor U30419 (N_30419,N_20715,N_23241);
nand U30420 (N_30420,N_22570,N_24077);
nor U30421 (N_30421,N_29023,N_23017);
xnor U30422 (N_30422,N_26370,N_26421);
or U30423 (N_30423,N_23942,N_22618);
and U30424 (N_30424,N_25726,N_20343);
nand U30425 (N_30425,N_23863,N_21522);
nand U30426 (N_30426,N_25919,N_22273);
or U30427 (N_30427,N_20073,N_23944);
and U30428 (N_30428,N_29294,N_29048);
nand U30429 (N_30429,N_27980,N_22807);
nor U30430 (N_30430,N_21302,N_29528);
and U30431 (N_30431,N_25407,N_23592);
xnor U30432 (N_30432,N_25609,N_25618);
or U30433 (N_30433,N_20557,N_23819);
xnor U30434 (N_30434,N_23014,N_20590);
nand U30435 (N_30435,N_21068,N_23832);
nand U30436 (N_30436,N_22360,N_24990);
nand U30437 (N_30437,N_28946,N_20265);
or U30438 (N_30438,N_24174,N_25275);
or U30439 (N_30439,N_29971,N_20651);
xnor U30440 (N_30440,N_23235,N_26190);
nand U30441 (N_30441,N_27603,N_20902);
nor U30442 (N_30442,N_29647,N_29231);
nand U30443 (N_30443,N_23754,N_28806);
and U30444 (N_30444,N_20233,N_20058);
or U30445 (N_30445,N_21950,N_24348);
nand U30446 (N_30446,N_24037,N_26579);
nand U30447 (N_30447,N_20573,N_28429);
or U30448 (N_30448,N_21744,N_20971);
or U30449 (N_30449,N_20618,N_23081);
nand U30450 (N_30450,N_21957,N_26926);
nand U30451 (N_30451,N_20282,N_23485);
or U30452 (N_30452,N_25755,N_20023);
nor U30453 (N_30453,N_27355,N_24336);
and U30454 (N_30454,N_28579,N_20292);
nand U30455 (N_30455,N_22728,N_26992);
xor U30456 (N_30456,N_29859,N_21517);
or U30457 (N_30457,N_27278,N_21621);
nor U30458 (N_30458,N_27697,N_22605);
and U30459 (N_30459,N_23894,N_27492);
nand U30460 (N_30460,N_25722,N_29519);
nand U30461 (N_30461,N_27223,N_26217);
nand U30462 (N_30462,N_27763,N_27522);
xor U30463 (N_30463,N_28611,N_25446);
nor U30464 (N_30464,N_21278,N_24062);
nor U30465 (N_30465,N_27427,N_25672);
and U30466 (N_30466,N_23786,N_20459);
xor U30467 (N_30467,N_21555,N_25877);
nand U30468 (N_30468,N_28942,N_21942);
and U30469 (N_30469,N_20218,N_25576);
and U30470 (N_30470,N_25192,N_28569);
nand U30471 (N_30471,N_27971,N_20382);
xor U30472 (N_30472,N_25884,N_20702);
nand U30473 (N_30473,N_27599,N_22286);
or U30474 (N_30474,N_20744,N_20617);
nor U30475 (N_30475,N_21988,N_24168);
or U30476 (N_30476,N_20297,N_29977);
and U30477 (N_30477,N_29409,N_22339);
nor U30478 (N_30478,N_28817,N_25436);
xnor U30479 (N_30479,N_20694,N_26011);
nor U30480 (N_30480,N_20750,N_21714);
nor U30481 (N_30481,N_27413,N_29447);
nor U30482 (N_30482,N_22324,N_21433);
xor U30483 (N_30483,N_21615,N_29824);
xor U30484 (N_30484,N_26086,N_29073);
xnor U30485 (N_30485,N_24300,N_21319);
nor U30486 (N_30486,N_28468,N_22703);
xnor U30487 (N_30487,N_29645,N_27300);
nand U30488 (N_30488,N_27514,N_24372);
or U30489 (N_30489,N_21603,N_23756);
nor U30490 (N_30490,N_21310,N_23354);
nor U30491 (N_30491,N_28245,N_21625);
or U30492 (N_30492,N_23414,N_29319);
xor U30493 (N_30493,N_20116,N_23097);
xor U30494 (N_30494,N_24148,N_21474);
or U30495 (N_30495,N_21832,N_26265);
nand U30496 (N_30496,N_26476,N_28968);
or U30497 (N_30497,N_24884,N_26460);
xor U30498 (N_30498,N_24736,N_29365);
xnor U30499 (N_30499,N_20408,N_21033);
xor U30500 (N_30500,N_23519,N_27585);
xnor U30501 (N_30501,N_29554,N_21377);
nand U30502 (N_30502,N_20909,N_23555);
and U30503 (N_30503,N_28350,N_25474);
nand U30504 (N_30504,N_21635,N_26034);
nor U30505 (N_30505,N_23551,N_23232);
nand U30506 (N_30506,N_27819,N_22492);
nor U30507 (N_30507,N_23427,N_25054);
nor U30508 (N_30508,N_22904,N_21069);
or U30509 (N_30509,N_24678,N_25739);
or U30510 (N_30510,N_23164,N_26872);
nand U30511 (N_30511,N_25365,N_26765);
xor U30512 (N_30512,N_25939,N_23028);
and U30513 (N_30513,N_25958,N_25793);
nand U30514 (N_30514,N_28829,N_29119);
xnor U30515 (N_30515,N_27861,N_26443);
nor U30516 (N_30516,N_24561,N_22104);
and U30517 (N_30517,N_27188,N_29540);
nand U30518 (N_30518,N_23022,N_25935);
nand U30519 (N_30519,N_21261,N_21495);
xnor U30520 (N_30520,N_27397,N_22884);
nor U30521 (N_30521,N_22643,N_27570);
nand U30522 (N_30522,N_22504,N_22371);
and U30523 (N_30523,N_22531,N_28848);
and U30524 (N_30524,N_23306,N_20808);
xnor U30525 (N_30525,N_20941,N_25122);
nor U30526 (N_30526,N_24832,N_20659);
or U30527 (N_30527,N_24524,N_27614);
and U30528 (N_30528,N_21844,N_27121);
and U30529 (N_30529,N_23943,N_25623);
nor U30530 (N_30530,N_22971,N_28189);
or U30531 (N_30531,N_20526,N_20792);
nor U30532 (N_30532,N_20684,N_28918);
and U30533 (N_30533,N_29093,N_22746);
and U30534 (N_30534,N_28529,N_27200);
nor U30535 (N_30535,N_27896,N_26779);
xor U30536 (N_30536,N_28954,N_26311);
and U30537 (N_30537,N_21165,N_29607);
and U30538 (N_30538,N_22146,N_26710);
or U30539 (N_30539,N_26414,N_22507);
and U30540 (N_30540,N_27874,N_25668);
nor U30541 (N_30541,N_22780,N_29732);
nand U30542 (N_30542,N_22448,N_22721);
nor U30543 (N_30543,N_29007,N_21004);
xnor U30544 (N_30544,N_22456,N_24619);
nor U30545 (N_30545,N_21502,N_26980);
nor U30546 (N_30546,N_21364,N_20356);
nand U30547 (N_30547,N_22913,N_26665);
nor U30548 (N_30548,N_29411,N_21861);
and U30549 (N_30549,N_29067,N_26834);
nand U30550 (N_30550,N_29085,N_25486);
nor U30551 (N_30551,N_28583,N_20558);
nor U30552 (N_30552,N_24754,N_27484);
xor U30553 (N_30553,N_26632,N_29962);
xor U30554 (N_30554,N_28349,N_25590);
nor U30555 (N_30555,N_26649,N_28186);
nand U30556 (N_30556,N_22175,N_21931);
xor U30557 (N_30557,N_26913,N_28766);
or U30558 (N_30558,N_29935,N_20838);
xor U30559 (N_30559,N_21851,N_20364);
nor U30560 (N_30560,N_20930,N_24294);
or U30561 (N_30561,N_25000,N_23529);
and U30562 (N_30562,N_21865,N_22417);
nor U30563 (N_30563,N_22016,N_22438);
xnor U30564 (N_30564,N_25283,N_25669);
or U30565 (N_30565,N_26628,N_21856);
nand U30566 (N_30566,N_27601,N_20352);
or U30567 (N_30567,N_29397,N_23712);
nor U30568 (N_30568,N_20463,N_20175);
nand U30569 (N_30569,N_22606,N_20097);
or U30570 (N_30570,N_24621,N_23666);
or U30571 (N_30571,N_23327,N_27923);
nand U30572 (N_30572,N_22449,N_23737);
xnor U30573 (N_30573,N_26022,N_20221);
xnor U30574 (N_30574,N_23076,N_29867);
nand U30575 (N_30575,N_23813,N_22115);
nor U30576 (N_30576,N_26640,N_21743);
nand U30577 (N_30577,N_23116,N_21765);
nor U30578 (N_30578,N_20104,N_25246);
or U30579 (N_30579,N_20330,N_21516);
nor U30580 (N_30580,N_21353,N_23456);
and U30581 (N_30581,N_26036,N_23574);
xor U30582 (N_30582,N_27634,N_20180);
and U30583 (N_30583,N_26985,N_20082);
nor U30584 (N_30584,N_24526,N_29398);
or U30585 (N_30585,N_23994,N_24120);
nor U30586 (N_30586,N_29026,N_21203);
xor U30587 (N_30587,N_29753,N_24448);
and U30588 (N_30588,N_21854,N_20595);
nor U30589 (N_30589,N_21822,N_27986);
xnor U30590 (N_30590,N_29535,N_25188);
or U30591 (N_30591,N_23590,N_24185);
and U30592 (N_30592,N_23563,N_27963);
nor U30593 (N_30593,N_25496,N_24643);
and U30594 (N_30594,N_23112,N_28965);
or U30595 (N_30595,N_26806,N_24378);
and U30596 (N_30596,N_21640,N_27490);
nand U30597 (N_30597,N_21870,N_22263);
xnor U30598 (N_30598,N_21016,N_27820);
or U30599 (N_30599,N_20018,N_24233);
nand U30600 (N_30600,N_22151,N_22727);
or U30601 (N_30601,N_26758,N_23387);
or U30602 (N_30602,N_20518,N_24985);
xor U30603 (N_30603,N_27326,N_23757);
and U30604 (N_30604,N_28347,N_24980);
nor U30605 (N_30605,N_27096,N_25874);
nand U30606 (N_30606,N_25964,N_26500);
nor U30607 (N_30607,N_23860,N_27470);
nor U30608 (N_30608,N_21820,N_24994);
and U30609 (N_30609,N_21951,N_25875);
nand U30610 (N_30610,N_25061,N_21327);
and U30611 (N_30611,N_23362,N_24279);
nand U30612 (N_30612,N_20080,N_29605);
nor U30613 (N_30613,N_26522,N_26815);
nor U30614 (N_30614,N_24831,N_20686);
nor U30615 (N_30615,N_24782,N_20260);
nand U30616 (N_30616,N_22559,N_20254);
nor U30617 (N_30617,N_26307,N_26246);
xnor U30618 (N_30618,N_21363,N_23540);
or U30619 (N_30619,N_20904,N_23101);
and U30620 (N_30620,N_20383,N_27390);
or U30621 (N_30621,N_27750,N_23403);
nor U30622 (N_30622,N_20083,N_25651);
xor U30623 (N_30623,N_20507,N_25099);
or U30624 (N_30624,N_21955,N_29498);
nand U30625 (N_30625,N_20725,N_22935);
nand U30626 (N_30626,N_23870,N_27172);
xor U30627 (N_30627,N_21070,N_29772);
and U30628 (N_30628,N_23141,N_23796);
and U30629 (N_30629,N_26892,N_28796);
xor U30630 (N_30630,N_22863,N_21894);
nor U30631 (N_30631,N_25859,N_21256);
and U30632 (N_30632,N_23490,N_22843);
or U30633 (N_30633,N_22743,N_27043);
nor U30634 (N_30634,N_27312,N_21529);
xnor U30635 (N_30635,N_29530,N_28295);
or U30636 (N_30636,N_22862,N_22614);
nor U30637 (N_30637,N_29504,N_24823);
nor U30638 (N_30638,N_28162,N_29358);
and U30639 (N_30639,N_27097,N_26785);
nand U30640 (N_30640,N_28853,N_26819);
xnor U30641 (N_30641,N_29879,N_28385);
nor U30642 (N_30642,N_20258,N_29013);
nor U30643 (N_30643,N_29857,N_29666);
xor U30644 (N_30644,N_25469,N_26198);
and U30645 (N_30645,N_25247,N_23173);
xnor U30646 (N_30646,N_20545,N_27702);
or U30647 (N_30647,N_26269,N_21766);
nor U30648 (N_30648,N_21992,N_24613);
nor U30649 (N_30649,N_27841,N_29208);
nand U30650 (N_30650,N_28371,N_25717);
nand U30651 (N_30651,N_26729,N_21489);
nor U30652 (N_30652,N_24386,N_27882);
nand U30653 (N_30653,N_21664,N_26373);
and U30654 (N_30654,N_21386,N_22004);
xnor U30655 (N_30655,N_22327,N_27632);
xnor U30656 (N_30656,N_27789,N_20828);
or U30657 (N_30657,N_22343,N_22783);
nand U30658 (N_30658,N_29370,N_23595);
or U30659 (N_30659,N_22670,N_20149);
nand U30660 (N_30660,N_24142,N_24525);
nor U30661 (N_30661,N_25055,N_24964);
nor U30662 (N_30662,N_26961,N_23562);
or U30663 (N_30663,N_24466,N_28340);
nor U30664 (N_30664,N_25796,N_24166);
and U30665 (N_30665,N_22921,N_26818);
nor U30666 (N_30666,N_25856,N_25917);
xnor U30667 (N_30667,N_27951,N_23698);
xor U30668 (N_30668,N_22951,N_28552);
and U30669 (N_30669,N_27523,N_29161);
xnor U30670 (N_30670,N_25406,N_26151);
nor U30671 (N_30671,N_23862,N_20354);
nor U30672 (N_30672,N_25167,N_28194);
nor U30673 (N_30673,N_24006,N_22159);
or U30674 (N_30674,N_20889,N_21459);
xor U30675 (N_30675,N_21533,N_21214);
and U30676 (N_30676,N_26309,N_27488);
xor U30677 (N_30677,N_27192,N_28958);
or U30678 (N_30678,N_29044,N_27521);
xnor U30679 (N_30679,N_21729,N_29754);
and U30680 (N_30680,N_25386,N_22056);
nor U30681 (N_30681,N_21983,N_29717);
or U30682 (N_30682,N_21061,N_20271);
or U30683 (N_30683,N_20273,N_22075);
and U30684 (N_30684,N_26439,N_21038);
or U30685 (N_30685,N_23891,N_25359);
nand U30686 (N_30686,N_26774,N_22357);
and U30687 (N_30687,N_23535,N_26606);
and U30688 (N_30688,N_28215,N_25762);
and U30689 (N_30689,N_25524,N_26353);
nand U30690 (N_30690,N_27064,N_27699);
and U30691 (N_30691,N_29758,N_24138);
xnor U30692 (N_30692,N_20871,N_22048);
xnor U30693 (N_30693,N_23772,N_28261);
or U30694 (N_30694,N_24260,N_25095);
xor U30695 (N_30695,N_28271,N_27912);
or U30696 (N_30696,N_24794,N_25139);
and U30697 (N_30697,N_29913,N_21079);
nand U30698 (N_30698,N_24638,N_22705);
nand U30699 (N_30699,N_28591,N_23518);
or U30700 (N_30700,N_20832,N_26138);
and U30701 (N_30701,N_28354,N_26227);
or U30702 (N_30702,N_29374,N_29352);
or U30703 (N_30703,N_24482,N_26784);
and U30704 (N_30704,N_27130,N_23769);
and U30705 (N_30705,N_24883,N_24979);
or U30706 (N_30706,N_25256,N_25257);
and U30707 (N_30707,N_22607,N_29129);
or U30708 (N_30708,N_22316,N_25649);
nor U30709 (N_30709,N_25499,N_21909);
nand U30710 (N_30710,N_24557,N_28983);
xor U30711 (N_30711,N_24889,N_20360);
xor U30712 (N_30712,N_28218,N_29675);
nand U30713 (N_30713,N_21332,N_26898);
nand U30714 (N_30714,N_23497,N_23879);
and U30715 (N_30715,N_24928,N_23997);
and U30716 (N_30716,N_20375,N_28627);
or U30717 (N_30717,N_22243,N_25040);
nor U30718 (N_30718,N_25916,N_20153);
xor U30719 (N_30719,N_29172,N_24462);
or U30720 (N_30720,N_25007,N_27027);
nand U30721 (N_30721,N_24109,N_21575);
xor U30722 (N_30722,N_24768,N_22894);
nand U30723 (N_30723,N_28235,N_22661);
xor U30724 (N_30724,N_26359,N_29376);
or U30725 (N_30725,N_24200,N_24687);
or U30726 (N_30726,N_27675,N_21042);
nand U30727 (N_30727,N_26082,N_28121);
xnor U30728 (N_30728,N_28632,N_29684);
xnor U30729 (N_30729,N_28692,N_25824);
xor U30730 (N_30730,N_28737,N_28604);
nor U30731 (N_30731,N_27001,N_27609);
and U30732 (N_30732,N_22836,N_27251);
and U30733 (N_30733,N_20777,N_20428);
or U30734 (N_30734,N_26180,N_20029);
nand U30735 (N_30735,N_23789,N_23340);
nand U30736 (N_30736,N_24726,N_21755);
xor U30737 (N_30737,N_29983,N_29542);
nand U30738 (N_30738,N_21284,N_25042);
and U30739 (N_30739,N_24588,N_24028);
or U30740 (N_30740,N_25716,N_24531);
xor U30741 (N_30741,N_20236,N_25262);
or U30742 (N_30742,N_26277,N_26643);
or U30743 (N_30743,N_28830,N_23524);
or U30744 (N_30744,N_21187,N_28013);
and U30745 (N_30745,N_28280,N_24059);
or U30746 (N_30746,N_27048,N_29562);
nor U30747 (N_30747,N_28602,N_26124);
nor U30748 (N_30748,N_24604,N_22143);
or U30749 (N_30749,N_27577,N_24637);
or U30750 (N_30750,N_25749,N_24091);
nand U30751 (N_30751,N_29696,N_27713);
or U30752 (N_30752,N_20819,N_24339);
nor U30753 (N_30753,N_24285,N_23439);
or U30754 (N_30754,N_22794,N_20975);
nor U30755 (N_30755,N_24467,N_25510);
xor U30756 (N_30756,N_26465,N_28476);
and U30757 (N_30757,N_24115,N_20321);
nor U30758 (N_30758,N_21088,N_26089);
or U30759 (N_30759,N_27801,N_22341);
or U30760 (N_30760,N_27802,N_22887);
and U30761 (N_30761,N_22880,N_23776);
xor U30762 (N_30762,N_22034,N_29369);
nand U30763 (N_30763,N_28222,N_27304);
or U30764 (N_30764,N_28355,N_27904);
nor U30765 (N_30765,N_26788,N_29745);
nand U30766 (N_30766,N_21878,N_21113);
xnor U30767 (N_30767,N_28097,N_21368);
nor U30768 (N_30768,N_24034,N_29672);
xnor U30769 (N_30769,N_20277,N_29662);
and U30770 (N_30770,N_29583,N_21811);
nor U30771 (N_30771,N_22540,N_25655);
or U30772 (N_30772,N_25839,N_23904);
nand U30773 (N_30773,N_28842,N_26631);
and U30774 (N_30774,N_20262,N_21023);
nand U30775 (N_30775,N_20509,N_25673);
xor U30776 (N_30776,N_22653,N_20927);
or U30777 (N_30777,N_22466,N_28216);
or U30778 (N_30778,N_21169,N_20200);
or U30779 (N_30779,N_29105,N_25197);
or U30780 (N_30780,N_26746,N_26511);
and U30781 (N_30781,N_28952,N_25866);
and U30782 (N_30782,N_28382,N_20947);
and U30783 (N_30783,N_24574,N_20969);
nor U30784 (N_30784,N_28662,N_21594);
nor U30785 (N_30785,N_21773,N_28282);
and U30786 (N_30786,N_26695,N_20075);
and U30787 (N_30787,N_23045,N_22183);
and U30788 (N_30788,N_27117,N_24767);
nor U30789 (N_30789,N_21352,N_29736);
nor U30790 (N_30790,N_22890,N_21021);
or U30791 (N_30791,N_25957,N_22778);
xor U30792 (N_30792,N_20174,N_27965);
or U30793 (N_30793,N_23276,N_23800);
nor U30794 (N_30794,N_27580,N_20219);
nand U30795 (N_30795,N_24310,N_27406);
and U30796 (N_30796,N_27969,N_22157);
and U30797 (N_30797,N_22014,N_20968);
nor U30798 (N_30798,N_29371,N_20789);
nor U30799 (N_30799,N_24536,N_29492);
nand U30800 (N_30800,N_21704,N_21721);
xnor U30801 (N_30801,N_25823,N_21994);
nand U30802 (N_30802,N_21127,N_23960);
xor U30803 (N_30803,N_21277,N_25885);
nor U30804 (N_30804,N_22113,N_25574);
nor U30805 (N_30805,N_28042,N_26742);
xor U30806 (N_30806,N_27022,N_26510);
nor U30807 (N_30807,N_24358,N_27751);
xor U30808 (N_30808,N_24555,N_24798);
xnor U30809 (N_30809,N_27851,N_25723);
xor U30810 (N_30810,N_28130,N_26901);
or U30811 (N_30811,N_24680,N_20559);
nor U30812 (N_30812,N_23099,N_29552);
or U30813 (N_30813,N_27550,N_23715);
nand U30814 (N_30814,N_21713,N_23651);
xnor U30815 (N_30815,N_26752,N_29140);
nand U30816 (N_30816,N_26237,N_28734);
xor U30817 (N_30817,N_22269,N_27979);
xor U30818 (N_30818,N_25733,N_22340);
xnor U30819 (N_30819,N_22308,N_23292);
xor U30820 (N_30820,N_21151,N_21428);
xor U30821 (N_30821,N_28972,N_20454);
and U30822 (N_30822,N_21567,N_25059);
xor U30823 (N_30823,N_20844,N_21568);
xor U30824 (N_30824,N_21448,N_21527);
or U30825 (N_30825,N_27786,N_29158);
nand U30826 (N_30826,N_29661,N_22203);
nor U30827 (N_30827,N_23278,N_29246);
or U30828 (N_30828,N_28929,N_24829);
nor U30829 (N_30829,N_20205,N_27924);
and U30830 (N_30830,N_21037,N_25827);
nor U30831 (N_30831,N_26248,N_25421);
or U30832 (N_30832,N_21752,N_22564);
or U30833 (N_30833,N_25696,N_29638);
and U30834 (N_30834,N_28154,N_29548);
and U30835 (N_30835,N_24069,N_22364);
nand U30836 (N_30836,N_28026,N_27082);
xor U30837 (N_30837,N_27333,N_23450);
and U30838 (N_30838,N_25766,N_24449);
xnor U30839 (N_30839,N_23102,N_26962);
or U30840 (N_30840,N_23274,N_29644);
or U30841 (N_30841,N_22463,N_23216);
nor U30842 (N_30842,N_22367,N_25741);
or U30843 (N_30843,N_24919,N_28359);
or U30844 (N_30844,N_29916,N_22350);
xnor U30845 (N_30845,N_25551,N_28789);
or U30846 (N_30846,N_25328,N_23384);
and U30847 (N_30847,N_27764,N_21705);
nand U30848 (N_30848,N_29247,N_24411);
nor U30849 (N_30849,N_21658,N_22931);
nand U30850 (N_30850,N_28750,N_24400);
xor U30851 (N_30851,N_27046,N_20849);
or U30852 (N_30852,N_28863,N_29820);
xnor U30853 (N_30853,N_23892,N_28869);
and U30854 (N_30854,N_26123,N_26920);
and U30855 (N_30855,N_25087,N_29125);
nand U30856 (N_30856,N_20973,N_20867);
and U30857 (N_30857,N_22954,N_23472);
nor U30858 (N_30858,N_29029,N_21875);
nor U30859 (N_30859,N_29333,N_21020);
and U30860 (N_30860,N_23194,N_25337);
nor U30861 (N_30861,N_25584,N_29868);
or U30862 (N_30862,N_20054,N_22495);
xnor U30863 (N_30863,N_25846,N_23910);
or U30864 (N_30864,N_25768,N_26663);
and U30865 (N_30865,N_26835,N_22895);
xor U30866 (N_30866,N_28836,N_27652);
and U30867 (N_30867,N_23912,N_27905);
nor U30868 (N_30868,N_27959,N_25030);
xor U30869 (N_30869,N_23935,N_22719);
or U30870 (N_30870,N_26780,N_26178);
or U30871 (N_30871,N_24143,N_28780);
xor U30872 (N_30872,N_28565,N_29490);
nor U30873 (N_30873,N_28666,N_23878);
xor U30874 (N_30874,N_26226,N_29494);
or U30875 (N_30875,N_22011,N_20735);
and U30876 (N_30876,N_28064,N_24591);
or U30877 (N_30877,N_21532,N_27687);
or U30878 (N_30878,N_21519,N_24916);
nor U30879 (N_30879,N_27376,N_22764);
xor U30880 (N_30880,N_29071,N_23947);
xor U30881 (N_30881,N_20177,N_26030);
nand U30882 (N_30882,N_29687,N_29256);
or U30883 (N_30883,N_21656,N_20541);
nand U30884 (N_30884,N_28533,N_23571);
nand U30885 (N_30885,N_24047,N_20059);
nand U30886 (N_30886,N_21445,N_29833);
nor U30887 (N_30887,N_29873,N_21223);
nand U30888 (N_30888,N_26676,N_26336);
and U30889 (N_30889,N_28981,N_21944);
nand U30890 (N_30890,N_26945,N_25915);
and U30891 (N_30891,N_25692,N_26279);
or U30892 (N_30892,N_22620,N_25222);
or U30893 (N_30893,N_26814,N_22097);
nand U30894 (N_30894,N_25753,N_26505);
and U30895 (N_30895,N_27805,N_29863);
or U30896 (N_30896,N_20521,N_20445);
or U30897 (N_30897,N_23259,N_26543);
or U30898 (N_30898,N_23092,N_21082);
and U30899 (N_30899,N_27009,N_22538);
nand U30900 (N_30900,N_24926,N_27370);
or U30901 (N_30901,N_20809,N_23810);
or U30902 (N_30902,N_23964,N_23750);
nand U30903 (N_30903,N_29564,N_28266);
or U30904 (N_30904,N_25563,N_23023);
and U30905 (N_30905,N_29808,N_28793);
xnor U30906 (N_30906,N_26891,N_26853);
nand U30907 (N_30907,N_25984,N_25016);
nand U30908 (N_30908,N_26378,N_27621);
or U30909 (N_30909,N_21961,N_29293);
and U30910 (N_30910,N_22479,N_21463);
and U30911 (N_30911,N_28966,N_24430);
nor U30912 (N_30912,N_20385,N_22566);
or U30913 (N_30913,N_24631,N_27070);
xnor U30914 (N_30914,N_23149,N_29914);
and U30915 (N_30915,N_24253,N_22493);
nand U30916 (N_30916,N_22116,N_28228);
or U30917 (N_30917,N_20793,N_23138);
or U30918 (N_30918,N_27929,N_27934);
nor U30919 (N_30919,N_20490,N_27645);
nor U30920 (N_30920,N_28277,N_22989);
xnor U30921 (N_30921,N_24407,N_21030);
nor U30922 (N_30922,N_24320,N_29778);
or U30923 (N_30923,N_25352,N_21745);
nor U30924 (N_30924,N_25702,N_21967);
and U30925 (N_30925,N_27622,N_22515);
xnor U30926 (N_30926,N_26650,N_21036);
nand U30927 (N_30927,N_26114,N_23683);
nor U30928 (N_30928,N_22304,N_29678);
nand U30929 (N_30929,N_29532,N_22815);
or U30930 (N_30930,N_26925,N_25043);
nand U30931 (N_30931,N_27007,N_20010);
or U30932 (N_30932,N_21466,N_27316);
and U30933 (N_30933,N_28590,N_28079);
nand U30934 (N_30934,N_26243,N_29529);
xor U30935 (N_30935,N_29936,N_25511);
xnor U30936 (N_30936,N_23839,N_21842);
nand U30937 (N_30937,N_24564,N_22005);
and U30938 (N_30938,N_25143,N_29920);
nand U30939 (N_30939,N_28061,N_26165);
nand U30940 (N_30940,N_27238,N_27138);
xor U30941 (N_30941,N_23883,N_20797);
or U30942 (N_30942,N_26521,N_23308);
xor U30943 (N_30943,N_22514,N_24405);
nor U30944 (N_30944,N_20957,N_20574);
nor U30945 (N_30945,N_21179,N_20338);
or U30946 (N_30946,N_23379,N_25903);
nor U30947 (N_30947,N_22398,N_22878);
nand U30948 (N_30948,N_27024,N_20546);
nor U30949 (N_30949,N_20629,N_24127);
and U30950 (N_30950,N_24128,N_20781);
nor U30951 (N_30951,N_25549,N_29715);
nand U30952 (N_30952,N_21915,N_29854);
nor U30953 (N_30953,N_26472,N_27021);
nand U30954 (N_30954,N_27371,N_26730);
nor U30955 (N_30955,N_25788,N_26201);
or U30956 (N_30956,N_26335,N_28192);
or U30957 (N_30957,N_21786,N_20040);
xnor U30958 (N_30958,N_21655,N_20940);
or U30959 (N_30959,N_20301,N_29641);
nor U30960 (N_30960,N_21056,N_25100);
and U30961 (N_30961,N_22471,N_27684);
and U30962 (N_30962,N_29200,N_21898);
and U30963 (N_30963,N_20015,N_23407);
and U30964 (N_30964,N_20424,N_29795);
and U30965 (N_30965,N_25891,N_23909);
nor U30966 (N_30966,N_27557,N_23917);
or U30967 (N_30967,N_23021,N_29080);
nand U30968 (N_30968,N_20641,N_20255);
or U30969 (N_30969,N_27105,N_20959);
nand U30970 (N_30970,N_22028,N_24261);
nand U30971 (N_30971,N_25410,N_25362);
and U30972 (N_30972,N_29180,N_25316);
nand U30973 (N_30973,N_20887,N_27107);
nor U30974 (N_30974,N_25769,N_21971);
nand U30975 (N_30975,N_20501,N_29493);
xor U30976 (N_30976,N_29126,N_29064);
and U30977 (N_30977,N_20090,N_22110);
or U30978 (N_30978,N_20311,N_21880);
nand U30979 (N_30979,N_21639,N_27853);
or U30980 (N_30980,N_21484,N_28786);
and U30981 (N_30981,N_20171,N_24073);
nand U30982 (N_30982,N_26481,N_28272);
nand U30983 (N_30983,N_25750,N_22964);
nand U30984 (N_30984,N_22804,N_26813);
or U30985 (N_30985,N_28940,N_25138);
nand U30986 (N_30986,N_21598,N_25206);
nand U30987 (N_30987,N_21728,N_28500);
xnor U30988 (N_30988,N_22869,N_22251);
nor U30989 (N_30989,N_22093,N_20875);
or U30990 (N_30990,N_29452,N_28263);
nand U30991 (N_30991,N_27095,N_29917);
xnor U30992 (N_30992,N_26344,N_22161);
nand U30993 (N_30993,N_24612,N_22599);
or U30994 (N_30994,N_23281,N_26877);
nand U30995 (N_30995,N_26541,N_28645);
and U30996 (N_30996,N_28680,N_29327);
xnor U30997 (N_30997,N_27738,N_22213);
or U30998 (N_30998,N_27981,N_24454);
nand U30999 (N_30999,N_26966,N_26206);
xnor U31000 (N_31000,N_26886,N_21071);
nor U31001 (N_31001,N_24227,N_26830);
xnor U31002 (N_31002,N_28770,N_22169);
xor U31003 (N_31003,N_27915,N_25452);
nor U31004 (N_31004,N_20025,N_28726);
and U31005 (N_31005,N_21181,N_29545);
or U31006 (N_31006,N_26209,N_28043);
xnor U31007 (N_31007,N_29340,N_22497);
nand U31008 (N_31008,N_22982,N_27480);
nor U31009 (N_31009,N_20497,N_28664);
nand U31010 (N_31010,N_29697,N_29958);
nand U31011 (N_31011,N_29550,N_22206);
and U31012 (N_31012,N_29905,N_20796);
nand U31013 (N_31013,N_22092,N_24949);
and U31014 (N_31014,N_20942,N_25155);
or U31015 (N_31015,N_26403,N_23532);
nor U31016 (N_31016,N_23129,N_29173);
or U31017 (N_31017,N_27511,N_24364);
nor U31018 (N_31018,N_20949,N_27358);
or U31019 (N_31019,N_23603,N_23294);
xor U31020 (N_31020,N_23142,N_24211);
nor U31021 (N_31021,N_20362,N_22688);
nor U31022 (N_31022,N_25215,N_27873);
and U31023 (N_31023,N_25266,N_25218);
nor U31024 (N_31024,N_23399,N_27903);
nand U31025 (N_31025,N_26608,N_27696);
and U31026 (N_31026,N_22120,N_26924);
and U31027 (N_31027,N_23069,N_29084);
nand U31028 (N_31028,N_24960,N_21683);
xnor U31029 (N_31029,N_24343,N_28482);
xnor U31030 (N_31030,N_25370,N_29615);
nor U31031 (N_31031,N_26934,N_20453);
xnor U31032 (N_31032,N_23855,N_25671);
and U31033 (N_31033,N_23201,N_25851);
nor U31034 (N_31034,N_20527,N_20530);
nand U31035 (N_31035,N_25005,N_25617);
nand U31036 (N_31036,N_23451,N_24932);
and U31037 (N_31037,N_20105,N_20993);
nand U31038 (N_31038,N_28931,N_27407);
nor U31039 (N_31039,N_25566,N_23075);
or U31040 (N_31040,N_28729,N_24187);
and U31041 (N_31041,N_29888,N_22323);
or U31042 (N_31042,N_29259,N_22274);
xnor U31043 (N_31043,N_28777,N_24251);
nor U31044 (N_31044,N_22429,N_28139);
xor U31045 (N_31045,N_22787,N_22855);
nor U31046 (N_31046,N_24967,N_25906);
nor U31047 (N_31047,N_28339,N_28801);
xnor U31048 (N_31048,N_26052,N_23109);
and U31049 (N_31049,N_21852,N_24901);
nor U31050 (N_31050,N_20537,N_27399);
xnor U31051 (N_31051,N_23841,N_29505);
and U31052 (N_31052,N_21663,N_21928);
and U31053 (N_31053,N_23743,N_29784);
nand U31054 (N_31054,N_26189,N_26447);
or U31055 (N_31055,N_28469,N_23505);
xnor U31056 (N_31056,N_27935,N_27846);
and U31057 (N_31057,N_27662,N_25375);
nand U31058 (N_31058,N_22851,N_24861);
xor U31059 (N_31059,N_27567,N_29897);
nor U31060 (N_31060,N_25530,N_29884);
or U31061 (N_31061,N_27176,N_27045);
nor U31062 (N_31062,N_24232,N_23137);
and U31063 (N_31063,N_28752,N_25160);
xnor U31064 (N_31064,N_20946,N_28781);
or U31065 (N_31065,N_27907,N_26188);
and U31066 (N_31066,N_25603,N_29892);
nor U31067 (N_31067,N_22561,N_22773);
and U31068 (N_31068,N_29975,N_21259);
xor U31069 (N_31069,N_21199,N_23305);
nand U31070 (N_31070,N_28629,N_29269);
and U31071 (N_31071,N_28012,N_27990);
nor U31072 (N_31072,N_21101,N_22602);
nor U31073 (N_31073,N_29227,N_20673);
and U31074 (N_31074,N_24171,N_25523);
nand U31075 (N_31075,N_25004,N_28430);
and U31076 (N_31076,N_21129,N_21978);
and U31077 (N_31077,N_24345,N_24933);
xor U31078 (N_31078,N_26076,N_20159);
or U31079 (N_31079,N_28107,N_28203);
nand U31080 (N_31080,N_24651,N_27363);
nor U31081 (N_31081,N_22598,N_23923);
and U31082 (N_31082,N_20635,N_21255);
and U31083 (N_31083,N_24506,N_27272);
xor U31084 (N_31084,N_23895,N_25751);
xnor U31085 (N_31085,N_28703,N_26694);
and U31086 (N_31086,N_24719,N_27218);
nor U31087 (N_31087,N_22459,N_20127);
xor U31088 (N_31088,N_21577,N_20627);
or U31089 (N_31089,N_24586,N_28109);
xor U31090 (N_31090,N_23161,N_28387);
nand U31091 (N_31091,N_23641,N_20624);
nand U31092 (N_31092,N_26664,N_22498);
nand U31093 (N_31093,N_23934,N_23768);
and U31094 (N_31094,N_28120,N_28440);
nand U31095 (N_31095,N_28641,N_27360);
nand U31096 (N_31096,N_26938,N_20711);
and U31097 (N_31097,N_26182,N_29391);
nand U31098 (N_31098,N_24943,N_21110);
nand U31099 (N_31099,N_27339,N_20806);
xnor U31100 (N_31100,N_29794,N_21171);
xnor U31101 (N_31101,N_26211,N_23198);
and U31102 (N_31102,N_29827,N_29127);
xnor U31103 (N_31103,N_25512,N_29710);
and U31104 (N_31104,N_29367,N_23036);
and U31105 (N_31105,N_21453,N_24770);
or U31106 (N_31106,N_20069,N_21608);
nor U31107 (N_31107,N_28095,N_20837);
and U31108 (N_31108,N_27832,N_25301);
nor U31109 (N_31109,N_25056,N_29618);
nand U31110 (N_31110,N_26104,N_27661);
xnor U31111 (N_31111,N_23170,N_20646);
or U31112 (N_31112,N_23348,N_22475);
xnor U31113 (N_31113,N_28790,N_25911);
nand U31114 (N_31114,N_25388,N_25931);
or U31115 (N_31115,N_21422,N_29258);
nor U31116 (N_31116,N_25272,N_28991);
nor U31117 (N_31117,N_20523,N_24254);
nor U31118 (N_31118,N_26204,N_21314);
or U31119 (N_31119,N_22219,N_28240);
nor U31120 (N_31120,N_22673,N_20589);
nor U31121 (N_31121,N_23481,N_29728);
or U31122 (N_31122,N_22991,N_22458);
nand U31123 (N_31123,N_24342,N_25791);
and U31124 (N_31124,N_24267,N_26684);
xnor U31125 (N_31125,N_27466,N_25263);
and U31126 (N_31126,N_22082,N_29444);
nand U31127 (N_31127,N_20279,N_29516);
nor U31128 (N_31128,N_21914,N_27732);
and U31129 (N_31129,N_21491,N_28531);
or U31130 (N_31130,N_25124,N_26492);
or U31131 (N_31131,N_26636,N_22754);
and U31132 (N_31132,N_24473,N_21965);
or U31133 (N_31133,N_29624,N_27057);
xnor U31134 (N_31134,N_29674,N_29348);
xor U31135 (N_31135,N_25349,N_28219);
and U31136 (N_31136,N_29755,N_25647);
and U31137 (N_31137,N_20987,N_20743);
or U31138 (N_31138,N_23449,N_23958);
xnor U31139 (N_31139,N_28214,N_24433);
xor U31140 (N_31140,N_25051,N_23421);
nor U31141 (N_31141,N_26653,N_26438);
or U31142 (N_31142,N_25084,N_20178);
and U31143 (N_31143,N_23240,N_25635);
and U31144 (N_31144,N_24136,N_24542);
nand U31145 (N_31145,N_23591,N_25638);
or U31146 (N_31146,N_25742,N_26146);
nand U31147 (N_31147,N_28017,N_20425);
and U31148 (N_31148,N_24455,N_20872);
or U31149 (N_31149,N_22315,N_25718);
nor U31150 (N_31150,N_27263,N_27545);
nand U31151 (N_31151,N_28659,N_26046);
xor U31152 (N_31152,N_26674,N_21630);
and U31153 (N_31153,N_20938,N_26681);
nand U31154 (N_31154,N_21400,N_26715);
nand U31155 (N_31155,N_20900,N_24365);
nand U31156 (N_31156,N_21649,N_22933);
nor U31157 (N_31157,N_21073,N_28631);
or U31158 (N_31158,N_25497,N_21905);
and U31159 (N_31159,N_20092,N_28669);
xor U31160 (N_31160,N_21881,N_26348);
and U31161 (N_31161,N_28204,N_20340);
nand U31162 (N_31162,N_25997,N_24202);
xnor U31163 (N_31163,N_24153,N_23444);
or U31164 (N_31164,N_20753,N_21136);
xor U31165 (N_31165,N_20420,N_20576);
or U31166 (N_31166,N_21378,N_28205);
nand U31167 (N_31167,N_21751,N_20861);
xor U31168 (N_31168,N_26191,N_29727);
xnor U31169 (N_31169,N_26270,N_20136);
or U31170 (N_31170,N_22524,N_27366);
xnor U31171 (N_31171,N_22469,N_29017);
or U31172 (N_31172,N_28665,N_20183);
nor U31173 (N_31173,N_28193,N_21190);
or U31174 (N_31174,N_28784,N_29779);
and U31175 (N_31175,N_23717,N_29386);
or U31176 (N_31176,N_20398,N_20924);
xnor U31177 (N_31177,N_24995,N_25719);
or U31178 (N_31178,N_26910,N_23183);
and U31179 (N_31179,N_22433,N_28575);
xor U31180 (N_31180,N_29094,N_26496);
and U31181 (N_31181,N_23252,N_23086);
nand U31182 (N_31182,N_29392,N_26097);
xor U31183 (N_31183,N_28819,N_28275);
nand U31184 (N_31184,N_26761,N_29077);
and U31185 (N_31185,N_26401,N_26696);
nand U31186 (N_31186,N_29388,N_27493);
nor U31187 (N_31187,N_22786,N_22600);
and U31188 (N_31188,N_21926,N_27646);
nand U31189 (N_31189,N_25683,N_27460);
nand U31190 (N_31190,N_28721,N_29010);
xor U31191 (N_31191,N_24853,N_24259);
xnor U31192 (N_31192,N_28564,N_28023);
xor U31193 (N_31193,N_26594,N_27429);
xnor U31194 (N_31194,N_22601,N_25460);
nand U31195 (N_31195,N_24677,N_24902);
nand U31196 (N_31196,N_29792,N_28585);
or U31197 (N_31197,N_23231,N_26749);
or U31198 (N_31198,N_23206,N_25178);
nor U31199 (N_31199,N_20726,N_20621);
nand U31200 (N_31200,N_29033,N_26133);
or U31201 (N_31201,N_25413,N_28390);
nor U31202 (N_31202,N_28810,N_25784);
and U31203 (N_31203,N_27680,N_25481);
and U31204 (N_31204,N_25567,N_29594);
xor U31205 (N_31205,N_20760,N_27756);
or U31206 (N_31206,N_28455,N_27340);
and U31207 (N_31207,N_24048,N_21839);
and U31208 (N_31208,N_29164,N_21475);
and U31209 (N_31209,N_27408,N_22544);
and U31210 (N_31210,N_22344,N_22303);
nand U31211 (N_31211,N_22918,N_25023);
or U31212 (N_31212,N_26612,N_29612);
xor U31213 (N_31213,N_22214,N_27445);
nor U31214 (N_31214,N_24589,N_28797);
nand U31215 (N_31215,N_24317,N_24897);
or U31216 (N_31216,N_27111,N_27930);
or U31217 (N_31217,N_23202,N_23263);
xor U31218 (N_31218,N_26020,N_25261);
xor U31219 (N_31219,N_20499,N_25562);
nand U31220 (N_31220,N_20870,N_21065);
or U31221 (N_31221,N_29691,N_22789);
and U31222 (N_31222,N_28268,N_22866);
nand U31223 (N_31223,N_22551,N_26252);
or U31224 (N_31224,N_29837,N_22623);
nand U31225 (N_31225,N_21796,N_23685);
or U31226 (N_31226,N_25849,N_23279);
xnor U31227 (N_31227,N_23833,N_20936);
nor U31228 (N_31228,N_26160,N_23412);
nor U31229 (N_31229,N_21827,N_20722);
and U31230 (N_31230,N_22795,N_25026);
xor U31231 (N_31231,N_22944,N_27014);
nor U31232 (N_31232,N_22545,N_27825);
xor U31233 (N_31233,N_23208,N_26486);
and U31234 (N_31234,N_24838,N_23434);
or U31235 (N_31235,N_22178,N_25773);
or U31236 (N_31236,N_26461,N_21406);
nor U31237 (N_31237,N_29360,N_28426);
nor U31238 (N_31238,N_25517,N_26549);
nand U31239 (N_31239,N_28065,N_20841);
xor U31240 (N_31240,N_28758,N_25189);
or U31241 (N_31241,N_21162,N_24126);
nor U31242 (N_31242,N_25921,N_21838);
nand U31243 (N_31243,N_24221,N_28778);
xnor U31244 (N_31244,N_22919,N_20814);
and U31245 (N_31245,N_20538,N_23607);
or U31246 (N_31246,N_23718,N_27435);
nor U31247 (N_31247,N_24915,N_25412);
xor U31248 (N_31248,N_20571,N_25487);
xnor U31249 (N_31249,N_26512,N_28610);
and U31250 (N_31250,N_27260,N_20296);
xnor U31251 (N_31251,N_22037,N_28246);
nand U31252 (N_31252,N_26876,N_25970);
or U31253 (N_31253,N_21228,N_20657);
nor U31254 (N_31254,N_24196,N_22499);
or U31255 (N_31255,N_21189,N_23047);
nor U31256 (N_31256,N_23849,N_21579);
nor U31257 (N_31257,N_26363,N_23264);
xor U31258 (N_31258,N_23417,N_21305);
or U31259 (N_31259,N_26470,N_27350);
nor U31260 (N_31260,N_22085,N_24450);
nor U31261 (N_31261,N_26978,N_27393);
xor U31262 (N_31262,N_29679,N_23701);
nand U31263 (N_31263,N_27347,N_26547);
nand U31264 (N_31264,N_20148,N_23516);
nor U31265 (N_31265,N_28562,N_20039);
nor U31266 (N_31266,N_20939,N_22941);
or U31267 (N_31267,N_28132,N_28614);
nand U31268 (N_31268,N_26387,N_23392);
xnor U31269 (N_31269,N_26708,N_27735);
nor U31270 (N_31270,N_23475,N_24011);
xor U31271 (N_31271,N_28345,N_25745);
nand U31272 (N_31272,N_29006,N_22984);
nor U31273 (N_31273,N_25994,N_22395);
nor U31274 (N_31274,N_25805,N_26974);
and U31275 (N_31275,N_22318,N_26651);
nand U31276 (N_31276,N_29864,N_29534);
nor U31277 (N_31277,N_27219,N_26590);
nand U31278 (N_31278,N_22985,N_20126);
xnor U31279 (N_31279,N_24532,N_21366);
xor U31280 (N_31280,N_20836,N_22080);
nor U31281 (N_31281,N_24888,N_23731);
xnor U31282 (N_31282,N_21072,N_20958);
nor U31283 (N_31283,N_21168,N_27734);
xor U31284 (N_31284,N_23052,N_26545);
nand U31285 (N_31285,N_26174,N_27357);
or U31286 (N_31286,N_24440,N_24539);
and U31287 (N_31287,N_25976,N_21873);
nor U31288 (N_31288,N_26504,N_26428);
nand U31289 (N_31289,N_21050,N_24844);
xnor U31290 (N_31290,N_26903,N_22613);
nor U31291 (N_31291,N_20591,N_21933);
xnor U31292 (N_31292,N_25688,N_24569);
nand U31293 (N_31293,N_25303,N_25505);
nor U31294 (N_31294,N_28320,N_27212);
and U31295 (N_31295,N_29565,N_20584);
and U31296 (N_31296,N_24403,N_21793);
or U31297 (N_31297,N_20728,N_24484);
and U31298 (N_31298,N_28328,N_25199);
nand U31299 (N_31299,N_21341,N_20772);
xnor U31300 (N_31300,N_24356,N_26942);
nor U31301 (N_31301,N_26155,N_28337);
nand U31302 (N_31302,N_26977,N_22336);
nand U31303 (N_31303,N_26683,N_29769);
nand U31304 (N_31304,N_26864,N_24470);
nand U31305 (N_31305,N_21315,N_27870);
nand U31306 (N_31306,N_24326,N_23502);
nand U31307 (N_31307,N_29115,N_24265);
nand U31308 (N_31308,N_21780,N_22814);
nor U31309 (N_31309,N_22955,N_25064);
nor U31310 (N_31310,N_27626,N_26291);
and U31311 (N_31311,N_25786,N_22761);
xnor U31312 (N_31312,N_23506,N_28776);
and U31313 (N_31313,N_22905,N_22900);
or U31314 (N_31314,N_26748,N_27348);
and U31315 (N_31315,N_23463,N_24180);
xnor U31316 (N_31316,N_25594,N_21604);
xnor U31317 (N_31317,N_25643,N_24081);
nor U31318 (N_31318,N_21112,N_27191);
or U31319 (N_31319,N_26603,N_27956);
nor U31320 (N_31320,N_29334,N_24360);
nor U31321 (N_31321,N_28912,N_29092);
or U31322 (N_31322,N_25162,N_25698);
nand U31323 (N_31323,N_21355,N_21607);
nand U31324 (N_31324,N_20303,N_27248);
nand U31325 (N_31325,N_20115,N_27587);
and U31326 (N_31326,N_23673,N_25767);
nor U31327 (N_31327,N_23581,N_23601);
and U31328 (N_31328,N_29924,N_28816);
nor U31329 (N_31329,N_27137,N_21936);
xor U31330 (N_31330,N_26448,N_26789);
and U31331 (N_31331,N_24934,N_29999);
and U31332 (N_31332,N_20227,N_25425);
nor U31333 (N_31333,N_27859,N_25710);
and U31334 (N_31334,N_22353,N_20326);
or U31335 (N_31335,N_23747,N_21338);
xnor U31336 (N_31336,N_29489,N_20035);
or U31337 (N_31337,N_21720,N_21150);
nand U31338 (N_31338,N_20826,N_23803);
and U31339 (N_31339,N_23632,N_28101);
or U31340 (N_31340,N_23724,N_20220);
and U31341 (N_31341,N_24443,N_29440);
and U31342 (N_31342,N_29881,N_28202);
nand U31343 (N_31343,N_26721,N_26347);
nand U31344 (N_31344,N_26701,N_22784);
nand U31345 (N_31345,N_28322,N_26098);
nand U31346 (N_31346,N_28044,N_22129);
nand U31347 (N_31347,N_21777,N_20976);
nor U31348 (N_31348,N_27516,N_27617);
or U31349 (N_31349,N_24016,N_21938);
or U31350 (N_31350,N_23383,N_28380);
or U31351 (N_31351,N_29848,N_29050);
or U31352 (N_31352,N_22040,N_20032);
nor U31353 (N_31353,N_24043,N_20005);
and U31354 (N_31354,N_26714,N_25665);
nor U31355 (N_31355,N_21580,N_29773);
nor U31356 (N_31356,N_29268,N_21597);
or U31357 (N_31357,N_25321,N_28606);
nand U31358 (N_31358,N_24367,N_24751);
and U31359 (N_31359,N_20446,N_29774);
xnor U31360 (N_31360,N_20189,N_26026);
and U31361 (N_31361,N_23404,N_28615);
nand U31362 (N_31362,N_26882,N_27818);
nor U31363 (N_31363,N_23767,N_27714);
or U31364 (N_31364,N_20201,N_29456);
nor U31365 (N_31365,N_20195,N_22608);
or U31366 (N_31366,N_24991,N_20859);
and U31367 (N_31367,N_27168,N_28188);
and U31368 (N_31368,N_25797,N_25103);
nor U31369 (N_31369,N_21017,N_20432);
xnor U31370 (N_31370,N_29335,N_20824);
nand U31371 (N_31371,N_22812,N_20483);
nand U31372 (N_31372,N_25323,N_23794);
nor U31373 (N_31373,N_21005,N_20655);
or U31374 (N_31374,N_21326,N_26351);
and U31375 (N_31375,N_27109,N_22404);
xor U31376 (N_31376,N_22868,N_23570);
and U31377 (N_31377,N_20517,N_24118);
xor U31378 (N_31378,N_22410,N_25605);
nand U31379 (N_31379,N_21733,N_20931);
and U31380 (N_31380,N_20378,N_24655);
nand U31381 (N_31381,N_28916,N_22779);
nand U31382 (N_31382,N_28607,N_29341);
xnor U31383 (N_31383,N_23406,N_20954);
nor U31384 (N_31384,N_20784,N_27798);
and U31385 (N_31385,N_21334,N_22430);
and U31386 (N_31386,N_22832,N_25983);
nor U31387 (N_31387,N_21783,N_26874);
xor U31388 (N_31388,N_23903,N_24639);
nor U31389 (N_31389,N_23072,N_29204);
and U31390 (N_31390,N_29196,N_21719);
nor U31391 (N_31391,N_26313,N_21818);
xnor U31392 (N_31392,N_22671,N_25628);
or U31393 (N_31393,N_23233,N_28882);
and U31394 (N_31394,N_25752,N_21331);
nand U31395 (N_31395,N_23579,N_28508);
or U31396 (N_31396,N_23242,N_24493);
nor U31397 (N_31397,N_28524,N_28499);
xor U31398 (N_31398,N_24243,N_28164);
nand U31399 (N_31399,N_24428,N_27149);
nand U31400 (N_31400,N_24394,N_23300);
and U31401 (N_31401,N_20845,N_28865);
nand U31402 (N_31402,N_29992,N_28943);
nand U31403 (N_31403,N_20937,N_27505);
and U31404 (N_31404,N_27817,N_28677);
or U31405 (N_31405,N_21525,N_26432);
or U31406 (N_31406,N_21530,N_26524);
and U31407 (N_31407,N_22025,N_27718);
or U31408 (N_31408,N_24731,N_22946);
and U31409 (N_31409,N_22720,N_26069);
nor U31410 (N_31410,N_28145,N_23496);
nor U31411 (N_31411,N_21866,N_29328);
nor U31412 (N_31412,N_21514,N_29314);
and U31413 (N_31413,N_24635,N_20613);
nand U31414 (N_31414,N_21684,N_20166);
xor U31415 (N_31415,N_27344,N_28670);
nor U31416 (N_31416,N_20287,N_23373);
nor U31417 (N_31417,N_25174,N_28481);
nand U31418 (N_31418,N_25494,N_22124);
nor U31419 (N_31419,N_23865,N_23900);
xnor U31420 (N_31420,N_28151,N_22525);
nor U31421 (N_31421,N_27468,N_20966);
xor U31422 (N_31422,N_22134,N_21921);
or U31423 (N_31423,N_24245,N_23956);
nand U31424 (N_31424,N_27415,N_28892);
or U31425 (N_31425,N_23030,N_22817);
and U31426 (N_31426,N_24753,N_27895);
nor U31427 (N_31427,N_26060,N_26208);
nand U31428 (N_31428,N_22708,N_23106);
nand U31429 (N_31429,N_24811,N_26705);
xnor U31430 (N_31430,N_26333,N_26254);
xnor U31431 (N_31431,N_20622,N_23644);
nand U31432 (N_31432,N_28067,N_23661);
xor U31433 (N_31433,N_22748,N_20873);
nand U31434 (N_31434,N_20512,N_23438);
nor U31435 (N_31435,N_23906,N_27500);
and U31436 (N_31436,N_21690,N_22403);
or U31437 (N_31437,N_27970,N_21547);
xor U31438 (N_31438,N_20783,N_26558);
nor U31439 (N_31439,N_22205,N_24562);
or U31440 (N_31440,N_29325,N_21987);
or U31441 (N_31441,N_27167,N_24772);
nor U31442 (N_31442,N_22901,N_21307);
nor U31443 (N_31443,N_23063,N_21237);
nor U31444 (N_31444,N_22610,N_24291);
or U31445 (N_31445,N_22271,N_20216);
nor U31446 (N_31446,N_25676,N_25777);
nand U31447 (N_31447,N_29284,N_21052);
nand U31448 (N_31448,N_24067,N_22225);
xor U31449 (N_31449,N_24477,N_26392);
xnor U31450 (N_31450,N_29128,N_21520);
or U31451 (N_31451,N_23061,N_29668);
nor U31452 (N_31452,N_25310,N_25154);
xnor U31453 (N_31453,N_28055,N_22938);
and U31454 (N_31454,N_23227,N_24481);
nor U31455 (N_31455,N_26795,N_26340);
or U31456 (N_31456,N_27555,N_23793);
xor U31457 (N_31457,N_21395,N_25075);
nor U31458 (N_31458,N_26843,N_24711);
nor U31459 (N_31459,N_29692,N_23687);
and U31460 (N_31460,N_24749,N_22375);
or U31461 (N_31461,N_26136,N_27775);
xnor U31462 (N_31462,N_25727,N_25561);
nand U31463 (N_31463,N_24581,N_25223);
or U31464 (N_31464,N_29844,N_27025);
or U31465 (N_31465,N_20246,N_21454);
or U31466 (N_31466,N_29904,N_27833);
nand U31467 (N_31467,N_28288,N_25770);
and U31468 (N_31468,N_21874,N_25185);
nor U31469 (N_31469,N_26614,N_23898);
or U31470 (N_31470,N_29932,N_26225);
nand U31471 (N_31471,N_20003,N_24909);
xor U31472 (N_31472,N_20913,N_25912);
xor U31473 (N_31473,N_23799,N_23725);
and U31474 (N_31474,N_23007,N_25857);
nand U31475 (N_31475,N_26673,N_27954);
or U31476 (N_31476,N_29965,N_21152);
or U31477 (N_31477,N_24836,N_25164);
nand U31478 (N_31478,N_25736,N_26154);
xnor U31479 (N_31479,N_24822,N_28011);
nor U31480 (N_31480,N_26890,N_29345);
and U31481 (N_31481,N_27703,N_20854);
xor U31482 (N_31482,N_29654,N_26354);
xnor U31483 (N_31483,N_27225,N_28413);
nor U31484 (N_31484,N_23016,N_20288);
xor U31485 (N_31485,N_24215,N_22386);
xor U31486 (N_31486,N_22859,N_24441);
nor U31487 (N_31487,N_25083,N_28710);
xor U31488 (N_31488,N_27295,N_22527);
nor U31489 (N_31489,N_26262,N_26061);
nor U31490 (N_31490,N_29141,N_20099);
or U31491 (N_31491,N_28207,N_22220);
or U31492 (N_31492,N_21029,N_26964);
nand U31493 (N_31493,N_28243,N_23046);
or U31494 (N_31494,N_23257,N_27291);
nor U31495 (N_31495,N_23066,N_25949);
xor U31496 (N_31496,N_24576,N_28616);
or U31497 (N_31497,N_29742,N_21401);
xnor U31498 (N_31498,N_20592,N_23530);
and U31499 (N_31499,N_29987,N_28818);
or U31500 (N_31500,N_20780,N_22849);
nand U31501 (N_31501,N_25013,N_20961);
nor U31502 (N_31502,N_26660,N_21415);
nand U31503 (N_31503,N_21831,N_28939);
nor U31504 (N_31504,N_24743,N_25881);
nand U31505 (N_31505,N_20665,N_24519);
or U31506 (N_31506,N_22230,N_23834);
nor U31507 (N_31507,N_29102,N_25779);
nor U31508 (N_31508,N_20505,N_21025);
nand U31509 (N_31509,N_20252,N_22745);
xnor U31510 (N_31510,N_24159,N_21959);
xnor U31511 (N_31511,N_27814,N_26745);
nand U31512 (N_31512,N_20847,N_25068);
xnor U31513 (N_31513,N_22284,N_23557);
or U31514 (N_31514,N_21694,N_21676);
and U31515 (N_31515,N_21272,N_28724);
xnor U31516 (N_31516,N_28911,N_25306);
nand U31517 (N_31517,N_23299,N_21009);
nand U31518 (N_31518,N_21350,N_20366);
xor U31519 (N_31519,N_29655,N_25368);
or U31520 (N_31520,N_24066,N_22306);
xnor U31521 (N_31521,N_22017,N_28316);
nand U31522 (N_31522,N_22298,N_23054);
xor U31523 (N_31523,N_27513,N_26852);
nand U31524 (N_31524,N_24584,N_26183);
nand U31525 (N_31525,N_24704,N_27085);
nand U31526 (N_31526,N_25121,N_29045);
or U31527 (N_31527,N_27017,N_24188);
and U31528 (N_31528,N_22619,N_24976);
nand U31529 (N_31529,N_20916,N_23467);
nor U31530 (N_31530,N_21560,N_27126);
or U31531 (N_31531,N_28890,N_22006);
xor U31532 (N_31532,N_20122,N_23019);
nand U31533 (N_31533,N_27148,N_29223);
and U31534 (N_31534,N_23103,N_28030);
or U31535 (N_31535,N_27384,N_20088);
or U31536 (N_31536,N_23378,N_24551);
xor U31537 (N_31537,N_20295,N_24122);
and U31538 (N_31538,N_23874,N_28841);
or U31539 (N_31539,N_22122,N_23510);
nor U31540 (N_31540,N_22604,N_21473);
and U31541 (N_31541,N_25829,N_25539);
and U31542 (N_31542,N_20638,N_23684);
xor U31543 (N_31543,N_25444,N_21847);
xor U31544 (N_31544,N_26544,N_26989);
and U31545 (N_31545,N_23365,N_28959);
and U31546 (N_31546,N_24476,N_27098);
or U31547 (N_31547,N_28824,N_24341);
nand U31548 (N_31548,N_20650,N_28809);
nor U31549 (N_31549,N_29266,N_22156);
nand U31550 (N_31550,N_27204,N_21303);
and U31551 (N_31551,N_28106,N_22636);
or U31552 (N_31552,N_29214,N_21293);
and U31553 (N_31553,N_29763,N_26108);
nor U31554 (N_31554,N_29787,N_22628);
or U31555 (N_31555,N_20705,N_26698);
nor U31556 (N_31556,N_23323,N_20890);
nor U31557 (N_31557,N_23599,N_20765);
nor U31558 (N_31558,N_23364,N_22387);
or U31559 (N_31559,N_22769,N_25442);
nor U31560 (N_31560,N_20671,N_25390);
nand U31561 (N_31561,N_28388,N_26241);
and U31562 (N_31562,N_25320,N_29270);
and U31563 (N_31563,N_21450,N_21929);
and U31564 (N_31564,N_27710,N_20776);
nand U31565 (N_31565,N_20290,N_25815);
and U31566 (N_31566,N_26559,N_28530);
nor U31567 (N_31567,N_20448,N_23657);
xnor U31568 (N_31568,N_21469,N_23782);
xor U31569 (N_31569,N_21232,N_20985);
xnor U31570 (N_31570,N_29590,N_29783);
and U31571 (N_31571,N_29984,N_25018);
or U31572 (N_31572,N_23823,N_25977);
and U31573 (N_31573,N_27229,N_27839);
nand U31574 (N_31574,N_29944,N_22252);
xnor U31575 (N_31575,N_26677,N_27239);
nand U31576 (N_31576,N_28080,N_29389);
nand U31577 (N_31577,N_26963,N_22548);
or U31578 (N_31578,N_24041,N_27600);
nor U31579 (N_31579,N_28443,N_25798);
nand U31580 (N_31580,N_23366,N_29243);
nand U31581 (N_31581,N_23907,N_23177);
or U31582 (N_31582,N_21177,N_21084);
nor U31583 (N_31583,N_24657,N_26163);
nand U31584 (N_31584,N_27244,N_26670);
nor U31585 (N_31585,N_23393,N_26609);
nand U31586 (N_31586,N_20821,N_29229);
and U31587 (N_31587,N_29228,N_29142);
and U31588 (N_31588,N_24938,N_25022);
xor U31589 (N_31589,N_25184,N_25967);
and U31590 (N_31590,N_29089,N_21536);
nand U31591 (N_31591,N_29473,N_29512);
nor U31592 (N_31592,N_20894,N_27386);
or U31593 (N_31593,N_29401,N_21468);
or U31594 (N_31594,N_24954,N_26051);
xor U31595 (N_31595,N_24578,N_22766);
xor U31596 (N_31596,N_21251,N_22046);
nor U31597 (N_31597,N_21627,N_26798);
nand U31598 (N_31598,N_22397,N_22476);
xor U31599 (N_31599,N_27203,N_20165);
nor U31600 (N_31600,N_29601,N_28510);
or U31601 (N_31601,N_22767,N_21606);
and U31602 (N_31602,N_22847,N_27462);
or U31603 (N_31603,N_21276,N_21227);
and U31604 (N_31604,N_25624,N_28657);
xnor U31605 (N_31605,N_22571,N_27000);
nand U31606 (N_31606,N_24459,N_21521);
nand U31607 (N_31607,N_28081,N_23395);
xor U31608 (N_31608,N_24624,N_27972);
nand U31609 (N_31609,N_20372,N_23397);
and U31610 (N_31610,N_27655,N_25435);
nand U31611 (N_31611,N_29282,N_20249);
nand U31612 (N_31612,N_22725,N_24106);
nand U31613 (N_31613,N_22883,N_21710);
and U31614 (N_31614,N_26648,N_27572);
or U31615 (N_31615,N_20363,N_21235);
xor U31616 (N_31616,N_23429,N_26050);
and U31617 (N_31617,N_27667,N_27075);
nand U31618 (N_31618,N_20017,N_24150);
nand U31619 (N_31619,N_21109,N_20393);
nand U31620 (N_31620,N_20852,N_27721);
or U31621 (N_31621,N_28213,N_20052);
and U31622 (N_31622,N_24898,N_27815);
nor U31623 (N_31623,N_24633,N_27685);
nand U31624 (N_31624,N_28444,N_26662);
nand U31625 (N_31625,N_21119,N_27591);
nand U31626 (N_31626,N_27960,N_28864);
xor U31627 (N_31627,N_26084,N_23729);
nor U31628 (N_31628,N_24541,N_23783);
and U31629 (N_31629,N_28715,N_24644);
or U31630 (N_31630,N_26697,N_24891);
xor U31631 (N_31631,N_26904,N_22629);
xor U31632 (N_31632,N_29497,N_26944);
nor U31633 (N_31633,N_29698,N_25021);
nand U31634 (N_31634,N_26699,N_29373);
and U31635 (N_31635,N_22624,N_28208);
or U31636 (N_31636,N_22038,N_29224);
nor U31637 (N_31637,N_24887,N_27241);
or U31638 (N_31638,N_20062,N_20123);
xnor U31639 (N_31639,N_22590,N_22172);
and U31640 (N_31640,N_28982,N_20339);
nor U31641 (N_31641,N_29695,N_27049);
or U31642 (N_31642,N_29309,N_24445);
xor U31643 (N_31643,N_26464,N_27886);
nor U31644 (N_31644,N_27264,N_24620);
nand U31645 (N_31645,N_23559,N_26388);
nor U31646 (N_31646,N_25049,N_23195);
nand U31647 (N_31647,N_21825,N_24961);
nand U31648 (N_31648,N_29592,N_22328);
and U31649 (N_31649,N_20358,N_24355);
nor U31650 (N_31650,N_24671,N_24053);
and U31651 (N_31651,N_25996,N_24375);
nor U31652 (N_31652,N_28656,N_20923);
xor U31653 (N_31653,N_25858,N_29982);
nand U31654 (N_31654,N_25062,N_29031);
or U31655 (N_31655,N_27375,N_25229);
nand U31656 (N_31656,N_24796,N_25923);
or U31657 (N_31657,N_26583,N_26918);
xor U31658 (N_31658,N_23171,N_26736);
or U31659 (N_31659,N_28338,N_28142);
nand U31660 (N_31660,N_24771,N_28873);
nor U31661 (N_31661,N_23950,N_27943);
nor U31662 (N_31662,N_23067,N_27367);
xnor U31663 (N_31663,N_20774,N_29339);
and U31664 (N_31664,N_22647,N_27332);
xor U31665 (N_31665,N_26419,N_25780);
xor U31666 (N_31666,N_27876,N_21419);
and U31667 (N_31667,N_22867,N_22023);
and U31668 (N_31668,N_29964,N_22701);
or U31669 (N_31669,N_24262,N_23710);
nand U31670 (N_31670,N_29018,N_24560);
and U31671 (N_31671,N_25765,N_27556);
or U31672 (N_31672,N_20678,N_25001);
xnor U31673 (N_31673,N_26256,N_22741);
nor U31674 (N_31674,N_23369,N_23111);
nand U31675 (N_31675,N_21986,N_29802);
nor U31676 (N_31676,N_20800,N_27420);
or U31677 (N_31677,N_20294,N_26949);
and U31678 (N_31678,N_23842,N_23405);
xnor U31679 (N_31679,N_27422,N_27606);
or U31680 (N_31680,N_26450,N_20747);
or U31681 (N_31681,N_27032,N_22434);
xnor U31682 (N_31682,N_29574,N_20044);
or U31683 (N_31683,N_26984,N_27884);
nand U31684 (N_31684,N_20495,N_24038);
nor U31685 (N_31685,N_20305,N_28521);
nand U31686 (N_31686,N_26343,N_25626);
and U31687 (N_31687,N_23940,N_25071);
or U31688 (N_31688,N_21257,N_25070);
or U31689 (N_31689,N_24306,N_29838);
nand U31690 (N_31690,N_24436,N_21439);
or U31691 (N_31691,N_25382,N_22064);
nand U31692 (N_31692,N_24835,N_22750);
and U31693 (N_31693,N_26253,N_20076);
and U31694 (N_31694,N_28745,N_23586);
nor U31695 (N_31695,N_26273,N_25309);
xnor U31696 (N_31696,N_28921,N_24295);
xor U31697 (N_31697,N_23918,N_27365);
and U31698 (N_31698,N_27361,N_24679);
and U31699 (N_31699,N_21229,N_23587);
nor U31700 (N_31700,N_29299,N_28096);
or U31701 (N_31701,N_25947,N_29737);
nand U31702 (N_31702,N_26716,N_25498);
nand U31703 (N_31703,N_29744,N_21897);
nand U31704 (N_31704,N_24090,N_24688);
nor U31705 (N_31705,N_29402,N_20412);
and U31706 (N_31706,N_27633,N_25701);
xor U31707 (N_31707,N_28384,N_20506);
nand U31708 (N_31708,N_27657,N_29677);
nand U31709 (N_31709,N_23056,N_29954);
xnor U31710 (N_31710,N_24533,N_20302);
nand U31711 (N_31711,N_27782,N_28477);
xor U31712 (N_31712,N_29459,N_20788);
nand U31713 (N_31713,N_24105,N_29683);
xor U31714 (N_31714,N_24847,N_22234);
nand U31715 (N_31715,N_28725,N_20241);
xor U31716 (N_31716,N_28872,N_25411);
nor U31717 (N_31717,N_24426,N_23048);
and U31718 (N_31718,N_29852,N_24019);
or U31719 (N_31719,N_20479,N_29377);
xor U31720 (N_31720,N_28767,N_23982);
xor U31721 (N_31721,N_26503,N_28697);
nor U31722 (N_31722,N_26444,N_26932);
nand U31723 (N_31723,N_22393,N_23286);
and U31724 (N_31724,N_26096,N_23071);
nand U31725 (N_31725,N_26661,N_27869);
and U31726 (N_31726,N_25888,N_25661);
or U31727 (N_31727,N_26720,N_26196);
nor U31728 (N_31728,N_27787,N_28792);
nand U31729 (N_31729,N_21380,N_25980);
nor U31730 (N_31730,N_23663,N_28375);
nor U31731 (N_31731,N_20400,N_24249);
nand U31732 (N_31732,N_27253,N_21158);
nor U31733 (N_31733,N_22043,N_22572);
nor U31734 (N_31734,N_26152,N_24925);
nand U31735 (N_31735,N_23234,N_27110);
nand U31736 (N_31736,N_25855,N_28626);
nand U31737 (N_31737,N_20324,N_21045);
nor U31738 (N_31738,N_24697,N_29271);
and U31739 (N_31739,N_27118,N_21376);
xnor U31740 (N_31740,N_21863,N_29310);
nand U31741 (N_31741,N_29525,N_25312);
xnor U31742 (N_31742,N_25526,N_23695);
xnor U31743 (N_31743,N_24035,N_24570);
nor U31744 (N_31744,N_21553,N_26261);
or U31745 (N_31745,N_20748,N_28024);
and U31746 (N_31746,N_28377,N_20825);
nand U31747 (N_31747,N_25987,N_21641);
xnor U31748 (N_31748,N_29210,N_25212);
nand U31749 (N_31749,N_21188,N_20315);
nor U31750 (N_31750,N_28970,N_26187);
and U31751 (N_31751,N_29203,N_27543);
and U31752 (N_31752,N_29429,N_25476);
nand U31753 (N_31753,N_20551,N_25419);
nand U31754 (N_31754,N_24290,N_22655);
and U31755 (N_31755,N_26181,N_23285);
and U31756 (N_31756,N_24179,N_29740);
xnor U31757 (N_31757,N_29599,N_28823);
nor U31758 (N_31758,N_22977,N_24978);
xnor U31759 (N_31759,N_21155,N_23229);
nor U31760 (N_31760,N_24070,N_29978);
nand U31761 (N_31761,N_27650,N_26297);
nand U31762 (N_31762,N_26972,N_28746);
xor U31763 (N_31763,N_25136,N_27259);
nor U31764 (N_31764,N_28414,N_29576);
nand U31765 (N_31765,N_27483,N_25032);
or U31766 (N_31766,N_24322,N_28050);
nor U31767 (N_31767,N_22103,N_26565);
nand U31768 (N_31768,N_25806,N_23636);
nand U31769 (N_31769,N_23480,N_29598);
xor U31770 (N_31770,N_24308,N_25656);
and U31771 (N_31771,N_28718,N_22394);
xnor U31772 (N_31772,N_28090,N_28184);
xor U31773 (N_31773,N_26743,N_20323);
xnor U31774 (N_31774,N_23088,N_22672);
or U31775 (N_31775,N_24099,N_22425);
or U31776 (N_31776,N_20129,N_26613);
xnor U31777 (N_31777,N_26689,N_29595);
nor U31778 (N_31778,N_24682,N_24837);
or U31779 (N_31779,N_24914,N_28016);
or U31780 (N_31780,N_28379,N_23275);
or U31781 (N_31781,N_29762,N_29752);
nand U31782 (N_31782,N_22297,N_21922);
xor U31783 (N_31783,N_25077,N_28687);
or U31784 (N_31784,N_29368,N_28904);
nor U31785 (N_31785,N_22908,N_28287);
and U31786 (N_31786,N_25109,N_28420);
nor U31787 (N_31787,N_28294,N_24843);
and U31788 (N_31788,N_25082,N_20664);
nor U31789 (N_31789,N_21275,N_23689);
xor U31790 (N_31790,N_27921,N_28446);
and U31791 (N_31791,N_29872,N_23144);
or U31792 (N_31792,N_27069,N_22658);
nor U31793 (N_31793,N_23556,N_23565);
and U31794 (N_31794,N_24788,N_21416);
xnor U31795 (N_31795,N_23974,N_21325);
nand U31796 (N_31796,N_21476,N_24025);
nand U31797 (N_31797,N_25895,N_23331);
or U31798 (N_31798,N_28082,N_26580);
nand U31799 (N_31799,N_27630,N_27510);
or U31800 (N_31800,N_21441,N_28714);
nor U31801 (N_31801,N_29135,N_27283);
nor U31802 (N_31802,N_24509,N_25532);
nor U31803 (N_31803,N_24676,N_25577);
and U31804 (N_31804,N_28975,N_23245);
nor U31805 (N_31805,N_23837,N_24333);
nand U31806 (N_31806,N_21420,N_29703);
and U31807 (N_31807,N_24875,N_20308);
nor U31808 (N_31808,N_20128,N_20030);
or U31809 (N_31809,N_21343,N_28598);
and U31810 (N_31810,N_23843,N_29317);
and U31811 (N_31811,N_26070,N_21093);
xnor U31812 (N_31812,N_26479,N_29909);
and U31813 (N_31813,N_24739,N_26494);
and U31814 (N_31814,N_20074,N_27074);
nor U31815 (N_31815,N_21173,N_25336);
xor U31816 (N_31816,N_29069,N_29261);
nand U31817 (N_31817,N_26499,N_29060);
nand U31818 (N_31818,N_26164,N_25934);
nor U31819 (N_31819,N_21747,N_29503);
or U31820 (N_31820,N_28519,N_25801);
or U31821 (N_31821,N_25183,N_21886);
xor U31822 (N_31822,N_25118,N_26850);
and U31823 (N_31823,N_27799,N_26858);
or U31824 (N_31824,N_28134,N_29709);
nand U31825 (N_31825,N_20009,N_26787);
or U31826 (N_31826,N_24787,N_29537);
nand U31827 (N_31827,N_23126,N_20891);
or U31828 (N_31828,N_24859,N_24830);
xnor U31829 (N_31829,N_24957,N_28812);
or U31830 (N_31830,N_26604,N_20674);
xnor U31831 (N_31831,N_22486,N_25046);
nand U31832 (N_31832,N_28029,N_27423);
xnor U31833 (N_31833,N_21287,N_23723);
nor U31834 (N_31834,N_22969,N_24114);
or U31835 (N_31835,N_29454,N_22290);
nand U31836 (N_31836,N_24691,N_29652);
xnor U31837 (N_31837,N_23145,N_23338);
nor U31838 (N_31838,N_25758,N_23408);
xnor U31839 (N_31839,N_23811,N_27062);
xnor U31840 (N_31840,N_25973,N_29746);
nor U31841 (N_31841,N_27369,N_26352);
and U31842 (N_31842,N_28772,N_29730);
and U31843 (N_31843,N_23826,N_24857);
nand U31844 (N_31844,N_22674,N_24416);
and U31845 (N_31845,N_22584,N_25324);
and U31846 (N_31846,N_29207,N_29238);
or U31847 (N_31847,N_29635,N_23359);
nor U31848 (N_31848,N_27528,N_29326);
and U31849 (N_31849,N_23968,N_20672);
nor U31850 (N_31850,N_26081,N_28775);
nand U31851 (N_31851,N_26330,N_28635);
xor U31852 (N_31852,N_24479,N_28028);
xor U31853 (N_31853,N_25130,N_20361);
nor U31854 (N_31854,N_20714,N_24102);
nor U31855 (N_31855,N_23139,N_28683);
nor U31856 (N_31856,N_27761,N_20532);
nor U31857 (N_31857,N_22666,N_22076);
or U31858 (N_31858,N_20199,N_24761);
nor U31859 (N_31859,N_27767,N_28756);
nand U31860 (N_31860,N_24468,N_27297);
and U31861 (N_31861,N_28279,N_23778);
nand U31862 (N_31862,N_22435,N_21198);
nor U31863 (N_31863,N_25462,N_23604);
nor U31864 (N_31864,N_24406,N_26623);
and U31865 (N_31865,N_27453,N_24893);
nor U31866 (N_31866,N_23588,N_21140);
and U31867 (N_31867,N_29725,N_23688);
or U31868 (N_31868,N_26171,N_20276);
or U31869 (N_31869,N_28719,N_23988);
xnor U31870 (N_31870,N_24051,N_25148);
xor U31871 (N_31871,N_29095,N_29175);
nand U31872 (N_31872,N_23886,N_23060);
xor U31873 (N_31873,N_28851,N_24855);
nand U31874 (N_31874,N_25377,N_22622);
or U31875 (N_31875,N_28117,N_24834);
nand U31876 (N_31876,N_27627,N_22589);
and U31877 (N_31877,N_20198,N_22212);
and U31878 (N_31878,N_24275,N_25180);
nand U31879 (N_31879,N_21600,N_22630);
nor U31880 (N_31880,N_25204,N_21945);
and U31881 (N_31881,N_23993,N_25235);
xnor U31882 (N_31882,N_26002,N_28884);
and U31883 (N_31883,N_22045,N_21611);
nor U31884 (N_31884,N_22792,N_24154);
or U31885 (N_31885,N_22637,N_25239);
nor U31886 (N_31886,N_21236,N_23010);
or U31887 (N_31887,N_22912,N_24463);
xnor U31888 (N_31888,N_21143,N_21966);
nor U31889 (N_31889,N_26599,N_22699);
nor U31890 (N_31890,N_29053,N_25253);
nor U31891 (N_31891,N_25404,N_24755);
and U31892 (N_31892,N_27101,N_23927);
nand U31893 (N_31893,N_24458,N_27290);
and U31894 (N_31894,N_22756,N_29194);
and U31895 (N_31895,N_28691,N_20730);
and U31896 (N_31896,N_21289,N_28534);
nand U31897 (N_31897,N_28960,N_20626);
nand U31898 (N_31898,N_22732,N_26840);
or U31899 (N_31899,N_26856,N_26919);
xnor U31900 (N_31900,N_27385,N_27196);
and U31901 (N_31901,N_22455,N_26561);
or U31902 (N_31902,N_26607,N_21754);
nor U31903 (N_31903,N_25342,N_21241);
xnor U31904 (N_31904,N_22820,N_20708);
nor U31905 (N_31905,N_25783,N_28152);
and U31906 (N_31906,N_25170,N_26475);
xor U31907 (N_31907,N_24408,N_29510);
xor U31908 (N_31908,N_22649,N_25627);
and U31909 (N_31909,N_21007,N_23703);
nand U31910 (N_31910,N_24975,N_29523);
and U31911 (N_31911,N_26369,N_29281);
xnor U31912 (N_31912,N_21860,N_25395);
nor U31913 (N_31913,N_20833,N_27909);
nor U31914 (N_31914,N_27607,N_29182);
xor U31915 (N_31915,N_21246,N_24966);
nand U31916 (N_31916,N_24218,N_22291);
and U31917 (N_31917,N_24779,N_29159);
xor U31918 (N_31918,N_27758,N_28085);
and U31919 (N_31919,N_26375,N_24653);
xnor U31920 (N_31920,N_27720,N_26639);
xnor U31921 (N_31921,N_25173,N_29831);
or U31922 (N_31922,N_23385,N_21545);
and U31923 (N_31923,N_25761,N_20160);
xnor U31924 (N_31924,N_28986,N_22197);
or U31925 (N_31925,N_29759,N_24998);
or U31926 (N_31926,N_20648,N_24699);
or U31927 (N_31927,N_22981,N_20831);
or U31928 (N_31928,N_24864,N_20972);
xnor U31929 (N_31929,N_28636,N_27994);
nor U31930 (N_31930,N_23752,N_23671);
xnor U31931 (N_31931,N_25076,N_24758);
nand U31932 (N_31932,N_21258,N_26184);
xnor U31933 (N_31933,N_27279,N_22682);
or U31934 (N_31934,N_21643,N_23136);
xor U31935 (N_31935,N_27381,N_21051);
and U31936 (N_31936,N_24594,N_29931);
and U31937 (N_31937,N_27222,N_23220);
xor U31938 (N_31938,N_27037,N_22305);
nor U31939 (N_31939,N_26857,N_22033);
nor U31940 (N_31940,N_26302,N_29518);
nor U31941 (N_31941,N_22747,N_29443);
and U31942 (N_31942,N_29342,N_28010);
or U31943 (N_31943,N_21252,N_22259);
nand U31944 (N_31944,N_25116,N_23851);
nor U31945 (N_31945,N_20456,N_29495);
and U31946 (N_31946,N_27019,N_24453);
and U31947 (N_31947,N_20112,N_20283);
and U31948 (N_31948,N_23822,N_25355);
or U31949 (N_31949,N_26529,N_29817);
or U31950 (N_31950,N_23283,N_21558);
or U31951 (N_31951,N_21107,N_27267);
and U31952 (N_31952,N_24421,N_21483);
nand U31953 (N_31953,N_22967,N_21081);
nor U31954 (N_31954,N_22422,N_20866);
nor U31955 (N_31955,N_27957,N_29585);
xnor U31956 (N_31956,N_22942,N_25242);
nor U31957 (N_31957,N_29449,N_21130);
xor U31958 (N_31958,N_24432,N_29219);
nand U31959 (N_31959,N_27120,N_25878);
and U31960 (N_31960,N_22374,N_21482);
xnor U31961 (N_31961,N_20230,N_25991);
xnor U31962 (N_31962,N_27689,N_23991);
and U31963 (N_31963,N_22055,N_23546);
xnor U31964 (N_31964,N_24129,N_28768);
and U31965 (N_31965,N_26868,N_28755);
xnor U31966 (N_31966,N_23781,N_22013);
nor U31967 (N_31967,N_28999,N_21682);
and U31968 (N_31968,N_27976,N_26095);
and U31969 (N_31969,N_22568,N_23605);
and U31970 (N_31970,N_25963,N_21399);
nand U31971 (N_31971,N_24690,N_29163);
and U31972 (N_31972,N_28732,N_21455);
nand U31973 (N_31973,N_26041,N_28545);
and U31974 (N_31974,N_27495,N_21083);
nand U31975 (N_31975,N_26557,N_29439);
and U31976 (N_31976,N_22793,N_28760);
and U31977 (N_31977,N_26508,N_23361);
and U31978 (N_31978,N_22680,N_26572);
and U31979 (N_31979,N_27659,N_29915);
and U31980 (N_31980,N_22321,N_29572);
nor U31981 (N_31981,N_20268,N_29484);
nand U31982 (N_31982,N_23932,N_23613);
and U31983 (N_31983,N_23468,N_28383);
nand U31984 (N_31984,N_29168,N_22412);
or U31985 (N_31985,N_26032,N_24815);
nor U31986 (N_31986,N_24607,N_20134);
nor U31987 (N_31987,N_21899,N_20925);
nor U31988 (N_31988,N_24207,N_27084);
nor U31989 (N_31989,N_24729,N_25340);
and U31990 (N_31990,N_20605,N_21879);
xnor U31991 (N_31991,N_20120,N_21653);
nand U31992 (N_31992,N_26220,N_27906);
nand U31993 (N_31993,N_28831,N_20712);
and U31994 (N_31994,N_24381,N_24498);
nor U31995 (N_31995,N_27450,N_29005);
and U31996 (N_31996,N_28694,N_26040);
or U31997 (N_31997,N_23847,N_22198);
and U31998 (N_31998,N_24989,N_22419);
and U31999 (N_31999,N_29461,N_22567);
and U32000 (N_32000,N_29764,N_26418);
nand U32001 (N_32001,N_27036,N_25258);
nand U32002 (N_32002,N_24031,N_28461);
xor U32003 (N_32003,N_27171,N_26621);
or U32004 (N_32004,N_29016,N_26327);
xnor U32005 (N_32005,N_23320,N_22995);
nand U32006 (N_32006,N_22248,N_22049);
xor U32007 (N_32007,N_26120,N_24848);
and U32008 (N_32008,N_29874,N_24152);
nor U32009 (N_32009,N_26264,N_26866);
or U32010 (N_32010,N_24328,N_29278);
nand U32011 (N_32011,N_23931,N_22105);
and U32012 (N_32012,N_27416,N_27741);
xor U32013 (N_32013,N_29796,N_21018);
xor U32014 (N_32014,N_24819,N_24054);
nand U32015 (N_32015,N_22342,N_27207);
or U32016 (N_32016,N_25557,N_21569);
and U32017 (N_32017,N_25503,N_21648);
nand U32018 (N_32018,N_29741,N_22007);
or U32019 (N_32019,N_27975,N_20211);
nor U32020 (N_32020,N_24390,N_26574);
nand U32021 (N_32021,N_25611,N_20620);
nor U32022 (N_32022,N_20566,N_25102);
and U32023 (N_32023,N_26734,N_20470);
nand U32024 (N_32024,N_23740,N_24565);
nand U32025 (N_32025,N_27791,N_29577);
xnor U32026 (N_32026,N_23462,N_20106);
or U32027 (N_32027,N_20187,N_21605);
xnor U32028 (N_32028,N_29821,N_28053);
or U32029 (N_32029,N_21365,N_27409);
and U32030 (N_32030,N_27154,N_23824);
nor U32031 (N_32031,N_25126,N_24948);
or U32032 (N_32032,N_27040,N_25790);
nor U32033 (N_32033,N_25575,N_22518);
or U32034 (N_32034,N_22997,N_21776);
nand U32035 (N_32035,N_26638,N_25237);
nand U32036 (N_32036,N_23755,N_20430);
and U32037 (N_32037,N_21096,N_23547);
or U32038 (N_32038,N_29663,N_20802);
nor U32039 (N_32039,N_22631,N_27224);
nand U32040 (N_32040,N_26109,N_22299);
nor U32041 (N_32041,N_26012,N_27668);
xor U32042 (N_32042,N_28633,N_26828);
nand U32043 (N_32043,N_24614,N_25820);
or U32044 (N_32044,N_26404,N_24795);
or U32045 (N_32045,N_28170,N_28418);
or U32046 (N_32046,N_20466,N_26004);
and U32047 (N_32047,N_21954,N_23363);
xor U32048 (N_32048,N_25842,N_27797);
and U32049 (N_32049,N_20716,N_24228);
xnor U32050 (N_32050,N_23643,N_22443);
and U32051 (N_32051,N_21286,N_21590);
nor U32052 (N_32052,N_26578,N_25066);
nor U32053 (N_32053,N_22099,N_26435);
nand U32054 (N_32054,N_22547,N_23435);
xnor U32055 (N_32055,N_22140,N_24882);
and U32056 (N_32056,N_22272,N_22224);
or U32057 (N_32057,N_23280,N_25203);
xnor U32058 (N_32058,N_29217,N_27725);
or U32059 (N_32059,N_20701,N_26523);
nand U32060 (N_32060,N_23185,N_21758);
and U32061 (N_32061,N_29997,N_29735);
xor U32062 (N_32062,N_29132,N_29551);
nor U32063 (N_32063,N_22911,N_22185);
nor U32064 (N_32064,N_28220,N_22400);
xor U32065 (N_32065,N_21620,N_26480);
nor U32066 (N_32066,N_26669,N_23156);
nor U32067 (N_32067,N_24744,N_22876);
xor U32068 (N_32068,N_29571,N_25652);
xor U32069 (N_32069,N_23721,N_25599);
nand U32070 (N_32070,N_22123,N_24314);
nor U32071 (N_32071,N_22039,N_27410);
xor U32072 (N_32072,N_25893,N_28370);
and U32073 (N_32073,N_24774,N_25400);
nand U32074 (N_32074,N_20426,N_22453);
xnor U32075 (N_32075,N_20051,N_21298);
nand U32076 (N_32076,N_27478,N_27898);
and U32077 (N_32077,N_26951,N_26306);
nor U32078 (N_32078,N_20544,N_25879);
nand U32079 (N_32079,N_23642,N_22333);
nand U32080 (N_32080,N_26179,N_29690);
nor U32081 (N_32081,N_23726,N_26630);
and U32082 (N_32082,N_25198,N_25072);
nor U32083 (N_32083,N_29081,N_20392);
xor U32084 (N_32084,N_24304,N_29937);
xor U32085 (N_32085,N_28989,N_26281);
nand U32086 (N_32086,N_29887,N_22960);
xor U32087 (N_32087,N_27144,N_27208);
nand U32088 (N_32088,N_24554,N_20746);
nor U32089 (N_32089,N_27443,N_20011);
nor U32090 (N_32090,N_21562,N_28988);
and U32091 (N_32091,N_26010,N_20614);
nor U32092 (N_32092,N_20423,N_24444);
or U32093 (N_32093,N_20688,N_22965);
nor U32094 (N_32094,N_29506,N_22996);
and U32095 (N_32095,N_21624,N_28811);
or U32096 (N_32096,N_26990,N_25399);
or U32097 (N_32097,N_28623,N_22302);
nor U32098 (N_32098,N_29237,N_23704);
nand U32099 (N_32099,N_28326,N_23610);
nor U32100 (N_32100,N_28517,N_27679);
nand U32101 (N_32101,N_21392,N_21253);
xor U32102 (N_32102,N_22634,N_28259);
or U32103 (N_32103,N_27235,N_22657);
or U32104 (N_32104,N_27551,N_21814);
and U32105 (N_32105,N_21121,N_24451);
nor U32106 (N_32106,N_29111,N_21330);
xor U32107 (N_32107,N_26274,N_24014);
nand U32108 (N_32108,N_20529,N_28655);
xnor U32109 (N_32109,N_25057,N_21645);
or U32110 (N_32110,N_24684,N_25731);
and U32111 (N_32111,N_20892,N_22999);
nor U32112 (N_32112,N_27707,N_20179);
nor U32113 (N_32113,N_27275,N_25326);
or U32114 (N_32114,N_23214,N_27183);
and U32115 (N_32115,N_26570,N_25845);
and U32116 (N_32116,N_24908,N_28332);
nand U32117 (N_32117,N_28341,N_27321);
nand U32118 (N_32118,N_28619,N_27472);
or U32119 (N_32119,N_29304,N_26808);
nor U32120 (N_32120,N_29573,N_25648);
nor U32121 (N_32121,N_22509,N_20100);
nor U32122 (N_32122,N_26704,N_28740);
xor U32123 (N_32123,N_28994,N_23221);
nand U32124 (N_32124,N_24055,N_23627);
or U32125 (N_32125,N_27227,N_26871);
nand U32126 (N_32126,N_23646,N_20154);
nand U32127 (N_32127,N_23316,N_22724);
and U32128 (N_32128,N_24374,N_21996);
xnor U32129 (N_32129,N_29408,N_21673);
nor U32130 (N_32130,N_26385,N_29568);
or U32131 (N_32131,N_27700,N_29883);
nand U32132 (N_32132,N_23622,N_23925);
xnor U32133 (N_32133,N_26861,N_26467);
nand U32134 (N_32134,N_23517,N_21715);
xnor U32135 (N_32135,N_22442,N_24648);
or U32136 (N_32136,N_28034,N_27838);
xor U32137 (N_32137,N_20369,N_29096);
nand U32138 (N_32138,N_23624,N_25363);
nand U32139 (N_32139,N_26053,N_29106);
and U32140 (N_32140,N_27477,N_28634);
or U32141 (N_32141,N_24534,N_27002);
nor U32142 (N_32142,N_29619,N_25105);
nor U32143 (N_32143,N_25484,N_20472);
xor U32144 (N_32144,N_20865,N_22244);
xnor U32145 (N_32145,N_22228,N_24748);
nand U32146 (N_32146,N_21249,N_20101);
nor U32147 (N_32147,N_22226,N_20103);
or U32148 (N_32148,N_28410,N_24630);
nor U32149 (N_32149,N_25098,N_26929);
and U32150 (N_32150,N_26822,N_29149);
nand U32151 (N_32151,N_26186,N_21505);
or U32152 (N_32152,N_29707,N_26518);
or U32153 (N_32153,N_20500,N_25317);
xnor U32154 (N_32154,N_26703,N_28068);
or U32155 (N_32155,N_23852,N_21488);
xor U32156 (N_32156,N_23154,N_23678);
and U32157 (N_32157,N_27590,N_21661);
xnor U32158 (N_32158,N_22844,N_23342);
or U32159 (N_32159,N_21570,N_25238);
or U32160 (N_32160,N_21937,N_26573);
xor U32161 (N_32161,N_22163,N_27296);
nand U32162 (N_32162,N_21835,N_20286);
or U32163 (N_32163,N_29609,N_29124);
nor U32164 (N_32164,N_21763,N_29877);
and U32165 (N_32165,N_29526,N_26894);
or U32166 (N_32166,N_23512,N_28398);
or U32167 (N_32167,N_20173,N_28833);
nor U32168 (N_32168,N_27615,N_22852);
xor U32169 (N_32169,N_21288,N_22382);
nor U32170 (N_32170,N_23270,N_24517);
and U32171 (N_32171,N_26288,N_23121);
or U32172 (N_32172,N_29770,N_23343);
nand U32173 (N_32173,N_28847,N_28950);
nand U32174 (N_32174,N_25292,N_22015);
nor U32175 (N_32175,N_22356,N_28472);
xnor U32176 (N_32176,N_28168,N_25965);
or U32177 (N_32177,N_26773,N_25615);
nand U32178 (N_32178,N_29251,N_29671);
nor U32179 (N_32179,N_24877,N_24715);
nor U32180 (N_32180,N_23272,N_28880);
and U32181 (N_32181,N_24247,N_21846);
or U32182 (N_32182,N_28438,N_20158);
nand U32183 (N_32183,N_20634,N_26455);
nor U32184 (N_32184,N_20596,N_26895);
nor U32185 (N_32185,N_27780,N_25700);
xnor U32186 (N_32186,N_21443,N_22517);
nand U32187 (N_32187,N_22790,N_25273);
xnor U32188 (N_32188,N_28791,N_23807);
xor U32189 (N_32189,N_20042,N_23948);
nand U32190 (N_32190,N_20061,N_26431);
nor U32191 (N_32191,N_20951,N_25787);
nand U32192 (N_32192,N_24201,N_23835);
or U32193 (N_32193,N_22998,N_23521);
nand U32194 (N_32194,N_25458,N_22091);
nor U32195 (N_32195,N_25314,N_21424);
xnor U32196 (N_32196,N_28639,N_24820);
and U32197 (N_32197,N_22088,N_24606);
xnor U32198 (N_32198,N_25606,N_28870);
nand U32199 (N_32199,N_26810,N_24511);
xor U32200 (N_32200,N_21267,N_22870);
and U32201 (N_32201,N_20929,N_22261);
nand U32202 (N_32202,N_21510,N_20795);
and U32203 (N_32203,N_29162,N_22494);
nand U32204 (N_32204,N_29777,N_26452);
nand U32205 (N_32205,N_28158,N_29832);
nand U32206 (N_32206,N_20417,N_21979);
nand U32207 (N_32207,N_28478,N_27119);
or U32208 (N_32208,N_28352,N_29148);
and U32209 (N_32209,N_23580,N_24940);
nand U32210 (N_32210,N_22352,N_23090);
nand U32211 (N_32211,N_23073,N_24427);
and U32212 (N_32212,N_22799,N_20981);
xnor U32213 (N_32213,N_25560,N_27112);
nand U32214 (N_32214,N_28933,N_25918);
xnor U32215 (N_32215,N_27100,N_27878);
nand U32216 (N_32216,N_26668,N_22069);
xnor U32217 (N_32217,N_25455,N_27736);
or U32218 (N_32218,N_23554,N_24958);
and U32219 (N_32219,N_28244,N_21980);
nand U32220 (N_32220,N_25644,N_28763);
and U32221 (N_32221,N_26493,N_24246);
and U32222 (N_32222,N_20565,N_26318);
and U32223 (N_32223,N_29355,N_26000);
and U32224 (N_32224,N_22980,N_25186);
or U32225 (N_32225,N_22280,N_25491);
or U32226 (N_32226,N_29617,N_29830);
xnor U32227 (N_32227,N_28074,N_29825);
or U32228 (N_32228,N_28563,N_29197);
and U32229 (N_32229,N_27739,N_22638);
xor U32230 (N_32230,N_22264,N_22835);
xor U32231 (N_32231,N_22262,N_28990);
or U32232 (N_32232,N_22166,N_23694);
nor U32233 (N_32233,N_28365,N_26569);
nand U32234 (N_32234,N_23341,N_24718);
nor U32235 (N_32235,N_24434,N_27318);
or U32236 (N_32236,N_29212,N_28612);
nor U32237 (N_32237,N_27777,N_25360);
and U32238 (N_32238,N_24184,N_22875);
nand U32239 (N_32239,N_25015,N_29511);
nand U32240 (N_32240,N_22520,N_22830);
xnor U32241 (N_32241,N_20243,N_26727);
nor U32242 (N_32242,N_22683,N_23939);
and U32243 (N_32243,N_25817,N_29667);
nand U32244 (N_32244,N_26236,N_27236);
nand U32245 (N_32245,N_27526,N_20598);
xnor U32246 (N_32246,N_27701,N_27498);
xnor U32247 (N_32247,N_25694,N_20442);
or U32248 (N_32248,N_28052,N_25868);
xor U32249 (N_32249,N_28181,N_23186);
and U32250 (N_32250,N_21970,N_21614);
nand U32251 (N_32251,N_28501,N_27827);
nand U32252 (N_32252,N_23664,N_21208);
nor U32253 (N_32253,N_23349,N_28495);
and U32254 (N_32254,N_21118,N_22952);
nor U32255 (N_32255,N_26016,N_20132);
xor U32256 (N_32256,N_26128,N_23953);
or U32257 (N_32257,N_22760,N_21659);
xor U32258 (N_32258,N_20093,N_22846);
nor U32259 (N_32259,N_22676,N_22841);
and U32260 (N_32260,N_20409,N_29775);
nand U32261 (N_32261,N_28700,N_24009);
nand U32262 (N_32262,N_26278,N_29726);
nand U32263 (N_32263,N_23880,N_26166);
xnor U32264 (N_32264,N_29991,N_22644);
nand U32265 (N_32265,N_25630,N_20709);
and U32266 (N_32266,N_25268,N_26881);
nor U32267 (N_32267,N_21679,N_22293);
or U32268 (N_32268,N_20717,N_23560);
nor U32269 (N_32269,N_28032,N_26538);
xnor U32270 (N_32270,N_22277,N_29479);
nand U32271 (N_32271,N_20948,N_29961);
nor U32272 (N_32272,N_28651,N_26121);
nor U32273 (N_32273,N_23196,N_26148);
nor U32274 (N_32274,N_20898,N_24404);
nor U32275 (N_32275,N_22675,N_26005);
or U32276 (N_32276,N_20640,N_26232);
nand U32277 (N_32277,N_26860,N_27128);
or U32278 (N_32278,N_22929,N_20787);
nor U32279 (N_32279,N_29353,N_24799);
and U32280 (N_32280,N_23318,N_21192);
xor U32281 (N_32281,N_20786,N_26445);
and U32282 (N_32282,N_28381,N_26560);
xnor U32283 (N_32283,N_21405,N_20754);
nor U32284 (N_32284,N_27717,N_23656);
nor U32285 (N_32285,N_25391,N_23207);
nor U32286 (N_32286,N_25350,N_23157);
xnor U32287 (N_32287,N_26581,N_27067);
or U32288 (N_32288,N_25356,N_20779);
nand U32289 (N_32289,N_23269,N_20021);
or U32290 (N_32290,N_21760,N_29199);
or U32291 (N_32291,N_24987,N_23476);
or U32292 (N_32292,N_21528,N_29720);
or U32293 (N_32293,N_29004,N_22577);
nor U32294 (N_32294,N_21161,N_22138);
xor U32295 (N_32295,N_21712,N_29090);
nand U32296 (N_32296,N_25134,N_23328);
or U32297 (N_32297,N_29405,N_26305);
nand U32298 (N_32298,N_26516,N_22036);
or U32299 (N_32299,N_25926,N_24351);
nand U32300 (N_32300,N_28448,N_21869);
nand U32301 (N_32301,N_28947,N_29059);
nor U32302 (N_32302,N_22231,N_24293);
and U32303 (N_32303,N_29323,N_21830);
and U32304 (N_32304,N_22008,N_23845);
xnor U32305 (N_32305,N_27449,N_27885);
and U32306 (N_32306,N_28435,N_29815);
nor U32307 (N_32307,N_26425,N_29955);
xor U32308 (N_32308,N_22943,N_25971);
nor U32309 (N_32309,N_25414,N_21973);
xnor U32310 (N_32310,N_26110,N_23952);
nand U32311 (N_32311,N_23728,N_28974);
nand U32312 (N_32312,N_23564,N_29248);
nand U32313 (N_32313,N_24098,N_23043);
and U32314 (N_32314,N_25343,N_26656);
nor U32315 (N_32315,N_25236,N_23401);
or U32316 (N_32316,N_25165,N_26215);
xnor U32317 (N_32317,N_26300,N_23732);
nand U32318 (N_32318,N_22685,N_29434);
nor U32319 (N_32319,N_28285,N_22137);
and U32320 (N_32320,N_28084,N_23693);
or U32321 (N_32321,N_29869,N_26268);
xnor U32322 (N_32322,N_20048,N_23861);
nand U32323 (N_32323,N_27757,N_23981);
and U32324 (N_32324,N_22210,N_28298);
or U32325 (N_32325,N_29559,N_23277);
nor U32326 (N_32326,N_27173,N_25137);
or U32327 (N_32327,N_28513,N_22669);
nand U32328 (N_32328,N_25759,N_22249);
xnor U32329 (N_32329,N_20164,N_25982);
or U32330 (N_32330,N_24777,N_28144);
nand U32331 (N_32331,N_24520,N_22024);
xnor U32332 (N_32332,N_25663,N_23499);
nor U32333 (N_32333,N_25364,N_20471);
or U32334 (N_32334,N_21122,N_28903);
nand U32335 (N_32335,N_26321,N_26339);
nand U32336 (N_32336,N_28538,N_29567);
and U32337 (N_32337,N_20773,N_25828);
or U32338 (N_32338,N_26449,N_22396);
or U32339 (N_32339,N_27809,N_20919);
or U32340 (N_32340,N_29622,N_25546);
xnor U32341 (N_32341,N_27941,N_29457);
nor U32342 (N_32342,N_28839,N_27016);
xor U32343 (N_32343,N_27461,N_24923);
xor U32344 (N_32344,N_23148,N_24252);
xor U32345 (N_32345,N_26601,N_27571);
xor U32346 (N_32346,N_28122,N_20963);
nor U32347 (N_32347,N_21972,N_24156);
nand U32348 (N_32348,N_20410,N_25193);
or U32349 (N_32349,N_20060,N_21128);
and U32350 (N_32350,N_21546,N_22639);
nand U32351 (N_32351,N_24713,N_27596);
and U32352 (N_32352,N_28917,N_20817);
nor U32353 (N_32353,N_27273,N_29648);
or U32354 (N_32354,N_22848,N_21233);
and U32355 (N_32355,N_26119,N_26764);
and U32356 (N_32356,N_29967,N_29466);
xnor U32357 (N_32357,N_29193,N_21539);
nand U32358 (N_32358,N_28087,N_20768);
and U32359 (N_32359,N_29876,N_20188);
or U32360 (N_32360,N_25305,N_23057);
nand U32361 (N_32361,N_27581,N_23482);
xnor U32362 (N_32362,N_25728,N_20477);
nor U32363 (N_32363,N_20842,N_26021);
nor U32364 (N_32364,N_27020,N_26842);
xor U32365 (N_32365,N_24165,N_21215);
nor U32366 (N_32366,N_25909,N_25772);
nand U32367 (N_32367,N_25819,N_24805);
nor U32368 (N_32368,N_29496,N_27755);
nand U32369 (N_32369,N_29750,N_25922);
nand U32370 (N_32370,N_29471,N_20485);
nor U32371 (N_32371,N_26142,N_24398);
xor U32372 (N_32372,N_29103,N_29272);
and U32373 (N_32373,N_21518,N_27860);
and U32374 (N_32374,N_20612,N_23504);
or U32375 (N_32375,N_25531,N_23033);
nand U32376 (N_32376,N_25339,N_22081);
or U32377 (N_32377,N_24550,N_23753);
or U32378 (N_32378,N_25123,N_21309);
xor U32379 (N_32379,N_28128,N_28133);
and U32380 (N_32380,N_29771,N_25448);
or U32381 (N_32381,N_22381,N_24556);
and U32382 (N_32382,N_23458,N_21930);
xnor U32383 (N_32383,N_23125,N_27442);
nand U32384 (N_32384,N_25631,N_26316);
xnor U32385 (N_32385,N_24182,N_23872);
xor U32386 (N_32386,N_29911,N_29886);
nor U32387 (N_32387,N_23873,N_21998);
and U32388 (N_32388,N_24231,N_23396);
nand U32389 (N_32389,N_23493,N_26817);
or U32390 (N_32390,N_24663,N_26899);
xor U32391 (N_32391,N_29994,N_24963);
or U32392 (N_32392,N_26760,N_27322);
xor U32393 (N_32393,N_20351,N_28436);
or U32394 (N_32394,N_27288,N_29790);
and U32395 (N_32395,N_26382,N_24716);
and U32396 (N_32396,N_20522,N_24095);
nor U32397 (N_32397,N_20812,N_28112);
nand U32398 (N_32398,N_29101,N_29290);
nand U32399 (N_32399,N_29739,N_25289);
nand U32400 (N_32400,N_23431,N_23514);
nand U32401 (N_32401,N_25014,N_28785);
and U32402 (N_32402,N_22755,N_23312);
xnor U32403 (N_32403,N_23933,N_21297);
nor U32404 (N_32404,N_21144,N_29527);
xnor U32405 (N_32405,N_29940,N_29040);
or U32406 (N_32406,N_21230,N_21810);
xnor U32407 (N_32407,N_28759,N_20110);
and U32408 (N_32408,N_21039,N_23541);
xnor U32409 (N_32409,N_27537,N_20611);
and U32410 (N_32410,N_23082,N_21977);
xor U32411 (N_32411,N_24175,N_27958);
or U32412 (N_32412,N_27451,N_27845);
and U32413 (N_32413,N_22788,N_27382);
and U32414 (N_32414,N_27642,N_25315);
xor U32415 (N_32415,N_22695,N_28866);
nand U32416 (N_32416,N_21549,N_22256);
and U32417 (N_32417,N_27270,N_24658);
nand U32418 (N_32418,N_27214,N_22072);
and U32419 (N_32419,N_26571,N_28559);
and U32420 (N_32420,N_21265,N_24334);
and U32421 (N_32421,N_29441,N_20462);
nor U32422 (N_32422,N_25601,N_27486);
and U32423 (N_32423,N_22242,N_20213);
or U32424 (N_32424,N_23222,N_21592);
nor U32425 (N_32425,N_24776,N_20979);
nand U32426 (N_32426,N_26379,N_20415);
xnor U32427 (N_32427,N_27623,N_29453);
or U32428 (N_32428,N_25132,N_25978);
nand U32429 (N_32429,N_20291,N_20508);
nand U32430 (N_32430,N_24483,N_23634);
nand U32431 (N_32431,N_26323,N_25579);
nand U32432 (N_32432,N_27249,N_26825);
nand U32433 (N_32433,N_27419,N_27586);
or U32434 (N_32434,N_24380,N_27123);
and U32435 (N_32435,N_28549,N_28927);
or U32436 (N_32436,N_27174,N_27065);
xor U32437 (N_32437,N_25181,N_25063);
and U32438 (N_32438,N_22389,N_28867);
or U32439 (N_32439,N_22583,N_23087);
and U32440 (N_32440,N_21172,N_20359);
xnor U32441 (N_32441,N_27908,N_26517);
nor U32442 (N_32442,N_22385,N_22426);
and U32443 (N_32443,N_21464,N_28934);
nor U32444 (N_32444,N_26267,N_23409);
or U32445 (N_32445,N_28747,N_25708);
nor U32446 (N_32446,N_20000,N_25608);
or U32447 (N_32447,N_28054,N_21907);
nor U32448 (N_32448,N_23254,N_24096);
and U32449 (N_32449,N_22446,N_20444);
nor U32450 (N_32450,N_21576,N_26228);
nand U32451 (N_32451,N_28233,N_21689);
and U32452 (N_32452,N_24076,N_29659);
or U32453 (N_32453,N_25490,N_22012);
xor U32454 (N_32454,N_26033,N_24628);
or U32455 (N_32455,N_20835,N_25610);
or U32456 (N_32456,N_21100,N_29416);
nor U32457 (N_32457,N_27071,N_26645);
nor U32458 (N_32458,N_24078,N_22179);
xor U32459 (N_32459,N_25207,N_24104);
and U32460 (N_32460,N_24786,N_27392);
xnor U32461 (N_32461,N_20231,N_26192);
or U32462 (N_32462,N_22856,N_20525);
or U32463 (N_32463,N_26491,N_26907);
nor U32464 (N_32464,N_27536,N_24698);
nand U32465 (N_32465,N_27704,N_23576);
nor U32466 (N_32466,N_22945,N_20041);
nand U32467 (N_32467,N_23816,N_20693);
and U32468 (N_32468,N_27858,N_26381);
xor U32469 (N_32469,N_28523,N_29451);
nor U32470 (N_32470,N_24474,N_26362);
and U32471 (N_32471,N_25277,N_27709);
nand U32472 (N_32472,N_23527,N_21035);
and U32473 (N_32473,N_23324,N_29826);
xor U32474 (N_32474,N_22257,N_28905);
and U32475 (N_32475,N_23042,N_22354);
or U32476 (N_32476,N_28596,N_24841);
and U32477 (N_32477,N_29930,N_26075);
xor U32478 (N_32478,N_23746,N_22528);
nor U32479 (N_32479,N_22145,N_22079);
xor U32480 (N_32480,N_26168,N_20882);
xnor U32481 (N_32481,N_20654,N_28875);
xor U32482 (N_32482,N_29781,N_23795);
xor U32483 (N_32483,N_25544,N_28570);
xnor U32484 (N_32484,N_27165,N_26079);
nand U32485 (N_32485,N_20407,N_27166);
xor U32486 (N_32486,N_27628,N_27821);
or U32487 (N_32487,N_27744,N_29515);
or U32488 (N_32488,N_28782,N_21435);
xor U32489 (N_32489,N_23936,N_28541);
and U32490 (N_32490,N_29426,N_21094);
and U32491 (N_32491,N_20157,N_23006);
xnor U32492 (N_32492,N_20450,N_23382);
or U32493 (N_32493,N_27840,N_22891);
and U32494 (N_32494,N_24327,N_27053);
nor U32495 (N_32495,N_26224,N_26355);
xnor U32496 (N_32496,N_23441,N_21771);
nor U32497 (N_32497,N_26916,N_27201);
or U32498 (N_32498,N_26719,N_22575);
xor U32499 (N_32499,N_22865,N_22549);
and U32500 (N_32500,N_22909,N_23032);
xnor U32501 (N_32501,N_28825,N_26803);
and U32502 (N_32502,N_20244,N_29556);
xor U32503 (N_32503,N_22233,N_27690);
xor U32504 (N_32504,N_24064,N_24264);
xor U32505 (N_32505,N_28348,N_23983);
nor U32506 (N_32506,N_25480,N_25598);
nor U32507 (N_32507,N_20934,N_21876);
or U32508 (N_32508,N_23858,N_24489);
or U32509 (N_32509,N_20181,N_23248);
and U32510 (N_32510,N_25245,N_23708);
xor U32511 (N_32511,N_28964,N_28883);
or U32512 (N_32512,N_20125,N_22379);
nor U32513 (N_32513,N_21887,N_28871);
xnor U32514 (N_32514,N_24900,N_26979);
nand U32515 (N_32515,N_27271,N_29421);
nand U32516 (N_32516,N_28496,N_25550);
xnor U32517 (N_32517,N_28230,N_28749);
and U32518 (N_32518,N_27293,N_24965);
or U32519 (N_32519,N_25443,N_22111);
nand U32520 (N_32520,N_20229,N_28217);
nand U32521 (N_32521,N_29712,N_26286);
nand U32522 (N_32522,N_22798,N_27937);
nor U32523 (N_32523,N_23998,N_20656);
nor U32524 (N_32524,N_26260,N_27773);
or U32525 (N_32525,N_22983,N_25158);
xnor U32526 (N_32526,N_21823,N_22073);
xnor U32527 (N_32527,N_22702,N_29039);
xnor U32528 (N_32528,N_23114,N_27533);
nor U32529 (N_32529,N_21736,N_27670);
xnor U32530 (N_32530,N_23714,N_26971);
xnor U32531 (N_32531,N_25264,N_29002);
nand U32532 (N_32532,N_27372,N_22491);
xnor U32533 (N_32533,N_20194,N_29570);
and U32534 (N_32534,N_27899,N_22121);
and U32535 (N_32535,N_27193,N_26312);
xor U32536 (N_32536,N_24863,N_27691);
and U32537 (N_32537,N_28937,N_28578);
nand U32538 (N_32538,N_26045,N_24324);
nand U32539 (N_32539,N_28149,N_20438);
nand U32540 (N_32540,N_22948,N_23464);
or U32541 (N_32541,N_23447,N_29136);
nand U32542 (N_32542,N_23150,N_28325);
or U32543 (N_32543,N_26943,N_24579);
and U32544 (N_32544,N_28312,N_27177);
nor U32545 (N_32545,N_21829,N_24167);
xor U32546 (N_32546,N_23775,N_28156);
nand U32547 (N_32547,N_26315,N_23668);
or U32548 (N_32548,N_25564,N_26596);
nor U32549 (N_32549,N_28009,N_28754);
xnor U32550 (N_32550,N_28031,N_24930);
nand U32551 (N_32551,N_21034,N_21003);
nor U32552 (N_32552,N_28160,N_27579);
nor U32553 (N_32553,N_25434,N_24885);
nand U32554 (N_32554,N_20543,N_25453);
xnor U32555 (N_32555,N_23537,N_28675);
nor U32556 (N_32556,N_25521,N_28242);
or U32557 (N_32557,N_23459,N_29215);
or U32558 (N_32558,N_22071,N_20698);
and U32559 (N_32559,N_28684,N_23567);
nor U32560 (N_32560,N_27604,N_22777);
nand U32561 (N_32561,N_26117,N_22424);
xnor U32562 (N_32562,N_21024,N_23055);
nor U32563 (N_32563,N_28358,N_25901);
or U32564 (N_32564,N_26625,N_23751);
nor U32565 (N_32565,N_23218,N_22771);
and U32566 (N_32566,N_20586,N_23815);
nand U32567 (N_32567,N_20016,N_26239);
nand U32568 (N_32568,N_22083,N_25541);
nor U32569 (N_32569,N_29785,N_24766);
or U32570 (N_32570,N_25554,N_29288);
and U32571 (N_32571,N_25654,N_21174);
nand U32572 (N_32572,N_25714,N_26535);
nor U32573 (N_32573,N_24640,N_25044);
or U32574 (N_32574,N_28321,N_28434);
nor U32575 (N_32575,N_20597,N_21947);
or U32576 (N_32576,N_23085,N_27368);
or U32577 (N_32577,N_26610,N_24546);
nand U32578 (N_32578,N_23817,N_21163);
or U32579 (N_32579,N_22100,N_28226);
xnor U32580 (N_32580,N_26769,N_27089);
nand U32581 (N_32581,N_24315,N_20484);
nor U32582 (N_32582,N_20285,N_25886);
xor U32583 (N_32583,N_23079,N_26118);
xor U32584 (N_32584,N_28453,N_24997);
or U32585 (N_32585,N_23949,N_21901);
or U32586 (N_32586,N_21407,N_23690);
xor U32587 (N_32587,N_23985,N_22781);
nand U32588 (N_32588,N_22029,N_23501);
and U32589 (N_32589,N_23779,N_22211);
xnor U32590 (N_32590,N_23120,N_29500);
xnor U32591 (N_32591,N_25276,N_29082);
or U32592 (N_32592,N_26025,N_25778);
nor U32593 (N_32593,N_21370,N_25117);
or U32594 (N_32594,N_28525,N_20906);
or U32595 (N_32595,N_23015,N_25933);
nor U32596 (N_32596,N_23026,N_23986);
nor U32597 (N_32597,N_27535,N_29042);
xnor U32598 (N_32598,N_24666,N_22481);
nand U32599 (N_32599,N_26728,N_24583);
nand U32600 (N_32600,N_22762,N_23333);
nor U32601 (N_32601,N_26993,N_26207);
or U32602 (N_32602,N_20562,N_27029);
nor U32603 (N_32603,N_21526,N_26939);
xnor U32604 (N_32604,N_27194,N_20983);
xor U32605 (N_32605,N_29273,N_23224);
or U32606 (N_32606,N_26229,N_26556);
or U32607 (N_32607,N_20270,N_25641);
or U32608 (N_32608,N_24452,N_24936);
nor U32609 (N_32609,N_23420,N_25848);
or U32610 (N_32610,N_23027,N_22359);
or U32611 (N_32611,N_24052,N_22802);
and U32612 (N_32612,N_26647,N_23686);
and U32613 (N_32613,N_26982,N_26093);
and U32614 (N_32614,N_25271,N_24827);
and U32615 (N_32615,N_27356,N_24049);
nand U32616 (N_32616,N_23461,N_22961);
xor U32617 (N_32617,N_27018,N_25732);
nand U32618 (N_32618,N_26451,N_23108);
and U32619 (N_32619,N_25809,N_29956);
and U32620 (N_32620,N_27566,N_23190);
or U32621 (N_32621,N_20619,N_21609);
xor U32622 (N_32622,N_25614,N_25432);
nand U32623 (N_32623,N_29563,N_23130);
nand U32624 (N_32624,N_26739,N_26790);
xnor U32625 (N_32625,N_24988,N_21220);
and U32626 (N_32626,N_29558,N_20474);
and U32627 (N_32627,N_29130,N_20846);
nor U32628 (N_32628,N_24927,N_22001);
and U32629 (N_32629,N_28751,N_25616);
and U32630 (N_32630,N_20822,N_28153);
and U32631 (N_32631,N_20376,N_28237);
and U32632 (N_32632,N_20461,N_28490);
nor U32633 (N_32633,N_25255,N_24986);
xnor U32634 (N_32634,N_28808,N_25081);
or U32635 (N_32635,N_29893,N_22924);
xnor U32636 (N_32636,N_25734,N_29030);
nand U32637 (N_32637,N_20755,N_21989);
and U32638 (N_32638,N_29947,N_29731);
xnor U32639 (N_32639,N_24244,N_20575);
xnor U32640 (N_32640,N_20318,N_29981);
nor U32641 (N_32641,N_28587,N_21571);
or U32642 (N_32642,N_28971,N_26066);
or U32643 (N_32643,N_29587,N_20885);
or U32644 (N_32644,N_24391,N_29642);
nand U32645 (N_32645,N_22652,N_22431);
xor U32646 (N_32646,N_22107,N_21864);
and U32647 (N_32647,N_29604,N_24826);
xor U32648 (N_32648,N_23614,N_28187);
and U32649 (N_32649,N_20758,N_25119);
xor U32650 (N_32650,N_23558,N_28257);
nor U32651 (N_32651,N_26582,N_23188);
nand U32652 (N_32652,N_25417,N_28554);
and U32653 (N_32653,N_21418,N_22506);
nor U32654 (N_32654,N_28788,N_26213);
nor U32655 (N_32655,N_28166,N_23321);
or U32656 (N_32656,N_21956,N_26845);
or U32657 (N_32657,N_29851,N_27268);
or U32658 (N_32658,N_20441,N_26328);
xnor U32659 (N_32659,N_28537,N_26234);
nor U32660 (N_32660,N_21145,N_29477);
xnor U32661 (N_32661,N_21670,N_29628);
nor U32662 (N_32662,N_29719,N_25384);
nor U32663 (N_32663,N_22632,N_28066);
nor U32664 (N_32664,N_23808,N_25251);
nand U32665 (N_32665,N_22543,N_20293);
xor U32666 (N_32666,N_26644,N_24598);
nor U32667 (N_32667,N_24756,N_26047);
xor U32668 (N_32668,N_25667,N_25224);
and U32669 (N_32669,N_29068,N_25426);
nand U32670 (N_32670,N_20310,N_27354);
nand U32671 (N_32671,N_26848,N_24087);
nand U32672 (N_32672,N_26515,N_25743);
or U32673 (N_32673,N_29724,N_28588);
xor U32674 (N_32674,N_22707,N_23844);
nand U32675 (N_32675,N_28459,N_27281);
nand U32676 (N_32676,N_28076,N_26384);
nand U32677 (N_32677,N_21895,N_23973);
nor U32678 (N_32678,N_24693,N_24500);
or U32679 (N_32679,N_27560,N_24641);
nand U32680 (N_32680,N_22405,N_24750);
nor U32681 (N_32681,N_26366,N_24660);
xnor U32682 (N_32682,N_28333,N_28548);
nand U32683 (N_32683,N_29633,N_23200);
and U32684 (N_32684,N_22833,N_27920);
xnor U32685 (N_32685,N_20272,N_24959);
xor U32686 (N_32686,N_21941,N_22910);
xnor U32687 (N_32687,N_25944,N_24664);
nor U32688 (N_32688,N_21767,N_21462);
nor U32689 (N_32689,N_27028,N_23635);
and U32690 (N_32690,N_28660,N_26873);
nor U32691 (N_32691,N_24058,N_23356);
nand U32692 (N_32692,N_26751,N_24763);
nand U32693 (N_32693,N_27829,N_27133);
nand U32694 (N_32694,N_21563,N_28542);
xnor U32695 (N_32695,N_28131,N_24487);
xnor U32696 (N_32696,N_25074,N_27169);
nor U32697 (N_32697,N_24340,N_28437);
and U32698 (N_32698,N_26399,N_21280);
or U32699 (N_32699,N_23924,N_23246);
and U32700 (N_32700,N_23498,N_23566);
or U32701 (N_32701,N_21599,N_22782);
nor U32702 (N_32702,N_26056,N_21739);
and U32703 (N_32703,N_27568,N_28712);
xnor U32704 (N_32704,N_23739,N_25592);
nor U32705 (N_32705,N_21707,N_28007);
xnor U32706 (N_32706,N_23830,N_26437);
nor U32707 (N_32707,N_20690,N_24270);
and U32708 (N_32708,N_26935,N_25405);
nand U32709 (N_32709,N_28709,N_21795);
nor U32710 (N_32710,N_27257,N_27254);
nand U32711 (N_32711,N_29011,N_23115);
xor U32712 (N_32712,N_24424,N_27985);
or U32713 (N_32713,N_20790,N_27573);
nand U32714 (N_32714,N_21716,N_27987);
or U32715 (N_32715,N_28951,N_23838);
or U32716 (N_32716,N_21792,N_27436);
xnor U32717 (N_32717,N_24974,N_21046);
nor U32718 (N_32718,N_20022,N_26672);
nand U32719 (N_32719,N_29807,N_29301);
and U32720 (N_32720,N_27346,N_23963);
nor U32721 (N_32721,N_26240,N_29117);
xor U32722 (N_32722,N_26885,N_24491);
xnor U32723 (N_32723,N_27215,N_25495);
xor U32724 (N_32724,N_26250,N_21761);
and U32725 (N_32725,N_24858,N_23070);
nand U32726 (N_32726,N_20028,N_24347);
nor U32727 (N_32727,N_27052,N_25910);
xnor U32728 (N_32728,N_20848,N_25938);
xnor U32729 (N_32729,N_24730,N_20429);
nor U32730 (N_32730,N_23334,N_29934);
and U32731 (N_32731,N_20996,N_29396);
nor U32732 (N_32732,N_24992,N_25706);
or U32733 (N_32733,N_26550,N_22712);
and U32734 (N_32734,N_21273,N_29653);
nand U32735 (N_32735,N_26054,N_24080);
or U32736 (N_32736,N_26014,N_25085);
and U32737 (N_32737,N_23621,N_27914);
xnor U32738 (N_32738,N_20312,N_29424);
or U32739 (N_32739,N_25596,N_22177);
and U32740 (N_32740,N_23391,N_22241);
or U32741 (N_32741,N_23975,N_25398);
and U32742 (N_32742,N_22155,N_28033);
nor U32743 (N_32743,N_28557,N_28020);
or U32744 (N_32744,N_23238,N_20874);
or U32745 (N_32745,N_25067,N_28374);
and U32746 (N_32746,N_28885,N_21738);
and U32747 (N_32747,N_20131,N_22825);
or U32748 (N_32748,N_24056,N_26956);
and U32749 (N_32749,N_26289,N_25620);
nand U32750 (N_32750,N_22635,N_21086);
or U32751 (N_32751,N_29230,N_24669);
nand U32752 (N_32752,N_28486,N_28834);
and U32753 (N_32753,N_21782,N_28895);
and U32754 (N_32754,N_22168,N_26921);
nor U32755 (N_32755,N_25073,N_22503);
or U32756 (N_32756,N_27740,N_20033);
or U32757 (N_32757,N_26490,N_27766);
and U32758 (N_32758,N_28681,N_22659);
nor U32759 (N_32759,N_23172,N_21540);
nor U32760 (N_32760,N_23742,N_27835);
or U32761 (N_32761,N_20794,N_26991);
and U32762 (N_32762,N_26409,N_29875);
and U32763 (N_32763,N_22128,N_22136);
or U32764 (N_32764,N_23762,N_25826);
nor U32765 (N_32765,N_24399,N_22871);
nand U32766 (N_32766,N_20333,N_24881);
or U32767 (N_32767,N_22307,N_24577);
and U32768 (N_32768,N_27491,N_26755);
and U32769 (N_32769,N_26575,N_21848);
or U32770 (N_32770,N_27280,N_27132);
or U32771 (N_32771,N_21821,N_23089);
and U32772 (N_32772,N_25899,N_29582);
nor U32773 (N_32773,N_24686,N_27457);
nand U32774 (N_32774,N_22106,N_27836);
nor U32775 (N_32775,N_21002,N_22881);
and U32776 (N_32776,N_27583,N_21804);
and U32777 (N_32777,N_22238,N_28686);
nand U32778 (N_32778,N_25534,N_26620);
or U32779 (N_32779,N_28963,N_29660);
or U32780 (N_32780,N_29849,N_27362);
xnor U32781 (N_32781,N_29629,N_26811);
and U32782 (N_32782,N_28463,N_23707);
nor U32783 (N_32783,N_20284,N_20864);
nor U32784 (N_32784,N_22834,N_26618);
and U32785 (N_32785,N_28308,N_29185);
and U32786 (N_32786,N_25737,N_23531);
xor U32787 (N_32787,N_23790,N_21613);
and U32788 (N_32788,N_21985,N_20896);
nand U32789 (N_32789,N_23119,N_20974);
and U32790 (N_32790,N_29189,N_27781);
and U32791 (N_32791,N_24282,N_22246);
or U32792 (N_32792,N_23199,N_21247);
nand U32793 (N_32793,N_27794,N_27309);
xor U32794 (N_32794,N_29862,N_24319);
nor U32795 (N_32795,N_26367,N_20264);
and U32796 (N_32796,N_20823,N_28957);
and U32797 (N_32797,N_21552,N_29621);
or U32798 (N_32798,N_25632,N_20752);
or U32799 (N_32799,N_21949,N_23389);
nand U32800 (N_32800,N_29349,N_20224);
nor U32801 (N_32801,N_24890,N_21014);
or U32802 (N_32802,N_26008,N_21843);
xnor U32803 (N_32803,N_21384,N_29561);
and U32804 (N_32804,N_20094,N_26685);
or U32805 (N_32805,N_26927,N_28967);
nand U32806 (N_32806,N_26776,N_25113);
nor U32807 (N_32807,N_28389,N_26777);
nor U32808 (N_32808,N_24790,N_29900);
xnor U32809 (N_32809,N_27778,N_28566);
and U32810 (N_32810,N_25821,N_28661);
nor U32811 (N_32811,N_21943,N_28062);
or U32812 (N_32812,N_29865,N_23095);
xnor U32813 (N_32813,N_22281,N_28528);
xnor U32814 (N_32814,N_25281,N_29312);
and U32815 (N_32815,N_20604,N_26111);
nand U32816 (N_32816,N_23168,N_23928);
or U32817 (N_32817,N_29091,N_28114);
nand U32818 (N_32818,N_24368,N_29113);
nand U32819 (N_32819,N_23124,N_23005);
nand U32820 (N_32820,N_22487,N_24632);
xnor U32821 (N_32821,N_24797,N_21175);
and U32822 (N_32822,N_22734,N_29699);
nand U32823 (N_32823,N_26257,N_28037);
nand U32824 (N_32824,N_23771,N_20991);
or U32825 (N_32825,N_24213,N_23122);
and U32826 (N_32826,N_28046,N_29508);
nand U32827 (N_32827,N_22923,N_26820);
nor U32828 (N_32828,N_20685,N_20214);
and U32829 (N_32829,N_27106,N_24920);
or U32830 (N_32830,N_28041,N_20064);
and U32831 (N_32831,N_21185,N_28618);
or U32832 (N_32832,N_25267,N_21802);
xor U32833 (N_32833,N_28307,N_25418);
nor U32834 (N_32834,N_29579,N_29378);
xor U32835 (N_32835,N_23618,N_20130);
or U32836 (N_32836,N_22715,N_26498);
and U32837 (N_32837,N_20208,N_21917);
and U32838 (N_32838,N_28484,N_25600);
xor U32839 (N_32839,N_21538,N_26959);
or U32840 (N_32840,N_23273,N_27760);
and U32841 (N_32841,N_21111,N_24266);
or U32842 (N_32842,N_20520,N_25595);
or U32843 (N_32843,N_28048,N_20895);
and U32844 (N_32844,N_23733,N_25744);
nand U32845 (N_32845,N_20345,N_29822);
and U32846 (N_32846,N_29038,N_26463);
and U32847 (N_32847,N_24705,N_23322);
xor U32848 (N_32848,N_26332,N_21534);
xnor U32849 (N_32849,N_20476,N_22245);
xnor U32850 (N_32850,N_25685,N_22009);
or U32851 (N_32851,N_29446,N_22580);
nor U32852 (N_32852,N_23158,N_24040);
or U32853 (N_32853,N_21953,N_21769);
nor U32854 (N_32854,N_28576,N_25571);
xor U32855 (N_32855,N_27364,N_22536);
nand U32856 (N_32856,N_20043,N_28707);
and U32857 (N_32857,N_25012,N_26975);
and U32858 (N_32858,N_25114,N_21572);
nand U32859 (N_32859,N_28223,N_21702);
nand U32860 (N_32860,N_22930,N_27175);
or U32861 (N_32861,N_26948,N_29800);
or U32862 (N_32862,N_27843,N_21952);
nor U32863 (N_32863,N_23440,N_26271);
or U32864 (N_32864,N_26035,N_24563);
nor U32865 (N_32865,N_22132,N_22366);
or U32866 (N_32866,N_23513,N_26263);
nor U32867 (N_32867,N_27992,N_26568);
and U32868 (N_32868,N_26085,N_22668);
xnor U32869 (N_32869,N_21225,N_26101);
nand U32870 (N_32870,N_26365,N_24496);
nand U32871 (N_32871,N_20952,N_26539);
nand U32872 (N_32872,N_28161,N_28877);
nand U32873 (N_32873,N_28648,N_25774);
nand U32874 (N_32874,N_26837,N_28369);
nand U32875 (N_32875,N_29151,N_26671);
nor U32876 (N_32876,N_26087,N_20691);
and U32877 (N_32877,N_20608,N_23699);
or U32878 (N_32878,N_26272,N_25522);
nand U32879 (N_32879,N_25191,N_28620);
nand U32880 (N_32880,N_21809,N_21581);
xor U32881 (N_32881,N_27900,N_22457);
nand U32882 (N_32882,N_28283,N_22229);
xnor U32883 (N_32883,N_20086,N_21393);
xnor U32884 (N_32884,N_22893,N_29075);
or U32885 (N_32885,N_25720,N_24956);
and U32886 (N_32886,N_26028,N_21301);
nor U32887 (N_32887,N_27530,N_23763);
nor U32888 (N_32888,N_21691,N_25439);
xnor U32889 (N_32889,N_25604,N_21205);
nand U32890 (N_32890,N_26185,N_27722);
xor U32891 (N_32891,N_20307,N_28506);
or U32892 (N_32892,N_20299,N_24065);
xor U32893 (N_32893,N_20117,N_27559);
nor U32894 (N_32894,N_26772,N_28803);
or U32895 (N_32895,N_27973,N_29351);
xor U32896 (N_32896,N_27552,N_21053);
xnor U32897 (N_32897,N_28828,N_26986);
or U32898 (N_32898,N_24545,N_28393);
and U32899 (N_32899,N_21740,N_23256);
nor U32900 (N_32900,N_20141,N_26299);
xnor U32901 (N_32901,N_23174,N_24512);
and U32902 (N_32902,N_29110,N_24164);
xor U32903 (N_32903,N_20720,N_21813);
or U32904 (N_32904,N_26700,N_25285);
nand U32905 (N_32905,N_27242,N_29245);
nand U32906 (N_32906,N_28296,N_28169);
nand U32907 (N_32907,N_24821,N_21564);
or U32908 (N_32908,N_21356,N_27888);
xor U32909 (N_32909,N_29926,N_26326);
nand U32910 (N_32910,N_20001,N_26566);
and U32911 (N_32911,N_25133,N_29205);
or U32912 (N_32912,N_22535,N_23598);
and U32913 (N_32913,N_21178,N_28733);
or U32914 (N_32914,N_27228,N_21087);
xor U32915 (N_32915,N_29015,N_24733);
and U32916 (N_32916,N_25211,N_21935);
and U32917 (N_32917,N_20414,N_21470);
nor U32918 (N_32918,N_27499,N_21414);
nor U32919 (N_32919,N_21885,N_23626);
nand U32920 (N_32920,N_21911,N_24746);
and U32921 (N_32921,N_20540,N_25423);
nand U32922 (N_32922,N_28961,N_27060);
nor U32923 (N_32923,N_26038,N_24371);
nand U32924 (N_32924,N_29131,N_23380);
xnor U32925 (N_32925,N_25433,N_27131);
nand U32926 (N_32926,N_25680,N_25662);
or U32927 (N_32927,N_27005,N_20433);
and U32928 (N_32928,N_25520,N_29569);
nor U32929 (N_32929,N_20087,N_21828);
nand U32930 (N_32930,N_23123,N_21685);
xnor U32931 (N_32931,N_27730,N_27871);
xor U32932 (N_32932,N_23630,N_29835);
xor U32933 (N_32933,N_24538,N_27810);
or U32934 (N_32934,N_22278,N_24335);
nand U32935 (N_32935,N_28127,N_25295);
or U32936 (N_32936,N_21359,N_23848);
nand U32937 (N_32937,N_26659,N_22873);
and U32938 (N_32938,N_28441,N_23155);
nand U32939 (N_32939,N_27124,N_27748);
or U32940 (N_32940,N_25205,N_23972);
or U32941 (N_32941,N_27608,N_21748);
nand U32942 (N_32942,N_28558,N_23293);
nor U32943 (N_32943,N_22805,N_29167);
or U32944 (N_32944,N_28713,N_21757);
or U32945 (N_32945,N_22926,N_21055);
xor U32946 (N_32946,N_22051,N_24670);
xnor U32947 (N_32947,N_21019,N_25357);
xnor U32948 (N_32948,N_25380,N_24357);
nand U32949 (N_32949,N_29240,N_28526);
xor U32950 (N_32950,N_27185,N_23313);
nand U32951 (N_32951,N_28150,N_25440);
or U32952 (N_32952,N_23037,N_24045);
nand U32953 (N_32953,N_25513,N_29153);
xnor U32954 (N_32954,N_24415,N_27352);
xnor U32955 (N_32955,N_29332,N_26597);
nor U32956 (N_32956,N_20932,N_21990);
or U32957 (N_32957,N_20869,N_20065);
and U32958 (N_32958,N_26725,N_21631);
xor U32959 (N_32959,N_27404,N_22821);
nand U32960 (N_32960,N_26308,N_21960);
xor U32961 (N_32961,N_23402,N_29218);
nand U32962 (N_32962,N_25936,N_27373);
nand U32963 (N_32963,N_22020,N_27122);
and U32964 (N_32964,N_26794,N_24258);
and U32965 (N_32965,N_29979,N_29705);
nor U32966 (N_32966,N_28073,N_20616);
xnor U32967 (N_32967,N_29455,N_25334);
nor U32968 (N_32968,N_29716,N_25286);
nand U32969 (N_32969,N_23984,N_26068);
or U32970 (N_32970,N_29366,N_24438);
or U32971 (N_32971,N_20579,N_29970);
nand U32972 (N_32972,N_25208,N_28568);
and U32973 (N_32973,N_21166,N_25792);
and U32974 (N_32974,N_26576,N_22335);
and U32975 (N_32975,N_22595,N_21191);
and U32976 (N_32976,N_22800,N_21361);
xnor U32977 (N_32977,N_29070,N_27430);
xor U32978 (N_32978,N_26836,N_23128);
or U32979 (N_32979,N_22162,N_20397);
nor U32980 (N_32980,N_27424,N_22733);
xnor U32981 (N_32981,N_25304,N_20349);
or U32982 (N_32982,N_23350,N_23336);
nor U32983 (N_32983,N_24765,N_27506);
nor U32984 (N_32984,N_20475,N_26143);
nand U32985 (N_32985,N_24846,N_24361);
and U32986 (N_32986,N_28110,N_21224);
or U32987 (N_32987,N_24610,N_28025);
and U32988 (N_32988,N_20639,N_24793);
and U32989 (N_32989,N_23846,N_25322);
nand U32990 (N_32990,N_23176,N_24092);
or U32991 (N_32991,N_25008,N_28072);
nand U32992 (N_32992,N_25161,N_25284);
or U32993 (N_32993,N_25307,N_29195);
or U32994 (N_32994,N_28913,N_28652);
xnor U32995 (N_32995,N_23893,N_22361);
nand U32996 (N_32996,N_20063,N_28147);
nand U32997 (N_32997,N_26497,N_23132);
or U32998 (N_32998,N_24527,N_22369);
nand U32999 (N_32999,N_25863,N_24839);
or U33000 (N_33000,N_26235,N_21918);
or U33001 (N_33001,N_25396,N_27663);
nor U33002 (N_33002,N_20569,N_29206);
xnor U33003 (N_33003,N_29933,N_28613);
nand U33004 (N_33004,N_23143,N_27847);
or U33005 (N_33005,N_24121,N_25177);
xor U33006 (N_33006,N_28914,N_28442);
and U33007 (N_33007,N_23360,N_27141);
nor U33008 (N_33008,N_22966,N_21741);
nand U33009 (N_33009,N_24937,N_20113);
xnor U33010 (N_33010,N_28273,N_25017);
or U33011 (N_33011,N_27476,N_22654);
and U33012 (N_33012,N_28346,N_20628);
nor U33013 (N_33013,N_28640,N_27345);
nand U33014 (N_33014,N_29553,N_20911);
nor U33015 (N_33015,N_26415,N_23660);
xor U33016 (N_33016,N_22332,N_29657);
and U33017 (N_33017,N_25830,N_20202);
or U33018 (N_33018,N_26113,N_24297);
nand U33019 (N_33019,N_27440,N_29276);
nor U33020 (N_33020,N_28331,N_28827);
nand U33021 (N_33021,N_27140,N_28881);
and U33022 (N_33022,N_23999,N_27999);
and U33023 (N_33023,N_22042,N_24910);
xor U33024 (N_33024,N_26039,N_21535);
nand U33025 (N_33025,N_24277,N_21628);
and U33026 (N_33026,N_27849,N_28984);
and U33027 (N_33027,N_21591,N_28178);
nand U33028 (N_33028,N_26018,N_28856);
or U33029 (N_33029,N_20737,N_22196);
and U33030 (N_33030,N_21737,N_21027);
and U33031 (N_33031,N_22648,N_27824);
nor U33032 (N_33032,N_29847,N_25249);
and U33033 (N_33033,N_22751,N_24044);
nand U33034 (N_33034,N_25152,N_28367);
or U33035 (N_33035,N_21090,N_20578);
xor U33036 (N_33036,N_29253,N_25092);
xnor U33037 (N_33037,N_29305,N_24373);
nand U33038 (N_33038,N_27746,N_23745);
or U33039 (N_33039,N_24808,N_22693);
and U33040 (N_33040,N_21672,N_27926);
or U33041 (N_33041,N_27266,N_20176);
nor U33042 (N_33042,N_20146,N_29324);
nand U33043 (N_33043,N_27854,N_21342);
and U33044 (N_33044,N_28452,N_28738);
nand U33045 (N_33045,N_29078,N_21397);
nand U33046 (N_33046,N_22193,N_28102);
and U33047 (N_33047,N_28466,N_25960);
xor U33048 (N_33048,N_22645,N_29651);
nand U33049 (N_33049,N_24240,N_29065);
xor U33050 (N_33050,N_28854,N_29311);
and U33051 (N_33051,N_26088,N_25730);
or U33052 (N_33052,N_20056,N_22925);
or U33053 (N_33053,N_22978,N_26970);
nor U33054 (N_33054,N_27919,N_29895);
nand U33055 (N_33055,N_27776,N_26454);
and U33056 (N_33056,N_27901,N_21840);
or U33057 (N_33057,N_29664,N_28532);
xnor U33058 (N_33058,N_20964,N_21362);
nand U33059 (N_33059,N_27961,N_21637);
xor U33060 (N_33060,N_28100,N_27686);
nor U33061 (N_33061,N_26078,N_26923);
or U33062 (N_33062,N_27816,N_21344);
xor U33063 (N_33063,N_24769,N_21882);
xnor U33064 (N_33064,N_26679,N_20978);
xnor U33065 (N_33065,N_21196,N_27026);
xnor U33066 (N_33066,N_25402,N_21116);
nor U33067 (N_33067,N_22957,N_28717);
and U33068 (N_33068,N_20813,N_22060);
and U33069 (N_33069,N_28315,N_22932);
nor U33070 (N_33070,N_21496,N_21499);
nor U33071 (N_33071,N_21666,N_21932);
or U33072 (N_33072,N_27576,N_29602);
nand U33073 (N_33073,N_25932,N_28667);
or U33074 (N_33074,N_24236,N_24465);
and U33075 (N_33075,N_21862,N_24464);
and U33076 (N_33076,N_25841,N_25376);
and U33077 (N_33077,N_29192,N_21001);
or U33078 (N_33078,N_25485,N_26690);
nor U33079 (N_33079,N_26501,N_21266);
nor U33080 (N_33080,N_21095,N_25431);
xnor U33081 (N_33081,N_22824,N_23419);
nand U33082 (N_33082,N_20834,N_26936);
and U33083 (N_33083,N_24151,N_25689);
nor U33084 (N_33084,N_23966,N_29046);
nor U33085 (N_33085,N_20380,N_23612);
xnor U33086 (N_33086,N_25619,N_23436);
nor U33087 (N_33087,N_24983,N_26199);
nand U33088 (N_33088,N_26624,N_26995);
nand U33089 (N_33089,N_28925,N_23250);
nand U33090 (N_33090,N_29993,N_22019);
xnor U33091 (N_33091,N_25041,N_22108);
or U33092 (N_33092,N_26205,N_29157);
nand U33093 (N_33093,N_28254,N_29543);
nor U33094 (N_33094,N_28644,N_22445);
and U33095 (N_33095,N_20804,N_27558);
and U33096 (N_33096,N_27433,N_21688);
or U33097 (N_33097,N_25383,N_22742);
and U33098 (N_33098,N_26615,N_21254);
and U33099 (N_33099,N_24299,N_23589);
nand U33100 (N_33100,N_26007,N_27868);
nand U33101 (N_33101,N_21853,N_28311);
xnor U33102 (N_33102,N_27875,N_20492);
nand U33103 (N_33103,N_29818,N_20884);
xor U33104 (N_33104,N_28200,N_24599);
nand U33105 (N_33105,N_28998,N_28773);
and U33106 (N_33106,N_26655,N_26259);
xnor U33107 (N_33107,N_27458,N_29379);
nand U33108 (N_33108,N_21345,N_26013);
or U33109 (N_33109,N_26598,N_25760);
and U33110 (N_33110,N_22372,N_27068);
xnor U33111 (N_33111,N_24575,N_27517);
or U33112 (N_33112,N_29460,N_21075);
nand U33113 (N_33113,N_20304,N_27519);
nor U33114 (N_33114,N_25836,N_27995);
nor U33115 (N_33115,N_26009,N_22958);
nor U33116 (N_33116,N_21711,N_26955);
or U33117 (N_33117,N_25800,N_24280);
nand U33118 (N_33118,N_20767,N_25634);
or U33119 (N_33119,N_28094,N_25347);
nand U33120 (N_33120,N_28919,N_28930);
nor U33121 (N_33121,N_23674,N_23921);
and U33122 (N_33122,N_28372,N_26396);
nor U33123 (N_33123,N_28035,N_28251);
xnor U33124 (N_33124,N_21554,N_24544);
or U33125 (N_33125,N_25629,N_29267);
nor U33126 (N_33126,N_25585,N_26356);
nand U33127 (N_33127,N_22897,N_27619);
xor U33128 (N_33128,N_20493,N_20468);
or U33129 (N_33129,N_26527,N_26766);
and U33130 (N_33130,N_21889,N_29329);
and U33131 (N_33131,N_21652,N_22320);
nor U33132 (N_33132,N_24709,N_25214);
or U33133 (N_33133,N_27636,N_28527);
nand U33134 (N_33134,N_26838,N_27998);
nor U33135 (N_33135,N_27006,N_25703);
nor U33136 (N_33136,N_25318,N_24376);
and U33137 (N_33137,N_29448,N_24255);
nand U33138 (N_33138,N_22221,N_22378);
nor U33139 (N_33139,N_20633,N_25366);
nand U33140 (N_33140,N_25151,N_29435);
nor U33141 (N_33141,N_25233,N_23237);
nor U33142 (N_33142,N_28597,N_22216);
nor U33143 (N_33143,N_26642,N_24325);
xor U33144 (N_33144,N_24558,N_27790);
and U33145 (N_33145,N_20739,N_20607);
or U33146 (N_33146,N_20451,N_24272);
xor U33147 (N_33147,N_29322,N_26441);
xnor U33148 (N_33148,N_23289,N_24773);
nor U33149 (N_33149,N_29766,N_23706);
nand U33150 (N_33150,N_25024,N_27209);
or U33151 (N_33151,N_26577,N_21239);
and U33152 (N_33152,N_24036,N_24689);
nand U33153 (N_33153,N_22626,N_20102);
xnor U33154 (N_33154,N_20055,N_22078);
and U33155 (N_33155,N_28487,N_25880);
or U33156 (N_33156,N_20439,N_20019);
nand U33157 (N_33157,N_26127,N_29433);
xnor U33158 (N_33158,N_24147,N_26763);
nor U33159 (N_33159,N_29845,N_21981);
or U33160 (N_33160,N_20531,N_21382);
xor U33161 (N_33161,N_27743,N_25636);
xor U33162 (N_33162,N_27479,N_26675);
nor U33163 (N_33163,N_29840,N_26552);
nand U33164 (N_33164,N_24287,N_26530);
and U33165 (N_33165,N_22697,N_29277);
nand U33166 (N_33166,N_29588,N_24993);
and U33167 (N_33167,N_28628,N_26485);
nor U33168 (N_33168,N_28421,N_26024);
or U33169 (N_33169,N_22373,N_23448);
nand U33170 (N_33170,N_28225,N_24759);
nand U33171 (N_33171,N_25697,N_24947);
or U33172 (N_33172,N_26688,N_25825);
and U33173 (N_33173,N_26218,N_26064);
nand U33174 (N_33174,N_21299,N_21511);
nand U33175 (N_33175,N_24344,N_26283);
nand U33176 (N_33176,N_20734,N_25518);
or U33177 (N_33177,N_25429,N_29346);
nand U33178 (N_33178,N_23616,N_26996);
nor U33179 (N_33179,N_27038,N_23989);
nand U33180 (N_33180,N_24071,N_25381);
xor U33181 (N_33181,N_22736,N_29782);
nand U33182 (N_33182,N_22656,N_28278);
nand U33183 (N_33183,N_27947,N_23640);
nor U33184 (N_33184,N_27889,N_20860);
nor U33185 (N_33185,N_24833,N_27811);
or U33186 (N_33186,N_25814,N_27162);
or U33187 (N_33187,N_20108,N_27933);
and U33188 (N_33188,N_26466,N_22968);
nand U33189 (N_33189,N_20980,N_22176);
nand U33190 (N_33190,N_28433,N_25330);
nor U33191 (N_33191,N_22355,N_27952);
and U33192 (N_33192,N_20516,N_29160);
xor U33193 (N_33193,N_26350,N_28173);
and U33194 (N_33194,N_22700,N_27088);
xnor U33195 (N_33195,N_28993,N_28424);
xor U33196 (N_33196,N_26593,N_23882);
and U33197 (N_33197,N_28599,N_28027);
or U33198 (N_33198,N_28544,N_25135);
nor U33199 (N_33199,N_20732,N_20759);
nor U33200 (N_33200,N_22331,N_21313);
and U33201 (N_33201,N_21756,N_20067);
nor U33202 (N_33202,N_23253,N_24907);
or U33203 (N_33203,N_22592,N_26420);
nor U33204 (N_33204,N_27575,N_25182);
and U33205 (N_33205,N_25771,N_23802);
and U33206 (N_33206,N_22201,N_27822);
xnor U33207 (N_33207,N_20593,N_28518);
and U33208 (N_33208,N_27913,N_25642);
or U33209 (N_33209,N_28265,N_27643);
nand U33210 (N_33210,N_26717,N_22501);
and U33211 (N_33211,N_28286,N_28111);
xor U33212 (N_33212,N_21669,N_23877);
xor U33213 (N_33213,N_25028,N_28555);
and U33214 (N_33214,N_23711,N_27726);
xor U33215 (N_33215,N_29517,N_23623);
xor U33216 (N_33216,N_24471,N_26507);
and U33217 (N_33217,N_26407,N_27252);
xnor U33218 (N_33218,N_27887,N_25639);
nor U33219 (N_33219,N_29274,N_22044);
nor U33220 (N_33220,N_20988,N_24593);
or U33221 (N_33221,N_29462,N_25516);
nand U33222 (N_33222,N_21819,N_23296);
or U33223 (N_33223,N_25445,N_28138);
nor U33224 (N_33224,N_20487,N_22003);
or U33225 (N_33225,N_27234,N_21995);
nand U33226 (N_33226,N_24029,N_24276);
nand U33227 (N_33227,N_29300,N_21447);
nand U33228 (N_33228,N_20337,N_24649);
or U33229 (N_33229,N_24490,N_27076);
xor U33230 (N_33230,N_20204,N_23543);
nand U33231 (N_33231,N_27379,N_24393);
or U33232 (N_33232,N_27862,N_29478);
xor U33233 (N_33233,N_27051,N_29482);
and U33234 (N_33234,N_27152,N_20600);
or U33235 (N_33235,N_27217,N_27893);
nand U33236 (N_33236,N_22714,N_28247);
nand U33237 (N_33237,N_22651,N_22950);
xor U33238 (N_33238,N_20210,N_24146);
nor U33239 (N_33239,N_24924,N_26144);
or U33240 (N_33240,N_29024,N_22579);
nand U33241 (N_33241,N_27842,N_24382);
xor U33242 (N_33242,N_29813,N_24316);
or U33243 (N_33243,N_24708,N_24116);
nand U33244 (N_33244,N_25120,N_21290);
or U33245 (N_33245,N_21131,N_21357);
nor U33246 (N_33246,N_21324,N_21279);
or U33247 (N_33247,N_21638,N_29757);
and U33248 (N_33248,N_26591,N_24074);
nor U33249 (N_33249,N_21619,N_28269);
or U33250 (N_33250,N_20818,N_23326);
and U33251 (N_33251,N_21799,N_26044);
xor U33252 (N_33252,N_26826,N_25500);
or U33253 (N_33253,N_25660,N_25715);
nand U33254 (N_33254,N_27890,N_29123);
xnor U33255 (N_33255,N_26412,N_20168);
nand U33256 (N_33256,N_24134,N_26027);
nand U33257 (N_33257,N_24338,N_29819);
nor U33258 (N_33258,N_29431,N_23792);
nor U33259 (N_33259,N_26564,N_26967);
nor U33260 (N_33260,N_20234,N_28698);
nand U33261 (N_33261,N_20095,N_24862);
or U33262 (N_33262,N_26732,N_27942);
xnor U33263 (N_33263,N_21816,N_21456);
nand U33264 (N_33264,N_28103,N_24953);
nand U33265 (N_33265,N_24801,N_28978);
nor U33266 (N_33266,N_25588,N_25972);
and U33267 (N_33267,N_20742,N_28356);
nor U33268 (N_33268,N_21180,N_26912);
xor U33269 (N_33269,N_24472,N_23780);
xnor U33270 (N_33270,N_28743,N_24503);
and U33271 (N_33271,N_26156,N_23575);
xor U33272 (N_33272,N_22370,N_27078);
or U33273 (N_33273,N_28637,N_24084);
nand U33274 (N_33274,N_22621,N_27883);
xor U33275 (N_33275,N_23675,N_25060);
or U33276 (N_33276,N_27147,N_27418);
nor U33277 (N_33277,N_20192,N_22927);
nand U33278 (N_33278,N_27108,N_26965);
and U33279 (N_33279,N_24366,N_25279);
or U33280 (N_33280,N_28135,N_20692);
or U33281 (N_33281,N_23178,N_27452);
nand U33282 (N_33282,N_20733,N_24567);
and U33283 (N_33283,N_24286,N_23511);
or U33284 (N_33284,N_22311,N_29546);
xor U33285 (N_33285,N_29676,N_29938);
or U33286 (N_33286,N_24752,N_27334);
and U33287 (N_33287,N_22519,N_21160);
nand U33288 (N_33288,N_23288,N_27302);
nor U33289 (N_33289,N_26083,N_20660);
and U33290 (N_33290,N_21857,N_22130);
and U33291 (N_33291,N_26702,N_22358);
xor U33292 (N_33292,N_23602,N_29898);
and U33293 (N_33293,N_28723,N_29951);
nand U33294 (N_33294,N_20440,N_22627);
nor U33295 (N_33295,N_21385,N_28137);
or U33296 (N_33296,N_23175,N_22237);
xor U33297 (N_33297,N_23302,N_21759);
xnor U33298 (N_33298,N_23639,N_26427);
nand U33299 (N_33299,N_27323,N_23788);
and U33300 (N_33300,N_23353,N_28368);
or U33301 (N_33301,N_25867,N_21794);
xnor U33302 (N_33302,N_29871,N_20421);
and U33303 (N_33303,N_21194,N_22391);
nand U33304 (N_33304,N_27724,N_26753);
or U33305 (N_33305,N_23388,N_21768);
xnor U33306 (N_33306,N_23528,N_26324);
nand U33307 (N_33307,N_22899,N_22772);
nand U33308 (N_33308,N_21665,N_20764);
nand U33309 (N_33309,N_21381,N_20404);
xnor U33310 (N_33310,N_29536,N_25998);
nor U33311 (N_33311,N_26429,N_26141);
nand U33312 (N_33312,N_25735,N_28609);
xnor U33313 (N_33313,N_27187,N_27529);
and U33314 (N_33314,N_20689,N_29722);
and U33315 (N_33315,N_28843,N_20377);
xnor U33316 (N_33316,N_20713,N_20880);
nor U33317 (N_33317,N_27104,N_28654);
or U33318 (N_33318,N_26968,N_20935);
nand U33319 (N_33319,N_29116,N_21411);
and U33320 (N_33320,N_29816,N_28475);
nor U33321 (N_33321,N_24193,N_25058);
or U33322 (N_33322,N_25966,N_25202);
nand U33323 (N_33323,N_28505,N_29646);
nor U33324 (N_33324,N_26878,N_24802);
nand U33325 (N_33325,N_24008,N_27210);
nand U33326 (N_33326,N_29885,N_29150);
or U33327 (N_33327,N_27387,N_23371);
nand U33328 (N_33328,N_20464,N_25027);
and U33329 (N_33329,N_28987,N_28941);
or U33330 (N_33330,N_22692,N_21141);
and U33331 (N_33331,N_23978,N_21274);
or U33332 (N_33332,N_21908,N_24722);
xor U33333 (N_33333,N_22753,N_23544);
xor U33334 (N_33334,N_25725,N_23453);
nand U33335 (N_33335,N_24728,N_22500);
or U33336 (N_33336,N_29555,N_26377);
nor U33337 (N_33337,N_23871,N_27475);
xnor U33338 (N_33338,N_24181,N_22288);
and U33339 (N_33339,N_23655,N_26829);
nand U33340 (N_33340,N_27808,N_23670);
nand U33341 (N_33341,N_26946,N_27035);
and U33342 (N_33342,N_20419,N_24379);
xnor U33343 (N_33343,N_22774,N_26483);
xor U33344 (N_33344,N_20037,N_20405);
nand U33345 (N_33345,N_20186,N_26161);
nor U33346 (N_33346,N_24972,N_23307);
nand U33347 (N_33347,N_20567,N_23335);
and U33348 (N_33348,N_27269,N_29680);
xor U33349 (N_33349,N_24278,N_24158);
nor U33350 (N_33350,N_21417,N_20883);
or U33351 (N_33351,N_28742,N_28783);
or U33352 (N_33352,N_20956,N_23432);
nor U33353 (N_33353,N_28688,N_20510);
nor U33354 (N_33354,N_21601,N_20636);
nor U33355 (N_33355,N_29810,N_24000);
nor U33356 (N_33356,N_22035,N_20344);
and U33357 (N_33357,N_28318,N_29990);
xor U33358 (N_33358,N_23473,N_26153);
nand U33359 (N_33359,N_24804,N_20413);
nand U33360 (N_33360,N_24311,N_29706);
xnor U33361 (N_33361,N_21651,N_20757);
and U33362 (N_33362,N_29381,N_26953);
nor U33363 (N_33363,N_29919,N_20184);
nand U33364 (N_33364,N_21726,N_21486);
nor U33365 (N_33365,N_22376,N_21790);
nor U33366 (N_33366,N_20266,N_28815);
xor U33367 (N_33367,N_26357,N_27338);
and U33368 (N_33368,N_28992,N_25248);
and U33369 (N_33369,N_22489,N_20007);
or U33370 (N_33370,N_28336,N_23035);
or U33371 (N_33371,N_28622,N_29985);
or U33372 (N_33372,N_27918,N_28323);
nand U33373 (N_33373,N_28605,N_29718);
and U33374 (N_33374,N_22522,N_27727);
xnor U33375 (N_33375,N_23315,N_27426);
or U33376 (N_33376,N_22541,N_25478);
nand U33377 (N_33377,N_21028,N_26422);
nor U33378 (N_33378,N_24140,N_20632);
nand U33379 (N_33379,N_29689,N_21138);
nand U33380 (N_33380,N_23658,N_22523);
nand U33381 (N_33381,N_20652,N_24057);
nand U33382 (N_33382,N_26781,N_21687);
or U33383 (N_33383,N_24192,N_25461);
and U33384 (N_33384,N_29776,N_21311);
or U33385 (N_33385,N_29356,N_27330);
or U33386 (N_33386,N_29143,N_22642);
or U33387 (N_33387,N_23596,N_24149);
nand U33388 (N_33388,N_22940,N_27240);
and U33389 (N_33389,N_24502,N_22723);
xnor U33390 (N_33390,N_29297,N_27534);
xnor U33391 (N_33391,N_22096,N_21927);
and U33392 (N_33392,N_22947,N_24905);
nand U33393 (N_33393,N_21934,N_28805);
nand U33394 (N_33394,N_23375,N_26851);
or U33395 (N_33395,N_26266,N_26426);
or U33396 (N_33396,N_20237,N_22440);
and U33397 (N_33397,N_22827,N_28798);
nor U33398 (N_33398,N_28258,N_29918);
or U33399 (N_33399,N_26733,N_29178);
nand U33400 (N_33400,N_20903,N_20775);
xnor U33401 (N_33401,N_24296,N_23159);
nand U33402 (N_33402,N_24597,N_28250);
or U33403 (N_33403,N_22283,N_25296);
and U33404 (N_33404,N_20240,N_29344);
nor U33405 (N_33405,N_26869,N_24026);
nor U33406 (N_33406,N_29801,N_28795);
xor U33407 (N_33407,N_29188,N_22776);
nor U33408 (N_33408,N_20666,N_21896);
nor U33409 (N_33409,N_23677,N_22578);
nand U33410 (N_33410,N_28467,N_21182);
and U33411 (N_33411,N_29406,N_27631);
and U33412 (N_33412,N_22268,N_20542);
nand U33413 (N_33413,N_26285,N_26799);
nand U33414 (N_33414,N_25658,N_20238);
nor U33415 (N_33415,N_23515,N_28183);
nor U33416 (N_33416,N_28838,N_24194);
nor U33417 (N_33417,N_22488,N_23836);
and U33418 (N_33418,N_29463,N_20418);
and U33419 (N_33419,N_25019,N_28509);
and U33420 (N_33420,N_24780,N_23261);
nand U33421 (N_33421,N_24225,N_26423);
nor U33422 (N_33422,N_25319,N_21841);
or U33423 (N_33423,N_23487,N_28573);
or U33424 (N_33424,N_26863,N_27677);
xnor U33425 (N_33425,N_23169,N_23381);
nand U33426 (N_33426,N_23774,N_25950);
nand U33427 (N_33427,N_28005,N_27769);
nand U33428 (N_33428,N_24675,N_29812);
and U33429 (N_33429,N_21374,N_28126);
and U33430 (N_33430,N_29287,N_25975);
or U33431 (N_33431,N_29009,N_27625);
or U33432 (N_33432,N_27245,N_23969);
xor U33433 (N_33433,N_21157,N_24741);
or U33434 (N_33434,N_27437,N_21561);
xnor U33435 (N_33435,N_29640,N_25493);
and U33436 (N_33436,N_28401,N_28069);
nand U33437 (N_33437,N_24778,N_25864);
and U33438 (N_33438,N_23979,N_21409);
and U33439 (N_33439,N_26055,N_24738);
xor U33440 (N_33440,N_23100,N_20367);
or U33441 (N_33441,N_28089,N_25999);
and U33442 (N_33442,N_21681,N_29803);
or U33443 (N_33443,N_20535,N_25677);
and U33444 (N_33444,N_28887,N_29383);
xnor U33445 (N_33445,N_29620,N_22558);
nand U33446 (N_33446,N_24867,N_29836);
nor U33447 (N_33447,N_25687,N_26122);
xnor U33448 (N_33448,N_20524,N_25287);
nor U33449 (N_33449,N_28019,N_26132);
and U33450 (N_33450,N_27574,N_29923);
nor U33451 (N_33451,N_25990,N_23425);
nand U33452 (N_33452,N_24389,N_24220);
nand U33453 (N_33453,N_20955,N_25581);
nand U33454 (N_33454,N_27079,N_20077);
or U33455 (N_33455,N_29986,N_25738);
xor U33456 (N_33456,N_24945,N_27314);
nor U33457 (N_33457,N_27796,N_21060);
nand U33458 (N_33458,N_28949,N_28018);
nand U33459 (N_33459,N_29669,N_24580);
nand U33460 (N_33460,N_27547,N_21770);
nand U33461 (N_33461,N_23890,N_28704);
nor U33462 (N_33462,N_22667,N_29177);
or U33463 (N_33463,N_25466,N_27647);
or U33464 (N_33464,N_21774,N_24412);
xnor U33465 (N_33465,N_27944,N_20662);
xnor U33466 (N_33466,N_27771,N_21402);
xnor U33467 (N_33467,N_26400,N_26744);
or U33468 (N_33468,N_20853,N_27471);
xor U33469 (N_33469,N_23410,N_21176);
xor U33470 (N_33470,N_29858,N_26417);
xnor U33471 (N_33471,N_25580,N_26888);
and U33472 (N_33472,N_27823,N_23765);
and U33473 (N_33473,N_25394,N_28826);
nor U33474 (N_33474,N_29420,N_29404);
and U33475 (N_33475,N_23691,N_26195);
and U33476 (N_33476,N_22054,N_21067);
nor U33477 (N_33477,N_28902,N_29487);
nor U33478 (N_33478,N_25693,N_25298);
xor U33479 (N_33479,N_21958,N_27063);
nand U33480 (N_33480,N_22874,N_22609);
xnor U33481 (N_33481,N_20555,N_26915);
xor U33482 (N_33482,N_25096,N_25226);
and U33483 (N_33483,N_21066,N_20389);
or U33484 (N_33484,N_20683,N_24552);
or U33485 (N_33485,N_27664,N_23920);
xnor U33486 (N_33486,N_23025,N_24289);
or U33487 (N_33487,N_23486,N_20977);
and U33488 (N_33488,N_27374,N_24571);
or U33489 (N_33489,N_27531,N_28119);
or U33490 (N_33490,N_29331,N_20447);
nor U33491 (N_33491,N_27793,N_20253);
xnor U33492 (N_33492,N_23857,N_28416);
nand U33493 (N_33493,N_28862,N_28802);
or U33494 (N_33494,N_20257,N_23376);
nor U33495 (N_33495,N_21480,N_28922);
xnor U33496 (N_33496,N_20965,N_23901);
and U33497 (N_33497,N_22864,N_25131);
xor U33498 (N_33498,N_29650,N_20577);
xnor U33499 (N_33499,N_29152,N_29283);
xnor U33500 (N_33500,N_22063,N_20247);
nor U33501 (N_33501,N_23437,N_22296);
xnor U33502 (N_33502,N_27673,N_21170);
and U33503 (N_33503,N_21734,N_24535);
and U33504 (N_33504,N_25711,N_23488);
xor U33505 (N_33505,N_23013,N_27335);
or U33506 (N_33506,N_27161,N_27864);
nor U33507 (N_33507,N_23191,N_26812);
xnor U33508 (N_33508,N_24032,N_25217);
and U33509 (N_33509,N_20736,N_27145);
and U33510 (N_33510,N_22526,N_22026);
nand U33511 (N_33511,N_28302,N_24139);
xor U33512 (N_33512,N_24634,N_27158);
xor U33513 (N_33513,N_28248,N_21647);
xnor U33514 (N_33514,N_27438,N_24337);
and U33515 (N_33515,N_29028,N_21701);
or U33516 (N_33516,N_26371,N_20072);
nor U33517 (N_33517,N_28584,N_28757);
xor U33518 (N_33518,N_20914,N_23152);
and U33519 (N_33519,N_27058,N_22451);
xor U33520 (N_33520,N_23741,N_21154);
and U33521 (N_33521,N_20810,N_23443);
nor U33522 (N_33522,N_21585,N_20550);
or U33523 (N_33523,N_22973,N_22478);
or U33524 (N_33524,N_21775,N_25803);
nor U33525 (N_33525,N_26304,N_26859);
nand U33526 (N_33526,N_21206,N_28679);
nand U33527 (N_33527,N_24248,N_24323);
nand U33528 (N_33528,N_24235,N_23805);
xnor U33529 (N_33529,N_21243,N_29834);
and U33530 (N_33530,N_20710,N_26048);
xor U33531 (N_33531,N_24626,N_28364);
nor U33532 (N_33532,N_23029,N_29395);
and U33533 (N_33533,N_28300,N_23298);
xnor U33534 (N_33534,N_24177,N_23866);
or U33535 (N_33535,N_29957,N_28852);
nand U33536 (N_33536,N_26930,N_20027);
nor U33537 (N_33537,N_24402,N_27588);
nand U33538 (N_33538,N_23962,N_20855);
nor U33539 (N_33539,N_24530,N_28594);
and U33540 (N_33540,N_25270,N_24868);
nand U33541 (N_33541,N_27083,N_25740);
and U33542 (N_33542,N_26824,N_20350);
nor U33543 (N_33543,N_25804,N_25187);
nor U33544 (N_33544,N_20960,N_22801);
nor U33545 (N_33545,N_26754,N_22141);
nor U33546 (N_33546,N_28899,N_22454);
xnor U33547 (N_33547,N_24810,N_20435);
and U33548 (N_33548,N_23455,N_23987);
nand U33549 (N_33549,N_28898,N_23147);
and U33550 (N_33550,N_24100,N_25802);
and U33551 (N_33551,N_23209,N_21438);
or U33552 (N_33552,N_23853,N_28199);
xnor U33553 (N_33553,N_26759,N_27284);
and U33554 (N_33554,N_25775,N_28507);
and U33555 (N_33555,N_22363,N_27011);
nand U33556 (N_33556,N_21436,N_22227);
and U33557 (N_33557,N_20275,N_24971);
nor U33558 (N_33558,N_22737,N_22421);
nor U33559 (N_33559,N_21008,N_29222);
or U33560 (N_33560,N_22260,N_21320);
nor U33561 (N_33561,N_24781,N_28274);
xor U33562 (N_33562,N_25475,N_28860);
xnor U33563 (N_33563,N_25646,N_23337);
nand U33564 (N_33564,N_21423,N_28191);
nor U33565 (N_33565,N_26807,N_29394);
nor U33566 (N_33566,N_27261,N_25489);
nand U33567 (N_33567,N_20992,N_27405);
nor U33568 (N_33568,N_29407,N_22266);
or U33569 (N_33569,N_29133,N_24757);
nor U33570 (N_33570,N_23295,N_22740);
or U33571 (N_33571,N_28901,N_29811);
xnor U33572 (N_33572,N_21764,N_27737);
and U33573 (N_33573,N_28996,N_22294);
nor U33574 (N_33574,N_29681,N_21826);
nand U33575 (N_33575,N_29255,N_28404);
nor U33576 (N_33576,N_25695,N_28753);
nand U33577 (N_33577,N_21139,N_25090);
nand U33578 (N_33578,N_24101,N_20206);
and U33579 (N_33579,N_27779,N_24880);
nor U33580 (N_33580,N_22279,N_21867);
and U33581 (N_33581,N_28617,N_27287);
nand U33582 (N_33582,N_29704,N_25190);
or U33583 (N_33583,N_29524,N_27785);
nand U33584 (N_33584,N_27139,N_22087);
nand U33585 (N_33585,N_22270,N_29611);
xor U33586 (N_33586,N_20365,N_25149);
nor U33587 (N_33587,N_22872,N_25558);
nand U33588 (N_33588,N_27996,N_24460);
xnor U33589 (N_33589,N_26276,N_25053);
nand U33590 (N_33590,N_26197,N_25101);
or U33591 (N_33591,N_22877,N_22588);
and U33592 (N_33592,N_20480,N_26831);
nand U33593 (N_33593,N_20387,N_29850);
and U33594 (N_33594,N_20668,N_27465);
and U33595 (N_33595,N_21389,N_27190);
xnor U33596 (N_33596,N_22806,N_29062);
and U33597 (N_33597,N_27863,N_28821);
nor U33598 (N_33598,N_23303,N_28837);
xnor U33599 (N_33599,N_23672,N_21735);
nor U33600 (N_33600,N_26554,N_26413);
or U33601 (N_33601,N_24155,N_28924);
or U33602 (N_33602,N_22819,N_22187);
xor U33603 (N_33603,N_24007,N_26150);
nor U33604 (N_33604,N_24611,N_21788);
and U33605 (N_33605,N_21153,N_29890);
nor U33606 (N_33606,N_20811,N_29001);
nand U33607 (N_33607,N_21013,N_24133);
nand U33608 (N_33608,N_21492,N_23619);
and U33609 (N_33609,N_28330,N_28059);
and U33610 (N_33610,N_24627,N_22922);
nand U33611 (N_33611,N_29021,N_28148);
nor U33612 (N_33612,N_23351,N_24219);
and U33613 (N_33613,N_22917,N_26741);
and U33614 (N_33614,N_23692,N_20306);
and U33615 (N_33615,N_26303,N_29943);
xor U33616 (N_33616,N_26723,N_28450);
and U33617 (N_33617,N_21487,N_24292);
xnor U33618 (N_33618,N_27391,N_20370);
xnor U33619 (N_33619,N_21040,N_21789);
or U33620 (N_33620,N_26922,N_23577);
xor U33621 (N_33621,N_24203,N_21317);
nand U33622 (N_33622,N_21281,N_23084);
nand U33623 (N_33623,N_27055,N_28706);
xnor U33624 (N_33624,N_24587,N_22236);
or U33625 (N_33625,N_29616,N_20162);
nor U33626 (N_33626,N_27848,N_21329);
xnor U33627 (N_33627,N_24392,N_21321);
nand U33628 (N_33628,N_29054,N_26911);
or U33629 (N_33629,N_28520,N_25816);
or U33630 (N_33630,N_28722,N_29946);
nor U33631 (N_33631,N_26718,N_26176);
and U33632 (N_33632,N_24480,N_20858);
and U33633 (N_33633,N_20161,N_21367);
nand U33634 (N_33634,N_25447,N_29049);
xor U33635 (N_33635,N_23181,N_21779);
and U33636 (N_33636,N_23226,N_20667);
xnor U33637 (N_33637,N_24735,N_26528);
xor U33638 (N_33638,N_26107,N_29688);
nor U33639 (N_33639,N_23424,N_26430);
xor U33640 (N_33640,N_24005,N_21085);
nand U33641 (N_33641,N_26458,N_20057);
and U33642 (N_33642,N_22450,N_29711);
xnor U33643 (N_33643,N_29522,N_24030);
nand U33644 (N_33644,N_23193,N_24257);
nand U33645 (N_33645,N_22010,N_22427);
nor U33646 (N_33646,N_20771,N_21512);
and U33647 (N_33647,N_23990,N_25094);
or U33648 (N_33648,N_22207,N_25467);
nand U33649 (N_33649,N_28551,N_26090);
xor U33650 (N_33650,N_27336,N_22310);
nand U33651 (N_33651,N_24307,N_20336);
or U33652 (N_33652,N_26969,N_23044);
xor U33653 (N_33653,N_26950,N_20564);
and U33654 (N_33654,N_24516,N_24429);
nand U33655 (N_33655,N_22972,N_25992);
xnor U33656 (N_33656,N_27770,N_23187);
xnor U33657 (N_33657,N_24072,N_25389);
nand U33658 (N_33658,N_21285,N_22532);
and U33659 (N_33659,N_23211,N_24950);
nor U33660 (N_33660,N_25969,N_28378);
and U33661 (N_33661,N_27050,N_27784);
and U33662 (N_33662,N_27783,N_20135);
xnor U33663 (N_33663,N_22557,N_21548);
or U33664 (N_33664,N_29969,N_23050);
nand U33665 (N_33665,N_20881,N_29899);
or U33666 (N_33666,N_21730,N_21425);
and U33667 (N_33667,N_26802,N_25456);
and U33668 (N_33668,N_25031,N_28699);
or U33669 (N_33669,N_23992,N_23869);
xnor U33670 (N_33670,N_27496,N_27091);
nand U33671 (N_33671,N_27592,N_22482);
or U33672 (N_33672,N_21054,N_27226);
or U33673 (N_33673,N_22831,N_24422);
or U33674 (N_33674,N_24079,N_25789);
nand U33675 (N_33675,N_21940,N_25583);
nor U33676 (N_33676,N_25860,N_27325);
xnor U33677 (N_33677,N_26214,N_26247);
nor U33678 (N_33678,N_20741,N_27143);
xnor U33679 (N_33679,N_29922,N_29003);
xnor U33680 (N_33680,N_24595,N_22070);
nor U33681 (N_33681,N_22142,N_29950);
nand U33682 (N_33682,N_24775,N_23418);
or U33683 (N_33683,N_23875,N_20594);
or U33684 (N_33684,N_22047,N_25869);
or U33685 (N_33685,N_25241,N_28304);
nand U33686 (N_33686,N_21142,N_29154);
nor U33687 (N_33687,N_21108,N_27474);
and U33688 (N_33688,N_20196,N_22347);
nand U33689 (N_33689,N_28077,N_23163);
and U33690 (N_33690,N_28589,N_26800);
nand U33691 (N_33691,N_25852,N_26137);
nand U33692 (N_33692,N_20138,N_27582);
nor U33693 (N_33693,N_21753,N_23545);
xor U33694 (N_33694,N_20982,N_25904);
and U33695 (N_33695,N_29499,N_22513);
xnor U33696 (N_33696,N_22002,N_29878);
xor U33697 (N_33697,N_27186,N_29315);
nor U33698 (N_33698,N_24499,N_20944);
nor U33699 (N_33699,N_29968,N_29058);
or U33700 (N_33700,N_28540,N_25260);
xnor U33701 (N_33701,N_27569,N_21283);
nand U33702 (N_33702,N_26941,N_28649);
nand U33703 (N_33703,N_24878,N_25200);
or U33704 (N_33704,N_25454,N_22090);
xor U33705 (N_33705,N_29291,N_23009);
nand U33706 (N_33706,N_25176,N_23568);
nand U33707 (N_33707,N_20317,N_22368);
nor U33708 (N_33708,N_26295,N_23301);
nor U33709 (N_33709,N_24195,N_29415);
or U33710 (N_33710,N_24173,N_22838);
and U33711 (N_33711,N_28392,N_29187);
and U33712 (N_33712,N_24384,N_26408);
xor U33713 (N_33713,N_28303,N_25033);
nor U33714 (N_33714,N_28593,N_22617);
or U33715 (N_33715,N_21797,N_22139);
or U33716 (N_33716,N_23735,N_20910);
or U33717 (N_33717,N_23332,N_28705);
xor U33718 (N_33718,N_27774,N_25010);
nand U33719 (N_33719,N_20151,N_20319);
xnor U33720 (N_33720,N_20856,N_23730);
xor U33721 (N_33721,N_26001,N_24425);
and U33722 (N_33722,N_28720,N_25582);
nor U33723 (N_33723,N_22411,N_24169);
or U33724 (N_33724,N_27728,N_27061);
xor U33725 (N_33725,N_26747,N_20676);
and U33726 (N_33726,N_21633,N_21503);
nor U33727 (N_33727,N_29165,N_23135);
and U33728 (N_33728,N_28422,N_25025);
xor U33729 (N_33729,N_21268,N_29155);
nor U33730 (N_33730,N_23665,N_23696);
xor U33731 (N_33731,N_26960,N_20334);
or U33732 (N_33732,N_28976,N_22402);
xnor U33733 (N_33733,N_22275,N_23098);
nor U33734 (N_33734,N_24962,N_21369);
or U33735 (N_33735,N_29076,N_24283);
or U33736 (N_33736,N_27136,N_21493);
and U33737 (N_33737,N_26003,N_25519);
xnor U33738 (N_33738,N_21868,N_28319);
nor U33739 (N_33739,N_22993,N_21076);
nand U33740 (N_33740,N_22330,N_27949);
and U33741 (N_33741,N_26981,N_22326);
and U33742 (N_33742,N_25956,N_27978);
and U33743 (N_33743,N_25822,N_24922);
and U33744 (N_33744,N_22797,N_26738);
nand U33745 (N_33745,N_23416,N_21693);
or U33746 (N_33746,N_22641,N_26889);
and U33747 (N_33747,N_25038,N_24615);
or U33748 (N_33748,N_22898,N_28485);
nor U33749 (N_33749,N_21333,N_28051);
or U33750 (N_33750,N_25843,N_25230);
or U33751 (N_33751,N_20357,N_25940);
and U33752 (N_33752,N_23654,N_25896);
nand U33753 (N_33753,N_21778,N_28260);
nor U33754 (N_33754,N_22718,N_25146);
xnor U33755 (N_33755,N_21421,N_26832);
nand U33756 (N_33756,N_20840,N_24540);
nand U33757 (N_33757,N_23548,N_28146);
and U33758 (N_33758,N_27648,N_24659);
nor U33759 (N_33759,N_26796,N_24094);
xor U33760 (N_33760,N_24205,N_28249);
or U33761 (N_33761,N_28457,N_24617);
nor U33762 (N_33762,N_21888,N_21644);
and U33763 (N_33763,N_28962,N_20269);
or U33764 (N_33764,N_24107,N_21430);
or U33765 (N_33765,N_28668,N_22109);
and U33766 (N_33766,N_29202,N_29701);
nand U33767 (N_33767,N_26442,N_25905);
nor U33768 (N_33768,N_23507,N_25280);
and U33769 (N_33769,N_20805,N_29626);
or U33770 (N_33770,N_29216,N_22420);
or U33771 (N_33771,N_26080,N_23970);
nor U33772 (N_33772,N_21497,N_25799);
nor U33773 (N_33773,N_26666,N_21432);
nand U33774 (N_33774,N_28571,N_29989);
nor U33775 (N_33775,N_27762,N_29104);
nand U33776 (N_33776,N_20228,N_26976);
xor U33777 (N_33777,N_21125,N_23062);
or U33778 (N_33778,N_24981,N_26616);
and U33779 (N_33779,N_20658,N_27142);
xor U33780 (N_33780,N_23825,N_28329);
and U33781 (N_33781,N_29382,N_20091);
nor U33782 (N_33782,N_22325,N_29949);
nor U33783 (N_33783,N_23961,N_28179);
or U33784 (N_33784,N_25535,N_23110);
or U33785 (N_33785,N_22687,N_26478);
nand U33786 (N_33786,N_26477,N_20050);
xnor U33787 (N_33787,N_27877,N_24418);
xnor U33788 (N_33788,N_22094,N_27099);
xnor U33789 (N_33789,N_29953,N_26380);
or U33790 (N_33790,N_28185,N_29789);
or U33791 (N_33791,N_25589,N_24349);
or U33792 (N_33792,N_21850,N_29702);
xor U33793 (N_33793,N_23094,N_26440);
and U33794 (N_33794,N_22167,N_25515);
and U33795 (N_33795,N_29713,N_29966);
and U33796 (N_33796,N_27431,N_25810);
or U33797 (N_33797,N_20147,N_28716);
or U33798 (N_33798,N_26410,N_27867);
and U33799 (N_33799,N_23759,N_20843);
nand U33800 (N_33800,N_25463,N_20274);
nand U33801 (N_33801,N_27202,N_25294);
xor U33802 (N_33802,N_25408,N_24977);
nor U33803 (N_33803,N_21479,N_27656);
nand U33804 (N_33804,N_22576,N_20609);
nand U33805 (N_33805,N_29738,N_28343);
nor U33806 (N_33806,N_27620,N_21578);
xnor U33807 (N_33807,N_22406,N_27881);
nand U33808 (N_33808,N_22889,N_22101);
or U33809 (N_33809,N_23959,N_25201);
xnor U33810 (N_33810,N_22646,N_21923);
xor U33811 (N_33811,N_24383,N_21207);
xnor U33812 (N_33812,N_20197,N_21593);
or U33813 (N_33813,N_29025,N_28419);
nand U33814 (N_33814,N_29380,N_29665);
nor U33815 (N_33815,N_23534,N_23040);
nand U33816 (N_33816,N_23814,N_22058);
nand U33817 (N_33817,N_27795,N_27310);
xnor U33818 (N_33818,N_26680,N_29302);
nand U33819 (N_33819,N_20723,N_25009);
xnor U33820 (N_33820,N_22474,N_28955);
xnor U33821 (N_33821,N_29780,N_23131);
nand U33822 (N_33822,N_24942,N_22791);
xnor U33823 (N_33823,N_25946,N_20803);
and U33824 (N_33824,N_23859,N_26692);
nor U33825 (N_33825,N_20427,N_21133);
and U33826 (N_33826,N_21200,N_26735);
nor U33827 (N_33827,N_27826,N_23249);
nor U33828 (N_33828,N_21408,N_20687);
xnor U33829 (N_33829,N_23804,N_29387);
or U33830 (N_33830,N_27894,N_27695);
or U33831 (N_33831,N_25927,N_22803);
nor U33832 (N_33832,N_23489,N_23317);
or U33833 (N_33833,N_25781,N_27359);
xnor U33834 (N_33834,N_22763,N_23058);
nand U33835 (N_33835,N_24172,N_22550);
xor U33836 (N_33836,N_20457,N_20649);
or U33837 (N_33837,N_24504,N_25914);
and U33838 (N_33838,N_24650,N_27681);
xor U33839 (N_33839,N_23008,N_20630);
nand U33840 (N_33840,N_27178,N_29856);
and U33841 (N_33841,N_27102,N_21210);
and U33842 (N_33842,N_20761,N_27197);
or U33843 (N_33843,N_24982,N_25897);
and U33844 (N_33844,N_28948,N_20681);
nand U33845 (N_33845,N_23413,N_24103);
or U33846 (N_33846,N_27448,N_29176);
and U33847 (N_33847,N_29610,N_24042);
or U33848 (N_33848,N_28091,N_25565);
xnor U33849 (N_33849,N_22770,N_21612);
nor U33850 (N_33850,N_26908,N_29903);
and U33851 (N_33851,N_21295,N_27637);
xor U33852 (N_33852,N_26884,N_21636);
or U33853 (N_33853,N_26509,N_21091);
nor U33854 (N_33854,N_21449,N_21446);
xor U33855 (N_33855,N_20416,N_23477);
nor U33856 (N_33856,N_25228,N_22684);
and U33857 (N_33857,N_26280,N_27982);
and U33858 (N_33858,N_23266,N_27653);
and U33859 (N_33859,N_25378,N_26862);
xor U33860 (N_33860,N_20528,N_28878);
nor U33861 (N_33861,N_21494,N_24061);
or U33862 (N_33862,N_21674,N_29521);
xor U33863 (N_33863,N_26775,N_25625);
nand U33864 (N_33864,N_26242,N_21123);
nand U33865 (N_33865,N_27389,N_25140);
xor U33866 (N_33866,N_24021,N_29670);
nor U33867 (N_33867,N_25477,N_26158);
nor U33868 (N_33868,N_24241,N_23339);
nand U33869 (N_33869,N_26345,N_24222);
or U33870 (N_33870,N_23749,N_23219);
xnor U33871 (N_33871,N_24618,N_29428);
or U33872 (N_33872,N_24645,N_27539);
xor U33873 (N_33873,N_22086,N_25065);
xor U33874 (N_33874,N_24083,N_21801);
nand U33875 (N_33875,N_26896,N_28547);
nand U33876 (N_33876,N_23980,N_25543);
xor U33877 (N_33877,N_29603,N_27256);
xnor U33878 (N_33878,N_26562,N_27865);
nor U33879 (N_33879,N_26130,N_28682);
xnor U33880 (N_33880,N_29485,N_29839);
or U33881 (N_33881,N_28386,N_26337);
or U33882 (N_33882,N_28098,N_22986);
or U33883 (N_33883,N_29714,N_26553);
nor U33884 (N_33884,N_26325,N_25387);
nor U33885 (N_33885,N_25252,N_27844);
and U33886 (N_33886,N_26194,N_25078);
and U33887 (N_33887,N_26793,N_23204);
or U33888 (N_33888,N_24162,N_22190);
or U33889 (N_33889,N_23223,N_24605);
or U33890 (N_33890,N_26633,N_21358);
nor U33891 (N_33891,N_29079,N_22351);
nor U33892 (N_33892,N_24284,N_24817);
or U33893 (N_33893,N_22067,N_23282);
or U33894 (N_33894,N_29584,N_29052);
or U33895 (N_33895,N_25125,N_23818);
xnor U33896 (N_33896,N_20756,N_22314);
or U33897 (N_33897,N_25704,N_23637);
nand U33898 (N_33898,N_29233,N_26126);
xnor U33899 (N_33899,N_25995,N_20386);
xor U33900 (N_33900,N_21444,N_22319);
or U33901 (N_33901,N_25951,N_21498);
nor U33902 (N_33902,N_28425,N_22390);
and U33903 (N_33903,N_25892,N_25942);
nand U33904 (N_33904,N_25573,N_21403);
nand U33905 (N_33905,N_23525,N_29734);
and U33906 (N_33906,N_26459,N_22253);
nor U33907 (N_33907,N_26731,N_20251);
nand U33908 (N_33908,N_21391,N_21686);
xnor U33909 (N_33909,N_21700,N_25039);
or U33910 (N_33910,N_20769,N_24160);
xor U33911 (N_33911,N_21557,N_22539);
xor U33912 (N_33912,N_21099,N_24602);
nor U33913 (N_33913,N_24918,N_20857);
and U33914 (N_33914,N_21244,N_24712);
and U33915 (N_33915,N_25006,N_22468);
xnor U33916 (N_33916,N_20489,N_22858);
xnor U33917 (N_33917,N_24701,N_23268);
xor U33918 (N_33918,N_27666,N_25379);
nand U33919 (N_33919,N_22285,N_22258);
or U33920 (N_33920,N_20491,N_21900);
or U33921 (N_33921,N_22860,N_22153);
nor U33922 (N_33922,N_21410,N_26058);
and U33923 (N_33923,N_22554,N_24622);
xnor U33924 (N_33924,N_22117,N_20926);
xnor U33925 (N_33925,N_22521,N_22915);
nor U33926 (N_33926,N_22467,N_23469);
and U33927 (N_33927,N_23368,N_29896);
and U33928 (N_33928,N_27812,N_20498);
xnor U33929 (N_33929,N_28264,N_28503);
or U33930 (N_33930,N_21883,N_29442);
and U33931 (N_33931,N_27879,N_27004);
nand U33932 (N_33932,N_27181,N_24456);
nand U33933 (N_33933,N_20223,N_28514);
nor U33934 (N_33934,N_25313,N_20203);
or U33935 (N_33935,N_21323,N_21322);
xnor U33936 (N_33936,N_20513,N_27651);
xnor U33937 (N_33937,N_27644,N_21596);
nand U33938 (N_33938,N_23059,N_29221);
or U33939 (N_33939,N_27205,N_22663);
and U33940 (N_33940,N_27481,N_23553);
xnor U33941 (N_33941,N_20006,N_27503);
or U33942 (N_33942,N_28771,N_24204);
or U33943 (N_33943,N_24012,N_27974);
or U33944 (N_33944,N_23965,N_26691);
xnor U33945 (N_33945,N_27658,N_27563);
xor U33946 (N_33946,N_20024,N_25220);
nor U33947 (N_33947,N_22533,N_29260);
and U33948 (N_33948,N_28480,N_29027);
or U33949 (N_33949,N_25299,N_29748);
nor U33950 (N_33950,N_29520,N_25088);
nand U33951 (N_33951,N_23727,N_24665);
and U33952 (N_33952,N_23166,N_27164);
and U33953 (N_33953,N_26071,N_23615);
nor U33954 (N_33954,N_25754,N_27343);
or U33955 (N_33955,N_29036,N_23452);
or U33956 (N_33956,N_27654,N_28049);
and U33957 (N_33957,N_27094,N_21910);
and U33958 (N_33958,N_21413,N_28859);
xor U33959 (N_33959,N_25259,N_21375);
and U33960 (N_33960,N_25441,N_28299);
xnor U33961 (N_33961,N_20496,N_26782);
and U33962 (N_33962,N_20391,N_23955);
xnor U33963 (N_33963,N_28078,N_27565);
and U33964 (N_33964,N_24996,N_22738);
or U33965 (N_33965,N_25392,N_26360);
nor U33966 (N_33966,N_21300,N_26627);
nand U33967 (N_33967,N_22857,N_28373);
or U33968 (N_33968,N_20182,N_21642);
nand U33969 (N_33969,N_22822,N_20342);
nand U33970 (N_33970,N_23738,N_27432);
or U33971 (N_33971,N_29468,N_22556);
and U33972 (N_33972,N_26502,N_26386);
nor U33973 (N_33973,N_27403,N_22247);
nor U33974 (N_33974,N_20399,N_24720);
or U33975 (N_33975,N_23442,N_28407);
nand U33976 (N_33976,N_21460,N_21262);
nor U33977 (N_33977,N_25141,N_27856);
or U33978 (N_33978,N_20329,N_22542);
or U33979 (N_33979,N_22555,N_24033);
and U33980 (N_33980,N_21893,N_22739);
and U33981 (N_33981,N_28309,N_24896);
and U33982 (N_33982,N_23561,N_21306);
or U33983 (N_33983,N_26473,N_23287);
nor U33984 (N_33984,N_28601,N_27425);
or U33985 (N_33985,N_27660,N_24747);
and U33986 (N_33986,N_25508,N_23758);
and U33987 (N_33987,N_24329,N_28281);
or U33988 (N_33988,N_26402,N_28291);
or U33989 (N_33989,N_28224,N_20807);
xor U33990 (N_33990,N_27953,N_27589);
and U33991 (N_33991,N_29798,N_21650);
or U33992 (N_33992,N_26513,N_28813);
xor U33993 (N_33993,N_23083,N_26329);
nor U33994 (N_33994,N_29643,N_20549);
nor U33995 (N_33995,N_22990,N_22149);
and U33996 (N_33996,N_26909,N_24486);
and U33997 (N_33997,N_23911,N_21877);
and U33998 (N_33998,N_23068,N_27151);
xor U33999 (N_33999,N_28764,N_20647);
or U34000 (N_34000,N_21209,N_26756);
nand U34001 (N_34001,N_24485,N_24785);
and U34002 (N_34002,N_29976,N_27672);
xnor U34003 (N_34003,N_27243,N_22439);
xor U34004 (N_34004,N_24256,N_29432);
or U34005 (N_34005,N_21427,N_26801);
nor U34006 (N_34006,N_29034,N_28489);
and U34007 (N_34007,N_22569,N_29375);
nand U34008 (N_34008,N_21383,N_27962);
nor U34009 (N_34009,N_26629,N_21226);
and U34010 (N_34010,N_26883,N_25482);
nor U34011 (N_34011,N_26737,N_21749);
xor U34012 (N_34012,N_23134,N_23611);
nand U34013 (N_34013,N_20250,N_25367);
or U34014 (N_34014,N_22886,N_26693);
nand U34015 (N_34015,N_22377,N_24899);
nand U34016 (N_34016,N_27467,N_26839);
nand U34017 (N_34017,N_29581,N_27624);
or U34018 (N_34018,N_23041,N_22195);
or U34019 (N_34019,N_23167,N_23347);
nand U34020 (N_34020,N_26394,N_27258);
nor U34021 (N_34021,N_22882,N_28083);
and U34022 (N_34022,N_29385,N_29364);
and U34023 (N_34023,N_28289,N_29275);
nand U34024 (N_34024,N_21812,N_27305);
xnor U34025 (N_34025,N_21732,N_22068);
and U34026 (N_34026,N_26149,N_28001);
and U34027 (N_34027,N_20905,N_28211);
and U34028 (N_34028,N_28483,N_24385);
xnor U34029 (N_34029,N_22472,N_29100);
or U34030 (N_34030,N_22218,N_20912);
xnor U34031 (N_34031,N_22934,N_28909);
xor U34032 (N_34032,N_22691,N_25955);
nor U34033 (N_34033,N_22189,N_26029);
or U34034 (N_34034,N_29072,N_23192);
and U34035 (N_34035,N_23649,N_20829);
or U34036 (N_34036,N_20026,N_20548);
and U34037 (N_34037,N_21699,N_21250);
and U34038 (N_34038,N_26115,N_22970);
nand U34039 (N_34039,N_22816,N_21270);
nor U34040 (N_34040,N_20791,N_23074);
nand U34041 (N_34041,N_27693,N_21216);
xnor U34042 (N_34042,N_23538,N_27602);
and U34043 (N_34043,N_20879,N_22516);
xor U34044 (N_34044,N_23902,N_25538);
nor U34045 (N_34045,N_27246,N_27494);
nor U34046 (N_34046,N_23821,N_28995);
xor U34047 (N_34047,N_20031,N_21426);
nand U34048 (N_34048,N_28159,N_22118);
nor U34049 (N_34049,N_20436,N_24732);
xor U34050 (N_34050,N_21124,N_25265);
nand U34051 (N_34051,N_29306,N_24845);
nor U34052 (N_34052,N_21565,N_21156);
nor U34053 (N_34053,N_29412,N_27916);
nand U34054 (N_34054,N_20917,N_29927);
and U34055 (N_34055,N_23372,N_28176);
xnor U34056 (N_34056,N_25509,N_21105);
or U34057 (N_34057,N_29035,N_27564);
or U34058 (N_34058,N_24117,N_24740);
and U34059 (N_34059,N_28093,N_28327);
and U34060 (N_34060,N_20801,N_22460);
and U34061 (N_34061,N_23151,N_28708);
or U34062 (N_34062,N_24410,N_28536);
nor U34063 (N_34063,N_23127,N_21556);
nor U34064 (N_34064,N_26173,N_28861);
nand U34065 (N_34065,N_29486,N_20004);
or U34066 (N_34066,N_23829,N_24132);
nand U34067 (N_34067,N_20989,N_24590);
xor U34068 (N_34068,N_29107,N_27274);
xor U34069 (N_34069,N_20239,N_29606);
nor U34070 (N_34070,N_27464,N_25091);
nor U34071 (N_34071,N_27671,N_29945);
nor U34072 (N_34072,N_22171,N_22416);
nand U34073 (N_34073,N_25675,N_22436);
nor U34074 (N_34074,N_23748,N_24944);
or U34075 (N_34075,N_21106,N_27380);
and U34076 (N_34076,N_28894,N_25142);
xnor U34077 (N_34077,N_25288,N_27182);
or U34078 (N_34078,N_21102,N_24110);
or U34079 (N_34079,N_21372,N_25666);
and U34080 (N_34080,N_29252,N_22660);
xnor U34081 (N_34081,N_21962,N_23265);
nor U34082 (N_34082,N_26364,N_24737);
nand U34083 (N_34083,N_21282,N_22287);
nor U34084 (N_34084,N_29303,N_24439);
nand U34085 (N_34085,N_26849,N_28908);
nor U34086 (N_34086,N_28553,N_20816);
or U34087 (N_34087,N_26405,N_20830);
nor U34088 (N_34088,N_29169,N_24734);
or U34089 (N_34089,N_21371,N_26023);
or U34090 (N_34090,N_25449,N_23346);
nand U34091 (N_34091,N_24601,N_21316);
and U34092 (N_34092,N_24387,N_28846);
nand U34093 (N_34093,N_25853,N_27308);
nand U34094 (N_34094,N_20631,N_28334);
and U34095 (N_34095,N_20281,N_22987);
or U34096 (N_34096,N_27282,N_26900);
nand U34097 (N_34097,N_25989,N_29491);
nor U34098 (N_34098,N_27388,N_22709);
xor U34099 (N_34099,N_23584,N_29464);
xor U34100 (N_34100,N_29241,N_29637);
and U34101 (N_34101,N_25961,N_21785);
nand U34102 (N_34102,N_23179,N_27341);
xnor U34103 (N_34103,N_25358,N_23617);
or U34104 (N_34104,N_29959,N_23422);
and U34105 (N_34105,N_23153,N_22974);
xnor U34106 (N_34106,N_21654,N_28057);
or U34107 (N_34107,N_25291,N_27665);
xor U34108 (N_34108,N_29632,N_23230);
nand U34109 (N_34109,N_22963,N_25645);
nand U34110 (N_34110,N_24849,N_22276);
xor U34111 (N_34111,N_20422,N_24876);
and U34112 (N_34112,N_28671,N_22949);
xor U34113 (N_34113,N_23760,N_21339);
or U34114 (N_34114,N_20034,N_29320);
and U34115 (N_34115,N_28071,N_22711);
nand U34116 (N_34116,N_24840,N_20124);
and U34117 (N_34117,N_25650,N_21586);
xor U34118 (N_34118,N_20878,N_20990);
nand U34119 (N_34119,N_21234,N_24931);
or U34120 (N_34120,N_21762,N_23096);
or U34121 (N_34121,N_20899,N_28979);
nor U34122 (N_34122,N_25873,N_20718);
or U34123 (N_34123,N_26587,N_27396);
xor U34124 (N_34124,N_28731,N_26255);
and U34125 (N_34125,N_25902,N_24984);
or U34126 (N_34126,N_28400,N_26823);
nand U34127 (N_34127,N_21806,N_21242);
xor U34128 (N_34128,N_23929,N_23133);
nor U34129 (N_34129,N_25172,N_23508);
and U34130 (N_34130,N_21011,N_26770);
or U34131 (N_34131,N_22173,N_21750);
nor U34132 (N_34132,N_29285,N_24157);
and U34133 (N_34133,N_29088,N_27421);
and U34134 (N_34134,N_23957,N_26275);
or U34135 (N_34135,N_27277,N_20519);
nor U34136 (N_34136,N_29063,N_20242);
xor U34137 (N_34137,N_25900,N_24895);
or U34138 (N_34138,N_27803,N_20997);
or U34139 (N_34139,N_22265,N_26514);
xor U34140 (N_34140,N_23262,N_22594);
or U34141 (N_34141,N_26563,N_21524);
and U34142 (N_34142,N_24288,N_22920);
and U34143 (N_34143,N_28663,N_29226);
xor U34144 (N_34144,N_29236,N_22127);
or U34145 (N_34145,N_22758,N_27509);
or U34146 (N_34146,N_23850,N_24917);
and U34147 (N_34147,N_23638,N_29608);
and U34148 (N_34148,N_23430,N_26106);
nand U34149 (N_34149,N_24646,N_27447);
nand U34150 (N_34150,N_26983,N_24870);
or U34151 (N_34151,N_26875,N_27880);
xor U34152 (N_34152,N_28056,N_22407);
or U34153 (N_34153,N_25127,N_21336);
nor U34154 (N_34154,N_28206,N_20193);
xnor U34155 (N_34155,N_22444,N_21360);
or U34156 (N_34156,N_22861,N_23812);
xnor U34157 (N_34157,N_29929,N_22686);
nand U34158 (N_34158,N_25832,N_23465);
xor U34159 (N_34159,N_26395,N_23736);
or U34160 (N_34160,N_28608,N_23867);
nor U34161 (N_34161,N_29547,N_26865);
and U34162 (N_34162,N_23734,N_28088);
nor U34163 (N_34163,N_26221,N_28741);
nand U34164 (N_34164,N_24674,N_24446);
or U34165 (N_34165,N_22976,N_29112);
nor U34166 (N_34166,N_24723,N_26177);
nand U34167 (N_34167,N_22222,N_28456);
or U34168 (N_34168,N_23483,N_20232);
xnor U34169 (N_34169,N_23669,N_24800);
nor U34170 (N_34170,N_25794,N_22796);
xor U34171 (N_34171,N_27857,N_23189);
or U34172 (N_34172,N_28621,N_24616);
or U34173 (N_34173,N_21566,N_22191);
and U34174 (N_34174,N_25894,N_21312);
or U34175 (N_34175,N_20740,N_23971);
nor U34176 (N_34176,N_23827,N_20156);
or U34177 (N_34177,N_24600,N_21328);
nor U34178 (N_34178,N_20799,N_23702);
xor U34179 (N_34179,N_24046,N_25979);
nand U34180 (N_34180,N_26816,N_24303);
xor U34181 (N_34181,N_23180,N_29625);
nand U34182 (N_34182,N_26457,N_25533);
xnor U34183 (N_34183,N_27708,N_27087);
nand U34184 (N_34184,N_21833,N_21467);
and U34185 (N_34185,N_20185,N_26804);
xor U34186 (N_34186,N_24935,N_26233);
nand U34187 (N_34187,N_28945,N_20763);
nor U34188 (N_34188,N_26533,N_27719);
nand U34189 (N_34189,N_29146,N_20738);
nand U34190 (N_34190,N_27377,N_23000);
xor U34191 (N_34191,N_20707,N_23091);
nor U34192 (N_34192,N_27313,N_29995);
xor U34193 (N_34193,N_29450,N_20118);
xor U34194 (N_34194,N_21472,N_28209);
nand U34195 (N_34195,N_29430,N_25464);
xnor U34196 (N_34196,N_28116,N_21248);
and U34197 (N_34197,N_28172,N_22150);
nand U34198 (N_34198,N_27610,N_28711);
or U34199 (N_34199,N_27250,N_24879);
or U34200 (N_34200,N_23770,N_23937);
xor U34201 (N_34201,N_22470,N_28317);
nor U34202 (N_34202,N_20045,N_26805);
nor U34203 (N_34203,N_26931,N_27911);
nor U34204 (N_34204,N_24332,N_28306);
xnor U34205 (N_34205,N_28363,N_21134);
and U34206 (N_34206,N_22640,N_25861);
and U34207 (N_34207,N_26740,N_26125);
or U34208 (N_34208,N_26532,N_27073);
nor U34209 (N_34209,N_22916,N_22334);
and U34210 (N_34210,N_26147,N_25385);
xnor U34211 (N_34211,N_26786,N_20766);
nand U34212 (N_34212,N_23648,N_25335);
and U34213 (N_34213,N_23766,N_21481);
and U34214 (N_34214,N_21815,N_21022);
xor U34215 (N_34215,N_27459,N_27412);
xnor U34216 (N_34216,N_27593,N_26855);
xor U34217 (N_34217,N_21884,N_21394);
nor U34218 (N_34218,N_22089,N_25929);
nand U34219 (N_34219,N_23018,N_25547);
nand U34220 (N_34220,N_20314,N_24668);
or U34221 (N_34221,N_29190,N_24999);
xnor U34222 (N_34222,N_22704,N_28305);
xnor U34223 (N_34223,N_28858,N_26893);
nor U34224 (N_34224,N_25345,N_28857);
or U34225 (N_34225,N_21617,N_24872);
nand U34226 (N_34226,N_27977,N_28580);
or U34227 (N_34227,N_29557,N_20568);
nor U34228 (N_34228,N_26389,N_28653);
or U34229 (N_34229,N_20994,N_20411);
nand U34230 (N_34230,N_20603,N_27159);
or U34231 (N_34231,N_24513,N_22186);
xnor U34232 (N_34232,N_28624,N_25681);
nand U34233 (N_34233,N_23002,N_28231);
or U34234 (N_34234,N_23633,N_22992);
nor U34235 (N_34235,N_27233,N_27331);
and U34236 (N_34236,N_26099,N_20680);
nand U34237 (N_34237,N_29362,N_27549);
or U34238 (N_34238,N_22432,N_28595);
and U34239 (N_34239,N_20046,N_27473);
xor U34240 (N_34240,N_22582,N_22907);
and U34241 (N_34241,N_24234,N_26103);
nor U34242 (N_34242,N_25653,N_26707);
or U34243 (N_34243,N_23454,N_26251);
nand U34244 (N_34244,N_27501,N_29279);
or U34245 (N_34245,N_20140,N_25937);
nor U34246 (N_34246,N_28582,N_27641);
or U34247 (N_34247,N_27047,N_20150);
xor U34248 (N_34248,N_27649,N_27747);
and U34249 (N_34249,N_21221,N_21387);
xor U34250 (N_34250,N_21183,N_21078);
nor U34251 (N_34251,N_29866,N_24237);
xor U34252 (N_34252,N_25269,N_26453);
or U34253 (N_34253,N_24010,N_23954);
xnor U34254 (N_34254,N_28451,N_20547);
nand U34255 (N_34255,N_24661,N_28502);
or U34256 (N_34256,N_29330,N_29097);
nor U34257 (N_34257,N_28897,N_22854);
nor U34258 (N_34258,N_23840,N_26841);
nor U34259 (N_34259,N_27113,N_25196);
and U34260 (N_34260,N_23897,N_25459);
and U34261 (N_34261,N_20661,N_20700);
and U34262 (N_34262,N_25346,N_27694);
xor U34263 (N_34263,N_29249,N_26791);
or U34264 (N_34264,N_25570,N_21032);
xor U34265 (N_34265,N_22975,N_26293);
xor U34266 (N_34266,N_24865,N_29337);
nor U34267 (N_34267,N_27012,N_28402);
xor U34268 (N_34268,N_29749,N_28396);
and U34269 (N_34269,N_24642,N_24423);
and U34270 (N_34270,N_21589,N_24582);
and U34271 (N_34271,N_20111,N_28690);
and U34272 (N_34272,N_25811,N_22818);
and U34273 (N_34273,N_24814,N_25079);
and U34274 (N_34274,N_22462,N_28301);
or U34275 (N_34275,N_22962,N_27247);
nor U34276 (N_34276,N_24969,N_25925);
nor U34277 (N_34277,N_25597,N_24911);
and U34278 (N_34278,N_23162,N_26374);
and U34279 (N_34279,N_21803,N_28695);
and U34280 (N_34280,N_24354,N_26928);
xor U34281 (N_34281,N_29733,N_20481);
xor U34282 (N_34282,N_20642,N_21680);
or U34283 (N_34283,N_22383,N_25153);
nor U34284 (N_34284,N_27401,N_21573);
nand U34285 (N_34285,N_29393,N_24238);
nor U34286 (N_34286,N_24363,N_28417);
nor U34287 (N_34287,N_26203,N_27711);
or U34288 (N_34288,N_24022,N_23801);
or U34289 (N_34289,N_23093,N_28002);
nor U34290 (N_34290,N_27984,N_20278);
nor U34291 (N_34291,N_25416,N_20984);
nor U34292 (N_34292,N_22418,N_22254);
nand U34293 (N_34293,N_27262,N_28494);
nor U34294 (N_34294,N_21787,N_27938);
nand U34295 (N_34295,N_28886,N_26542);
nand U34296 (N_34296,N_21304,N_28045);
xnor U34297 (N_34297,N_26006,N_25540);
nand U34298 (N_34298,N_25529,N_29156);
nand U34299 (N_34299,N_24572,N_21457);
nand U34300 (N_34300,N_20079,N_24696);
nor U34301 (N_34301,N_23182,N_21452);
or U34302 (N_34302,N_27507,N_27932);
nor U34303 (N_34303,N_23051,N_25254);
or U34304 (N_34304,N_21148,N_22710);
or U34305 (N_34305,N_29087,N_23433);
xor U34306 (N_34306,N_27578,N_21351);
nor U34307 (N_34307,N_28003,N_21465);
nand U34308 (N_34308,N_27134,N_21708);
nand U34309 (N_34309,N_22065,N_20355);
nand U34310 (N_34310,N_29842,N_28252);
or U34311 (N_34311,N_20615,N_27772);
or U34312 (N_34312,N_27198,N_28674);
and U34313 (N_34313,N_21212,N_26436);
nor U34314 (N_34314,N_29403,N_26170);
and U34315 (N_34315,N_26433,N_24789);
xnor U34316 (N_34316,N_29201,N_21626);
nor U34317 (N_34317,N_27806,N_27525);
nor U34318 (N_34318,N_22181,N_28953);
or U34319 (N_34319,N_26997,N_26223);
xor U34320 (N_34320,N_24522,N_28787);
and U34321 (N_34321,N_25684,N_25050);
or U34322 (N_34322,N_24596,N_23930);
nor U34323 (N_34323,N_24312,N_28267);
nand U34324 (N_34324,N_29580,N_25374);
xor U34325 (N_34325,N_27706,N_20402);
and U34326 (N_34326,N_26768,N_21872);
or U34327 (N_34327,N_20511,N_24667);
xor U34328 (N_34328,N_25179,N_27231);
xor U34329 (N_34329,N_26987,N_29014);
xor U34330 (N_34330,N_23809,N_25166);
xor U34331 (N_34331,N_28342,N_24039);
nand U34332 (N_34332,N_20554,N_25209);
xor U34333 (N_34333,N_25401,N_27150);
nor U34334 (N_34334,N_25746,N_22148);
nand U34335 (N_34335,N_22511,N_20145);
nand U34336 (N_34336,N_29788,N_25840);
or U34337 (N_34337,N_20967,N_22689);
and U34338 (N_34338,N_21059,N_27745);
or U34339 (N_34339,N_29191,N_28458);
or U34340 (N_34340,N_23325,N_21412);
nor U34341 (N_34341,N_20606,N_28058);
nand U34342 (N_34342,N_25945,N_20534);
nor U34343 (N_34343,N_20552,N_23345);
xnor U34344 (N_34344,N_29470,N_28036);
nand U34345 (N_34345,N_22603,N_27584);
nand U34346 (N_34346,N_26589,N_20862);
nor U34347 (N_34347,N_26957,N_24866);
xnor U34348 (N_34348,N_23828,N_28021);
xor U34349 (N_34349,N_25219,N_28190);
nor U34350 (N_34350,N_23676,N_25150);
nor U34351 (N_34351,N_20133,N_27230);
xor U34352 (N_34352,N_28238,N_24921);
and U34353 (N_34353,N_20390,N_26880);
xnor U34354 (N_34354,N_27524,N_22839);
or U34355 (N_34355,N_24001,N_25465);
xor U34356 (N_34356,N_28879,N_24492);
or U34357 (N_34357,N_29313,N_29693);
nor U34358 (N_34358,N_26548,N_22349);
nand U34359 (N_34359,N_22292,N_24762);
nand U34360 (N_34360,N_29921,N_21471);
nor U34361 (N_34361,N_26534,N_22022);
xor U34362 (N_34362,N_22465,N_28464);
xor U34363 (N_34363,N_20155,N_21404);
nor U34364 (N_34364,N_26059,N_26292);
and U34365 (N_34365,N_27285,N_26488);
or U34366 (N_34366,N_23578,N_24523);
xnor U34367 (N_34367,N_24951,N_27688);
nand U34368 (N_34368,N_20070,N_20368);
and U34369 (N_34369,N_28896,N_20328);
and U34370 (N_34370,N_24725,N_28774);
nand U34371 (N_34371,N_26722,N_28197);
nor U34372 (N_34372,N_27692,N_21346);
or U34373 (N_34373,N_25104,N_20706);
nor U34374 (N_34374,N_25691,N_25591);
xnor U34375 (N_34375,N_20970,N_27788);
nand U34376 (N_34376,N_27712,N_24229);
nor U34377 (N_34377,N_25871,N_26222);
nand U34378 (N_34378,N_21537,N_22050);
and U34379 (N_34379,N_27237,N_25048);
and U34380 (N_34380,N_21559,N_25479);
nor U34381 (N_34381,N_22665,N_22031);
nand U34382 (N_34382,N_20908,N_26169);
and U34383 (N_34383,N_28473,N_29539);
and U34384 (N_34384,N_22757,N_29804);
nor U34385 (N_34385,N_21137,N_27395);
nor U34386 (N_34386,N_22512,N_28171);
nand U34387 (N_34387,N_23916,N_20002);
xnor U34388 (N_34388,N_24488,N_27276);
and U34389 (N_34389,N_23479,N_21784);
xor U34390 (N_34390,N_29436,N_20727);
xnor U34391 (N_34391,N_27553,N_24714);
nor U34392 (N_34392,N_20212,N_29476);
and U34393 (N_34393,N_22845,N_24301);
nand U34394 (N_34394,N_25128,N_20897);
nand U34395 (N_34395,N_27997,N_23291);
nor U34396 (N_34396,N_27463,N_28125);
or U34397 (N_34397,N_25344,N_27394);
nor U34398 (N_34398,N_20503,N_21062);
and U34399 (N_34399,N_22837,N_25278);
nor U34400 (N_34400,N_27294,N_29972);
and U34401 (N_34401,N_22114,N_29685);
xnor U34402 (N_34402,N_26767,N_21097);
xor U34403 (N_34403,N_24652,N_22612);
nor U34404 (N_34404,N_27030,N_27255);
xnor U34405 (N_34405,N_22235,N_28515);
or U34406 (N_34406,N_21507,N_24417);
or U34407 (N_34407,N_24189,N_21703);
and U34408 (N_34408,N_22322,N_22953);
and U34409 (N_34409,N_23922,N_23919);
or U34410 (N_34410,N_21582,N_21204);
nor U34411 (N_34411,N_20697,N_23217);
or U34412 (N_34412,N_21500,N_20679);
nand U34413 (N_34413,N_29841,N_25221);
or U34414 (N_34414,N_27759,N_22098);
and U34415 (N_34415,N_28070,N_27800);
nor U34416 (N_34416,N_20460,N_24968);
and U34417 (N_34417,N_29413,N_24683);
nand U34418 (N_34418,N_21706,N_23284);
xnor U34419 (N_34419,N_21292,N_28543);
xnor U34420 (N_34420,N_26657,N_23329);
and U34421 (N_34421,N_25504,N_26320);
nand U34422 (N_34422,N_20068,N_29074);
xor U34423 (N_34423,N_23031,N_29828);
and U34424 (N_34424,N_20114,N_22896);
nor U34425 (N_34425,N_25954,N_29480);
or U34426 (N_34426,N_24250,N_22597);
xor U34427 (N_34427,N_20643,N_28977);
or U34428 (N_34428,N_25492,N_26116);
or U34429 (N_34429,N_20098,N_23681);
xor U34430 (N_34430,N_24873,N_28876);
nand U34431 (N_34431,N_26212,N_20724);
or U34432 (N_34432,N_23426,N_29907);
nor U34433 (N_34433,N_23820,N_29656);
and U34434 (N_34434,N_25699,N_20839);
nor U34435 (N_34435,N_23213,N_29445);
nand U34436 (N_34436,N_29597,N_22164);
and U34437 (N_34437,N_27541,N_24783);
xnor U34438 (N_34438,N_27792,N_25373);
xor U34439 (N_34439,N_22057,N_23526);
nand U34440 (N_34440,N_27508,N_26536);
or U34441 (N_34441,N_20300,N_22530);
and U34442 (N_34442,N_27317,N_27917);
nor U34443 (N_34443,N_26906,N_26131);
nor U34444 (N_34444,N_22826,N_25785);
and U34445 (N_34445,N_26605,N_21147);
or U34446 (N_34446,N_26342,N_21574);
or U34447 (N_34447,N_29636,N_22731);
and U34448 (N_34448,N_24274,N_21058);
nor U34449 (N_34449,N_25047,N_27678);
nor U34450 (N_34450,N_29578,N_27910);
nor U34451 (N_34451,N_25908,N_20107);
nand U34452 (N_34452,N_25112,N_20047);
or U34453 (N_34453,N_25438,N_22170);
xor U34454 (N_34454,N_21167,N_26635);
and U34455 (N_34455,N_22441,N_20570);
nand U34456 (N_34456,N_22730,N_29988);
and U34457 (N_34457,N_28022,N_23645);
or U34458 (N_34458,N_23719,N_28165);
and U34459 (N_34459,N_26139,N_26446);
nor U34460 (N_34460,N_28581,N_24625);
xor U34461 (N_34461,N_23977,N_25709);
xor U34462 (N_34462,N_28136,N_22690);
or U34463 (N_34463,N_23117,N_25020);
nor U34464 (N_34464,N_23243,N_24929);
nor U34465 (N_34465,N_23020,N_22560);
or U34466 (N_34466,N_24745,N_21434);
nor U34467 (N_34467,N_29099,N_22365);
nand U34468 (N_34468,N_21186,N_28658);
nand U34469 (N_34469,N_23908,N_24760);
and U34470 (N_34470,N_26019,N_22662);
and U34471 (N_34471,N_20536,N_24724);
and U34472 (N_34472,N_26626,N_24068);
nor U34473 (N_34473,N_26998,N_28761);
or U34474 (N_34474,N_24903,N_27180);
nor U34475 (N_34475,N_25457,N_29120);
xor U34476 (N_34476,N_25108,N_25865);
nor U34477 (N_34477,N_20096,N_22586);
and U34478 (N_34478,N_24273,N_28600);
and U34479 (N_34479,N_20119,N_20316);
nand U34480 (N_34480,N_22696,N_26902);
nand U34481 (N_34481,N_29086,N_29174);
and U34482 (N_34482,N_27179,N_26468);
or U34483 (N_34483,N_21968,N_25808);
nor U34484 (N_34484,N_26555,N_29475);
or U34485 (N_34485,N_26210,N_28105);
and U34486 (N_34486,N_27540,N_25712);
xor U34487 (N_34487,N_20169,N_25483);
or U34488 (N_34488,N_29338,N_22809);
nand U34489 (N_34489,N_26245,N_26622);
nand U34490 (N_34490,N_24813,N_21723);
xor U34491 (N_34491,N_20514,N_22184);
nor U34492 (N_34492,N_20962,N_23509);
or U34493 (N_34493,N_27402,N_23679);
or U34494 (N_34494,N_24692,N_29118);
nor U34495 (N_34495,N_24015,N_24647);
or U34496 (N_34496,N_28428,N_26112);
xnor U34497 (N_34497,N_24609,N_26077);
and U34498 (N_34498,N_21509,N_25002);
nor U34499 (N_34499,N_21902,N_29814);
nand U34500 (N_34500,N_27988,N_27086);
nor U34501 (N_34501,N_27613,N_22813);
xnor U34502 (N_34502,N_28141,N_29020);
and U34503 (N_34503,N_20553,N_29531);
and U34504 (N_34504,N_29098,N_25213);
nand U34505 (N_34505,N_29721,N_25372);
or U34506 (N_34506,N_29600,N_20371);
nor U34507 (N_34507,N_26611,N_24497);
nand U34508 (N_34508,N_27213,N_20625);
and U34509 (N_34509,N_27042,N_21696);
nor U34510 (N_34510,N_24559,N_24710);
nand U34511 (N_34511,N_21543,N_23606);
or U34512 (N_34512,N_23239,N_28814);
nand U34513 (N_34513,N_22126,N_20888);
and U34514 (N_34514,N_27554,N_29066);
nand U34515 (N_34515,N_25568,N_28956);
xor U34516 (N_34516,N_28736,N_28351);
nand U34517 (N_34517,N_28255,N_29952);
nand U34518 (N_34518,N_21195,N_25156);
and U34519 (N_34519,N_26135,N_26216);
nor U34520 (N_34520,N_21347,N_21193);
nor U34521 (N_34521,N_20449,N_29889);
and U34522 (N_34522,N_28935,N_25093);
nand U34523 (N_34523,N_27512,N_28938);
xnor U34524 (N_34524,N_20731,N_24707);
xnor U34525 (N_34525,N_21240,N_20388);
or U34526 (N_34526,N_24023,N_21925);
and U34527 (N_34527,N_26175,N_23967);
and U34528 (N_34528,N_23650,N_25713);
and U34529 (N_34529,N_29472,N_23478);
or U34530 (N_34530,N_27807,N_24537);
or U34531 (N_34531,N_25243,N_25327);
or U34532 (N_34532,N_21294,N_22563);
and U34533 (N_34533,N_22362,N_28678);
nor U34534 (N_34534,N_21271,N_22553);
xnor U34535 (N_34535,N_20245,N_25556);
nand U34536 (N_34536,N_23460,N_21049);
and U34537 (N_34537,N_24856,N_22027);
or U34538 (N_34538,N_24706,N_28324);
nand U34539 (N_34539,N_25274,N_29673);
and U34540 (N_34540,N_25721,N_20749);
or U34541 (N_34541,N_27044,N_29384);
and U34542 (N_34542,N_26847,N_25831);
nand U34543 (N_34543,N_29614,N_27813);
or U34544 (N_34544,N_27674,N_29483);
and U34545 (N_34545,N_27081,N_29134);
and U34546 (N_34546,N_20226,N_27232);
nor U34547 (N_34547,N_27378,N_22312);
nand U34548 (N_34548,N_29289,N_23549);
nand U34549 (N_34549,N_22477,N_20515);
and U34550 (N_34550,N_26298,N_23374);
nor U34551 (N_34551,N_28310,N_24629);
nand U34552 (N_34552,N_27639,N_25948);
nor U34553 (N_34553,N_27328,N_20876);
and U34554 (N_34554,N_23428,N_23355);
nor U34555 (N_34555,N_22534,N_23446);
nand U34556 (N_34556,N_24673,N_22565);
and U34557 (N_34557,N_25835,N_23609);
and U34558 (N_34558,N_21667,N_29166);
nor U34559 (N_34559,N_27129,N_21632);
nand U34560 (N_34560,N_29829,N_23080);
or U34561 (N_34561,N_26091,N_23358);
nand U34562 (N_34562,N_27945,N_24851);
nand U34563 (N_34563,N_25707,N_23260);
and U34564 (N_34564,N_28177,N_28835);
nand U34565 (N_34565,N_28985,N_23236);
nand U34566 (N_34566,N_27157,N_24568);
nand U34567 (N_34567,N_26641,N_29902);
or U34568 (N_34568,N_29694,N_29414);
nand U34569 (N_34569,N_24727,N_29630);
nor U34570 (N_34570,N_23647,N_22309);
nor U34571 (N_34571,N_28893,N_21718);
and U34572 (N_34572,N_24457,N_21584);
xor U34573 (N_34573,N_25240,N_29225);
nand U34574 (N_34574,N_21114,N_21043);
xnor U34575 (N_34575,N_22125,N_20556);
and U34576 (N_34576,N_27561,N_24904);
xor U34577 (N_34577,N_24131,N_22345);
and U34578 (N_34578,N_22202,N_29760);
and U34579 (N_34579,N_24178,N_27015);
and U34580 (N_34580,N_27753,N_20217);
nand U34581 (N_34581,N_26652,N_21245);
nand U34582 (N_34582,N_21318,N_28403);
nand U34583 (N_34583,N_26637,N_23806);
nand U34584 (N_34584,N_29488,N_22133);
xnor U34585 (N_34585,N_27605,N_29894);
or U34586 (N_34586,N_29361,N_26678);
and U34587 (N_34587,N_27635,N_27039);
xor U34588 (N_34588,N_21477,N_25371);
xor U34589 (N_34589,N_21015,N_21997);
xnor U34590 (N_34590,N_29400,N_28479);
nand U34591 (N_34591,N_22698,N_22892);
and U34592 (N_34592,N_23258,N_24495);
and U34593 (N_34593,N_28470,N_28769);
nand U34594 (N_34594,N_20327,N_24860);
xor U34595 (N_34595,N_24018,N_29357);
nor U34596 (N_34596,N_26162,N_25679);
nor U34597 (N_34597,N_27299,N_24475);
nand U34598 (N_34598,N_21724,N_27292);
nor U34599 (N_34599,N_22729,N_22956);
or U34600 (N_34600,N_21924,N_25157);
xnor U34601 (N_34601,N_20560,N_22775);
and U34602 (N_34602,N_27456,N_24163);
nand U34603 (N_34603,N_25528,N_23165);
or U34604 (N_34604,N_24510,N_20084);
nor U34605 (N_34605,N_26526,N_28262);
nand U34606 (N_34606,N_24784,N_28560);
and U34607 (N_34607,N_28104,N_28891);
nor U34608 (N_34608,N_22633,N_25555);
nand U34609 (N_34609,N_22208,N_24352);
xor U34610 (N_34610,N_22077,N_27968);
and U34611 (N_34611,N_24331,N_25194);
nand U34612 (N_34612,N_24623,N_20347);
nor U34613 (N_34613,N_21982,N_25129);
nand U34614 (N_34614,N_21906,N_24161);
and U34615 (N_34615,N_24214,N_26520);
nor U34616 (N_34616,N_26067,N_29418);
xor U34617 (N_34617,N_25351,N_23926);
or U34618 (N_34618,N_26658,N_21478);
nor U34619 (N_34619,N_21791,N_26471);
nand U34620 (N_34620,N_29198,N_20998);
xnor U34621 (N_34621,N_24359,N_23797);
and U34622 (N_34622,N_28344,N_21440);
nand U34623 (N_34623,N_25300,N_22759);
nor U34624 (N_34624,N_28014,N_26102);
nor U34625 (N_34625,N_27532,N_26619);
xor U34626 (N_34626,N_23913,N_28234);
and U34627 (N_34627,N_27948,N_21523);
nand U34628 (N_34628,N_20704,N_23709);
and U34629 (N_34629,N_20785,N_21662);
and U34630 (N_34630,N_25889,N_27093);
nand U34631 (N_34631,N_29316,N_29639);
nand U34632 (N_34632,N_29756,N_21618);
xor U34633 (N_34633,N_20215,N_20248);
and U34634 (N_34634,N_28498,N_25586);
or U34635 (N_34635,N_25428,N_23104);
and U34636 (N_34636,N_25169,N_27487);
nor U34637 (N_34637,N_22061,N_25052);
nand U34638 (N_34638,N_26317,N_27411);
nand U34639 (N_34639,N_20406,N_25757);
or U34640 (N_34640,N_25559,N_20335);
nor U34641 (N_34641,N_24603,N_22496);
xor U34642 (N_34642,N_20682,N_28113);
or U34643 (N_34643,N_25776,N_22939);
and U34644 (N_34644,N_23720,N_25232);
or U34645 (N_34645,N_28221,N_20452);
or U34646 (N_34646,N_20762,N_22735);
nand U34647 (N_34647,N_27964,N_27455);
or U34648 (N_34648,N_22480,N_24515);
nand U34649 (N_34649,N_25450,N_27966);
nand U34650 (N_34650,N_24362,N_21120);
nor U34651 (N_34651,N_26588,N_27072);
and U34652 (N_34652,N_26063,N_25807);
xnor U34653 (N_34653,N_21531,N_25225);
or U34654 (N_34654,N_20139,N_20921);
or U34655 (N_34655,N_20280,N_21892);
nor U34656 (N_34656,N_28290,N_29363);
nor U34657 (N_34657,N_24353,N_23542);
nand U34658 (N_34658,N_29910,N_29882);
or U34659 (N_34659,N_20396,N_29239);
or U34660 (N_34660,N_25907,N_24271);
and U34661 (N_34661,N_29264,N_28063);
or U34662 (N_34662,N_25369,N_27454);
nand U34663 (N_34663,N_26482,N_27765);
and U34664 (N_34664,N_22853,N_27398);
nor U34665 (N_34665,N_29925,N_20322);
xnor U34666 (N_34666,N_28335,N_29438);
nand U34667 (N_34667,N_20209,N_25397);
nand U34668 (N_34668,N_22529,N_26073);
nand U34669 (N_34669,N_28195,N_27991);
nor U34670 (N_34670,N_21544,N_22348);
or U34671 (N_34671,N_21976,N_23569);
nor U34672 (N_34672,N_28270,N_21098);
nor U34673 (N_34673,N_29560,N_23938);
nor U34674 (N_34674,N_24112,N_23885);
nand U34675 (N_34675,N_29786,N_29262);
nand U34676 (N_34676,N_24955,N_25833);
and U34677 (N_34677,N_21975,N_26905);
xnor U34678 (N_34678,N_21698,N_24973);
or U34679 (N_34679,N_20144,N_21541);
and U34680 (N_34680,N_22152,N_29083);
and U34681 (N_34681,N_24198,N_27527);
or U34682 (N_34682,N_22823,N_21126);
and U34683 (N_34683,N_22625,N_26489);
and U34684 (N_34684,N_21077,N_21164);
or U34685 (N_34685,N_21080,N_29390);
nand U34686 (N_34686,N_22131,N_27834);
xor U34687 (N_34687,N_29939,N_22452);
and U34688 (N_34688,N_24004,N_24656);
nor U34689 (N_34689,N_28140,N_20137);
nor U34690 (N_34690,N_26792,N_21731);
and U34691 (N_34691,N_24085,N_29514);
nand U34692 (N_34692,N_24401,N_24566);
or U34693 (N_34693,N_27546,N_29846);
and U34694 (N_34694,N_28923,N_28800);
and U34695 (N_34695,N_28465,N_22301);
and U34696 (N_34696,N_21602,N_20877);
xor U34697 (N_34697,N_28511,N_27337);
xnor U34698 (N_34698,N_25552,N_25250);
xnor U34699 (N_34699,N_21132,N_25325);
or U34700 (N_34700,N_28314,N_23039);
nor U34701 (N_34701,N_26072,N_24505);
xnor U34702 (N_34702,N_28642,N_28807);
and U34703 (N_34703,N_21388,N_22937);
nand U34704 (N_34704,N_29631,N_21349);
nand U34705 (N_34705,N_20670,N_29410);
nand U34706 (N_34706,N_27189,N_27742);
nor U34707 (N_34707,N_25952,N_21725);
nand U34708 (N_34708,N_20583,N_23012);
and U34709 (N_34709,N_25338,N_29700);
and U34710 (N_34710,N_20401,N_23951);
nand U34711 (N_34711,N_25569,N_22144);
nor U34712 (N_34712,N_21501,N_25657);
nand U34713 (N_34713,N_28397,N_25472);
nor U34714 (N_34714,N_23370,N_28673);
nand U34715 (N_34715,N_28689,N_20585);
nand U34716 (N_34716,N_28574,N_22679);
and U34717 (N_34717,N_23247,N_23787);
nor U34718 (N_34718,N_27327,N_20267);
or U34719 (N_34719,N_21781,N_21159);
or U34720 (N_34720,N_28928,N_26100);
and U34721 (N_34721,N_20675,N_23713);
xnor U34722 (N_34722,N_23680,N_24941);
and U34723 (N_34723,N_24871,N_28522);
nand U34724 (N_34724,N_26159,N_29928);
nand U34725 (N_34725,N_29321,N_29055);
xor U34726 (N_34726,N_23445,N_26167);
nand U34727 (N_34727,N_29575,N_24854);
nor U34728 (N_34728,N_21442,N_20020);
xor U34729 (N_34729,N_29791,N_27155);
or U34730 (N_34730,N_29509,N_26391);
xnor U34731 (N_34731,N_23304,N_28920);
and U34732 (N_34732,N_23484,N_21431);
xor U34733 (N_34733,N_25107,N_28118);
nand U34734 (N_34734,N_24223,N_23523);
xnor U34735 (N_34735,N_25089,N_23352);
and U34736 (N_34736,N_28236,N_25545);
nor U34737 (N_34737,N_29566,N_21115);
and U34738 (N_34738,N_24396,N_22694);
and U34739 (N_34739,N_23594,N_22840);
or U34740 (N_34740,N_20868,N_26778);
nand U34741 (N_34741,N_29122,N_23652);
nand U34742 (N_34742,N_22484,N_27160);
xnor U34743 (N_34743,N_20953,N_25302);
and U34744 (N_34744,N_20581,N_23905);
or U34745 (N_34745,N_27080,N_26567);
nand U34746 (N_34746,N_25144,N_21849);
nand U34747 (N_34747,N_26973,N_28556);
xnor U34748 (N_34748,N_21871,N_24702);
and U34749 (N_34749,N_20395,N_20572);
nor U34750 (N_34750,N_25968,N_22903);
nor U34751 (N_34751,N_29109,N_29658);
nand U34752 (N_34752,N_28744,N_24176);
or U34753 (N_34753,N_28727,N_27939);
or U34754 (N_34754,N_21595,N_25354);
nor U34755 (N_34755,N_29032,N_24216);
and U34756 (N_34756,N_22084,N_24298);
and U34757 (N_34757,N_27116,N_25430);
nor U34758 (N_34758,N_22317,N_27940);
or U34759 (N_34759,N_23398,N_26319);
xor U34760 (N_34760,N_26988,N_22713);
nor U34761 (N_34761,N_22611,N_29425);
nand U34762 (N_34762,N_27502,N_23140);
and U34763 (N_34763,N_22850,N_24514);
nor U34764 (N_34764,N_29286,N_20599);
nand U34765 (N_34765,N_28039,N_26334);
and U34766 (N_34766,N_29507,N_26368);
nor U34767 (N_34767,N_20602,N_29963);
xor U34768 (N_34768,N_29823,N_22289);
or U34769 (N_34769,N_22906,N_24397);
nor U34770 (N_34770,N_25111,N_23309);
and U34771 (N_34771,N_22581,N_20163);
or U34772 (N_34772,N_21041,N_24970);
and U34773 (N_34773,N_24469,N_28577);
or U34774 (N_34774,N_23415,N_27315);
or U34775 (N_34775,N_24501,N_27640);
nor U34776 (N_34776,N_25409,N_28157);
nand U34777 (N_34777,N_23582,N_22447);
xor U34778 (N_34778,N_22749,N_24063);
xor U34779 (N_34779,N_23024,N_26646);
nand U34780 (N_34780,N_29912,N_21396);
and U34781 (N_34781,N_26879,N_26654);
and U34782 (N_34782,N_27515,N_28849);
and U34783 (N_34783,N_24816,N_23011);
or U34784 (N_34784,N_29853,N_22888);
xor U34785 (N_34785,N_23470,N_25290);
and U34786 (N_34786,N_25029,N_27729);
or U34787 (N_34787,N_25988,N_25415);
nor U34788 (N_34788,N_20945,N_28406);
nor U34789 (N_34789,N_21623,N_26551);
or U34790 (N_34790,N_29137,N_27597);
and U34791 (N_34791,N_29307,N_26157);
or U34792 (N_34792,N_21858,N_21587);
and U34793 (N_34793,N_28196,N_25876);
nor U34794 (N_34794,N_29474,N_29145);
nand U34795 (N_34795,N_26713,N_28638);
or U34796 (N_34796,N_29417,N_20696);
xor U34797 (N_34797,N_22250,N_25422);
nand U34798 (N_34798,N_24124,N_24125);
xor U34799 (N_34799,N_24939,N_25403);
nor U34800 (N_34800,N_26406,N_25329);
nor U34801 (N_34801,N_21746,N_29232);
or U34802 (N_34802,N_27090,N_26506);
nor U34803 (N_34803,N_20331,N_26338);
nand U34804 (N_34804,N_24141,N_23631);
nand U34805 (N_34805,N_29870,N_20053);
xnor U34806 (N_34806,N_23049,N_24803);
and U34807 (N_34807,N_21485,N_24494);
or U34808 (N_34808,N_22428,N_26031);
nand U34809 (N_34809,N_28060,N_27993);
nor U34810 (N_34810,N_26238,N_20263);
nor U34811 (N_34811,N_24350,N_20482);
nand U34812 (N_34812,N_25282,N_25818);
nand U34813 (N_34813,N_20191,N_29220);
or U34814 (N_34814,N_20928,N_28284);
nand U34815 (N_34815,N_20469,N_24097);
xnor U34816 (N_34816,N_22282,N_28488);
or U34817 (N_34817,N_24518,N_23491);
or U34818 (N_34818,N_29544,N_20013);
and U34819 (N_34819,N_28376,N_24309);
nor U34820 (N_34820,N_29179,N_28889);
or U34821 (N_34821,N_27414,N_21202);
or U34822 (N_34822,N_29056,N_21671);
or U34823 (N_34823,N_29747,N_28592);
or U34824 (N_34824,N_24119,N_24230);
xnor U34825 (N_34825,N_25145,N_27504);
or U34826 (N_34826,N_24210,N_24894);
and U34827 (N_34827,N_29901,N_25470);
xor U34828 (N_34828,N_22842,N_26687);
xor U34829 (N_34829,N_22678,N_28229);
nand U34830 (N_34830,N_23583,N_23390);
nand U34831 (N_34831,N_28115,N_28366);
xnor U34832 (N_34832,N_29767,N_23798);
and U34833 (N_34833,N_27831,N_22928);
xor U34834 (N_34834,N_27927,N_22413);
nand U34835 (N_34835,N_25872,N_23003);
xnor U34836 (N_34836,N_27013,N_28239);
or U34837 (N_34837,N_26202,N_24807);
and U34838 (N_34838,N_27754,N_21506);
or U34839 (N_34839,N_26042,N_20943);
or U34840 (N_34840,N_25834,N_27594);
nor U34841 (N_34841,N_28844,N_29941);
or U34842 (N_34842,N_21508,N_28907);
nand U34843 (N_34843,N_26686,N_20563);
xnor U34844 (N_34844,N_22188,N_24528);
nand U34845 (N_34845,N_24850,N_23915);
and U34846 (N_34846,N_25587,N_24809);
nand U34847 (N_34847,N_28647,N_23716);
or U34848 (N_34848,N_29729,N_23550);
nand U34849 (N_34849,N_23184,N_25924);
xor U34850 (N_34850,N_23495,N_22979);
nand U34851 (N_34851,N_28888,N_25887);
or U34852 (N_34852,N_21920,N_27195);
nand U34853 (N_34853,N_27892,N_23881);
nand U34854 (N_34854,N_26600,N_23077);
or U34855 (N_34855,N_27216,N_29235);
nor U34856 (N_34856,N_24224,N_24190);
or U34857 (N_34857,N_25764,N_28493);
nand U34858 (N_34858,N_22768,N_24027);
or U34859 (N_34859,N_21772,N_26372);
and U34860 (N_34860,N_22041,N_27324);
and U34861 (N_34861,N_27731,N_20851);
nor U34862 (N_34862,N_25502,N_24086);
or U34863 (N_34863,N_29298,N_27298);
xnor U34864 (N_34864,N_21238,N_28926);
nand U34865 (N_34865,N_23310,N_26062);
xor U34866 (N_34866,N_21551,N_22885);
xnor U34867 (N_34867,N_29973,N_20886);
or U34868 (N_34868,N_27723,N_25488);
and U34869 (N_34869,N_20261,N_24199);
or U34870 (N_34870,N_23572,N_24717);
xnor U34871 (N_34871,N_20332,N_21946);
nor U34872 (N_34872,N_27319,N_29998);
nand U34873 (N_34873,N_27852,N_27056);
xnor U34874 (N_34874,N_25548,N_24003);
or U34875 (N_34875,N_27562,N_26854);
xnor U34876 (N_34876,N_29265,N_29211);
nand U34877 (N_34877,N_27211,N_21974);
nor U34878 (N_34878,N_28936,N_28167);
and U34879 (N_34879,N_20235,N_24435);
nor U34880 (N_34880,N_29295,N_26393);
nand U34881 (N_34881,N_25986,N_29974);
or U34882 (N_34882,N_20325,N_23212);
nand U34883 (N_34883,N_23888,N_28395);
nor U34884 (N_34884,N_21903,N_27538);
nor U34885 (N_34885,N_23697,N_24269);
nand U34886 (N_34886,N_21588,N_28399);
nand U34887 (N_34887,N_25572,N_21515);
nor U34888 (N_34888,N_28357,N_20582);
or U34889 (N_34889,N_21074,N_20121);
and U34890 (N_34890,N_26846,N_21657);
and U34891 (N_34891,N_28460,N_25003);
xor U34892 (N_34892,N_29181,N_28702);
xor U34893 (N_34893,N_23311,N_24263);
nand U34894 (N_34894,N_28822,N_24013);
or U34895 (N_34895,N_27031,N_22052);
xor U34896 (N_34896,N_21219,N_27439);
xnor U34897 (N_34897,N_28092,N_22591);
and U34898 (N_34898,N_25633,N_20374);
xor U34899 (N_34899,N_22392,N_21807);
nand U34900 (N_34900,N_25473,N_22914);
and U34901 (N_34901,N_23244,N_28567);
nand U34902 (N_34902,N_21916,N_27320);
or U34903 (N_34903,N_29139,N_28182);
and U34904 (N_34904,N_21919,N_21913);
or U34905 (N_34905,N_20778,N_22199);
nand U34906 (N_34906,N_25882,N_22502);
nand U34907 (N_34907,N_23761,N_25981);
nand U34908 (N_34908,N_25913,N_22473);
nand U34909 (N_34909,N_28447,N_22408);
xor U34910 (N_34910,N_27676,N_25536);
xor U34911 (N_34911,N_24547,N_29586);
or U34912 (N_34912,N_27752,N_25686);
nand U34913 (N_34913,N_29708,N_28572);
and U34914 (N_34914,N_22587,N_25069);
nor U34915 (N_34915,N_22409,N_23064);
nor U34916 (N_34916,N_23290,N_24186);
nor U34917 (N_34917,N_29336,N_27983);
or U34918 (N_34918,N_20922,N_24892);
or U34919 (N_34919,N_25227,N_22147);
and U34920 (N_34920,N_21201,N_24395);
nand U34921 (N_34921,N_28180,N_22112);
or U34922 (N_34922,N_25163,N_28391);
xor U34923 (N_34923,N_23876,N_28276);
xor U34924 (N_34924,N_26301,N_23267);
and U34925 (N_34925,N_20827,N_26947);
and U34926 (N_34926,N_26383,N_27077);
or U34927 (N_34927,N_25837,N_29502);
nor U34928 (N_34928,N_25097,N_24242);
or U34929 (N_34929,N_24852,N_26797);
nand U34930 (N_34930,N_20313,N_29308);
or U34931 (N_34931,N_20309,N_23225);
and U34932 (N_34932,N_27698,N_25812);
and U34933 (N_34933,N_28086,N_21583);
and U34934 (N_34934,N_23662,N_21461);
and U34935 (N_34935,N_22204,N_29422);
and U34936 (N_34936,N_22664,N_29843);
and U34937 (N_34937,N_29047,N_23034);
nand U34938 (N_34938,N_29061,N_25110);
nand U34939 (N_34939,N_21337,N_29634);
nand U34940 (N_34940,N_26484,N_21390);
or U34941 (N_34941,N_20601,N_23251);
or U34942 (N_34942,N_26462,N_25659);
or U34943 (N_34943,N_23945,N_28474);
xnor U34944 (N_34944,N_21340,N_22180);
and U34945 (N_34945,N_23889,N_20289);
nand U34946 (N_34946,N_23004,N_28915);
and U34947 (N_34947,N_26140,N_28163);
nand U34948 (N_34948,N_20863,N_25195);
nand U34949 (N_34949,N_27003,N_28539);
xnor U34950 (N_34950,N_26015,N_24212);
xor U34951 (N_34951,N_26057,N_26474);
nand U34952 (N_34952,N_29942,N_28256);
nor U34953 (N_34953,N_29799,N_25621);
and U34954 (N_34954,N_21634,N_26711);
and U34955 (N_34955,N_25664,N_20580);
and U34956 (N_34956,N_21984,N_25341);
nand U34957 (N_34957,N_29855,N_29761);
nor U34958 (N_34958,N_25670,N_26994);
nor U34959 (N_34959,N_22508,N_25930);
nand U34960 (N_34960,N_22677,N_21717);
and U34961 (N_34961,N_22388,N_26917);
nor U34962 (N_34962,N_21437,N_27548);
nor U34963 (N_34963,N_28471,N_27383);
nand U34964 (N_34964,N_27482,N_24913);
nand U34965 (N_34965,N_29184,N_29596);
xor U34966 (N_34966,N_25959,N_21348);
and U34967 (N_34967,N_20143,N_25159);
xor U34968 (N_34968,N_21458,N_23552);
nor U34969 (N_34969,N_29296,N_23600);
xor U34970 (N_34970,N_27715,N_22717);
xor U34971 (N_34971,N_23520,N_24447);
or U34972 (N_34972,N_21859,N_28550);
xor U34973 (N_34973,N_20729,N_23078);
and U34974 (N_34974,N_26726,N_21969);
xnor U34975 (N_34975,N_21855,N_20637);
nor U34976 (N_34976,N_21044,N_27544);
nor U34977 (N_34977,N_27928,N_20222);
nor U34978 (N_34978,N_23868,N_26397);
or U34979 (N_34979,N_29423,N_21939);
and U34980 (N_34980,N_27705,N_20920);
nor U34981 (N_34981,N_22744,N_20353);
or U34982 (N_34982,N_27417,N_25613);
or U34983 (N_34983,N_28075,N_29213);
xnor U34984 (N_34984,N_26999,N_27033);
xor U34985 (N_34985,N_28015,N_27922);
nand U34986 (N_34986,N_28832,N_20078);
xor U34987 (N_34987,N_21197,N_28491);
xor U34988 (N_34988,N_21805,N_25036);
nor U34989 (N_34989,N_26282,N_24636);
xor U34990 (N_34990,N_28672,N_27595);
xor U34991 (N_34991,N_22810,N_29765);
xnor U34992 (N_34992,N_21964,N_29234);
and U34993 (N_34993,N_20918,N_24437);
nand U34994 (N_34994,N_28210,N_29012);
or U34995 (N_34995,N_26017,N_25507);
nand U34996 (N_34996,N_20623,N_26346);
xor U34997 (N_34997,N_23667,N_29399);
nor U34998 (N_34998,N_28362,N_28910);
xor U34999 (N_34999,N_20458,N_21379);
xnor U35000 (N_35000,N_28981,N_27689);
xnor U35001 (N_35001,N_22753,N_21995);
nor U35002 (N_35002,N_24692,N_24821);
or U35003 (N_35003,N_23392,N_23152);
and U35004 (N_35004,N_27902,N_26388);
xor U35005 (N_35005,N_20035,N_27803);
nand U35006 (N_35006,N_23042,N_24271);
xnor U35007 (N_35007,N_29076,N_29847);
nand U35008 (N_35008,N_21709,N_25307);
nor U35009 (N_35009,N_25100,N_20285);
or U35010 (N_35010,N_23657,N_27081);
nor U35011 (N_35011,N_21895,N_29908);
nor U35012 (N_35012,N_26675,N_21098);
or U35013 (N_35013,N_24696,N_28988);
nand U35014 (N_35014,N_21590,N_25360);
or U35015 (N_35015,N_29783,N_22027);
nand U35016 (N_35016,N_22745,N_29507);
and U35017 (N_35017,N_21263,N_21083);
nor U35018 (N_35018,N_22326,N_27348);
and U35019 (N_35019,N_27053,N_22687);
nand U35020 (N_35020,N_23309,N_27671);
or U35021 (N_35021,N_28155,N_20827);
nor U35022 (N_35022,N_24477,N_27218);
and U35023 (N_35023,N_24804,N_20113);
xor U35024 (N_35024,N_24434,N_26187);
xnor U35025 (N_35025,N_26744,N_21241);
xor U35026 (N_35026,N_25525,N_29343);
or U35027 (N_35027,N_21915,N_20419);
xnor U35028 (N_35028,N_27927,N_24955);
nor U35029 (N_35029,N_21616,N_23681);
nand U35030 (N_35030,N_26602,N_28410);
xor U35031 (N_35031,N_29034,N_27784);
or U35032 (N_35032,N_27595,N_24787);
nor U35033 (N_35033,N_26649,N_25836);
or U35034 (N_35034,N_26388,N_20077);
or U35035 (N_35035,N_21864,N_21145);
nand U35036 (N_35036,N_29267,N_25203);
nand U35037 (N_35037,N_25672,N_29989);
nor U35038 (N_35038,N_22049,N_27283);
nand U35039 (N_35039,N_23762,N_24047);
nand U35040 (N_35040,N_22612,N_21058);
or U35041 (N_35041,N_29397,N_26882);
xor U35042 (N_35042,N_29874,N_28340);
xor U35043 (N_35043,N_28360,N_22452);
xor U35044 (N_35044,N_27921,N_29490);
and U35045 (N_35045,N_27566,N_29883);
nand U35046 (N_35046,N_20541,N_28521);
nand U35047 (N_35047,N_21592,N_21461);
nand U35048 (N_35048,N_28032,N_27241);
nand U35049 (N_35049,N_23150,N_24759);
nand U35050 (N_35050,N_22270,N_23807);
and U35051 (N_35051,N_28679,N_28345);
xor U35052 (N_35052,N_22882,N_25419);
and U35053 (N_35053,N_26480,N_22987);
nor U35054 (N_35054,N_22991,N_28322);
nor U35055 (N_35055,N_23781,N_24874);
or U35056 (N_35056,N_26984,N_23130);
nand U35057 (N_35057,N_28585,N_25041);
nand U35058 (N_35058,N_22682,N_29913);
and U35059 (N_35059,N_25285,N_29120);
nor U35060 (N_35060,N_20850,N_28926);
nor U35061 (N_35061,N_28537,N_26999);
and U35062 (N_35062,N_22276,N_29951);
or U35063 (N_35063,N_26166,N_23801);
xor U35064 (N_35064,N_22144,N_28448);
or U35065 (N_35065,N_21257,N_25302);
xor U35066 (N_35066,N_22391,N_28960);
nand U35067 (N_35067,N_20946,N_23895);
and U35068 (N_35068,N_28773,N_25452);
nand U35069 (N_35069,N_24193,N_21463);
nand U35070 (N_35070,N_29176,N_28538);
xnor U35071 (N_35071,N_22505,N_21974);
nand U35072 (N_35072,N_26814,N_28739);
nand U35073 (N_35073,N_21085,N_26845);
and U35074 (N_35074,N_23155,N_21613);
nor U35075 (N_35075,N_26819,N_28868);
nor U35076 (N_35076,N_22424,N_22662);
or U35077 (N_35077,N_22738,N_25248);
and U35078 (N_35078,N_25684,N_28164);
or U35079 (N_35079,N_27846,N_28077);
and U35080 (N_35080,N_23129,N_28030);
or U35081 (N_35081,N_26206,N_22916);
and U35082 (N_35082,N_25479,N_23624);
nand U35083 (N_35083,N_25946,N_28799);
xor U35084 (N_35084,N_29962,N_27629);
and U35085 (N_35085,N_27979,N_25171);
xnor U35086 (N_35086,N_22153,N_20639);
nor U35087 (N_35087,N_28074,N_26009);
or U35088 (N_35088,N_21994,N_28295);
or U35089 (N_35089,N_21577,N_24118);
and U35090 (N_35090,N_27949,N_20858);
and U35091 (N_35091,N_27988,N_22778);
nand U35092 (N_35092,N_28474,N_24737);
nand U35093 (N_35093,N_23532,N_28880);
nor U35094 (N_35094,N_20725,N_28479);
or U35095 (N_35095,N_26805,N_28010);
or U35096 (N_35096,N_22410,N_22438);
xnor U35097 (N_35097,N_22360,N_28411);
nor U35098 (N_35098,N_23368,N_21807);
or U35099 (N_35099,N_21483,N_22178);
or U35100 (N_35100,N_21937,N_26088);
and U35101 (N_35101,N_23223,N_20752);
or U35102 (N_35102,N_21017,N_27345);
nor U35103 (N_35103,N_23872,N_27402);
xor U35104 (N_35104,N_23947,N_24644);
xor U35105 (N_35105,N_29077,N_28526);
and U35106 (N_35106,N_26055,N_28948);
or U35107 (N_35107,N_21563,N_21083);
and U35108 (N_35108,N_23340,N_26752);
nand U35109 (N_35109,N_26323,N_24886);
and U35110 (N_35110,N_28797,N_28022);
xor U35111 (N_35111,N_26749,N_29121);
nor U35112 (N_35112,N_23894,N_27973);
nor U35113 (N_35113,N_28825,N_27943);
xor U35114 (N_35114,N_29144,N_20748);
and U35115 (N_35115,N_23028,N_28937);
or U35116 (N_35116,N_27447,N_29047);
xnor U35117 (N_35117,N_22350,N_20429);
nand U35118 (N_35118,N_24618,N_28432);
or U35119 (N_35119,N_23703,N_28676);
nand U35120 (N_35120,N_22452,N_20438);
nand U35121 (N_35121,N_25619,N_26926);
xnor U35122 (N_35122,N_27888,N_20049);
nand U35123 (N_35123,N_29435,N_21436);
and U35124 (N_35124,N_26007,N_26147);
or U35125 (N_35125,N_28108,N_20084);
xnor U35126 (N_35126,N_21598,N_27181);
xnor U35127 (N_35127,N_23025,N_28308);
xor U35128 (N_35128,N_24389,N_26023);
nand U35129 (N_35129,N_25811,N_22526);
and U35130 (N_35130,N_29319,N_28662);
or U35131 (N_35131,N_21646,N_23346);
xor U35132 (N_35132,N_21619,N_26871);
and U35133 (N_35133,N_20856,N_22856);
and U35134 (N_35134,N_27661,N_23793);
or U35135 (N_35135,N_23838,N_24359);
and U35136 (N_35136,N_28490,N_27058);
nor U35137 (N_35137,N_26755,N_23332);
or U35138 (N_35138,N_22961,N_23001);
or U35139 (N_35139,N_24217,N_22192);
xnor U35140 (N_35140,N_29535,N_25895);
nor U35141 (N_35141,N_28937,N_22413);
nand U35142 (N_35142,N_29360,N_25457);
or U35143 (N_35143,N_24653,N_23438);
nand U35144 (N_35144,N_20738,N_20643);
xor U35145 (N_35145,N_23079,N_25205);
or U35146 (N_35146,N_21594,N_27224);
or U35147 (N_35147,N_26446,N_21998);
nor U35148 (N_35148,N_29571,N_27995);
or U35149 (N_35149,N_22920,N_25913);
xnor U35150 (N_35150,N_29320,N_20848);
nand U35151 (N_35151,N_25090,N_27893);
and U35152 (N_35152,N_27995,N_20895);
nand U35153 (N_35153,N_21783,N_21520);
or U35154 (N_35154,N_24465,N_21370);
nand U35155 (N_35155,N_25384,N_21306);
nand U35156 (N_35156,N_29305,N_27618);
nand U35157 (N_35157,N_21883,N_27333);
xnor U35158 (N_35158,N_21792,N_23735);
or U35159 (N_35159,N_28658,N_21421);
nor U35160 (N_35160,N_25304,N_26476);
and U35161 (N_35161,N_26391,N_23508);
nor U35162 (N_35162,N_22605,N_23799);
xnor U35163 (N_35163,N_25665,N_28904);
or U35164 (N_35164,N_27961,N_26033);
xor U35165 (N_35165,N_29507,N_27960);
nand U35166 (N_35166,N_29900,N_24786);
xor U35167 (N_35167,N_21023,N_29431);
or U35168 (N_35168,N_24835,N_24338);
nand U35169 (N_35169,N_24743,N_23921);
and U35170 (N_35170,N_21997,N_27795);
nand U35171 (N_35171,N_21190,N_29370);
nor U35172 (N_35172,N_29636,N_26605);
or U35173 (N_35173,N_22724,N_29988);
xnor U35174 (N_35174,N_27131,N_21934);
nor U35175 (N_35175,N_28021,N_24644);
xnor U35176 (N_35176,N_22817,N_22511);
nor U35177 (N_35177,N_26109,N_21014);
nand U35178 (N_35178,N_28515,N_24867);
xor U35179 (N_35179,N_29999,N_24476);
nand U35180 (N_35180,N_29063,N_23292);
xor U35181 (N_35181,N_23655,N_23068);
xnor U35182 (N_35182,N_20886,N_28499);
nand U35183 (N_35183,N_23642,N_25295);
nor U35184 (N_35184,N_22075,N_24939);
xnor U35185 (N_35185,N_24187,N_28922);
and U35186 (N_35186,N_27594,N_29702);
nand U35187 (N_35187,N_25672,N_23200);
nor U35188 (N_35188,N_28760,N_28721);
and U35189 (N_35189,N_26315,N_23057);
or U35190 (N_35190,N_29880,N_21031);
nand U35191 (N_35191,N_21496,N_25629);
xnor U35192 (N_35192,N_22357,N_25161);
nand U35193 (N_35193,N_28760,N_27593);
xor U35194 (N_35194,N_28169,N_26811);
nor U35195 (N_35195,N_27485,N_23398);
nand U35196 (N_35196,N_23932,N_27886);
nor U35197 (N_35197,N_27135,N_24258);
or U35198 (N_35198,N_25089,N_20276);
xnor U35199 (N_35199,N_25875,N_23490);
xnor U35200 (N_35200,N_26691,N_25119);
and U35201 (N_35201,N_21565,N_26210);
nor U35202 (N_35202,N_27596,N_26416);
or U35203 (N_35203,N_28316,N_25062);
xor U35204 (N_35204,N_21972,N_20384);
nand U35205 (N_35205,N_27142,N_23652);
and U35206 (N_35206,N_26715,N_26902);
xor U35207 (N_35207,N_21559,N_28988);
nor U35208 (N_35208,N_27626,N_26494);
and U35209 (N_35209,N_25982,N_28503);
xor U35210 (N_35210,N_22607,N_26370);
and U35211 (N_35211,N_28416,N_22594);
and U35212 (N_35212,N_28406,N_28033);
or U35213 (N_35213,N_23139,N_22774);
nand U35214 (N_35214,N_22562,N_27481);
and U35215 (N_35215,N_24956,N_27115);
nor U35216 (N_35216,N_23191,N_23934);
xor U35217 (N_35217,N_23124,N_25225);
or U35218 (N_35218,N_23665,N_29538);
or U35219 (N_35219,N_23244,N_29389);
nor U35220 (N_35220,N_26856,N_21980);
nand U35221 (N_35221,N_27626,N_29272);
and U35222 (N_35222,N_24190,N_24246);
nor U35223 (N_35223,N_20567,N_23686);
nand U35224 (N_35224,N_20991,N_26437);
or U35225 (N_35225,N_27891,N_20807);
or U35226 (N_35226,N_23243,N_27602);
xor U35227 (N_35227,N_20507,N_24473);
nand U35228 (N_35228,N_23180,N_28497);
nor U35229 (N_35229,N_28162,N_23684);
xor U35230 (N_35230,N_22597,N_29354);
xor U35231 (N_35231,N_27113,N_23129);
or U35232 (N_35232,N_29919,N_28769);
or U35233 (N_35233,N_27851,N_28941);
nor U35234 (N_35234,N_27110,N_20991);
or U35235 (N_35235,N_23630,N_20882);
xor U35236 (N_35236,N_24481,N_28168);
and U35237 (N_35237,N_29177,N_25557);
nor U35238 (N_35238,N_28771,N_25598);
or U35239 (N_35239,N_25784,N_21249);
or U35240 (N_35240,N_26751,N_29520);
nor U35241 (N_35241,N_26773,N_22182);
or U35242 (N_35242,N_27201,N_27453);
nand U35243 (N_35243,N_25442,N_22621);
nand U35244 (N_35244,N_26563,N_28198);
or U35245 (N_35245,N_21900,N_25800);
nand U35246 (N_35246,N_25781,N_24785);
nand U35247 (N_35247,N_24181,N_23154);
and U35248 (N_35248,N_21554,N_23451);
and U35249 (N_35249,N_29207,N_28575);
or U35250 (N_35250,N_24272,N_24713);
nand U35251 (N_35251,N_26256,N_20560);
nor U35252 (N_35252,N_26717,N_20217);
nand U35253 (N_35253,N_24903,N_26815);
and U35254 (N_35254,N_20671,N_27849);
or U35255 (N_35255,N_22075,N_24322);
xnor U35256 (N_35256,N_26479,N_20862);
and U35257 (N_35257,N_24071,N_21782);
and U35258 (N_35258,N_29024,N_23663);
nor U35259 (N_35259,N_27809,N_29581);
xnor U35260 (N_35260,N_24858,N_20257);
xor U35261 (N_35261,N_20737,N_28983);
nor U35262 (N_35262,N_24642,N_21231);
xor U35263 (N_35263,N_20875,N_26305);
and U35264 (N_35264,N_22293,N_22097);
and U35265 (N_35265,N_23757,N_27484);
or U35266 (N_35266,N_28215,N_24449);
or U35267 (N_35267,N_25080,N_26090);
nor U35268 (N_35268,N_20071,N_29102);
nand U35269 (N_35269,N_24872,N_25978);
xnor U35270 (N_35270,N_24113,N_20041);
or U35271 (N_35271,N_27881,N_26074);
nor U35272 (N_35272,N_23143,N_21982);
xnor U35273 (N_35273,N_29887,N_24008);
nand U35274 (N_35274,N_28511,N_21764);
and U35275 (N_35275,N_29913,N_26169);
and U35276 (N_35276,N_26957,N_21062);
or U35277 (N_35277,N_26381,N_29453);
nor U35278 (N_35278,N_27980,N_22366);
nand U35279 (N_35279,N_28835,N_26776);
and U35280 (N_35280,N_23593,N_27930);
nand U35281 (N_35281,N_28276,N_24670);
or U35282 (N_35282,N_20815,N_25354);
or U35283 (N_35283,N_26192,N_20826);
or U35284 (N_35284,N_26144,N_21665);
xnor U35285 (N_35285,N_21195,N_29032);
nand U35286 (N_35286,N_25560,N_28997);
or U35287 (N_35287,N_25532,N_22663);
nor U35288 (N_35288,N_28792,N_27198);
xnor U35289 (N_35289,N_23951,N_21953);
or U35290 (N_35290,N_24480,N_22491);
and U35291 (N_35291,N_29177,N_25767);
nor U35292 (N_35292,N_21382,N_23827);
xor U35293 (N_35293,N_26514,N_20432);
xor U35294 (N_35294,N_21855,N_27365);
xor U35295 (N_35295,N_22400,N_23494);
and U35296 (N_35296,N_28504,N_29112);
xor U35297 (N_35297,N_22755,N_25131);
or U35298 (N_35298,N_24354,N_23229);
or U35299 (N_35299,N_25434,N_29299);
nand U35300 (N_35300,N_27591,N_20204);
and U35301 (N_35301,N_22168,N_25579);
xnor U35302 (N_35302,N_20430,N_27907);
nor U35303 (N_35303,N_22375,N_24020);
and U35304 (N_35304,N_21560,N_27144);
nor U35305 (N_35305,N_22821,N_21300);
xor U35306 (N_35306,N_28372,N_25179);
or U35307 (N_35307,N_26638,N_27425);
nand U35308 (N_35308,N_22634,N_26630);
xor U35309 (N_35309,N_27900,N_20614);
and U35310 (N_35310,N_22248,N_28147);
xor U35311 (N_35311,N_20890,N_22112);
or U35312 (N_35312,N_23425,N_24497);
nor U35313 (N_35313,N_25043,N_25178);
nand U35314 (N_35314,N_29677,N_28970);
and U35315 (N_35315,N_23612,N_27877);
xor U35316 (N_35316,N_29211,N_26251);
or U35317 (N_35317,N_25686,N_20868);
nor U35318 (N_35318,N_24078,N_23224);
and U35319 (N_35319,N_21097,N_21485);
and U35320 (N_35320,N_29078,N_20269);
and U35321 (N_35321,N_26064,N_29587);
xor U35322 (N_35322,N_25174,N_22239);
and U35323 (N_35323,N_27216,N_25709);
xor U35324 (N_35324,N_24078,N_25979);
nor U35325 (N_35325,N_27654,N_27338);
and U35326 (N_35326,N_25544,N_25223);
nand U35327 (N_35327,N_20663,N_23884);
or U35328 (N_35328,N_22120,N_22721);
and U35329 (N_35329,N_23641,N_25659);
or U35330 (N_35330,N_27594,N_25242);
xnor U35331 (N_35331,N_24134,N_21013);
or U35332 (N_35332,N_29173,N_24037);
xor U35333 (N_35333,N_21936,N_29939);
and U35334 (N_35334,N_21692,N_20236);
xor U35335 (N_35335,N_20294,N_20157);
xor U35336 (N_35336,N_20185,N_20850);
xor U35337 (N_35337,N_29634,N_27920);
and U35338 (N_35338,N_29026,N_20506);
nor U35339 (N_35339,N_26785,N_23693);
nand U35340 (N_35340,N_22325,N_29967);
or U35341 (N_35341,N_24459,N_20948);
nand U35342 (N_35342,N_23870,N_21775);
xor U35343 (N_35343,N_23108,N_25792);
nor U35344 (N_35344,N_20348,N_27988);
nor U35345 (N_35345,N_21264,N_23307);
and U35346 (N_35346,N_26250,N_29320);
xnor U35347 (N_35347,N_20026,N_24703);
or U35348 (N_35348,N_29506,N_29348);
xnor U35349 (N_35349,N_25810,N_28761);
and U35350 (N_35350,N_24295,N_26743);
or U35351 (N_35351,N_21589,N_24192);
nor U35352 (N_35352,N_25627,N_22022);
and U35353 (N_35353,N_23865,N_23202);
nand U35354 (N_35354,N_28201,N_29068);
and U35355 (N_35355,N_20913,N_28689);
and U35356 (N_35356,N_20593,N_29934);
or U35357 (N_35357,N_26353,N_28492);
nor U35358 (N_35358,N_25660,N_24883);
and U35359 (N_35359,N_27445,N_28052);
or U35360 (N_35360,N_29464,N_24511);
nand U35361 (N_35361,N_28503,N_20537);
nor U35362 (N_35362,N_29623,N_22623);
xor U35363 (N_35363,N_23407,N_21173);
or U35364 (N_35364,N_24652,N_20503);
xnor U35365 (N_35365,N_21491,N_29949);
xnor U35366 (N_35366,N_27332,N_25133);
and U35367 (N_35367,N_26709,N_23833);
and U35368 (N_35368,N_29233,N_20442);
or U35369 (N_35369,N_29371,N_28607);
nor U35370 (N_35370,N_24387,N_27210);
xor U35371 (N_35371,N_24758,N_25884);
nor U35372 (N_35372,N_21008,N_28587);
nand U35373 (N_35373,N_26744,N_26739);
xnor U35374 (N_35374,N_21368,N_23647);
xor U35375 (N_35375,N_29044,N_28126);
nor U35376 (N_35376,N_22541,N_20647);
nand U35377 (N_35377,N_24775,N_21976);
or U35378 (N_35378,N_20965,N_24681);
nor U35379 (N_35379,N_28407,N_23410);
xor U35380 (N_35380,N_29865,N_25150);
nand U35381 (N_35381,N_27135,N_28918);
xor U35382 (N_35382,N_23673,N_20074);
or U35383 (N_35383,N_27342,N_29576);
xnor U35384 (N_35384,N_27069,N_29917);
xor U35385 (N_35385,N_29413,N_29780);
or U35386 (N_35386,N_22294,N_21453);
nor U35387 (N_35387,N_28044,N_23813);
and U35388 (N_35388,N_24741,N_24996);
or U35389 (N_35389,N_24094,N_22901);
and U35390 (N_35390,N_26308,N_20219);
nand U35391 (N_35391,N_23123,N_23881);
xnor U35392 (N_35392,N_22003,N_20753);
nor U35393 (N_35393,N_26343,N_20457);
or U35394 (N_35394,N_21477,N_21853);
nand U35395 (N_35395,N_21001,N_27187);
xor U35396 (N_35396,N_26132,N_24526);
nor U35397 (N_35397,N_22036,N_25680);
and U35398 (N_35398,N_29765,N_28030);
nor U35399 (N_35399,N_21985,N_23444);
nor U35400 (N_35400,N_25658,N_23310);
or U35401 (N_35401,N_20115,N_21967);
xor U35402 (N_35402,N_23816,N_25045);
or U35403 (N_35403,N_27038,N_21887);
xnor U35404 (N_35404,N_22323,N_26800);
or U35405 (N_35405,N_23207,N_27312);
or U35406 (N_35406,N_23570,N_22011);
nor U35407 (N_35407,N_23733,N_28701);
xnor U35408 (N_35408,N_24562,N_21840);
xor U35409 (N_35409,N_29871,N_25738);
nand U35410 (N_35410,N_20404,N_24422);
or U35411 (N_35411,N_20447,N_27241);
or U35412 (N_35412,N_24940,N_21442);
and U35413 (N_35413,N_29836,N_20256);
or U35414 (N_35414,N_24980,N_23516);
xnor U35415 (N_35415,N_29399,N_21904);
nor U35416 (N_35416,N_27999,N_27136);
xor U35417 (N_35417,N_26654,N_21085);
xnor U35418 (N_35418,N_21008,N_24056);
and U35419 (N_35419,N_20016,N_25334);
nor U35420 (N_35420,N_22153,N_22025);
nand U35421 (N_35421,N_22796,N_22871);
and U35422 (N_35422,N_24080,N_26039);
nor U35423 (N_35423,N_25310,N_26631);
or U35424 (N_35424,N_23565,N_29854);
xor U35425 (N_35425,N_22787,N_27489);
nor U35426 (N_35426,N_26092,N_28900);
and U35427 (N_35427,N_24009,N_25582);
nor U35428 (N_35428,N_27136,N_27335);
nor U35429 (N_35429,N_21679,N_24872);
xor U35430 (N_35430,N_26284,N_27828);
nor U35431 (N_35431,N_20110,N_25326);
xnor U35432 (N_35432,N_22287,N_21136);
xnor U35433 (N_35433,N_29357,N_28176);
and U35434 (N_35434,N_22318,N_26000);
or U35435 (N_35435,N_24561,N_20287);
and U35436 (N_35436,N_29110,N_22493);
xor U35437 (N_35437,N_26998,N_29038);
nand U35438 (N_35438,N_21719,N_21828);
nor U35439 (N_35439,N_26795,N_22293);
and U35440 (N_35440,N_25576,N_22592);
nor U35441 (N_35441,N_24582,N_22595);
nand U35442 (N_35442,N_21796,N_29272);
and U35443 (N_35443,N_20910,N_23532);
or U35444 (N_35444,N_29435,N_29120);
and U35445 (N_35445,N_27662,N_25359);
nor U35446 (N_35446,N_20865,N_20260);
or U35447 (N_35447,N_21812,N_20097);
or U35448 (N_35448,N_25126,N_25691);
xnor U35449 (N_35449,N_26697,N_28243);
and U35450 (N_35450,N_20517,N_25439);
xnor U35451 (N_35451,N_29367,N_23532);
nand U35452 (N_35452,N_21683,N_27823);
nand U35453 (N_35453,N_28855,N_22500);
and U35454 (N_35454,N_28457,N_29401);
and U35455 (N_35455,N_23290,N_20677);
and U35456 (N_35456,N_23734,N_27169);
xnor U35457 (N_35457,N_20054,N_26596);
and U35458 (N_35458,N_29889,N_20066);
and U35459 (N_35459,N_25628,N_21321);
or U35460 (N_35460,N_28485,N_25772);
or U35461 (N_35461,N_21674,N_24653);
xor U35462 (N_35462,N_26848,N_28385);
xor U35463 (N_35463,N_22077,N_25580);
or U35464 (N_35464,N_20391,N_25602);
or U35465 (N_35465,N_24785,N_28222);
nand U35466 (N_35466,N_27301,N_20633);
and U35467 (N_35467,N_24040,N_24057);
xnor U35468 (N_35468,N_25872,N_21947);
nand U35469 (N_35469,N_26923,N_29403);
or U35470 (N_35470,N_24028,N_25816);
and U35471 (N_35471,N_27366,N_20462);
nor U35472 (N_35472,N_21692,N_28505);
and U35473 (N_35473,N_27897,N_26185);
or U35474 (N_35474,N_21614,N_28592);
nand U35475 (N_35475,N_25093,N_29831);
or U35476 (N_35476,N_23780,N_25969);
and U35477 (N_35477,N_22262,N_20141);
nand U35478 (N_35478,N_23278,N_27982);
xor U35479 (N_35479,N_25596,N_24687);
xor U35480 (N_35480,N_26414,N_22783);
xor U35481 (N_35481,N_28924,N_22413);
nor U35482 (N_35482,N_21688,N_21090);
and U35483 (N_35483,N_24331,N_20067);
or U35484 (N_35484,N_21211,N_25451);
nand U35485 (N_35485,N_28339,N_20721);
nor U35486 (N_35486,N_28585,N_20877);
nor U35487 (N_35487,N_25114,N_29595);
nand U35488 (N_35488,N_28700,N_26069);
xor U35489 (N_35489,N_24658,N_24656);
or U35490 (N_35490,N_21286,N_26231);
nor U35491 (N_35491,N_29400,N_23772);
nor U35492 (N_35492,N_26724,N_26990);
xnor U35493 (N_35493,N_29779,N_21523);
and U35494 (N_35494,N_23930,N_21895);
or U35495 (N_35495,N_22584,N_27749);
nand U35496 (N_35496,N_24651,N_22438);
xor U35497 (N_35497,N_28698,N_22818);
nor U35498 (N_35498,N_29700,N_20387);
and U35499 (N_35499,N_20829,N_26099);
and U35500 (N_35500,N_24471,N_25525);
or U35501 (N_35501,N_24066,N_20550);
nand U35502 (N_35502,N_27141,N_28339);
xnor U35503 (N_35503,N_29535,N_27528);
and U35504 (N_35504,N_26168,N_21522);
or U35505 (N_35505,N_20893,N_25345);
nand U35506 (N_35506,N_21628,N_22837);
xnor U35507 (N_35507,N_29842,N_21658);
nand U35508 (N_35508,N_27149,N_28079);
and U35509 (N_35509,N_24084,N_21954);
or U35510 (N_35510,N_28464,N_24359);
nand U35511 (N_35511,N_25472,N_20473);
or U35512 (N_35512,N_28232,N_25070);
xnor U35513 (N_35513,N_21572,N_20561);
and U35514 (N_35514,N_29785,N_23682);
nor U35515 (N_35515,N_23039,N_28510);
xnor U35516 (N_35516,N_20738,N_21897);
or U35517 (N_35517,N_25606,N_29636);
xor U35518 (N_35518,N_20780,N_29575);
xor U35519 (N_35519,N_27029,N_24963);
nor U35520 (N_35520,N_26372,N_24065);
xor U35521 (N_35521,N_27243,N_29595);
or U35522 (N_35522,N_20875,N_24164);
nor U35523 (N_35523,N_22951,N_23380);
nor U35524 (N_35524,N_22935,N_25163);
and U35525 (N_35525,N_21478,N_27849);
nor U35526 (N_35526,N_25328,N_23872);
nand U35527 (N_35527,N_20173,N_20497);
xnor U35528 (N_35528,N_26199,N_27383);
xor U35529 (N_35529,N_27530,N_20300);
or U35530 (N_35530,N_29871,N_24885);
or U35531 (N_35531,N_25196,N_29955);
nand U35532 (N_35532,N_23056,N_21179);
xor U35533 (N_35533,N_25889,N_20711);
and U35534 (N_35534,N_28208,N_29718);
or U35535 (N_35535,N_23132,N_24188);
nor U35536 (N_35536,N_27211,N_28682);
nand U35537 (N_35537,N_22631,N_22177);
xnor U35538 (N_35538,N_22152,N_29263);
nand U35539 (N_35539,N_25532,N_20320);
nor U35540 (N_35540,N_25257,N_26223);
xor U35541 (N_35541,N_26545,N_27175);
xnor U35542 (N_35542,N_28360,N_25713);
nor U35543 (N_35543,N_27254,N_21453);
and U35544 (N_35544,N_23025,N_25382);
or U35545 (N_35545,N_29618,N_22186);
xor U35546 (N_35546,N_25201,N_20519);
nand U35547 (N_35547,N_20483,N_20136);
xor U35548 (N_35548,N_20723,N_22582);
nand U35549 (N_35549,N_24717,N_25686);
and U35550 (N_35550,N_20783,N_24144);
and U35551 (N_35551,N_24631,N_20507);
or U35552 (N_35552,N_28364,N_28264);
nand U35553 (N_35553,N_24337,N_28719);
and U35554 (N_35554,N_27326,N_27940);
or U35555 (N_35555,N_25936,N_26651);
or U35556 (N_35556,N_29333,N_22767);
nand U35557 (N_35557,N_25247,N_21655);
nor U35558 (N_35558,N_25544,N_26527);
and U35559 (N_35559,N_25820,N_21710);
or U35560 (N_35560,N_26604,N_27652);
nor U35561 (N_35561,N_22343,N_23110);
nand U35562 (N_35562,N_29994,N_28812);
or U35563 (N_35563,N_26461,N_28442);
or U35564 (N_35564,N_28997,N_26676);
nor U35565 (N_35565,N_24332,N_23200);
nor U35566 (N_35566,N_25313,N_21009);
xnor U35567 (N_35567,N_20793,N_24778);
nand U35568 (N_35568,N_27280,N_24100);
and U35569 (N_35569,N_24870,N_20053);
xor U35570 (N_35570,N_21220,N_21315);
xor U35571 (N_35571,N_25076,N_27070);
or U35572 (N_35572,N_20557,N_22340);
or U35573 (N_35573,N_20050,N_25901);
nand U35574 (N_35574,N_28065,N_20306);
or U35575 (N_35575,N_23129,N_26623);
nor U35576 (N_35576,N_23870,N_23177);
xor U35577 (N_35577,N_21709,N_21026);
xnor U35578 (N_35578,N_29945,N_26303);
xnor U35579 (N_35579,N_22561,N_29844);
and U35580 (N_35580,N_27648,N_23240);
nor U35581 (N_35581,N_26667,N_21377);
xnor U35582 (N_35582,N_20014,N_29923);
nand U35583 (N_35583,N_29455,N_21558);
xor U35584 (N_35584,N_22990,N_22181);
xnor U35585 (N_35585,N_25027,N_20010);
or U35586 (N_35586,N_26761,N_29828);
nor U35587 (N_35587,N_21339,N_23447);
nor U35588 (N_35588,N_23713,N_21258);
or U35589 (N_35589,N_25728,N_23218);
xnor U35590 (N_35590,N_29436,N_20666);
nand U35591 (N_35591,N_24433,N_29004);
and U35592 (N_35592,N_20632,N_28037);
or U35593 (N_35593,N_23233,N_21313);
xor U35594 (N_35594,N_29395,N_22172);
and U35595 (N_35595,N_26899,N_25757);
nand U35596 (N_35596,N_21210,N_24888);
nor U35597 (N_35597,N_24415,N_29868);
and U35598 (N_35598,N_28910,N_26258);
xor U35599 (N_35599,N_28330,N_25080);
and U35600 (N_35600,N_27529,N_23561);
or U35601 (N_35601,N_29470,N_29879);
and U35602 (N_35602,N_23402,N_24234);
or U35603 (N_35603,N_27600,N_21798);
and U35604 (N_35604,N_26914,N_20164);
and U35605 (N_35605,N_27930,N_25303);
or U35606 (N_35606,N_26387,N_20882);
nor U35607 (N_35607,N_28479,N_24594);
nor U35608 (N_35608,N_20746,N_22003);
and U35609 (N_35609,N_21869,N_20299);
xnor U35610 (N_35610,N_24341,N_26897);
nor U35611 (N_35611,N_25636,N_20624);
nand U35612 (N_35612,N_27457,N_20288);
and U35613 (N_35613,N_21332,N_24859);
nor U35614 (N_35614,N_22027,N_29467);
and U35615 (N_35615,N_27878,N_27023);
nor U35616 (N_35616,N_29434,N_28822);
and U35617 (N_35617,N_26988,N_23920);
nor U35618 (N_35618,N_25222,N_29606);
or U35619 (N_35619,N_29638,N_21671);
or U35620 (N_35620,N_21800,N_29926);
nand U35621 (N_35621,N_28261,N_23702);
xnor U35622 (N_35622,N_21166,N_29857);
nand U35623 (N_35623,N_27485,N_23342);
or U35624 (N_35624,N_24432,N_29601);
and U35625 (N_35625,N_24099,N_27847);
nor U35626 (N_35626,N_26467,N_27890);
nand U35627 (N_35627,N_28712,N_23606);
nand U35628 (N_35628,N_21876,N_20421);
nor U35629 (N_35629,N_28755,N_23866);
nor U35630 (N_35630,N_21719,N_27082);
nor U35631 (N_35631,N_22910,N_29498);
nor U35632 (N_35632,N_26549,N_26288);
nor U35633 (N_35633,N_26028,N_26218);
xnor U35634 (N_35634,N_25499,N_28351);
and U35635 (N_35635,N_20172,N_23919);
nand U35636 (N_35636,N_25280,N_20830);
xor U35637 (N_35637,N_27462,N_20799);
or U35638 (N_35638,N_23466,N_24460);
nor U35639 (N_35639,N_27702,N_21624);
or U35640 (N_35640,N_29382,N_25059);
nor U35641 (N_35641,N_28630,N_29831);
xor U35642 (N_35642,N_20508,N_29919);
nand U35643 (N_35643,N_26518,N_29708);
or U35644 (N_35644,N_29742,N_20406);
or U35645 (N_35645,N_23630,N_27795);
or U35646 (N_35646,N_21224,N_28626);
xnor U35647 (N_35647,N_28368,N_24370);
or U35648 (N_35648,N_27543,N_20984);
nor U35649 (N_35649,N_25534,N_23780);
or U35650 (N_35650,N_23487,N_21534);
and U35651 (N_35651,N_27133,N_21533);
xor U35652 (N_35652,N_26963,N_22535);
nor U35653 (N_35653,N_27938,N_22191);
nand U35654 (N_35654,N_20419,N_24671);
nor U35655 (N_35655,N_27111,N_24391);
nand U35656 (N_35656,N_25497,N_25828);
nor U35657 (N_35657,N_27887,N_25573);
nor U35658 (N_35658,N_20550,N_24152);
xnor U35659 (N_35659,N_28051,N_20517);
nor U35660 (N_35660,N_20360,N_20517);
and U35661 (N_35661,N_25875,N_25164);
nor U35662 (N_35662,N_28051,N_26742);
nand U35663 (N_35663,N_27041,N_26451);
or U35664 (N_35664,N_29858,N_25043);
or U35665 (N_35665,N_24890,N_27499);
or U35666 (N_35666,N_22002,N_26085);
or U35667 (N_35667,N_25500,N_26490);
xnor U35668 (N_35668,N_28862,N_20713);
and U35669 (N_35669,N_24259,N_23988);
nor U35670 (N_35670,N_20832,N_28790);
or U35671 (N_35671,N_20679,N_23296);
nor U35672 (N_35672,N_28380,N_28603);
and U35673 (N_35673,N_29860,N_23279);
or U35674 (N_35674,N_20244,N_20320);
or U35675 (N_35675,N_22410,N_26894);
nand U35676 (N_35676,N_21306,N_27189);
or U35677 (N_35677,N_25603,N_25574);
nor U35678 (N_35678,N_20218,N_27754);
or U35679 (N_35679,N_28318,N_29984);
nand U35680 (N_35680,N_23141,N_21649);
nand U35681 (N_35681,N_24157,N_20812);
xor U35682 (N_35682,N_20597,N_26134);
nand U35683 (N_35683,N_25755,N_24551);
nor U35684 (N_35684,N_24178,N_20631);
nand U35685 (N_35685,N_27329,N_22385);
nand U35686 (N_35686,N_27669,N_29995);
xnor U35687 (N_35687,N_29496,N_22274);
nor U35688 (N_35688,N_25527,N_23519);
xnor U35689 (N_35689,N_26294,N_20523);
nor U35690 (N_35690,N_23160,N_20136);
xnor U35691 (N_35691,N_29205,N_28604);
and U35692 (N_35692,N_23176,N_23307);
nand U35693 (N_35693,N_21432,N_23495);
and U35694 (N_35694,N_23251,N_28517);
nor U35695 (N_35695,N_22038,N_27705);
xor U35696 (N_35696,N_20763,N_21703);
nand U35697 (N_35697,N_24438,N_28533);
nor U35698 (N_35698,N_25467,N_26115);
nor U35699 (N_35699,N_29584,N_27994);
and U35700 (N_35700,N_20891,N_29521);
and U35701 (N_35701,N_27757,N_24357);
or U35702 (N_35702,N_23452,N_25398);
nand U35703 (N_35703,N_23605,N_26810);
xor U35704 (N_35704,N_22143,N_23001);
nand U35705 (N_35705,N_24266,N_23851);
nand U35706 (N_35706,N_24143,N_24162);
or U35707 (N_35707,N_26777,N_26416);
xnor U35708 (N_35708,N_28630,N_28151);
or U35709 (N_35709,N_20466,N_20842);
nor U35710 (N_35710,N_29632,N_29638);
xor U35711 (N_35711,N_24331,N_27171);
nand U35712 (N_35712,N_21774,N_25450);
or U35713 (N_35713,N_21015,N_24432);
nor U35714 (N_35714,N_24692,N_24960);
nand U35715 (N_35715,N_23543,N_28945);
nand U35716 (N_35716,N_22377,N_21318);
and U35717 (N_35717,N_22282,N_26185);
nand U35718 (N_35718,N_20040,N_25227);
nor U35719 (N_35719,N_24905,N_27718);
nor U35720 (N_35720,N_27184,N_25091);
nand U35721 (N_35721,N_28777,N_23977);
xnor U35722 (N_35722,N_24313,N_29832);
nand U35723 (N_35723,N_21652,N_27319);
nor U35724 (N_35724,N_28951,N_27246);
xor U35725 (N_35725,N_23872,N_21126);
nor U35726 (N_35726,N_26260,N_27726);
or U35727 (N_35727,N_22371,N_29965);
nor U35728 (N_35728,N_22206,N_24808);
xor U35729 (N_35729,N_29394,N_24067);
or U35730 (N_35730,N_25355,N_21910);
nor U35731 (N_35731,N_22058,N_20414);
or U35732 (N_35732,N_23448,N_23967);
nand U35733 (N_35733,N_24883,N_27762);
nor U35734 (N_35734,N_25646,N_29979);
xnor U35735 (N_35735,N_28119,N_23804);
nand U35736 (N_35736,N_29864,N_27791);
or U35737 (N_35737,N_28317,N_26321);
xnor U35738 (N_35738,N_26898,N_24652);
nor U35739 (N_35739,N_28807,N_24773);
or U35740 (N_35740,N_21849,N_26579);
nand U35741 (N_35741,N_29383,N_20698);
and U35742 (N_35742,N_21047,N_27381);
nor U35743 (N_35743,N_23009,N_20845);
and U35744 (N_35744,N_25022,N_20277);
xnor U35745 (N_35745,N_25171,N_24786);
nand U35746 (N_35746,N_26657,N_23416);
xor U35747 (N_35747,N_24934,N_26848);
nand U35748 (N_35748,N_26730,N_24123);
xnor U35749 (N_35749,N_24734,N_25893);
xnor U35750 (N_35750,N_28313,N_24066);
nand U35751 (N_35751,N_22783,N_20014);
xor U35752 (N_35752,N_28496,N_22608);
nand U35753 (N_35753,N_28154,N_26356);
nand U35754 (N_35754,N_29520,N_28281);
nand U35755 (N_35755,N_21576,N_23051);
nand U35756 (N_35756,N_24291,N_22998);
nand U35757 (N_35757,N_26541,N_26201);
nand U35758 (N_35758,N_23949,N_25747);
xnor U35759 (N_35759,N_20282,N_26442);
or U35760 (N_35760,N_27124,N_23597);
and U35761 (N_35761,N_28877,N_24717);
nand U35762 (N_35762,N_27690,N_29698);
nand U35763 (N_35763,N_29197,N_22474);
and U35764 (N_35764,N_21179,N_29807);
xnor U35765 (N_35765,N_24125,N_25782);
or U35766 (N_35766,N_23024,N_28464);
xor U35767 (N_35767,N_24729,N_20068);
and U35768 (N_35768,N_24065,N_27305);
nand U35769 (N_35769,N_26541,N_20416);
xor U35770 (N_35770,N_26636,N_20439);
xor U35771 (N_35771,N_23154,N_28756);
xnor U35772 (N_35772,N_22078,N_26492);
and U35773 (N_35773,N_25428,N_28767);
nand U35774 (N_35774,N_21236,N_26235);
nand U35775 (N_35775,N_24033,N_26834);
or U35776 (N_35776,N_22209,N_24816);
and U35777 (N_35777,N_21935,N_20743);
and U35778 (N_35778,N_29860,N_20490);
xnor U35779 (N_35779,N_23416,N_21958);
or U35780 (N_35780,N_21984,N_20120);
nand U35781 (N_35781,N_29666,N_21665);
nand U35782 (N_35782,N_29081,N_20471);
or U35783 (N_35783,N_24384,N_22256);
xnor U35784 (N_35784,N_29936,N_21479);
nor U35785 (N_35785,N_28074,N_28305);
or U35786 (N_35786,N_25220,N_29361);
and U35787 (N_35787,N_23364,N_24248);
or U35788 (N_35788,N_28752,N_26817);
xor U35789 (N_35789,N_27276,N_29652);
xnor U35790 (N_35790,N_23251,N_26853);
nand U35791 (N_35791,N_22419,N_29710);
nand U35792 (N_35792,N_21328,N_20142);
xnor U35793 (N_35793,N_25813,N_22514);
and U35794 (N_35794,N_27958,N_21346);
nand U35795 (N_35795,N_28532,N_24839);
nor U35796 (N_35796,N_27513,N_24714);
nor U35797 (N_35797,N_23041,N_28730);
and U35798 (N_35798,N_22516,N_26826);
xnor U35799 (N_35799,N_25238,N_23545);
and U35800 (N_35800,N_21532,N_29626);
nand U35801 (N_35801,N_26893,N_25619);
and U35802 (N_35802,N_21625,N_22203);
nor U35803 (N_35803,N_28642,N_25643);
and U35804 (N_35804,N_23075,N_24802);
and U35805 (N_35805,N_28365,N_27953);
nand U35806 (N_35806,N_21012,N_24255);
xor U35807 (N_35807,N_27337,N_26528);
nand U35808 (N_35808,N_29169,N_29598);
nand U35809 (N_35809,N_27909,N_20222);
or U35810 (N_35810,N_22701,N_28973);
or U35811 (N_35811,N_21284,N_24675);
xnor U35812 (N_35812,N_20043,N_24518);
xor U35813 (N_35813,N_26966,N_23257);
nand U35814 (N_35814,N_24480,N_21418);
or U35815 (N_35815,N_27324,N_20131);
xor U35816 (N_35816,N_21627,N_25229);
or U35817 (N_35817,N_21159,N_26861);
or U35818 (N_35818,N_29212,N_29073);
or U35819 (N_35819,N_26338,N_26657);
nand U35820 (N_35820,N_21785,N_20464);
nor U35821 (N_35821,N_20813,N_23127);
nor U35822 (N_35822,N_22006,N_23489);
nand U35823 (N_35823,N_27620,N_25504);
and U35824 (N_35824,N_21425,N_25535);
or U35825 (N_35825,N_25730,N_26519);
nor U35826 (N_35826,N_27236,N_28890);
xnor U35827 (N_35827,N_29786,N_23906);
nor U35828 (N_35828,N_25522,N_23065);
xor U35829 (N_35829,N_24780,N_24547);
and U35830 (N_35830,N_27624,N_22518);
nor U35831 (N_35831,N_21423,N_22747);
xor U35832 (N_35832,N_24153,N_24836);
xor U35833 (N_35833,N_27269,N_29892);
nor U35834 (N_35834,N_28765,N_25504);
or U35835 (N_35835,N_26198,N_28542);
xor U35836 (N_35836,N_27963,N_24965);
xnor U35837 (N_35837,N_28734,N_22987);
nand U35838 (N_35838,N_22849,N_20492);
or U35839 (N_35839,N_26426,N_29880);
xor U35840 (N_35840,N_21051,N_22469);
or U35841 (N_35841,N_20354,N_28186);
nand U35842 (N_35842,N_20080,N_20625);
nor U35843 (N_35843,N_20305,N_23971);
xnor U35844 (N_35844,N_29527,N_25601);
nand U35845 (N_35845,N_21740,N_24450);
nand U35846 (N_35846,N_24768,N_29047);
or U35847 (N_35847,N_26166,N_23668);
xor U35848 (N_35848,N_20151,N_23208);
nand U35849 (N_35849,N_20339,N_27774);
or U35850 (N_35850,N_27498,N_21609);
xor U35851 (N_35851,N_20543,N_28103);
or U35852 (N_35852,N_23167,N_26669);
nand U35853 (N_35853,N_25939,N_21442);
nand U35854 (N_35854,N_22219,N_20599);
or U35855 (N_35855,N_27494,N_20208);
and U35856 (N_35856,N_27860,N_20550);
nor U35857 (N_35857,N_22763,N_21952);
nor U35858 (N_35858,N_29057,N_28224);
and U35859 (N_35859,N_28590,N_21907);
nand U35860 (N_35860,N_21676,N_23472);
nand U35861 (N_35861,N_27397,N_21831);
nand U35862 (N_35862,N_28258,N_24685);
and U35863 (N_35863,N_25460,N_26230);
xnor U35864 (N_35864,N_21247,N_24471);
and U35865 (N_35865,N_20914,N_27722);
or U35866 (N_35866,N_27850,N_21018);
or U35867 (N_35867,N_20364,N_25584);
or U35868 (N_35868,N_20874,N_22494);
xor U35869 (N_35869,N_26744,N_23132);
or U35870 (N_35870,N_29979,N_28599);
nor U35871 (N_35871,N_21261,N_21367);
xnor U35872 (N_35872,N_28495,N_27690);
and U35873 (N_35873,N_29233,N_22373);
nand U35874 (N_35874,N_26836,N_22006);
xnor U35875 (N_35875,N_23313,N_22634);
nor U35876 (N_35876,N_24760,N_24273);
nand U35877 (N_35877,N_21019,N_29201);
and U35878 (N_35878,N_25230,N_28781);
and U35879 (N_35879,N_29814,N_23479);
nor U35880 (N_35880,N_29356,N_25243);
nor U35881 (N_35881,N_22777,N_28635);
nor U35882 (N_35882,N_20989,N_29141);
xnor U35883 (N_35883,N_26978,N_25302);
or U35884 (N_35884,N_22288,N_27012);
nand U35885 (N_35885,N_29887,N_23910);
nand U35886 (N_35886,N_25692,N_26780);
xnor U35887 (N_35887,N_28606,N_23886);
nor U35888 (N_35888,N_29593,N_29851);
xor U35889 (N_35889,N_23076,N_23555);
xor U35890 (N_35890,N_29552,N_25305);
or U35891 (N_35891,N_29142,N_25244);
or U35892 (N_35892,N_24209,N_20865);
nor U35893 (N_35893,N_20047,N_21960);
or U35894 (N_35894,N_27996,N_22159);
nand U35895 (N_35895,N_23374,N_21102);
nor U35896 (N_35896,N_27513,N_26803);
and U35897 (N_35897,N_22316,N_25295);
xnor U35898 (N_35898,N_21573,N_21970);
xor U35899 (N_35899,N_20610,N_23394);
nand U35900 (N_35900,N_23012,N_25384);
nor U35901 (N_35901,N_21841,N_28535);
or U35902 (N_35902,N_29574,N_29232);
nor U35903 (N_35903,N_25811,N_22443);
xor U35904 (N_35904,N_25005,N_21232);
or U35905 (N_35905,N_20323,N_23421);
and U35906 (N_35906,N_25727,N_22821);
and U35907 (N_35907,N_22713,N_25453);
nand U35908 (N_35908,N_24755,N_26283);
or U35909 (N_35909,N_29877,N_26640);
and U35910 (N_35910,N_26525,N_28710);
nor U35911 (N_35911,N_28967,N_21863);
nand U35912 (N_35912,N_23138,N_25326);
nand U35913 (N_35913,N_21915,N_29097);
or U35914 (N_35914,N_22300,N_20658);
xor U35915 (N_35915,N_21060,N_28458);
or U35916 (N_35916,N_25036,N_20428);
nand U35917 (N_35917,N_26897,N_24977);
nand U35918 (N_35918,N_22321,N_26790);
or U35919 (N_35919,N_25873,N_29196);
nand U35920 (N_35920,N_23132,N_28430);
nand U35921 (N_35921,N_21191,N_29042);
nor U35922 (N_35922,N_21586,N_27888);
xnor U35923 (N_35923,N_20611,N_26091);
nand U35924 (N_35924,N_26588,N_20101);
or U35925 (N_35925,N_24095,N_25309);
xnor U35926 (N_35926,N_21327,N_22271);
xnor U35927 (N_35927,N_28090,N_27173);
xnor U35928 (N_35928,N_27639,N_22445);
xnor U35929 (N_35929,N_25181,N_27950);
nor U35930 (N_35930,N_22111,N_20773);
or U35931 (N_35931,N_22629,N_27180);
and U35932 (N_35932,N_21584,N_22331);
nor U35933 (N_35933,N_29204,N_21150);
or U35934 (N_35934,N_21289,N_20768);
and U35935 (N_35935,N_28258,N_27957);
nand U35936 (N_35936,N_23580,N_26944);
xnor U35937 (N_35937,N_26947,N_23947);
or U35938 (N_35938,N_25842,N_29293);
or U35939 (N_35939,N_23306,N_26767);
xor U35940 (N_35940,N_29728,N_23046);
nor U35941 (N_35941,N_25168,N_23099);
nor U35942 (N_35942,N_28696,N_29088);
xnor U35943 (N_35943,N_21281,N_26512);
xor U35944 (N_35944,N_26004,N_24073);
nand U35945 (N_35945,N_22964,N_24848);
xnor U35946 (N_35946,N_20921,N_24246);
xnor U35947 (N_35947,N_28556,N_27909);
nand U35948 (N_35948,N_28430,N_20477);
or U35949 (N_35949,N_22659,N_26271);
and U35950 (N_35950,N_26995,N_28460);
xor U35951 (N_35951,N_28072,N_28832);
xor U35952 (N_35952,N_24959,N_20989);
and U35953 (N_35953,N_22625,N_24558);
nand U35954 (N_35954,N_25478,N_23618);
and U35955 (N_35955,N_26854,N_26235);
xnor U35956 (N_35956,N_23291,N_25715);
and U35957 (N_35957,N_25020,N_22314);
or U35958 (N_35958,N_26822,N_27062);
or U35959 (N_35959,N_28739,N_28593);
nand U35960 (N_35960,N_24041,N_25192);
nor U35961 (N_35961,N_24053,N_27821);
and U35962 (N_35962,N_26306,N_22202);
nand U35963 (N_35963,N_29589,N_28683);
or U35964 (N_35964,N_22744,N_29220);
nand U35965 (N_35965,N_28283,N_26563);
and U35966 (N_35966,N_20539,N_21926);
nand U35967 (N_35967,N_21006,N_20299);
nand U35968 (N_35968,N_24255,N_21868);
nand U35969 (N_35969,N_26040,N_23898);
xor U35970 (N_35970,N_29461,N_25377);
and U35971 (N_35971,N_27620,N_22487);
xnor U35972 (N_35972,N_23714,N_29762);
or U35973 (N_35973,N_28712,N_26816);
and U35974 (N_35974,N_22314,N_27551);
nor U35975 (N_35975,N_29580,N_20715);
xnor U35976 (N_35976,N_21148,N_26987);
nand U35977 (N_35977,N_28388,N_22959);
nand U35978 (N_35978,N_26267,N_23926);
nor U35979 (N_35979,N_27248,N_23731);
nand U35980 (N_35980,N_22483,N_22167);
nand U35981 (N_35981,N_25134,N_28714);
and U35982 (N_35982,N_29713,N_27891);
nor U35983 (N_35983,N_22966,N_20793);
nand U35984 (N_35984,N_25271,N_23662);
xor U35985 (N_35985,N_27968,N_24709);
or U35986 (N_35986,N_26964,N_22863);
nor U35987 (N_35987,N_28229,N_23100);
nor U35988 (N_35988,N_28549,N_29770);
nand U35989 (N_35989,N_24908,N_21161);
and U35990 (N_35990,N_25237,N_20068);
nand U35991 (N_35991,N_20563,N_25107);
xnor U35992 (N_35992,N_28013,N_22912);
nor U35993 (N_35993,N_25871,N_22188);
xor U35994 (N_35994,N_27828,N_21259);
or U35995 (N_35995,N_26463,N_25751);
or U35996 (N_35996,N_29263,N_26893);
nand U35997 (N_35997,N_25129,N_23597);
nand U35998 (N_35998,N_26501,N_22828);
nand U35999 (N_35999,N_26063,N_28061);
nand U36000 (N_36000,N_20080,N_28762);
or U36001 (N_36001,N_21948,N_25942);
and U36002 (N_36002,N_21848,N_24279);
nor U36003 (N_36003,N_21254,N_28005);
and U36004 (N_36004,N_29267,N_26959);
xnor U36005 (N_36005,N_28047,N_23943);
nand U36006 (N_36006,N_26251,N_24028);
xnor U36007 (N_36007,N_29954,N_27105);
nor U36008 (N_36008,N_25878,N_20076);
and U36009 (N_36009,N_28050,N_27053);
and U36010 (N_36010,N_21507,N_21909);
and U36011 (N_36011,N_23973,N_28726);
xor U36012 (N_36012,N_20604,N_25357);
nor U36013 (N_36013,N_23227,N_21974);
xnor U36014 (N_36014,N_26116,N_20512);
or U36015 (N_36015,N_20964,N_28060);
or U36016 (N_36016,N_29135,N_20832);
xnor U36017 (N_36017,N_26318,N_20639);
nor U36018 (N_36018,N_29538,N_29643);
nand U36019 (N_36019,N_28237,N_20764);
and U36020 (N_36020,N_28380,N_20637);
xor U36021 (N_36021,N_24464,N_22635);
and U36022 (N_36022,N_21469,N_23322);
or U36023 (N_36023,N_25387,N_20597);
or U36024 (N_36024,N_26325,N_25815);
and U36025 (N_36025,N_29229,N_22488);
or U36026 (N_36026,N_24632,N_23960);
or U36027 (N_36027,N_21885,N_25744);
nor U36028 (N_36028,N_26844,N_21520);
and U36029 (N_36029,N_23869,N_20456);
nand U36030 (N_36030,N_26181,N_23321);
xor U36031 (N_36031,N_26517,N_22994);
or U36032 (N_36032,N_27036,N_29655);
or U36033 (N_36033,N_25422,N_29029);
and U36034 (N_36034,N_24474,N_26408);
nand U36035 (N_36035,N_25544,N_29713);
nand U36036 (N_36036,N_28298,N_20039);
nor U36037 (N_36037,N_24244,N_25041);
or U36038 (N_36038,N_24976,N_22876);
xnor U36039 (N_36039,N_23708,N_27263);
and U36040 (N_36040,N_22608,N_25025);
or U36041 (N_36041,N_20372,N_20100);
nand U36042 (N_36042,N_24811,N_23260);
and U36043 (N_36043,N_23034,N_22463);
nand U36044 (N_36044,N_29783,N_28969);
nor U36045 (N_36045,N_23047,N_28833);
xor U36046 (N_36046,N_25901,N_23856);
and U36047 (N_36047,N_27766,N_26588);
nor U36048 (N_36048,N_26372,N_29851);
xnor U36049 (N_36049,N_28478,N_22642);
xnor U36050 (N_36050,N_23197,N_28141);
nor U36051 (N_36051,N_22175,N_27393);
xnor U36052 (N_36052,N_24955,N_24234);
and U36053 (N_36053,N_24571,N_24569);
or U36054 (N_36054,N_26774,N_20064);
xor U36055 (N_36055,N_27125,N_22596);
nor U36056 (N_36056,N_29184,N_20607);
nor U36057 (N_36057,N_28804,N_20668);
xnor U36058 (N_36058,N_23261,N_28161);
or U36059 (N_36059,N_20067,N_22943);
and U36060 (N_36060,N_29953,N_25626);
or U36061 (N_36061,N_23237,N_29352);
nor U36062 (N_36062,N_26567,N_24728);
or U36063 (N_36063,N_26746,N_21636);
nand U36064 (N_36064,N_28704,N_28654);
nor U36065 (N_36065,N_27168,N_22728);
xor U36066 (N_36066,N_20153,N_21052);
nand U36067 (N_36067,N_22856,N_25665);
and U36068 (N_36068,N_22866,N_27147);
nor U36069 (N_36069,N_28723,N_27853);
or U36070 (N_36070,N_29112,N_21858);
or U36071 (N_36071,N_25460,N_29226);
or U36072 (N_36072,N_25669,N_24200);
xor U36073 (N_36073,N_22393,N_24491);
or U36074 (N_36074,N_20552,N_21336);
nor U36075 (N_36075,N_20959,N_29317);
nand U36076 (N_36076,N_25466,N_22485);
nand U36077 (N_36077,N_24559,N_22377);
xor U36078 (N_36078,N_27635,N_24102);
nor U36079 (N_36079,N_26448,N_23045);
nand U36080 (N_36080,N_27930,N_20331);
nor U36081 (N_36081,N_25031,N_22852);
nor U36082 (N_36082,N_20817,N_26236);
and U36083 (N_36083,N_28832,N_23088);
nand U36084 (N_36084,N_23336,N_27993);
or U36085 (N_36085,N_27628,N_23670);
xnor U36086 (N_36086,N_25328,N_22568);
nand U36087 (N_36087,N_27434,N_21932);
nor U36088 (N_36088,N_22201,N_28575);
xnor U36089 (N_36089,N_26055,N_26103);
nand U36090 (N_36090,N_27407,N_26525);
nand U36091 (N_36091,N_28000,N_26901);
nand U36092 (N_36092,N_26446,N_23031);
xor U36093 (N_36093,N_21722,N_27838);
nor U36094 (N_36094,N_24573,N_20777);
nand U36095 (N_36095,N_25219,N_20625);
nor U36096 (N_36096,N_24531,N_27864);
or U36097 (N_36097,N_27081,N_26902);
xor U36098 (N_36098,N_26799,N_27499);
and U36099 (N_36099,N_26501,N_20063);
or U36100 (N_36100,N_20564,N_29568);
xnor U36101 (N_36101,N_21098,N_20316);
nor U36102 (N_36102,N_21558,N_29010);
nand U36103 (N_36103,N_22601,N_23381);
xor U36104 (N_36104,N_23109,N_28930);
xnor U36105 (N_36105,N_27449,N_23753);
nor U36106 (N_36106,N_23570,N_20283);
nand U36107 (N_36107,N_29997,N_22782);
nor U36108 (N_36108,N_21543,N_20755);
and U36109 (N_36109,N_28555,N_24160);
and U36110 (N_36110,N_28040,N_24557);
nand U36111 (N_36111,N_29798,N_23476);
xor U36112 (N_36112,N_25639,N_21563);
and U36113 (N_36113,N_26637,N_29544);
nand U36114 (N_36114,N_28538,N_22279);
and U36115 (N_36115,N_22306,N_25678);
nor U36116 (N_36116,N_28863,N_28078);
or U36117 (N_36117,N_26630,N_25734);
nand U36118 (N_36118,N_20454,N_23922);
and U36119 (N_36119,N_29906,N_27203);
xor U36120 (N_36120,N_21569,N_21765);
nor U36121 (N_36121,N_27318,N_25052);
nor U36122 (N_36122,N_21431,N_22679);
or U36123 (N_36123,N_20437,N_21071);
or U36124 (N_36124,N_22683,N_22233);
and U36125 (N_36125,N_22302,N_29713);
and U36126 (N_36126,N_20695,N_20879);
nand U36127 (N_36127,N_21294,N_29509);
nand U36128 (N_36128,N_25494,N_26112);
nor U36129 (N_36129,N_28768,N_22857);
and U36130 (N_36130,N_27178,N_23644);
and U36131 (N_36131,N_26982,N_26453);
nand U36132 (N_36132,N_28955,N_26270);
and U36133 (N_36133,N_27155,N_25386);
and U36134 (N_36134,N_25377,N_29995);
xor U36135 (N_36135,N_27703,N_26513);
nor U36136 (N_36136,N_23048,N_29938);
nand U36137 (N_36137,N_23199,N_25639);
or U36138 (N_36138,N_21836,N_21543);
or U36139 (N_36139,N_22733,N_26064);
and U36140 (N_36140,N_21348,N_29509);
xor U36141 (N_36141,N_28191,N_23785);
nor U36142 (N_36142,N_29326,N_23185);
xnor U36143 (N_36143,N_25446,N_28595);
nand U36144 (N_36144,N_27060,N_24679);
or U36145 (N_36145,N_29974,N_21207);
nor U36146 (N_36146,N_29173,N_26243);
nor U36147 (N_36147,N_27575,N_24373);
and U36148 (N_36148,N_25316,N_24891);
and U36149 (N_36149,N_29431,N_21942);
nor U36150 (N_36150,N_26620,N_22990);
nor U36151 (N_36151,N_23225,N_22043);
nor U36152 (N_36152,N_29979,N_24142);
and U36153 (N_36153,N_24974,N_25360);
xor U36154 (N_36154,N_25579,N_22453);
and U36155 (N_36155,N_22224,N_27279);
xnor U36156 (N_36156,N_22373,N_22943);
xnor U36157 (N_36157,N_20469,N_29480);
xor U36158 (N_36158,N_28036,N_24317);
or U36159 (N_36159,N_25655,N_24719);
nor U36160 (N_36160,N_22776,N_26680);
or U36161 (N_36161,N_26694,N_26458);
and U36162 (N_36162,N_29122,N_28132);
and U36163 (N_36163,N_28568,N_23673);
nand U36164 (N_36164,N_21681,N_25110);
or U36165 (N_36165,N_26555,N_21842);
xnor U36166 (N_36166,N_21894,N_23551);
nand U36167 (N_36167,N_22148,N_24486);
nor U36168 (N_36168,N_26107,N_25559);
nand U36169 (N_36169,N_22525,N_27817);
xnor U36170 (N_36170,N_26178,N_27380);
xor U36171 (N_36171,N_24983,N_28119);
nand U36172 (N_36172,N_23986,N_24213);
and U36173 (N_36173,N_20305,N_25596);
xnor U36174 (N_36174,N_23417,N_28331);
nor U36175 (N_36175,N_27567,N_24555);
or U36176 (N_36176,N_21078,N_20575);
or U36177 (N_36177,N_21114,N_20074);
or U36178 (N_36178,N_24514,N_21350);
or U36179 (N_36179,N_21662,N_24354);
or U36180 (N_36180,N_28913,N_28577);
nand U36181 (N_36181,N_29252,N_27671);
and U36182 (N_36182,N_27654,N_21994);
xor U36183 (N_36183,N_23616,N_23022);
xor U36184 (N_36184,N_20772,N_29581);
xnor U36185 (N_36185,N_20337,N_27223);
or U36186 (N_36186,N_20768,N_28841);
or U36187 (N_36187,N_24351,N_24424);
xnor U36188 (N_36188,N_29691,N_28979);
xnor U36189 (N_36189,N_28961,N_25136);
and U36190 (N_36190,N_24002,N_25861);
xnor U36191 (N_36191,N_27196,N_22406);
xor U36192 (N_36192,N_21055,N_21957);
and U36193 (N_36193,N_22618,N_27931);
nand U36194 (N_36194,N_21463,N_25125);
nand U36195 (N_36195,N_27394,N_28905);
or U36196 (N_36196,N_29565,N_27459);
and U36197 (N_36197,N_28565,N_21806);
and U36198 (N_36198,N_23799,N_23985);
or U36199 (N_36199,N_20621,N_25984);
or U36200 (N_36200,N_28477,N_23533);
nand U36201 (N_36201,N_28555,N_25440);
nand U36202 (N_36202,N_20169,N_26151);
nor U36203 (N_36203,N_23755,N_27233);
and U36204 (N_36204,N_22168,N_23110);
nand U36205 (N_36205,N_25376,N_20645);
or U36206 (N_36206,N_26075,N_23339);
and U36207 (N_36207,N_28348,N_23628);
xnor U36208 (N_36208,N_20081,N_24984);
nand U36209 (N_36209,N_26880,N_28906);
xor U36210 (N_36210,N_22286,N_20334);
nor U36211 (N_36211,N_28589,N_29201);
xor U36212 (N_36212,N_21635,N_20815);
or U36213 (N_36213,N_20911,N_22842);
and U36214 (N_36214,N_29597,N_23977);
and U36215 (N_36215,N_25839,N_25802);
nand U36216 (N_36216,N_26718,N_20243);
nor U36217 (N_36217,N_25608,N_24410);
and U36218 (N_36218,N_23354,N_27521);
and U36219 (N_36219,N_21095,N_28099);
and U36220 (N_36220,N_21002,N_26503);
and U36221 (N_36221,N_22967,N_20072);
xnor U36222 (N_36222,N_24311,N_27799);
or U36223 (N_36223,N_27159,N_25092);
nor U36224 (N_36224,N_24988,N_20445);
and U36225 (N_36225,N_22421,N_24206);
or U36226 (N_36226,N_25760,N_24672);
or U36227 (N_36227,N_29252,N_26600);
nand U36228 (N_36228,N_27328,N_25613);
nor U36229 (N_36229,N_20687,N_27606);
xnor U36230 (N_36230,N_21625,N_20196);
and U36231 (N_36231,N_21686,N_25218);
xnor U36232 (N_36232,N_27885,N_24567);
nand U36233 (N_36233,N_28389,N_22318);
nand U36234 (N_36234,N_20063,N_23108);
nor U36235 (N_36235,N_21288,N_22781);
nand U36236 (N_36236,N_25829,N_25567);
and U36237 (N_36237,N_25943,N_24182);
and U36238 (N_36238,N_21552,N_25019);
nor U36239 (N_36239,N_24499,N_26703);
and U36240 (N_36240,N_26569,N_23424);
nand U36241 (N_36241,N_21419,N_25496);
nand U36242 (N_36242,N_23330,N_21999);
and U36243 (N_36243,N_22328,N_22792);
or U36244 (N_36244,N_22219,N_24067);
or U36245 (N_36245,N_25376,N_25068);
or U36246 (N_36246,N_20995,N_23860);
nor U36247 (N_36247,N_24569,N_21627);
xor U36248 (N_36248,N_23832,N_21756);
nand U36249 (N_36249,N_21890,N_26404);
and U36250 (N_36250,N_23184,N_26761);
and U36251 (N_36251,N_25295,N_24164);
nand U36252 (N_36252,N_21210,N_25666);
xor U36253 (N_36253,N_25621,N_28519);
nor U36254 (N_36254,N_20221,N_26529);
and U36255 (N_36255,N_24093,N_26586);
nor U36256 (N_36256,N_20756,N_22872);
xnor U36257 (N_36257,N_27363,N_29122);
or U36258 (N_36258,N_26517,N_24848);
and U36259 (N_36259,N_20891,N_26348);
nand U36260 (N_36260,N_22153,N_21397);
nor U36261 (N_36261,N_26428,N_29671);
and U36262 (N_36262,N_29517,N_26573);
xor U36263 (N_36263,N_20732,N_23808);
and U36264 (N_36264,N_22317,N_21108);
and U36265 (N_36265,N_20079,N_29198);
or U36266 (N_36266,N_21321,N_29421);
xnor U36267 (N_36267,N_23485,N_22459);
nand U36268 (N_36268,N_29123,N_25191);
nor U36269 (N_36269,N_25261,N_22085);
xor U36270 (N_36270,N_24530,N_21817);
xnor U36271 (N_36271,N_27529,N_22427);
xor U36272 (N_36272,N_28033,N_28870);
xnor U36273 (N_36273,N_22704,N_28145);
nor U36274 (N_36274,N_25531,N_25807);
and U36275 (N_36275,N_23620,N_24235);
nor U36276 (N_36276,N_27648,N_29663);
or U36277 (N_36277,N_20064,N_26439);
nor U36278 (N_36278,N_29277,N_26379);
nor U36279 (N_36279,N_21561,N_21265);
xnor U36280 (N_36280,N_26634,N_21419);
nand U36281 (N_36281,N_29033,N_20473);
nor U36282 (N_36282,N_27081,N_25699);
or U36283 (N_36283,N_29781,N_24583);
xor U36284 (N_36284,N_23367,N_27478);
and U36285 (N_36285,N_25483,N_21187);
nor U36286 (N_36286,N_26809,N_26068);
xnor U36287 (N_36287,N_22959,N_29534);
and U36288 (N_36288,N_24737,N_25839);
nand U36289 (N_36289,N_20814,N_28949);
xnor U36290 (N_36290,N_24135,N_20773);
nand U36291 (N_36291,N_22666,N_24197);
nand U36292 (N_36292,N_23594,N_24758);
and U36293 (N_36293,N_21928,N_27076);
and U36294 (N_36294,N_27594,N_29474);
nor U36295 (N_36295,N_21919,N_26079);
and U36296 (N_36296,N_27629,N_20787);
xor U36297 (N_36297,N_23858,N_23846);
or U36298 (N_36298,N_22731,N_25173);
nor U36299 (N_36299,N_26267,N_22358);
and U36300 (N_36300,N_25315,N_20851);
nor U36301 (N_36301,N_27875,N_28786);
nand U36302 (N_36302,N_20553,N_27455);
nor U36303 (N_36303,N_25622,N_23721);
nand U36304 (N_36304,N_27206,N_24005);
nor U36305 (N_36305,N_29782,N_28387);
and U36306 (N_36306,N_25112,N_28168);
nor U36307 (N_36307,N_21730,N_20748);
xnor U36308 (N_36308,N_22933,N_22562);
or U36309 (N_36309,N_21076,N_26573);
nor U36310 (N_36310,N_27642,N_21847);
or U36311 (N_36311,N_29143,N_26209);
or U36312 (N_36312,N_26878,N_22744);
or U36313 (N_36313,N_28259,N_24679);
nand U36314 (N_36314,N_22049,N_22749);
nand U36315 (N_36315,N_27829,N_24584);
xnor U36316 (N_36316,N_23279,N_25256);
nor U36317 (N_36317,N_24050,N_22102);
nor U36318 (N_36318,N_25068,N_24949);
xor U36319 (N_36319,N_20596,N_20144);
or U36320 (N_36320,N_28292,N_21542);
or U36321 (N_36321,N_21667,N_23150);
xor U36322 (N_36322,N_26908,N_28777);
and U36323 (N_36323,N_21550,N_27399);
nor U36324 (N_36324,N_29620,N_24333);
nand U36325 (N_36325,N_23551,N_29592);
and U36326 (N_36326,N_23867,N_20906);
xnor U36327 (N_36327,N_23604,N_24834);
or U36328 (N_36328,N_29352,N_26683);
nor U36329 (N_36329,N_23814,N_27644);
nand U36330 (N_36330,N_20026,N_22609);
nor U36331 (N_36331,N_21223,N_23758);
nand U36332 (N_36332,N_23428,N_25841);
nor U36333 (N_36333,N_24638,N_22288);
or U36334 (N_36334,N_21871,N_21844);
or U36335 (N_36335,N_22768,N_24945);
nor U36336 (N_36336,N_28485,N_24397);
nor U36337 (N_36337,N_27857,N_27629);
nor U36338 (N_36338,N_20645,N_22298);
or U36339 (N_36339,N_25076,N_20476);
nor U36340 (N_36340,N_23466,N_28824);
nor U36341 (N_36341,N_29226,N_28075);
or U36342 (N_36342,N_23611,N_26126);
nor U36343 (N_36343,N_23039,N_23628);
nand U36344 (N_36344,N_24853,N_25842);
and U36345 (N_36345,N_29158,N_26793);
or U36346 (N_36346,N_21812,N_21896);
nor U36347 (N_36347,N_27513,N_23733);
xnor U36348 (N_36348,N_25613,N_29730);
or U36349 (N_36349,N_20023,N_20709);
nor U36350 (N_36350,N_26996,N_24592);
or U36351 (N_36351,N_28367,N_22620);
xor U36352 (N_36352,N_29660,N_20722);
nand U36353 (N_36353,N_25849,N_25510);
nand U36354 (N_36354,N_28228,N_25755);
nand U36355 (N_36355,N_21395,N_25421);
or U36356 (N_36356,N_20197,N_24115);
or U36357 (N_36357,N_22125,N_28056);
nor U36358 (N_36358,N_26614,N_24529);
and U36359 (N_36359,N_23007,N_24356);
xnor U36360 (N_36360,N_21653,N_25642);
nand U36361 (N_36361,N_24806,N_27151);
nor U36362 (N_36362,N_24024,N_20459);
xnor U36363 (N_36363,N_24381,N_23430);
nand U36364 (N_36364,N_26443,N_26557);
nand U36365 (N_36365,N_20790,N_23260);
nor U36366 (N_36366,N_29431,N_23996);
or U36367 (N_36367,N_29930,N_24456);
xor U36368 (N_36368,N_24198,N_25811);
or U36369 (N_36369,N_21150,N_24583);
xor U36370 (N_36370,N_26847,N_26794);
and U36371 (N_36371,N_20582,N_24955);
nand U36372 (N_36372,N_20394,N_23403);
and U36373 (N_36373,N_24302,N_28166);
and U36374 (N_36374,N_24495,N_29487);
and U36375 (N_36375,N_23418,N_23785);
nand U36376 (N_36376,N_24506,N_25523);
or U36377 (N_36377,N_24107,N_22493);
xnor U36378 (N_36378,N_21258,N_25127);
nand U36379 (N_36379,N_23370,N_20620);
nor U36380 (N_36380,N_21781,N_21244);
or U36381 (N_36381,N_26609,N_28818);
xnor U36382 (N_36382,N_22814,N_24421);
xor U36383 (N_36383,N_20543,N_29171);
nor U36384 (N_36384,N_25772,N_20466);
or U36385 (N_36385,N_21368,N_20397);
nand U36386 (N_36386,N_29988,N_20605);
nor U36387 (N_36387,N_28102,N_27333);
nand U36388 (N_36388,N_27203,N_24193);
nand U36389 (N_36389,N_29144,N_25875);
and U36390 (N_36390,N_24948,N_28697);
xor U36391 (N_36391,N_29461,N_22795);
or U36392 (N_36392,N_22997,N_22945);
and U36393 (N_36393,N_24411,N_23278);
or U36394 (N_36394,N_20731,N_21129);
xor U36395 (N_36395,N_23462,N_22003);
and U36396 (N_36396,N_29887,N_22926);
and U36397 (N_36397,N_20793,N_20504);
nand U36398 (N_36398,N_27749,N_24280);
nand U36399 (N_36399,N_26047,N_28432);
xor U36400 (N_36400,N_28862,N_23053);
xnor U36401 (N_36401,N_27517,N_28229);
and U36402 (N_36402,N_22179,N_26922);
or U36403 (N_36403,N_27411,N_22603);
xor U36404 (N_36404,N_25201,N_20387);
nor U36405 (N_36405,N_20714,N_21291);
nor U36406 (N_36406,N_29626,N_23858);
or U36407 (N_36407,N_22524,N_29116);
nor U36408 (N_36408,N_20649,N_20136);
or U36409 (N_36409,N_24399,N_27706);
nor U36410 (N_36410,N_22247,N_28157);
nor U36411 (N_36411,N_27428,N_23450);
or U36412 (N_36412,N_22656,N_24102);
xor U36413 (N_36413,N_29484,N_26375);
and U36414 (N_36414,N_27591,N_22539);
nand U36415 (N_36415,N_24029,N_22030);
or U36416 (N_36416,N_21001,N_27583);
nand U36417 (N_36417,N_27746,N_24084);
nor U36418 (N_36418,N_28012,N_26644);
xor U36419 (N_36419,N_28447,N_24239);
nor U36420 (N_36420,N_28377,N_25666);
and U36421 (N_36421,N_25385,N_21426);
or U36422 (N_36422,N_25315,N_26963);
nor U36423 (N_36423,N_27882,N_26339);
nor U36424 (N_36424,N_23302,N_26753);
or U36425 (N_36425,N_25275,N_22812);
nand U36426 (N_36426,N_24078,N_25318);
nand U36427 (N_36427,N_20861,N_27642);
or U36428 (N_36428,N_26584,N_29513);
and U36429 (N_36429,N_25614,N_20271);
and U36430 (N_36430,N_28948,N_27108);
nor U36431 (N_36431,N_20659,N_24296);
nand U36432 (N_36432,N_28659,N_26126);
xnor U36433 (N_36433,N_23202,N_24995);
and U36434 (N_36434,N_22287,N_23325);
nor U36435 (N_36435,N_27705,N_23787);
xor U36436 (N_36436,N_20230,N_24775);
nor U36437 (N_36437,N_25005,N_28190);
nand U36438 (N_36438,N_29821,N_22637);
nand U36439 (N_36439,N_22107,N_26160);
nand U36440 (N_36440,N_28264,N_25964);
nor U36441 (N_36441,N_29191,N_26057);
nor U36442 (N_36442,N_24216,N_29248);
and U36443 (N_36443,N_21534,N_23255);
or U36444 (N_36444,N_25493,N_20810);
or U36445 (N_36445,N_21484,N_22497);
and U36446 (N_36446,N_22348,N_28543);
nand U36447 (N_36447,N_21134,N_28192);
and U36448 (N_36448,N_28289,N_20996);
nor U36449 (N_36449,N_20427,N_28880);
and U36450 (N_36450,N_24580,N_22985);
nand U36451 (N_36451,N_21423,N_25981);
or U36452 (N_36452,N_25038,N_24528);
nand U36453 (N_36453,N_28870,N_21744);
xnor U36454 (N_36454,N_26145,N_24503);
and U36455 (N_36455,N_23749,N_24717);
xnor U36456 (N_36456,N_25129,N_20354);
xnor U36457 (N_36457,N_27644,N_23611);
xnor U36458 (N_36458,N_24249,N_26869);
and U36459 (N_36459,N_25512,N_24588);
nor U36460 (N_36460,N_26462,N_26950);
or U36461 (N_36461,N_26623,N_29787);
nor U36462 (N_36462,N_26609,N_25002);
and U36463 (N_36463,N_25165,N_21457);
nor U36464 (N_36464,N_22202,N_28445);
nand U36465 (N_36465,N_22585,N_26434);
xnor U36466 (N_36466,N_24878,N_23038);
or U36467 (N_36467,N_20362,N_27649);
nor U36468 (N_36468,N_20402,N_29089);
and U36469 (N_36469,N_22032,N_24104);
nor U36470 (N_36470,N_25962,N_25335);
xor U36471 (N_36471,N_28196,N_27967);
and U36472 (N_36472,N_25221,N_27388);
nand U36473 (N_36473,N_26132,N_28634);
or U36474 (N_36474,N_28231,N_21459);
xor U36475 (N_36475,N_22902,N_24689);
nand U36476 (N_36476,N_28924,N_24559);
and U36477 (N_36477,N_24015,N_27436);
or U36478 (N_36478,N_24370,N_23156);
nand U36479 (N_36479,N_23785,N_23866);
nor U36480 (N_36480,N_24891,N_22309);
nor U36481 (N_36481,N_25803,N_20645);
and U36482 (N_36482,N_26961,N_27423);
xor U36483 (N_36483,N_28211,N_29373);
nor U36484 (N_36484,N_26932,N_25800);
nor U36485 (N_36485,N_28123,N_25034);
nor U36486 (N_36486,N_20145,N_28649);
and U36487 (N_36487,N_27265,N_27867);
nand U36488 (N_36488,N_22943,N_22474);
and U36489 (N_36489,N_26184,N_24255);
and U36490 (N_36490,N_25816,N_28710);
nor U36491 (N_36491,N_22334,N_28399);
or U36492 (N_36492,N_27919,N_24584);
nand U36493 (N_36493,N_23530,N_22883);
xor U36494 (N_36494,N_29393,N_29319);
nor U36495 (N_36495,N_21106,N_21154);
xor U36496 (N_36496,N_26668,N_21681);
or U36497 (N_36497,N_23980,N_23113);
nand U36498 (N_36498,N_24433,N_26651);
or U36499 (N_36499,N_27803,N_21962);
nor U36500 (N_36500,N_26586,N_28166);
xor U36501 (N_36501,N_22140,N_25390);
or U36502 (N_36502,N_27357,N_25601);
xor U36503 (N_36503,N_25938,N_21677);
or U36504 (N_36504,N_24320,N_22213);
and U36505 (N_36505,N_21789,N_28353);
or U36506 (N_36506,N_28993,N_23576);
or U36507 (N_36507,N_20598,N_20568);
xor U36508 (N_36508,N_29729,N_23172);
nor U36509 (N_36509,N_28889,N_25809);
nor U36510 (N_36510,N_23752,N_22447);
xnor U36511 (N_36511,N_28747,N_22274);
and U36512 (N_36512,N_22682,N_21999);
xor U36513 (N_36513,N_28778,N_21200);
or U36514 (N_36514,N_24283,N_29950);
nor U36515 (N_36515,N_28807,N_29140);
nor U36516 (N_36516,N_21274,N_26664);
nor U36517 (N_36517,N_23268,N_26829);
and U36518 (N_36518,N_23609,N_22798);
and U36519 (N_36519,N_29507,N_20647);
nand U36520 (N_36520,N_25611,N_20234);
or U36521 (N_36521,N_28389,N_23745);
xnor U36522 (N_36522,N_29627,N_24028);
and U36523 (N_36523,N_26316,N_28291);
xnor U36524 (N_36524,N_23629,N_23671);
or U36525 (N_36525,N_21344,N_25377);
nor U36526 (N_36526,N_21102,N_26433);
nand U36527 (N_36527,N_25977,N_22831);
and U36528 (N_36528,N_22204,N_27739);
xnor U36529 (N_36529,N_28203,N_29367);
xnor U36530 (N_36530,N_21200,N_26659);
nand U36531 (N_36531,N_29247,N_21678);
xor U36532 (N_36532,N_26463,N_23142);
nand U36533 (N_36533,N_26148,N_24517);
nor U36534 (N_36534,N_23309,N_20851);
nor U36535 (N_36535,N_24706,N_21513);
and U36536 (N_36536,N_25870,N_22426);
and U36537 (N_36537,N_29283,N_29018);
nand U36538 (N_36538,N_22191,N_25600);
nand U36539 (N_36539,N_21771,N_23480);
and U36540 (N_36540,N_28349,N_27972);
nor U36541 (N_36541,N_20428,N_27698);
and U36542 (N_36542,N_29700,N_29036);
and U36543 (N_36543,N_21375,N_22326);
xnor U36544 (N_36544,N_24789,N_21249);
nand U36545 (N_36545,N_29200,N_26527);
or U36546 (N_36546,N_27484,N_20966);
and U36547 (N_36547,N_24423,N_26341);
nand U36548 (N_36548,N_21780,N_20812);
and U36549 (N_36549,N_23596,N_20141);
nand U36550 (N_36550,N_28857,N_28676);
nor U36551 (N_36551,N_23347,N_25288);
or U36552 (N_36552,N_25940,N_27913);
nand U36553 (N_36553,N_21500,N_28289);
and U36554 (N_36554,N_27035,N_24309);
and U36555 (N_36555,N_27721,N_20396);
nand U36556 (N_36556,N_20044,N_24739);
and U36557 (N_36557,N_23077,N_29022);
nor U36558 (N_36558,N_26121,N_20919);
or U36559 (N_36559,N_28701,N_24950);
or U36560 (N_36560,N_25824,N_21994);
nand U36561 (N_36561,N_20467,N_28508);
nand U36562 (N_36562,N_26386,N_24998);
and U36563 (N_36563,N_29949,N_21742);
xor U36564 (N_36564,N_22486,N_28237);
or U36565 (N_36565,N_21700,N_26488);
nor U36566 (N_36566,N_22121,N_28872);
xnor U36567 (N_36567,N_27680,N_23016);
or U36568 (N_36568,N_24247,N_29132);
nor U36569 (N_36569,N_26087,N_29405);
nor U36570 (N_36570,N_20968,N_21389);
and U36571 (N_36571,N_28003,N_27899);
xnor U36572 (N_36572,N_24384,N_28786);
and U36573 (N_36573,N_29167,N_21910);
or U36574 (N_36574,N_25253,N_21355);
xor U36575 (N_36575,N_20345,N_26095);
xor U36576 (N_36576,N_29379,N_22049);
xnor U36577 (N_36577,N_25301,N_23566);
nor U36578 (N_36578,N_20223,N_26862);
nand U36579 (N_36579,N_25079,N_20732);
or U36580 (N_36580,N_23227,N_24965);
nor U36581 (N_36581,N_24212,N_25757);
xor U36582 (N_36582,N_21238,N_23829);
xor U36583 (N_36583,N_21312,N_25730);
xor U36584 (N_36584,N_25572,N_25068);
nor U36585 (N_36585,N_28055,N_22510);
nand U36586 (N_36586,N_29356,N_25275);
and U36587 (N_36587,N_27608,N_22827);
nand U36588 (N_36588,N_26025,N_20003);
and U36589 (N_36589,N_28805,N_21038);
or U36590 (N_36590,N_21491,N_23836);
nand U36591 (N_36591,N_25101,N_28795);
nand U36592 (N_36592,N_27552,N_21336);
nand U36593 (N_36593,N_29050,N_20347);
or U36594 (N_36594,N_21450,N_23796);
and U36595 (N_36595,N_23935,N_26472);
or U36596 (N_36596,N_26247,N_28309);
nor U36597 (N_36597,N_23035,N_23946);
and U36598 (N_36598,N_23422,N_20845);
nor U36599 (N_36599,N_28472,N_23656);
nand U36600 (N_36600,N_27418,N_29493);
or U36601 (N_36601,N_22923,N_20978);
or U36602 (N_36602,N_21305,N_21248);
xor U36603 (N_36603,N_22523,N_29975);
nor U36604 (N_36604,N_23486,N_24236);
xor U36605 (N_36605,N_21729,N_26945);
xor U36606 (N_36606,N_27091,N_23632);
or U36607 (N_36607,N_25197,N_23726);
nor U36608 (N_36608,N_22488,N_21721);
nand U36609 (N_36609,N_27646,N_23518);
xnor U36610 (N_36610,N_23978,N_22576);
or U36611 (N_36611,N_21385,N_25987);
xor U36612 (N_36612,N_21572,N_22913);
or U36613 (N_36613,N_29828,N_28267);
nand U36614 (N_36614,N_26681,N_26146);
xor U36615 (N_36615,N_21481,N_28643);
xnor U36616 (N_36616,N_20467,N_20327);
xor U36617 (N_36617,N_27266,N_22793);
nor U36618 (N_36618,N_26926,N_28782);
nor U36619 (N_36619,N_26487,N_20774);
xnor U36620 (N_36620,N_28032,N_28948);
and U36621 (N_36621,N_21812,N_23213);
nand U36622 (N_36622,N_25703,N_29242);
xnor U36623 (N_36623,N_26291,N_23368);
or U36624 (N_36624,N_21812,N_20440);
and U36625 (N_36625,N_22292,N_27153);
nand U36626 (N_36626,N_29562,N_28176);
or U36627 (N_36627,N_27187,N_21883);
xnor U36628 (N_36628,N_26038,N_28414);
nand U36629 (N_36629,N_22662,N_23554);
nand U36630 (N_36630,N_25441,N_24866);
and U36631 (N_36631,N_25654,N_26507);
nand U36632 (N_36632,N_24142,N_26642);
or U36633 (N_36633,N_28096,N_29353);
or U36634 (N_36634,N_25680,N_22872);
or U36635 (N_36635,N_25951,N_28789);
xor U36636 (N_36636,N_28042,N_23866);
or U36637 (N_36637,N_28870,N_29848);
nand U36638 (N_36638,N_23920,N_20820);
xnor U36639 (N_36639,N_27840,N_28401);
xor U36640 (N_36640,N_21823,N_23557);
nor U36641 (N_36641,N_25817,N_25055);
xnor U36642 (N_36642,N_21243,N_29595);
and U36643 (N_36643,N_25249,N_21018);
nand U36644 (N_36644,N_26354,N_20691);
and U36645 (N_36645,N_20262,N_23268);
nor U36646 (N_36646,N_22929,N_20459);
and U36647 (N_36647,N_22029,N_28847);
nor U36648 (N_36648,N_25668,N_28630);
xnor U36649 (N_36649,N_20106,N_24100);
xnor U36650 (N_36650,N_23554,N_24288);
nand U36651 (N_36651,N_27031,N_23359);
and U36652 (N_36652,N_22162,N_20662);
or U36653 (N_36653,N_28839,N_20750);
or U36654 (N_36654,N_25471,N_20928);
nor U36655 (N_36655,N_27796,N_28964);
or U36656 (N_36656,N_25893,N_25364);
or U36657 (N_36657,N_20742,N_20208);
nor U36658 (N_36658,N_21855,N_24641);
xor U36659 (N_36659,N_22828,N_27381);
or U36660 (N_36660,N_21289,N_24481);
or U36661 (N_36661,N_22166,N_25077);
and U36662 (N_36662,N_21488,N_21790);
and U36663 (N_36663,N_29073,N_21423);
and U36664 (N_36664,N_27319,N_29500);
nor U36665 (N_36665,N_29619,N_20624);
xor U36666 (N_36666,N_24281,N_28986);
xnor U36667 (N_36667,N_25282,N_20159);
nor U36668 (N_36668,N_27688,N_28044);
xnor U36669 (N_36669,N_21738,N_24186);
or U36670 (N_36670,N_20873,N_27934);
xor U36671 (N_36671,N_22579,N_22414);
nor U36672 (N_36672,N_20442,N_22736);
nand U36673 (N_36673,N_22063,N_23291);
and U36674 (N_36674,N_22525,N_28977);
and U36675 (N_36675,N_22461,N_28457);
and U36676 (N_36676,N_22615,N_29827);
xnor U36677 (N_36677,N_29988,N_24832);
or U36678 (N_36678,N_24376,N_25330);
or U36679 (N_36679,N_25345,N_20267);
xnor U36680 (N_36680,N_28185,N_22808);
or U36681 (N_36681,N_25887,N_20164);
or U36682 (N_36682,N_20210,N_29731);
nor U36683 (N_36683,N_26458,N_26686);
nand U36684 (N_36684,N_21418,N_26184);
and U36685 (N_36685,N_26782,N_29679);
xnor U36686 (N_36686,N_26766,N_29778);
nand U36687 (N_36687,N_26198,N_26387);
xor U36688 (N_36688,N_29741,N_25248);
nor U36689 (N_36689,N_27409,N_26726);
xnor U36690 (N_36690,N_25198,N_20480);
or U36691 (N_36691,N_20391,N_27563);
xor U36692 (N_36692,N_23827,N_28222);
nor U36693 (N_36693,N_24814,N_27108);
or U36694 (N_36694,N_22826,N_21224);
nor U36695 (N_36695,N_27408,N_25641);
nor U36696 (N_36696,N_24014,N_24028);
or U36697 (N_36697,N_20056,N_20398);
nor U36698 (N_36698,N_27040,N_29512);
nor U36699 (N_36699,N_29050,N_25330);
xor U36700 (N_36700,N_29545,N_22625);
nor U36701 (N_36701,N_27068,N_22504);
or U36702 (N_36702,N_27930,N_22175);
nor U36703 (N_36703,N_28395,N_27731);
and U36704 (N_36704,N_23900,N_27343);
or U36705 (N_36705,N_24009,N_24229);
and U36706 (N_36706,N_27157,N_29593);
or U36707 (N_36707,N_26151,N_25292);
nor U36708 (N_36708,N_25051,N_23289);
or U36709 (N_36709,N_24632,N_24586);
xnor U36710 (N_36710,N_25442,N_25137);
nor U36711 (N_36711,N_23903,N_25744);
nand U36712 (N_36712,N_20187,N_20091);
or U36713 (N_36713,N_24721,N_27412);
and U36714 (N_36714,N_25090,N_21903);
xnor U36715 (N_36715,N_25209,N_22860);
xnor U36716 (N_36716,N_27436,N_27291);
and U36717 (N_36717,N_22000,N_29464);
nor U36718 (N_36718,N_22375,N_27458);
and U36719 (N_36719,N_29677,N_21716);
nand U36720 (N_36720,N_29711,N_24938);
xnor U36721 (N_36721,N_23711,N_25582);
nand U36722 (N_36722,N_26357,N_24661);
nand U36723 (N_36723,N_23410,N_22881);
nor U36724 (N_36724,N_25220,N_27617);
xnor U36725 (N_36725,N_21721,N_28600);
nand U36726 (N_36726,N_22125,N_25366);
and U36727 (N_36727,N_20175,N_26079);
or U36728 (N_36728,N_23224,N_26506);
or U36729 (N_36729,N_24866,N_23514);
xnor U36730 (N_36730,N_24766,N_20178);
or U36731 (N_36731,N_21577,N_21208);
nor U36732 (N_36732,N_20876,N_29068);
nand U36733 (N_36733,N_23124,N_20978);
or U36734 (N_36734,N_20293,N_21602);
nand U36735 (N_36735,N_28929,N_23704);
xor U36736 (N_36736,N_28950,N_21981);
nor U36737 (N_36737,N_26297,N_23088);
xnor U36738 (N_36738,N_28987,N_22838);
nor U36739 (N_36739,N_22753,N_22939);
nand U36740 (N_36740,N_24992,N_27940);
xnor U36741 (N_36741,N_29927,N_25028);
nand U36742 (N_36742,N_20517,N_21548);
or U36743 (N_36743,N_22758,N_26965);
and U36744 (N_36744,N_22487,N_29596);
nand U36745 (N_36745,N_20940,N_25664);
nand U36746 (N_36746,N_28510,N_20691);
nand U36747 (N_36747,N_29032,N_27007);
xnor U36748 (N_36748,N_28962,N_26126);
xnor U36749 (N_36749,N_25122,N_28621);
or U36750 (N_36750,N_25478,N_27750);
and U36751 (N_36751,N_29489,N_25725);
nand U36752 (N_36752,N_27210,N_22049);
and U36753 (N_36753,N_28270,N_28686);
nand U36754 (N_36754,N_24775,N_22010);
xnor U36755 (N_36755,N_21058,N_23951);
nand U36756 (N_36756,N_23030,N_22553);
nand U36757 (N_36757,N_27610,N_20087);
xor U36758 (N_36758,N_20503,N_21753);
and U36759 (N_36759,N_26860,N_28509);
nand U36760 (N_36760,N_20658,N_29402);
nand U36761 (N_36761,N_26349,N_29503);
nand U36762 (N_36762,N_23327,N_26058);
xnor U36763 (N_36763,N_25526,N_23319);
nand U36764 (N_36764,N_25320,N_29031);
and U36765 (N_36765,N_29617,N_27402);
and U36766 (N_36766,N_25763,N_29536);
nor U36767 (N_36767,N_27333,N_24110);
and U36768 (N_36768,N_29721,N_26996);
or U36769 (N_36769,N_23071,N_28738);
or U36770 (N_36770,N_24467,N_25143);
nand U36771 (N_36771,N_20614,N_28713);
and U36772 (N_36772,N_24885,N_28714);
nand U36773 (N_36773,N_20794,N_21872);
nor U36774 (N_36774,N_29475,N_27668);
and U36775 (N_36775,N_29192,N_25521);
or U36776 (N_36776,N_22750,N_24575);
or U36777 (N_36777,N_22244,N_21456);
xnor U36778 (N_36778,N_28393,N_20021);
nor U36779 (N_36779,N_25739,N_24828);
nand U36780 (N_36780,N_27534,N_25212);
xnor U36781 (N_36781,N_21723,N_24392);
xor U36782 (N_36782,N_27063,N_20018);
nor U36783 (N_36783,N_21740,N_27107);
xor U36784 (N_36784,N_25727,N_25196);
and U36785 (N_36785,N_23063,N_24572);
nor U36786 (N_36786,N_26872,N_29475);
nand U36787 (N_36787,N_24027,N_20532);
and U36788 (N_36788,N_22270,N_29301);
nor U36789 (N_36789,N_29305,N_24477);
and U36790 (N_36790,N_25350,N_24365);
nand U36791 (N_36791,N_28453,N_27034);
nand U36792 (N_36792,N_28492,N_21513);
and U36793 (N_36793,N_26645,N_25106);
or U36794 (N_36794,N_27448,N_21153);
xor U36795 (N_36795,N_29198,N_25474);
nor U36796 (N_36796,N_22303,N_21950);
or U36797 (N_36797,N_21522,N_23677);
xnor U36798 (N_36798,N_21736,N_20248);
nand U36799 (N_36799,N_21043,N_20015);
xor U36800 (N_36800,N_22121,N_21916);
or U36801 (N_36801,N_28468,N_24106);
nor U36802 (N_36802,N_22108,N_20596);
or U36803 (N_36803,N_21229,N_23289);
xnor U36804 (N_36804,N_25350,N_24209);
nor U36805 (N_36805,N_28505,N_26834);
nor U36806 (N_36806,N_28085,N_25204);
and U36807 (N_36807,N_24766,N_24196);
xor U36808 (N_36808,N_20957,N_22284);
nand U36809 (N_36809,N_23569,N_22673);
and U36810 (N_36810,N_21871,N_20834);
xnor U36811 (N_36811,N_21792,N_27091);
nor U36812 (N_36812,N_22488,N_25964);
nor U36813 (N_36813,N_20822,N_24620);
xnor U36814 (N_36814,N_26482,N_29766);
nor U36815 (N_36815,N_26779,N_27002);
nor U36816 (N_36816,N_23925,N_29589);
or U36817 (N_36817,N_28906,N_24125);
or U36818 (N_36818,N_29822,N_26530);
xnor U36819 (N_36819,N_28596,N_27661);
xor U36820 (N_36820,N_23953,N_26622);
and U36821 (N_36821,N_21477,N_27620);
xor U36822 (N_36822,N_29775,N_27955);
and U36823 (N_36823,N_27741,N_21000);
and U36824 (N_36824,N_25390,N_25518);
and U36825 (N_36825,N_27884,N_22198);
or U36826 (N_36826,N_25468,N_25863);
xnor U36827 (N_36827,N_27866,N_22681);
or U36828 (N_36828,N_20974,N_24460);
and U36829 (N_36829,N_23731,N_29587);
xnor U36830 (N_36830,N_28310,N_27179);
nor U36831 (N_36831,N_25890,N_28953);
nor U36832 (N_36832,N_23575,N_20086);
nand U36833 (N_36833,N_26885,N_29781);
nor U36834 (N_36834,N_29875,N_28156);
or U36835 (N_36835,N_29293,N_24997);
or U36836 (N_36836,N_26661,N_23652);
nor U36837 (N_36837,N_27601,N_26416);
xnor U36838 (N_36838,N_21715,N_24785);
nor U36839 (N_36839,N_28127,N_20842);
nor U36840 (N_36840,N_26332,N_24686);
xor U36841 (N_36841,N_29616,N_26334);
and U36842 (N_36842,N_26100,N_20612);
or U36843 (N_36843,N_20519,N_22942);
nand U36844 (N_36844,N_26587,N_29816);
nor U36845 (N_36845,N_29547,N_20126);
or U36846 (N_36846,N_27301,N_26253);
xor U36847 (N_36847,N_23433,N_27004);
xnor U36848 (N_36848,N_29715,N_23419);
nand U36849 (N_36849,N_29736,N_25583);
or U36850 (N_36850,N_29485,N_28715);
nand U36851 (N_36851,N_25171,N_28649);
nor U36852 (N_36852,N_24670,N_21435);
or U36853 (N_36853,N_21966,N_22063);
or U36854 (N_36854,N_26135,N_24144);
xor U36855 (N_36855,N_20560,N_21775);
or U36856 (N_36856,N_21233,N_24892);
or U36857 (N_36857,N_28810,N_21129);
xor U36858 (N_36858,N_25369,N_24255);
xor U36859 (N_36859,N_26759,N_21471);
nand U36860 (N_36860,N_26496,N_20180);
nor U36861 (N_36861,N_21950,N_23668);
and U36862 (N_36862,N_29108,N_28979);
xnor U36863 (N_36863,N_28703,N_24147);
nand U36864 (N_36864,N_20622,N_29094);
nor U36865 (N_36865,N_25917,N_26613);
or U36866 (N_36866,N_27652,N_20004);
nand U36867 (N_36867,N_26358,N_21506);
nor U36868 (N_36868,N_23316,N_28340);
xor U36869 (N_36869,N_23786,N_26757);
nor U36870 (N_36870,N_20086,N_28600);
xnor U36871 (N_36871,N_25545,N_29986);
and U36872 (N_36872,N_21974,N_28932);
nand U36873 (N_36873,N_20905,N_20500);
nand U36874 (N_36874,N_28103,N_28314);
xnor U36875 (N_36875,N_22509,N_29956);
xor U36876 (N_36876,N_22376,N_25549);
nand U36877 (N_36877,N_21504,N_28458);
and U36878 (N_36878,N_27397,N_20342);
and U36879 (N_36879,N_21056,N_20205);
and U36880 (N_36880,N_20160,N_21838);
nor U36881 (N_36881,N_29211,N_27637);
or U36882 (N_36882,N_29344,N_28187);
or U36883 (N_36883,N_29925,N_21112);
nand U36884 (N_36884,N_26099,N_25241);
nor U36885 (N_36885,N_22417,N_25448);
or U36886 (N_36886,N_28693,N_28139);
and U36887 (N_36887,N_22919,N_22474);
xor U36888 (N_36888,N_20422,N_21829);
or U36889 (N_36889,N_29552,N_20020);
xor U36890 (N_36890,N_21013,N_29033);
nor U36891 (N_36891,N_27849,N_24932);
xnor U36892 (N_36892,N_28654,N_27436);
nor U36893 (N_36893,N_27927,N_29315);
or U36894 (N_36894,N_23357,N_27738);
nor U36895 (N_36895,N_28250,N_24036);
nand U36896 (N_36896,N_24539,N_20576);
nor U36897 (N_36897,N_28457,N_29995);
nor U36898 (N_36898,N_24054,N_23793);
nand U36899 (N_36899,N_23588,N_29196);
xnor U36900 (N_36900,N_21287,N_23931);
nor U36901 (N_36901,N_27556,N_21506);
and U36902 (N_36902,N_25295,N_29201);
nand U36903 (N_36903,N_21017,N_24853);
or U36904 (N_36904,N_24439,N_27563);
nand U36905 (N_36905,N_22203,N_21393);
nor U36906 (N_36906,N_25962,N_22327);
nand U36907 (N_36907,N_28495,N_29825);
nor U36908 (N_36908,N_27036,N_23917);
nor U36909 (N_36909,N_29237,N_27439);
nor U36910 (N_36910,N_20401,N_24190);
nor U36911 (N_36911,N_28448,N_23697);
or U36912 (N_36912,N_23795,N_23965);
or U36913 (N_36913,N_25075,N_24848);
nor U36914 (N_36914,N_26788,N_25898);
nand U36915 (N_36915,N_23461,N_25306);
nand U36916 (N_36916,N_28528,N_29268);
xor U36917 (N_36917,N_29159,N_20818);
and U36918 (N_36918,N_20639,N_23046);
nor U36919 (N_36919,N_24818,N_28459);
or U36920 (N_36920,N_24100,N_27876);
or U36921 (N_36921,N_23393,N_24453);
nand U36922 (N_36922,N_26052,N_21410);
nor U36923 (N_36923,N_24313,N_23656);
nor U36924 (N_36924,N_24347,N_20112);
or U36925 (N_36925,N_20290,N_25617);
or U36926 (N_36926,N_28801,N_26355);
nor U36927 (N_36927,N_29649,N_22752);
nor U36928 (N_36928,N_23192,N_29063);
nor U36929 (N_36929,N_25413,N_20657);
nor U36930 (N_36930,N_21677,N_28735);
xnor U36931 (N_36931,N_23698,N_27841);
nand U36932 (N_36932,N_23222,N_21963);
nand U36933 (N_36933,N_24774,N_28773);
xor U36934 (N_36934,N_27086,N_22618);
nor U36935 (N_36935,N_21977,N_29874);
and U36936 (N_36936,N_23402,N_21486);
nor U36937 (N_36937,N_24990,N_22593);
nor U36938 (N_36938,N_20888,N_26017);
nand U36939 (N_36939,N_25122,N_28830);
nand U36940 (N_36940,N_25576,N_29422);
and U36941 (N_36941,N_23654,N_29644);
or U36942 (N_36942,N_27637,N_29347);
and U36943 (N_36943,N_26283,N_26939);
xnor U36944 (N_36944,N_26070,N_24532);
nor U36945 (N_36945,N_28805,N_23962);
nand U36946 (N_36946,N_20023,N_26130);
and U36947 (N_36947,N_29778,N_26610);
nand U36948 (N_36948,N_25887,N_25767);
xnor U36949 (N_36949,N_22652,N_24493);
xnor U36950 (N_36950,N_27257,N_29422);
or U36951 (N_36951,N_25448,N_26214);
and U36952 (N_36952,N_26707,N_23015);
nor U36953 (N_36953,N_29583,N_23112);
nor U36954 (N_36954,N_23691,N_21697);
xnor U36955 (N_36955,N_27405,N_27909);
or U36956 (N_36956,N_22664,N_21685);
nor U36957 (N_36957,N_22236,N_24786);
or U36958 (N_36958,N_26709,N_26714);
and U36959 (N_36959,N_25551,N_26287);
or U36960 (N_36960,N_26826,N_23956);
xor U36961 (N_36961,N_28552,N_26615);
and U36962 (N_36962,N_24393,N_23418);
and U36963 (N_36963,N_20578,N_22938);
and U36964 (N_36964,N_25122,N_28948);
or U36965 (N_36965,N_26473,N_28600);
xnor U36966 (N_36966,N_27078,N_24243);
or U36967 (N_36967,N_21914,N_22145);
and U36968 (N_36968,N_29377,N_28611);
and U36969 (N_36969,N_29576,N_25605);
xnor U36970 (N_36970,N_22575,N_24236);
xnor U36971 (N_36971,N_20791,N_25706);
nand U36972 (N_36972,N_21659,N_22793);
xor U36973 (N_36973,N_29838,N_29328);
xnor U36974 (N_36974,N_28534,N_29528);
nand U36975 (N_36975,N_22348,N_27360);
xnor U36976 (N_36976,N_21321,N_20967);
and U36977 (N_36977,N_28983,N_23283);
and U36978 (N_36978,N_27721,N_21670);
nor U36979 (N_36979,N_22611,N_29231);
and U36980 (N_36980,N_21686,N_21394);
xor U36981 (N_36981,N_27007,N_25954);
or U36982 (N_36982,N_20908,N_21822);
nor U36983 (N_36983,N_27834,N_22102);
xnor U36984 (N_36984,N_21017,N_23653);
nand U36985 (N_36985,N_25799,N_24945);
xor U36986 (N_36986,N_24603,N_27212);
xor U36987 (N_36987,N_23829,N_20330);
and U36988 (N_36988,N_25288,N_21549);
nand U36989 (N_36989,N_24803,N_28996);
nand U36990 (N_36990,N_24428,N_25870);
or U36991 (N_36991,N_29855,N_24399);
or U36992 (N_36992,N_21676,N_24204);
and U36993 (N_36993,N_26259,N_24868);
xnor U36994 (N_36994,N_28206,N_29994);
xnor U36995 (N_36995,N_24485,N_20745);
and U36996 (N_36996,N_26706,N_26778);
xor U36997 (N_36997,N_21531,N_24111);
or U36998 (N_36998,N_24129,N_20155);
or U36999 (N_36999,N_24265,N_29066);
and U37000 (N_37000,N_25267,N_20125);
or U37001 (N_37001,N_29667,N_21873);
nand U37002 (N_37002,N_20865,N_28519);
or U37003 (N_37003,N_26540,N_28102);
nor U37004 (N_37004,N_26989,N_29770);
xnor U37005 (N_37005,N_21939,N_20058);
or U37006 (N_37006,N_21221,N_23033);
xor U37007 (N_37007,N_27284,N_22808);
xnor U37008 (N_37008,N_21447,N_27472);
or U37009 (N_37009,N_26778,N_23632);
nand U37010 (N_37010,N_27656,N_25630);
nand U37011 (N_37011,N_26057,N_25818);
or U37012 (N_37012,N_24346,N_22423);
and U37013 (N_37013,N_26848,N_29012);
or U37014 (N_37014,N_25439,N_26546);
or U37015 (N_37015,N_22123,N_21600);
nor U37016 (N_37016,N_23226,N_29414);
and U37017 (N_37017,N_25111,N_28653);
or U37018 (N_37018,N_20790,N_28536);
nor U37019 (N_37019,N_26610,N_23732);
or U37020 (N_37020,N_26198,N_23090);
nor U37021 (N_37021,N_20461,N_28047);
or U37022 (N_37022,N_25361,N_25572);
and U37023 (N_37023,N_20955,N_21002);
or U37024 (N_37024,N_28210,N_28007);
xnor U37025 (N_37025,N_27944,N_29896);
nor U37026 (N_37026,N_23720,N_28494);
xor U37027 (N_37027,N_28384,N_29168);
or U37028 (N_37028,N_29157,N_21051);
nor U37029 (N_37029,N_20559,N_28313);
or U37030 (N_37030,N_23725,N_28864);
nand U37031 (N_37031,N_25961,N_20501);
xor U37032 (N_37032,N_20381,N_20172);
nand U37033 (N_37033,N_29893,N_26225);
or U37034 (N_37034,N_20148,N_21263);
nor U37035 (N_37035,N_22446,N_25195);
nand U37036 (N_37036,N_27034,N_21673);
xnor U37037 (N_37037,N_29597,N_27505);
xnor U37038 (N_37038,N_21984,N_24740);
or U37039 (N_37039,N_20988,N_21727);
and U37040 (N_37040,N_27140,N_20717);
or U37041 (N_37041,N_25552,N_25816);
or U37042 (N_37042,N_26322,N_23231);
and U37043 (N_37043,N_26556,N_21248);
nand U37044 (N_37044,N_28341,N_27830);
nand U37045 (N_37045,N_29964,N_24465);
nor U37046 (N_37046,N_23332,N_27138);
nand U37047 (N_37047,N_22217,N_23142);
nand U37048 (N_37048,N_27546,N_20516);
nor U37049 (N_37049,N_29442,N_27790);
nand U37050 (N_37050,N_23045,N_26278);
nand U37051 (N_37051,N_25871,N_29721);
and U37052 (N_37052,N_28329,N_25219);
or U37053 (N_37053,N_23125,N_27471);
or U37054 (N_37054,N_26353,N_24039);
xor U37055 (N_37055,N_28579,N_25047);
xnor U37056 (N_37056,N_29469,N_25296);
nand U37057 (N_37057,N_28810,N_26366);
xor U37058 (N_37058,N_29323,N_26007);
or U37059 (N_37059,N_22860,N_21508);
or U37060 (N_37060,N_29695,N_27831);
xor U37061 (N_37061,N_23819,N_26182);
and U37062 (N_37062,N_24914,N_22607);
xor U37063 (N_37063,N_28819,N_21486);
xnor U37064 (N_37064,N_25649,N_26300);
nand U37065 (N_37065,N_21964,N_23773);
and U37066 (N_37066,N_23475,N_23068);
or U37067 (N_37067,N_20890,N_29531);
nand U37068 (N_37068,N_21828,N_23204);
nand U37069 (N_37069,N_28581,N_29470);
nor U37070 (N_37070,N_26833,N_23659);
and U37071 (N_37071,N_29519,N_26020);
and U37072 (N_37072,N_23080,N_28492);
nor U37073 (N_37073,N_20220,N_23352);
or U37074 (N_37074,N_29999,N_26181);
xnor U37075 (N_37075,N_21550,N_27717);
nand U37076 (N_37076,N_20547,N_29776);
and U37077 (N_37077,N_26546,N_27725);
and U37078 (N_37078,N_25472,N_28543);
nand U37079 (N_37079,N_23573,N_20603);
nand U37080 (N_37080,N_29709,N_20289);
nand U37081 (N_37081,N_24764,N_29919);
nand U37082 (N_37082,N_20099,N_27706);
xnor U37083 (N_37083,N_22998,N_23305);
nor U37084 (N_37084,N_23460,N_26136);
nor U37085 (N_37085,N_27934,N_23401);
or U37086 (N_37086,N_20443,N_23526);
nand U37087 (N_37087,N_26945,N_21535);
xor U37088 (N_37088,N_20098,N_23890);
and U37089 (N_37089,N_22254,N_23168);
nand U37090 (N_37090,N_20857,N_27611);
nor U37091 (N_37091,N_22864,N_29701);
nand U37092 (N_37092,N_25981,N_21924);
nor U37093 (N_37093,N_29411,N_29348);
nor U37094 (N_37094,N_23457,N_23698);
nor U37095 (N_37095,N_22708,N_26630);
or U37096 (N_37096,N_23343,N_23491);
xor U37097 (N_37097,N_26930,N_24897);
xnor U37098 (N_37098,N_20336,N_21939);
xor U37099 (N_37099,N_25330,N_27090);
or U37100 (N_37100,N_20471,N_21836);
nor U37101 (N_37101,N_25887,N_27332);
nor U37102 (N_37102,N_29127,N_20152);
or U37103 (N_37103,N_28867,N_28762);
and U37104 (N_37104,N_20402,N_29778);
or U37105 (N_37105,N_28404,N_23548);
and U37106 (N_37106,N_28905,N_29010);
nor U37107 (N_37107,N_20242,N_21348);
xnor U37108 (N_37108,N_25760,N_24522);
and U37109 (N_37109,N_26739,N_29876);
nand U37110 (N_37110,N_22364,N_20306);
nor U37111 (N_37111,N_22795,N_29756);
xnor U37112 (N_37112,N_21630,N_25790);
or U37113 (N_37113,N_27252,N_25516);
nand U37114 (N_37114,N_21847,N_29475);
nand U37115 (N_37115,N_27459,N_29664);
or U37116 (N_37116,N_27412,N_26471);
nor U37117 (N_37117,N_27755,N_21349);
nor U37118 (N_37118,N_29588,N_29937);
or U37119 (N_37119,N_29212,N_23467);
or U37120 (N_37120,N_26372,N_28113);
or U37121 (N_37121,N_20458,N_27262);
and U37122 (N_37122,N_22513,N_26157);
xor U37123 (N_37123,N_21312,N_20617);
and U37124 (N_37124,N_22096,N_23207);
nor U37125 (N_37125,N_21088,N_26465);
xnor U37126 (N_37126,N_27343,N_22410);
xnor U37127 (N_37127,N_22637,N_27554);
and U37128 (N_37128,N_22578,N_22884);
nand U37129 (N_37129,N_20372,N_20964);
nand U37130 (N_37130,N_23323,N_25352);
nor U37131 (N_37131,N_25925,N_27924);
nand U37132 (N_37132,N_24880,N_28556);
nand U37133 (N_37133,N_29027,N_23201);
xnor U37134 (N_37134,N_28493,N_24592);
xnor U37135 (N_37135,N_20092,N_22809);
or U37136 (N_37136,N_25657,N_27981);
nand U37137 (N_37137,N_23940,N_28703);
or U37138 (N_37138,N_22594,N_29399);
nor U37139 (N_37139,N_28730,N_25425);
xor U37140 (N_37140,N_21070,N_21505);
and U37141 (N_37141,N_23047,N_21062);
xor U37142 (N_37142,N_21208,N_20482);
and U37143 (N_37143,N_27736,N_26621);
nor U37144 (N_37144,N_22345,N_25848);
or U37145 (N_37145,N_26268,N_29134);
nand U37146 (N_37146,N_27765,N_26210);
nor U37147 (N_37147,N_29606,N_23362);
or U37148 (N_37148,N_20571,N_27720);
and U37149 (N_37149,N_24927,N_20245);
nor U37150 (N_37150,N_23979,N_22768);
or U37151 (N_37151,N_21935,N_29199);
and U37152 (N_37152,N_21396,N_22125);
and U37153 (N_37153,N_21404,N_27588);
or U37154 (N_37154,N_26706,N_29098);
or U37155 (N_37155,N_24095,N_27336);
nor U37156 (N_37156,N_27459,N_26894);
xnor U37157 (N_37157,N_24410,N_24574);
nand U37158 (N_37158,N_21259,N_21998);
xnor U37159 (N_37159,N_21776,N_23660);
nor U37160 (N_37160,N_24351,N_22783);
nand U37161 (N_37161,N_20642,N_22067);
nor U37162 (N_37162,N_20527,N_26690);
or U37163 (N_37163,N_25965,N_29698);
or U37164 (N_37164,N_21858,N_21670);
nand U37165 (N_37165,N_22639,N_29263);
nand U37166 (N_37166,N_28587,N_29360);
nor U37167 (N_37167,N_29886,N_25104);
or U37168 (N_37168,N_21110,N_28942);
xor U37169 (N_37169,N_22858,N_29059);
xnor U37170 (N_37170,N_29773,N_24627);
nor U37171 (N_37171,N_29764,N_25692);
nand U37172 (N_37172,N_27213,N_29548);
xnor U37173 (N_37173,N_28622,N_23968);
and U37174 (N_37174,N_29402,N_25231);
nand U37175 (N_37175,N_21091,N_29895);
or U37176 (N_37176,N_28228,N_25822);
xor U37177 (N_37177,N_22895,N_22163);
nor U37178 (N_37178,N_29333,N_25100);
and U37179 (N_37179,N_28480,N_26584);
nor U37180 (N_37180,N_23727,N_27198);
nor U37181 (N_37181,N_20902,N_29837);
or U37182 (N_37182,N_21520,N_21072);
nand U37183 (N_37183,N_28760,N_22495);
and U37184 (N_37184,N_22041,N_24260);
and U37185 (N_37185,N_21918,N_21530);
and U37186 (N_37186,N_23076,N_29739);
and U37187 (N_37187,N_28150,N_26798);
nand U37188 (N_37188,N_24155,N_21870);
nand U37189 (N_37189,N_27580,N_24369);
xnor U37190 (N_37190,N_25236,N_29332);
xor U37191 (N_37191,N_27134,N_26106);
or U37192 (N_37192,N_24416,N_24829);
or U37193 (N_37193,N_21706,N_26347);
nand U37194 (N_37194,N_25299,N_24283);
and U37195 (N_37195,N_29942,N_23346);
xor U37196 (N_37196,N_29134,N_20108);
or U37197 (N_37197,N_26089,N_28222);
and U37198 (N_37198,N_27953,N_28887);
xor U37199 (N_37199,N_22511,N_29689);
xnor U37200 (N_37200,N_28394,N_25910);
nand U37201 (N_37201,N_24011,N_20626);
or U37202 (N_37202,N_20845,N_29886);
or U37203 (N_37203,N_29847,N_28473);
xor U37204 (N_37204,N_25331,N_28064);
xor U37205 (N_37205,N_20195,N_25983);
and U37206 (N_37206,N_23085,N_26317);
xnor U37207 (N_37207,N_26374,N_21935);
or U37208 (N_37208,N_22800,N_22151);
xor U37209 (N_37209,N_28367,N_22583);
and U37210 (N_37210,N_23686,N_27623);
and U37211 (N_37211,N_24475,N_27188);
and U37212 (N_37212,N_22137,N_23724);
or U37213 (N_37213,N_21636,N_28403);
nand U37214 (N_37214,N_28005,N_20971);
and U37215 (N_37215,N_21743,N_29523);
or U37216 (N_37216,N_27544,N_23546);
nor U37217 (N_37217,N_28455,N_27654);
xor U37218 (N_37218,N_25352,N_28893);
or U37219 (N_37219,N_26531,N_21839);
xnor U37220 (N_37220,N_27438,N_22214);
or U37221 (N_37221,N_21806,N_26178);
nor U37222 (N_37222,N_25319,N_29442);
nor U37223 (N_37223,N_25685,N_27820);
or U37224 (N_37224,N_27579,N_24507);
and U37225 (N_37225,N_29596,N_22320);
nand U37226 (N_37226,N_26603,N_29652);
nor U37227 (N_37227,N_24232,N_21569);
and U37228 (N_37228,N_25623,N_29761);
nor U37229 (N_37229,N_22924,N_20145);
xor U37230 (N_37230,N_20632,N_22862);
nand U37231 (N_37231,N_28016,N_27070);
or U37232 (N_37232,N_29092,N_27201);
nand U37233 (N_37233,N_23898,N_23494);
or U37234 (N_37234,N_24283,N_21036);
xnor U37235 (N_37235,N_24200,N_25569);
nand U37236 (N_37236,N_22264,N_28919);
and U37237 (N_37237,N_20558,N_21532);
xnor U37238 (N_37238,N_25651,N_29127);
and U37239 (N_37239,N_29968,N_23006);
nor U37240 (N_37240,N_23435,N_22584);
and U37241 (N_37241,N_21905,N_26167);
and U37242 (N_37242,N_25675,N_23904);
nand U37243 (N_37243,N_28583,N_22209);
or U37244 (N_37244,N_23932,N_26979);
nand U37245 (N_37245,N_28964,N_29116);
or U37246 (N_37246,N_29403,N_27270);
nand U37247 (N_37247,N_29450,N_27107);
and U37248 (N_37248,N_24480,N_23118);
nor U37249 (N_37249,N_28666,N_26696);
and U37250 (N_37250,N_21838,N_27986);
nand U37251 (N_37251,N_23549,N_28252);
xnor U37252 (N_37252,N_26982,N_24444);
and U37253 (N_37253,N_25550,N_27345);
xor U37254 (N_37254,N_26826,N_23681);
or U37255 (N_37255,N_29382,N_22687);
nand U37256 (N_37256,N_24451,N_22752);
xnor U37257 (N_37257,N_27143,N_25198);
nor U37258 (N_37258,N_22418,N_28054);
nand U37259 (N_37259,N_27767,N_25575);
nand U37260 (N_37260,N_21318,N_21333);
nand U37261 (N_37261,N_22593,N_20685);
or U37262 (N_37262,N_27910,N_24347);
nand U37263 (N_37263,N_20495,N_28110);
and U37264 (N_37264,N_27278,N_20862);
or U37265 (N_37265,N_20668,N_20887);
nand U37266 (N_37266,N_29976,N_28175);
nor U37267 (N_37267,N_27740,N_24884);
xor U37268 (N_37268,N_24119,N_27359);
xnor U37269 (N_37269,N_25391,N_27989);
nor U37270 (N_37270,N_29868,N_29149);
or U37271 (N_37271,N_28494,N_21397);
nand U37272 (N_37272,N_29470,N_29678);
nor U37273 (N_37273,N_29560,N_21504);
or U37274 (N_37274,N_20832,N_26526);
nor U37275 (N_37275,N_21096,N_24736);
or U37276 (N_37276,N_22367,N_26237);
xor U37277 (N_37277,N_23604,N_25267);
nor U37278 (N_37278,N_27439,N_28869);
or U37279 (N_37279,N_23798,N_29055);
xnor U37280 (N_37280,N_27729,N_26459);
nand U37281 (N_37281,N_29843,N_27104);
xor U37282 (N_37282,N_21307,N_25271);
or U37283 (N_37283,N_21638,N_26918);
xnor U37284 (N_37284,N_29055,N_28432);
nor U37285 (N_37285,N_22012,N_22034);
xnor U37286 (N_37286,N_27789,N_25484);
nand U37287 (N_37287,N_28015,N_25443);
and U37288 (N_37288,N_21909,N_23437);
and U37289 (N_37289,N_29965,N_26305);
nor U37290 (N_37290,N_27585,N_24971);
nor U37291 (N_37291,N_25647,N_26970);
nor U37292 (N_37292,N_26009,N_24166);
nand U37293 (N_37293,N_24364,N_23391);
xnor U37294 (N_37294,N_23728,N_29175);
or U37295 (N_37295,N_23969,N_26044);
and U37296 (N_37296,N_23530,N_27641);
nand U37297 (N_37297,N_29023,N_29171);
nor U37298 (N_37298,N_29125,N_22908);
and U37299 (N_37299,N_22292,N_20563);
and U37300 (N_37300,N_26181,N_27791);
or U37301 (N_37301,N_23046,N_21102);
and U37302 (N_37302,N_24002,N_23460);
xnor U37303 (N_37303,N_25637,N_28794);
nand U37304 (N_37304,N_29750,N_23403);
and U37305 (N_37305,N_29799,N_29481);
or U37306 (N_37306,N_28175,N_28943);
and U37307 (N_37307,N_26980,N_20621);
nor U37308 (N_37308,N_25835,N_29045);
xor U37309 (N_37309,N_27571,N_29500);
or U37310 (N_37310,N_22308,N_26471);
or U37311 (N_37311,N_23022,N_28622);
xor U37312 (N_37312,N_22764,N_21579);
nand U37313 (N_37313,N_21911,N_26285);
or U37314 (N_37314,N_28642,N_20745);
nand U37315 (N_37315,N_21247,N_23347);
or U37316 (N_37316,N_28205,N_27182);
or U37317 (N_37317,N_26149,N_23045);
xnor U37318 (N_37318,N_23975,N_25356);
nand U37319 (N_37319,N_24880,N_21047);
or U37320 (N_37320,N_21029,N_27254);
xor U37321 (N_37321,N_20025,N_20367);
xor U37322 (N_37322,N_24548,N_24534);
and U37323 (N_37323,N_29546,N_24278);
or U37324 (N_37324,N_26778,N_23135);
or U37325 (N_37325,N_21713,N_25936);
xnor U37326 (N_37326,N_29388,N_22804);
nand U37327 (N_37327,N_23531,N_25574);
and U37328 (N_37328,N_25483,N_24781);
or U37329 (N_37329,N_27478,N_23404);
xnor U37330 (N_37330,N_26361,N_21395);
nand U37331 (N_37331,N_23457,N_23056);
nor U37332 (N_37332,N_20408,N_20784);
xor U37333 (N_37333,N_24294,N_27198);
nor U37334 (N_37334,N_22932,N_23649);
or U37335 (N_37335,N_24417,N_23132);
xor U37336 (N_37336,N_24888,N_27234);
nand U37337 (N_37337,N_25652,N_27184);
nor U37338 (N_37338,N_24410,N_24658);
xnor U37339 (N_37339,N_21481,N_28791);
or U37340 (N_37340,N_21860,N_24576);
nand U37341 (N_37341,N_20140,N_27149);
nand U37342 (N_37342,N_23298,N_21530);
nor U37343 (N_37343,N_29933,N_25413);
nor U37344 (N_37344,N_25276,N_29118);
nor U37345 (N_37345,N_29096,N_29839);
xnor U37346 (N_37346,N_23422,N_21483);
nand U37347 (N_37347,N_24479,N_28810);
and U37348 (N_37348,N_22396,N_22499);
nor U37349 (N_37349,N_20384,N_26001);
nand U37350 (N_37350,N_27736,N_25120);
xor U37351 (N_37351,N_25778,N_21832);
and U37352 (N_37352,N_22980,N_21028);
xor U37353 (N_37353,N_23046,N_21736);
nand U37354 (N_37354,N_22963,N_24913);
nand U37355 (N_37355,N_25475,N_26435);
xnor U37356 (N_37356,N_21789,N_27576);
nand U37357 (N_37357,N_23159,N_28967);
xor U37358 (N_37358,N_26356,N_28922);
and U37359 (N_37359,N_22349,N_25116);
xor U37360 (N_37360,N_26664,N_23241);
xnor U37361 (N_37361,N_23197,N_24702);
and U37362 (N_37362,N_25711,N_26934);
nand U37363 (N_37363,N_23980,N_28625);
or U37364 (N_37364,N_22510,N_29697);
or U37365 (N_37365,N_21120,N_24624);
nand U37366 (N_37366,N_26603,N_21809);
xor U37367 (N_37367,N_28683,N_20054);
or U37368 (N_37368,N_28370,N_27022);
or U37369 (N_37369,N_27316,N_26500);
and U37370 (N_37370,N_27079,N_22481);
xnor U37371 (N_37371,N_23479,N_29582);
nor U37372 (N_37372,N_29116,N_24735);
nor U37373 (N_37373,N_22197,N_26240);
xnor U37374 (N_37374,N_27288,N_27016);
xor U37375 (N_37375,N_23717,N_28803);
or U37376 (N_37376,N_24765,N_22419);
or U37377 (N_37377,N_20549,N_25285);
and U37378 (N_37378,N_25576,N_22595);
or U37379 (N_37379,N_20549,N_22774);
xnor U37380 (N_37380,N_29567,N_27829);
xor U37381 (N_37381,N_20705,N_22758);
or U37382 (N_37382,N_26892,N_22293);
or U37383 (N_37383,N_29956,N_28630);
or U37384 (N_37384,N_25695,N_22430);
nand U37385 (N_37385,N_20511,N_25197);
and U37386 (N_37386,N_21460,N_24133);
xnor U37387 (N_37387,N_22624,N_29129);
xnor U37388 (N_37388,N_27968,N_28077);
or U37389 (N_37389,N_25437,N_28253);
nor U37390 (N_37390,N_25794,N_23532);
xor U37391 (N_37391,N_27801,N_22349);
xor U37392 (N_37392,N_22332,N_26831);
or U37393 (N_37393,N_28878,N_28810);
nand U37394 (N_37394,N_28673,N_26024);
nor U37395 (N_37395,N_24060,N_20494);
xor U37396 (N_37396,N_21836,N_22214);
and U37397 (N_37397,N_24898,N_26114);
xnor U37398 (N_37398,N_22557,N_22861);
nand U37399 (N_37399,N_26230,N_23428);
or U37400 (N_37400,N_27278,N_20048);
or U37401 (N_37401,N_27197,N_29261);
and U37402 (N_37402,N_27660,N_20374);
xor U37403 (N_37403,N_20072,N_27397);
xnor U37404 (N_37404,N_23611,N_22598);
nor U37405 (N_37405,N_24616,N_24890);
and U37406 (N_37406,N_24704,N_24532);
or U37407 (N_37407,N_25035,N_22506);
xor U37408 (N_37408,N_29703,N_22036);
and U37409 (N_37409,N_22236,N_21664);
and U37410 (N_37410,N_25233,N_20947);
and U37411 (N_37411,N_21677,N_26368);
xor U37412 (N_37412,N_26080,N_20183);
and U37413 (N_37413,N_29005,N_28750);
or U37414 (N_37414,N_29524,N_25819);
and U37415 (N_37415,N_29926,N_23967);
nor U37416 (N_37416,N_23251,N_23556);
or U37417 (N_37417,N_25497,N_26278);
or U37418 (N_37418,N_21171,N_25542);
nand U37419 (N_37419,N_23208,N_29679);
nand U37420 (N_37420,N_26137,N_28331);
nor U37421 (N_37421,N_20404,N_20488);
or U37422 (N_37422,N_25245,N_25998);
nor U37423 (N_37423,N_29368,N_20145);
nor U37424 (N_37424,N_21920,N_20253);
nor U37425 (N_37425,N_29091,N_28107);
or U37426 (N_37426,N_24862,N_22434);
and U37427 (N_37427,N_28861,N_25157);
and U37428 (N_37428,N_27273,N_29281);
nand U37429 (N_37429,N_26638,N_22392);
or U37430 (N_37430,N_21117,N_21566);
or U37431 (N_37431,N_29410,N_20087);
xnor U37432 (N_37432,N_21619,N_27350);
nor U37433 (N_37433,N_29792,N_27081);
nand U37434 (N_37434,N_21746,N_23270);
nand U37435 (N_37435,N_22979,N_25752);
nor U37436 (N_37436,N_23856,N_29345);
xnor U37437 (N_37437,N_24542,N_28198);
nand U37438 (N_37438,N_23421,N_22686);
xnor U37439 (N_37439,N_23692,N_27151);
and U37440 (N_37440,N_29419,N_26242);
or U37441 (N_37441,N_22337,N_25467);
or U37442 (N_37442,N_22964,N_29066);
and U37443 (N_37443,N_24710,N_29754);
or U37444 (N_37444,N_25420,N_22627);
or U37445 (N_37445,N_25754,N_25270);
nor U37446 (N_37446,N_25270,N_27057);
and U37447 (N_37447,N_29622,N_21265);
or U37448 (N_37448,N_26079,N_20971);
nor U37449 (N_37449,N_26719,N_27467);
xnor U37450 (N_37450,N_23226,N_22398);
nand U37451 (N_37451,N_28981,N_25792);
xnor U37452 (N_37452,N_23501,N_28213);
or U37453 (N_37453,N_24059,N_22132);
nor U37454 (N_37454,N_29364,N_20834);
and U37455 (N_37455,N_27857,N_23072);
xnor U37456 (N_37456,N_22592,N_25390);
nor U37457 (N_37457,N_21089,N_28458);
xnor U37458 (N_37458,N_26989,N_26622);
or U37459 (N_37459,N_20774,N_25416);
xor U37460 (N_37460,N_23047,N_27577);
nand U37461 (N_37461,N_23278,N_25823);
xor U37462 (N_37462,N_20434,N_25551);
nand U37463 (N_37463,N_28296,N_22291);
nor U37464 (N_37464,N_25817,N_22133);
and U37465 (N_37465,N_23953,N_24900);
nor U37466 (N_37466,N_27723,N_27758);
nand U37467 (N_37467,N_28817,N_28260);
nand U37468 (N_37468,N_25501,N_26576);
or U37469 (N_37469,N_20878,N_28165);
or U37470 (N_37470,N_25320,N_26723);
nor U37471 (N_37471,N_21285,N_26921);
nor U37472 (N_37472,N_24197,N_28264);
xor U37473 (N_37473,N_29832,N_29553);
xnor U37474 (N_37474,N_21864,N_25773);
and U37475 (N_37475,N_28370,N_22007);
xor U37476 (N_37476,N_22556,N_29025);
or U37477 (N_37477,N_21779,N_29774);
or U37478 (N_37478,N_21347,N_22206);
nand U37479 (N_37479,N_24915,N_24051);
nor U37480 (N_37480,N_27320,N_27595);
or U37481 (N_37481,N_23438,N_26913);
xor U37482 (N_37482,N_22251,N_23233);
or U37483 (N_37483,N_23790,N_20904);
nor U37484 (N_37484,N_28888,N_24304);
xnor U37485 (N_37485,N_26603,N_21071);
nor U37486 (N_37486,N_27426,N_28389);
nor U37487 (N_37487,N_25345,N_24267);
xnor U37488 (N_37488,N_24112,N_27601);
nand U37489 (N_37489,N_25928,N_29151);
and U37490 (N_37490,N_25578,N_20761);
and U37491 (N_37491,N_28663,N_29060);
xnor U37492 (N_37492,N_20255,N_24325);
or U37493 (N_37493,N_21012,N_26547);
nor U37494 (N_37494,N_26461,N_25911);
nand U37495 (N_37495,N_21796,N_29522);
nand U37496 (N_37496,N_20922,N_21117);
xor U37497 (N_37497,N_22613,N_24226);
nand U37498 (N_37498,N_26011,N_28775);
xnor U37499 (N_37499,N_28357,N_21748);
nor U37500 (N_37500,N_24622,N_28984);
and U37501 (N_37501,N_21647,N_22065);
nand U37502 (N_37502,N_21634,N_29278);
and U37503 (N_37503,N_22908,N_24493);
and U37504 (N_37504,N_28735,N_27245);
nor U37505 (N_37505,N_22774,N_21141);
and U37506 (N_37506,N_21256,N_22916);
xor U37507 (N_37507,N_22090,N_26844);
xnor U37508 (N_37508,N_25772,N_25058);
or U37509 (N_37509,N_21030,N_28161);
and U37510 (N_37510,N_25563,N_24213);
nand U37511 (N_37511,N_21530,N_29030);
or U37512 (N_37512,N_24790,N_22902);
or U37513 (N_37513,N_20778,N_21116);
and U37514 (N_37514,N_25661,N_27466);
nand U37515 (N_37515,N_25496,N_29214);
and U37516 (N_37516,N_21816,N_22212);
nor U37517 (N_37517,N_21496,N_20631);
and U37518 (N_37518,N_21721,N_23142);
and U37519 (N_37519,N_25159,N_24933);
nor U37520 (N_37520,N_26202,N_25802);
nand U37521 (N_37521,N_25763,N_28551);
and U37522 (N_37522,N_21092,N_21746);
xnor U37523 (N_37523,N_29186,N_24202);
and U37524 (N_37524,N_29100,N_23658);
nand U37525 (N_37525,N_27464,N_21236);
nor U37526 (N_37526,N_27376,N_24751);
nand U37527 (N_37527,N_26137,N_26172);
or U37528 (N_37528,N_22897,N_21892);
nor U37529 (N_37529,N_27975,N_23717);
nand U37530 (N_37530,N_25109,N_27688);
nor U37531 (N_37531,N_28791,N_21845);
nor U37532 (N_37532,N_25622,N_25291);
or U37533 (N_37533,N_25951,N_29139);
or U37534 (N_37534,N_28629,N_25556);
nand U37535 (N_37535,N_20829,N_26940);
nor U37536 (N_37536,N_21910,N_23860);
or U37537 (N_37537,N_23533,N_21680);
or U37538 (N_37538,N_25358,N_26031);
nand U37539 (N_37539,N_27205,N_24586);
and U37540 (N_37540,N_25268,N_25726);
or U37541 (N_37541,N_26451,N_21313);
xnor U37542 (N_37542,N_22554,N_28813);
or U37543 (N_37543,N_21269,N_25567);
or U37544 (N_37544,N_26259,N_24889);
and U37545 (N_37545,N_21453,N_25949);
or U37546 (N_37546,N_21118,N_28237);
nor U37547 (N_37547,N_28947,N_29540);
nand U37548 (N_37548,N_25822,N_26231);
and U37549 (N_37549,N_23958,N_27292);
or U37550 (N_37550,N_23643,N_24772);
or U37551 (N_37551,N_20665,N_20790);
nor U37552 (N_37552,N_25910,N_20928);
or U37553 (N_37553,N_25513,N_27868);
xnor U37554 (N_37554,N_28694,N_20630);
or U37555 (N_37555,N_28929,N_27574);
xor U37556 (N_37556,N_26384,N_28071);
nand U37557 (N_37557,N_24041,N_27637);
xnor U37558 (N_37558,N_24307,N_23859);
xor U37559 (N_37559,N_21743,N_27422);
nor U37560 (N_37560,N_29389,N_21536);
nand U37561 (N_37561,N_28747,N_20080);
xnor U37562 (N_37562,N_28161,N_28023);
xor U37563 (N_37563,N_25978,N_25316);
and U37564 (N_37564,N_28164,N_25535);
nand U37565 (N_37565,N_26321,N_26166);
or U37566 (N_37566,N_25370,N_24336);
nand U37567 (N_37567,N_28825,N_23003);
or U37568 (N_37568,N_29687,N_26534);
nor U37569 (N_37569,N_28432,N_27719);
nor U37570 (N_37570,N_20608,N_28924);
nand U37571 (N_37571,N_28298,N_26667);
and U37572 (N_37572,N_24255,N_26434);
or U37573 (N_37573,N_24607,N_25852);
xnor U37574 (N_37574,N_24301,N_28424);
xnor U37575 (N_37575,N_29079,N_29821);
nand U37576 (N_37576,N_21496,N_29390);
and U37577 (N_37577,N_22852,N_20401);
nand U37578 (N_37578,N_28093,N_27528);
or U37579 (N_37579,N_22009,N_21180);
xor U37580 (N_37580,N_29375,N_25353);
xor U37581 (N_37581,N_22457,N_23226);
nor U37582 (N_37582,N_20092,N_23865);
and U37583 (N_37583,N_29633,N_21878);
xor U37584 (N_37584,N_27395,N_22054);
and U37585 (N_37585,N_26380,N_26963);
xnor U37586 (N_37586,N_22479,N_27270);
xnor U37587 (N_37587,N_29431,N_24017);
or U37588 (N_37588,N_26282,N_25712);
nand U37589 (N_37589,N_22558,N_24296);
xnor U37590 (N_37590,N_20420,N_28828);
and U37591 (N_37591,N_24613,N_21995);
and U37592 (N_37592,N_26182,N_28691);
and U37593 (N_37593,N_25481,N_26839);
xnor U37594 (N_37594,N_27364,N_28994);
xor U37595 (N_37595,N_21697,N_29439);
nor U37596 (N_37596,N_28495,N_23865);
nand U37597 (N_37597,N_23818,N_21591);
nand U37598 (N_37598,N_29929,N_26749);
and U37599 (N_37599,N_24737,N_27843);
nor U37600 (N_37600,N_23354,N_29460);
nor U37601 (N_37601,N_20217,N_20031);
and U37602 (N_37602,N_28409,N_21906);
nor U37603 (N_37603,N_29287,N_27147);
or U37604 (N_37604,N_26969,N_23079);
and U37605 (N_37605,N_23378,N_24218);
xnor U37606 (N_37606,N_27161,N_21791);
xor U37607 (N_37607,N_20925,N_22564);
nor U37608 (N_37608,N_20027,N_29550);
nor U37609 (N_37609,N_29511,N_29896);
nand U37610 (N_37610,N_23326,N_21105);
xnor U37611 (N_37611,N_23510,N_26312);
and U37612 (N_37612,N_21135,N_20170);
nand U37613 (N_37613,N_25949,N_29291);
nand U37614 (N_37614,N_21314,N_28988);
nand U37615 (N_37615,N_25495,N_24067);
nor U37616 (N_37616,N_29184,N_25179);
or U37617 (N_37617,N_28796,N_29275);
or U37618 (N_37618,N_25183,N_27000);
xnor U37619 (N_37619,N_20476,N_26770);
and U37620 (N_37620,N_26605,N_28922);
nand U37621 (N_37621,N_24121,N_28225);
nor U37622 (N_37622,N_25840,N_28914);
or U37623 (N_37623,N_25853,N_22256);
xnor U37624 (N_37624,N_24749,N_22005);
nor U37625 (N_37625,N_29949,N_22998);
and U37626 (N_37626,N_26380,N_28320);
nand U37627 (N_37627,N_24783,N_21043);
nor U37628 (N_37628,N_26475,N_25254);
or U37629 (N_37629,N_20342,N_22161);
nand U37630 (N_37630,N_29618,N_27032);
or U37631 (N_37631,N_26721,N_23314);
or U37632 (N_37632,N_23470,N_26972);
and U37633 (N_37633,N_26892,N_25670);
nor U37634 (N_37634,N_29796,N_21469);
or U37635 (N_37635,N_25900,N_22585);
and U37636 (N_37636,N_26828,N_22435);
and U37637 (N_37637,N_26333,N_29307);
nand U37638 (N_37638,N_27901,N_28729);
or U37639 (N_37639,N_25219,N_26471);
nand U37640 (N_37640,N_26673,N_25403);
or U37641 (N_37641,N_25111,N_25584);
or U37642 (N_37642,N_20099,N_27698);
or U37643 (N_37643,N_21774,N_24843);
nor U37644 (N_37644,N_26139,N_21478);
or U37645 (N_37645,N_20517,N_27632);
xnor U37646 (N_37646,N_23487,N_23309);
nand U37647 (N_37647,N_25073,N_29744);
nor U37648 (N_37648,N_26990,N_23692);
and U37649 (N_37649,N_21733,N_22114);
and U37650 (N_37650,N_26557,N_24303);
and U37651 (N_37651,N_23636,N_21402);
nand U37652 (N_37652,N_27855,N_24359);
and U37653 (N_37653,N_20911,N_23168);
nand U37654 (N_37654,N_29469,N_24156);
nand U37655 (N_37655,N_28764,N_25874);
xor U37656 (N_37656,N_21670,N_25976);
and U37657 (N_37657,N_24038,N_20361);
xor U37658 (N_37658,N_26698,N_29709);
xor U37659 (N_37659,N_25846,N_23137);
nand U37660 (N_37660,N_25535,N_28877);
xnor U37661 (N_37661,N_25741,N_21490);
nand U37662 (N_37662,N_23138,N_22329);
and U37663 (N_37663,N_29354,N_20953);
nand U37664 (N_37664,N_20692,N_26387);
or U37665 (N_37665,N_22264,N_27666);
xor U37666 (N_37666,N_24977,N_21573);
or U37667 (N_37667,N_21302,N_22388);
and U37668 (N_37668,N_21452,N_24455);
nor U37669 (N_37669,N_22131,N_24400);
nand U37670 (N_37670,N_23141,N_26179);
or U37671 (N_37671,N_22734,N_24531);
and U37672 (N_37672,N_29368,N_23471);
nor U37673 (N_37673,N_28548,N_21585);
or U37674 (N_37674,N_25029,N_25546);
nor U37675 (N_37675,N_25899,N_22675);
nor U37676 (N_37676,N_29272,N_24699);
nor U37677 (N_37677,N_21045,N_20622);
or U37678 (N_37678,N_21246,N_29840);
nor U37679 (N_37679,N_28878,N_24080);
xor U37680 (N_37680,N_26299,N_21864);
nand U37681 (N_37681,N_23515,N_21103);
or U37682 (N_37682,N_24229,N_28128);
xor U37683 (N_37683,N_26106,N_29756);
or U37684 (N_37684,N_25619,N_24120);
xnor U37685 (N_37685,N_20525,N_25464);
and U37686 (N_37686,N_25946,N_24521);
nand U37687 (N_37687,N_25128,N_25224);
nand U37688 (N_37688,N_24781,N_21567);
and U37689 (N_37689,N_26827,N_24860);
nand U37690 (N_37690,N_26019,N_27581);
nand U37691 (N_37691,N_27911,N_23966);
nor U37692 (N_37692,N_21100,N_29051);
nor U37693 (N_37693,N_21850,N_28564);
xor U37694 (N_37694,N_26640,N_27190);
or U37695 (N_37695,N_20736,N_29801);
and U37696 (N_37696,N_29315,N_22272);
and U37697 (N_37697,N_24016,N_27920);
and U37698 (N_37698,N_21186,N_25188);
or U37699 (N_37699,N_27286,N_24310);
or U37700 (N_37700,N_21238,N_28097);
nor U37701 (N_37701,N_25441,N_29259);
nand U37702 (N_37702,N_24335,N_24023);
xor U37703 (N_37703,N_29277,N_27594);
nor U37704 (N_37704,N_23176,N_22697);
xnor U37705 (N_37705,N_24768,N_24495);
xor U37706 (N_37706,N_23973,N_23954);
xnor U37707 (N_37707,N_29577,N_24527);
nor U37708 (N_37708,N_26376,N_28732);
and U37709 (N_37709,N_22215,N_21616);
or U37710 (N_37710,N_27472,N_21245);
and U37711 (N_37711,N_24780,N_23963);
nand U37712 (N_37712,N_21173,N_20847);
and U37713 (N_37713,N_27793,N_23414);
xnor U37714 (N_37714,N_27508,N_27251);
xnor U37715 (N_37715,N_21584,N_23365);
and U37716 (N_37716,N_20546,N_28391);
nor U37717 (N_37717,N_29043,N_28159);
nor U37718 (N_37718,N_25386,N_23426);
and U37719 (N_37719,N_23200,N_25762);
nor U37720 (N_37720,N_28121,N_21674);
nand U37721 (N_37721,N_27737,N_28880);
nand U37722 (N_37722,N_25371,N_25182);
nor U37723 (N_37723,N_23881,N_27376);
or U37724 (N_37724,N_20857,N_27162);
and U37725 (N_37725,N_29581,N_26365);
nor U37726 (N_37726,N_28245,N_29404);
and U37727 (N_37727,N_22373,N_24606);
and U37728 (N_37728,N_25479,N_22724);
or U37729 (N_37729,N_23907,N_20234);
nor U37730 (N_37730,N_27319,N_21322);
nand U37731 (N_37731,N_27645,N_20248);
nand U37732 (N_37732,N_22911,N_26760);
or U37733 (N_37733,N_28450,N_22899);
nand U37734 (N_37734,N_25579,N_24508);
or U37735 (N_37735,N_25052,N_24226);
or U37736 (N_37736,N_20681,N_21146);
and U37737 (N_37737,N_20798,N_28173);
and U37738 (N_37738,N_26570,N_28092);
or U37739 (N_37739,N_29922,N_22749);
nand U37740 (N_37740,N_25158,N_26980);
nand U37741 (N_37741,N_23721,N_27183);
nor U37742 (N_37742,N_27496,N_23193);
or U37743 (N_37743,N_29461,N_24076);
and U37744 (N_37744,N_21996,N_21438);
or U37745 (N_37745,N_27860,N_26967);
and U37746 (N_37746,N_27517,N_20087);
or U37747 (N_37747,N_24906,N_29803);
xor U37748 (N_37748,N_29325,N_29912);
nor U37749 (N_37749,N_29870,N_26538);
and U37750 (N_37750,N_20530,N_27158);
nor U37751 (N_37751,N_28479,N_26357);
nand U37752 (N_37752,N_26609,N_28094);
nand U37753 (N_37753,N_23665,N_23679);
nor U37754 (N_37754,N_23551,N_20309);
or U37755 (N_37755,N_20937,N_26988);
xor U37756 (N_37756,N_26439,N_21425);
nand U37757 (N_37757,N_27338,N_29272);
nor U37758 (N_37758,N_29124,N_22847);
xnor U37759 (N_37759,N_28436,N_22848);
nand U37760 (N_37760,N_22941,N_29981);
or U37761 (N_37761,N_21075,N_22147);
and U37762 (N_37762,N_22240,N_23459);
or U37763 (N_37763,N_26894,N_26068);
nor U37764 (N_37764,N_23618,N_29091);
and U37765 (N_37765,N_28764,N_29160);
nand U37766 (N_37766,N_22667,N_21546);
and U37767 (N_37767,N_28275,N_25811);
nor U37768 (N_37768,N_26364,N_24314);
nor U37769 (N_37769,N_28995,N_26974);
or U37770 (N_37770,N_21399,N_24789);
nor U37771 (N_37771,N_29362,N_22042);
nor U37772 (N_37772,N_26112,N_25304);
xor U37773 (N_37773,N_20374,N_25841);
nand U37774 (N_37774,N_24173,N_24771);
or U37775 (N_37775,N_20939,N_28261);
nor U37776 (N_37776,N_22233,N_29040);
nand U37777 (N_37777,N_23990,N_27529);
xnor U37778 (N_37778,N_20866,N_21400);
xor U37779 (N_37779,N_22022,N_21807);
and U37780 (N_37780,N_28760,N_22704);
and U37781 (N_37781,N_29074,N_20275);
nor U37782 (N_37782,N_29960,N_29911);
nor U37783 (N_37783,N_24031,N_27472);
or U37784 (N_37784,N_27680,N_28432);
nand U37785 (N_37785,N_29707,N_23754);
and U37786 (N_37786,N_26345,N_25410);
and U37787 (N_37787,N_22065,N_23844);
or U37788 (N_37788,N_27217,N_21272);
xnor U37789 (N_37789,N_27089,N_29609);
nand U37790 (N_37790,N_29511,N_23945);
nand U37791 (N_37791,N_25256,N_20476);
xor U37792 (N_37792,N_28722,N_25029);
nand U37793 (N_37793,N_21662,N_27299);
xor U37794 (N_37794,N_24350,N_24259);
or U37795 (N_37795,N_20646,N_29241);
or U37796 (N_37796,N_20748,N_28618);
or U37797 (N_37797,N_27068,N_20342);
and U37798 (N_37798,N_20340,N_25133);
and U37799 (N_37799,N_24198,N_21942);
and U37800 (N_37800,N_25854,N_23602);
nand U37801 (N_37801,N_26814,N_27156);
xor U37802 (N_37802,N_27729,N_24258);
nand U37803 (N_37803,N_27739,N_27841);
or U37804 (N_37804,N_23195,N_26690);
and U37805 (N_37805,N_21685,N_26863);
nand U37806 (N_37806,N_28134,N_26429);
nor U37807 (N_37807,N_28335,N_27401);
nor U37808 (N_37808,N_22998,N_26927);
nand U37809 (N_37809,N_22661,N_28098);
nor U37810 (N_37810,N_22120,N_23623);
or U37811 (N_37811,N_21879,N_23850);
or U37812 (N_37812,N_27386,N_26595);
nand U37813 (N_37813,N_20932,N_23812);
and U37814 (N_37814,N_26147,N_20561);
nand U37815 (N_37815,N_27273,N_21214);
and U37816 (N_37816,N_21041,N_28015);
nor U37817 (N_37817,N_29311,N_20619);
nand U37818 (N_37818,N_20123,N_28706);
nor U37819 (N_37819,N_29793,N_24801);
nor U37820 (N_37820,N_21583,N_28050);
xor U37821 (N_37821,N_27480,N_22368);
xor U37822 (N_37822,N_28840,N_22547);
nand U37823 (N_37823,N_21163,N_24183);
or U37824 (N_37824,N_22762,N_22663);
xor U37825 (N_37825,N_24903,N_25586);
and U37826 (N_37826,N_21976,N_27196);
xor U37827 (N_37827,N_26045,N_25507);
or U37828 (N_37828,N_29349,N_24147);
xnor U37829 (N_37829,N_22391,N_21530);
and U37830 (N_37830,N_27068,N_21633);
xnor U37831 (N_37831,N_29469,N_20958);
and U37832 (N_37832,N_25717,N_21615);
xnor U37833 (N_37833,N_22191,N_24943);
nand U37834 (N_37834,N_24171,N_21276);
nor U37835 (N_37835,N_25885,N_23041);
and U37836 (N_37836,N_20036,N_28552);
nor U37837 (N_37837,N_22798,N_29710);
or U37838 (N_37838,N_26806,N_20525);
or U37839 (N_37839,N_26424,N_26985);
and U37840 (N_37840,N_22471,N_24126);
xnor U37841 (N_37841,N_27037,N_29671);
or U37842 (N_37842,N_26801,N_21468);
and U37843 (N_37843,N_26092,N_27814);
nor U37844 (N_37844,N_22063,N_28353);
or U37845 (N_37845,N_25865,N_20169);
nand U37846 (N_37846,N_22661,N_21447);
xnor U37847 (N_37847,N_26327,N_21808);
xor U37848 (N_37848,N_27117,N_20561);
nor U37849 (N_37849,N_27003,N_24628);
and U37850 (N_37850,N_29960,N_27534);
xor U37851 (N_37851,N_20441,N_26460);
xor U37852 (N_37852,N_28157,N_25045);
or U37853 (N_37853,N_25415,N_25189);
and U37854 (N_37854,N_25966,N_20870);
xnor U37855 (N_37855,N_26024,N_24241);
xnor U37856 (N_37856,N_28668,N_21523);
nand U37857 (N_37857,N_21369,N_23067);
xnor U37858 (N_37858,N_26897,N_25386);
nor U37859 (N_37859,N_25153,N_24638);
or U37860 (N_37860,N_27295,N_20392);
and U37861 (N_37861,N_26360,N_28369);
xor U37862 (N_37862,N_23549,N_20577);
or U37863 (N_37863,N_27844,N_25389);
nand U37864 (N_37864,N_26554,N_22909);
xnor U37865 (N_37865,N_21285,N_20099);
xor U37866 (N_37866,N_22475,N_28559);
nor U37867 (N_37867,N_25104,N_26509);
or U37868 (N_37868,N_28089,N_29368);
nand U37869 (N_37869,N_29929,N_23400);
and U37870 (N_37870,N_26859,N_20916);
xor U37871 (N_37871,N_26276,N_27108);
or U37872 (N_37872,N_20360,N_29723);
xor U37873 (N_37873,N_27156,N_27999);
nand U37874 (N_37874,N_21836,N_25634);
nand U37875 (N_37875,N_24087,N_21984);
nor U37876 (N_37876,N_26580,N_23779);
or U37877 (N_37877,N_26078,N_27547);
nand U37878 (N_37878,N_23384,N_28302);
or U37879 (N_37879,N_22133,N_22467);
and U37880 (N_37880,N_20729,N_20988);
nand U37881 (N_37881,N_27500,N_21884);
xor U37882 (N_37882,N_27316,N_27711);
xor U37883 (N_37883,N_23477,N_25849);
xor U37884 (N_37884,N_26177,N_27554);
nand U37885 (N_37885,N_21510,N_26064);
nor U37886 (N_37886,N_23986,N_25963);
or U37887 (N_37887,N_29889,N_24941);
and U37888 (N_37888,N_29571,N_24311);
nor U37889 (N_37889,N_21031,N_29891);
xnor U37890 (N_37890,N_29017,N_26812);
nand U37891 (N_37891,N_26640,N_25332);
nor U37892 (N_37892,N_21847,N_24738);
or U37893 (N_37893,N_26183,N_26229);
xor U37894 (N_37894,N_27426,N_25268);
and U37895 (N_37895,N_28454,N_28648);
nor U37896 (N_37896,N_23382,N_22001);
nand U37897 (N_37897,N_20754,N_20116);
nand U37898 (N_37898,N_20952,N_20211);
nand U37899 (N_37899,N_20970,N_21432);
xor U37900 (N_37900,N_27726,N_29201);
nand U37901 (N_37901,N_26050,N_24007);
or U37902 (N_37902,N_20462,N_26723);
xnor U37903 (N_37903,N_20026,N_29959);
or U37904 (N_37904,N_26025,N_29009);
or U37905 (N_37905,N_23206,N_24989);
nor U37906 (N_37906,N_21254,N_26880);
or U37907 (N_37907,N_26525,N_27798);
xor U37908 (N_37908,N_24319,N_22979);
nor U37909 (N_37909,N_25318,N_24742);
or U37910 (N_37910,N_24311,N_25481);
nor U37911 (N_37911,N_22315,N_25539);
and U37912 (N_37912,N_25495,N_20900);
xnor U37913 (N_37913,N_23647,N_28492);
xnor U37914 (N_37914,N_25203,N_21332);
and U37915 (N_37915,N_24817,N_29079);
nor U37916 (N_37916,N_28178,N_23066);
and U37917 (N_37917,N_21076,N_21808);
or U37918 (N_37918,N_20326,N_28246);
or U37919 (N_37919,N_24707,N_25544);
or U37920 (N_37920,N_26648,N_26129);
or U37921 (N_37921,N_29331,N_26382);
xnor U37922 (N_37922,N_21410,N_25541);
and U37923 (N_37923,N_25583,N_21214);
or U37924 (N_37924,N_28240,N_22656);
and U37925 (N_37925,N_26644,N_29170);
and U37926 (N_37926,N_26685,N_27925);
xor U37927 (N_37927,N_27830,N_20893);
nand U37928 (N_37928,N_21517,N_28463);
or U37929 (N_37929,N_25583,N_23536);
and U37930 (N_37930,N_23317,N_20014);
and U37931 (N_37931,N_22073,N_26147);
or U37932 (N_37932,N_27809,N_24403);
or U37933 (N_37933,N_28300,N_25863);
xnor U37934 (N_37934,N_23353,N_20457);
nand U37935 (N_37935,N_23306,N_26342);
or U37936 (N_37936,N_23249,N_29243);
or U37937 (N_37937,N_25442,N_29070);
nor U37938 (N_37938,N_25026,N_26712);
xor U37939 (N_37939,N_25943,N_29029);
nor U37940 (N_37940,N_21965,N_21616);
xor U37941 (N_37941,N_29112,N_23134);
nand U37942 (N_37942,N_28894,N_20009);
and U37943 (N_37943,N_27058,N_28363);
xnor U37944 (N_37944,N_20319,N_24475);
or U37945 (N_37945,N_28977,N_26590);
nand U37946 (N_37946,N_22984,N_22169);
or U37947 (N_37947,N_29337,N_23450);
nor U37948 (N_37948,N_26405,N_24746);
or U37949 (N_37949,N_24560,N_28696);
and U37950 (N_37950,N_21943,N_23622);
nand U37951 (N_37951,N_29087,N_23511);
or U37952 (N_37952,N_23046,N_25416);
nand U37953 (N_37953,N_20898,N_24437);
xor U37954 (N_37954,N_26536,N_23959);
or U37955 (N_37955,N_29034,N_26622);
xor U37956 (N_37956,N_20984,N_27347);
xnor U37957 (N_37957,N_23023,N_29558);
or U37958 (N_37958,N_24366,N_21811);
or U37959 (N_37959,N_28995,N_22492);
nand U37960 (N_37960,N_28848,N_23209);
and U37961 (N_37961,N_29138,N_21244);
xor U37962 (N_37962,N_24119,N_22593);
nor U37963 (N_37963,N_27510,N_29380);
nand U37964 (N_37964,N_28687,N_28360);
and U37965 (N_37965,N_27789,N_27453);
nor U37966 (N_37966,N_23029,N_21354);
and U37967 (N_37967,N_24727,N_23034);
nand U37968 (N_37968,N_27135,N_27432);
nor U37969 (N_37969,N_20258,N_28941);
or U37970 (N_37970,N_24342,N_27716);
nor U37971 (N_37971,N_29543,N_23083);
nor U37972 (N_37972,N_21771,N_22555);
or U37973 (N_37973,N_20507,N_22020);
nor U37974 (N_37974,N_27820,N_27234);
xnor U37975 (N_37975,N_22554,N_22820);
and U37976 (N_37976,N_28698,N_22727);
nor U37977 (N_37977,N_27799,N_24064);
xor U37978 (N_37978,N_21542,N_21201);
nand U37979 (N_37979,N_22127,N_27025);
and U37980 (N_37980,N_25679,N_21531);
and U37981 (N_37981,N_25615,N_29906);
nor U37982 (N_37982,N_29699,N_25126);
nor U37983 (N_37983,N_27526,N_22771);
nor U37984 (N_37984,N_26405,N_26874);
xor U37985 (N_37985,N_22333,N_28124);
and U37986 (N_37986,N_26307,N_20474);
and U37987 (N_37987,N_27103,N_28085);
nand U37988 (N_37988,N_23311,N_23540);
or U37989 (N_37989,N_26801,N_27798);
nor U37990 (N_37990,N_24731,N_25849);
xor U37991 (N_37991,N_23771,N_21491);
or U37992 (N_37992,N_29602,N_22204);
and U37993 (N_37993,N_25494,N_22572);
xor U37994 (N_37994,N_25866,N_28405);
and U37995 (N_37995,N_28030,N_23672);
nor U37996 (N_37996,N_24723,N_21278);
xnor U37997 (N_37997,N_29334,N_24782);
and U37998 (N_37998,N_28163,N_20350);
and U37999 (N_37999,N_23012,N_24951);
nand U38000 (N_38000,N_22343,N_28059);
or U38001 (N_38001,N_25515,N_26896);
nor U38002 (N_38002,N_24166,N_26675);
nand U38003 (N_38003,N_24835,N_25813);
and U38004 (N_38004,N_26295,N_25016);
xor U38005 (N_38005,N_21744,N_23621);
nand U38006 (N_38006,N_25270,N_29443);
nor U38007 (N_38007,N_29133,N_20144);
or U38008 (N_38008,N_22020,N_26860);
xnor U38009 (N_38009,N_27486,N_22438);
and U38010 (N_38010,N_23109,N_20218);
nor U38011 (N_38011,N_21500,N_22515);
nor U38012 (N_38012,N_24453,N_22444);
or U38013 (N_38013,N_29082,N_26488);
xor U38014 (N_38014,N_29323,N_23403);
nor U38015 (N_38015,N_24975,N_21406);
xnor U38016 (N_38016,N_28610,N_23422);
or U38017 (N_38017,N_27824,N_20837);
nand U38018 (N_38018,N_23610,N_29512);
nand U38019 (N_38019,N_21120,N_24955);
and U38020 (N_38020,N_26019,N_25407);
xnor U38021 (N_38021,N_24718,N_22842);
and U38022 (N_38022,N_29545,N_24792);
xnor U38023 (N_38023,N_21200,N_23141);
nand U38024 (N_38024,N_20375,N_29382);
nor U38025 (N_38025,N_27292,N_27974);
or U38026 (N_38026,N_22079,N_23573);
xnor U38027 (N_38027,N_26276,N_26094);
and U38028 (N_38028,N_29277,N_27064);
and U38029 (N_38029,N_20950,N_24617);
xnor U38030 (N_38030,N_28356,N_20847);
nand U38031 (N_38031,N_24092,N_20182);
xnor U38032 (N_38032,N_27619,N_28864);
xor U38033 (N_38033,N_29090,N_23901);
xor U38034 (N_38034,N_21331,N_23615);
and U38035 (N_38035,N_21555,N_20183);
or U38036 (N_38036,N_29845,N_25263);
and U38037 (N_38037,N_22861,N_23721);
and U38038 (N_38038,N_28333,N_24850);
or U38039 (N_38039,N_20894,N_24151);
and U38040 (N_38040,N_20803,N_27487);
and U38041 (N_38041,N_24694,N_28848);
xnor U38042 (N_38042,N_25748,N_29985);
xnor U38043 (N_38043,N_28983,N_23631);
xnor U38044 (N_38044,N_24992,N_26061);
or U38045 (N_38045,N_28299,N_29453);
or U38046 (N_38046,N_23612,N_24516);
or U38047 (N_38047,N_22841,N_28383);
xnor U38048 (N_38048,N_25743,N_25614);
or U38049 (N_38049,N_24588,N_25996);
and U38050 (N_38050,N_26427,N_23358);
nor U38051 (N_38051,N_29763,N_25618);
and U38052 (N_38052,N_24397,N_24697);
or U38053 (N_38053,N_28653,N_23540);
and U38054 (N_38054,N_23708,N_25442);
or U38055 (N_38055,N_21864,N_27739);
and U38056 (N_38056,N_27710,N_20421);
nor U38057 (N_38057,N_21557,N_29597);
and U38058 (N_38058,N_28009,N_26073);
or U38059 (N_38059,N_21139,N_20879);
nand U38060 (N_38060,N_21555,N_26023);
and U38061 (N_38061,N_22811,N_23683);
or U38062 (N_38062,N_20990,N_21405);
nand U38063 (N_38063,N_26306,N_29819);
xnor U38064 (N_38064,N_24668,N_28362);
xor U38065 (N_38065,N_25667,N_26824);
nor U38066 (N_38066,N_29756,N_24544);
xor U38067 (N_38067,N_26868,N_20614);
and U38068 (N_38068,N_26142,N_24061);
and U38069 (N_38069,N_20826,N_20155);
and U38070 (N_38070,N_24355,N_22626);
nand U38071 (N_38071,N_26684,N_23914);
xor U38072 (N_38072,N_20421,N_21440);
xnor U38073 (N_38073,N_28922,N_21104);
and U38074 (N_38074,N_27401,N_22326);
or U38075 (N_38075,N_25255,N_29999);
nor U38076 (N_38076,N_29648,N_24250);
xor U38077 (N_38077,N_26682,N_28880);
nand U38078 (N_38078,N_24253,N_20210);
nand U38079 (N_38079,N_20951,N_22501);
or U38080 (N_38080,N_25597,N_29740);
xnor U38081 (N_38081,N_22150,N_28498);
xor U38082 (N_38082,N_23037,N_21888);
nand U38083 (N_38083,N_20353,N_21990);
xor U38084 (N_38084,N_22627,N_29534);
and U38085 (N_38085,N_24521,N_28382);
nand U38086 (N_38086,N_29107,N_29992);
nand U38087 (N_38087,N_28797,N_20037);
nand U38088 (N_38088,N_22346,N_27363);
or U38089 (N_38089,N_29910,N_20802);
xnor U38090 (N_38090,N_28190,N_20557);
xor U38091 (N_38091,N_24730,N_23130);
and U38092 (N_38092,N_20111,N_27729);
nand U38093 (N_38093,N_21493,N_23767);
xor U38094 (N_38094,N_23601,N_24905);
xnor U38095 (N_38095,N_21582,N_29886);
and U38096 (N_38096,N_27568,N_22254);
nand U38097 (N_38097,N_23247,N_26800);
or U38098 (N_38098,N_20664,N_24378);
nor U38099 (N_38099,N_21080,N_22765);
nand U38100 (N_38100,N_22303,N_28710);
or U38101 (N_38101,N_23803,N_29830);
nand U38102 (N_38102,N_26248,N_28310);
xnor U38103 (N_38103,N_24277,N_20551);
nor U38104 (N_38104,N_27867,N_20730);
nor U38105 (N_38105,N_22307,N_22435);
and U38106 (N_38106,N_25118,N_20268);
or U38107 (N_38107,N_20217,N_22170);
xor U38108 (N_38108,N_25689,N_28265);
xnor U38109 (N_38109,N_28531,N_23639);
or U38110 (N_38110,N_25982,N_27946);
nor U38111 (N_38111,N_26924,N_24377);
or U38112 (N_38112,N_24440,N_22721);
xnor U38113 (N_38113,N_27724,N_29926);
or U38114 (N_38114,N_26370,N_23223);
or U38115 (N_38115,N_20914,N_25199);
nand U38116 (N_38116,N_25315,N_23361);
and U38117 (N_38117,N_23946,N_28325);
nand U38118 (N_38118,N_26095,N_27398);
nor U38119 (N_38119,N_24907,N_29558);
and U38120 (N_38120,N_24213,N_22537);
nor U38121 (N_38121,N_25973,N_24198);
and U38122 (N_38122,N_22972,N_24353);
xor U38123 (N_38123,N_29003,N_24688);
or U38124 (N_38124,N_21267,N_27004);
nand U38125 (N_38125,N_22379,N_20802);
nand U38126 (N_38126,N_29291,N_23699);
or U38127 (N_38127,N_27746,N_24724);
and U38128 (N_38128,N_21093,N_29817);
nor U38129 (N_38129,N_28564,N_26243);
xnor U38130 (N_38130,N_28463,N_23795);
and U38131 (N_38131,N_29277,N_24251);
xnor U38132 (N_38132,N_24405,N_23075);
nor U38133 (N_38133,N_21221,N_23866);
or U38134 (N_38134,N_25401,N_22176);
xnor U38135 (N_38135,N_29085,N_26966);
and U38136 (N_38136,N_26910,N_29912);
nor U38137 (N_38137,N_23676,N_29864);
nand U38138 (N_38138,N_27451,N_27671);
or U38139 (N_38139,N_20677,N_22553);
xor U38140 (N_38140,N_27089,N_25215);
xnor U38141 (N_38141,N_26427,N_23218);
xnor U38142 (N_38142,N_26082,N_29519);
nand U38143 (N_38143,N_24397,N_23489);
and U38144 (N_38144,N_27953,N_21127);
xor U38145 (N_38145,N_20352,N_24151);
and U38146 (N_38146,N_24825,N_27441);
or U38147 (N_38147,N_29401,N_21449);
xnor U38148 (N_38148,N_22341,N_26831);
nor U38149 (N_38149,N_20370,N_21921);
nand U38150 (N_38150,N_23113,N_26412);
and U38151 (N_38151,N_27968,N_25026);
and U38152 (N_38152,N_22154,N_22727);
nand U38153 (N_38153,N_21840,N_22929);
xor U38154 (N_38154,N_22967,N_29392);
or U38155 (N_38155,N_25604,N_23702);
xnor U38156 (N_38156,N_26587,N_27979);
nor U38157 (N_38157,N_28571,N_28706);
xor U38158 (N_38158,N_26008,N_22539);
nand U38159 (N_38159,N_27345,N_25188);
xnor U38160 (N_38160,N_29780,N_28120);
nand U38161 (N_38161,N_26819,N_24288);
or U38162 (N_38162,N_20294,N_20893);
nand U38163 (N_38163,N_24148,N_23272);
nor U38164 (N_38164,N_21748,N_28099);
or U38165 (N_38165,N_27444,N_29259);
nand U38166 (N_38166,N_28647,N_21240);
xnor U38167 (N_38167,N_20894,N_21926);
or U38168 (N_38168,N_23673,N_21134);
or U38169 (N_38169,N_24244,N_20668);
nor U38170 (N_38170,N_22107,N_25737);
nand U38171 (N_38171,N_25216,N_28681);
xor U38172 (N_38172,N_28581,N_24376);
nand U38173 (N_38173,N_20635,N_20643);
xnor U38174 (N_38174,N_20758,N_24922);
nand U38175 (N_38175,N_24897,N_20017);
nand U38176 (N_38176,N_29233,N_25940);
and U38177 (N_38177,N_27359,N_24224);
xor U38178 (N_38178,N_28289,N_26240);
xnor U38179 (N_38179,N_20871,N_24079);
nor U38180 (N_38180,N_26467,N_22306);
xor U38181 (N_38181,N_26490,N_20557);
nand U38182 (N_38182,N_28827,N_23157);
or U38183 (N_38183,N_25331,N_20439);
nor U38184 (N_38184,N_29320,N_26445);
or U38185 (N_38185,N_21547,N_22367);
nor U38186 (N_38186,N_22736,N_20692);
nor U38187 (N_38187,N_26387,N_29166);
nand U38188 (N_38188,N_26915,N_27096);
and U38189 (N_38189,N_20536,N_23876);
nor U38190 (N_38190,N_27194,N_25432);
nor U38191 (N_38191,N_22793,N_25318);
and U38192 (N_38192,N_23281,N_22288);
nand U38193 (N_38193,N_21962,N_29030);
nor U38194 (N_38194,N_28345,N_23776);
xnor U38195 (N_38195,N_28139,N_20458);
and U38196 (N_38196,N_27368,N_20870);
or U38197 (N_38197,N_25588,N_21321);
or U38198 (N_38198,N_20056,N_29099);
nor U38199 (N_38199,N_27219,N_24330);
nor U38200 (N_38200,N_29971,N_21763);
nor U38201 (N_38201,N_23150,N_24381);
and U38202 (N_38202,N_28489,N_27005);
or U38203 (N_38203,N_27479,N_26297);
and U38204 (N_38204,N_26623,N_24891);
xor U38205 (N_38205,N_28714,N_23480);
xor U38206 (N_38206,N_29959,N_23245);
and U38207 (N_38207,N_23753,N_25127);
nor U38208 (N_38208,N_24801,N_21773);
nand U38209 (N_38209,N_23079,N_26476);
or U38210 (N_38210,N_29560,N_28573);
or U38211 (N_38211,N_23260,N_25010);
and U38212 (N_38212,N_26237,N_21279);
and U38213 (N_38213,N_29746,N_29424);
and U38214 (N_38214,N_23275,N_22238);
or U38215 (N_38215,N_27154,N_20370);
and U38216 (N_38216,N_20454,N_25308);
and U38217 (N_38217,N_22133,N_24420);
xor U38218 (N_38218,N_20622,N_21837);
nand U38219 (N_38219,N_28016,N_26990);
and U38220 (N_38220,N_29003,N_23608);
xor U38221 (N_38221,N_25840,N_21542);
nor U38222 (N_38222,N_25529,N_25816);
and U38223 (N_38223,N_28396,N_27876);
nand U38224 (N_38224,N_20092,N_29892);
nor U38225 (N_38225,N_22104,N_23122);
xnor U38226 (N_38226,N_23232,N_25687);
or U38227 (N_38227,N_26582,N_29608);
and U38228 (N_38228,N_24653,N_24435);
xnor U38229 (N_38229,N_29542,N_20374);
or U38230 (N_38230,N_20759,N_22847);
nand U38231 (N_38231,N_25535,N_20211);
nor U38232 (N_38232,N_26232,N_20251);
and U38233 (N_38233,N_23285,N_26591);
xor U38234 (N_38234,N_28328,N_27961);
xor U38235 (N_38235,N_28646,N_21718);
or U38236 (N_38236,N_22933,N_27562);
nand U38237 (N_38237,N_22225,N_23032);
xor U38238 (N_38238,N_22435,N_20381);
or U38239 (N_38239,N_22841,N_24548);
and U38240 (N_38240,N_23278,N_28783);
nand U38241 (N_38241,N_26397,N_25074);
nand U38242 (N_38242,N_25530,N_23940);
nand U38243 (N_38243,N_23503,N_20267);
nand U38244 (N_38244,N_24336,N_21447);
xor U38245 (N_38245,N_24044,N_21023);
or U38246 (N_38246,N_23572,N_20415);
nand U38247 (N_38247,N_24882,N_28343);
nor U38248 (N_38248,N_24115,N_28283);
nand U38249 (N_38249,N_24736,N_21565);
nand U38250 (N_38250,N_24192,N_26416);
nand U38251 (N_38251,N_22986,N_25411);
or U38252 (N_38252,N_23368,N_23178);
xor U38253 (N_38253,N_20990,N_24034);
or U38254 (N_38254,N_25295,N_23426);
nand U38255 (N_38255,N_27622,N_29038);
nor U38256 (N_38256,N_21093,N_21416);
nand U38257 (N_38257,N_24055,N_27096);
or U38258 (N_38258,N_28251,N_22725);
xnor U38259 (N_38259,N_25993,N_22716);
nand U38260 (N_38260,N_20937,N_24810);
xor U38261 (N_38261,N_20407,N_23871);
and U38262 (N_38262,N_27678,N_21081);
and U38263 (N_38263,N_20385,N_28469);
nand U38264 (N_38264,N_22082,N_22042);
nand U38265 (N_38265,N_26680,N_21462);
and U38266 (N_38266,N_21860,N_21498);
or U38267 (N_38267,N_20348,N_26658);
nor U38268 (N_38268,N_29949,N_21581);
xor U38269 (N_38269,N_28440,N_21505);
xnor U38270 (N_38270,N_24704,N_26517);
xor U38271 (N_38271,N_22570,N_27446);
nand U38272 (N_38272,N_29290,N_28341);
nor U38273 (N_38273,N_21758,N_25500);
xnor U38274 (N_38274,N_29898,N_29931);
xor U38275 (N_38275,N_26988,N_24306);
and U38276 (N_38276,N_26507,N_25074);
xor U38277 (N_38277,N_22388,N_26366);
or U38278 (N_38278,N_28725,N_26852);
and U38279 (N_38279,N_22088,N_20835);
and U38280 (N_38280,N_24817,N_21969);
nor U38281 (N_38281,N_22095,N_29401);
and U38282 (N_38282,N_26109,N_21353);
nor U38283 (N_38283,N_24657,N_27470);
nor U38284 (N_38284,N_28581,N_28031);
nand U38285 (N_38285,N_25508,N_26993);
nand U38286 (N_38286,N_23963,N_21885);
nand U38287 (N_38287,N_24731,N_26284);
nand U38288 (N_38288,N_25318,N_22852);
nor U38289 (N_38289,N_21195,N_25884);
and U38290 (N_38290,N_29280,N_22441);
or U38291 (N_38291,N_28317,N_27659);
nand U38292 (N_38292,N_20802,N_20568);
and U38293 (N_38293,N_24290,N_20744);
and U38294 (N_38294,N_21603,N_23514);
and U38295 (N_38295,N_26340,N_29193);
nand U38296 (N_38296,N_22385,N_25553);
or U38297 (N_38297,N_23543,N_20203);
xor U38298 (N_38298,N_20345,N_23714);
or U38299 (N_38299,N_24449,N_26770);
or U38300 (N_38300,N_22892,N_22404);
xnor U38301 (N_38301,N_21847,N_27131);
or U38302 (N_38302,N_25354,N_25490);
xor U38303 (N_38303,N_23337,N_21595);
or U38304 (N_38304,N_22378,N_22840);
nor U38305 (N_38305,N_20105,N_23229);
nand U38306 (N_38306,N_27909,N_25367);
and U38307 (N_38307,N_20786,N_23598);
nand U38308 (N_38308,N_23943,N_25245);
and U38309 (N_38309,N_28585,N_23192);
nor U38310 (N_38310,N_23244,N_20522);
and U38311 (N_38311,N_24300,N_25759);
xnor U38312 (N_38312,N_28576,N_28591);
xnor U38313 (N_38313,N_25154,N_27996);
xnor U38314 (N_38314,N_26684,N_28584);
xnor U38315 (N_38315,N_27961,N_25038);
xnor U38316 (N_38316,N_29637,N_29268);
xor U38317 (N_38317,N_25421,N_29058);
xnor U38318 (N_38318,N_26080,N_29806);
nand U38319 (N_38319,N_27774,N_29333);
and U38320 (N_38320,N_22105,N_22690);
xor U38321 (N_38321,N_22823,N_24592);
nor U38322 (N_38322,N_25551,N_22436);
and U38323 (N_38323,N_23141,N_22822);
nor U38324 (N_38324,N_24845,N_29320);
nand U38325 (N_38325,N_25938,N_23672);
nand U38326 (N_38326,N_21822,N_22710);
nor U38327 (N_38327,N_21118,N_28737);
or U38328 (N_38328,N_25115,N_25384);
or U38329 (N_38329,N_21920,N_20119);
nor U38330 (N_38330,N_23920,N_20727);
xor U38331 (N_38331,N_22576,N_24691);
and U38332 (N_38332,N_20577,N_27787);
nor U38333 (N_38333,N_29142,N_24658);
and U38334 (N_38334,N_20621,N_28700);
or U38335 (N_38335,N_20800,N_29689);
nand U38336 (N_38336,N_28342,N_23379);
and U38337 (N_38337,N_23163,N_29106);
nor U38338 (N_38338,N_24595,N_21269);
or U38339 (N_38339,N_20680,N_22760);
or U38340 (N_38340,N_27370,N_21574);
and U38341 (N_38341,N_23145,N_28335);
or U38342 (N_38342,N_28655,N_24588);
and U38343 (N_38343,N_25883,N_23302);
nor U38344 (N_38344,N_22066,N_28908);
and U38345 (N_38345,N_21245,N_20103);
xnor U38346 (N_38346,N_20549,N_24449);
or U38347 (N_38347,N_22649,N_25960);
or U38348 (N_38348,N_23875,N_29053);
xor U38349 (N_38349,N_25665,N_26319);
xnor U38350 (N_38350,N_25792,N_23966);
nor U38351 (N_38351,N_25064,N_28258);
and U38352 (N_38352,N_21116,N_27625);
xor U38353 (N_38353,N_27691,N_26382);
or U38354 (N_38354,N_22952,N_26463);
and U38355 (N_38355,N_22545,N_24530);
nand U38356 (N_38356,N_20822,N_22008);
xnor U38357 (N_38357,N_27995,N_27900);
or U38358 (N_38358,N_20475,N_23005);
xnor U38359 (N_38359,N_24148,N_29915);
nor U38360 (N_38360,N_20882,N_27548);
and U38361 (N_38361,N_20549,N_29133);
or U38362 (N_38362,N_22865,N_27314);
and U38363 (N_38363,N_23877,N_24953);
or U38364 (N_38364,N_26221,N_20515);
nand U38365 (N_38365,N_21837,N_29899);
nor U38366 (N_38366,N_23405,N_26798);
nand U38367 (N_38367,N_28479,N_26189);
nor U38368 (N_38368,N_28245,N_22251);
and U38369 (N_38369,N_22807,N_23399);
or U38370 (N_38370,N_21035,N_29908);
or U38371 (N_38371,N_24348,N_25975);
nor U38372 (N_38372,N_26333,N_28391);
xnor U38373 (N_38373,N_24846,N_20356);
and U38374 (N_38374,N_24842,N_22634);
and U38375 (N_38375,N_20220,N_22637);
nand U38376 (N_38376,N_20101,N_26707);
xnor U38377 (N_38377,N_26779,N_25183);
nand U38378 (N_38378,N_29558,N_24609);
and U38379 (N_38379,N_22117,N_20403);
nand U38380 (N_38380,N_26708,N_29333);
xor U38381 (N_38381,N_26428,N_21831);
nor U38382 (N_38382,N_20478,N_26642);
and U38383 (N_38383,N_28754,N_28277);
or U38384 (N_38384,N_25551,N_28774);
nand U38385 (N_38385,N_24559,N_20435);
nor U38386 (N_38386,N_23693,N_24628);
and U38387 (N_38387,N_23383,N_27309);
and U38388 (N_38388,N_24816,N_25834);
and U38389 (N_38389,N_25586,N_21023);
or U38390 (N_38390,N_28500,N_26724);
or U38391 (N_38391,N_27194,N_26960);
and U38392 (N_38392,N_26019,N_23342);
nor U38393 (N_38393,N_28918,N_20822);
nand U38394 (N_38394,N_23585,N_24242);
nor U38395 (N_38395,N_22203,N_25755);
and U38396 (N_38396,N_20746,N_25467);
xnor U38397 (N_38397,N_24858,N_25300);
nand U38398 (N_38398,N_21588,N_28970);
nor U38399 (N_38399,N_23659,N_24526);
or U38400 (N_38400,N_27532,N_28389);
and U38401 (N_38401,N_24870,N_23491);
and U38402 (N_38402,N_21744,N_28328);
or U38403 (N_38403,N_28902,N_21262);
nand U38404 (N_38404,N_28564,N_24047);
nand U38405 (N_38405,N_29173,N_22913);
and U38406 (N_38406,N_24192,N_29677);
nand U38407 (N_38407,N_27924,N_28029);
and U38408 (N_38408,N_28215,N_23987);
or U38409 (N_38409,N_27945,N_22164);
nor U38410 (N_38410,N_27720,N_24720);
nand U38411 (N_38411,N_26037,N_21608);
xor U38412 (N_38412,N_28666,N_26799);
nand U38413 (N_38413,N_24022,N_20401);
nand U38414 (N_38414,N_23348,N_25321);
xnor U38415 (N_38415,N_29757,N_22618);
nand U38416 (N_38416,N_22782,N_27567);
xor U38417 (N_38417,N_26154,N_21826);
nor U38418 (N_38418,N_21455,N_20222);
or U38419 (N_38419,N_21628,N_26570);
or U38420 (N_38420,N_20717,N_29110);
nor U38421 (N_38421,N_20141,N_25648);
nand U38422 (N_38422,N_28130,N_20293);
and U38423 (N_38423,N_29468,N_29834);
or U38424 (N_38424,N_25692,N_29521);
and U38425 (N_38425,N_25696,N_22133);
and U38426 (N_38426,N_27745,N_20712);
and U38427 (N_38427,N_27599,N_23779);
xnor U38428 (N_38428,N_22717,N_20439);
xor U38429 (N_38429,N_27857,N_25425);
and U38430 (N_38430,N_21873,N_22804);
nor U38431 (N_38431,N_26646,N_26314);
xnor U38432 (N_38432,N_28158,N_29744);
nand U38433 (N_38433,N_20035,N_22947);
xnor U38434 (N_38434,N_29617,N_23069);
nor U38435 (N_38435,N_28094,N_21248);
or U38436 (N_38436,N_25594,N_25897);
nand U38437 (N_38437,N_24656,N_23027);
nor U38438 (N_38438,N_24987,N_27867);
xor U38439 (N_38439,N_22768,N_24830);
nor U38440 (N_38440,N_27209,N_22906);
nand U38441 (N_38441,N_20868,N_20297);
or U38442 (N_38442,N_26994,N_28698);
nor U38443 (N_38443,N_24973,N_27312);
nand U38444 (N_38444,N_26401,N_29588);
or U38445 (N_38445,N_28890,N_24481);
nand U38446 (N_38446,N_26959,N_22569);
nor U38447 (N_38447,N_20644,N_26256);
nand U38448 (N_38448,N_23212,N_26288);
or U38449 (N_38449,N_24828,N_23534);
and U38450 (N_38450,N_27592,N_25798);
and U38451 (N_38451,N_23282,N_20276);
nand U38452 (N_38452,N_27168,N_27078);
and U38453 (N_38453,N_20044,N_22303);
or U38454 (N_38454,N_20859,N_25198);
nand U38455 (N_38455,N_28709,N_20471);
nand U38456 (N_38456,N_27757,N_20026);
nor U38457 (N_38457,N_23251,N_25048);
xor U38458 (N_38458,N_29881,N_26156);
and U38459 (N_38459,N_26108,N_22959);
xnor U38460 (N_38460,N_24229,N_24937);
xnor U38461 (N_38461,N_29341,N_23818);
nor U38462 (N_38462,N_21976,N_22337);
and U38463 (N_38463,N_23995,N_28168);
nor U38464 (N_38464,N_23656,N_20135);
nor U38465 (N_38465,N_24013,N_29444);
and U38466 (N_38466,N_26557,N_23429);
and U38467 (N_38467,N_21264,N_22496);
or U38468 (N_38468,N_25028,N_20674);
or U38469 (N_38469,N_23197,N_24578);
nand U38470 (N_38470,N_26669,N_28134);
xnor U38471 (N_38471,N_23329,N_23591);
and U38472 (N_38472,N_26630,N_23029);
or U38473 (N_38473,N_26758,N_25343);
nand U38474 (N_38474,N_23549,N_21310);
or U38475 (N_38475,N_26497,N_24260);
nand U38476 (N_38476,N_26563,N_25120);
nand U38477 (N_38477,N_29668,N_22083);
nor U38478 (N_38478,N_23543,N_22385);
xor U38479 (N_38479,N_26117,N_29187);
and U38480 (N_38480,N_21445,N_27514);
nand U38481 (N_38481,N_25268,N_20472);
xor U38482 (N_38482,N_23388,N_27043);
nor U38483 (N_38483,N_21820,N_20791);
and U38484 (N_38484,N_21285,N_29619);
or U38485 (N_38485,N_28503,N_27134);
nand U38486 (N_38486,N_27215,N_24816);
nor U38487 (N_38487,N_28648,N_28852);
or U38488 (N_38488,N_24385,N_26488);
and U38489 (N_38489,N_20755,N_24082);
nand U38490 (N_38490,N_26608,N_20596);
and U38491 (N_38491,N_22849,N_27759);
nand U38492 (N_38492,N_22470,N_27968);
xor U38493 (N_38493,N_26290,N_22208);
nand U38494 (N_38494,N_28657,N_29900);
or U38495 (N_38495,N_23333,N_27107);
or U38496 (N_38496,N_21540,N_22816);
xnor U38497 (N_38497,N_20692,N_20874);
nor U38498 (N_38498,N_20706,N_24857);
nand U38499 (N_38499,N_20112,N_21294);
nor U38500 (N_38500,N_23450,N_28997);
xor U38501 (N_38501,N_25242,N_25787);
nand U38502 (N_38502,N_24180,N_25306);
or U38503 (N_38503,N_29542,N_27381);
and U38504 (N_38504,N_25462,N_28029);
and U38505 (N_38505,N_20457,N_25299);
and U38506 (N_38506,N_20267,N_29105);
and U38507 (N_38507,N_21474,N_29891);
or U38508 (N_38508,N_27022,N_25469);
or U38509 (N_38509,N_23510,N_26468);
or U38510 (N_38510,N_26158,N_23512);
or U38511 (N_38511,N_21098,N_26466);
and U38512 (N_38512,N_27387,N_26518);
and U38513 (N_38513,N_21917,N_22329);
nand U38514 (N_38514,N_28840,N_25334);
and U38515 (N_38515,N_23532,N_28975);
nor U38516 (N_38516,N_23504,N_20273);
nand U38517 (N_38517,N_24116,N_20639);
or U38518 (N_38518,N_21976,N_21706);
nand U38519 (N_38519,N_27511,N_20793);
and U38520 (N_38520,N_20578,N_26176);
xnor U38521 (N_38521,N_22618,N_25201);
xnor U38522 (N_38522,N_26118,N_24189);
nand U38523 (N_38523,N_26413,N_24749);
and U38524 (N_38524,N_28081,N_27690);
or U38525 (N_38525,N_23194,N_25815);
or U38526 (N_38526,N_26033,N_28780);
nand U38527 (N_38527,N_26660,N_23305);
xor U38528 (N_38528,N_20405,N_27735);
or U38529 (N_38529,N_24055,N_26134);
or U38530 (N_38530,N_20269,N_29545);
nand U38531 (N_38531,N_20856,N_24433);
and U38532 (N_38532,N_21217,N_25022);
and U38533 (N_38533,N_21278,N_25358);
or U38534 (N_38534,N_24300,N_20022);
and U38535 (N_38535,N_22103,N_27589);
or U38536 (N_38536,N_24394,N_20583);
nor U38537 (N_38537,N_27802,N_29365);
or U38538 (N_38538,N_22230,N_24201);
and U38539 (N_38539,N_24310,N_22315);
nor U38540 (N_38540,N_29257,N_24534);
xor U38541 (N_38541,N_27612,N_22892);
nor U38542 (N_38542,N_23825,N_27796);
nor U38543 (N_38543,N_25863,N_20325);
xnor U38544 (N_38544,N_27585,N_26816);
and U38545 (N_38545,N_24303,N_25002);
or U38546 (N_38546,N_24979,N_28703);
nand U38547 (N_38547,N_23832,N_23303);
or U38548 (N_38548,N_23403,N_28629);
or U38549 (N_38549,N_20855,N_27615);
xor U38550 (N_38550,N_25676,N_20920);
and U38551 (N_38551,N_20319,N_20713);
nand U38552 (N_38552,N_26300,N_26444);
nor U38553 (N_38553,N_23111,N_25376);
nor U38554 (N_38554,N_29005,N_27563);
nand U38555 (N_38555,N_25475,N_23566);
or U38556 (N_38556,N_23618,N_29312);
or U38557 (N_38557,N_23025,N_26828);
or U38558 (N_38558,N_24766,N_23413);
or U38559 (N_38559,N_21400,N_20371);
and U38560 (N_38560,N_23498,N_24979);
xor U38561 (N_38561,N_21856,N_25979);
nor U38562 (N_38562,N_22666,N_27200);
xnor U38563 (N_38563,N_24459,N_26427);
or U38564 (N_38564,N_21453,N_23524);
nand U38565 (N_38565,N_26250,N_21189);
nor U38566 (N_38566,N_20710,N_29736);
xor U38567 (N_38567,N_28532,N_22599);
nand U38568 (N_38568,N_29610,N_27901);
nor U38569 (N_38569,N_27655,N_28905);
xnor U38570 (N_38570,N_22724,N_24356);
xnor U38571 (N_38571,N_23173,N_23210);
and U38572 (N_38572,N_26789,N_22558);
nand U38573 (N_38573,N_26639,N_23556);
nand U38574 (N_38574,N_23977,N_23589);
or U38575 (N_38575,N_28083,N_23862);
nor U38576 (N_38576,N_28706,N_28421);
nand U38577 (N_38577,N_21106,N_27233);
xor U38578 (N_38578,N_23867,N_20573);
and U38579 (N_38579,N_22309,N_23166);
nand U38580 (N_38580,N_24666,N_29076);
nor U38581 (N_38581,N_23887,N_23001);
or U38582 (N_38582,N_26936,N_29230);
and U38583 (N_38583,N_24601,N_27541);
nor U38584 (N_38584,N_25769,N_27042);
xor U38585 (N_38585,N_21224,N_26568);
xnor U38586 (N_38586,N_29277,N_22361);
nand U38587 (N_38587,N_27618,N_22484);
or U38588 (N_38588,N_23336,N_25569);
nor U38589 (N_38589,N_23916,N_26277);
nand U38590 (N_38590,N_29162,N_21861);
or U38591 (N_38591,N_29150,N_28609);
and U38592 (N_38592,N_20637,N_24074);
nor U38593 (N_38593,N_20829,N_28546);
nor U38594 (N_38594,N_24060,N_23303);
and U38595 (N_38595,N_27586,N_21875);
or U38596 (N_38596,N_20751,N_25048);
nand U38597 (N_38597,N_27039,N_23221);
xnor U38598 (N_38598,N_24854,N_24949);
xnor U38599 (N_38599,N_28052,N_28600);
nand U38600 (N_38600,N_25134,N_26227);
and U38601 (N_38601,N_23099,N_22417);
nand U38602 (N_38602,N_24957,N_28120);
xor U38603 (N_38603,N_22108,N_27818);
nor U38604 (N_38604,N_26146,N_28646);
xor U38605 (N_38605,N_21141,N_26109);
nand U38606 (N_38606,N_29162,N_20308);
nor U38607 (N_38607,N_20230,N_22034);
nand U38608 (N_38608,N_27218,N_22081);
or U38609 (N_38609,N_29794,N_21731);
nand U38610 (N_38610,N_26374,N_27486);
xor U38611 (N_38611,N_25062,N_25508);
xor U38612 (N_38612,N_29907,N_21452);
and U38613 (N_38613,N_23097,N_20169);
and U38614 (N_38614,N_22198,N_27072);
nand U38615 (N_38615,N_20327,N_25493);
or U38616 (N_38616,N_26472,N_29291);
nand U38617 (N_38617,N_26393,N_21266);
nand U38618 (N_38618,N_22090,N_26654);
nor U38619 (N_38619,N_26382,N_25069);
nand U38620 (N_38620,N_23114,N_23950);
nand U38621 (N_38621,N_24200,N_21187);
xnor U38622 (N_38622,N_21434,N_24204);
or U38623 (N_38623,N_24500,N_24710);
and U38624 (N_38624,N_25201,N_29882);
nand U38625 (N_38625,N_28335,N_21740);
nand U38626 (N_38626,N_26787,N_26869);
and U38627 (N_38627,N_24053,N_24251);
xnor U38628 (N_38628,N_26269,N_29330);
xnor U38629 (N_38629,N_29346,N_21999);
or U38630 (N_38630,N_26091,N_29706);
nor U38631 (N_38631,N_23521,N_24537);
and U38632 (N_38632,N_22808,N_22793);
nor U38633 (N_38633,N_28280,N_23155);
xor U38634 (N_38634,N_20971,N_26378);
and U38635 (N_38635,N_22145,N_23538);
nand U38636 (N_38636,N_25461,N_27053);
and U38637 (N_38637,N_26899,N_22893);
xnor U38638 (N_38638,N_29299,N_28927);
and U38639 (N_38639,N_25404,N_21004);
or U38640 (N_38640,N_22029,N_24688);
xnor U38641 (N_38641,N_24216,N_26701);
xnor U38642 (N_38642,N_26014,N_24542);
or U38643 (N_38643,N_26753,N_23624);
nor U38644 (N_38644,N_20655,N_20737);
xor U38645 (N_38645,N_29112,N_26159);
nand U38646 (N_38646,N_25093,N_27826);
nor U38647 (N_38647,N_24980,N_21508);
or U38648 (N_38648,N_24843,N_20985);
nand U38649 (N_38649,N_26048,N_23526);
and U38650 (N_38650,N_25145,N_25686);
or U38651 (N_38651,N_27714,N_26238);
nor U38652 (N_38652,N_22762,N_21629);
nand U38653 (N_38653,N_24218,N_28513);
nor U38654 (N_38654,N_26631,N_20330);
nand U38655 (N_38655,N_24164,N_25378);
nand U38656 (N_38656,N_25526,N_21446);
nor U38657 (N_38657,N_22731,N_23599);
xnor U38658 (N_38658,N_24713,N_24413);
and U38659 (N_38659,N_23486,N_28393);
nand U38660 (N_38660,N_20817,N_24256);
nor U38661 (N_38661,N_20649,N_22550);
or U38662 (N_38662,N_29584,N_20862);
xnor U38663 (N_38663,N_20115,N_23812);
nand U38664 (N_38664,N_28658,N_23130);
xnor U38665 (N_38665,N_28587,N_23448);
and U38666 (N_38666,N_25898,N_28882);
or U38667 (N_38667,N_25768,N_22834);
or U38668 (N_38668,N_20893,N_24880);
or U38669 (N_38669,N_21872,N_24791);
nor U38670 (N_38670,N_27945,N_24771);
xnor U38671 (N_38671,N_25196,N_23835);
and U38672 (N_38672,N_22869,N_22710);
xor U38673 (N_38673,N_24563,N_27478);
nor U38674 (N_38674,N_27811,N_29483);
xnor U38675 (N_38675,N_29330,N_28304);
or U38676 (N_38676,N_28579,N_23319);
or U38677 (N_38677,N_29801,N_29896);
xnor U38678 (N_38678,N_22744,N_29383);
nand U38679 (N_38679,N_28584,N_29698);
or U38680 (N_38680,N_28151,N_28946);
or U38681 (N_38681,N_28765,N_24774);
and U38682 (N_38682,N_27782,N_22758);
or U38683 (N_38683,N_26665,N_28296);
nand U38684 (N_38684,N_28908,N_22784);
and U38685 (N_38685,N_28712,N_20429);
nor U38686 (N_38686,N_23436,N_29060);
nor U38687 (N_38687,N_22065,N_29198);
xor U38688 (N_38688,N_27230,N_29468);
or U38689 (N_38689,N_27880,N_23111);
nor U38690 (N_38690,N_28299,N_26322);
xor U38691 (N_38691,N_29505,N_20847);
xor U38692 (N_38692,N_28680,N_21296);
nor U38693 (N_38693,N_24549,N_24408);
nor U38694 (N_38694,N_23940,N_26428);
xor U38695 (N_38695,N_22178,N_27148);
nand U38696 (N_38696,N_29445,N_23786);
nand U38697 (N_38697,N_29475,N_26653);
xnor U38698 (N_38698,N_26639,N_29687);
nand U38699 (N_38699,N_23262,N_27500);
nand U38700 (N_38700,N_22479,N_24236);
xor U38701 (N_38701,N_20188,N_24607);
xnor U38702 (N_38702,N_29823,N_21250);
or U38703 (N_38703,N_28111,N_21427);
or U38704 (N_38704,N_27029,N_23966);
xor U38705 (N_38705,N_26890,N_23917);
nand U38706 (N_38706,N_24284,N_27932);
nand U38707 (N_38707,N_28259,N_29005);
and U38708 (N_38708,N_29535,N_26431);
nand U38709 (N_38709,N_24360,N_29728);
or U38710 (N_38710,N_25394,N_21714);
nand U38711 (N_38711,N_27529,N_24221);
and U38712 (N_38712,N_29710,N_27473);
xnor U38713 (N_38713,N_26646,N_28686);
nor U38714 (N_38714,N_20278,N_21455);
or U38715 (N_38715,N_26074,N_23771);
or U38716 (N_38716,N_21175,N_25496);
or U38717 (N_38717,N_29247,N_23342);
or U38718 (N_38718,N_29106,N_21249);
nor U38719 (N_38719,N_20739,N_27347);
xnor U38720 (N_38720,N_25082,N_25467);
nor U38721 (N_38721,N_20955,N_29810);
xnor U38722 (N_38722,N_24127,N_27090);
xor U38723 (N_38723,N_27251,N_22274);
nand U38724 (N_38724,N_25100,N_26169);
and U38725 (N_38725,N_23328,N_25634);
or U38726 (N_38726,N_24668,N_21040);
nor U38727 (N_38727,N_27862,N_22674);
nor U38728 (N_38728,N_23836,N_26063);
nand U38729 (N_38729,N_28508,N_20095);
nand U38730 (N_38730,N_25007,N_27268);
nand U38731 (N_38731,N_29689,N_28342);
or U38732 (N_38732,N_24492,N_20316);
xnor U38733 (N_38733,N_25510,N_21695);
and U38734 (N_38734,N_20164,N_29278);
or U38735 (N_38735,N_23262,N_22743);
or U38736 (N_38736,N_22134,N_24413);
or U38737 (N_38737,N_28359,N_26776);
xor U38738 (N_38738,N_24167,N_22553);
or U38739 (N_38739,N_26817,N_24941);
and U38740 (N_38740,N_29014,N_25023);
or U38741 (N_38741,N_23070,N_22420);
or U38742 (N_38742,N_23502,N_22199);
nor U38743 (N_38743,N_28448,N_27859);
nand U38744 (N_38744,N_20554,N_20918);
or U38745 (N_38745,N_25394,N_24624);
nor U38746 (N_38746,N_29389,N_24467);
and U38747 (N_38747,N_28079,N_28945);
or U38748 (N_38748,N_22041,N_24707);
nand U38749 (N_38749,N_29920,N_27352);
nor U38750 (N_38750,N_24790,N_21867);
nand U38751 (N_38751,N_21214,N_27042);
and U38752 (N_38752,N_22366,N_23663);
or U38753 (N_38753,N_26611,N_28263);
nand U38754 (N_38754,N_28670,N_28364);
or U38755 (N_38755,N_28956,N_22404);
and U38756 (N_38756,N_29598,N_25340);
and U38757 (N_38757,N_24937,N_21044);
xor U38758 (N_38758,N_20206,N_26531);
nor U38759 (N_38759,N_29575,N_23143);
xor U38760 (N_38760,N_26152,N_27208);
xor U38761 (N_38761,N_20652,N_29342);
or U38762 (N_38762,N_25251,N_26202);
nand U38763 (N_38763,N_27322,N_20376);
nor U38764 (N_38764,N_22851,N_27359);
or U38765 (N_38765,N_29222,N_20745);
nand U38766 (N_38766,N_20346,N_20816);
nand U38767 (N_38767,N_21225,N_26479);
xnor U38768 (N_38768,N_29724,N_25523);
xnor U38769 (N_38769,N_27160,N_22521);
xor U38770 (N_38770,N_24989,N_26187);
or U38771 (N_38771,N_22760,N_21460);
nand U38772 (N_38772,N_20030,N_21949);
and U38773 (N_38773,N_21702,N_20871);
or U38774 (N_38774,N_28975,N_23723);
nor U38775 (N_38775,N_26319,N_28475);
and U38776 (N_38776,N_24948,N_27520);
and U38777 (N_38777,N_28920,N_25639);
and U38778 (N_38778,N_23293,N_22826);
and U38779 (N_38779,N_22020,N_21896);
nand U38780 (N_38780,N_29366,N_28876);
nand U38781 (N_38781,N_22537,N_29706);
nand U38782 (N_38782,N_24653,N_21117);
and U38783 (N_38783,N_26120,N_20393);
or U38784 (N_38784,N_24858,N_23481);
xor U38785 (N_38785,N_26953,N_25818);
nand U38786 (N_38786,N_23818,N_23103);
and U38787 (N_38787,N_21108,N_23390);
nor U38788 (N_38788,N_23546,N_21916);
or U38789 (N_38789,N_25870,N_24568);
nand U38790 (N_38790,N_27353,N_24330);
nor U38791 (N_38791,N_26620,N_24453);
and U38792 (N_38792,N_28245,N_20434);
and U38793 (N_38793,N_22589,N_24824);
nand U38794 (N_38794,N_21958,N_28005);
and U38795 (N_38795,N_29326,N_25199);
nor U38796 (N_38796,N_20920,N_22746);
nor U38797 (N_38797,N_22787,N_27052);
and U38798 (N_38798,N_25971,N_27414);
xnor U38799 (N_38799,N_24172,N_27402);
and U38800 (N_38800,N_26388,N_28545);
xnor U38801 (N_38801,N_23066,N_22022);
xnor U38802 (N_38802,N_22764,N_28953);
nand U38803 (N_38803,N_23163,N_28307);
nand U38804 (N_38804,N_28750,N_22508);
nand U38805 (N_38805,N_27019,N_28532);
nand U38806 (N_38806,N_26339,N_29493);
nand U38807 (N_38807,N_23396,N_23292);
nand U38808 (N_38808,N_20857,N_25113);
xnor U38809 (N_38809,N_28728,N_22723);
or U38810 (N_38810,N_21239,N_29180);
nand U38811 (N_38811,N_27856,N_28180);
nor U38812 (N_38812,N_22915,N_20676);
nand U38813 (N_38813,N_25473,N_29022);
and U38814 (N_38814,N_23377,N_22532);
nand U38815 (N_38815,N_24268,N_23598);
nor U38816 (N_38816,N_23776,N_25029);
and U38817 (N_38817,N_21391,N_23881);
and U38818 (N_38818,N_25243,N_28565);
nor U38819 (N_38819,N_20442,N_28713);
nand U38820 (N_38820,N_22650,N_20277);
xnor U38821 (N_38821,N_28538,N_25086);
or U38822 (N_38822,N_26612,N_23728);
xnor U38823 (N_38823,N_25758,N_20901);
and U38824 (N_38824,N_22720,N_25477);
nor U38825 (N_38825,N_20200,N_20123);
xnor U38826 (N_38826,N_26313,N_26287);
and U38827 (N_38827,N_25884,N_28003);
xor U38828 (N_38828,N_26615,N_24018);
xnor U38829 (N_38829,N_28706,N_24338);
xor U38830 (N_38830,N_26049,N_29668);
or U38831 (N_38831,N_24043,N_27735);
or U38832 (N_38832,N_21870,N_22580);
and U38833 (N_38833,N_29894,N_23572);
xnor U38834 (N_38834,N_21550,N_24300);
or U38835 (N_38835,N_28619,N_26216);
xor U38836 (N_38836,N_29217,N_26120);
and U38837 (N_38837,N_21710,N_29469);
and U38838 (N_38838,N_24303,N_27601);
nor U38839 (N_38839,N_26097,N_26065);
nand U38840 (N_38840,N_25926,N_29849);
and U38841 (N_38841,N_20404,N_29145);
and U38842 (N_38842,N_26787,N_20500);
or U38843 (N_38843,N_28674,N_22042);
nand U38844 (N_38844,N_26678,N_20378);
xnor U38845 (N_38845,N_23601,N_26512);
and U38846 (N_38846,N_24644,N_27866);
nor U38847 (N_38847,N_27665,N_20135);
nand U38848 (N_38848,N_21330,N_21282);
nor U38849 (N_38849,N_27755,N_24229);
xnor U38850 (N_38850,N_29188,N_24830);
and U38851 (N_38851,N_28687,N_25766);
and U38852 (N_38852,N_21062,N_26697);
or U38853 (N_38853,N_25159,N_27798);
xnor U38854 (N_38854,N_28963,N_23513);
nor U38855 (N_38855,N_26645,N_24566);
and U38856 (N_38856,N_23186,N_20641);
and U38857 (N_38857,N_23424,N_23028);
nand U38858 (N_38858,N_24484,N_23151);
or U38859 (N_38859,N_22808,N_22691);
and U38860 (N_38860,N_27509,N_26486);
xor U38861 (N_38861,N_27993,N_28213);
xor U38862 (N_38862,N_29303,N_25869);
or U38863 (N_38863,N_29509,N_23171);
or U38864 (N_38864,N_21842,N_28134);
or U38865 (N_38865,N_27745,N_23518);
or U38866 (N_38866,N_26493,N_29518);
nand U38867 (N_38867,N_22393,N_26151);
or U38868 (N_38868,N_28104,N_26322);
nor U38869 (N_38869,N_25411,N_22668);
xnor U38870 (N_38870,N_24640,N_23457);
or U38871 (N_38871,N_29957,N_20153);
or U38872 (N_38872,N_25247,N_21599);
xor U38873 (N_38873,N_27539,N_29731);
nor U38874 (N_38874,N_24794,N_27372);
or U38875 (N_38875,N_20987,N_23284);
or U38876 (N_38876,N_23388,N_21078);
nand U38877 (N_38877,N_21160,N_21372);
nor U38878 (N_38878,N_26020,N_27370);
or U38879 (N_38879,N_23909,N_25918);
or U38880 (N_38880,N_24260,N_23543);
or U38881 (N_38881,N_25200,N_20758);
xor U38882 (N_38882,N_24738,N_28569);
xor U38883 (N_38883,N_28835,N_24772);
xor U38884 (N_38884,N_22185,N_23339);
and U38885 (N_38885,N_22804,N_21064);
nor U38886 (N_38886,N_23574,N_28126);
xnor U38887 (N_38887,N_27292,N_22210);
or U38888 (N_38888,N_23938,N_25460);
nor U38889 (N_38889,N_25400,N_29408);
nand U38890 (N_38890,N_22013,N_26634);
xor U38891 (N_38891,N_26247,N_23720);
or U38892 (N_38892,N_28524,N_26963);
or U38893 (N_38893,N_27862,N_25325);
or U38894 (N_38894,N_27683,N_28580);
nand U38895 (N_38895,N_22871,N_21484);
or U38896 (N_38896,N_23682,N_25561);
nor U38897 (N_38897,N_27272,N_23197);
nand U38898 (N_38898,N_27852,N_20090);
or U38899 (N_38899,N_27785,N_22578);
or U38900 (N_38900,N_29913,N_22787);
or U38901 (N_38901,N_22542,N_21141);
xor U38902 (N_38902,N_24149,N_24958);
or U38903 (N_38903,N_24984,N_21914);
nor U38904 (N_38904,N_24070,N_23884);
xnor U38905 (N_38905,N_29457,N_26920);
xor U38906 (N_38906,N_20957,N_26049);
and U38907 (N_38907,N_25772,N_29497);
nor U38908 (N_38908,N_24486,N_23369);
xnor U38909 (N_38909,N_27162,N_23347);
nand U38910 (N_38910,N_26603,N_20834);
nor U38911 (N_38911,N_24144,N_28688);
nand U38912 (N_38912,N_23450,N_20944);
or U38913 (N_38913,N_22638,N_25819);
and U38914 (N_38914,N_27665,N_20009);
and U38915 (N_38915,N_28508,N_23986);
or U38916 (N_38916,N_20043,N_22900);
and U38917 (N_38917,N_26845,N_25571);
and U38918 (N_38918,N_22118,N_21817);
xnor U38919 (N_38919,N_27383,N_22827);
xnor U38920 (N_38920,N_23658,N_25093);
nor U38921 (N_38921,N_28363,N_23932);
nor U38922 (N_38922,N_21587,N_24710);
or U38923 (N_38923,N_25407,N_21434);
or U38924 (N_38924,N_23049,N_25705);
or U38925 (N_38925,N_26335,N_26885);
xor U38926 (N_38926,N_21930,N_29741);
xnor U38927 (N_38927,N_26700,N_25651);
and U38928 (N_38928,N_21688,N_27065);
nor U38929 (N_38929,N_24991,N_21162);
xnor U38930 (N_38930,N_25679,N_22317);
xor U38931 (N_38931,N_27985,N_24632);
xnor U38932 (N_38932,N_21325,N_28662);
or U38933 (N_38933,N_28087,N_25350);
and U38934 (N_38934,N_28095,N_21725);
and U38935 (N_38935,N_27106,N_20681);
nand U38936 (N_38936,N_28293,N_21554);
xnor U38937 (N_38937,N_21538,N_26060);
nor U38938 (N_38938,N_28813,N_22558);
nor U38939 (N_38939,N_20178,N_22589);
xnor U38940 (N_38940,N_20413,N_23062);
and U38941 (N_38941,N_25180,N_22569);
or U38942 (N_38942,N_27424,N_24544);
and U38943 (N_38943,N_20509,N_25778);
or U38944 (N_38944,N_27947,N_24740);
nor U38945 (N_38945,N_27459,N_27500);
nor U38946 (N_38946,N_22567,N_27116);
nor U38947 (N_38947,N_25974,N_28086);
or U38948 (N_38948,N_22064,N_23459);
nand U38949 (N_38949,N_25939,N_27523);
nand U38950 (N_38950,N_25506,N_28255);
nor U38951 (N_38951,N_21003,N_22578);
nor U38952 (N_38952,N_22265,N_29758);
nor U38953 (N_38953,N_22116,N_27791);
xor U38954 (N_38954,N_23800,N_27974);
or U38955 (N_38955,N_24486,N_24214);
nor U38956 (N_38956,N_24867,N_26175);
nand U38957 (N_38957,N_22971,N_24858);
and U38958 (N_38958,N_20575,N_28536);
and U38959 (N_38959,N_27516,N_22187);
or U38960 (N_38960,N_23426,N_29543);
nand U38961 (N_38961,N_28270,N_28070);
or U38962 (N_38962,N_25862,N_23813);
xor U38963 (N_38963,N_26568,N_22525);
xnor U38964 (N_38964,N_27399,N_21496);
nand U38965 (N_38965,N_27523,N_23584);
xnor U38966 (N_38966,N_23761,N_25307);
or U38967 (N_38967,N_24246,N_24641);
and U38968 (N_38968,N_20931,N_29520);
or U38969 (N_38969,N_27598,N_28527);
nor U38970 (N_38970,N_25528,N_20879);
xnor U38971 (N_38971,N_25012,N_24096);
xnor U38972 (N_38972,N_29141,N_24929);
nor U38973 (N_38973,N_26844,N_29941);
xnor U38974 (N_38974,N_27988,N_28899);
nand U38975 (N_38975,N_29307,N_20087);
or U38976 (N_38976,N_23644,N_21837);
and U38977 (N_38977,N_29495,N_21054);
or U38978 (N_38978,N_23979,N_25351);
or U38979 (N_38979,N_22027,N_28319);
nor U38980 (N_38980,N_25258,N_28190);
xor U38981 (N_38981,N_26917,N_20260);
or U38982 (N_38982,N_28597,N_29878);
nor U38983 (N_38983,N_24243,N_20951);
or U38984 (N_38984,N_23093,N_27023);
or U38985 (N_38985,N_28126,N_23221);
or U38986 (N_38986,N_25676,N_25037);
nor U38987 (N_38987,N_29889,N_22018);
nor U38988 (N_38988,N_27539,N_25452);
nor U38989 (N_38989,N_27377,N_25781);
and U38990 (N_38990,N_29308,N_20874);
and U38991 (N_38991,N_21425,N_20628);
or U38992 (N_38992,N_26020,N_24376);
xnor U38993 (N_38993,N_21551,N_24609);
and U38994 (N_38994,N_21943,N_28458);
nand U38995 (N_38995,N_25156,N_24169);
nor U38996 (N_38996,N_20890,N_23704);
nor U38997 (N_38997,N_25357,N_21361);
or U38998 (N_38998,N_20167,N_24800);
or U38999 (N_38999,N_22436,N_21455);
nor U39000 (N_39000,N_20328,N_29240);
xnor U39001 (N_39001,N_26682,N_26153);
xor U39002 (N_39002,N_22169,N_27024);
or U39003 (N_39003,N_29976,N_21830);
nor U39004 (N_39004,N_26711,N_26121);
or U39005 (N_39005,N_22772,N_22029);
nand U39006 (N_39006,N_24074,N_22761);
or U39007 (N_39007,N_26572,N_21111);
or U39008 (N_39008,N_24721,N_22416);
nor U39009 (N_39009,N_22035,N_26659);
and U39010 (N_39010,N_21750,N_26202);
nand U39011 (N_39011,N_22492,N_21843);
nor U39012 (N_39012,N_23097,N_23264);
and U39013 (N_39013,N_24032,N_20723);
nand U39014 (N_39014,N_29024,N_22103);
xnor U39015 (N_39015,N_27565,N_27591);
nor U39016 (N_39016,N_22073,N_26036);
or U39017 (N_39017,N_28264,N_29185);
nor U39018 (N_39018,N_22779,N_22742);
nor U39019 (N_39019,N_26365,N_23380);
nor U39020 (N_39020,N_25607,N_28202);
and U39021 (N_39021,N_26253,N_23555);
nor U39022 (N_39022,N_23862,N_24388);
nand U39023 (N_39023,N_24644,N_22037);
xor U39024 (N_39024,N_25424,N_25931);
and U39025 (N_39025,N_22152,N_27633);
nor U39026 (N_39026,N_23418,N_23805);
nor U39027 (N_39027,N_21959,N_22024);
nand U39028 (N_39028,N_23196,N_25338);
nand U39029 (N_39029,N_26949,N_24541);
xor U39030 (N_39030,N_29087,N_25190);
and U39031 (N_39031,N_25719,N_25091);
or U39032 (N_39032,N_21006,N_28468);
and U39033 (N_39033,N_29450,N_22506);
nand U39034 (N_39034,N_28569,N_28253);
and U39035 (N_39035,N_26812,N_28453);
nor U39036 (N_39036,N_29914,N_27207);
nor U39037 (N_39037,N_23043,N_29815);
xor U39038 (N_39038,N_24036,N_24178);
and U39039 (N_39039,N_24921,N_25712);
nand U39040 (N_39040,N_27444,N_28992);
xor U39041 (N_39041,N_21440,N_28345);
or U39042 (N_39042,N_28410,N_26791);
and U39043 (N_39043,N_20612,N_22272);
and U39044 (N_39044,N_28664,N_29468);
nor U39045 (N_39045,N_20405,N_27889);
nand U39046 (N_39046,N_22657,N_25233);
or U39047 (N_39047,N_24700,N_24355);
xnor U39048 (N_39048,N_23169,N_22163);
xor U39049 (N_39049,N_29025,N_22678);
nand U39050 (N_39050,N_28351,N_23093);
or U39051 (N_39051,N_24725,N_28500);
xnor U39052 (N_39052,N_28973,N_26113);
and U39053 (N_39053,N_20649,N_26028);
xor U39054 (N_39054,N_25191,N_22080);
or U39055 (N_39055,N_26234,N_21033);
nor U39056 (N_39056,N_22092,N_29633);
xor U39057 (N_39057,N_28153,N_22867);
and U39058 (N_39058,N_20285,N_22632);
nand U39059 (N_39059,N_25314,N_23705);
and U39060 (N_39060,N_23431,N_26430);
nand U39061 (N_39061,N_21810,N_25777);
nand U39062 (N_39062,N_21783,N_26574);
and U39063 (N_39063,N_21412,N_20151);
and U39064 (N_39064,N_24278,N_28535);
nand U39065 (N_39065,N_25325,N_22435);
nor U39066 (N_39066,N_25800,N_28107);
nor U39067 (N_39067,N_24990,N_25061);
nor U39068 (N_39068,N_26110,N_24863);
nand U39069 (N_39069,N_21777,N_23724);
or U39070 (N_39070,N_25014,N_23274);
or U39071 (N_39071,N_24866,N_24705);
or U39072 (N_39072,N_24401,N_24709);
xor U39073 (N_39073,N_27411,N_21577);
nor U39074 (N_39074,N_21631,N_20674);
and U39075 (N_39075,N_28770,N_26850);
nor U39076 (N_39076,N_24772,N_23769);
nand U39077 (N_39077,N_27903,N_20245);
nor U39078 (N_39078,N_21741,N_27236);
or U39079 (N_39079,N_25147,N_20734);
nand U39080 (N_39080,N_26873,N_29283);
or U39081 (N_39081,N_28657,N_25761);
nand U39082 (N_39082,N_21342,N_23011);
xor U39083 (N_39083,N_26230,N_29941);
xor U39084 (N_39084,N_24559,N_21585);
xnor U39085 (N_39085,N_27397,N_22583);
or U39086 (N_39086,N_20162,N_25538);
nor U39087 (N_39087,N_26904,N_27532);
nor U39088 (N_39088,N_22217,N_21342);
nor U39089 (N_39089,N_26302,N_23754);
and U39090 (N_39090,N_20247,N_28877);
xnor U39091 (N_39091,N_20787,N_28173);
nor U39092 (N_39092,N_21584,N_21500);
xor U39093 (N_39093,N_24772,N_23135);
nand U39094 (N_39094,N_29389,N_22796);
nor U39095 (N_39095,N_24914,N_29957);
nand U39096 (N_39096,N_29746,N_22235);
xor U39097 (N_39097,N_23699,N_20390);
xor U39098 (N_39098,N_24616,N_25510);
nor U39099 (N_39099,N_26115,N_21277);
nor U39100 (N_39100,N_20527,N_28731);
nor U39101 (N_39101,N_26655,N_22915);
nand U39102 (N_39102,N_22664,N_24057);
xor U39103 (N_39103,N_28503,N_24636);
and U39104 (N_39104,N_28441,N_24771);
xor U39105 (N_39105,N_20792,N_27035);
and U39106 (N_39106,N_27249,N_29158);
or U39107 (N_39107,N_23629,N_28234);
nand U39108 (N_39108,N_21996,N_21982);
nor U39109 (N_39109,N_26802,N_23281);
nor U39110 (N_39110,N_22407,N_27395);
nand U39111 (N_39111,N_20345,N_22202);
nand U39112 (N_39112,N_25072,N_28407);
and U39113 (N_39113,N_24030,N_20513);
nand U39114 (N_39114,N_27046,N_27794);
or U39115 (N_39115,N_28172,N_24660);
nand U39116 (N_39116,N_20067,N_26998);
and U39117 (N_39117,N_26480,N_24173);
and U39118 (N_39118,N_20499,N_26647);
or U39119 (N_39119,N_22728,N_28532);
and U39120 (N_39120,N_21576,N_29811);
nand U39121 (N_39121,N_23446,N_29863);
and U39122 (N_39122,N_26098,N_27462);
or U39123 (N_39123,N_25274,N_22467);
nor U39124 (N_39124,N_29962,N_25357);
or U39125 (N_39125,N_20601,N_20519);
or U39126 (N_39126,N_24763,N_22550);
or U39127 (N_39127,N_20341,N_22127);
nor U39128 (N_39128,N_25902,N_27022);
nand U39129 (N_39129,N_29793,N_26521);
or U39130 (N_39130,N_21433,N_21395);
or U39131 (N_39131,N_21328,N_26618);
or U39132 (N_39132,N_29127,N_26317);
or U39133 (N_39133,N_22967,N_23190);
and U39134 (N_39134,N_21154,N_24912);
xnor U39135 (N_39135,N_29854,N_28121);
xnor U39136 (N_39136,N_22379,N_27154);
nand U39137 (N_39137,N_22449,N_20967);
xnor U39138 (N_39138,N_20665,N_25131);
nor U39139 (N_39139,N_27405,N_21183);
nor U39140 (N_39140,N_29239,N_25960);
and U39141 (N_39141,N_21850,N_27193);
and U39142 (N_39142,N_26669,N_27558);
nor U39143 (N_39143,N_26200,N_22269);
and U39144 (N_39144,N_22850,N_29307);
and U39145 (N_39145,N_20391,N_26097);
nor U39146 (N_39146,N_27356,N_23059);
xor U39147 (N_39147,N_27196,N_26421);
nor U39148 (N_39148,N_26431,N_28035);
nand U39149 (N_39149,N_26644,N_21996);
nand U39150 (N_39150,N_20180,N_24883);
nand U39151 (N_39151,N_28590,N_20968);
nand U39152 (N_39152,N_29766,N_21210);
nor U39153 (N_39153,N_27648,N_21015);
and U39154 (N_39154,N_21996,N_22274);
nand U39155 (N_39155,N_28525,N_20675);
nor U39156 (N_39156,N_26944,N_27112);
or U39157 (N_39157,N_27066,N_29550);
and U39158 (N_39158,N_21875,N_29901);
xnor U39159 (N_39159,N_22372,N_23571);
or U39160 (N_39160,N_23103,N_20683);
nand U39161 (N_39161,N_27814,N_22876);
nor U39162 (N_39162,N_21772,N_20259);
and U39163 (N_39163,N_27597,N_22947);
nor U39164 (N_39164,N_29970,N_20073);
nor U39165 (N_39165,N_27051,N_21571);
nor U39166 (N_39166,N_20949,N_22808);
nor U39167 (N_39167,N_29496,N_26019);
xnor U39168 (N_39168,N_20888,N_24155);
or U39169 (N_39169,N_27201,N_20826);
or U39170 (N_39170,N_21399,N_26573);
xor U39171 (N_39171,N_23692,N_26618);
xnor U39172 (N_39172,N_20124,N_26852);
or U39173 (N_39173,N_29256,N_26682);
nand U39174 (N_39174,N_25386,N_24555);
xor U39175 (N_39175,N_23375,N_22027);
nand U39176 (N_39176,N_28338,N_25284);
or U39177 (N_39177,N_24378,N_29426);
nand U39178 (N_39178,N_26890,N_25509);
and U39179 (N_39179,N_24541,N_28901);
nand U39180 (N_39180,N_20608,N_27526);
nor U39181 (N_39181,N_28401,N_25559);
or U39182 (N_39182,N_29919,N_21286);
xnor U39183 (N_39183,N_26558,N_27261);
nor U39184 (N_39184,N_26224,N_25975);
nor U39185 (N_39185,N_28576,N_23197);
and U39186 (N_39186,N_23643,N_20197);
nor U39187 (N_39187,N_22207,N_20085);
xor U39188 (N_39188,N_22037,N_28485);
xnor U39189 (N_39189,N_21880,N_27587);
xor U39190 (N_39190,N_24170,N_24072);
nor U39191 (N_39191,N_28292,N_26173);
or U39192 (N_39192,N_25420,N_26162);
or U39193 (N_39193,N_28555,N_21010);
nor U39194 (N_39194,N_28106,N_24929);
or U39195 (N_39195,N_21744,N_20914);
nand U39196 (N_39196,N_28674,N_26793);
nor U39197 (N_39197,N_28134,N_20017);
or U39198 (N_39198,N_21382,N_21675);
nand U39199 (N_39199,N_27114,N_20891);
nand U39200 (N_39200,N_22736,N_25031);
or U39201 (N_39201,N_29049,N_27031);
and U39202 (N_39202,N_28183,N_29378);
xnor U39203 (N_39203,N_26232,N_27645);
and U39204 (N_39204,N_26350,N_26057);
nand U39205 (N_39205,N_29131,N_29151);
xor U39206 (N_39206,N_24218,N_28327);
or U39207 (N_39207,N_26533,N_29695);
or U39208 (N_39208,N_20957,N_25412);
nor U39209 (N_39209,N_28102,N_22802);
nor U39210 (N_39210,N_23684,N_29453);
nand U39211 (N_39211,N_21067,N_20295);
nor U39212 (N_39212,N_23239,N_22055);
xnor U39213 (N_39213,N_20883,N_23983);
or U39214 (N_39214,N_24746,N_24120);
xor U39215 (N_39215,N_23995,N_26771);
and U39216 (N_39216,N_23398,N_24025);
nand U39217 (N_39217,N_21925,N_25462);
or U39218 (N_39218,N_21667,N_28495);
nor U39219 (N_39219,N_28986,N_29874);
nor U39220 (N_39220,N_21435,N_27803);
nor U39221 (N_39221,N_28719,N_23935);
xor U39222 (N_39222,N_29183,N_21885);
nor U39223 (N_39223,N_23869,N_24946);
nor U39224 (N_39224,N_27003,N_29004);
nand U39225 (N_39225,N_28496,N_23830);
nand U39226 (N_39226,N_26971,N_27156);
and U39227 (N_39227,N_25119,N_24978);
xnor U39228 (N_39228,N_28035,N_21102);
nor U39229 (N_39229,N_28783,N_26121);
and U39230 (N_39230,N_27763,N_28969);
and U39231 (N_39231,N_26594,N_21577);
nand U39232 (N_39232,N_22514,N_24466);
or U39233 (N_39233,N_28503,N_21463);
and U39234 (N_39234,N_28986,N_24453);
xor U39235 (N_39235,N_24685,N_23117);
nor U39236 (N_39236,N_26095,N_28722);
xnor U39237 (N_39237,N_20207,N_26110);
nand U39238 (N_39238,N_29231,N_29658);
nor U39239 (N_39239,N_20978,N_28906);
nand U39240 (N_39240,N_21838,N_25071);
xor U39241 (N_39241,N_23127,N_23052);
nor U39242 (N_39242,N_23269,N_22376);
xor U39243 (N_39243,N_20094,N_23912);
and U39244 (N_39244,N_29814,N_27960);
nand U39245 (N_39245,N_29832,N_20425);
nor U39246 (N_39246,N_26166,N_20301);
xor U39247 (N_39247,N_25388,N_23595);
nor U39248 (N_39248,N_25690,N_20288);
xnor U39249 (N_39249,N_26226,N_23878);
and U39250 (N_39250,N_24020,N_28872);
nor U39251 (N_39251,N_20972,N_21766);
or U39252 (N_39252,N_27481,N_22392);
and U39253 (N_39253,N_23256,N_25866);
nand U39254 (N_39254,N_21617,N_22835);
xnor U39255 (N_39255,N_24933,N_24716);
and U39256 (N_39256,N_23376,N_22823);
xor U39257 (N_39257,N_25093,N_28587);
or U39258 (N_39258,N_27410,N_23703);
nor U39259 (N_39259,N_20565,N_26240);
xnor U39260 (N_39260,N_21256,N_26113);
nand U39261 (N_39261,N_24473,N_23655);
xor U39262 (N_39262,N_23748,N_29739);
or U39263 (N_39263,N_20766,N_27599);
and U39264 (N_39264,N_22676,N_29629);
nand U39265 (N_39265,N_24142,N_29149);
nand U39266 (N_39266,N_25742,N_29417);
nor U39267 (N_39267,N_28066,N_22529);
nand U39268 (N_39268,N_26461,N_29608);
and U39269 (N_39269,N_23798,N_20738);
xnor U39270 (N_39270,N_25557,N_27662);
nand U39271 (N_39271,N_27026,N_23306);
or U39272 (N_39272,N_22271,N_24286);
nand U39273 (N_39273,N_24367,N_27549);
and U39274 (N_39274,N_27814,N_27131);
xnor U39275 (N_39275,N_27684,N_25802);
nor U39276 (N_39276,N_27935,N_23169);
and U39277 (N_39277,N_24340,N_29963);
xor U39278 (N_39278,N_21830,N_26163);
nor U39279 (N_39279,N_28727,N_22109);
and U39280 (N_39280,N_26700,N_28895);
nand U39281 (N_39281,N_22564,N_29528);
nand U39282 (N_39282,N_26485,N_22338);
nor U39283 (N_39283,N_25494,N_27889);
or U39284 (N_39284,N_25803,N_21838);
or U39285 (N_39285,N_20468,N_20141);
xor U39286 (N_39286,N_24123,N_21628);
xnor U39287 (N_39287,N_26978,N_26366);
nor U39288 (N_39288,N_22351,N_27762);
nor U39289 (N_39289,N_20074,N_20378);
or U39290 (N_39290,N_23349,N_21175);
and U39291 (N_39291,N_29802,N_20955);
xnor U39292 (N_39292,N_20156,N_28716);
and U39293 (N_39293,N_22678,N_24808);
nand U39294 (N_39294,N_26818,N_22473);
nand U39295 (N_39295,N_28108,N_29930);
and U39296 (N_39296,N_29013,N_25260);
nand U39297 (N_39297,N_24079,N_22822);
nand U39298 (N_39298,N_20990,N_28227);
or U39299 (N_39299,N_21229,N_29762);
nor U39300 (N_39300,N_23278,N_29838);
nand U39301 (N_39301,N_25072,N_29504);
nor U39302 (N_39302,N_28281,N_22611);
or U39303 (N_39303,N_20072,N_23978);
and U39304 (N_39304,N_26010,N_23827);
and U39305 (N_39305,N_24846,N_28394);
nand U39306 (N_39306,N_22618,N_25484);
and U39307 (N_39307,N_29236,N_28603);
and U39308 (N_39308,N_27450,N_20930);
and U39309 (N_39309,N_27786,N_27366);
nand U39310 (N_39310,N_28810,N_27150);
nand U39311 (N_39311,N_28641,N_24119);
xnor U39312 (N_39312,N_25674,N_25006);
or U39313 (N_39313,N_23731,N_27835);
nand U39314 (N_39314,N_25877,N_20774);
xnor U39315 (N_39315,N_25041,N_24678);
nand U39316 (N_39316,N_29035,N_25809);
xor U39317 (N_39317,N_22666,N_21930);
nand U39318 (N_39318,N_21171,N_28123);
and U39319 (N_39319,N_24356,N_27078);
and U39320 (N_39320,N_22906,N_26882);
and U39321 (N_39321,N_25363,N_21973);
or U39322 (N_39322,N_25661,N_29843);
or U39323 (N_39323,N_21435,N_28620);
nand U39324 (N_39324,N_29533,N_20441);
nand U39325 (N_39325,N_28096,N_28171);
nor U39326 (N_39326,N_24674,N_21646);
or U39327 (N_39327,N_28241,N_24408);
nor U39328 (N_39328,N_25447,N_29359);
xor U39329 (N_39329,N_26218,N_21619);
xnor U39330 (N_39330,N_29933,N_20014);
nand U39331 (N_39331,N_24424,N_27192);
and U39332 (N_39332,N_28360,N_21522);
nor U39333 (N_39333,N_27796,N_21661);
and U39334 (N_39334,N_20740,N_23264);
or U39335 (N_39335,N_21103,N_25626);
and U39336 (N_39336,N_29683,N_26100);
nor U39337 (N_39337,N_22665,N_22317);
nand U39338 (N_39338,N_20935,N_21131);
nor U39339 (N_39339,N_29339,N_27746);
nand U39340 (N_39340,N_21759,N_27935);
nand U39341 (N_39341,N_24987,N_20436);
nand U39342 (N_39342,N_20414,N_24884);
and U39343 (N_39343,N_29178,N_21695);
nand U39344 (N_39344,N_24665,N_27040);
nor U39345 (N_39345,N_21133,N_27800);
or U39346 (N_39346,N_20949,N_23427);
xnor U39347 (N_39347,N_21822,N_23754);
nand U39348 (N_39348,N_26142,N_21257);
xor U39349 (N_39349,N_22245,N_26900);
nor U39350 (N_39350,N_28937,N_25154);
xor U39351 (N_39351,N_25693,N_26574);
nor U39352 (N_39352,N_21071,N_26441);
and U39353 (N_39353,N_29044,N_27772);
or U39354 (N_39354,N_20956,N_26258);
nand U39355 (N_39355,N_21082,N_20410);
and U39356 (N_39356,N_24107,N_28118);
nand U39357 (N_39357,N_28883,N_25256);
nand U39358 (N_39358,N_26577,N_23298);
and U39359 (N_39359,N_26653,N_20869);
xor U39360 (N_39360,N_22803,N_20621);
nor U39361 (N_39361,N_25388,N_28710);
or U39362 (N_39362,N_28114,N_21086);
or U39363 (N_39363,N_24065,N_29723);
nand U39364 (N_39364,N_22065,N_26768);
xor U39365 (N_39365,N_22987,N_23910);
nand U39366 (N_39366,N_24234,N_22447);
xor U39367 (N_39367,N_28519,N_29188);
nor U39368 (N_39368,N_22639,N_25746);
nand U39369 (N_39369,N_29329,N_27898);
xnor U39370 (N_39370,N_28004,N_22153);
and U39371 (N_39371,N_23330,N_28859);
or U39372 (N_39372,N_27922,N_20367);
and U39373 (N_39373,N_26433,N_21846);
xnor U39374 (N_39374,N_22993,N_23043);
nand U39375 (N_39375,N_25734,N_27214);
nand U39376 (N_39376,N_21969,N_20697);
nand U39377 (N_39377,N_28580,N_20298);
and U39378 (N_39378,N_27671,N_28533);
or U39379 (N_39379,N_22268,N_21466);
xnor U39380 (N_39380,N_20870,N_24127);
nor U39381 (N_39381,N_20970,N_26475);
nor U39382 (N_39382,N_27542,N_23839);
and U39383 (N_39383,N_27089,N_21034);
or U39384 (N_39384,N_27025,N_27877);
nand U39385 (N_39385,N_24772,N_29324);
nor U39386 (N_39386,N_26460,N_28315);
or U39387 (N_39387,N_27461,N_23198);
nand U39388 (N_39388,N_24897,N_25444);
or U39389 (N_39389,N_22826,N_22052);
and U39390 (N_39390,N_20165,N_25644);
or U39391 (N_39391,N_26536,N_23545);
and U39392 (N_39392,N_25732,N_22513);
or U39393 (N_39393,N_20111,N_25259);
nor U39394 (N_39394,N_22806,N_20623);
nor U39395 (N_39395,N_24194,N_29631);
or U39396 (N_39396,N_23468,N_29474);
and U39397 (N_39397,N_26999,N_23190);
and U39398 (N_39398,N_25671,N_28772);
nand U39399 (N_39399,N_29351,N_23037);
nand U39400 (N_39400,N_28518,N_28120);
nand U39401 (N_39401,N_22637,N_24958);
nand U39402 (N_39402,N_21229,N_29531);
and U39403 (N_39403,N_29774,N_27572);
nand U39404 (N_39404,N_23527,N_22394);
or U39405 (N_39405,N_29882,N_26635);
xnor U39406 (N_39406,N_26158,N_27778);
nand U39407 (N_39407,N_24002,N_22565);
xnor U39408 (N_39408,N_22713,N_22304);
xor U39409 (N_39409,N_29058,N_22382);
xnor U39410 (N_39410,N_25860,N_26774);
xnor U39411 (N_39411,N_29917,N_21146);
nor U39412 (N_39412,N_22294,N_29485);
xnor U39413 (N_39413,N_24641,N_27410);
xnor U39414 (N_39414,N_26560,N_26729);
nand U39415 (N_39415,N_20250,N_27168);
nand U39416 (N_39416,N_25119,N_22413);
nand U39417 (N_39417,N_24880,N_23115);
or U39418 (N_39418,N_29629,N_27795);
nand U39419 (N_39419,N_27071,N_22620);
or U39420 (N_39420,N_23108,N_21922);
and U39421 (N_39421,N_20397,N_29879);
xnor U39422 (N_39422,N_23723,N_25917);
xnor U39423 (N_39423,N_26774,N_26388);
nor U39424 (N_39424,N_21291,N_26128);
xor U39425 (N_39425,N_28578,N_26870);
nor U39426 (N_39426,N_22821,N_25902);
and U39427 (N_39427,N_27973,N_25861);
xor U39428 (N_39428,N_25645,N_26771);
nand U39429 (N_39429,N_26286,N_21252);
or U39430 (N_39430,N_24804,N_24198);
nor U39431 (N_39431,N_22327,N_29520);
or U39432 (N_39432,N_24322,N_26923);
or U39433 (N_39433,N_20147,N_26321);
nor U39434 (N_39434,N_23913,N_28629);
xor U39435 (N_39435,N_26026,N_26674);
nand U39436 (N_39436,N_29039,N_24330);
nor U39437 (N_39437,N_24710,N_24331);
nor U39438 (N_39438,N_26030,N_22349);
or U39439 (N_39439,N_28941,N_21698);
xnor U39440 (N_39440,N_24876,N_23975);
or U39441 (N_39441,N_28298,N_29191);
and U39442 (N_39442,N_27814,N_25505);
xor U39443 (N_39443,N_23560,N_27318);
or U39444 (N_39444,N_29494,N_23335);
and U39445 (N_39445,N_21037,N_22150);
nor U39446 (N_39446,N_21320,N_25055);
or U39447 (N_39447,N_24133,N_25447);
or U39448 (N_39448,N_21629,N_25138);
and U39449 (N_39449,N_22288,N_29724);
and U39450 (N_39450,N_27068,N_26157);
and U39451 (N_39451,N_22618,N_20113);
nor U39452 (N_39452,N_22628,N_21636);
and U39453 (N_39453,N_29463,N_27691);
nor U39454 (N_39454,N_25358,N_23982);
nand U39455 (N_39455,N_27067,N_22855);
and U39456 (N_39456,N_23965,N_24350);
xnor U39457 (N_39457,N_21246,N_23293);
xnor U39458 (N_39458,N_28576,N_26679);
nand U39459 (N_39459,N_25079,N_21838);
nor U39460 (N_39460,N_28721,N_27943);
nand U39461 (N_39461,N_24099,N_24642);
nand U39462 (N_39462,N_23810,N_22535);
xor U39463 (N_39463,N_21833,N_20153);
nand U39464 (N_39464,N_27148,N_28775);
nand U39465 (N_39465,N_23517,N_28144);
nand U39466 (N_39466,N_29718,N_28423);
nor U39467 (N_39467,N_25192,N_20794);
xor U39468 (N_39468,N_25898,N_22796);
or U39469 (N_39469,N_22483,N_26096);
xnor U39470 (N_39470,N_29775,N_25117);
or U39471 (N_39471,N_25647,N_23120);
xnor U39472 (N_39472,N_28073,N_20483);
or U39473 (N_39473,N_25364,N_25095);
and U39474 (N_39474,N_27271,N_24061);
nor U39475 (N_39475,N_22526,N_28115);
nand U39476 (N_39476,N_25792,N_25150);
and U39477 (N_39477,N_22178,N_28770);
and U39478 (N_39478,N_29966,N_22166);
or U39479 (N_39479,N_21467,N_29398);
and U39480 (N_39480,N_22749,N_25978);
nor U39481 (N_39481,N_28671,N_24242);
nor U39482 (N_39482,N_28476,N_29435);
nor U39483 (N_39483,N_23106,N_22138);
nand U39484 (N_39484,N_27536,N_22433);
xnor U39485 (N_39485,N_27094,N_28418);
nor U39486 (N_39486,N_28743,N_20563);
nor U39487 (N_39487,N_25511,N_27512);
nand U39488 (N_39488,N_20042,N_26173);
nor U39489 (N_39489,N_22473,N_23206);
and U39490 (N_39490,N_21326,N_24639);
or U39491 (N_39491,N_22409,N_28857);
and U39492 (N_39492,N_26033,N_25065);
or U39493 (N_39493,N_22483,N_25362);
and U39494 (N_39494,N_22372,N_25688);
and U39495 (N_39495,N_26133,N_23318);
xor U39496 (N_39496,N_24543,N_26237);
and U39497 (N_39497,N_23950,N_21837);
and U39498 (N_39498,N_25111,N_22086);
or U39499 (N_39499,N_20904,N_25107);
nand U39500 (N_39500,N_29401,N_23189);
and U39501 (N_39501,N_27825,N_28982);
and U39502 (N_39502,N_29905,N_27215);
nand U39503 (N_39503,N_25256,N_26513);
and U39504 (N_39504,N_26426,N_20464);
nor U39505 (N_39505,N_28672,N_23558);
nor U39506 (N_39506,N_25999,N_22958);
or U39507 (N_39507,N_20265,N_22630);
xor U39508 (N_39508,N_26813,N_24421);
nor U39509 (N_39509,N_23954,N_28129);
xor U39510 (N_39510,N_27553,N_21745);
xnor U39511 (N_39511,N_20209,N_21166);
or U39512 (N_39512,N_29613,N_23843);
or U39513 (N_39513,N_26342,N_27628);
and U39514 (N_39514,N_22836,N_23913);
nor U39515 (N_39515,N_29023,N_23067);
xnor U39516 (N_39516,N_27416,N_28948);
nand U39517 (N_39517,N_20434,N_22691);
nor U39518 (N_39518,N_28949,N_24520);
nand U39519 (N_39519,N_26971,N_22228);
xor U39520 (N_39520,N_23381,N_25194);
nand U39521 (N_39521,N_20006,N_26291);
and U39522 (N_39522,N_28308,N_27119);
nand U39523 (N_39523,N_21184,N_22130);
xnor U39524 (N_39524,N_27808,N_29835);
and U39525 (N_39525,N_22805,N_23526);
xnor U39526 (N_39526,N_26835,N_20325);
or U39527 (N_39527,N_20205,N_25744);
nand U39528 (N_39528,N_22952,N_28930);
and U39529 (N_39529,N_24095,N_27388);
xor U39530 (N_39530,N_28472,N_28004);
or U39531 (N_39531,N_23749,N_21138);
and U39532 (N_39532,N_27618,N_22444);
and U39533 (N_39533,N_20832,N_28613);
nor U39534 (N_39534,N_28887,N_29841);
or U39535 (N_39535,N_27845,N_22331);
xor U39536 (N_39536,N_23326,N_28290);
xnor U39537 (N_39537,N_22670,N_21503);
and U39538 (N_39538,N_23399,N_23756);
xor U39539 (N_39539,N_27583,N_25684);
xnor U39540 (N_39540,N_26272,N_28946);
or U39541 (N_39541,N_27806,N_25040);
nor U39542 (N_39542,N_28439,N_25777);
nor U39543 (N_39543,N_24730,N_21106);
nor U39544 (N_39544,N_27689,N_25123);
nand U39545 (N_39545,N_25960,N_21825);
or U39546 (N_39546,N_29507,N_21021);
xnor U39547 (N_39547,N_25256,N_25417);
nand U39548 (N_39548,N_23197,N_28725);
or U39549 (N_39549,N_20840,N_28545);
xor U39550 (N_39550,N_23044,N_26145);
nor U39551 (N_39551,N_25822,N_26354);
nor U39552 (N_39552,N_29287,N_29218);
xnor U39553 (N_39553,N_26466,N_22052);
xor U39554 (N_39554,N_23396,N_24818);
nand U39555 (N_39555,N_26018,N_20777);
nor U39556 (N_39556,N_20626,N_28131);
nand U39557 (N_39557,N_25341,N_29099);
nand U39558 (N_39558,N_27556,N_23083);
xor U39559 (N_39559,N_22463,N_28844);
nor U39560 (N_39560,N_29660,N_20363);
nor U39561 (N_39561,N_25193,N_20434);
nand U39562 (N_39562,N_28285,N_23942);
nor U39563 (N_39563,N_27509,N_26194);
and U39564 (N_39564,N_23427,N_29431);
nor U39565 (N_39565,N_26229,N_22365);
xor U39566 (N_39566,N_21134,N_28821);
nor U39567 (N_39567,N_26994,N_23091);
and U39568 (N_39568,N_20273,N_20309);
or U39569 (N_39569,N_25079,N_26085);
or U39570 (N_39570,N_28719,N_27776);
or U39571 (N_39571,N_23389,N_23166);
and U39572 (N_39572,N_20496,N_25276);
nor U39573 (N_39573,N_26906,N_27228);
and U39574 (N_39574,N_27370,N_26697);
nor U39575 (N_39575,N_26602,N_26505);
nand U39576 (N_39576,N_21040,N_21607);
or U39577 (N_39577,N_24611,N_20977);
nand U39578 (N_39578,N_21990,N_25440);
xor U39579 (N_39579,N_24729,N_21180);
xor U39580 (N_39580,N_26720,N_28554);
xor U39581 (N_39581,N_20664,N_23154);
and U39582 (N_39582,N_27069,N_20347);
nor U39583 (N_39583,N_24419,N_24817);
xnor U39584 (N_39584,N_20783,N_27928);
xor U39585 (N_39585,N_20765,N_25652);
xor U39586 (N_39586,N_27182,N_23459);
nor U39587 (N_39587,N_25014,N_24117);
or U39588 (N_39588,N_22847,N_28693);
or U39589 (N_39589,N_25239,N_25745);
and U39590 (N_39590,N_27094,N_21794);
and U39591 (N_39591,N_25972,N_29522);
nor U39592 (N_39592,N_22351,N_20480);
xnor U39593 (N_39593,N_28099,N_29432);
or U39594 (N_39594,N_22952,N_22923);
nor U39595 (N_39595,N_29187,N_22196);
or U39596 (N_39596,N_26463,N_27959);
xor U39597 (N_39597,N_23516,N_29449);
nand U39598 (N_39598,N_22671,N_26945);
nor U39599 (N_39599,N_22368,N_25607);
and U39600 (N_39600,N_22817,N_20303);
xor U39601 (N_39601,N_23830,N_21980);
xor U39602 (N_39602,N_26754,N_21430);
nand U39603 (N_39603,N_21143,N_27373);
nand U39604 (N_39604,N_29949,N_24511);
nor U39605 (N_39605,N_27084,N_24021);
or U39606 (N_39606,N_25003,N_24630);
nor U39607 (N_39607,N_21539,N_21435);
nand U39608 (N_39608,N_29136,N_24072);
nand U39609 (N_39609,N_29501,N_25283);
nand U39610 (N_39610,N_29746,N_23548);
nor U39611 (N_39611,N_27735,N_21975);
or U39612 (N_39612,N_22912,N_23597);
nand U39613 (N_39613,N_22968,N_28966);
nand U39614 (N_39614,N_26921,N_24784);
and U39615 (N_39615,N_22314,N_22221);
nor U39616 (N_39616,N_24927,N_27983);
or U39617 (N_39617,N_28411,N_23016);
xnor U39618 (N_39618,N_23526,N_25035);
nor U39619 (N_39619,N_26674,N_27336);
nand U39620 (N_39620,N_28743,N_24930);
nand U39621 (N_39621,N_26185,N_25869);
nor U39622 (N_39622,N_27992,N_20488);
nor U39623 (N_39623,N_27353,N_23162);
or U39624 (N_39624,N_20082,N_28862);
and U39625 (N_39625,N_24497,N_26406);
or U39626 (N_39626,N_22057,N_24591);
or U39627 (N_39627,N_21851,N_23294);
nand U39628 (N_39628,N_23065,N_27705);
and U39629 (N_39629,N_21301,N_27822);
xor U39630 (N_39630,N_29549,N_29057);
and U39631 (N_39631,N_26745,N_26198);
or U39632 (N_39632,N_22661,N_26389);
nor U39633 (N_39633,N_23369,N_22154);
or U39634 (N_39634,N_24763,N_26584);
nor U39635 (N_39635,N_21851,N_29065);
nand U39636 (N_39636,N_21673,N_26325);
and U39637 (N_39637,N_26087,N_27197);
xnor U39638 (N_39638,N_26625,N_28057);
nand U39639 (N_39639,N_20635,N_20113);
and U39640 (N_39640,N_22827,N_24853);
or U39641 (N_39641,N_22947,N_20682);
or U39642 (N_39642,N_22176,N_20543);
and U39643 (N_39643,N_29784,N_22161);
nand U39644 (N_39644,N_29236,N_28756);
nand U39645 (N_39645,N_25759,N_20350);
nor U39646 (N_39646,N_22967,N_22958);
xor U39647 (N_39647,N_28048,N_21356);
and U39648 (N_39648,N_20915,N_23616);
nor U39649 (N_39649,N_25217,N_21868);
and U39650 (N_39650,N_26967,N_29591);
and U39651 (N_39651,N_29265,N_28747);
nand U39652 (N_39652,N_20699,N_25051);
nor U39653 (N_39653,N_27627,N_20445);
or U39654 (N_39654,N_26221,N_28079);
and U39655 (N_39655,N_23817,N_21800);
or U39656 (N_39656,N_20086,N_22253);
nand U39657 (N_39657,N_24125,N_28516);
nand U39658 (N_39658,N_20361,N_24786);
and U39659 (N_39659,N_24457,N_26910);
nor U39660 (N_39660,N_24488,N_24828);
and U39661 (N_39661,N_28316,N_29463);
and U39662 (N_39662,N_29599,N_28986);
and U39663 (N_39663,N_26930,N_20692);
nor U39664 (N_39664,N_28841,N_26099);
or U39665 (N_39665,N_20832,N_28827);
or U39666 (N_39666,N_26459,N_24128);
nand U39667 (N_39667,N_22390,N_21873);
xor U39668 (N_39668,N_21136,N_20804);
nor U39669 (N_39669,N_28218,N_25926);
xnor U39670 (N_39670,N_20689,N_29377);
or U39671 (N_39671,N_20919,N_23220);
nor U39672 (N_39672,N_27818,N_24125);
nor U39673 (N_39673,N_20890,N_26538);
and U39674 (N_39674,N_28686,N_28150);
or U39675 (N_39675,N_22235,N_22191);
and U39676 (N_39676,N_26108,N_27813);
xnor U39677 (N_39677,N_27567,N_25994);
nor U39678 (N_39678,N_28372,N_20471);
nand U39679 (N_39679,N_29066,N_20805);
or U39680 (N_39680,N_23910,N_26799);
xnor U39681 (N_39681,N_20621,N_27533);
or U39682 (N_39682,N_26734,N_29877);
nor U39683 (N_39683,N_25162,N_22449);
or U39684 (N_39684,N_27305,N_22743);
and U39685 (N_39685,N_23047,N_27849);
nand U39686 (N_39686,N_23029,N_29086);
nor U39687 (N_39687,N_21141,N_27565);
nor U39688 (N_39688,N_27875,N_28682);
or U39689 (N_39689,N_25379,N_26022);
nor U39690 (N_39690,N_28250,N_20953);
nand U39691 (N_39691,N_23380,N_28154);
nor U39692 (N_39692,N_20157,N_27807);
xor U39693 (N_39693,N_24367,N_24723);
xnor U39694 (N_39694,N_24519,N_29150);
nand U39695 (N_39695,N_26673,N_22464);
nand U39696 (N_39696,N_22781,N_29641);
xnor U39697 (N_39697,N_25838,N_28077);
or U39698 (N_39698,N_25821,N_27948);
nand U39699 (N_39699,N_23831,N_27541);
nor U39700 (N_39700,N_22182,N_21212);
and U39701 (N_39701,N_21431,N_20189);
and U39702 (N_39702,N_22939,N_22378);
xnor U39703 (N_39703,N_20441,N_25275);
and U39704 (N_39704,N_26590,N_26714);
nand U39705 (N_39705,N_21969,N_21132);
and U39706 (N_39706,N_27509,N_26918);
nor U39707 (N_39707,N_24071,N_21372);
nor U39708 (N_39708,N_26298,N_27398);
nor U39709 (N_39709,N_24483,N_23323);
xor U39710 (N_39710,N_21741,N_20613);
nor U39711 (N_39711,N_20742,N_22869);
and U39712 (N_39712,N_24589,N_24608);
or U39713 (N_39713,N_23862,N_26253);
and U39714 (N_39714,N_28372,N_23041);
and U39715 (N_39715,N_22847,N_27852);
or U39716 (N_39716,N_26117,N_28867);
nand U39717 (N_39717,N_20423,N_25975);
nor U39718 (N_39718,N_23181,N_27840);
xnor U39719 (N_39719,N_22837,N_27093);
and U39720 (N_39720,N_20597,N_23254);
nor U39721 (N_39721,N_26107,N_29992);
and U39722 (N_39722,N_21386,N_25787);
nor U39723 (N_39723,N_25463,N_28549);
and U39724 (N_39724,N_26332,N_25832);
nand U39725 (N_39725,N_24410,N_20452);
and U39726 (N_39726,N_22099,N_23281);
and U39727 (N_39727,N_22969,N_21959);
or U39728 (N_39728,N_24976,N_28092);
nor U39729 (N_39729,N_23569,N_20870);
nor U39730 (N_39730,N_20987,N_26285);
nand U39731 (N_39731,N_28130,N_23107);
and U39732 (N_39732,N_25159,N_20733);
nand U39733 (N_39733,N_29507,N_29604);
nand U39734 (N_39734,N_20000,N_25144);
or U39735 (N_39735,N_20764,N_29263);
or U39736 (N_39736,N_25387,N_27487);
or U39737 (N_39737,N_22524,N_21196);
xor U39738 (N_39738,N_28567,N_21959);
and U39739 (N_39739,N_23420,N_24832);
xnor U39740 (N_39740,N_25717,N_27981);
nand U39741 (N_39741,N_23400,N_28496);
xnor U39742 (N_39742,N_26674,N_23453);
xnor U39743 (N_39743,N_23701,N_27041);
or U39744 (N_39744,N_24635,N_26822);
xor U39745 (N_39745,N_25255,N_22974);
nor U39746 (N_39746,N_29528,N_24880);
nor U39747 (N_39747,N_25653,N_22153);
or U39748 (N_39748,N_20103,N_22134);
or U39749 (N_39749,N_22285,N_24143);
or U39750 (N_39750,N_23200,N_26069);
xor U39751 (N_39751,N_21009,N_24589);
and U39752 (N_39752,N_29113,N_21716);
xnor U39753 (N_39753,N_24524,N_21386);
or U39754 (N_39754,N_23988,N_23932);
nand U39755 (N_39755,N_27454,N_28100);
and U39756 (N_39756,N_29447,N_20919);
nor U39757 (N_39757,N_28365,N_28488);
or U39758 (N_39758,N_29236,N_20813);
nor U39759 (N_39759,N_26083,N_24521);
nor U39760 (N_39760,N_28542,N_27134);
xor U39761 (N_39761,N_29522,N_29569);
xnor U39762 (N_39762,N_22861,N_21530);
nor U39763 (N_39763,N_26648,N_25317);
and U39764 (N_39764,N_21991,N_23311);
nand U39765 (N_39765,N_29351,N_27401);
xor U39766 (N_39766,N_25408,N_20348);
nor U39767 (N_39767,N_22537,N_26213);
and U39768 (N_39768,N_24519,N_29941);
xnor U39769 (N_39769,N_24049,N_26645);
xor U39770 (N_39770,N_28852,N_20700);
xnor U39771 (N_39771,N_24897,N_20525);
or U39772 (N_39772,N_23711,N_26944);
nor U39773 (N_39773,N_22126,N_26066);
or U39774 (N_39774,N_23985,N_28373);
and U39775 (N_39775,N_25005,N_21968);
and U39776 (N_39776,N_21138,N_29753);
or U39777 (N_39777,N_27407,N_25788);
nand U39778 (N_39778,N_20533,N_24143);
or U39779 (N_39779,N_23541,N_22213);
nand U39780 (N_39780,N_26122,N_24254);
or U39781 (N_39781,N_29700,N_22402);
or U39782 (N_39782,N_24258,N_27051);
nand U39783 (N_39783,N_26739,N_26175);
nand U39784 (N_39784,N_21317,N_22700);
or U39785 (N_39785,N_21116,N_20739);
or U39786 (N_39786,N_23768,N_26141);
and U39787 (N_39787,N_23025,N_29981);
and U39788 (N_39788,N_20635,N_28029);
xor U39789 (N_39789,N_25742,N_26983);
xnor U39790 (N_39790,N_22308,N_23434);
xnor U39791 (N_39791,N_24796,N_26701);
nor U39792 (N_39792,N_23636,N_20574);
and U39793 (N_39793,N_29241,N_26055);
or U39794 (N_39794,N_27910,N_28693);
and U39795 (N_39795,N_26432,N_28462);
nor U39796 (N_39796,N_28987,N_23364);
xnor U39797 (N_39797,N_21053,N_20962);
xnor U39798 (N_39798,N_20483,N_24712);
nor U39799 (N_39799,N_24654,N_20013);
xor U39800 (N_39800,N_24576,N_20332);
nand U39801 (N_39801,N_27991,N_24632);
nor U39802 (N_39802,N_26378,N_24968);
or U39803 (N_39803,N_22956,N_27266);
or U39804 (N_39804,N_24967,N_29623);
and U39805 (N_39805,N_20883,N_29946);
nor U39806 (N_39806,N_20405,N_25770);
and U39807 (N_39807,N_27663,N_20840);
nand U39808 (N_39808,N_26595,N_20267);
or U39809 (N_39809,N_27640,N_21162);
nand U39810 (N_39810,N_22145,N_29966);
or U39811 (N_39811,N_26482,N_20799);
or U39812 (N_39812,N_23315,N_23600);
nor U39813 (N_39813,N_24388,N_23387);
xor U39814 (N_39814,N_24992,N_27302);
or U39815 (N_39815,N_27182,N_28369);
nor U39816 (N_39816,N_23018,N_26927);
xor U39817 (N_39817,N_29287,N_26781);
xnor U39818 (N_39818,N_20047,N_27381);
nor U39819 (N_39819,N_25649,N_28214);
nor U39820 (N_39820,N_27548,N_20917);
nand U39821 (N_39821,N_27759,N_20562);
nand U39822 (N_39822,N_21919,N_27323);
or U39823 (N_39823,N_23066,N_28152);
xnor U39824 (N_39824,N_25808,N_25405);
or U39825 (N_39825,N_28499,N_21707);
or U39826 (N_39826,N_22397,N_23148);
or U39827 (N_39827,N_29821,N_24527);
xor U39828 (N_39828,N_22370,N_26563);
nor U39829 (N_39829,N_28102,N_26321);
xor U39830 (N_39830,N_29811,N_29777);
nor U39831 (N_39831,N_21380,N_22910);
or U39832 (N_39832,N_20471,N_26662);
or U39833 (N_39833,N_21688,N_22542);
or U39834 (N_39834,N_28281,N_25036);
or U39835 (N_39835,N_29925,N_20523);
or U39836 (N_39836,N_20843,N_22009);
xnor U39837 (N_39837,N_26315,N_20723);
and U39838 (N_39838,N_27772,N_27245);
nand U39839 (N_39839,N_22244,N_22180);
nor U39840 (N_39840,N_23722,N_23312);
xor U39841 (N_39841,N_24603,N_23309);
nand U39842 (N_39842,N_28383,N_25011);
xor U39843 (N_39843,N_20002,N_26496);
and U39844 (N_39844,N_28275,N_23645);
or U39845 (N_39845,N_26532,N_26118);
nor U39846 (N_39846,N_26645,N_22585);
or U39847 (N_39847,N_20642,N_20689);
and U39848 (N_39848,N_28427,N_25500);
or U39849 (N_39849,N_24460,N_23057);
nand U39850 (N_39850,N_23114,N_25434);
nand U39851 (N_39851,N_20252,N_22097);
and U39852 (N_39852,N_23183,N_23807);
xor U39853 (N_39853,N_27972,N_24687);
and U39854 (N_39854,N_23376,N_22158);
nand U39855 (N_39855,N_25764,N_23008);
nor U39856 (N_39856,N_22703,N_28845);
and U39857 (N_39857,N_25750,N_23908);
nand U39858 (N_39858,N_26962,N_20791);
nor U39859 (N_39859,N_23526,N_27151);
nand U39860 (N_39860,N_26180,N_26094);
nor U39861 (N_39861,N_29849,N_20880);
or U39862 (N_39862,N_22937,N_25106);
or U39863 (N_39863,N_23580,N_23069);
nor U39864 (N_39864,N_23699,N_20774);
nor U39865 (N_39865,N_23366,N_21189);
nor U39866 (N_39866,N_20857,N_21278);
and U39867 (N_39867,N_20339,N_27233);
nor U39868 (N_39868,N_26869,N_24926);
nor U39869 (N_39869,N_27413,N_22852);
nand U39870 (N_39870,N_23286,N_26390);
xnor U39871 (N_39871,N_24968,N_26883);
nor U39872 (N_39872,N_29898,N_26914);
or U39873 (N_39873,N_27704,N_24940);
and U39874 (N_39874,N_21646,N_28118);
and U39875 (N_39875,N_26822,N_27750);
nor U39876 (N_39876,N_20887,N_23370);
and U39877 (N_39877,N_26471,N_23496);
nand U39878 (N_39878,N_26837,N_21054);
nor U39879 (N_39879,N_29930,N_23995);
or U39880 (N_39880,N_20318,N_23347);
nand U39881 (N_39881,N_29251,N_29097);
nand U39882 (N_39882,N_26050,N_25463);
and U39883 (N_39883,N_23821,N_27360);
and U39884 (N_39884,N_26141,N_20261);
nand U39885 (N_39885,N_21079,N_21027);
or U39886 (N_39886,N_23991,N_23307);
xor U39887 (N_39887,N_21199,N_22333);
nor U39888 (N_39888,N_24930,N_24761);
xor U39889 (N_39889,N_23242,N_23902);
nand U39890 (N_39890,N_24260,N_24265);
nand U39891 (N_39891,N_29838,N_28937);
nand U39892 (N_39892,N_24566,N_25572);
nand U39893 (N_39893,N_22026,N_27242);
or U39894 (N_39894,N_27236,N_25087);
and U39895 (N_39895,N_20870,N_26636);
and U39896 (N_39896,N_29847,N_20732);
or U39897 (N_39897,N_23916,N_20410);
xnor U39898 (N_39898,N_27429,N_25025);
nand U39899 (N_39899,N_26738,N_27461);
or U39900 (N_39900,N_28095,N_27706);
and U39901 (N_39901,N_22518,N_24230);
xor U39902 (N_39902,N_27598,N_27547);
and U39903 (N_39903,N_23822,N_28669);
xnor U39904 (N_39904,N_26229,N_27679);
nand U39905 (N_39905,N_24271,N_22258);
and U39906 (N_39906,N_23596,N_22945);
nand U39907 (N_39907,N_24464,N_27274);
nand U39908 (N_39908,N_21162,N_25603);
and U39909 (N_39909,N_20899,N_29082);
nor U39910 (N_39910,N_23729,N_24298);
or U39911 (N_39911,N_23885,N_20978);
and U39912 (N_39912,N_24648,N_22467);
nor U39913 (N_39913,N_20403,N_21550);
nand U39914 (N_39914,N_22755,N_20797);
and U39915 (N_39915,N_26809,N_24042);
nor U39916 (N_39916,N_24119,N_29475);
and U39917 (N_39917,N_25855,N_20576);
and U39918 (N_39918,N_23878,N_22075);
and U39919 (N_39919,N_22924,N_24540);
and U39920 (N_39920,N_25137,N_25851);
nand U39921 (N_39921,N_27216,N_23702);
and U39922 (N_39922,N_24956,N_24455);
or U39923 (N_39923,N_28234,N_27951);
nor U39924 (N_39924,N_22468,N_23430);
or U39925 (N_39925,N_26407,N_22906);
xor U39926 (N_39926,N_20607,N_29571);
nor U39927 (N_39927,N_24400,N_21603);
or U39928 (N_39928,N_29634,N_23025);
nand U39929 (N_39929,N_20531,N_20793);
xor U39930 (N_39930,N_29082,N_21833);
nand U39931 (N_39931,N_24898,N_20483);
or U39932 (N_39932,N_27891,N_23346);
or U39933 (N_39933,N_22817,N_23913);
nor U39934 (N_39934,N_20942,N_26410);
or U39935 (N_39935,N_22572,N_22744);
nor U39936 (N_39936,N_23847,N_23273);
nor U39937 (N_39937,N_22758,N_26190);
or U39938 (N_39938,N_29611,N_23192);
nand U39939 (N_39939,N_28834,N_27744);
nor U39940 (N_39940,N_22014,N_26929);
xnor U39941 (N_39941,N_23288,N_20860);
or U39942 (N_39942,N_25443,N_22002);
xnor U39943 (N_39943,N_27282,N_23230);
nor U39944 (N_39944,N_27633,N_22237);
nand U39945 (N_39945,N_26200,N_23768);
and U39946 (N_39946,N_28897,N_27054);
nor U39947 (N_39947,N_25240,N_27321);
nand U39948 (N_39948,N_24873,N_20368);
or U39949 (N_39949,N_25011,N_29984);
xor U39950 (N_39950,N_28277,N_25640);
nand U39951 (N_39951,N_25220,N_25112);
or U39952 (N_39952,N_24795,N_27386);
nor U39953 (N_39953,N_26262,N_28257);
or U39954 (N_39954,N_28975,N_26251);
xor U39955 (N_39955,N_28581,N_24374);
nand U39956 (N_39956,N_21474,N_23528);
nand U39957 (N_39957,N_21847,N_26045);
or U39958 (N_39958,N_24218,N_24274);
and U39959 (N_39959,N_28215,N_26652);
or U39960 (N_39960,N_23681,N_27523);
nand U39961 (N_39961,N_20780,N_29270);
nand U39962 (N_39962,N_21029,N_23773);
nor U39963 (N_39963,N_23425,N_29760);
nand U39964 (N_39964,N_21553,N_25750);
or U39965 (N_39965,N_27587,N_27533);
and U39966 (N_39966,N_23298,N_26636);
and U39967 (N_39967,N_23253,N_21229);
nor U39968 (N_39968,N_24881,N_23661);
and U39969 (N_39969,N_25313,N_22663);
nor U39970 (N_39970,N_27440,N_25251);
xnor U39971 (N_39971,N_22446,N_23180);
and U39972 (N_39972,N_22127,N_24347);
and U39973 (N_39973,N_23089,N_29191);
nor U39974 (N_39974,N_20074,N_21480);
nand U39975 (N_39975,N_24502,N_27945);
nand U39976 (N_39976,N_22267,N_29647);
xnor U39977 (N_39977,N_26627,N_28797);
nand U39978 (N_39978,N_21373,N_24995);
or U39979 (N_39979,N_22251,N_21360);
xor U39980 (N_39980,N_27394,N_20949);
and U39981 (N_39981,N_29196,N_22120);
nand U39982 (N_39982,N_24486,N_22571);
or U39983 (N_39983,N_21536,N_20020);
nand U39984 (N_39984,N_21501,N_24404);
nor U39985 (N_39985,N_27205,N_26787);
nand U39986 (N_39986,N_22756,N_21525);
xnor U39987 (N_39987,N_21035,N_22475);
or U39988 (N_39988,N_26176,N_21113);
or U39989 (N_39989,N_21830,N_22315);
nand U39990 (N_39990,N_20492,N_28147);
nand U39991 (N_39991,N_24530,N_23612);
xor U39992 (N_39992,N_22150,N_20669);
xor U39993 (N_39993,N_22914,N_28990);
nor U39994 (N_39994,N_27415,N_29773);
nor U39995 (N_39995,N_27873,N_25055);
nand U39996 (N_39996,N_26610,N_26787);
or U39997 (N_39997,N_29402,N_22183);
xnor U39998 (N_39998,N_27646,N_29013);
xor U39999 (N_39999,N_24324,N_20952);
nor U40000 (N_40000,N_38233,N_39868);
xnor U40001 (N_40001,N_37856,N_38489);
xnor U40002 (N_40002,N_39138,N_34814);
nand U40003 (N_40003,N_30494,N_33068);
and U40004 (N_40004,N_32166,N_34154);
and U40005 (N_40005,N_35190,N_33019);
nor U40006 (N_40006,N_33841,N_35726);
and U40007 (N_40007,N_30067,N_34585);
or U40008 (N_40008,N_35698,N_36514);
nor U40009 (N_40009,N_37109,N_33315);
and U40010 (N_40010,N_30016,N_38649);
xor U40011 (N_40011,N_32896,N_32149);
nor U40012 (N_40012,N_30648,N_36965);
or U40013 (N_40013,N_38668,N_34685);
nand U40014 (N_40014,N_36688,N_34436);
and U40015 (N_40015,N_38847,N_31439);
nor U40016 (N_40016,N_31029,N_36443);
or U40017 (N_40017,N_38890,N_39132);
nor U40018 (N_40018,N_31742,N_36936);
and U40019 (N_40019,N_39476,N_35624);
nor U40020 (N_40020,N_32176,N_33235);
and U40021 (N_40021,N_38943,N_36609);
nor U40022 (N_40022,N_30337,N_35393);
or U40023 (N_40023,N_35936,N_32475);
nand U40024 (N_40024,N_31339,N_32131);
and U40025 (N_40025,N_35806,N_35203);
nand U40026 (N_40026,N_32290,N_31984);
or U40027 (N_40027,N_38258,N_38633);
or U40028 (N_40028,N_30239,N_30947);
nand U40029 (N_40029,N_36819,N_30764);
nor U40030 (N_40030,N_37031,N_32384);
and U40031 (N_40031,N_32954,N_32917);
nand U40032 (N_40032,N_34198,N_36738);
and U40033 (N_40033,N_37790,N_36914);
nor U40034 (N_40034,N_39991,N_37019);
and U40035 (N_40035,N_36218,N_32926);
xnor U40036 (N_40036,N_32945,N_32338);
and U40037 (N_40037,N_39439,N_35609);
nor U40038 (N_40038,N_36845,N_35439);
or U40039 (N_40039,N_30826,N_35569);
xor U40040 (N_40040,N_34260,N_30715);
nor U40041 (N_40041,N_31510,N_36347);
xnor U40042 (N_40042,N_35909,N_33392);
xor U40043 (N_40043,N_31309,N_34225);
nand U40044 (N_40044,N_38113,N_33554);
nor U40045 (N_40045,N_32367,N_34803);
nor U40046 (N_40046,N_34243,N_35181);
or U40047 (N_40047,N_35183,N_35602);
and U40048 (N_40048,N_32456,N_34210);
xnor U40049 (N_40049,N_32786,N_32471);
and U40050 (N_40050,N_34168,N_35968);
nand U40051 (N_40051,N_30877,N_30362);
xnor U40052 (N_40052,N_34067,N_33510);
nand U40053 (N_40053,N_36360,N_39222);
or U40054 (N_40054,N_31115,N_37386);
nand U40055 (N_40055,N_36850,N_31422);
nor U40056 (N_40056,N_34603,N_36289);
xor U40057 (N_40057,N_39905,N_33916);
nor U40058 (N_40058,N_31361,N_37393);
and U40059 (N_40059,N_39520,N_33327);
xnor U40060 (N_40060,N_34238,N_32611);
nand U40061 (N_40061,N_36250,N_39725);
xnor U40062 (N_40062,N_30476,N_34794);
and U40063 (N_40063,N_35350,N_32869);
nand U40064 (N_40064,N_34460,N_38672);
or U40065 (N_40065,N_31239,N_32282);
nand U40066 (N_40066,N_37780,N_37760);
and U40067 (N_40067,N_38375,N_33240);
xor U40068 (N_40068,N_35591,N_38423);
nand U40069 (N_40069,N_33982,N_38920);
xor U40070 (N_40070,N_34458,N_34720);
xor U40071 (N_40071,N_39238,N_31694);
xnor U40072 (N_40072,N_30772,N_38033);
nor U40073 (N_40073,N_32960,N_33662);
nand U40074 (N_40074,N_38590,N_37000);
or U40075 (N_40075,N_36026,N_36883);
nand U40076 (N_40076,N_35051,N_36916);
nor U40077 (N_40077,N_33179,N_33350);
nor U40078 (N_40078,N_38146,N_37890);
nand U40079 (N_40079,N_31637,N_30962);
or U40080 (N_40080,N_35037,N_30457);
xor U40081 (N_40081,N_34221,N_36253);
nor U40082 (N_40082,N_31921,N_35911);
or U40083 (N_40083,N_32705,N_38108);
nor U40084 (N_40084,N_37088,N_34641);
and U40085 (N_40085,N_35039,N_39206);
nor U40086 (N_40086,N_33170,N_30769);
nor U40087 (N_40087,N_35021,N_35402);
and U40088 (N_40088,N_34783,N_33022);
nand U40089 (N_40089,N_30680,N_38287);
xnor U40090 (N_40090,N_34751,N_30987);
nand U40091 (N_40091,N_36411,N_31167);
or U40092 (N_40092,N_35633,N_36752);
nor U40093 (N_40093,N_34982,N_39647);
or U40094 (N_40094,N_30612,N_31892);
or U40095 (N_40095,N_36869,N_38817);
nand U40096 (N_40096,N_37273,N_39140);
or U40097 (N_40097,N_34099,N_32362);
nand U40098 (N_40098,N_33529,N_36586);
nand U40099 (N_40099,N_34676,N_36406);
nand U40100 (N_40100,N_34507,N_34438);
and U40101 (N_40101,N_37551,N_35866);
and U40102 (N_40102,N_31389,N_34935);
or U40103 (N_40103,N_34249,N_39244);
and U40104 (N_40104,N_34505,N_34715);
and U40105 (N_40105,N_37538,N_36398);
xor U40106 (N_40106,N_38475,N_39605);
or U40107 (N_40107,N_31477,N_35538);
or U40108 (N_40108,N_33706,N_31311);
nand U40109 (N_40109,N_31137,N_35138);
nor U40110 (N_40110,N_34234,N_31601);
nor U40111 (N_40111,N_39954,N_33214);
xnor U40112 (N_40112,N_36113,N_31121);
nor U40113 (N_40113,N_37134,N_31142);
nand U40114 (N_40114,N_32915,N_39886);
or U40115 (N_40115,N_32759,N_31472);
nand U40116 (N_40116,N_31245,N_30647);
nand U40117 (N_40117,N_31990,N_38560);
xnor U40118 (N_40118,N_35060,N_35695);
or U40119 (N_40119,N_38265,N_37496);
nand U40120 (N_40120,N_37243,N_34555);
and U40121 (N_40121,N_35234,N_39943);
xor U40122 (N_40122,N_33990,N_34677);
and U40123 (N_40123,N_39553,N_36383);
or U40124 (N_40124,N_30874,N_37422);
or U40125 (N_40125,N_33857,N_35781);
xor U40126 (N_40126,N_31809,N_33863);
and U40127 (N_40127,N_32267,N_35425);
or U40128 (N_40128,N_31242,N_33588);
or U40129 (N_40129,N_36654,N_32928);
or U40130 (N_40130,N_37618,N_33285);
nor U40131 (N_40131,N_33267,N_33246);
xnor U40132 (N_40132,N_30713,N_36891);
xor U40133 (N_40133,N_39075,N_31816);
or U40134 (N_40134,N_38190,N_30072);
and U40135 (N_40135,N_39154,N_35783);
nor U40136 (N_40136,N_34078,N_35292);
xor U40137 (N_40137,N_37535,N_32665);
or U40138 (N_40138,N_39374,N_35755);
nor U40139 (N_40139,N_35071,N_31112);
xor U40140 (N_40140,N_33698,N_32146);
nor U40141 (N_40141,N_30336,N_34472);
and U40142 (N_40142,N_37991,N_34030);
or U40143 (N_40143,N_39980,N_37762);
and U40144 (N_40144,N_38861,N_38088);
or U40145 (N_40145,N_36039,N_37146);
nor U40146 (N_40146,N_39761,N_36774);
nand U40147 (N_40147,N_34039,N_35644);
xor U40148 (N_40148,N_37455,N_32527);
xor U40149 (N_40149,N_38786,N_38019);
or U40150 (N_40150,N_38568,N_38179);
nand U40151 (N_40151,N_32368,N_39939);
xor U40152 (N_40152,N_35958,N_38050);
xnor U40153 (N_40153,N_32407,N_36479);
or U40154 (N_40154,N_33561,N_39455);
and U40155 (N_40155,N_37728,N_38855);
or U40156 (N_40156,N_36804,N_32667);
and U40157 (N_40157,N_32138,N_32593);
and U40158 (N_40158,N_35450,N_36622);
xor U40159 (N_40159,N_39900,N_36651);
and U40160 (N_40160,N_30298,N_39107);
nand U40161 (N_40161,N_36298,N_33424);
and U40162 (N_40162,N_37521,N_39544);
xnor U40163 (N_40163,N_31032,N_37903);
xor U40164 (N_40164,N_38009,N_31876);
and U40165 (N_40165,N_37794,N_38788);
xor U40166 (N_40166,N_39371,N_32518);
or U40167 (N_40167,N_31075,N_38820);
or U40168 (N_40168,N_36970,N_35740);
and U40169 (N_40169,N_39670,N_31712);
nor U40170 (N_40170,N_37705,N_39551);
or U40171 (N_40171,N_31583,N_30477);
or U40172 (N_40172,N_39349,N_31359);
nand U40173 (N_40173,N_34850,N_36451);
nand U40174 (N_40174,N_32343,N_38770);
or U40175 (N_40175,N_30415,N_30423);
and U40176 (N_40176,N_39250,N_34787);
nor U40177 (N_40177,N_30940,N_30427);
nand U40178 (N_40178,N_37124,N_30500);
or U40179 (N_40179,N_31114,N_30075);
nand U40180 (N_40180,N_34601,N_30810);
nor U40181 (N_40181,N_30777,N_31053);
xnor U40182 (N_40182,N_33248,N_37465);
or U40183 (N_40183,N_39624,N_37061);
nand U40184 (N_40184,N_39085,N_39136);
or U40185 (N_40185,N_32326,N_34267);
nor U40186 (N_40186,N_39273,N_39828);
or U40187 (N_40187,N_36069,N_32971);
and U40188 (N_40188,N_38882,N_37044);
nor U40189 (N_40189,N_33448,N_31399);
nor U40190 (N_40190,N_37796,N_39674);
nor U40191 (N_40191,N_33385,N_32460);
nand U40192 (N_40192,N_33276,N_36710);
or U40193 (N_40193,N_39762,N_39470);
nor U40194 (N_40194,N_31039,N_37433);
or U40195 (N_40195,N_37605,N_30756);
or U40196 (N_40196,N_31341,N_37201);
xor U40197 (N_40197,N_36226,N_35990);
or U40198 (N_40198,N_37964,N_33570);
and U40199 (N_40199,N_36001,N_33941);
nor U40200 (N_40200,N_32724,N_38246);
and U40201 (N_40201,N_37288,N_31141);
or U40202 (N_40202,N_32752,N_31171);
and U40203 (N_40203,N_35570,N_31005);
xnor U40204 (N_40204,N_31286,N_36273);
and U40205 (N_40205,N_30552,N_38018);
or U40206 (N_40206,N_34333,N_39073);
nor U40207 (N_40207,N_32871,N_35555);
and U40208 (N_40208,N_39740,N_37557);
and U40209 (N_40209,N_33663,N_33013);
or U40210 (N_40210,N_32271,N_30884);
nand U40211 (N_40211,N_39743,N_34919);
and U40212 (N_40212,N_31549,N_34911);
nor U40213 (N_40213,N_30089,N_38413);
nand U40214 (N_40214,N_31230,N_31046);
xor U40215 (N_40215,N_37450,N_32428);
nor U40216 (N_40216,N_38397,N_31902);
nor U40217 (N_40217,N_35403,N_30311);
and U40218 (N_40218,N_31554,N_38309);
xnor U40219 (N_40219,N_34964,N_33270);
xor U40220 (N_40220,N_33932,N_35734);
or U40221 (N_40221,N_35691,N_39744);
nor U40222 (N_40222,N_36396,N_30235);
or U40223 (N_40223,N_36574,N_35006);
xnor U40224 (N_40224,N_35153,N_31219);
nand U40225 (N_40225,N_31837,N_39189);
and U40226 (N_40226,N_34877,N_32336);
and U40227 (N_40227,N_34960,N_34971);
nand U40228 (N_40228,N_39949,N_36865);
nor U40229 (N_40229,N_34204,N_30246);
nor U40230 (N_40230,N_39513,N_33413);
nand U40231 (N_40231,N_38099,N_38778);
and U40232 (N_40232,N_32785,N_30357);
or U40233 (N_40233,N_38735,N_37920);
or U40234 (N_40234,N_31739,N_35091);
nor U40235 (N_40235,N_30922,N_30852);
nand U40236 (N_40236,N_32615,N_31002);
nand U40237 (N_40237,N_30687,N_34366);
and U40238 (N_40238,N_32200,N_38254);
xnor U40239 (N_40239,N_33035,N_34388);
nand U40240 (N_40240,N_30578,N_35358);
and U40241 (N_40241,N_34371,N_32897);
nor U40242 (N_40242,N_37581,N_37381);
or U40243 (N_40243,N_38277,N_39519);
nand U40244 (N_40244,N_38355,N_39072);
nand U40245 (N_40245,N_33360,N_39607);
nand U40246 (N_40246,N_32463,N_34923);
nor U40247 (N_40247,N_38046,N_30272);
nor U40248 (N_40248,N_36177,N_37307);
or U40249 (N_40249,N_37841,N_33719);
and U40250 (N_40250,N_35194,N_37274);
nor U40251 (N_40251,N_38462,N_36367);
nor U40252 (N_40252,N_36811,N_37498);
xor U40253 (N_40253,N_39254,N_31486);
or U40254 (N_40254,N_33247,N_35387);
and U40255 (N_40255,N_35080,N_38272);
and U40256 (N_40256,N_39281,N_32633);
xor U40257 (N_40257,N_33571,N_30328);
and U40258 (N_40258,N_30491,N_39533);
or U40259 (N_40259,N_32644,N_35949);
and U40260 (N_40260,N_38961,N_36335);
nor U40261 (N_40261,N_32693,N_35798);
xor U40262 (N_40262,N_33381,N_37167);
nor U40263 (N_40263,N_38056,N_37731);
xnor U40264 (N_40264,N_31686,N_39277);
or U40265 (N_40265,N_39153,N_31778);
xor U40266 (N_40266,N_34189,N_30860);
xnor U40267 (N_40267,N_34931,N_32868);
or U40268 (N_40268,N_37143,N_31456);
nor U40269 (N_40269,N_39894,N_32266);
xor U40270 (N_40270,N_33044,N_36709);
xnor U40271 (N_40271,N_38203,N_34311);
nor U40272 (N_40272,N_32543,N_31267);
nor U40273 (N_40273,N_30448,N_30236);
nand U40274 (N_40274,N_39611,N_30260);
and U40275 (N_40275,N_37305,N_37036);
and U40276 (N_40276,N_35529,N_36402);
xnor U40277 (N_40277,N_35662,N_38352);
nand U40278 (N_40278,N_35852,N_32668);
nor U40279 (N_40279,N_34824,N_35433);
nor U40280 (N_40280,N_35581,N_34018);
nand U40281 (N_40281,N_32302,N_37816);
nor U40282 (N_40282,N_32046,N_38438);
nand U40283 (N_40283,N_34266,N_38814);
nand U40284 (N_40284,N_32060,N_36392);
nor U40285 (N_40285,N_37468,N_32062);
nand U40286 (N_40286,N_36087,N_33676);
nor U40287 (N_40287,N_30224,N_31275);
and U40288 (N_40288,N_37162,N_36745);
nor U40289 (N_40289,N_34227,N_30579);
and U40290 (N_40290,N_33707,N_33902);
nor U40291 (N_40291,N_33136,N_39305);
xor U40292 (N_40292,N_38694,N_31363);
xnor U40293 (N_40293,N_36134,N_39203);
or U40294 (N_40294,N_31836,N_33202);
xor U40295 (N_40295,N_32030,N_39695);
and U40296 (N_40296,N_33813,N_38754);
xnor U40297 (N_40297,N_31128,N_30694);
or U40298 (N_40298,N_32755,N_32016);
and U40299 (N_40299,N_31299,N_33630);
and U40300 (N_40300,N_39962,N_35354);
and U40301 (N_40301,N_33258,N_36687);
or U40302 (N_40302,N_30917,N_30542);
nand U40303 (N_40303,N_38999,N_31026);
or U40304 (N_40304,N_30291,N_32841);
or U40305 (N_40305,N_37436,N_32956);
xor U40306 (N_40306,N_34553,N_34009);
xnor U40307 (N_40307,N_36433,N_34322);
or U40308 (N_40308,N_37364,N_39580);
nand U40309 (N_40309,N_34978,N_38634);
or U40310 (N_40310,N_32637,N_33249);
or U40311 (N_40311,N_38874,N_35147);
nor U40312 (N_40312,N_39266,N_33727);
nand U40313 (N_40313,N_38115,N_30946);
or U40314 (N_40314,N_31703,N_39229);
xnor U40315 (N_40315,N_39411,N_38952);
nand U40316 (N_40316,N_37908,N_38889);
xor U40317 (N_40317,N_33898,N_30114);
nand U40318 (N_40318,N_35573,N_39663);
xor U40319 (N_40319,N_31704,N_33298);
nand U40320 (N_40320,N_36143,N_32605);
nand U40321 (N_40321,N_33810,N_35562);
nand U40322 (N_40322,N_33884,N_31869);
nand U40323 (N_40323,N_33809,N_30540);
and U40324 (N_40324,N_36927,N_33130);
and U40325 (N_40325,N_38981,N_34413);
xnor U40326 (N_40326,N_33295,N_36426);
nand U40327 (N_40327,N_33799,N_31807);
nor U40328 (N_40328,N_33769,N_31130);
nand U40329 (N_40329,N_30014,N_36959);
and U40330 (N_40330,N_30264,N_39158);
and U40331 (N_40331,N_30591,N_32329);
nand U40332 (N_40332,N_37980,N_39155);
and U40333 (N_40333,N_33187,N_33736);
nand U40334 (N_40334,N_33604,N_35255);
nand U40335 (N_40335,N_34337,N_31256);
or U40336 (N_40336,N_31159,N_32183);
xnor U40337 (N_40337,N_39854,N_38350);
nand U40338 (N_40338,N_36613,N_38774);
nor U40339 (N_40339,N_35957,N_30804);
nor U40340 (N_40340,N_39756,N_34359);
nand U40341 (N_40341,N_34593,N_35647);
and U40342 (N_40342,N_34456,N_39881);
or U40343 (N_40343,N_34374,N_38026);
or U40344 (N_40344,N_37778,N_38122);
nor U40345 (N_40345,N_36837,N_31280);
nand U40346 (N_40346,N_37598,N_30021);
nor U40347 (N_40347,N_30570,N_32311);
and U40348 (N_40348,N_39709,N_37101);
or U40349 (N_40349,N_34949,N_35200);
or U40350 (N_40350,N_30693,N_35811);
nor U40351 (N_40351,N_39387,N_38111);
or U40352 (N_40352,N_31711,N_32491);
nor U40353 (N_40353,N_35047,N_39822);
nor U40354 (N_40354,N_35337,N_38683);
xnor U40355 (N_40355,N_31706,N_38296);
nor U40356 (N_40356,N_37139,N_35092);
xnor U40357 (N_40357,N_33182,N_38541);
xnor U40358 (N_40358,N_34755,N_36728);
nor U40359 (N_40359,N_36708,N_35373);
and U40360 (N_40360,N_35437,N_35085);
nor U40361 (N_40361,N_36390,N_38704);
nand U40362 (N_40362,N_31860,N_37449);
or U40363 (N_40363,N_31343,N_39495);
nor U40364 (N_40364,N_36748,N_36921);
nor U40365 (N_40365,N_30001,N_32067);
nor U40366 (N_40366,N_32563,N_35696);
xor U40367 (N_40367,N_38414,N_39036);
and U40368 (N_40368,N_33256,N_36422);
xnor U40369 (N_40369,N_33271,N_36155);
xor U40370 (N_40370,N_31191,N_38592);
and U40371 (N_40371,N_38665,N_30341);
nor U40372 (N_40372,N_31063,N_36773);
xnor U40373 (N_40373,N_38734,N_35064);
and U40374 (N_40374,N_37713,N_30100);
nand U40375 (N_40375,N_31088,N_35222);
nand U40376 (N_40376,N_34790,N_34652);
or U40377 (N_40377,N_36189,N_32119);
nor U40378 (N_40378,N_30041,N_34180);
nand U40379 (N_40379,N_33610,N_31293);
xnor U40380 (N_40380,N_37302,N_30516);
nand U40381 (N_40381,N_30430,N_38726);
nor U40382 (N_40382,N_32419,N_32620);
and U40383 (N_40383,N_39948,N_30938);
nor U40384 (N_40384,N_30018,N_36193);
nand U40385 (N_40385,N_36064,N_36278);
xnor U40386 (N_40386,N_30678,N_37905);
or U40387 (N_40387,N_33948,N_30546);
or U40388 (N_40388,N_32347,N_38176);
xor U40389 (N_40389,N_38196,N_33127);
xnor U40390 (N_40390,N_35704,N_35083);
or U40391 (N_40391,N_30285,N_32624);
nand U40392 (N_40392,N_34177,N_30143);
and U40393 (N_40393,N_35599,N_36864);
xor U40394 (N_40394,N_35684,N_35802);
and U40395 (N_40395,N_36307,N_35854);
and U40396 (N_40396,N_35478,N_34797);
and U40397 (N_40397,N_33687,N_36697);
or U40398 (N_40398,N_37111,N_31423);
nor U40399 (N_40399,N_35414,N_33312);
xor U40400 (N_40400,N_34868,N_38432);
nand U40401 (N_40401,N_32320,N_32660);
xor U40402 (N_40402,N_33504,N_33671);
nor U40403 (N_40403,N_38412,N_30253);
nor U40404 (N_40404,N_30963,N_30558);
and U40405 (N_40405,N_38337,N_33917);
nor U40406 (N_40406,N_32949,N_35687);
xor U40407 (N_40407,N_30805,N_34749);
and U40408 (N_40408,N_36279,N_30327);
nand U40409 (N_40409,N_32001,N_32211);
nand U40410 (N_40410,N_37332,N_38699);
nor U40411 (N_40411,N_37203,N_35188);
nor U40412 (N_40412,N_30729,N_35232);
and U40413 (N_40413,N_37370,N_34182);
xnor U40414 (N_40414,N_30205,N_38135);
and U40415 (N_40415,N_39121,N_34286);
nand U40416 (N_40416,N_38079,N_36917);
nor U40417 (N_40417,N_34729,N_31730);
nand U40418 (N_40418,N_37893,N_38869);
nand U40419 (N_40419,N_36540,N_36236);
or U40420 (N_40420,N_37572,N_35679);
xor U40421 (N_40421,N_35423,N_31524);
nand U40422 (N_40422,N_34402,N_34918);
and U40423 (N_40423,N_32465,N_35828);
and U40424 (N_40424,N_38727,N_37089);
nand U40425 (N_40425,N_35572,N_32650);
and U40426 (N_40426,N_34075,N_39361);
nand U40427 (N_40427,N_34002,N_34951);
nor U40428 (N_40428,N_35861,N_39299);
xnor U40429 (N_40429,N_37529,N_38429);
xnor U40430 (N_40430,N_33176,N_33865);
nor U40431 (N_40431,N_37859,N_38676);
nand U40432 (N_40432,N_35473,N_33363);
nor U40433 (N_40433,N_39440,N_33404);
nand U40434 (N_40434,N_32369,N_36024);
and U40435 (N_40435,N_31721,N_33649);
and U40436 (N_40436,N_32588,N_34823);
nor U40437 (N_40437,N_32026,N_30058);
nor U40438 (N_40438,N_32074,N_39983);
and U40439 (N_40439,N_31094,N_31960);
xnor U40440 (N_40440,N_39546,N_33152);
or U40441 (N_40441,N_37073,N_30742);
or U40442 (N_40442,N_38958,N_31173);
nor U40443 (N_40443,N_33343,N_38746);
or U40444 (N_40444,N_32127,N_39007);
xor U40445 (N_40445,N_34459,N_37029);
and U40446 (N_40446,N_31751,N_34372);
or U40447 (N_40447,N_31584,N_35162);
nor U40448 (N_40448,N_38776,N_31880);
and U40449 (N_40449,N_36513,N_39882);
nor U40450 (N_40450,N_39481,N_35163);
or U40451 (N_40451,N_37764,N_38224);
xor U40452 (N_40452,N_32412,N_30712);
nand U40453 (N_40453,N_36757,N_39052);
nor U40454 (N_40454,N_31365,N_37403);
nand U40455 (N_40455,N_38101,N_33396);
or U40456 (N_40456,N_33626,N_38671);
nor U40457 (N_40457,N_33303,N_33429);
xnor U40458 (N_40458,N_32700,N_39282);
nor U40459 (N_40459,N_39050,N_35673);
or U40460 (N_40460,N_34389,N_34491);
xor U40461 (N_40461,N_34721,N_32036);
or U40462 (N_40462,N_35179,N_36625);
xnor U40463 (N_40463,N_34791,N_32743);
nand U40464 (N_40464,N_39726,N_33241);
nand U40465 (N_40465,N_36665,N_36399);
and U40466 (N_40466,N_39407,N_30836);
nor U40467 (N_40467,N_39554,N_32510);
and U40468 (N_40468,N_30774,N_31765);
and U40469 (N_40469,N_39641,N_35978);
or U40470 (N_40470,N_39212,N_31530);
nand U40471 (N_40471,N_30644,N_36611);
nand U40472 (N_40472,N_39175,N_31125);
or U40473 (N_40473,N_33960,N_32052);
or U40474 (N_40474,N_33839,N_36624);
and U40475 (N_40475,N_35542,N_36681);
or U40476 (N_40476,N_31935,N_34616);
nor U40477 (N_40477,N_33837,N_34361);
and U40478 (N_40478,N_33503,N_31487);
nand U40479 (N_40479,N_36284,N_33376);
nor U40480 (N_40480,N_38178,N_30656);
nand U40481 (N_40481,N_34090,N_30345);
nand U40482 (N_40482,N_35801,N_32629);
and U40483 (N_40483,N_34280,N_37060);
xnor U40484 (N_40484,N_35728,N_33164);
or U40485 (N_40485,N_32494,N_35767);
nor U40486 (N_40486,N_39433,N_31193);
nand U40487 (N_40487,N_31769,N_39532);
xnor U40488 (N_40488,N_36594,N_32358);
or U40489 (N_40489,N_35355,N_32316);
and U40490 (N_40490,N_33597,N_33617);
xor U40491 (N_40491,N_35191,N_37566);
nand U40492 (N_40492,N_38660,N_33511);
or U40493 (N_40493,N_38312,N_36018);
and U40494 (N_40494,N_34921,N_32998);
xor U40495 (N_40495,N_39542,N_32064);
xor U40496 (N_40496,N_37136,N_36491);
nor U40497 (N_40497,N_35744,N_39745);
nand U40498 (N_40498,N_30377,N_36702);
and U40499 (N_40499,N_34520,N_34289);
nand U40500 (N_40500,N_31255,N_37532);
xor U40501 (N_40501,N_35084,N_30390);
nand U40502 (N_40502,N_37401,N_32228);
nand U40503 (N_40503,N_32704,N_39069);
and U40504 (N_40504,N_37802,N_38362);
and U40505 (N_40505,N_35263,N_37059);
or U40506 (N_40506,N_30893,N_32215);
nor U40507 (N_40507,N_38801,N_33752);
xor U40508 (N_40508,N_35258,N_36458);
nand U40509 (N_40509,N_33382,N_33582);
and U40510 (N_40510,N_37834,N_34736);
and U40511 (N_40511,N_34347,N_33641);
xor U40512 (N_40512,N_31986,N_31673);
xnor U40513 (N_40513,N_33682,N_34745);
or U40514 (N_40514,N_32125,N_38327);
and U40515 (N_40515,N_30355,N_36438);
nand U40516 (N_40516,N_34469,N_32532);
nand U40517 (N_40517,N_38476,N_38338);
nand U40518 (N_40518,N_39182,N_31631);
xnor U40519 (N_40519,N_36414,N_31183);
or U40520 (N_40520,N_30966,N_31682);
and U40521 (N_40521,N_32858,N_37392);
nor U40522 (N_40522,N_36371,N_34999);
nand U40523 (N_40523,N_34080,N_37216);
and U40524 (N_40524,N_32691,N_37596);
nand U40525 (N_40525,N_36151,N_34480);
xnor U40526 (N_40526,N_35946,N_39379);
xor U40527 (N_40527,N_31384,N_36338);
nand U40528 (N_40528,N_36992,N_35565);
or U40529 (N_40529,N_37625,N_33168);
nand U40530 (N_40530,N_36052,N_31260);
and U40531 (N_40531,N_30146,N_30149);
nand U40532 (N_40532,N_38532,N_35556);
nand U40533 (N_40533,N_38910,N_38791);
or U40534 (N_40534,N_30164,N_39319);
and U40535 (N_40535,N_39497,N_39741);
and U40536 (N_40536,N_30740,N_33347);
xor U40537 (N_40537,N_34944,N_39522);
or U40538 (N_40538,N_33577,N_39101);
nand U40539 (N_40539,N_39561,N_37079);
and U40540 (N_40540,N_36904,N_34316);
and U40541 (N_40541,N_36867,N_32772);
nor U40542 (N_40542,N_38340,N_35134);
nand U40543 (N_40543,N_39099,N_38667);
nor U40544 (N_40544,N_38709,N_30853);
xor U40545 (N_40545,N_30824,N_35730);
and U40546 (N_40546,N_33342,N_34220);
nand U40547 (N_40547,N_35554,N_33756);
and U40548 (N_40548,N_38566,N_35523);
and U40549 (N_40549,N_32889,N_39657);
or U40550 (N_40550,N_36868,N_34159);
xnor U40551 (N_40551,N_30974,N_34183);
nand U40552 (N_40552,N_39797,N_37934);
or U40553 (N_40553,N_31527,N_32781);
and U40554 (N_40554,N_34429,N_32466);
nand U40555 (N_40555,N_30333,N_31322);
nand U40556 (N_40556,N_37775,N_32378);
nor U40557 (N_40557,N_33485,N_37090);
and U40558 (N_40558,N_30068,N_35316);
nand U40559 (N_40559,N_39342,N_38673);
or U40560 (N_40560,N_32340,N_37667);
xnor U40561 (N_40561,N_37617,N_36597);
nand U40562 (N_40562,N_34500,N_39162);
nand U40563 (N_40563,N_32737,N_38530);
xor U40564 (N_40564,N_34060,N_39569);
or U40565 (N_40565,N_36138,N_31052);
nand U40566 (N_40566,N_38409,N_38184);
and U40567 (N_40567,N_36259,N_30614);
xor U40568 (N_40568,N_37607,N_39995);
nor U40569 (N_40569,N_34156,N_32009);
or U40570 (N_40570,N_31186,N_35210);
and U40571 (N_40571,N_35130,N_32315);
nor U40572 (N_40572,N_36517,N_36034);
nand U40573 (N_40573,N_31690,N_38798);
nand U40574 (N_40574,N_32421,N_32108);
xnor U40575 (N_40575,N_37540,N_31151);
nor U40576 (N_40576,N_36793,N_33742);
nand U40577 (N_40577,N_37198,N_30807);
nor U40578 (N_40578,N_32337,N_39722);
nand U40579 (N_40579,N_30732,N_35873);
nor U40580 (N_40580,N_37810,N_31887);
or U40581 (N_40581,N_39872,N_34882);
xnor U40582 (N_40582,N_31226,N_33879);
nand U40583 (N_40583,N_37426,N_35754);
and U40584 (N_40584,N_38339,N_39139);
and U40585 (N_40585,N_35160,N_36099);
and U40586 (N_40586,N_33095,N_37851);
nor U40587 (N_40587,N_31789,N_30698);
nand U40588 (N_40588,N_34167,N_38015);
or U40589 (N_40589,N_39823,N_31475);
and U40590 (N_40590,N_34406,N_30174);
nand U40591 (N_40591,N_34993,N_37842);
and U40592 (N_40592,N_34261,N_36325);
or U40593 (N_40593,N_30761,N_36198);
and U40594 (N_40594,N_32033,N_35773);
and U40595 (N_40595,N_34717,N_39089);
nor U40596 (N_40596,N_32754,N_32497);
xnor U40597 (N_40597,N_31969,N_36790);
nand U40598 (N_40598,N_37317,N_38942);
nor U40599 (N_40599,N_34735,N_38925);
xnor U40600 (N_40600,N_38784,N_39738);
or U40601 (N_40601,N_34258,N_35849);
or U40602 (N_40602,N_32892,N_36723);
xor U40603 (N_40603,N_38074,N_31369);
nor U40604 (N_40604,N_30984,N_36410);
xor U40605 (N_40605,N_37161,N_31496);
nand U40606 (N_40606,N_36675,N_39248);
nand U40607 (N_40607,N_36108,N_39770);
or U40608 (N_40608,N_35997,N_38769);
xor U40609 (N_40609,N_34409,N_33470);
nand U40610 (N_40610,N_33123,N_31815);
or U40611 (N_40611,N_34345,N_38702);
nand U40612 (N_40612,N_33491,N_36830);
or U40613 (N_40613,N_34375,N_30123);
and U40614 (N_40614,N_37440,N_35750);
nand U40615 (N_40615,N_30703,N_32546);
nor U40616 (N_40616,N_34544,N_34961);
xnor U40617 (N_40617,N_31627,N_37456);
or U40618 (N_40618,N_30059,N_35032);
and U40619 (N_40619,N_35923,N_31517);
nor U40620 (N_40620,N_37464,N_30889);
and U40621 (N_40621,N_31215,N_38017);
nor U40622 (N_40622,N_39168,N_34068);
nor U40623 (N_40623,N_35295,N_36575);
and U40624 (N_40624,N_30878,N_39176);
nor U40625 (N_40625,N_35118,N_36776);
nor U40626 (N_40626,N_31908,N_33608);
nor U40627 (N_40627,N_38039,N_32760);
nand U40628 (N_40628,N_39157,N_37133);
xnor U40629 (N_40629,N_31907,N_39893);
nor U40630 (N_40630,N_32161,N_30706);
xor U40631 (N_40631,N_32547,N_36008);
and U40632 (N_40632,N_32521,N_37582);
and U40633 (N_40633,N_38471,N_35380);
and U40634 (N_40634,N_33581,N_32366);
nor U40635 (N_40635,N_38097,N_39926);
or U40636 (N_40636,N_36703,N_36870);
nor U40637 (N_40637,N_37281,N_32703);
nor U40638 (N_40638,N_34471,N_35532);
nand U40639 (N_40639,N_37484,N_31557);
xor U40640 (N_40640,N_34554,N_30073);
xor U40641 (N_40641,N_37628,N_33487);
nand U40642 (N_40642,N_30126,N_36375);
nor U40643 (N_40643,N_30730,N_38659);
xnor U40644 (N_40644,N_38411,N_31893);
nor U40645 (N_40645,N_34661,N_37724);
nand U40646 (N_40646,N_31597,N_39537);
or U40647 (N_40647,N_30196,N_30047);
xnor U40648 (N_40648,N_32232,N_37152);
nor U40649 (N_40649,N_34955,N_33049);
xnor U40650 (N_40650,N_39518,N_31506);
nand U40651 (N_40651,N_30566,N_35914);
or U40652 (N_40652,N_31972,N_34511);
nand U40653 (N_40653,N_39635,N_35384);
or U40654 (N_40654,N_39693,N_35048);
xor U40655 (N_40655,N_37237,N_37262);
and U40656 (N_40656,N_36014,N_32782);
or U40657 (N_40657,N_31076,N_31296);
nor U40658 (N_40658,N_32087,N_30822);
xnor U40659 (N_40659,N_30469,N_35335);
and U40660 (N_40660,N_35671,N_34354);
and U40661 (N_40661,N_36179,N_32435);
and U40662 (N_40662,N_38005,N_39651);
xnor U40663 (N_40663,N_31511,N_33148);
and U40664 (N_40664,N_30851,N_37439);
or U40665 (N_40665,N_34123,N_31340);
and U40666 (N_40666,N_32927,N_35078);
xor U40667 (N_40667,N_30219,N_31304);
or U40668 (N_40668,N_38436,N_34487);
and U40669 (N_40669,N_38864,N_32410);
or U40670 (N_40670,N_39634,N_39105);
nand U40671 (N_40671,N_39691,N_38567);
nand U40672 (N_40672,N_32722,N_39906);
or U40673 (N_40673,N_36027,N_33000);
nand U40674 (N_40674,N_34119,N_39829);
xnor U40675 (N_40675,N_38956,N_35205);
xnor U40676 (N_40676,N_35590,N_38062);
nor U40677 (N_40677,N_31977,N_32598);
or U40678 (N_40678,N_39463,N_32658);
xnor U40679 (N_40679,N_35543,N_30879);
or U40680 (N_40680,N_32736,N_35702);
and U40681 (N_40681,N_34605,N_31174);
nor U40682 (N_40682,N_37339,N_37726);
or U40683 (N_40683,N_33535,N_37246);
or U40684 (N_40684,N_33814,N_35157);
or U40685 (N_40685,N_31308,N_31643);
nor U40686 (N_40686,N_34207,N_32765);
or U40687 (N_40687,N_35792,N_37027);
xnor U40688 (N_40688,N_35003,N_39703);
or U40689 (N_40689,N_39813,N_34895);
and U40690 (N_40690,N_33543,N_30023);
or U40691 (N_40691,N_32870,N_36543);
and U40692 (N_40692,N_38330,N_36301);
or U40693 (N_40693,N_34262,N_35331);
nand U40694 (N_40694,N_34321,N_35116);
and U40695 (N_40695,N_34792,N_33089);
nor U40696 (N_40696,N_33269,N_34810);
nand U40697 (N_40697,N_33772,N_32542);
nor U40698 (N_40698,N_39268,N_31056);
nor U40699 (N_40699,N_32349,N_30218);
or U40700 (N_40700,N_31714,N_33478);
xnor U40701 (N_40701,N_36722,N_36539);
nor U40702 (N_40702,N_37138,N_36958);
or U40703 (N_40703,N_33915,N_35023);
nor U40704 (N_40704,N_35882,N_38407);
nand U40705 (N_40705,N_32888,N_33644);
or U40706 (N_40706,N_32810,N_36663);
nand U40707 (N_40707,N_35509,N_33097);
nor U40708 (N_40708,N_32069,N_30555);
nor U40709 (N_40709,N_31886,N_34737);
and U40710 (N_40710,N_37941,N_33425);
or U40711 (N_40711,N_39877,N_34802);
xnor U40712 (N_40712,N_32287,N_34135);
nor U40713 (N_40713,N_39308,N_30910);
and U40714 (N_40714,N_39128,N_35951);
xor U40715 (N_40715,N_32238,N_36114);
or U40716 (N_40716,N_37938,N_30886);
xnor U40717 (N_40717,N_39398,N_38450);
nor U40718 (N_40718,N_30171,N_30212);
xnor U40719 (N_40719,N_35847,N_33105);
and U40720 (N_40720,N_30854,N_31196);
nand U40721 (N_40721,N_35935,N_38511);
nor U40722 (N_40722,N_39527,N_35836);
nor U40723 (N_40723,N_35002,N_36182);
or U40724 (N_40724,N_32303,N_36887);
or U40725 (N_40725,N_37389,N_31190);
and U40726 (N_40726,N_30553,N_39907);
xor U40727 (N_40727,N_30900,N_31504);
nor U40728 (N_40728,N_33895,N_35278);
xor U40729 (N_40729,N_38029,N_38748);
xor U40730 (N_40730,N_38160,N_32488);
or U40731 (N_40731,N_39746,N_31620);
nand U40732 (N_40732,N_39875,N_30451);
xor U40733 (N_40733,N_36305,N_36508);
nand U40734 (N_40734,N_37531,N_39895);
or U40735 (N_40735,N_33226,N_36145);
xnor U40736 (N_40736,N_34360,N_35108);
nor U40737 (N_40737,N_30627,N_35743);
or U40738 (N_40738,N_39448,N_37554);
xor U40739 (N_40739,N_39773,N_38593);
or U40740 (N_40740,N_31246,N_36059);
xnor U40741 (N_40741,N_37984,N_31064);
nor U40742 (N_40742,N_30222,N_39771);
nor U40743 (N_40743,N_34350,N_30310);
or U40744 (N_40744,N_31050,N_34501);
or U40745 (N_40745,N_36853,N_38169);
nor U40746 (N_40746,N_30633,N_33473);
nand U40747 (N_40747,N_36472,N_33294);
nand U40748 (N_40748,N_39112,N_38997);
xor U40749 (N_40749,N_36158,N_38939);
or U40750 (N_40750,N_38285,N_30452);
nand U40751 (N_40751,N_32351,N_32195);
nor U40752 (N_40752,N_32996,N_36918);
xor U40753 (N_40753,N_31348,N_33726);
nand U40754 (N_40754,N_37710,N_34750);
and U40755 (N_40755,N_31574,N_38523);
or U40756 (N_40756,N_33459,N_38761);
xnor U40757 (N_40757,N_33894,N_31345);
xnor U40758 (N_40758,N_38758,N_31350);
or U40759 (N_40759,N_33838,N_30407);
nand U40760 (N_40760,N_37263,N_35016);
or U40761 (N_40761,N_33299,N_35338);
nand U40762 (N_40762,N_31016,N_30118);
and U40763 (N_40763,N_31702,N_33669);
and U40764 (N_40764,N_31335,N_32091);
and U40765 (N_40765,N_39256,N_30331);
and U40766 (N_40766,N_30104,N_35982);
nor U40767 (N_40767,N_31478,N_32356);
nand U40768 (N_40768,N_38730,N_30631);
nand U40769 (N_40769,N_37335,N_39545);
nor U40770 (N_40770,N_32216,N_34138);
xnor U40771 (N_40771,N_39243,N_38637);
or U40772 (N_40772,N_36265,N_35019);
nor U40773 (N_40773,N_35615,N_36956);
nand U40774 (N_40774,N_33980,N_31233);
and U40775 (N_40775,N_39062,N_39810);
nand U40776 (N_40776,N_31263,N_38928);
and U40777 (N_40777,N_31870,N_37253);
and U40778 (N_40778,N_30667,N_39638);
xor U40779 (N_40779,N_38822,N_32991);
and U40780 (N_40780,N_36760,N_39993);
nand U40781 (N_40781,N_32004,N_31287);
xnor U40782 (N_40782,N_36419,N_31618);
and U40783 (N_40783,N_36542,N_32389);
nor U40784 (N_40784,N_33645,N_37295);
nand U40785 (N_40785,N_37098,N_37782);
xor U40786 (N_40786,N_37973,N_32513);
nor U40787 (N_40787,N_36818,N_33070);
xnor U40788 (N_40788,N_32044,N_36569);
xor U40789 (N_40789,N_37080,N_39838);
or U40790 (N_40790,N_37149,N_32043);
or U40791 (N_40791,N_31208,N_38969);
or U40792 (N_40792,N_35328,N_39736);
or U40793 (N_40793,N_33334,N_30308);
nor U40794 (N_40794,N_34185,N_33180);
or U40795 (N_40795,N_32914,N_39523);
xnor U40796 (N_40796,N_34157,N_39260);
nand U40797 (N_40797,N_33969,N_38829);
nor U40798 (N_40798,N_37536,N_33796);
xnor U40799 (N_40799,N_33701,N_39093);
or U40800 (N_40800,N_38972,N_39734);
nand U40801 (N_40801,N_37963,N_36439);
nor U40802 (N_40802,N_36136,N_31199);
nand U40803 (N_40803,N_35834,N_32829);
and U40804 (N_40804,N_30110,N_31512);
or U40805 (N_40805,N_38826,N_35353);
or U40806 (N_40806,N_34025,N_31494);
or U40807 (N_40807,N_36063,N_32780);
xor U40808 (N_40808,N_38158,N_31734);
nand U40809 (N_40809,N_30658,N_34659);
nor U40810 (N_40810,N_38150,N_33001);
xnor U40811 (N_40811,N_33354,N_31678);
and U40812 (N_40812,N_34175,N_37398);
xnor U40813 (N_40813,N_39639,N_34149);
nor U40814 (N_40814,N_37825,N_35782);
nand U40815 (N_40815,N_35454,N_36729);
nand U40816 (N_40816,N_37579,N_37649);
xnor U40817 (N_40817,N_39599,N_37653);
nor U40818 (N_40818,N_34328,N_38427);
xnor U40819 (N_40819,N_34137,N_36612);
xor U40820 (N_40820,N_38027,N_34195);
or U40821 (N_40821,N_30641,N_31430);
or U40822 (N_40822,N_36263,N_37925);
xnor U40823 (N_40823,N_35984,N_35940);
xnor U40824 (N_40824,N_33057,N_32436);
or U40825 (N_40825,N_32999,N_34326);
xnor U40826 (N_40826,N_39040,N_33530);
and U40827 (N_40827,N_32092,N_35044);
and U40828 (N_40828,N_37567,N_33435);
or U40829 (N_40829,N_36358,N_36548);
nand U40830 (N_40830,N_32253,N_39751);
xnor U40831 (N_40831,N_30424,N_34692);
xnor U40832 (N_40832,N_36094,N_30916);
xnor U40833 (N_40833,N_33081,N_32824);
or U40834 (N_40834,N_32401,N_35129);
or U40835 (N_40835,N_32324,N_39899);
nand U40836 (N_40836,N_34448,N_30654);
nand U40837 (N_40837,N_37615,N_32822);
nand U40838 (N_40838,N_30720,N_35456);
and U40839 (N_40839,N_36401,N_31630);
or U40840 (N_40840,N_39711,N_31840);
nor U40841 (N_40841,N_39916,N_34208);
or U40842 (N_40842,N_36469,N_35681);
or U40843 (N_40843,N_38237,N_38846);
xnor U40844 (N_40844,N_39748,N_39129);
and U40845 (N_40845,N_33056,N_34519);
nor U40846 (N_40846,N_39869,N_35017);
xor U40847 (N_40847,N_37561,N_34858);
xor U40848 (N_40848,N_34642,N_38257);
nor U40849 (N_40849,N_30923,N_34950);
nor U40850 (N_40850,N_33684,N_33519);
nor U40851 (N_40851,N_32749,N_38663);
nor U40852 (N_40852,N_36683,N_33945);
xor U40853 (N_40853,N_35211,N_38938);
and U40854 (N_40854,N_35551,N_30825);
and U40855 (N_40855,N_31735,N_38832);
nor U40856 (N_40856,N_39412,N_36932);
or U40857 (N_40857,N_34726,N_39324);
or U40858 (N_40858,N_33207,N_36091);
nand U40859 (N_40859,N_31970,N_30857);
and U40860 (N_40860,N_31535,N_38415);
nor U40861 (N_40861,N_38191,N_30788);
and U40862 (N_40862,N_39715,N_37424);
nor U40863 (N_40863,N_38851,N_36254);
nor U40864 (N_40864,N_33889,N_37697);
nand U40865 (N_40865,N_33725,N_37001);
nand U40866 (N_40866,N_37819,N_30843);
and U40867 (N_40867,N_37677,N_37771);
or U40868 (N_40868,N_37127,N_30688);
nor U40869 (N_40869,N_39621,N_37522);
xnor U40870 (N_40870,N_34566,N_33874);
or U40871 (N_40871,N_38332,N_37245);
nor U40872 (N_40872,N_38173,N_35359);
xnor U40873 (N_40873,N_39253,N_32573);
nand U40874 (N_40874,N_30334,N_39491);
nand U40875 (N_40875,N_36892,N_30180);
nand U40876 (N_40876,N_31225,N_39148);
xnor U40877 (N_40877,N_39086,N_32441);
nor U40878 (N_40878,N_34213,N_36487);
xnor U40879 (N_40879,N_37861,N_32946);
nor U40880 (N_40880,N_39265,N_33003);
or U40881 (N_40881,N_38859,N_37377);
or U40882 (N_40882,N_39335,N_30903);
xor U40883 (N_40883,N_33171,N_35199);
xnor U40884 (N_40884,N_31433,N_30117);
nor U40885 (N_40885,N_38336,N_35114);
and U40886 (N_40886,N_33471,N_32963);
nor U40887 (N_40887,N_37914,N_39632);
nor U40888 (N_40888,N_30671,N_39598);
xor U40889 (N_40889,N_33355,N_37866);
xnor U40890 (N_40890,N_37330,N_36698);
or U40891 (N_40891,N_39493,N_34972);
and U40892 (N_40892,N_38982,N_31607);
and U40893 (N_40893,N_36620,N_31458);
or U40894 (N_40894,N_38109,N_38698);
and U40895 (N_40895,N_36836,N_32088);
xor U40896 (N_40896,N_37608,N_32710);
nand U40897 (N_40897,N_37057,N_34263);
and U40898 (N_40898,N_38664,N_38437);
nand U40899 (N_40899,N_37006,N_38206);
xnor U40900 (N_40900,N_35649,N_33593);
nor U40901 (N_40901,N_32570,N_33541);
nor U40902 (N_40902,N_31479,N_37995);
xnor U40903 (N_40903,N_35651,N_36532);
nand U40904 (N_40904,N_37547,N_33850);
nor U40905 (N_40905,N_30132,N_37597);
and U40906 (N_40906,N_31352,N_32229);
and U40907 (N_40907,N_34146,N_30225);
nor U40908 (N_40908,N_34275,N_37373);
nor U40909 (N_40909,N_30895,N_35912);
xnor U40910 (N_40910,N_36211,N_31222);
and U40911 (N_40911,N_32258,N_38420);
nor U40912 (N_40912,N_39973,N_38573);
xor U40913 (N_40913,N_34384,N_35076);
and U40914 (N_40914,N_38616,N_33920);
or U40915 (N_40915,N_32015,N_31446);
and U40916 (N_40916,N_38760,N_35186);
nor U40917 (N_40917,N_39310,N_38845);
or U40918 (N_40918,N_32508,N_37704);
xnor U40919 (N_40919,N_33599,N_33989);
or U40920 (N_40920,N_36288,N_33321);
or U40921 (N_40921,N_34427,N_34560);
and U40922 (N_40922,N_35430,N_36601);
nand U40923 (N_40923,N_30199,N_36445);
nor U40924 (N_40924,N_39910,N_37259);
nand U40925 (N_40925,N_32163,N_39779);
nor U40926 (N_40926,N_32913,N_32344);
and U40927 (N_40927,N_37415,N_31342);
or U40928 (N_40928,N_39223,N_31483);
xnor U40929 (N_40929,N_39990,N_38410);
nand U40930 (N_40930,N_31598,N_37142);
nor U40931 (N_40931,N_34807,N_37686);
and U40932 (N_40932,N_38918,N_39167);
and U40933 (N_40933,N_33329,N_31927);
nor U40934 (N_40934,N_35619,N_36999);
and U40935 (N_40935,N_33546,N_35213);
or U40936 (N_40936,N_31541,N_33388);
or U40937 (N_40937,N_32214,N_37665);
nor U40938 (N_40938,N_38755,N_33789);
and U40939 (N_40939,N_34046,N_34731);
nand U40940 (N_40940,N_34716,N_36277);
xnor U40941 (N_40941,N_38454,N_32239);
or U40942 (N_40942,N_39331,N_31391);
nand U40943 (N_40943,N_36504,N_36907);
nor U40944 (N_40944,N_30228,N_37899);
nor U40945 (N_40945,N_35204,N_31872);
and U40946 (N_40946,N_32032,N_32531);
or U40947 (N_40947,N_33587,N_39903);
or U40948 (N_40948,N_32318,N_36050);
nand U40949 (N_40949,N_38098,N_35999);
and U40950 (N_40950,N_37663,N_32923);
or U40951 (N_40951,N_36676,N_34547);
and U40952 (N_40952,N_33859,N_32153);
nand U40953 (N_40953,N_36963,N_32424);
nor U40954 (N_40954,N_31492,N_36882);
or U40955 (N_40955,N_36156,N_35262);
nand U40956 (N_40956,N_35122,N_31123);
xnor U40957 (N_40957,N_39078,N_33836);
and U40958 (N_40958,N_36925,N_31165);
nor U40959 (N_40959,N_38976,N_35011);
xnor U40960 (N_40960,N_31124,N_32286);
nand U40961 (N_40961,N_39498,N_38863);
nand U40962 (N_40962,N_38661,N_38187);
xnor U40963 (N_40963,N_35207,N_36515);
xnor U40964 (N_40964,N_32929,N_31641);
nand U40965 (N_40965,N_37915,N_37301);
xor U40966 (N_40966,N_38935,N_31120);
and U40967 (N_40967,N_36337,N_34074);
or U40968 (N_40968,N_36122,N_31657);
xor U40969 (N_40969,N_30478,N_36785);
xor U40970 (N_40970,N_39567,N_35714);
xor U40971 (N_40971,N_37940,N_36957);
nand U40972 (N_40972,N_36331,N_34818);
nand U40973 (N_40973,N_35307,N_33844);
or U40974 (N_40974,N_31386,N_30735);
xnor U40975 (N_40975,N_31201,N_39124);
nand U40976 (N_40976,N_36429,N_32285);
nand U40977 (N_40977,N_38815,N_37362);
xnor U40978 (N_40978,N_32816,N_37753);
nand U40979 (N_40979,N_39336,N_37331);
nor U40980 (N_40980,N_30652,N_39969);
nand U40981 (N_40981,N_31045,N_31300);
nand U40982 (N_40982,N_32089,N_38499);
or U40983 (N_40983,N_37592,N_32973);
nor U40984 (N_40984,N_31978,N_33483);
nand U40985 (N_40985,N_35309,N_31132);
xnor U40986 (N_40986,N_32859,N_31912);
or U40987 (N_40987,N_39483,N_39974);
xor U40988 (N_40988,N_34889,N_32662);
and U40989 (N_40989,N_38435,N_33339);
nor U40990 (N_40990,N_32906,N_35618);
or U40991 (N_40991,N_34842,N_31971);
xor U40992 (N_40992,N_31459,N_32426);
nand U40993 (N_40993,N_34217,N_36704);
and U40994 (N_40994,N_32376,N_36987);
nand U40995 (N_40995,N_33536,N_37338);
or U40996 (N_40996,N_38966,N_33775);
nor U40997 (N_40997,N_35519,N_30335);
xnor U40998 (N_40998,N_32235,N_31877);
xor U40999 (N_40999,N_37737,N_33311);
and U41000 (N_41000,N_32955,N_32081);
xor U41001 (N_41001,N_37774,N_38880);
or U41002 (N_41002,N_34339,N_39631);
nand U41003 (N_41003,N_38486,N_39985);
nand U41004 (N_41004,N_33456,N_32509);
or U41005 (N_41005,N_36875,N_35877);
or U41006 (N_41006,N_33693,N_39697);
or U41007 (N_41007,N_32943,N_33322);
nor U41008 (N_41008,N_30124,N_33197);
and U41009 (N_41009,N_35154,N_33181);
nor U41010 (N_41010,N_34580,N_33611);
nor U41011 (N_41011,N_37227,N_30955);
nor U41012 (N_41012,N_30699,N_39104);
xor U41013 (N_41013,N_34191,N_39798);
xor U41014 (N_41014,N_38116,N_33112);
and U41015 (N_41015,N_33565,N_38975);
nand U41016 (N_41016,N_34678,N_37865);
nor U41017 (N_41017,N_32528,N_37319);
nor U41018 (N_41018,N_35458,N_34247);
nand U41019 (N_41019,N_39247,N_36148);
nor U41020 (N_41020,N_31792,N_32304);
nand U41021 (N_41021,N_37636,N_36903);
nor U41022 (N_41022,N_37766,N_37675);
xor U41023 (N_41023,N_31680,N_35747);
xor U41024 (N_41024,N_30898,N_33014);
xor U41025 (N_41025,N_37967,N_34658);
xnor U41026 (N_41026,N_38290,N_39660);
or U41027 (N_41027,N_39326,N_37247);
nand U41028 (N_41028,N_32587,N_37931);
nor U41029 (N_41029,N_36035,N_33807);
xnor U41030 (N_41030,N_30738,N_37904);
nand U41031 (N_41031,N_35853,N_34581);
nand U41032 (N_41032,N_36013,N_35126);
xnor U41033 (N_41033,N_38780,N_33635);
and U41034 (N_41034,N_30806,N_33128);
or U41035 (N_41035,N_38112,N_30173);
xnor U41036 (N_41036,N_39111,N_36292);
nand U41037 (N_41037,N_38904,N_30677);
nand U41038 (N_41038,N_34324,N_37375);
nor U41039 (N_41039,N_32209,N_39700);
nand U41040 (N_41040,N_35260,N_36339);
or U41041 (N_41041,N_30924,N_39309);
or U41042 (N_41042,N_36368,N_31515);
nor U41043 (N_41043,N_38585,N_38463);
and U41044 (N_41044,N_39529,N_32159);
or U41045 (N_41045,N_31996,N_38025);
nand U41046 (N_41046,N_31258,N_37876);
or U41047 (N_41047,N_37702,N_30618);
and U41048 (N_41048,N_30685,N_31788);
and U41049 (N_41049,N_37871,N_32133);
or U41050 (N_41050,N_35986,N_31760);
nor U41051 (N_41051,N_33711,N_39055);
or U41052 (N_41052,N_34718,N_31732);
and U41053 (N_41053,N_32901,N_38868);
nor U41054 (N_41054,N_32851,N_37033);
or U41055 (N_41055,N_38701,N_39889);
nand U41056 (N_41056,N_34155,N_31347);
nand U41057 (N_41057,N_31316,N_30858);
nand U41058 (N_41058,N_32657,N_32500);
or U41059 (N_41059,N_38022,N_38558);
and U41060 (N_41060,N_34827,N_34199);
nor U41061 (N_41061,N_34704,N_35511);
xor U41062 (N_41062,N_31014,N_36245);
nand U41063 (N_41063,N_38241,N_39383);
nand U41064 (N_41064,N_35838,N_32129);
and U41065 (N_41065,N_30957,N_36194);
and U41066 (N_41066,N_36309,N_33042);
and U41067 (N_41067,N_33434,N_30592);
and U41068 (N_41068,N_37604,N_34334);
nor U41069 (N_41069,N_39640,N_32863);
xnor U41070 (N_41070,N_34924,N_32550);
and U41071 (N_41071,N_34319,N_39556);
and U41072 (N_41072,N_30312,N_32493);
nand U41073 (N_41073,N_37360,N_33673);
nor U41074 (N_41074,N_37776,N_38553);
nand U41075 (N_41075,N_37968,N_37289);
nand U41076 (N_41076,N_32268,N_38376);
nor U41077 (N_41077,N_39034,N_33675);
nor U41078 (N_41078,N_35408,N_36686);
xor U41079 (N_41079,N_30832,N_32619);
and U41080 (N_41080,N_33308,N_35925);
nand U41081 (N_41081,N_36522,N_38194);
and U41082 (N_41082,N_32123,N_36592);
xor U41083 (N_41083,N_33882,N_30406);
and U41084 (N_41084,N_33177,N_39848);
nor U41085 (N_41085,N_38494,N_31107);
nand U41086 (N_41086,N_32594,N_36139);
xor U41087 (N_41087,N_31797,N_34452);
and U41088 (N_41088,N_34625,N_33208);
xor U41089 (N_41089,N_39301,N_30508);
nor U41090 (N_41090,N_36626,N_31826);
xnor U41091 (N_41091,N_30665,N_31404);
nor U41092 (N_41092,N_35758,N_39946);
xor U41093 (N_41093,N_36499,N_31198);
or U41094 (N_41094,N_34398,N_32902);
xor U41095 (N_41095,N_37328,N_35598);
nand U41096 (N_41096,N_39707,N_34970);
nand U41097 (N_41097,N_37336,N_35371);
nand U41098 (N_41098,N_38977,N_39311);
and U41099 (N_41099,N_38329,N_35915);
and U41100 (N_41100,N_35664,N_37092);
nor U41101 (N_41101,N_33640,N_32799);
nor U41102 (N_41102,N_35352,N_32397);
or U41103 (N_41103,N_35327,N_34465);
nand U41104 (N_41104,N_31528,N_36938);
or U41105 (N_41105,N_30899,N_33741);
and U41106 (N_41106,N_30758,N_35460);
or U41107 (N_41107,N_32473,N_36900);
nand U41108 (N_41108,N_33237,N_38422);
nand U41109 (N_41109,N_30145,N_36777);
and U41110 (N_41110,N_39982,N_37750);
xor U41111 (N_41111,N_32348,N_33988);
xnor U41112 (N_41112,N_37313,N_34615);
xnor U41113 (N_41113,N_39384,N_34181);
or U41114 (N_41114,N_35521,N_30601);
nand U41115 (N_41115,N_37979,N_36744);
nor U41116 (N_41116,N_34064,N_33211);
nor U41117 (N_41117,N_37633,N_39789);
or U41118 (N_41118,N_30799,N_34098);
and U41119 (N_41119,N_34069,N_33508);
and U41120 (N_41120,N_37684,N_30257);
nor U41121 (N_41121,N_39283,N_33942);
nor U41122 (N_41122,N_32438,N_33791);
or U41123 (N_41123,N_32310,N_30979);
nor U41124 (N_41124,N_33114,N_37489);
nor U41125 (N_41125,N_33275,N_35357);
and U41126 (N_41126,N_38643,N_30289);
and U41127 (N_41127,N_39817,N_34994);
or U41128 (N_41128,N_37545,N_39922);
or U41129 (N_41129,N_37242,N_35074);
nand U41130 (N_41130,N_33904,N_34396);
and U41131 (N_41131,N_35778,N_30930);
xnor U41132 (N_41132,N_36066,N_35139);
and U41133 (N_41133,N_32012,N_36714);
xnor U41134 (N_41134,N_35452,N_37125);
xnor U41135 (N_41135,N_39438,N_35461);
or U41136 (N_41136,N_33949,N_34115);
and U41137 (N_41137,N_39271,N_36005);
xor U41138 (N_41138,N_31676,N_39343);
and U41139 (N_41139,N_39921,N_33494);
xor U41140 (N_41140,N_37506,N_31563);
or U41141 (N_41141,N_31846,N_30309);
or U41142 (N_41142,N_31273,N_32010);
or U41143 (N_41143,N_30466,N_36356);
or U41144 (N_41144,N_30829,N_36086);
or U41145 (N_41145,N_33578,N_38298);
xor U41146 (N_41146,N_38878,N_34559);
nand U41147 (N_41147,N_34047,N_39620);
nand U41148 (N_41148,N_37220,N_30714);
or U41149 (N_41149,N_31360,N_39061);
xnor U41150 (N_41150,N_34315,N_38517);
nand U41151 (N_41151,N_32800,N_37432);
and U41152 (N_41152,N_35229,N_31552);
or U41153 (N_41153,N_31808,N_30084);
or U41154 (N_41154,N_38653,N_39214);
and U41155 (N_41155,N_30623,N_31411);
nor U41156 (N_41156,N_31693,N_31272);
or U41157 (N_41157,N_30234,N_30045);
or U41158 (N_41158,N_35700,N_32248);
xor U41159 (N_41159,N_38313,N_35070);
nor U41160 (N_41160,N_31943,N_37945);
and U41161 (N_41161,N_39678,N_34522);
nor U41162 (N_41162,N_31095,N_37451);
nand U41163 (N_41163,N_38789,N_32028);
xnor U41164 (N_41164,N_31991,N_38806);
and U41165 (N_41165,N_38842,N_39263);
nand U41166 (N_41166,N_37349,N_32965);
or U41167 (N_41167,N_38060,N_31001);
and U41168 (N_41168,N_38835,N_39018);
or U41169 (N_41169,N_30931,N_34148);
nor U41170 (N_41170,N_31204,N_34916);
or U41171 (N_41171,N_35795,N_32218);
nand U41172 (N_41172,N_38706,N_32053);
xor U41173 (N_41173,N_37443,N_31406);
xor U41174 (N_41174,N_38119,N_32855);
or U41175 (N_41175,N_36413,N_38768);
xor U41176 (N_41176,N_38912,N_38253);
nand U41177 (N_41177,N_38460,N_30941);
nand U41178 (N_41178,N_38466,N_31945);
xor U41179 (N_41179,N_37387,N_36343);
and U41180 (N_41180,N_30701,N_35582);
xor U41181 (N_41181,N_32170,N_36041);
xor U41182 (N_41182,N_39688,N_35913);
nand U41183 (N_41183,N_35585,N_35228);
nor U41184 (N_41184,N_38149,N_32687);
nor U41185 (N_41185,N_30231,N_35719);
nand U41186 (N_41186,N_32808,N_39262);
xor U41187 (N_41187,N_33417,N_35779);
xor U41188 (N_41188,N_32072,N_39512);
and U41189 (N_41189,N_30409,N_34980);
nor U41190 (N_41190,N_39563,N_32893);
nand U41191 (N_41191,N_37912,N_31814);
nand U41192 (N_41192,N_33301,N_39106);
or U41193 (N_41193,N_37671,N_37526);
or U41194 (N_41194,N_31102,N_30636);
nor U41195 (N_41195,N_39360,N_36863);
nand U41196 (N_41196,N_33993,N_35012);
nand U41197 (N_41197,N_33251,N_31418);
nand U41198 (N_41198,N_32003,N_36610);
xnor U41199 (N_41199,N_31428,N_30554);
xnor U41200 (N_41200,N_39205,N_35890);
and U41201 (N_41201,N_39051,N_35690);
nand U41202 (N_41202,N_31058,N_32621);
nor U41203 (N_41203,N_33196,N_35884);
xor U41204 (N_41204,N_33041,N_32155);
or U41205 (N_41205,N_32697,N_30426);
and U41206 (N_41206,N_34494,N_38537);
xnor U41207 (N_41207,N_30584,N_37345);
nand U41208 (N_41208,N_33880,N_34214);
nor U41209 (N_41209,N_34528,N_37975);
and U41210 (N_41210,N_38345,N_39446);
xor U41211 (N_41211,N_32084,N_31903);
or U41212 (N_41212,N_38295,N_35009);
xor U41213 (N_41213,N_32933,N_32846);
or U41214 (N_41214,N_39327,N_32097);
and U41215 (N_41215,N_36944,N_31662);
and U41216 (N_41216,N_32365,N_33009);
nor U41217 (N_41217,N_33655,N_39902);
nand U41218 (N_41218,N_39027,N_32322);
xor U41219 (N_41219,N_34355,N_36240);
and U41220 (N_41220,N_31162,N_34144);
xnor U41221 (N_41221,N_33499,N_31312);
and U41222 (N_41222,N_39482,N_38816);
nor U41223 (N_41223,N_32795,N_34773);
xor U41224 (N_41224,N_37321,N_37958);
xor U41225 (N_41225,N_37447,N_33658);
nand U41226 (N_41226,N_32423,N_33512);
xor U41227 (N_41227,N_34437,N_39045);
nor U41228 (N_41228,N_32444,N_34357);
and U41229 (N_41229,N_35159,N_30991);
xor U41230 (N_41230,N_39274,N_37707);
and U41231 (N_41231,N_39019,N_31203);
nand U41232 (N_41232,N_32115,N_34848);
nor U41233 (N_41233,N_31065,N_35980);
xor U41234 (N_41234,N_37168,N_32468);
xor U41235 (N_41235,N_30266,N_33195);
and U41236 (N_41236,N_31849,N_37038);
nor U41237 (N_41237,N_30669,N_33970);
or U41238 (N_41238,N_32980,N_32600);
and U41239 (N_41239,N_36484,N_30412);
nor U41240 (N_41240,N_32681,N_38235);
nand U41241 (N_41241,N_31942,N_31786);
nor U41242 (N_41242,N_39307,N_32312);
or U41243 (N_41243,N_39912,N_35663);
or U41244 (N_41244,N_34524,N_30049);
and U41245 (N_41245,N_33274,N_33912);
nand U41246 (N_41246,N_31999,N_32392);
nand U41247 (N_41247,N_37474,N_38380);
nor U41248 (N_41248,N_32812,N_34169);
nand U41249 (N_41249,N_34000,N_35976);
and U41250 (N_41250,N_37378,N_38473);
nor U41251 (N_41251,N_33330,N_32690);
or U41252 (N_41252,N_38425,N_32107);
nor U41253 (N_41253,N_34444,N_31025);
nor U41254 (N_41254,N_35220,N_33856);
nor U41255 (N_41255,N_38714,N_37955);
or U41256 (N_41256,N_34541,N_34548);
xnor U41257 (N_41257,N_39672,N_34570);
nor U41258 (N_41258,N_34335,N_38656);
nor U41259 (N_41259,N_30765,N_30044);
xor U41260 (N_41260,N_30534,N_32485);
nor U41261 (N_41261,N_32013,N_31665);
or U41262 (N_41262,N_31930,N_37721);
nor U41263 (N_41263,N_31759,N_33409);
nor U41264 (N_41264,N_30821,N_34071);
and U41265 (N_41265,N_37923,N_36618);
nand U41266 (N_41266,N_38536,N_30095);
and U41267 (N_41267,N_32000,N_39847);
nand U41268 (N_41268,N_36447,N_35640);
and U41269 (N_41269,N_36384,N_36362);
and U41270 (N_41270,N_31987,N_37258);
nand U41271 (N_41271,N_32210,N_35189);
xnor U41272 (N_41272,N_36079,N_35657);
nand U41273 (N_41273,N_32762,N_37048);
and U41274 (N_41274,N_35409,N_36677);
xor U41275 (N_41275,N_34235,N_38651);
xor U41276 (N_41276,N_32203,N_37954);
or U41277 (N_41277,N_33522,N_39270);
or U41278 (N_41278,N_31269,N_35692);
nor U41279 (N_41279,N_34410,N_38848);
nand U41280 (N_41280,N_37610,N_38057);
xor U41281 (N_41281,N_39445,N_33926);
and U41282 (N_41282,N_33639,N_30217);
and U41283 (N_41283,N_39145,N_37395);
nor U41284 (N_41284,N_31292,N_32301);
and U41285 (N_41285,N_35623,N_34240);
or U41286 (N_41286,N_34241,N_36822);
and U41287 (N_41287,N_38197,N_32154);
nor U41288 (N_41288,N_34110,N_30522);
or U41289 (N_41289,N_39547,N_39080);
nor U41290 (N_41290,N_36326,N_34709);
nor U41291 (N_41291,N_30006,N_39981);
and U41292 (N_41292,N_33134,N_36185);
or U41293 (N_41293,N_35722,N_33931);
nor U41294 (N_41294,N_32592,N_32458);
and U41295 (N_41295,N_33348,N_35952);
and U41296 (N_41296,N_38598,N_34040);
and U41297 (N_41297,N_30789,N_36909);
nor U41298 (N_41298,N_31378,N_32270);
and U41299 (N_41299,N_33297,N_34561);
nand U41300 (N_41300,N_30022,N_32968);
xor U41301 (N_41301,N_33082,N_38279);
nand U41302 (N_41302,N_39332,N_36510);
xnor U41303 (N_41303,N_31899,N_32355);
xor U41304 (N_41304,N_31184,N_38551);
xor U41305 (N_41305,N_30587,N_39356);
or U41306 (N_41306,N_31370,N_37239);
and U41307 (N_41307,N_34774,N_32199);
or U41308 (N_41308,N_34962,N_39750);
xor U41309 (N_41309,N_36644,N_38932);
nand U41310 (N_41310,N_34651,N_32739);
or U41311 (N_41311,N_34056,N_32103);
and U41312 (N_41312,N_38431,N_34562);
and U41313 (N_41313,N_31317,N_39716);
or U41314 (N_41314,N_39068,N_37729);
xor U41315 (N_41315,N_31205,N_34830);
and U41316 (N_41316,N_36242,N_35196);
and U41317 (N_41317,N_39908,N_36424);
nand U41318 (N_41318,N_38610,N_38448);
nor U41319 (N_41319,N_30052,N_37068);
nand U41320 (N_41320,N_31328,N_35518);
nor U41321 (N_41321,N_30973,N_35273);
xnor U41322 (N_41322,N_35251,N_37651);
and U41323 (N_41323,N_39298,N_34629);
and U41324 (N_41324,N_37112,N_33757);
nor U41325 (N_41325,N_36795,N_31264);
xnor U41326 (N_41326,N_34526,N_36828);
and U41327 (N_41327,N_36536,N_38373);
nor U41328 (N_41328,N_33996,N_31481);
nor U41329 (N_41329,N_37367,N_34424);
xor U41330 (N_41330,N_35382,N_33864);
xnor U41331 (N_41331,N_35686,N_32082);
nand U41332 (N_41332,N_36666,N_37679);
and U41333 (N_41333,N_36641,N_30323);
nand U41334 (N_41334,N_30364,N_33935);
nand U41335 (N_41335,N_32696,N_37218);
xor U41336 (N_41336,N_39637,N_34205);
xor U41337 (N_41337,N_38888,N_36205);
and U41338 (N_41338,N_37145,N_37460);
or U41339 (N_41339,N_37419,N_39727);
nor U41340 (N_41340,N_36731,N_33300);
xnor U41341 (N_41341,N_38812,N_38950);
xor U41342 (N_41342,N_36690,N_38354);
and U41343 (N_41343,N_32319,N_33689);
and U41344 (N_41344,N_31249,N_39321);
or U41345 (N_41345,N_38404,N_32758);
or U41346 (N_41346,N_35534,N_38086);
nor U41347 (N_41347,N_32692,N_31551);
xnor U41348 (N_41348,N_31746,N_39940);
and U41349 (N_41349,N_36202,N_31424);
nor U41350 (N_41350,N_37490,N_36905);
xnor U41351 (N_41351,N_35459,N_37024);
nor U41352 (N_41352,N_38189,N_30020);
nor U41353 (N_41353,N_37366,N_32958);
and U41354 (N_41354,N_37388,N_33452);
xnor U41355 (N_41355,N_35737,N_36871);
xnor U41356 (N_41356,N_38171,N_35531);
xor U41357 (N_41357,N_38990,N_37751);
and U41358 (N_41358,N_38589,N_39541);
nand U41359 (N_41359,N_37534,N_34084);
xor U41360 (N_41360,N_38512,N_32796);
xor U41361 (N_41361,N_32771,N_33825);
nand U41362 (N_41362,N_37570,N_32459);
nor U41363 (N_41363,N_33162,N_36407);
nor U41364 (N_41364,N_37703,N_35628);
and U41365 (N_41365,N_31337,N_30287);
or U41366 (N_41366,N_31349,N_33045);
xor U41367 (N_41367,N_37756,N_35346);
and U41368 (N_41368,N_35385,N_39408);
nor U41369 (N_41369,N_35015,N_35223);
nor U41370 (N_41370,N_36979,N_32584);
nor U41371 (N_41371,N_31017,N_37268);
nor U41372 (N_41372,N_39488,N_32034);
nor U41373 (N_41373,N_34131,N_32924);
or U41374 (N_41374,N_37507,N_30745);
and U41375 (N_41375,N_31490,N_38032);
xnor U41376 (N_41376,N_36352,N_30085);
nand U41377 (N_41377,N_32884,N_38733);
or U41378 (N_41378,N_37907,N_34387);
and U41379 (N_41379,N_31452,N_39851);
xnor U41380 (N_41380,N_39012,N_32682);
or U41381 (N_41381,N_33680,N_37909);
and U41382 (N_41382,N_33423,N_38810);
nor U41383 (N_41383,N_35500,N_30972);
nor U41384 (N_41384,N_39765,N_38873);
nand U41385 (N_41385,N_35642,N_34385);
xnor U41386 (N_41386,N_35589,N_35840);
xnor U41387 (N_41387,N_33893,N_31832);
nand U41388 (N_41388,N_35865,N_34821);
nand U41389 (N_41389,N_39346,N_31231);
xor U41390 (N_41390,N_39091,N_36471);
xor U41391 (N_41391,N_32843,N_30718);
nand U41392 (N_41392,N_38011,N_38434);
nor U41393 (N_41393,N_35835,N_31994);
or U41394 (N_41394,N_32684,N_36369);
or U41395 (N_41395,N_34671,N_38402);
nor U41396 (N_41396,N_34282,N_39788);
and U41397 (N_41397,N_34670,N_33336);
and U41398 (N_41398,N_30950,N_37256);
or U41399 (N_41399,N_32090,N_31084);
or U41400 (N_41400,N_31683,N_32698);
nand U41401 (N_41401,N_36653,N_38038);
and U41402 (N_41402,N_37458,N_31152);
nor U41403 (N_41403,N_31654,N_33967);
and U41404 (N_41404,N_38654,N_31770);
and U41405 (N_41405,N_36363,N_35010);
nor U41406 (N_41406,N_32908,N_30838);
or U41407 (N_41407,N_30352,N_33395);
nor U41408 (N_41408,N_34636,N_31762);
xor U41409 (N_41409,N_33410,N_36308);
nor U41410 (N_41410,N_38860,N_36418);
nand U41411 (N_41411,N_38343,N_30280);
nor U41412 (N_41412,N_39237,N_36558);
and U41413 (N_41413,N_39839,N_33072);
or U41414 (N_41414,N_32202,N_32530);
nor U41415 (N_41415,N_30662,N_37985);
xor U41416 (N_41416,N_32490,N_31925);
nor U41417 (N_41417,N_30186,N_30642);
nand U41418 (N_41418,N_38601,N_38054);
nand U41419 (N_41419,N_35667,N_39654);
nor U41420 (N_41420,N_33443,N_33685);
nand U41421 (N_41421,N_31664,N_38294);
xor U41422 (N_41422,N_30581,N_38625);
and U41423 (N_41423,N_37135,N_36933);
or U41424 (N_41424,N_39568,N_33950);
nor U41425 (N_41425,N_33475,N_37182);
xnor U41426 (N_41426,N_32875,N_32885);
and U41427 (N_41427,N_39487,N_30447);
or U41428 (N_41428,N_30394,N_33712);
nand U41429 (N_41429,N_33773,N_34673);
xnor U41430 (N_41430,N_31061,N_37300);
nand U41431 (N_41431,N_34005,N_35583);
nor U41432 (N_41432,N_35817,N_34805);
and U41433 (N_41433,N_33985,N_30563);
nand U41434 (N_41434,N_30061,N_37074);
nand U41435 (N_41435,N_38273,N_31189);
nor U41436 (N_41436,N_37156,N_39218);
nor U41437 (N_41437,N_37107,N_36991);
nor U41438 (N_41438,N_36071,N_30025);
nor U41439 (N_41439,N_32694,N_35245);
or U41440 (N_41440,N_36912,N_31077);
nor U41441 (N_41441,N_38917,N_35381);
or U41442 (N_41442,N_32190,N_39960);
or U41443 (N_41443,N_31234,N_34975);
or U41444 (N_41444,N_32568,N_32022);
xor U41445 (N_41445,N_34695,N_35985);
nor U41446 (N_41446,N_38251,N_32295);
and U41447 (N_41447,N_38899,N_38250);
nand U41448 (N_41448,N_32745,N_36885);
nand U41449 (N_41449,N_36168,N_30517);
nor U41450 (N_41450,N_32457,N_32655);
and U41451 (N_41451,N_31964,N_35956);
nor U41452 (N_41452,N_31457,N_31085);
nand U41453 (N_41453,N_38270,N_30097);
and U41454 (N_41454,N_30828,N_35910);
nand U41455 (N_41455,N_31491,N_35685);
and U41456 (N_41456,N_37658,N_35495);
or U41457 (N_41457,N_37712,N_35850);
nor U41458 (N_41458,N_38229,N_32577);
or U41459 (N_41459,N_38955,N_35029);
or U41460 (N_41460,N_37399,N_30484);
xor U41461 (N_41461,N_37599,N_31380);
or U41462 (N_41462,N_38556,N_34878);
and U41463 (N_41463,N_36898,N_34956);
or U41464 (N_41464,N_38542,N_36341);
nor U41465 (N_41465,N_34910,N_32596);
and U41466 (N_41466,N_33010,N_35992);
or U41467 (N_41467,N_35033,N_33420);
xor U41468 (N_41468,N_37452,N_39033);
and U41469 (N_41469,N_32713,N_32916);
or U41470 (N_41470,N_31178,N_33526);
nand U41471 (N_41471,N_37150,N_39216);
or U41472 (N_41472,N_35948,N_31731);
xnor U41473 (N_41473,N_33732,N_34644);
and U41474 (N_41474,N_37509,N_33272);
or U41475 (N_41475,N_32784,N_38833);
or U41476 (N_41476,N_34902,N_35247);
nand U41477 (N_41477,N_30812,N_30932);
xor U41478 (N_41478,N_39415,N_39665);
nor U41479 (N_41479,N_37556,N_37678);
nor U41480 (N_41480,N_35319,N_36967);
and U41481 (N_41481,N_38849,N_31822);
xor U41482 (N_41482,N_39293,N_36489);
xnor U41483 (N_41483,N_37662,N_37919);
nor U41484 (N_41484,N_36685,N_36427);
xnor U41485 (N_41485,N_31336,N_39892);
nor U41486 (N_41486,N_33848,N_36886);
xor U41487 (N_41487,N_31247,N_36058);
nor U41488 (N_41488,N_37108,N_31667);
and U41489 (N_41489,N_37404,N_34854);
and U41490 (N_41490,N_30660,N_30670);
nand U41491 (N_41491,N_36553,N_39425);
nand U41492 (N_41492,N_36741,N_31096);
and U41493 (N_41493,N_31897,N_36208);
nand U41494 (N_41494,N_37163,N_38472);
and U41495 (N_41495,N_34881,N_37002);
nand U41496 (N_41496,N_36417,N_36649);
or U41497 (N_41497,N_38974,N_39159);
nor U41498 (N_41498,N_36980,N_38579);
nor U41499 (N_41499,N_34863,N_38937);
xor U41500 (N_41500,N_36270,N_36468);
or U41501 (N_41501,N_34338,N_39661);
nand U41502 (N_41502,N_34510,N_35739);
nand U41503 (N_41503,N_35942,N_36947);
xor U41504 (N_41504,N_39367,N_31842);
and U41505 (N_41505,N_34551,N_37176);
nor U41506 (N_41506,N_36978,N_30388);
xor U41507 (N_41507,N_33449,N_30716);
nand U41508 (N_41508,N_37497,N_37949);
nand U41509 (N_41509,N_38451,N_36910);
or U41510 (N_41510,N_35208,N_32430);
and U41511 (N_41511,N_33674,N_37616);
and U41512 (N_41512,N_39059,N_38782);
xnor U41513 (N_41513,N_34296,N_35301);
or U41514 (N_41514,N_39914,N_36952);
or U41515 (N_41515,N_35368,N_38286);
xor U41516 (N_41516,N_34602,N_34163);
nor U41517 (N_41517,N_38582,N_34229);
nor U41518 (N_41518,N_35202,N_39373);
or U41519 (N_41519,N_35567,N_38193);
and U41520 (N_41520,N_34738,N_38392);
xnor U41521 (N_41521,N_38021,N_36408);
or U41522 (N_41522,N_32194,N_31357);
nand U41523 (N_41523,N_33263,N_33930);
nor U41524 (N_41524,N_37960,N_31324);
or U41525 (N_41525,N_37071,N_34648);
nand U41526 (N_41526,N_38144,N_32386);
or U41527 (N_41527,N_32648,N_36530);
nand U41528 (N_41528,N_33380,N_30613);
nor U41529 (N_41529,N_35345,N_39233);
nand U41530 (N_41530,N_39063,N_30325);
or U41531 (N_41531,N_32417,N_33636);
or U41532 (N_41532,N_35034,N_38777);
nor U41533 (N_41533,N_35383,N_36486);
and U41534 (N_41534,N_39338,N_31602);
nand U41535 (N_41535,N_38979,N_39600);
nor U41536 (N_41536,N_38914,N_38168);
or U41537 (N_41537,N_36937,N_35955);
or U41538 (N_41538,N_31353,N_33192);
nand U41539 (N_41539,N_35947,N_34381);
nor U41540 (N_41540,N_39883,N_32080);
or U41541 (N_41541,N_35785,N_31810);
and U41542 (N_41542,N_31279,N_39975);
nor U41543 (N_41543,N_33115,N_39172);
xor U41544 (N_41544,N_35412,N_32360);
xnor U41545 (N_41545,N_36546,N_31963);
and U41546 (N_41546,N_32599,N_31829);
nor U41547 (N_41547,N_35620,N_36706);
and U41548 (N_41548,N_35377,N_32627);
or U41549 (N_41549,N_32217,N_36460);
nor U41550 (N_41550,N_31841,N_32860);
xnor U41551 (N_41551,N_35808,N_37180);
xor U41552 (N_41552,N_39375,N_36825);
or U41553 (N_41553,N_34043,N_38262);
nand U41554 (N_41554,N_39290,N_33690);
or U41555 (N_41555,N_34052,N_38640);
and U41556 (N_41556,N_39777,N_38691);
xnor U41557 (N_41557,N_32054,N_35055);
xor U41558 (N_41558,N_39372,N_39084);
nand U41559 (N_41559,N_35127,N_33183);
xnor U41560 (N_41560,N_34051,N_36633);
or U41561 (N_41561,N_30936,N_30259);
and U41562 (N_41562,N_34197,N_37622);
and U41563 (N_41563,N_33495,N_36518);
nor U41564 (N_41564,N_39185,N_33055);
xor U41565 (N_41565,N_31593,N_37342);
nand U41566 (N_41566,N_39350,N_36551);
nand U41567 (N_41567,N_37548,N_39996);
nor U41568 (N_41568,N_30400,N_30543);
or U41569 (N_41569,N_30464,N_34873);
xor U41570 (N_41570,N_37249,N_38107);
xor U41571 (N_41571,N_38614,N_32821);
nor U41572 (N_41572,N_35136,N_39003);
nand U41573 (N_41573,N_32899,N_36565);
or U41574 (N_41574,N_34186,N_36174);
nand U41575 (N_41575,N_32741,N_31626);
and U41576 (N_41576,N_32580,N_34798);
nor U41577 (N_41577,N_33375,N_32962);
xor U41578 (N_41578,N_34222,N_38587);
and U41579 (N_41579,N_35825,N_31692);
or U41580 (N_41580,N_33316,N_32047);
nor U41581 (N_41581,N_30150,N_35448);
nand U41582 (N_41582,N_38828,N_39786);
nor U41583 (N_41583,N_33069,N_37318);
and U41584 (N_41584,N_36187,N_32478);
or U41585 (N_41585,N_32730,N_38795);
and U41586 (N_41586,N_33928,N_31998);
and U41587 (N_41587,N_36577,N_36100);
xor U41588 (N_41588,N_33591,N_33465);
or U41589 (N_41589,N_39049,N_39083);
or U41590 (N_41590,N_35465,N_33509);
nor U41591 (N_41591,N_30258,N_35760);
xor U41592 (N_41592,N_33900,N_30723);
nor U41593 (N_41593,N_35605,N_33173);
nor U41594 (N_41594,N_38323,N_34281);
xnor U41595 (N_41595,N_39898,N_38752);
nor U41596 (N_41596,N_38161,N_36377);
or U41597 (N_41597,N_39841,N_32501);
xor U41598 (N_41598,N_32969,N_35934);
nor U41599 (N_41599,N_39760,N_35300);
nor U41600 (N_41600,N_37817,N_37343);
nand U41601 (N_41601,N_35763,N_31738);
or U41602 (N_41602,N_31718,N_31485);
xor U41603 (N_41603,N_32045,N_37718);
and U41604 (N_41604,N_37350,N_36068);
xor U41605 (N_41605,N_36019,N_38689);
or U41606 (N_41606,N_37966,N_36759);
xnor U41607 (N_41607,N_38562,N_34976);
and U41608 (N_41608,N_35604,N_30191);
nor U41609 (N_41609,N_35063,N_35789);
xnor U41610 (N_41610,N_32167,N_38403);
nand U41611 (N_41611,N_33160,N_32334);
xnor U41612 (N_41612,N_31556,N_35757);
nand U41613 (N_41613,N_34845,N_36074);
nand U41614 (N_41614,N_35376,N_35318);
and U41615 (N_41615,N_30392,N_30369);
and U41616 (N_41616,N_36839,N_31055);
xor U41617 (N_41617,N_39385,N_37412);
or U41618 (N_41618,N_39937,N_38428);
nand U41619 (N_41619,N_31956,N_32947);
xnor U41620 (N_41620,N_33528,N_37546);
xor U41621 (N_41621,N_36133,N_35918);
nor U41622 (N_41622,N_33679,N_37648);
nand U41623 (N_41623,N_37055,N_30026);
xnor U41624 (N_41624,N_36961,N_32566);
nand U41625 (N_41625,N_36090,N_35677);
nand U41626 (N_41626,N_32418,N_33924);
nand U41627 (N_41627,N_35356,N_38324);
nor U41628 (N_41628,N_33939,N_32121);
and U41629 (N_41629,N_34178,N_37503);
nor U41630 (N_41630,N_32098,N_35656);
nor U41631 (N_41631,N_33287,N_31802);
or U41632 (N_41632,N_36191,N_36689);
nand U41633 (N_41633,N_38040,N_32051);
nand U41634 (N_41634,N_37252,N_35858);
nor U41635 (N_41635,N_39410,N_35236);
nand U41636 (N_41636,N_34432,N_34171);
or U41637 (N_41637,N_31188,N_31071);
xnor U41638 (N_41638,N_34536,N_30664);
nor U41639 (N_41639,N_33476,N_33729);
nor U41640 (N_41640,N_33598,N_38137);
or U41641 (N_41641,N_38642,N_35054);
or U41642 (N_41642,N_34122,N_36072);
nand U41643 (N_41643,N_34026,N_37674);
and U41644 (N_41644,N_31008,N_33759);
or U41645 (N_41645,N_32109,N_33717);
nand U41646 (N_41646,N_35639,N_35486);
xnor U41647 (N_41647,N_36670,N_33090);
or U41648 (N_41648,N_33439,N_38620);
or U41649 (N_41649,N_33426,N_38936);
nand U41650 (N_41650,N_32814,N_38803);
nor U41651 (N_41651,N_35170,N_38496);
xnor U41652 (N_41652,N_31768,N_31688);
xnor U41653 (N_41653,N_31644,N_34073);
nor U41654 (N_41654,N_32670,N_33830);
nor U41655 (N_41655,N_33580,N_33681);
nor U41656 (N_41656,N_33559,N_37563);
or U41657 (N_41657,N_38215,N_38571);
nor U41658 (N_41658,N_39150,N_35180);
xnor U41659 (N_41659,N_34006,N_30704);
xor U41660 (N_41660,N_39066,N_32567);
nor U41661 (N_41661,N_30621,N_33899);
nor U41662 (N_41662,N_31431,N_38152);
and U41663 (N_41663,N_35974,N_33243);
nand U41664 (N_41664,N_32883,N_33643);
and U41665 (N_41665,N_39402,N_30210);
xnor U41666 (N_41666,N_37892,N_37860);
and U41667 (N_41667,N_35455,N_33953);
and U41668 (N_41668,N_35395,N_31772);
xnor U41669 (N_41669,N_32330,N_37337);
and U41670 (N_41670,N_33532,N_32143);
xor U41671 (N_41671,N_33966,N_36547);
xnor U41672 (N_41672,N_30307,N_39351);
or U41673 (N_41673,N_37550,N_30628);
or U41674 (N_41674,N_33954,N_34246);
xnor U41675 (N_41675,N_32160,N_35187);
and U41676 (N_41676,N_31090,N_33524);
xnor U41677 (N_41677,N_37895,N_34886);
and U41678 (N_41678,N_38204,N_31030);
or U41679 (N_41679,N_37846,N_34066);
nand U41680 (N_41680,N_38901,N_35396);
nor U41681 (N_41681,N_36820,N_34264);
or U41682 (N_41682,N_39671,N_37340);
nand U41683 (N_41683,N_32357,N_39381);
nor U41684 (N_41684,N_33795,N_30292);
or U41685 (N_41685,N_34517,N_39961);
or U41686 (N_41686,N_37312,N_35506);
xor U41687 (N_41687,N_36598,N_32607);
nand U41688 (N_41688,N_39333,N_32221);
xnor U41689 (N_41689,N_33631,N_35392);
nand U41690 (N_41690,N_39836,N_35841);
or U41691 (N_41691,N_38615,N_31617);
nor U41692 (N_41692,N_32236,N_34336);
nand U41693 (N_41693,N_38690,N_36470);
xor U41694 (N_41694,N_38513,N_35266);
or U41695 (N_41695,N_31905,N_39188);
or U41696 (N_41696,N_32548,N_32645);
nand U41697 (N_41697,N_30293,N_37715);
and U41698 (N_41698,N_39930,N_34843);
xor U41699 (N_41699,N_38255,N_33067);
and U41700 (N_41700,N_31949,N_33318);
or U41701 (N_41701,N_37087,N_35723);
or U41702 (N_41702,N_32939,N_33026);
or U41703 (N_41703,N_33677,N_39449);
nand U41704 (N_41704,N_33927,N_38662);
nor U41705 (N_41705,N_31879,N_38383);
nor U41706 (N_41706,N_32413,N_33386);
xnor U41707 (N_41707,N_31214,N_38715);
nand U41708 (N_41708,N_31806,N_36968);
and U41709 (N_41709,N_36248,N_30582);
or U41710 (N_41710,N_34706,N_37857);
or U41711 (N_41711,N_33820,N_38036);
nand U41712 (N_41712,N_31164,N_31965);
nand U41713 (N_41713,N_39723,N_37900);
nand U41714 (N_41714,N_35501,N_36953);
xor U41715 (N_41715,N_38012,N_32313);
and U41716 (N_41716,N_36260,N_33422);
and U41717 (N_41717,N_31864,N_38406);
or U41718 (N_41718,N_38248,N_39230);
and U41719 (N_41719,N_30198,N_37442);
nor U41720 (N_41720,N_37207,N_30366);
nand U41721 (N_41721,N_32747,N_36578);
or U41722 (N_41722,N_33616,N_37308);
nor U41723 (N_41723,N_35793,N_39318);
nand U41724 (N_41724,N_31608,N_32279);
nand U41725 (N_41725,N_36824,N_36631);
nand U41726 (N_41726,N_39474,N_39264);
and U41727 (N_41727,N_38572,N_38041);
or U41728 (N_41728,N_34660,N_38480);
or U41729 (N_41729,N_33492,N_37639);
and U41730 (N_41730,N_38268,N_37946);
nand U41731 (N_41731,N_32061,N_37614);
xor U41732 (N_41732,N_32951,N_37664);
xor U41733 (N_41733,N_35254,N_36679);
nor U41734 (N_41734,N_36082,N_30548);
nand U41735 (N_41735,N_31419,N_34653);
nand U41736 (N_41736,N_34669,N_30535);
or U41737 (N_41737,N_32122,N_33139);
and U41738 (N_41738,N_36494,N_38522);
xor U41739 (N_41739,N_38739,N_39573);
xor U41740 (N_41740,N_31489,N_35571);
nand U41741 (N_41741,N_30842,N_32907);
xor U41742 (N_41742,N_39368,N_34490);
nor U41743 (N_41743,N_38353,N_36872);
xnor U41744 (N_41744,N_38650,N_39496);
and U41745 (N_41745,N_32716,N_30397);
nand U41746 (N_41746,N_30296,N_37240);
and U41747 (N_41747,N_38387,N_36615);
or U41748 (N_41748,N_33223,N_32764);
nand U41749 (N_41749,N_30529,N_35276);
nor U41750 (N_41750,N_37654,N_34591);
nor U41751 (N_41751,N_35246,N_34608);
and U41752 (N_41752,N_36724,N_31605);
or U41753 (N_41753,N_31153,N_33740);
or U41754 (N_41754,N_31622,N_30455);
xnor U41755 (N_41755,N_35113,N_38783);
and U41756 (N_41756,N_36563,N_33975);
or U41757 (N_41757,N_37504,N_33092);
xor U41758 (N_41758,N_37777,N_36423);
nand U41759 (N_41759,N_34885,N_30113);
and U41760 (N_41760,N_35564,N_37030);
or U41761 (N_41761,N_33743,N_35831);
or U41762 (N_41762,N_34711,N_38217);
nor U41763 (N_41763,N_34007,N_32243);
and U41764 (N_41764,N_37815,N_38502);
nor U41765 (N_41765,N_35837,N_39504);
nor U41766 (N_41766,N_30037,N_34567);
xor U41767 (N_41767,N_39712,N_30249);
nor U41768 (N_41768,N_32470,N_32307);
and U41769 (N_41769,N_32240,N_39090);
and U41770 (N_41770,N_30303,N_30036);
xnor U41771 (N_41771,N_38389,N_37327);
and U41772 (N_41772,N_38167,N_35219);
nand U41773 (N_41773,N_38740,N_36251);
nand U41774 (N_41774,N_30184,N_30360);
or U41775 (N_41775,N_39430,N_33169);
xor U41776 (N_41776,N_39514,N_34529);
and U41777 (N_41777,N_36707,N_39364);
and U41778 (N_41778,N_31371,N_31929);
xor U41779 (N_41779,N_35682,N_31571);
or U41780 (N_41780,N_34049,N_38185);
or U41781 (N_41781,N_38973,N_37533);
nor U41782 (N_41782,N_39116,N_34136);
or U41783 (N_41783,N_36684,N_35198);
nand U41784 (N_41784,N_36370,N_33870);
nor U41785 (N_41785,N_31070,N_31805);
nor U41786 (N_41786,N_33234,N_38655);
nor U41787 (N_41787,N_35871,N_31187);
nor U41788 (N_41788,N_37266,N_35305);
or U41789 (N_41789,N_31953,N_36599);
nor U41790 (N_41790,N_34309,N_34369);
and U41791 (N_41791,N_36184,N_31791);
nor U41792 (N_41792,N_39165,N_39494);
nand U41793 (N_41793,N_32539,N_30645);
or U41794 (N_41794,N_36919,N_30992);
nand U41795 (N_41795,N_39584,N_35547);
or U41796 (N_41796,N_33372,N_32823);
nand U41797 (N_41797,N_37896,N_32265);
nor U41798 (N_41798,N_34539,N_36784);
or U41799 (N_41799,N_38399,N_31629);
xnor U41800 (N_41800,N_34399,N_34543);
xor U41801 (N_41801,N_31277,N_30928);
xnor U41802 (N_41802,N_30513,N_36285);
xor U41803 (N_41803,N_35413,N_31346);
xnor U41804 (N_41804,N_30127,N_31591);
nand U41805 (N_41805,N_33951,N_36282);
or U41806 (N_41806,N_31827,N_33107);
xor U41807 (N_41807,N_35315,N_36365);
xor U41808 (N_41808,N_37254,N_31405);
nand U41809 (N_41809,N_37725,N_33015);
nand U41810 (N_41810,N_39521,N_35404);
and U41811 (N_41811,N_37638,N_31579);
xor U41812 (N_41812,N_39669,N_31904);
or U41813 (N_41813,N_33100,N_32744);
nand U41814 (N_41814,N_36843,N_37194);
or U41815 (N_41815,N_32479,N_39195);
nor U41816 (N_41816,N_38365,N_30989);
xnor U41817 (N_41817,N_39131,N_32204);
nor U41818 (N_41818,N_30275,N_31091);
xnor U41819 (N_41819,N_30453,N_38946);
or U41820 (N_41820,N_38316,N_31974);
nor U41821 (N_41821,N_30163,N_30413);
nand U41822 (N_41822,N_36336,N_32224);
nor U41823 (N_41823,N_39227,N_30046);
xor U41824 (N_41824,N_36966,N_31848);
nand U41825 (N_41825,N_31533,N_36053);
or U41826 (N_41826,N_34739,N_34765);
and U41827 (N_41827,N_32976,N_34746);
and U41828 (N_41828,N_30144,N_39289);
or U41829 (N_41829,N_38297,N_38514);
nand U41830 (N_41830,N_39221,N_31212);
and U41831 (N_41831,N_34534,N_39234);
nand U41832 (N_41832,N_31538,N_38020);
xor U41833 (N_41833,N_31268,N_32005);
or U41834 (N_41834,N_33238,N_32979);
or U41835 (N_41835,N_34476,N_32886);
nor U41836 (N_41836,N_30598,N_30505);
nand U41837 (N_41837,N_31434,N_35991);
and U41838 (N_41838,N_38628,N_39967);
xor U41839 (N_41839,N_32727,N_36798);
xnor U41840 (N_41840,N_37969,N_39710);
nand U41841 (N_41841,N_35324,N_30349);
or U41842 (N_41842,N_36778,N_37689);
nand U41843 (N_41843,N_31103,N_33805);
and U41844 (N_41844,N_34874,N_36976);
or U41845 (N_41845,N_38092,N_34896);
nor U41846 (N_41846,N_34152,N_37717);
or U41847 (N_41847,N_31129,N_38516);
xnor U41848 (N_41848,N_33040,N_37140);
nor U41849 (N_41849,N_33433,N_31833);
or U41850 (N_41850,N_38087,N_37656);
or U41851 (N_41851,N_35283,N_33445);
xnor U41852 (N_41852,N_32476,N_31900);
and U41853 (N_41853,N_31649,N_37553);
nor U41854 (N_41854,N_31895,N_38838);
or U41855 (N_41855,N_37050,N_30247);
xnor U41856 (N_41856,N_33023,N_30610);
and U41857 (N_41857,N_35314,N_38723);
or U41858 (N_41858,N_34579,N_37996);
or U41859 (N_41859,N_39787,N_39629);
and U41860 (N_41860,N_38289,N_34778);
xnor U41861 (N_41861,N_32025,N_32134);
xnor U41862 (N_41862,N_37681,N_35669);
nand U41863 (N_41863,N_34150,N_34020);
or U41864 (N_41864,N_31868,N_38070);
nand U41865 (N_41865,N_34081,N_38675);
nand U41866 (N_41866,N_30128,N_31482);
nor U41867 (N_41867,N_39931,N_36483);
nand U41868 (N_41868,N_32641,N_37891);
nor U41869 (N_41869,N_32178,N_33907);
xnor U41870 (N_41870,N_30190,N_38308);
xnor U41871 (N_41871,N_30528,N_34766);
nor U41872 (N_41872,N_39858,N_34575);
or U41873 (N_41873,N_32677,N_31060);
nand U41874 (N_41874,N_37118,N_39022);
xor U41875 (N_41875,N_34906,N_39944);
nor U41876 (N_41876,N_30499,N_32964);
nor U41877 (N_41877,N_39453,N_32241);
xnor U41878 (N_41878,N_30547,N_38132);
nor U41879 (N_41879,N_35175,N_31828);
nor U41880 (N_41880,N_35969,N_38547);
nor U41881 (N_41881,N_36141,N_33454);
nand U41882 (N_41882,N_39696,N_35446);
xor U41883 (N_41883,N_38577,N_30919);
nand U41884 (N_41884,N_36634,N_37286);
xor U41885 (N_41885,N_33046,N_30401);
nand U41886 (N_41886,N_38764,N_34506);
and U41887 (N_41887,N_39314,N_33440);
xor U41888 (N_41888,N_39792,N_33236);
and U41889 (N_41889,N_32689,N_33573);
xor U41890 (N_41890,N_30418,N_38013);
nor U41891 (N_41891,N_36038,N_34817);
and U41892 (N_41892,N_35720,N_37368);
or U41893 (N_41893,N_38379,N_31503);
and U41894 (N_41894,N_36656,N_32688);
xor U41895 (N_41895,N_30775,N_38703);
or U41896 (N_41896,N_36031,N_35221);
xor U41897 (N_41897,N_32728,N_37100);
nor U41898 (N_41898,N_39988,N_37850);
and U41899 (N_41899,N_36220,N_38695);
or U41900 (N_41900,N_34992,N_39340);
nand U41901 (N_41901,N_31985,N_34597);
nand U41902 (N_41902,N_36043,N_33043);
and U41903 (N_41903,N_31086,N_34604);
xnor U41904 (N_41904,N_39303,N_33607);
or U41905 (N_41905,N_34279,N_31603);
or U41906 (N_41906,N_31134,N_38504);
or U41907 (N_41907,N_39957,N_38809);
and U41908 (N_41908,N_33357,N_35293);
or U41909 (N_41909,N_31202,N_31465);
or U41910 (N_41910,N_36228,N_35087);
and U41911 (N_41911,N_33369,N_38125);
or U41912 (N_41912,N_30597,N_39754);
and U41913 (N_41913,N_32094,N_36842);
and U41914 (N_41914,N_39341,N_33761);
or U41915 (N_41915,N_30010,N_31857);
xnor U41916 (N_41916,N_36295,N_32289);
or U41917 (N_41917,N_36022,N_34725);
and U41918 (N_41918,N_30178,N_37114);
xor U41919 (N_41919,N_34270,N_36566);
nand U41920 (N_41920,N_38259,N_31795);
nand U41921 (N_41921,N_36105,N_36747);
nand U41922 (N_41922,N_36023,N_33490);
and U41923 (N_41923,N_34752,N_30179);
or U41924 (N_41924,N_31722,N_39118);
or U41925 (N_41925,N_32333,N_31621);
and U41926 (N_41926,N_33103,N_38535);
nand U41927 (N_41927,N_38629,N_30434);
and U41928 (N_41928,N_33124,N_34341);
nor U41929 (N_41929,N_36455,N_37645);
nor U41930 (N_41930,N_35943,N_32499);
xnor U41931 (N_41931,N_37527,N_35440);
and U41932 (N_41932,N_34095,N_34609);
or U41933 (N_41933,N_36078,N_37642);
or U41934 (N_41934,N_31625,N_37779);
or U41935 (N_41935,N_33036,N_32184);
and U41936 (N_41936,N_31469,N_39690);
xor U41937 (N_41937,N_37017,N_35510);
nand U41938 (N_41938,N_30428,N_32610);
nor U41939 (N_41939,N_35013,N_39466);
or U41940 (N_41940,N_31368,N_37847);
and U41941 (N_41941,N_34537,N_32181);
and U41942 (N_41942,N_33647,N_36792);
or U41943 (N_41943,N_39811,N_32842);
or U41944 (N_41944,N_33451,N_39867);
or U41945 (N_41945,N_35680,N_31754);
or U41946 (N_41946,N_31117,N_34024);
or U41947 (N_41947,N_39252,N_34323);
xor U41948 (N_41948,N_36951,N_35906);
and U41949 (N_41949,N_39006,N_37213);
nand U41950 (N_41950,N_39833,N_36763);
nor U41951 (N_41951,N_39802,N_35983);
nand U41952 (N_41952,N_39613,N_33280);
and U41953 (N_41953,N_37584,N_31244);
nand U41954 (N_41954,N_35751,N_37159);
nor U41955 (N_41955,N_35967,N_35627);
or U41956 (N_41956,N_31144,N_39224);
nand U41957 (N_41957,N_39642,N_31366);
nand U41958 (N_41958,N_30131,N_38639);
nand U41959 (N_41959,N_38045,N_36234);
nor U41960 (N_41960,N_33296,N_31285);
nor U41961 (N_41961,N_37867,N_30978);
nor U41962 (N_41962,N_33709,N_30986);
and U41963 (N_41963,N_35786,N_36801);
xor U41964 (N_41964,N_39704,N_38103);
nor U41965 (N_41965,N_37997,N_32733);
nand U41966 (N_41966,N_30793,N_30850);
or U41967 (N_41967,N_35197,N_36827);
nand U41968 (N_41968,N_39347,N_36303);
xor U41969 (N_41969,N_39201,N_38947);
nand U41970 (N_41970,N_35014,N_34875);
and U41971 (N_41971,N_37448,N_36652);
or U41972 (N_41972,N_37826,N_38807);
or U41973 (N_41973,N_36740,N_35348);
nand U41974 (N_41974,N_30778,N_33324);
nand U41975 (N_41975,N_32685,N_37873);
or U41976 (N_41976,N_32557,N_31410);
xnor U41977 (N_41977,N_35508,N_36345);
xnor U41978 (N_41978,N_33358,N_31133);
and U41979 (N_41979,N_32300,N_30949);
or U41980 (N_41980,N_32102,N_39047);
and U41981 (N_41981,N_33200,N_33292);
xor U41982 (N_41982,N_38276,N_38371);
xnor U41983 (N_41983,N_34855,N_34573);
nand U41984 (N_41984,N_37277,N_30538);
nand U41985 (N_41985,N_32966,N_31993);
xor U41986 (N_41986,N_30906,N_33713);
and U41987 (N_41987,N_31038,N_39589);
or U41988 (N_41988,N_37773,N_31388);
or U41989 (N_41989,N_32431,N_36545);
nor U41990 (N_41990,N_38477,N_35332);
or U41991 (N_41991,N_35724,N_31695);
nor U41992 (N_41992,N_36405,N_30655);
and U41993 (N_41993,N_31236,N_37018);
nand U41994 (N_41994,N_34368,N_34781);
nor U41995 (N_41995,N_33745,N_36699);
or U41996 (N_41996,N_37894,N_37970);
and U41997 (N_41997,N_37637,N_35020);
or U41998 (N_41998,N_38360,N_37347);
and U41999 (N_41999,N_36606,N_39422);
nor U42000 (N_42000,N_39200,N_39447);
xor U42001 (N_42001,N_34675,N_35839);
nand U42002 (N_42002,N_37206,N_31126);
nand U42003 (N_42003,N_30242,N_34957);
or U42004 (N_42004,N_32020,N_35800);
or U42005 (N_42005,N_37832,N_30416);
and U42006 (N_42006,N_39475,N_33218);
nand U42007 (N_42007,N_32711,N_37478);
nand U42008 (N_42008,N_33797,N_34407);
nand U42009 (N_42009,N_37917,N_36758);
or U42010 (N_42010,N_36691,N_34330);
xnor U42011 (N_42011,N_37416,N_30365);
nor U42012 (N_42012,N_33028,N_32831);
nor U42013 (N_42013,N_35711,N_38773);
or U42014 (N_42014,N_37406,N_36328);
xor U42015 (N_42015,N_35447,N_36593);
xor U42016 (N_42016,N_32622,N_38139);
or U42017 (N_42017,N_34694,N_32449);
nand U42018 (N_42018,N_33793,N_39721);
or U42019 (N_42019,N_31898,N_31550);
nand U42020 (N_42020,N_30322,N_33469);
or U42021 (N_42021,N_31416,N_34606);
or U42022 (N_42022,N_31420,N_32942);
nand U42023 (N_42023,N_38188,N_33007);
or U42024 (N_42024,N_39808,N_39478);
nor U42025 (N_42025,N_33876,N_39692);
and U42026 (N_42026,N_31500,N_31049);
and U42027 (N_42027,N_38762,N_39419);
and U42028 (N_42028,N_38501,N_31745);
or U42029 (N_42029,N_36006,N_34813);
or U42030 (N_42030,N_31288,N_37105);
and U42031 (N_42031,N_34846,N_33622);
nor U42032 (N_42032,N_31798,N_37023);
nand U42033 (N_42033,N_34201,N_36595);
xor U42034 (N_42034,N_38143,N_32932);
nand U42035 (N_42035,N_34278,N_34230);
and U42036 (N_42036,N_35845,N_36354);
nor U42037 (N_42037,N_30490,N_37476);
and U42038 (N_42038,N_37228,N_32095);
and U42039 (N_42039,N_36587,N_31057);
or U42040 (N_42040,N_36661,N_36512);
nand U42041 (N_42041,N_31502,N_30302);
nand U42042 (N_42042,N_39887,N_35892);
nor U42043 (N_42043,N_30780,N_34607);
nor U42044 (N_42044,N_35672,N_37383);
nor U42045 (N_42045,N_35629,N_30238);
nand U42046 (N_42046,N_39005,N_33215);
and U42047 (N_42047,N_36879,N_31271);
or U42048 (N_42048,N_39752,N_33623);
or U42049 (N_42049,N_32276,N_34936);
xnor U42050 (N_42050,N_35351,N_36781);
nand U42051 (N_42051,N_36880,N_35727);
nor U42052 (N_42052,N_33356,N_35901);
nand U42053 (N_42053,N_35115,N_35444);
nor U42054 (N_42054,N_34393,N_39649);
xor U42055 (N_42055,N_30431,N_35765);
or U42056 (N_42056,N_32498,N_38037);
and U42057 (N_42057,N_34612,N_30092);
and U42058 (N_42058,N_37993,N_34756);
nand U42059 (N_42059,N_30343,N_33766);
nor U42060 (N_42060,N_34741,N_32656);
and U42061 (N_42061,N_34382,N_31440);
nand U42062 (N_42062,N_33653,N_37875);
nand U42063 (N_42063,N_37714,N_38269);
xor U42064 (N_42064,N_37505,N_37429);
nand U42065 (N_42065,N_31240,N_33851);
nand U42066 (N_42066,N_32534,N_37808);
or U42067 (N_42067,N_34306,N_32244);
and U42068 (N_42068,N_36621,N_32353);
nand U42069 (N_42069,N_38405,N_38481);
and U42070 (N_42070,N_34442,N_32117);
or U42071 (N_42071,N_39484,N_31647);
nor U42072 (N_42072,N_37164,N_36580);
nor U42073 (N_42073,N_31871,N_30317);
xor U42074 (N_42074,N_34887,N_32803);
and U42075 (N_42075,N_32626,N_36416);
nor U42076 (N_42076,N_37514,N_31392);
xor U42077 (N_42077,N_30790,N_33764);
nor U42078 (N_42078,N_31270,N_37376);
nor U42079 (N_42079,N_30286,N_32595);
or U42080 (N_42080,N_31051,N_39831);
nor U42081 (N_42081,N_31831,N_31207);
or U42082 (N_42082,N_33282,N_37353);
nand U42083 (N_42083,N_30496,N_30404);
or U42084 (N_42084,N_39098,N_35748);
nor U42085 (N_42085,N_39884,N_36346);
and U42086 (N_42086,N_31351,N_37372);
or U42087 (N_42087,N_37510,N_38482);
or U42088 (N_42088,N_37326,N_30827);
nor U42089 (N_42089,N_31435,N_31109);
xnor U42090 (N_42090,N_39403,N_38010);
nor U42091 (N_42091,N_37519,N_31906);
or U42092 (N_42092,N_37396,N_36452);
and U42093 (N_42093,N_35498,N_36188);
nor U42094 (N_42094,N_39048,N_36552);
nor U42095 (N_42095,N_32904,N_39183);
or U42096 (N_42096,N_35594,N_32227);
or U42097 (N_42097,N_36481,N_32484);
nand U42098 (N_42098,N_36607,N_33747);
xnor U42099 (N_42099,N_33986,N_34620);
or U42100 (N_42100,N_34663,N_35541);
nor U42101 (N_42101,N_32944,N_33142);
nor U42102 (N_42102,N_38930,N_31539);
nand U42103 (N_42103,N_31466,N_30705);
nor U42104 (N_42104,N_33031,N_33147);
xor U42105 (N_42105,N_33908,N_35225);
or U42106 (N_42106,N_33823,N_33349);
nor U42107 (N_42107,N_37621,N_36926);
nor U42108 (N_42108,N_39258,N_39755);
xnor U42109 (N_42109,N_35333,N_32516);
xor U42110 (N_42110,N_31913,N_32255);
and U42111 (N_42111,N_36441,N_38570);
or U42112 (N_42112,N_38608,N_38827);
xor U42113 (N_42113,N_39557,N_37022);
nand U42114 (N_42114,N_31729,N_31101);
xor U42115 (N_42115,N_39202,N_36436);
and U42116 (N_42116,N_31685,N_31228);
or U42117 (N_42117,N_31131,N_37062);
or U42118 (N_42118,N_35470,N_39087);
and U42119 (N_42119,N_39215,N_32179);
and U42120 (N_42120,N_31632,N_34421);
xor U42121 (N_42121,N_33328,N_38106);
and U42122 (N_42122,N_30980,N_30380);
and U42123 (N_42123,N_30233,N_34538);
or U42124 (N_42124,N_31139,N_35655);
nand U42125 (N_42125,N_36998,N_33940);
and U42126 (N_42126,N_38230,N_30635);
nand U42127 (N_42127,N_36204,N_38361);
nand U42128 (N_42128,N_39020,N_35843);
nor U42129 (N_42129,N_39160,N_31150);
nor U42130 (N_42130,N_31628,N_36800);
or U42131 (N_42131,N_33788,N_34689);
nand U42132 (N_42132,N_39730,N_38382);
and U42133 (N_42133,N_33800,N_35296);
nor U42134 (N_42134,N_35386,N_30214);
or U42135 (N_42135,N_30276,N_30796);
and U42136 (N_42136,N_39560,N_35429);
nand U42137 (N_42137,N_31387,N_38491);
xor U42138 (N_42138,N_30419,N_32403);
nand U42139 (N_42139,N_33368,N_35960);
xor U42140 (N_42140,N_36268,N_33533);
or U42141 (N_42141,N_34033,N_32941);
and U42142 (N_42142,N_34367,N_34594);
or U42143 (N_42143,N_35195,N_32536);
or U42144 (N_42144,N_39352,N_37589);
and U42145 (N_42145,N_35797,N_33320);
or U42146 (N_42146,N_31315,N_33411);
or U42147 (N_42147,N_33978,N_31813);
nand U42148 (N_42148,N_35653,N_33250);
nor U42149 (N_42149,N_35075,N_33683);
nand U42150 (N_42150,N_38444,N_34184);
nand U42151 (N_42151,N_32729,N_38349);
nor U42152 (N_42152,N_33190,N_39380);
xor U42153 (N_42153,N_34687,N_31408);
nand U42154 (N_42154,N_35491,N_32281);
xor U42155 (N_42155,N_35648,N_32614);
nor U42156 (N_42156,N_37211,N_31407);
and U42157 (N_42157,N_33060,N_38221);
or U42158 (N_42158,N_31413,N_31262);
or U42159 (N_42159,N_34364,N_39406);
or U42160 (N_42160,N_30595,N_33259);
and U42161 (N_42161,N_37515,N_32807);
nand U42162 (N_42162,N_38738,N_34719);
and U42163 (N_42163,N_34212,N_39816);
or U42164 (N_42164,N_38886,N_32856);
or U42165 (N_42165,N_38114,N_30381);
nor U42166 (N_42166,N_39555,N_38300);
or U42167 (N_42167,N_35073,N_33763);
and U42168 (N_42168,N_32766,N_33442);
or U42169 (N_42169,N_30462,N_37438);
or U42170 (N_42170,N_37172,N_36327);
nor U42171 (N_42171,N_30600,N_35670);
or U42172 (N_42172,N_38388,N_30556);
or U42173 (N_42173,N_37290,N_35370);
and U42174 (N_42174,N_30048,N_36739);
nor U42175 (N_42175,N_32391,N_37064);
and U42176 (N_42176,N_39378,N_39702);
nor U42177 (N_42177,N_35803,N_36359);
nand U42178 (N_42178,N_37650,N_39143);
nand U42179 (N_42179,N_34378,N_33659);
xor U42180 (N_42180,N_38527,N_34633);
xor U42181 (N_42181,N_39391,N_36196);
or U42182 (N_42182,N_31723,N_30488);
nor U42183 (N_42183,N_34856,N_31944);
and U42184 (N_42184,N_38772,N_31962);
nor U42185 (N_42185,N_34174,N_37537);
nand U42186 (N_42186,N_31559,N_33421);
and U42187 (N_42187,N_32277,N_36989);
nor U42188 (N_42188,N_33102,N_30862);
xnor U42189 (N_42189,N_39682,N_30078);
and U42190 (N_42190,N_36355,N_37910);
and U42191 (N_42191,N_39739,N_39142);
and U42192 (N_42192,N_37972,N_30120);
xor U42193 (N_42193,N_35883,N_35527);
nor U42194 (N_42194,N_33106,N_38971);
xor U42195 (N_42195,N_32207,N_37512);
nor U42196 (N_42196,N_39198,N_32597);
and U42197 (N_42197,N_36895,N_37010);
nor U42198 (N_42198,N_30819,N_36866);
or U42199 (N_42199,N_38692,N_31661);
or U42200 (N_42200,N_36498,N_34038);
nor U42201 (N_42201,N_39909,N_30571);
nand U42202 (N_42202,N_33245,N_34254);
and U42203 (N_42203,N_33869,N_37939);
and U42204 (N_42204,N_35496,N_34974);
or U42205 (N_42205,N_38678,N_37354);
or U42206 (N_42206,N_38080,N_33802);
nor U42207 (N_42207,N_38602,N_39919);
and U42208 (N_42208,N_30301,N_37397);
nand U42209 (N_42209,N_36349,N_34953);
nand U42210 (N_42210,N_32106,N_31884);
nor U42211 (N_42211,N_35334,N_32583);
nand U42212 (N_42212,N_34433,N_33592);
nor U42213 (N_42213,N_37795,N_36000);
xor U42214 (N_42214,N_37962,N_33340);
and U42215 (N_42215,N_30532,N_33447);
or U42216 (N_42216,N_30975,N_35481);
nor U42217 (N_42217,N_32538,N_37210);
nor U42218 (N_42218,N_36102,N_36089);
and U42219 (N_42219,N_33815,N_37423);
xor U42220 (N_42220,N_34777,N_33637);
nand U42221 (N_42221,N_37626,N_35035);
nor U42222 (N_42222,N_39767,N_36669);
nand U42223 (N_42223,N_33458,N_38963);
and U42224 (N_42224,N_32150,N_30188);
and U42225 (N_42225,N_30267,N_30463);
or U42226 (N_42226,N_33572,N_32715);
and U42227 (N_42227,N_38636,N_38307);
xor U42228 (N_42228,N_31395,N_32136);
xor U42229 (N_42229,N_31358,N_39348);
nor U42230 (N_42230,N_30442,N_37748);
nand U42231 (N_42231,N_37730,N_31367);
nor U42232 (N_42232,N_38967,N_38626);
or U42233 (N_42233,N_31938,N_31217);
and U42234 (N_42234,N_37384,N_32345);
nand U42235 (N_42235,N_33029,N_32794);
nor U42236 (N_42236,N_36590,N_37693);
xnor U42237 (N_42237,N_36928,N_34294);
nand U42238 (N_42238,N_33758,N_36036);
and U42239 (N_42239,N_39100,N_31480);
nand U42240 (N_42240,N_37524,N_34209);
nor U42241 (N_42241,N_30082,N_34112);
nand U42242 (N_42242,N_39163,N_38488);
and U42243 (N_42243,N_36003,N_31374);
and U42244 (N_42244,N_33595,N_37293);
xor U42245 (N_42245,N_33366,N_33204);
and U42246 (N_42246,N_35788,N_39581);
or U42247 (N_42247,N_31259,N_38916);
nand U42248 (N_42248,N_33463,N_35921);
xnor U42249 (N_42249,N_39173,N_38635);
nand U42250 (N_42250,N_38756,N_39718);
or U42251 (N_42251,N_39873,N_33544);
nand U42252 (N_42252,N_37977,N_30757);
nand U42253 (N_42253,N_34291,N_34681);
and U42254 (N_42254,N_31007,N_35612);
nand U42255 (N_42255,N_39000,N_39998);
nor U42256 (N_42256,N_37767,N_38372);
xnor U42257 (N_42257,N_34884,N_31580);
xor U42258 (N_42258,N_31855,N_37063);
nand U42259 (N_42259,N_31509,N_38965);
xnor U42260 (N_42260,N_34453,N_31513);
or U42261 (N_42261,N_34461,N_37668);
and U42262 (N_42262,N_30593,N_33126);
or U42263 (N_42263,N_36095,N_36262);
xnor U42264 (N_42264,N_34111,N_32789);
xnor U42265 (N_42265,N_38317,N_33158);
or U42266 (N_42266,N_30848,N_30278);
or U42267 (N_42267,N_38799,N_34320);
nand U42268 (N_42268,N_34532,N_30108);
or U42269 (N_42269,N_33638,N_33150);
nand U42270 (N_42270,N_30151,N_33584);
and U42271 (N_42271,N_39382,N_31801);
nand U42272 (N_42272,N_30952,N_39457);
nand U42273 (N_42273,N_35859,N_33341);
xor U42274 (N_42274,N_30468,N_39650);
nand U42275 (N_42275,N_32274,N_37066);
nor U42276 (N_42276,N_31426,N_38210);
xor U42277 (N_42277,N_34053,N_36183);
xor U42278 (N_42278,N_37197,N_34010);
or U42279 (N_42279,N_36751,N_39452);
and U42280 (N_42280,N_37942,N_31213);
nor U42281 (N_42281,N_33853,N_30814);
and U42282 (N_42282,N_35096,N_38696);
or U42283 (N_42283,N_35652,N_30344);
and U42284 (N_42284,N_37113,N_38280);
xor U42285 (N_42285,N_37357,N_34116);
nor U42286 (N_42286,N_37641,N_34587);
nor U42287 (N_42287,N_31592,N_37444);
nand U42288 (N_42288,N_32586,N_35022);
or U42289 (N_42289,N_30450,N_36457);
and U42290 (N_42290,N_32114,N_30057);
and U42291 (N_42291,N_31013,N_35693);
xnor U42292 (N_42292,N_38174,N_32206);
or U42293 (N_42293,N_39737,N_30580);
nor U42294 (N_42294,N_31224,N_36737);
and U42295 (N_42295,N_33345,N_37683);
and U42296 (N_42296,N_34108,N_36149);
and U42297 (N_42297,N_39017,N_30771);
xnor U42298 (N_42298,N_39137,N_35218);
xor U42299 (N_42299,N_39413,N_31394);
and U42300 (N_42300,N_36137,N_32254);
xnor U42301 (N_42301,N_38175,N_34851);
nor U42302 (N_42302,N_31040,N_30675);
nor U42303 (N_42303,N_38811,N_38208);
and U42304 (N_42304,N_33971,N_37755);
nand U42305 (N_42305,N_36831,N_33834);
xnor U42306 (N_42306,N_37632,N_33718);
or U42307 (N_42307,N_35512,N_35975);
nor U42308 (N_42308,N_34173,N_33175);
nor U42309 (N_42309,N_36712,N_30945);
nand U42310 (N_42310,N_30185,N_37157);
nand U42311 (N_42311,N_33482,N_30223);
xor U42312 (N_42312,N_32101,N_35889);
nand U42313 (N_42313,N_35515,N_33585);
xor U42314 (N_42314,N_34089,N_33771);
or U42315 (N_42315,N_35344,N_36322);
nand U42316 (N_42316,N_38843,N_35741);
nor U42317 (N_42317,N_32535,N_32416);
and U42318 (N_42318,N_39913,N_35584);
xor U42319 (N_42319,N_34513,N_33390);
xor U42320 (N_42320,N_38091,N_37306);
xnor U42321 (N_42321,N_39785,N_33909);
and U42322 (N_42322,N_34245,N_32623);
or U42323 (N_42323,N_31715,N_30681);
and U42324 (N_42324,N_35650,N_32572);
and U42325 (N_42325,N_39578,N_38333);
nand U42326 (N_42326,N_34610,N_36555);
and U42327 (N_42327,N_35484,N_33867);
nand U42328 (N_42328,N_35659,N_36249);
and U42329 (N_42329,N_36152,N_31229);
nor U42330 (N_42330,N_32720,N_35856);
nand U42331 (N_42331,N_33633,N_33527);
or U42332 (N_42332,N_39192,N_30982);
or U42333 (N_42333,N_35759,N_30439);
xnor U42334 (N_42334,N_39888,N_39749);
nor U42335 (N_42335,N_39236,N_35904);
and U42336 (N_42336,N_34475,N_36826);
or U42337 (N_42337,N_38374,N_37278);
nor U42338 (N_42338,N_31582,N_34557);
and U42339 (N_42339,N_38334,N_34428);
nand U42340 (N_42340,N_33206,N_31733);
nor U42341 (N_42341,N_31329,N_38708);
nand U42342 (N_42342,N_33672,N_31565);
nand U42343 (N_42343,N_33319,N_31838);
nand U42344 (N_42344,N_35888,N_38674);
xor U42345 (N_42345,N_39876,N_32370);
nor U42346 (N_42346,N_37304,N_38282);
xnor U42347 (N_42347,N_30169,N_31867);
and U42348 (N_42348,N_37132,N_38677);
xor U42349 (N_42349,N_32352,N_37215);
nor U42350 (N_42350,N_34966,N_35632);
nand U42351 (N_42351,N_37257,N_33614);
nand U42352 (N_42352,N_34097,N_31854);
nor U42353 (N_42353,N_33910,N_31068);
and U42354 (N_42354,N_37054,N_33974);
nor U42355 (N_42355,N_39427,N_30996);
xor U42356 (N_42356,N_33174,N_30690);
and U42357 (N_42357,N_34857,N_30531);
nand U42358 (N_42358,N_38130,N_34379);
xor U42359 (N_42359,N_35566,N_32997);
nand U42360 (N_42360,N_34934,N_38611);
nand U42361 (N_42361,N_36446,N_33981);
or U42362 (N_42362,N_38805,N_35416);
xor U42363 (N_42363,N_32994,N_30368);
or U42364 (N_42364,N_31122,N_34365);
nand U42365 (N_42365,N_35819,N_31507);
or U42366 (N_42366,N_35340,N_34509);
xnor U42367 (N_42367,N_34904,N_30683);
or U42368 (N_42368,N_35699,N_38581);
or U42369 (N_42369,N_33922,N_32533);
nand U42370 (N_42370,N_34130,N_38823);
xnor U42371 (N_42371,N_37698,N_30892);
xor U42372 (N_42372,N_30330,N_31532);
and U42373 (N_42373,N_34268,N_30398);
or U42374 (N_42374,N_39079,N_35322);
and U42375 (N_42375,N_38321,N_39417);
and U42376 (N_42376,N_32469,N_30707);
nand U42377 (N_42377,N_31931,N_34866);
nand U42378 (N_42378,N_32422,N_37166);
nor U42379 (N_42379,N_34085,N_39662);
and U42380 (N_42380,N_30166,N_33083);
or U42381 (N_42381,N_34925,N_31136);
or U42382 (N_42382,N_36127,N_30208);
nor U42383 (N_42383,N_39122,N_34308);
and U42384 (N_42384,N_35443,N_30766);
nand U42385 (N_42385,N_35290,N_38219);
or U42386 (N_42386,N_38445,N_39240);
and U42387 (N_42387,N_36311,N_37014);
and U42388 (N_42388,N_34457,N_36509);
nor U42389 (N_42389,N_30603,N_35822);
nand U42390 (N_42390,N_31570,N_37983);
nor U42391 (N_42391,N_38729,N_39008);
and U42392 (N_42392,N_38439,N_30691);
or U42393 (N_42393,N_39220,N_37202);
xnor U42394 (N_42394,N_38603,N_33378);
nand U42395 (N_42395,N_34390,N_39511);
or U42396 (N_42396,N_37334,N_30435);
nand U42397 (N_42397,N_33032,N_31761);
or U42398 (N_42398,N_38836,N_34613);
xnor U42399 (N_42399,N_32372,N_31701);
and U42400 (N_42400,N_31146,N_38223);
nor U42401 (N_42401,N_30156,N_30027);
nand U42402 (N_42402,N_36004,N_31355);
and U42403 (N_42403,N_36996,N_36007);
or U42404 (N_42404,N_30607,N_31743);
nand U42405 (N_42405,N_30561,N_38234);
nand U42406 (N_42406,N_32198,N_32680);
or U42407 (N_42407,N_32454,N_34710);
nand U42408 (N_42408,N_37541,N_32676);
xor U42409 (N_42409,N_34998,N_32408);
xor U42410 (N_42410,N_38913,N_36735);
nand U42411 (N_42411,N_32642,N_33307);
nand U42412 (N_42412,N_30387,N_34617);
and U42413 (N_42413,N_34454,N_37056);
and U42414 (N_42414,N_38157,N_32938);
xor U42415 (N_42415,N_37097,N_32825);
xor U42416 (N_42416,N_34940,N_31750);
or U42417 (N_42417,N_39742,N_35869);
xnor U42418 (N_42418,N_34549,N_35996);
nand U42419 (N_42419,N_35206,N_31720);
xnor U42420 (N_42420,N_32643,N_38131);
and U42421 (N_42421,N_36899,N_30596);
nand U42422 (N_42422,N_32909,N_35874);
nor U42423 (N_42423,N_32249,N_36519);
nor U42424 (N_42424,N_39245,N_34826);
nor U42425 (N_42425,N_30515,N_33468);
xnor U42426 (N_42426,N_35544,N_36960);
nand U42427 (N_42427,N_39938,N_32411);
or U42428 (N_42428,N_36209,N_37647);
nor U42429 (N_42429,N_32048,N_37880);
nor U42430 (N_42430,N_33783,N_37670);
nor U42431 (N_42431,N_36997,N_31283);
or U42432 (N_42432,N_33030,N_37445);
and U42433 (N_42433,N_37284,N_30818);
xor U42434 (N_42434,N_31716,N_34293);
xnor U42435 (N_42435,N_39950,N_33629);
xnor U42436 (N_42436,N_31412,N_36297);
or U42437 (N_42437,N_36477,N_31381);
or U42438 (N_42438,N_35349,N_32756);
nor U42439 (N_42439,N_36450,N_36873);
or U42440 (N_42440,N_39577,N_34239);
xnor U42441 (N_42441,N_35257,N_34416);
and U42442 (N_42442,N_30846,N_35855);
or U42443 (N_42443,N_35796,N_36449);
or U42444 (N_42444,N_33244,N_39885);
and U42445 (N_42445,N_34688,N_32007);
nor U42446 (N_42446,N_35089,N_36783);
xnor U42447 (N_42447,N_32425,N_30855);
and U42448 (N_42448,N_33415,N_39772);
nor U42449 (N_42449,N_34939,N_34440);
and U42450 (N_42450,N_36286,N_35306);
or U42451 (N_42451,N_36964,N_39442);
nand U42452 (N_42452,N_31325,N_39583);
xnor U42453 (N_42453,N_35557,N_33212);
or U42454 (N_42454,N_34441,N_35528);
xnor U42455 (N_42455,N_36834,N_30384);
and U42456 (N_42456,N_39450,N_35065);
xnor U42457 (N_42457,N_35069,N_38034);
nor U42458 (N_42458,N_30420,N_37234);
nand U42459 (N_42459,N_37801,N_36727);
and U42460 (N_42460,N_38449,N_33531);
xnor U42461 (N_42461,N_37845,N_34179);
nand U42462 (N_42462,N_31658,N_33479);
xnor U42463 (N_42463,N_34637,N_30890);
or U42464 (N_42464,N_32995,N_34515);
xor U42465 (N_42465,N_30465,N_38133);
xor U42466 (N_42466,N_32405,N_31520);
and U42467 (N_42467,N_34162,N_38359);
or U42468 (N_42468,N_39935,N_38830);
xor U42469 (N_42469,N_35424,N_33293);
and U42470 (N_42470,N_38390,N_38574);
xnor U42471 (N_42471,N_34707,N_33956);
nand U42472 (N_42472,N_34380,N_35289);
or U42473 (N_42473,N_39594,N_34498);
xor U42474 (N_42474,N_36846,N_31811);
and U42475 (N_42475,N_39592,N_33724);
nor U42476 (N_42476,N_39590,N_37084);
nor U42477 (N_42477,N_37303,N_36550);
xnor U42478 (N_42478,N_38657,N_30237);
and U42479 (N_42479,N_36400,N_39409);
xor U42480 (N_42480,N_37555,N_34901);
nand U42481 (N_42481,N_37879,N_35716);
nor U42482 (N_42482,N_31638,N_31508);
and U42483 (N_42483,N_37820,N_35678);
xor U42484 (N_42484,N_35449,N_38561);
nand U42485 (N_42485,N_31108,N_31989);
nand U42486 (N_42486,N_39503,N_37315);
nand U42487 (N_42487,N_34839,N_30015);
nand U42488 (N_42488,N_31289,N_33734);
nand U42489 (N_42489,N_37501,N_39462);
nand U42490 (N_42490,N_36172,N_31047);
or U42491 (N_42491,N_35588,N_31331);
xnor U42492 (N_42492,N_36881,N_35777);
and U42493 (N_42493,N_34050,N_36192);
or U42494 (N_42494,N_35226,N_31651);
and U42495 (N_42495,N_35525,N_39286);
xor U42496 (N_42496,N_39046,N_34545);
xor U42497 (N_42497,N_35706,N_32171);
and U42498 (N_42498,N_30213,N_33552);
or U42499 (N_42499,N_36954,N_34114);
nor U42500 (N_42500,N_32259,N_32328);
and U42501 (N_42501,N_39843,N_31310);
nor U42502 (N_42502,N_37046,N_35291);
xor U42503 (N_42503,N_39288,N_30795);
nand U42504 (N_42504,N_36165,N_35361);
nand U42505 (N_42505,N_34527,N_32864);
or U42506 (N_42506,N_39117,N_30408);
xnor U42507 (N_42507,N_34952,N_37611);
nand U42508 (N_42508,N_33338,N_38003);
nor U42509 (N_42509,N_36718,N_31294);
xor U42510 (N_42510,N_32035,N_33460);
nand U42511 (N_42511,N_37192,N_33721);
and U42512 (N_42512,N_35282,N_34054);
and U42513 (N_42513,N_36655,N_36173);
nor U42514 (N_42514,N_36485,N_30230);
nand U42515 (N_42515,N_36098,N_30983);
or U42516 (N_42516,N_33620,N_33534);
nand U42517 (N_42517,N_37311,N_34699);
xnor U42518 (N_42518,N_31771,N_36560);
or U42519 (N_42519,N_36425,N_35093);
or U42520 (N_42520,N_37174,N_32674);
xor U42521 (N_42521,N_31319,N_39987);
nand U42522 (N_42522,N_35749,N_39530);
or U42523 (N_42523,N_34128,N_38679);
and U42524 (N_42524,N_35876,N_36464);
xor U42525 (N_42525,N_38793,N_32269);
and U42526 (N_42526,N_36329,N_37823);
nand U42527 (N_42527,N_34101,N_39942);
and U42528 (N_42528,N_38314,N_33843);
nand U42529 (N_42529,N_39857,N_32299);
nor U42530 (N_42530,N_39177,N_30347);
nand U42531 (N_42531,N_37888,N_30211);
and U42532 (N_42532,N_35045,N_37803);
or U42533 (N_42533,N_38363,N_35833);
nor U42534 (N_42534,N_37539,N_39316);
and U42535 (N_42535,N_35621,N_39587);
and U42536 (N_42536,N_35622,N_36222);
xnor U42537 (N_42537,N_30379,N_39147);
nor U42538 (N_42538,N_30066,N_32647);
xnor U42539 (N_42539,N_31033,N_30215);
nor U42540 (N_42540,N_36016,N_36444);
nor U42541 (N_42541,N_38870,N_30013);
or U42542 (N_42542,N_34327,N_33654);
xnor U42543 (N_42543,N_32433,N_39076);
nand U42544 (N_42544,N_32582,N_36753);
nor U42545 (N_42545,N_35090,N_33803);
or U42546 (N_42546,N_35320,N_37868);
nor U42547 (N_42547,N_39339,N_38627);
and U42548 (N_42548,N_33852,N_35745);
nand U42549 (N_42549,N_37661,N_31041);
and U42550 (N_42550,N_33521,N_38199);
or U42551 (N_42551,N_34502,N_35269);
nor U42552 (N_42552,N_31044,N_37371);
and U42553 (N_42553,N_36181,N_34139);
nor U42554 (N_42554,N_33540,N_37178);
nor U42555 (N_42555,N_35824,N_31441);
xor U42556 (N_42556,N_31800,N_38077);
and U42557 (N_42557,N_38559,N_30964);
or U42558 (N_42558,N_30254,N_37913);
xor U42559 (N_42559,N_32056,N_38858);
nor U42560 (N_42560,N_31301,N_34586);
nor U42561 (N_42561,N_39588,N_34106);
nand U42562 (N_42562,N_38682,N_32602);
xor U42563 (N_42563,N_31820,N_31356);
nor U42564 (N_42564,N_36186,N_38732);
nand U42565 (N_42565,N_32559,N_33714);
xnor U42566 (N_42566,N_31794,N_39097);
nand U42567 (N_42567,N_32037,N_36583);
nor U42568 (N_42568,N_39161,N_35881);
or U42569 (N_42569,N_33609,N_38850);
nand U42570 (N_42570,N_38508,N_35535);
or U42571 (N_42571,N_36600,N_38016);
and U42572 (N_42572,N_38520,N_38421);
xnor U42573 (N_42573,N_39429,N_35868);
or U42574 (N_42574,N_36283,N_37402);
nor U42575 (N_42575,N_38515,N_32553);
xnor U42576 (N_42576,N_31787,N_36858);
nand U42577 (N_42577,N_30786,N_37185);
nand U42578 (N_42578,N_36382,N_39184);
nand U42579 (N_42579,N_34062,N_38854);
xnor U42580 (N_42580,N_33826,N_32104);
nand U42581 (N_42581,N_33306,N_32579);
and U42582 (N_42582,N_34664,N_30034);
or U42583 (N_42583,N_39849,N_30405);
xor U42584 (N_42584,N_30881,N_33723);
xnor U42585 (N_42585,N_32861,N_37797);
or U42586 (N_42586,N_36080,N_34190);
nand U42587 (N_42587,N_34202,N_38166);
xor U42588 (N_42588,N_38862,N_39261);
xnor U42589 (N_42589,N_34474,N_32019);
and U42590 (N_42590,N_36153,N_37188);
nor U42591 (N_42591,N_37805,N_32790);
nand U42592 (N_42592,N_31163,N_37994);
nor U42593 (N_42593,N_37613,N_31914);
nor U42594 (N_42594,N_32164,N_30403);
xnor U42595 (N_42595,N_34109,N_31567);
xor U42596 (N_42596,N_30926,N_38346);
xnor U42597 (N_42597,N_33346,N_39597);
or U42598 (N_42598,N_35025,N_35059);
and U42599 (N_42599,N_33071,N_30422);
nor U42600 (N_42600,N_31947,N_39302);
or U42601 (N_42601,N_35513,N_38840);
nand U42602 (N_42602,N_30599,N_36135);
or U42603 (N_42603,N_35539,N_39026);
nand U42604 (N_42604,N_34482,N_39735);
xor U42605 (N_42605,N_33414,N_36225);
and U42606 (N_42606,N_38922,N_33225);
and U42607 (N_42607,N_32021,N_38865);
nor U42608 (N_42608,N_30871,N_38198);
and U42609 (N_42609,N_34928,N_37223);
nand U42610 (N_42610,N_37095,N_30261);
xnor U42611 (N_42611,N_32162,N_32339);
or U42612 (N_42612,N_32686,N_32008);
nor U42613 (N_42613,N_31206,N_35277);
nor U42614 (N_42614,N_31866,N_35173);
xor U42615 (N_42615,N_38595,N_38292);
nor U42616 (N_42616,N_37025,N_32910);
nor U42617 (N_42617,N_38500,N_38725);
nor U42618 (N_42618,N_32813,N_39190);
or U42619 (N_42619,N_39287,N_37320);
and U42620 (N_42620,N_30182,N_32205);
nand U42621 (N_42621,N_36694,N_39862);
nor U42622 (N_42622,N_39294,N_37807);
or U42623 (N_42623,N_30902,N_39596);
nand U42624 (N_42624,N_33079,N_30339);
nand U42625 (N_42625,N_33921,N_30514);
and U42626 (N_42626,N_30497,N_38344);
nor U42627 (N_42627,N_38058,N_35027);
xnor U42628 (N_42628,N_32659,N_31158);
and U42629 (N_42629,N_36851,N_38172);
and U42630 (N_42630,N_35462,N_35746);
xnor U42631 (N_42631,N_32278,N_35043);
and U42632 (N_42632,N_35079,N_38164);
nand U42633 (N_42633,N_31785,N_34203);
or U42634 (N_42634,N_34758,N_36476);
or U42635 (N_42635,N_36915,N_34277);
nor U42636 (N_42636,N_33947,N_38305);
and U42637 (N_42637,N_36854,N_32145);
or U42638 (N_42638,N_32472,N_36463);
nor U42639 (N_42639,N_35095,N_34986);
nor U42640 (N_42640,N_36730,N_34048);
xor U42641 (N_42641,N_31639,N_39758);
xnor U42642 (N_42642,N_39065,N_36981);
xnor U42643 (N_42643,N_34027,N_37434);
xnor U42644 (N_42644,N_36224,N_34666);
nand U42645 (N_42645,N_31454,N_33694);
nand U42646 (N_42646,N_37513,N_32256);
xor U42647 (N_42647,N_38531,N_31796);
nand U42648 (N_42648,N_32017,N_34514);
or U42649 (N_42649,N_39643,N_37578);
nor U42650 (N_42650,N_32464,N_37787);
nor U42651 (N_42651,N_34120,N_31069);
or U42652 (N_42652,N_31305,N_30512);
nor U42653 (N_42653,N_30281,N_31265);
xor U42654 (N_42654,N_38707,N_35807);
and U42655 (N_42655,N_33104,N_38418);
or U42656 (N_42656,N_39377,N_34761);
nand U42657 (N_42657,N_32507,N_37558);
nor U42658 (N_42658,N_34959,N_39292);
and U42659 (N_42659,N_36934,N_34419);
and U42660 (N_42660,N_31078,N_38968);
and U42661 (N_42661,N_38787,N_31636);
xor U42662 (N_42662,N_39362,N_37431);
xor U42663 (N_42663,N_30773,N_34650);
or U42664 (N_42664,N_35028,N_34525);
and U42665 (N_42665,N_37827,N_35614);
and U42666 (N_42666,N_39295,N_34251);
xor U42667 (N_42667,N_32630,N_30611);
or U42668 (N_42668,N_34008,N_32872);
nand U42669 (N_42669,N_30619,N_39747);
or U42670 (N_42670,N_30885,N_33058);
nor U42671 (N_42671,N_31928,N_31804);
nor U42672 (N_42672,N_37660,N_35987);
or U42673 (N_42673,N_33520,N_38599);
and U42674 (N_42674,N_36775,N_31089);
or U42675 (N_42675,N_33720,N_30009);
nor U42676 (N_42676,N_36142,N_38929);
xnor U42677 (N_42677,N_32653,N_39043);
nand U42678 (N_42678,N_30867,N_31012);
and U42679 (N_42679,N_31321,N_31119);
nand U42680 (N_42680,N_31581,N_35150);
or U42681 (N_42681,N_33405,N_34446);
nor U42682 (N_42682,N_34464,N_36762);
xor U42683 (N_42683,N_34732,N_34894);
or U42684 (N_42684,N_36348,N_34727);
nor U42685 (N_42685,N_37569,N_33113);
nor U42686 (N_42686,N_31755,N_39418);
or U42687 (N_42687,N_35863,N_36238);
xnor U42688 (N_42688,N_36474,N_31889);
or U42689 (N_42689,N_30617,N_31560);
and U42690 (N_42690,N_32817,N_34680);
xnor U42691 (N_42691,N_35926,N_37217);
nor U42692 (N_42692,N_37358,N_35645);
or U42693 (N_42693,N_37634,N_32552);
nor U42694 (N_42694,N_30470,N_30492);
xor U42695 (N_42695,N_39984,N_31237);
nand U42696 (N_42696,N_33822,N_37462);
and U42697 (N_42697,N_35217,N_38065);
nand U42698 (N_42698,N_37952,N_34888);
and U42699 (N_42699,N_30106,N_32213);
xor U42700 (N_42700,N_34023,N_32989);
or U42701 (N_42701,N_36387,N_38306);
xor U42702 (N_42702,N_38455,N_38326);
xor U42703 (N_42703,N_34782,N_31932);
and U42704 (N_42704,N_34418,N_34914);
nand U42705 (N_42705,N_30537,N_31097);
nor U42706 (N_42706,N_38226,N_37872);
nand U42707 (N_42707,N_38749,N_35264);
xor U42708 (N_42708,N_35762,N_32375);
and U42709 (N_42709,N_32604,N_38507);
xnor U42710 (N_42710,N_36940,N_39799);
or U42711 (N_42711,N_30686,N_33278);
nand U42712 (N_42712,N_39393,N_36902);
xor U42713 (N_42713,N_37652,N_34624);
and U42714 (N_42714,N_35879,N_34161);
and U42715 (N_42715,N_38995,N_31179);
and U42716 (N_42716,N_33840,N_31048);
nor U42717 (N_42717,N_34086,N_36212);
nand U42718 (N_42718,N_38461,N_35144);
nand U42719 (N_42719,N_32305,N_37085);
xor U42720 (N_42720,N_33325,N_38430);
nor U42721 (N_42721,N_36350,N_38796);
nor U42722 (N_42722,N_39645,N_34269);
and U42723 (N_42723,N_31027,N_34117);
and U42724 (N_42724,N_38697,N_31451);
xnor U42725 (N_42725,N_30912,N_30055);
and U42726 (N_42726,N_32231,N_32174);
nor U42727 (N_42727,N_37722,N_30320);
and U42728 (N_42728,N_37128,N_31023);
nand U42729 (N_42729,N_30383,N_39622);
nand U42730 (N_42730,N_36847,N_32777);
nor U42731 (N_42731,N_30040,N_34806);
nand U42732 (N_42732,N_32483,N_34632);
and U42733 (N_42733,N_32830,N_30794);
xor U42734 (N_42734,N_31756,N_35635);
or U42735 (N_42735,N_36893,N_39480);
xor U42736 (N_42736,N_36829,N_36535);
nor U42737 (N_42737,N_35548,N_34129);
nor U42738 (N_42738,N_30905,N_37978);
nor U42739 (N_42739,N_30956,N_37761);
nand U42740 (N_42740,N_31116,N_35270);
nand U42741 (N_42741,N_31939,N_32380);
and U42742 (N_42742,N_32526,N_32128);
nand U42743 (N_42743,N_30475,N_34445);
xor U42744 (N_42744,N_35176,N_38138);
nand U42745 (N_42745,N_34405,N_31168);
and U42746 (N_42746,N_31081,N_30868);
nor U42747 (N_42747,N_32055,N_30753);
or U42748 (N_42748,N_37624,N_32525);
xor U42749 (N_42749,N_36619,N_32839);
nand U42750 (N_42750,N_32978,N_32361);
or U42751 (N_42751,N_35343,N_31973);
and U42752 (N_42752,N_38753,N_30299);
and U42753 (N_42753,N_31072,N_39687);
and U42754 (N_42754,N_36456,N_36659);
or U42755 (N_42755,N_30880,N_35694);
and U42756 (N_42756,N_34762,N_37341);
xnor U42757 (N_42757,N_38006,N_35631);
nand U42758 (N_42758,N_30999,N_33222);
xor U42759 (N_42759,N_37836,N_31495);
nand U42760 (N_42760,N_32757,N_31920);
and U42761 (N_42761,N_34226,N_33589);
nand U42762 (N_42762,N_36180,N_35005);
nor U42763 (N_42763,N_33437,N_39337);
and U42764 (N_42764,N_36808,N_30270);
xnor U42765 (N_42765,N_37005,N_35140);
or U42766 (N_42766,N_35731,N_37076);
and U42767 (N_42767,N_34598,N_33063);
or U42768 (N_42768,N_32721,N_32331);
nand U42769 (N_42769,N_37212,N_33484);
and U42770 (N_42770,N_37974,N_34463);
nand U42771 (N_42771,N_31313,N_30125);
and U42772 (N_42772,N_32342,N_37916);
xor U42773 (N_42773,N_35898,N_30948);
and U42774 (N_42774,N_37047,N_37502);
nor U42775 (N_42775,N_32986,N_34990);
nand U42776 (N_42776,N_34656,N_37700);
and U42777 (N_42777,N_38214,N_38200);
nor U42778 (N_42778,N_33612,N_30473);
or U42779 (N_42779,N_30207,N_36388);
nor U42780 (N_42780,N_36293,N_35451);
nand U42781 (N_42781,N_34223,N_36357);
xor U42782 (N_42782,N_30523,N_36814);
nand U42783 (N_42783,N_36977,N_32006);
xnor U42784 (N_42784,N_32561,N_38528);
nor U42785 (N_42785,N_36048,N_37390);
and U42786 (N_42786,N_37619,N_31526);
nand U42787 (N_42787,N_37738,N_31585);
nand U42788 (N_42788,N_35497,N_33264);
nor U42789 (N_42789,N_31209,N_30062);
or U42790 (N_42790,N_31959,N_32982);
xnor U42791 (N_42791,N_34933,N_39728);
and U42792 (N_42792,N_38007,N_37144);
or U42793 (N_42793,N_35891,N_36219);
or U42794 (N_42794,N_38004,N_32974);
nand U42795 (N_42795,N_30911,N_33455);
or U42796 (N_42796,N_32937,N_38875);
and U42797 (N_42797,N_32293,N_34784);
or U42798 (N_42798,N_31344,N_39458);
nor U42799 (N_42799,N_37789,N_36150);
nor U42800 (N_42800,N_39395,N_34898);
and U42801 (N_42801,N_39151,N_37854);
nand U42802 (N_42802,N_37012,N_33625);
nor U42803 (N_42803,N_39508,N_32847);
xnor U42804 (N_42804,N_34930,N_34363);
xor U42805 (N_42805,N_34233,N_34879);
and U42806 (N_42806,N_35399,N_33887);
nor U42807 (N_42807,N_32382,N_30882);
and U42808 (N_42808,N_34091,N_35312);
nand U42809 (N_42809,N_37833,N_34833);
and U42810 (N_42810,N_31059,N_31555);
nand U42811 (N_42811,N_39146,N_30031);
nand U42812 (N_42812,N_36461,N_35102);
xnor U42813 (N_42813,N_39804,N_35812);
nand U42814 (N_42814,N_37309,N_32589);
and U42815 (N_42815,N_33025,N_32317);
nor U42816 (N_42816,N_37122,N_32836);
nand U42817 (N_42817,N_30727,N_32144);
or U42818 (N_42818,N_37086,N_38328);
xor U42819 (N_42819,N_37275,N_37673);
and U42820 (N_42820,N_31333,N_38906);
nand U42821 (N_42821,N_39071,N_37577);
nand U42822 (N_42822,N_37248,N_39394);
nand U42823 (N_42823,N_37906,N_31182);
nor U42824 (N_42824,N_38583,N_36042);
xor U42825 (N_42825,N_35504,N_34134);
xor U42826 (N_42826,N_31708,N_33518);
and U42827 (N_42827,N_31436,N_34742);
nor U42828 (N_42828,N_30056,N_39801);
nor U42829 (N_42829,N_31425,N_36906);
nand U42830 (N_42830,N_38876,N_37067);
xnor U42831 (N_42831,N_39004,N_35428);
xor U42832 (N_42832,N_31824,N_33011);
nand U42833 (N_42833,N_36160,N_30634);
or U42834 (N_42834,N_38819,N_32451);
nor U42835 (N_42835,N_31518,N_35553);
nor U42836 (N_42836,N_39673,N_30284);
nand U42837 (N_42837,N_32116,N_30003);
xor U42838 (N_42838,N_30630,N_38002);
xnor U42839 (N_42839,N_38900,N_33286);
xor U42840 (N_42840,N_34572,N_37075);
xnor U42841 (N_42841,N_32651,N_33563);
nor U42842 (N_42842,N_37733,N_33873);
nor U42843 (N_42843,N_33846,N_37287);
nand U42844 (N_42844,N_32432,N_37848);
or U42845 (N_42845,N_33474,N_39502);
or U42846 (N_42846,N_39781,N_36662);
and U42847 (N_42847,N_30167,N_36267);
nand U42848 (N_42848,N_33550,N_30710);
nor U42849 (N_42849,N_31790,N_38209);
and U42850 (N_42850,N_37886,N_38881);
xor U42851 (N_42851,N_37292,N_34313);
nor U42852 (N_42852,N_30839,N_35922);
xnor U42853 (N_42853,N_37936,N_31498);
or U42854 (N_42854,N_34093,N_39732);
or U42855 (N_42855,N_31464,N_32635);
and U42856 (N_42856,N_31476,N_35050);
nor U42857 (N_42857,N_36832,N_39606);
nand U42858 (N_42858,N_31221,N_39780);
nand U42859 (N_42859,N_37041,N_35480);
xnor U42860 (N_42860,N_33201,N_33691);
nand U42861 (N_42861,N_39056,N_36462);
nor U42862 (N_42862,N_31291,N_38303);
xnor U42863 (N_42863,N_34849,N_38905);
or U42864 (N_42864,N_37141,N_36379);
nand U42865 (N_42865,N_38781,N_30000);
nor U42866 (N_42866,N_37999,N_31004);
nor U42867 (N_42867,N_33391,N_33937);
or U42868 (N_42868,N_32049,N_39970);
xor U42869 (N_42869,N_37792,N_36428);
nand U42870 (N_42870,N_36316,N_34793);
xnor U42871 (N_42871,N_34430,N_36046);
or U42872 (N_42872,N_32701,N_33359);
or U42873 (N_42873,N_34478,N_33239);
or U42874 (N_42874,N_31677,N_38117);
nand U42875 (N_42875,N_34479,N_36949);
nor U42876 (N_42876,N_38148,N_36223);
and U42877 (N_42877,N_37049,N_34840);
xnor U42878 (N_42878,N_37930,N_37265);
nor U42879 (N_42879,N_37924,N_34583);
or U42880 (N_42880,N_35274,N_37687);
nor U42881 (N_42881,N_35977,N_33964);
nor U42882 (N_42882,N_38073,N_32504);
nor U42883 (N_42883,N_38666,N_33737);
xor U42884 (N_42884,N_37021,N_31611);
and U42885 (N_42885,N_37768,N_38260);
nand U42886 (N_42886,N_36067,N_39766);
nor U42887 (N_42887,N_31127,N_38008);
xor U42888 (N_42888,N_30399,N_39586);
nand U42889 (N_42889,N_32556,N_38879);
and U42890 (N_42890,N_30402,N_33958);
or U42891 (N_42891,N_34493,N_35240);
nand U42892 (N_42892,N_37487,N_32158);
and U42893 (N_42893,N_34253,N_31830);
or U42894 (N_42894,N_34192,N_39113);
nand U42895 (N_42895,N_37646,N_31919);
nor U42896 (N_42896,N_32308,N_30209);
or U42897 (N_42897,N_35326,N_36232);
xor U42898 (N_42898,N_36884,N_38722);
xnor U42899 (N_42899,N_31681,N_34867);
nand U42900 (N_42900,N_38357,N_35950);
and U42901 (N_42901,N_31852,N_35098);
nand U42902 (N_42902,N_33353,N_30676);
and U42903 (N_42903,N_39032,N_35902);
xor U42904 (N_42904,N_35537,N_37351);
and U42905 (N_42905,N_30090,N_39135);
xnor U42906 (N_42906,N_30162,N_30525);
nand U42907 (N_42907,N_34708,N_33678);
or U42908 (N_42908,N_34967,N_39471);
nand U42909 (N_42909,N_31546,N_34804);
or U42910 (N_42910,N_37463,N_38554);
nor U42911 (N_42911,N_37982,N_32364);
nor U42912 (N_42912,N_34200,N_34016);
or U42913 (N_42913,N_37154,N_34425);
nand U42914 (N_42914,N_32891,N_36782);
or U42915 (N_42915,N_39543,N_32173);
or U42916 (N_42916,N_34015,N_33232);
nand U42917 (N_42917,N_32014,N_30459);
and U42918 (N_42918,N_34484,N_30960);
or U42919 (N_42919,N_36294,N_32779);
nor U42920 (N_42920,N_34118,N_31988);
nand U42921 (N_42921,N_35177,N_32879);
xnor U42922 (N_42922,N_35842,N_38331);
and U42923 (N_42923,N_39467,N_39601);
nand U42924 (N_42924,N_32925,N_34466);
nor U42925 (N_42925,N_32294,N_36658);
or U42926 (N_42926,N_37405,N_31306);
nand U42927 (N_42927,N_30545,N_32774);
nor U42928 (N_42928,N_39130,N_35297);
xnor U42929 (N_42929,N_32524,N_34092);
xor U42930 (N_42930,N_33146,N_30318);
xor U42931 (N_42931,N_34395,N_34822);
nand U42932 (N_42932,N_37629,N_31140);
or U42933 (N_42933,N_35971,N_32260);
xnor U42934 (N_42934,N_32565,N_32612);
nand U42935 (N_42935,N_37655,N_35930);
xnor U42936 (N_42936,N_36701,N_31211);
nand U42937 (N_42937,N_30115,N_32959);
nand U42938 (N_42938,N_36002,N_30220);
nand U42939 (N_42939,N_36946,N_35962);
nor U42940 (N_42940,N_31961,N_32709);
nor U42941 (N_42941,N_38867,N_37701);
or U42942 (N_42942,N_37884,N_36404);
nor U42943 (N_42943,N_30250,N_30183);
xor U42944 (N_42944,N_33583,N_39437);
nand U42945 (N_42945,N_36975,N_33785);
nand U42946 (N_42946,N_38712,N_35502);
xnor U42947 (N_42947,N_30929,N_37961);
or U42948 (N_42948,N_35209,N_36011);
nor U42949 (N_42949,N_36076,N_31009);
nor U42950 (N_42950,N_35124,N_30937);
xnor U42951 (N_42951,N_38123,N_34657);
nor U42952 (N_42952,N_35146,N_32222);
xnor U42953 (N_42953,N_31461,N_30432);
xnor U42954 (N_42954,N_36856,N_31156);
nor U42955 (N_42955,N_39904,N_38978);
or U42956 (N_42956,N_36962,N_38310);
nand U42957 (N_42957,N_36802,N_37045);
and U42958 (N_42958,N_38578,N_33816);
nor U42959 (N_42959,N_37609,N_35477);
or U42960 (N_42960,N_31274,N_33656);
or U42961 (N_42961,N_30091,N_39729);
xor U42962 (N_42962,N_30748,N_39322);
and U42963 (N_42963,N_38934,N_39077);
xnor U42964 (N_42964,N_36876,N_30338);
nand U42965 (N_42965,N_33979,N_34785);
or U42966 (N_42966,N_32273,N_31777);
nand U42967 (N_42967,N_31599,N_31882);
xnor U42968 (N_42968,N_37898,N_35867);
nor U42969 (N_42969,N_34733,N_32585);
xnor U42970 (N_42970,N_33501,N_30759);
nor U42971 (N_42971,N_34121,N_34187);
xnor U42972 (N_42972,N_39896,N_37719);
and U42973 (N_42973,N_38470,N_32866);
nand U42974 (N_42974,N_32725,N_32135);
nor U42975 (N_42975,N_30841,N_38539);
nor U42976 (N_42976,N_30894,N_39819);
or U42977 (N_42977,N_39655,N_34686);
or U42978 (N_42978,N_39134,N_34748);
or U42979 (N_42979,N_33229,N_38419);
nand U42980 (N_42980,N_35284,N_30134);
nand U42981 (N_42981,N_30834,N_39978);
xor U42982 (N_42982,N_35666,N_36380);
or U42983 (N_42983,N_39459,N_34285);
or U42984 (N_42984,N_39399,N_37119);
nand U42985 (N_42985,N_38275,N_36084);
nor U42986 (N_42986,N_33265,N_34141);
nor U42987 (N_42987,N_37500,N_35367);
xnor U42988 (N_42988,N_37096,N_39763);
xor U42989 (N_42989,N_33760,N_35244);
and U42990 (N_42990,N_36568,N_39992);
and U42991 (N_42991,N_37250,N_36761);
nor U42992 (N_42992,N_31043,N_39812);
or U42993 (N_42993,N_32663,N_35753);
xor U42994 (N_42994,N_33781,N_30139);
and U42995 (N_42995,N_39855,N_36157);
and U42996 (N_42996,N_31684,N_38391);
or U42997 (N_42997,N_37568,N_34343);
or U42998 (N_42998,N_33149,N_33652);
xor U42999 (N_42999,N_33903,N_32024);
nor U43000 (N_43000,N_34477,N_36506);
nand U43001 (N_43001,N_38687,N_39805);
nor U43002 (N_43002,N_31623,N_31534);
and U43003 (N_43003,N_38565,N_32066);
nor U43004 (N_43004,N_35814,N_31251);
xnor U43005 (N_43005,N_37838,N_32156);
nand U43006 (N_43006,N_34969,N_34634);
nand U43007 (N_43007,N_34237,N_36720);
or U43008 (N_43008,N_30024,N_38368);
nor U43009 (N_43009,N_37935,N_36028);
or U43010 (N_43010,N_32537,N_35117);
nand U43011 (N_43011,N_36230,N_31499);
nor U43012 (N_43012,N_34880,N_37885);
nor U43013 (N_43013,N_37241,N_30988);
nand U43014 (N_43014,N_37196,N_34408);
or U43015 (N_43015,N_30663,N_39259);
or U43016 (N_43016,N_35784,N_30436);
xnor U43017 (N_43017,N_39526,N_37408);
xor U43018 (N_43018,N_31726,N_31941);
and U43019 (N_43019,N_37181,N_38047);
nand U43020 (N_43020,N_31216,N_32988);
nor U43021 (N_43021,N_38278,N_34231);
xnor U43022 (N_43022,N_34808,N_31015);
xor U43023 (N_43023,N_31067,N_30122);
and U43024 (N_43024,N_38790,N_34550);
xor U43025 (N_43025,N_30324,N_35561);
and U43026 (N_43026,N_36385,N_34310);
nor U43027 (N_43027,N_34595,N_32189);
xnor U43028 (N_43028,N_31062,N_33961);
nor U43029 (N_43029,N_37457,N_36393);
nand U43030 (N_43030,N_31330,N_34941);
and U43031 (N_43031,N_38393,N_35374);
or U43032 (N_43032,N_35411,N_38871);
nor U43033 (N_43033,N_34165,N_32323);
nand U43034 (N_43034,N_32038,N_32152);
xor U43035 (N_43035,N_33076,N_39951);
or U43036 (N_43036,N_35171,N_33084);
nor U43037 (N_43037,N_39353,N_31022);
xnor U43038 (N_43038,N_33568,N_37160);
nor U43039 (N_43039,N_38638,N_38891);
and U43040 (N_43040,N_38319,N_35442);
nand U43041 (N_43041,N_39357,N_39932);
or U43042 (N_43042,N_37115,N_30389);
and U43043 (N_43043,N_36841,N_33178);
or U43044 (N_43044,N_33780,N_32683);
nand U43045 (N_43045,N_39604,N_38364);
xor U43046 (N_43046,N_32778,N_30751);
and U43047 (N_43047,N_31035,N_32522);
xor U43048 (N_43048,N_38446,N_32735);
xnor U43049 (N_43049,N_35638,N_30752);
and U43050 (N_43050,N_36541,N_30482);
nor U43051 (N_43051,N_31497,N_34302);
or U43052 (N_43052,N_35729,N_36266);
and U43053 (N_43053,N_30503,N_32058);
xor U43054 (N_43054,N_35299,N_37013);
nor U43055 (N_43055,N_39501,N_33398);
xor U43056 (N_43056,N_39566,N_38821);
xor U43057 (N_43057,N_32076,N_37989);
nand U43058 (N_43058,N_37003,N_39392);
nand U43059 (N_43059,N_35237,N_31471);
nor U43060 (N_43060,N_34083,N_37272);
or U43061 (N_43061,N_34705,N_30321);
and U43062 (N_43062,N_30872,N_39625);
nand U43063 (N_43063,N_35790,N_30373);
nand U43064 (N_43064,N_30524,N_39724);
nor U43065 (N_43065,N_33361,N_37316);
nor U43066 (N_43066,N_32068,N_39001);
nand U43067 (N_43067,N_38465,N_37052);
xor U43068 (N_43068,N_31982,N_37106);
nand U43069 (N_43069,N_34356,N_33198);
xnor U43070 (N_43070,N_32763,N_33145);
nand U43071 (N_43071,N_32634,N_36161);
nor U43072 (N_43072,N_31981,N_34786);
or U43073 (N_43073,N_33716,N_38884);
nand U43074 (N_43074,N_32523,N_30959);
or U43075 (N_43075,N_30817,N_38923);
nand U43076 (N_43076,N_33897,N_34351);
and U43077 (N_43077,N_36922,N_32564);
nor U43078 (N_43078,N_38304,N_36116);
nand U43079 (N_43079,N_33314,N_30863);
xor U43080 (N_43080,N_32529,N_38051);
nor U43081 (N_43081,N_36576,N_34455);
and U43082 (N_43082,N_36942,N_32400);
or U43083 (N_43083,N_33189,N_36888);
or U43084 (N_43084,N_32099,N_36635);
nand U43085 (N_43085,N_31066,N_33155);
or U43086 (N_43086,N_30161,N_39617);
xor U43087 (N_43087,N_30583,N_39400);
xnor U43088 (N_43088,N_31933,N_34892);
and U43089 (N_43089,N_33730,N_36203);
nor U43090 (N_43090,N_34764,N_32234);
xnor U43091 (N_43091,N_37454,N_37008);
nand U43092 (N_43092,N_33467,N_35489);
xnor U43093 (N_43093,N_37083,N_37562);
and U43094 (N_43094,N_39226,N_33847);
nand U43095 (N_43095,N_31724,N_33432);
and U43096 (N_43096,N_37877,N_39934);
or U43097 (N_43097,N_32439,N_38949);
and U43098 (N_43098,N_35366,N_34305);
xor U43099 (N_43099,N_32895,N_34504);
nand U43100 (N_43100,N_36207,N_33697);
nand U43101 (N_43101,N_39013,N_32905);
nor U43102 (N_43102,N_31858,N_31763);
or U43103 (N_43103,N_33806,N_34001);
xnor U43104 (N_43104,N_39126,N_38247);
and U43105 (N_43105,N_35764,N_30985);
xor U43106 (N_43106,N_32638,N_36213);
xor U43107 (N_43107,N_39366,N_34770);
and U43108 (N_43108,N_39685,N_34744);
or U43109 (N_43109,N_31997,N_37231);
or U43110 (N_43110,N_34862,N_34668);
nand U43111 (N_43111,N_38263,N_30350);
or U43112 (N_43112,N_37035,N_31937);
nand U43113 (N_43113,N_33053,N_36320);
or U43114 (N_43114,N_36020,N_31936);
or U43115 (N_43115,N_34963,N_38385);
nand U43116 (N_43116,N_33098,N_31596);
and U43117 (N_43117,N_35989,N_36627);
nand U43118 (N_43118,N_30385,N_34228);
or U43119 (N_43119,N_34158,N_35998);
xnor U43120 (N_43120,N_36314,N_36012);
xor U43121 (N_43121,N_36480,N_33135);
nor U43122 (N_43122,N_33943,N_39329);
nor U43123 (N_43123,N_30659,N_31257);
xor U43124 (N_43124,N_37992,N_35769);
nor U43125 (N_43125,N_35167,N_33538);
or U43126 (N_43126,N_33419,N_37491);
xnor U43127 (N_43127,N_32474,N_37769);
nand U43128 (N_43128,N_33094,N_37493);
xor U43129 (N_43129,N_39548,N_33515);
nor U43130 (N_43130,N_30802,N_34876);
and U43131 (N_43131,N_30458,N_35937);
nor U43132 (N_43132,N_36572,N_35592);
nor U43133 (N_43133,N_36695,N_34244);
or U43134 (N_43134,N_36466,N_30008);
or U43135 (N_43135,N_37840,N_35106);
and U43136 (N_43136,N_33991,N_32970);
xnor U43137 (N_43137,N_31819,N_33446);
and U43138 (N_43138,N_33946,N_31037);
or U43139 (N_43139,N_34170,N_30942);
xnor U43140 (N_43140,N_30536,N_37565);
nand U43141 (N_43141,N_36537,N_32732);
and U43142 (N_43142,N_32887,N_32487);
nand U43143 (N_43143,N_35057,N_35400);
or U43144 (N_43144,N_30673,N_37082);
xor U43145 (N_43145,N_33523,N_38609);
and U43146 (N_43146,N_38632,N_37657);
nand U43147 (N_43147,N_30864,N_35780);
nand U43148 (N_43148,N_36660,N_39656);
or U43149 (N_43149,N_36101,N_37165);
and U43150 (N_43150,N_36496,N_34236);
nand U43151 (N_43151,N_30252,N_36376);
and U43152 (N_43152,N_30141,N_39525);
or U43153 (N_43153,N_39428,N_31445);
nand U43154 (N_43154,N_32606,N_34412);
or U43155 (N_43155,N_36668,N_37839);
xor U43156 (N_43156,N_35052,N_34985);
and U43157 (N_43157,N_39389,N_33804);
or U43158 (N_43158,N_30017,N_32186);
nand U43159 (N_43159,N_37882,N_30177);
xor U43160 (N_43160,N_34643,N_39441);
or U43161 (N_43161,N_36591,N_30674);
nand U43162 (N_43162,N_35516,N_33163);
nand U43163 (N_43163,N_31699,N_33881);
nor U43164 (N_43164,N_33801,N_33039);
or U43165 (N_43165,N_34102,N_37746);
and U43166 (N_43166,N_35472,N_35577);
and U43167 (N_43167,N_34693,N_33193);
or U43168 (N_43168,N_39807,N_35917);
or U43169 (N_43169,N_36465,N_31218);
or U43170 (N_43170,N_37488,N_39070);
xnor U43171 (N_43171,N_30033,N_39506);
xor U43172 (N_43172,N_38447,N_33406);
nand U43173 (N_43173,N_34582,N_36047);
and U43174 (N_43174,N_36813,N_34096);
and U43175 (N_43175,N_30498,N_33157);
or U43176 (N_43176,N_30953,N_36617);
xor U43177 (N_43177,N_31624,N_31397);
and U43178 (N_43178,N_37990,N_31845);
nand U43179 (N_43179,N_35721,N_31946);
and U43180 (N_43180,N_37461,N_30559);
and U43181 (N_43181,N_39279,N_38993);
xnor U43182 (N_43182,N_37069,N_38183);
xnor U43183 (N_43183,N_36974,N_38647);
or U43184 (N_43184,N_35928,N_34344);
xor U43185 (N_43185,N_38894,N_39524);
nor U43186 (N_43186,N_31248,N_39764);
nand U43187 (N_43187,N_31645,N_35768);
nor U43188 (N_43188,N_38959,N_35732);
nor U43189 (N_43189,N_38994,N_30243);
or U43190 (N_43190,N_32811,N_30043);
and U43191 (N_43191,N_38853,N_32801);
and U43192 (N_43192,N_35311,N_37219);
nand U43193 (N_43193,N_32063,N_37459);
xor U43194 (N_43194,N_30332,N_32922);
nor U43195 (N_43195,N_32242,N_37414);
nor U43196 (N_43196,N_37692,N_37148);
nor U43197 (N_43197,N_32201,N_39465);
xnor U43198 (N_43198,N_34638,N_30065);
and U43199 (N_43199,N_39396,N_39092);
or U43200 (N_43200,N_33855,N_36911);
nand U43201 (N_43201,N_38897,N_33525);
nand U43202 (N_43202,N_35742,N_31393);
and U43203 (N_43203,N_39694,N_38141);
nor U43204 (N_43204,N_37310,N_34013);
nor U43205 (N_43205,N_34903,N_33333);
nand U43206 (N_43206,N_35526,N_30306);
nor U43207 (N_43207,N_37763,N_37189);
and U43208 (N_43208,N_35524,N_34467);
nand U43209 (N_43209,N_33228,N_39388);
and U43210 (N_43210,N_36614,N_30856);
xnor U43211 (N_43211,N_31105,N_34697);
xor U43212 (N_43212,N_35899,N_38766);
or U43213 (N_43213,N_38136,N_33335);
and U43214 (N_43214,N_32180,N_35155);
xor U43215 (N_43215,N_35303,N_33088);
and U43216 (N_43216,N_30815,N_30873);
nor U43217 (N_43217,N_33779,N_32646);
and U43218 (N_43218,N_35816,N_36119);
and U43219 (N_43219,N_33131,N_35718);
or U43220 (N_43220,N_37394,N_33829);
or U43221 (N_43221,N_30568,N_31254);
and U43222 (N_43222,N_38129,N_39231);
xnor U43223 (N_43223,N_38156,N_33047);
or U43224 (N_43224,N_31282,N_38053);
or U43225 (N_43225,N_32263,N_32314);
xnor U43226 (N_43226,N_38495,N_30342);
nor U43227 (N_43227,N_36353,N_31195);
and U43228 (N_43228,N_30933,N_35820);
xor U43229 (N_43229,N_39964,N_35813);
and U43230 (N_43230,N_35736,N_39141);
or U43231 (N_43231,N_31587,N_39030);
or U43232 (N_43232,N_34003,N_34257);
nor U43233 (N_43233,N_34082,N_30632);
and U43234 (N_43234,N_30282,N_32661);
nand U43235 (N_43235,N_35558,N_34041);
nand U43236 (N_43236,N_31562,N_32783);
and U43237 (N_43237,N_33754,N_36507);
nand U43238 (N_43238,N_34088,N_35082);
nor U43239 (N_43239,N_34132,N_30779);
or U43240 (N_43240,N_36351,N_36715);
or U43241 (N_43241,N_31916,N_36432);
xnor U43242 (N_43242,N_32079,N_30833);
and U43243 (N_43243,N_31276,N_31327);
nor U43244 (N_43244,N_32551,N_34767);
nor U43245 (N_43245,N_34621,N_32652);
nor U43246 (N_43246,N_33137,N_35249);
or U43247 (N_43247,N_31825,N_35008);
and U43248 (N_43248,N_34449,N_38440);
xnor U43249 (N_43249,N_37420,N_30255);
or U43250 (N_43250,N_37226,N_33542);
xnor U43251 (N_43251,N_30755,N_39879);
nor U43252 (N_43252,N_39653,N_36246);
and U43253 (N_43253,N_31799,N_35434);
or U43254 (N_43254,N_39272,N_34578);
nor U43255 (N_43255,N_36395,N_32673);
nor U43256 (N_43256,N_36342,N_37929);
or U43257 (N_43257,N_34376,N_37177);
and U43258 (N_43258,N_33831,N_34126);
or U43259 (N_43259,N_34646,N_36721);
and U43260 (N_43260,N_35885,N_30421);
nand U43261 (N_43261,N_35860,N_33765);
and U43262 (N_43262,N_37385,N_38951);
or U43263 (N_43263,N_31449,N_35310);
or U43264 (N_43264,N_37981,N_31442);
nor U43265 (N_43265,N_38170,N_36154);
nor U43266 (N_43266,N_32284,N_31003);
and U43267 (N_43267,N_35030,N_39768);
or U43268 (N_43268,N_34037,N_36816);
nand U43269 (N_43269,N_36454,N_35964);
and U43270 (N_43270,N_35552,N_38325);
xnor U43271 (N_43271,N_36584,N_31529);
nor U43272 (N_43272,N_38576,N_36075);
or U43273 (N_43273,N_30934,N_37590);
nand U43274 (N_43274,N_34348,N_32327);
and U43275 (N_43275,N_35242,N_39315);
nor U43276 (N_43276,N_30440,N_30977);
or U43277 (N_43277,N_35520,N_36815);
or U43278 (N_43278,N_31691,N_31911);
or U43279 (N_43279,N_30467,N_39986);
nor U43280 (N_43280,N_30921,N_35097);
and U43281 (N_43281,N_30943,N_31432);
and U43282 (N_43282,N_35420,N_32983);
nor U43283 (N_43283,N_37479,N_35418);
or U43284 (N_43284,N_33407,N_37844);
nor U43285 (N_43285,N_39686,N_32111);
or U43286 (N_43286,N_30526,N_35965);
and U43287 (N_43287,N_30626,N_35735);
nand U43288 (N_43288,N_32398,N_37441);
xor U43289 (N_43289,N_38575,N_34913);
nor U43290 (N_43290,N_37009,N_31648);
and U43291 (N_43291,N_33594,N_35068);
and U43292 (N_43292,N_33073,N_33744);
nand U43293 (N_43293,N_35616,N_35172);
and U43294 (N_43294,N_31758,N_39517);
xor U43295 (N_43295,N_34034,N_39576);
nor U43296 (N_43296,N_34295,N_34991);
and U43297 (N_43297,N_36755,N_39037);
nand U43298 (N_43298,N_39603,N_30227);
xor U43299 (N_43299,N_31650,N_31521);
xor U43300 (N_43300,N_35953,N_32027);
xnor U43301 (N_43301,N_36810,N_30200);
nor U43302 (N_43302,N_37757,N_37580);
xor U43303 (N_43303,N_32387,N_37081);
or U43304 (N_43304,N_32220,N_30510);
nand U43305 (N_43305,N_33438,N_37688);
and U43306 (N_43306,N_34599,N_36746);
nand U43307 (N_43307,N_38510,N_38902);
and U43308 (N_43308,N_33480,N_35973);
or U43309 (N_43309,N_35453,N_32555);
nor U43310 (N_43310,N_39431,N_35559);
xnor U43311 (N_43311,N_38090,N_31710);
xor U43312 (N_43312,N_30232,N_37965);
and U43313 (N_43313,N_32761,N_32208);
or U43314 (N_43314,N_34531,N_32672);
nand U43315 (N_43315,N_37225,N_36304);
nand U43316 (N_43316,N_31674,N_34828);
or U43317 (N_43317,N_32112,N_35848);
or U43318 (N_43318,N_39120,N_36941);
nor U43319 (N_43319,N_31812,N_35308);
or U43320 (N_43320,N_31372,N_39317);
or U43321 (N_43321,N_39284,N_36299);
nand U43322 (N_43322,N_32291,N_31553);
nor U43323 (N_43323,N_33860,N_35107);
nor U43324 (N_43324,N_33557,N_39081);
xnor U43325 (N_43325,N_30005,N_35505);
nor U43326 (N_43326,N_30063,N_32911);
and U43327 (N_43327,N_30168,N_33362);
and U43328 (N_43328,N_39783,N_30098);
xor U43329 (N_43329,N_34989,N_38908);
or U43330 (N_43330,N_32086,N_30606);
xnor U43331 (N_43331,N_37669,N_32603);
or U43332 (N_43332,N_39880,N_36734);
nor U43333 (N_43333,N_33952,N_38213);
or U43334 (N_43334,N_36639,N_36227);
nor U43335 (N_43335,N_30274,N_34780);
nor U43336 (N_43336,N_32948,N_39067);
or U43337 (N_43337,N_31705,N_30039);
nand U43338 (N_43338,N_34997,N_36112);
and U43339 (N_43339,N_36823,N_32157);
or U43340 (N_43340,N_34893,N_33281);
nor U43341 (N_43341,N_37065,N_30175);
or U43342 (N_43342,N_39296,N_31834);
xnor U43343 (N_43343,N_39538,N_33403);
or U43344 (N_43344,N_37593,N_33436);
nor U43345 (N_43345,N_36943,N_31741);
or U43346 (N_43346,N_34508,N_33186);
nand U43347 (N_43347,N_39191,N_37473);
and U43348 (N_43348,N_33819,N_38792);
nand U43349 (N_43349,N_32882,N_30909);
nor U43350 (N_43350,N_34838,N_31383);
xnor U43351 (N_43351,N_36531,N_39714);
nand U43352 (N_43352,N_37446,N_32105);
and U43353 (N_43353,N_31170,N_36650);
nor U43354 (N_43354,N_34451,N_34340);
nand U43355 (N_43355,N_37818,N_35469);
xor U43356 (N_43356,N_30935,N_31874);
nand U43357 (N_43357,N_31138,N_35201);
nor U43358 (N_43358,N_32734,N_30425);
nand U43359 (N_43359,N_37811,N_31757);
nand U43360 (N_43360,N_39778,N_34193);
xor U43361 (N_43361,N_36437,N_38543);
nor U43362 (N_43362,N_38118,N_30870);
xor U43363 (N_43363,N_35938,N_35578);
and U43364 (N_43364,N_33481,N_38367);
or U43365 (N_43365,N_32011,N_39627);
nor U43366 (N_43366,N_31320,N_38104);
or U43367 (N_43367,N_30319,N_39927);
and U43368 (N_43368,N_30297,N_38064);
nor U43369 (N_43369,N_38652,N_38095);
nand U43370 (N_43370,N_36159,N_38813);
and U43371 (N_43371,N_33603,N_31474);
nand U43372 (N_43372,N_37411,N_38228);
and U43373 (N_43373,N_36092,N_30925);
and U43374 (N_43374,N_34915,N_37852);
nand U43375 (N_43375,N_36117,N_36930);
or U43376 (N_43376,N_38518,N_35959);
or U43377 (N_43377,N_34063,N_30069);
or U43378 (N_43378,N_30456,N_34523);
nor U43379 (N_43379,N_33416,N_34299);
nand U43380 (N_43380,N_37417,N_35445);
and U43381 (N_43381,N_33323,N_36054);
and U43382 (N_43382,N_34492,N_32792);
xnor U43383 (N_43383,N_37595,N_30099);
nor U43384 (N_43384,N_32172,N_39636);
nor U43385 (N_43385,N_37011,N_35267);
or U43386 (N_43386,N_33430,N_33517);
xnor U43387 (N_43387,N_37214,N_32515);
nor U43388 (N_43388,N_33431,N_30112);
or U43389 (N_43389,N_32707,N_35574);
and U43390 (N_43390,N_30835,N_31200);
nand U43391 (N_43391,N_39827,N_30472);
nand U43392 (N_43392,N_33751,N_35120);
or U43393 (N_43393,N_37187,N_31675);
nand U43394 (N_43394,N_30615,N_36264);
and U43395 (N_43395,N_36163,N_33505);
and U43396 (N_43396,N_36554,N_32773);
or U43397 (N_43397,N_33077,N_34662);
xor U43398 (N_43398,N_30750,N_32876);
or U43399 (N_43399,N_36199,N_33119);
nor U43400 (N_43400,N_31958,N_35603);
or U43401 (N_43401,N_36009,N_35212);
or U43402 (N_43402,N_32649,N_39490);
nor U43403 (N_43403,N_30486,N_39628);
and U43404 (N_43404,N_33896,N_31414);
nand U43405 (N_43405,N_37103,N_35427);
and U43406 (N_43406,N_38458,N_30080);
and U43407 (N_43407,N_33891,N_36475);
nand U43408 (N_43408,N_32671,N_33514);
and U43409 (N_43409,N_33016,N_35929);
nand U43410 (N_43410,N_36787,N_38398);
and U43411 (N_43411,N_36200,N_33700);
xor U43412 (N_43412,N_34125,N_39038);
xnor U43413 (N_43413,N_36391,N_35610);
and U43414 (N_43414,N_38960,N_30116);
and U43415 (N_43415,N_36765,N_35826);
and U43416 (N_43416,N_37186,N_39369);
nor U43417 (N_43417,N_30746,N_30414);
or U43418 (N_43418,N_34401,N_38102);
nor U43419 (N_43419,N_36511,N_30268);
and U43420 (N_43420,N_30454,N_33052);
or U43421 (N_43421,N_30495,N_31460);
or U43422 (N_43422,N_36332,N_32246);
or U43423 (N_43423,N_34654,N_35407);
or U43424 (N_43424,N_30754,N_35844);
xor U43425 (N_43425,N_33034,N_36210);
nor U43426 (N_43426,N_36939,N_31082);
nand U43427 (N_43427,N_36106,N_31653);
nor U43428 (N_43428,N_33122,N_39753);
nand U43429 (N_43429,N_32292,N_30502);
nand U43430 (N_43430,N_35369,N_31154);
nand U43431 (N_43431,N_32826,N_32450);
nor U43432 (N_43432,N_37276,N_36167);
or U43433 (N_43433,N_39953,N_36321);
xnor U43434 (N_43434,N_31450,N_36779);
xor U43435 (N_43435,N_31865,N_36786);
nand U43436 (N_43436,N_37620,N_36623);
nor U43437 (N_43437,N_30201,N_39966);
and U43438 (N_43438,N_31364,N_32838);
or U43439 (N_43439,N_37428,N_35121);
nor U43440 (N_43440,N_30030,N_37495);
or U43441 (N_43441,N_33394,N_30970);
xor U43442 (N_43442,N_33310,N_33096);
xor U43443 (N_43443,N_33987,N_31080);
nor U43444 (N_43444,N_37950,N_36901);
or U43445 (N_43445,N_36229,N_34329);
or U43446 (N_43446,N_39492,N_37121);
nand U43447 (N_43447,N_39114,N_34224);
nor U43448 (N_43448,N_33811,N_30638);
nand U43449 (N_43449,N_35580,N_37744);
nand U43450 (N_43450,N_30608,N_35791);
and U43451 (N_43451,N_33755,N_32193);
xor U43452 (N_43452,N_30376,N_32085);
nor U43453 (N_43453,N_36501,N_35100);
or U43454 (N_43454,N_38320,N_34571);
or U43455 (N_43455,N_33861,N_31894);
or U43456 (N_43456,N_36374,N_36312);
nand U43457 (N_43457,N_30192,N_35688);
xor U43458 (N_43458,N_30354,N_38529);
nor U43459 (N_43459,N_33233,N_35823);
xnor U43460 (N_43460,N_36817,N_31672);
xnor U43461 (N_43461,N_32120,N_36323);
and U43462 (N_43462,N_30279,N_34832);
and U43463 (N_43463,N_31298,N_34730);
nor U43464 (N_43464,N_31783,N_36247);
or U43465 (N_43465,N_36733,N_34627);
and U43466 (N_43466,N_34485,N_33576);
nand U43467 (N_43467,N_32746,N_35733);
nand U43468 (N_43468,N_38416,N_36073);
nand U43469 (N_43469,N_32981,N_38469);
nand U43470 (N_43470,N_34628,N_31018);
or U43471 (N_43471,N_39401,N_39345);
nor U43472 (N_43472,N_33749,N_35625);
xor U43473 (N_43473,N_32903,N_30326);
xor U43474 (N_43474,N_31516,N_36493);
nor U43475 (N_43475,N_31752,N_38049);
nor U43476 (N_43476,N_34820,N_37348);
nor U43477 (N_43477,N_37798,N_32247);
and U43478 (N_43478,N_35007,N_39570);
xor U43479 (N_43479,N_33397,N_31851);
nor U43480 (N_43480,N_31307,N_31303);
xor U43481 (N_43481,N_32264,N_34346);
nor U43482 (N_43482,N_35601,N_35001);
nand U43483 (N_43483,N_31455,N_35707);
and U43484 (N_43484,N_33833,N_33220);
or U43485 (N_43485,N_30787,N_33389);
nand U43486 (N_43486,N_39929,N_30736);
and U43487 (N_43487,N_36711,N_39648);
or U43488 (N_43488,N_38394,N_33262);
nand U43489 (N_43489,N_37883,N_30277);
nand U43490 (N_43490,N_31569,N_33111);
and U43491 (N_43491,N_39999,N_38550);
and U43492 (N_43492,N_33558,N_30093);
xor U43493 (N_43493,N_35660,N_30245);
and U43494 (N_43494,N_32718,N_32936);
and U43495 (N_43495,N_35341,N_39680);
nor U43496 (N_43496,N_34871,N_33472);
and U43497 (N_43497,N_37708,N_31614);
nand U43498 (N_43498,N_31594,N_30002);
and U43499 (N_43499,N_34635,N_31707);
nor U43500 (N_43500,N_31314,N_38800);
and U43501 (N_43501,N_37881,N_31266);
nand U43502 (N_43502,N_35049,N_38085);
or U43503 (N_43503,N_31885,N_37099);
nor U43504 (N_43504,N_34422,N_38844);
and U43505 (N_43505,N_31421,N_31028);
nand U43506 (N_43506,N_34462,N_35347);
or U43507 (N_43507,N_31659,N_34801);
and U43508 (N_43508,N_36860,N_31890);
xnor U43509 (N_43509,N_35184,N_37104);
nor U43510 (N_43510,N_33033,N_33464);
nand U43511 (N_43511,N_33812,N_33133);
xor U43512 (N_43512,N_30918,N_38818);
and U43513 (N_43513,N_34420,N_31780);
nor U43514 (N_43514,N_39846,N_39824);
nand U43515 (N_43515,N_34890,N_36459);
nor U43516 (N_43516,N_36705,N_39609);
nor U43517 (N_43517,N_30572,N_37630);
and U43518 (N_43518,N_39108,N_34577);
and U43519 (N_43519,N_36973,N_32447);
nor U43520 (N_43520,N_37078,N_39125);
or U43521 (N_43521,N_37453,N_36128);
nand U43522 (N_43522,N_34019,N_35549);
xnor U43523 (N_43523,N_36920,N_33086);
and U43524 (N_43524,N_36237,N_33866);
xnor U43525 (N_43525,N_35302,N_32591);
nand U43526 (N_43526,N_35193,N_35596);
nor U43527 (N_43527,N_34872,N_32921);
and U43528 (N_43528,N_37467,N_35362);
nand U43529 (N_43529,N_33911,N_34242);
xor U43530 (N_43530,N_38100,N_33004);
xnor U43531 (N_43531,N_32545,N_37471);
nand U43532 (N_43532,N_37791,N_33549);
and U43533 (N_43533,N_34701,N_38921);
nor U43534 (N_43534,N_33695,N_30809);
or U43535 (N_43535,N_30577,N_31666);
or U43536 (N_43536,N_39249,N_38713);
and U43537 (N_43537,N_38591,N_30711);
or U43538 (N_43538,N_37706,N_31180);
xnor U43539 (N_43539,N_32002,N_31462);
xor U43540 (N_43540,N_34645,N_39806);
or U43541 (N_43541,N_36559,N_39239);
and U43542 (N_43542,N_35944,N_37926);
nor U43543 (N_43543,N_30830,N_36124);
nor U43544 (N_43544,N_36269,N_37482);
or U43545 (N_43545,N_33253,N_30064);
nand U43546 (N_43546,N_32862,N_37233);
nand U43547 (N_43547,N_31844,N_32618);
nor U43548 (N_43548,N_32554,N_33332);
nand U43549 (N_43549,N_32590,N_36109);
nand U43550 (N_43550,N_32177,N_37191);
or U43551 (N_43551,N_37921,N_31753);
or U43552 (N_43552,N_30719,N_33646);
nor U43553 (N_43553,N_30721,N_36693);
nand U43554 (N_43554,N_30993,N_30004);
xor U43555 (N_43555,N_37957,N_30481);
xnor U43556 (N_43556,N_30811,N_38342);
or U43557 (N_43557,N_36344,N_39677);
and U43558 (N_43558,N_30565,N_39666);
nor U43559 (N_43559,N_38044,N_33668);
nand U43560 (N_43560,N_36330,N_30051);
or U43561 (N_43561,N_32613,N_35703);
xor U43562 (N_43562,N_35941,N_34022);
or U43563 (N_43563,N_38291,N_39757);
and U43564 (N_43564,N_34497,N_32492);
or U43565 (N_43565,N_36638,N_38926);
and U43566 (N_43566,N_37824,N_35665);
xor U43567 (N_43567,N_32854,N_34036);
nor U43568 (N_43568,N_37573,N_38731);
nor U43569 (N_43569,N_32440,N_32628);
nor U43570 (N_43570,N_34533,N_30313);
nand U43571 (N_43571,N_32233,N_35995);
nor U43572 (N_43572,N_32849,N_36287);
and U43573 (N_43573,N_35342,N_38503);
and U43574 (N_43574,N_34908,N_32748);
nand U43575 (N_43575,N_34946,N_38192);
nand U43576 (N_43576,N_38293,N_33125);
or U43577 (N_43577,N_30140,N_31467);
nand U43578 (N_43578,N_39110,N_34072);
nand U43579 (N_43579,N_32298,N_34259);
and U43580 (N_43580,N_39911,N_39024);
and U43581 (N_43581,N_37170,N_31586);
nor U43582 (N_43582,N_36361,N_35133);
nor U43583 (N_43583,N_36239,N_32738);
or U43584 (N_43584,N_33399,N_31896);
and U43585 (N_43585,N_38261,N_38267);
and U43586 (N_43586,N_38617,N_39015);
nand U43587 (N_43587,N_38001,N_30121);
xnor U43588 (N_43588,N_33828,N_35597);
nand U43589 (N_43589,N_32050,N_32818);
nor U43590 (N_43590,N_32867,N_38464);
or U43591 (N_43591,N_33260,N_31362);
xnor U43592 (N_43592,N_38555,N_31856);
and U43593 (N_43593,N_34252,N_31934);
nand U43594 (N_43594,N_32769,N_38757);
xor U43595 (N_43595,N_37691,N_36490);
nor U43596 (N_43596,N_37427,N_34574);
nand U43597 (N_43597,N_31668,N_30666);
and U43598 (N_43598,N_32873,N_31302);
nand U43599 (N_43599,N_38763,N_36796);
and U43600 (N_43600,N_39376,N_36500);
or U43601 (N_43601,N_39464,N_38474);
and U43602 (N_43602,N_33412,N_38000);
and U43603 (N_43603,N_37709,N_32992);
and U43604 (N_43604,N_30509,N_33871);
or U43605 (N_43605,N_39323,N_32880);
xnor U43606 (N_43606,N_32415,N_39790);
nor U43607 (N_43607,N_30965,N_31261);
nor U43608 (N_43608,N_32972,N_39713);
nor U43609 (N_43609,N_39815,N_37346);
nand U43610 (N_43610,N_32549,N_31910);
xor U43611 (N_43611,N_38084,N_37110);
nor U43612 (N_43612,N_31024,N_39925);
or U43613 (N_43613,N_34397,N_39531);
and U43614 (N_43614,N_38619,N_35241);
nand U43615 (N_43615,N_38128,N_39591);
xnor U43616 (N_43616,N_34032,N_36862);
nand U43617 (N_43617,N_35676,N_30887);
xor U43618 (N_43618,N_34864,N_39011);
xnor U43619 (N_43619,N_34611,N_39602);
or U43620 (N_43620,N_34468,N_33762);
and U43621 (N_43621,N_35215,N_35606);
and U43622 (N_43622,N_31135,N_39840);
nand U43623 (N_43623,N_30562,N_39041);
nand U43624 (N_43624,N_37944,N_31736);
xnor U43625 (N_43625,N_31606,N_32609);
and U43626 (N_43626,N_36844,N_33489);
xor U43627 (N_43627,N_31220,N_35099);
xor U43628 (N_43628,N_35805,N_37560);
nor U43629 (N_43629,N_35970,N_38468);
xnor U43630 (N_43630,N_30616,N_33703);
xor U43631 (N_43631,N_38165,N_38180);
nor U43632 (N_43632,N_30551,N_36742);
or U43633 (N_43633,N_37516,N_32540);
nor U43634 (N_43634,N_30728,N_34698);
xnor U43635 (N_43635,N_38771,N_36768);
nand U43636 (N_43636,N_35056,N_34556);
nand U43637 (N_43637,N_38684,N_34434);
and U43638 (N_43638,N_33778,N_36010);
xnor U43639 (N_43639,N_36021,N_38288);
and U43640 (N_43640,N_33230,N_31536);
nor U43641 (N_43641,N_38944,N_37116);
and U43642 (N_43642,N_31197,N_34012);
xor U43643 (N_43643,N_31042,N_31099);
nor U43644 (N_43644,N_33141,N_34947);
or U43645 (N_43645,N_37190,N_38063);
and U43646 (N_43646,N_36716,N_36257);
and U43647 (N_43647,N_34014,N_35394);
nor U43648 (N_43648,N_35593,N_30361);
and U43649 (N_43649,N_37682,N_38794);
nand U43650 (N_43650,N_30594,N_37200);
xor U43651 (N_43651,N_31323,N_33849);
and U43652 (N_43652,N_32890,N_33006);
nand U43653 (N_43653,N_36637,N_35756);
or U43654 (N_43654,N_35111,N_30489);
and U43655 (N_43655,N_36403,N_33516);
nor U43656 (N_43656,N_35905,N_33393);
or U43657 (N_43657,N_38052,N_35185);
nand U43658 (N_43658,N_38964,N_37129);
nor U43659 (N_43659,N_33309,N_38068);
or U43660 (N_43660,N_30620,N_35294);
and U43661 (N_43661,N_33374,N_35271);
nand U43662 (N_43662,N_32569,N_32169);
xor U43663 (N_43663,N_37356,N_38741);
or U43664 (N_43664,N_33878,N_38242);
nor U43665 (N_43665,N_30700,N_36674);
xnor U43666 (N_43666,N_30575,N_34831);
nand U43667 (N_43667,N_34965,N_37720);
or U43668 (N_43668,N_39169,N_31576);
nor U43669 (N_43669,N_35466,N_30969);
xnor U43670 (N_43670,N_33770,N_35710);
xnor U43671 (N_43671,N_38883,N_31725);
and U43672 (N_43672,N_36664,N_31995);
nand U43673 (N_43673,N_38035,N_30573);
nor U43674 (N_43674,N_35611,N_36409);
nand U43675 (N_43675,N_33957,N_35931);
and U43676 (N_43676,N_32093,N_39574);
and U43677 (N_43677,N_36055,N_35487);
xnor U43678 (N_43678,N_32666,N_35907);
and U43679 (N_43679,N_37943,N_38957);
and U43680 (N_43680,N_33537,N_38540);
nand U43681 (N_43681,N_36923,N_32341);
or U43682 (N_43682,N_37007,N_35125);
or U43683 (N_43683,N_39291,N_34920);
nor U43684 (N_43684,N_35081,N_35815);
nor U43685 (N_43685,N_36274,N_33547);
or U43686 (N_43686,N_35717,N_38996);
or U43687 (N_43687,N_37472,N_34983);
nand U43688 (N_43688,N_31281,N_31290);
and U43689 (N_43689,N_39821,N_31522);
or U43690 (N_43690,N_34772,N_38607);
nor U43691 (N_43691,N_33704,N_39708);
nand U43692 (N_43692,N_37270,N_34423);
or U43693 (N_43693,N_35417,N_32819);
and U43694 (N_43694,N_32840,N_34700);
or U43695 (N_43695,N_38983,N_36060);
and U43696 (N_43696,N_30840,N_36503);
xnor U43697 (N_43697,N_39280,N_39719);
or U43698 (N_43698,N_32296,N_34987);
nor U43699 (N_43699,N_34400,N_39242);
or U43700 (N_43700,N_39994,N_30007);
xnor U43701 (N_43701,N_33194,N_35024);
nand U43702 (N_43702,N_35040,N_31332);
xor U43703 (N_43703,N_35752,N_31031);
nor U43704 (N_43704,N_31473,N_32059);
nand U43705 (N_43705,N_30976,N_32096);
nand U43706 (N_43706,N_30147,N_36993);
nand U43707 (N_43707,N_30847,N_34907);
nor U43708 (N_43708,N_39623,N_36971);
nand U43709 (N_43709,N_31073,N_30042);
and U43710 (N_43710,N_37470,N_36743);
xor U43711 (N_43711,N_38613,N_39186);
nor U43712 (N_43712,N_30888,N_36065);
or U43713 (N_43713,N_38909,N_39359);
xor U43714 (N_43714,N_31573,N_38487);
nor U43715 (N_43715,N_33283,N_39181);
xor U43716 (N_43716,N_36648,N_36520);
nor U43717 (N_43717,N_37208,N_33746);
nand U43718 (N_43718,N_32699,N_35426);
nor U43719 (N_43719,N_38072,N_37887);
xor U43720 (N_43720,N_34512,N_33934);
nand U43721 (N_43721,N_39021,N_32767);
xor U43722 (N_43722,N_30564,N_34377);
nor U43723 (N_43723,N_35939,N_30798);
nand U43724 (N_43724,N_38645,N_30129);
xnor U43725 (N_43725,N_36190,N_39897);
and U43726 (N_43726,N_34703,N_35192);
xor U43727 (N_43727,N_33185,N_31952);
nand U43728 (N_43728,N_31501,N_36524);
and U43729 (N_43729,N_39363,N_33892);
and U43730 (N_43730,N_38222,N_37948);
nand U43731 (N_43731,N_34775,N_32309);
nand U43732 (N_43732,N_36717,N_31670);
nand U43733 (N_43733,N_38685,N_30165);
and U43734 (N_43734,N_30096,N_30441);
xnor U43735 (N_43735,N_39039,N_30781);
nor U43736 (N_43736,N_30915,N_37269);
nor U43737 (N_43737,N_31172,N_32520);
or U43738 (N_43738,N_39776,N_34287);
nor U43739 (N_43739,N_38240,N_31232);
or U43740 (N_43740,N_33213,N_38456);
nor U43741 (N_43741,N_30204,N_37739);
nor U43742 (N_43742,N_35104,N_32625);
nor U43743 (N_43743,N_30356,N_38985);
and U43744 (N_43744,N_38498,N_34331);
and U43745 (N_43745,N_33020,N_33500);
and U43746 (N_43746,N_37559,N_35094);
or U43747 (N_43747,N_30417,N_36272);
nor U43748 (N_43748,N_39535,N_34143);
or U43749 (N_43749,N_35265,N_33722);
nor U43750 (N_43750,N_39834,N_38700);
and U43751 (N_43751,N_33087,N_33886);
nor U43752 (N_43752,N_37783,N_32437);
xor U43753 (N_43753,N_32280,N_33377);
or U43754 (N_43754,N_36049,N_34079);
and U43755 (N_43755,N_33387,N_33444);
nor U43756 (N_43756,N_32023,N_30820);
nand U43757 (N_43757,N_36589,N_36431);
nand U43758 (N_43758,N_38479,N_38524);
and U43759 (N_43759,N_38069,N_38646);
nand U43760 (N_43760,N_39208,N_39485);
or U43761 (N_43761,N_33883,N_30271);
xnor U43762 (N_43762,N_33151,N_39814);
and U43763 (N_43763,N_31873,N_36588);
xor U43764 (N_43764,N_32427,N_32332);
nand U43765 (N_43765,N_30695,N_36434);
nor U43766 (N_43766,N_38096,N_32018);
nand U43767 (N_43767,N_33827,N_39616);
or U43768 (N_43768,N_37736,N_30521);
xnor U43769 (N_43769,N_33600,N_32477);
and U43770 (N_43770,N_39405,N_30449);
nand U43771 (N_43771,N_33562,N_37232);
nand U43772 (N_43772,N_38378,N_30741);
nor U43773 (N_43773,N_37469,N_38093);
and U43774 (N_43774,N_32714,N_36123);
and U43775 (N_43775,N_30869,N_37754);
nand U43776 (N_43776,N_37800,N_32787);
nand U43777 (N_43777,N_39644,N_38318);
nor U43778 (N_43778,N_38301,N_33731);
xor U43779 (N_43779,N_35397,N_30845);
nor U43780 (N_43780,N_39275,N_35493);
nor U43781 (N_43781,N_33648,N_35772);
nand U43782 (N_43782,N_38546,N_30981);
and U43783 (N_43783,N_30800,N_33191);
nand U43784 (N_43784,N_36985,N_38067);
nand U43785 (N_43785,N_38151,N_37494);
or U43786 (N_43786,N_30391,N_39328);
or U43787 (N_43787,N_32857,N_35161);
nor U43788 (N_43788,N_36534,N_35643);
nor U43789 (N_43789,N_35903,N_33408);
nand U43790 (N_43790,N_32512,N_34563);
nor U43791 (N_43791,N_30256,N_39619);
or U43792 (N_43792,N_36833,N_35862);
and U43793 (N_43793,N_35086,N_34588);
or U43794 (N_43794,N_30866,N_36093);
nor U43795 (N_43795,N_37032,N_39423);
xnor U43796 (N_43796,N_33913,N_37480);
and U43797 (N_43797,N_36166,N_35494);
xor U43798 (N_43798,N_30148,N_38872);
and U43799 (N_43799,N_34759,N_35919);
and U43800 (N_43800,N_39461,N_34042);
nand U43801 (N_43801,N_30533,N_36118);
nor U43802 (N_43802,N_37323,N_36070);
or U43803 (N_43803,N_32742,N_38030);
xor U43804 (N_43804,N_32489,N_37329);
nand U43805 (N_43805,N_34304,N_33048);
or U43806 (N_43806,N_33627,N_30657);
or U43807 (N_43807,N_36121,N_31111);
xnor U43808 (N_43808,N_37352,N_37037);
xor U43809 (N_43809,N_37696,N_31883);
xnor U43810 (N_43810,N_37264,N_34352);
xnor U43811 (N_43811,N_31615,N_32791);
nor U43812 (N_43812,N_38751,N_38586);
nand U43813 (N_43813,N_33567,N_37261);
or U43814 (N_43814,N_39652,N_31092);
nand U43815 (N_43815,N_32775,N_35993);
xor U43816 (N_43816,N_34691,N_34937);
nand U43817 (N_43817,N_30501,N_39285);
or U43818 (N_43818,N_39871,N_36544);
xor U43819 (N_43819,N_39534,N_31966);
and U43820 (N_43820,N_38369,N_35419);
nand U43821 (N_43821,N_35279,N_39219);
xor U43822 (N_43822,N_33601,N_35766);
nor U43823 (N_43823,N_32070,N_36806);
nor U43824 (N_43824,N_37322,N_39235);
or U43825 (N_43825,N_37518,N_32377);
nand U43826 (N_43826,N_37806,N_34631);
nand U43827 (N_43827,N_36083,N_36235);
xor U43828 (N_43828,N_33777,N_32182);
and U43829 (N_43829,N_37959,N_31326);
and U43830 (N_43830,N_37285,N_33279);
xor U43831 (N_43831,N_33221,N_33268);
or U43832 (N_43832,N_30997,N_31918);
nand U43833 (N_43833,N_35658,N_38231);
nand U43834 (N_43834,N_31438,N_32073);
xor U43835 (N_43835,N_36030,N_35364);
or U43836 (N_43836,N_38370,N_39228);
and U43837 (N_43837,N_39416,N_36126);
xor U43838 (N_43838,N_35053,N_35401);
nand U43839 (N_43839,N_31238,N_38719);
nand U43840 (N_43840,N_35250,N_30813);
nor U43841 (N_43841,N_39199,N_34325);
and U43842 (N_43842,N_39733,N_33832);
xnor U43843 (N_43843,N_39803,N_35239);
or U43844 (N_43844,N_39509,N_30351);
nand U43845 (N_43845,N_35036,N_38606);
xnor U43846 (N_43846,N_30154,N_36616);
xor U43847 (N_43847,N_33161,N_39860);
nand U43848 (N_43848,N_32639,N_30142);
xor U43849 (N_43849,N_32453,N_31669);
nand U43850 (N_43850,N_35061,N_31679);
xor U43851 (N_43851,N_35560,N_33808);
xnor U43852 (N_43852,N_30372,N_33217);
nor U43853 (N_43853,N_34815,N_33686);
xor U43854 (N_43854,N_32132,N_30731);
and U43855 (N_43855,N_33768,N_37430);
and U43856 (N_43856,N_30221,N_30590);
or U43857 (N_43857,N_37004,N_37591);
and U43858 (N_43858,N_35683,N_36097);
nand U43859 (N_43859,N_39232,N_34124);
and U43860 (N_43860,N_32297,N_39516);
nor U43861 (N_43861,N_30958,N_36573);
or U43862 (N_43862,N_30609,N_32865);
and U43863 (N_43863,N_33735,N_37971);
or U43864 (N_43864,N_33188,N_38548);
nand U43865 (N_43865,N_34558,N_38804);
xnor U43866 (N_43866,N_31160,N_30367);
nand U43867 (N_43867,N_36990,N_37040);
or U43868 (N_43868,N_35517,N_37612);
or U43869 (N_43869,N_38747,N_33254);
nor U43870 (N_43870,N_36700,N_35761);
nor U43871 (N_43871,N_31157,N_37812);
and U43872 (N_43872,N_33506,N_36526);
and U43873 (N_43873,N_37822,N_30511);
nor U43874 (N_43874,N_30348,N_36538);
and U43875 (N_43875,N_35514,N_31640);
nand U43876 (N_43876,N_38544,N_36372);
nand U43877 (N_43877,N_39179,N_35360);
xor U43878 (N_43878,N_34133,N_32708);
nor U43879 (N_43879,N_33080,N_33118);
or U43880 (N_43880,N_36529,N_38145);
xor U43881 (N_43881,N_35256,N_38724);
nor U43882 (N_43882,N_32373,N_30797);
xor U43883 (N_43883,N_38140,N_38519);
or U43884 (N_43884,N_38940,N_38162);
and U43885 (N_43885,N_33065,N_32495);
nor U43886 (N_43886,N_35893,N_30643);
xor U43887 (N_43887,N_37282,N_34317);
nor U43888 (N_43888,N_31104,N_34841);
nor U43889 (N_43889,N_38341,N_32837);
or U43890 (N_43890,N_30995,N_33613);
xnor U43891 (N_43891,N_39209,N_36103);
and U43892 (N_43892,N_31967,N_31540);
or U43893 (N_43893,N_39127,N_35216);
xnor U43894 (N_43894,N_30625,N_37151);
nand U43895 (N_43895,N_38452,N_31992);
nor U43896 (N_43896,N_35897,N_38711);
nor U43897 (N_43897,N_35156,N_31453);
or U43898 (N_43898,N_39552,N_30346);
nand U43899 (N_43899,N_33400,N_33138);
or U43900 (N_43900,N_39965,N_32394);
and U43901 (N_43901,N_30624,N_30371);
nor U43902 (N_43902,N_30904,N_35485);
nor U43903 (N_43903,N_31635,N_34142);
or U43904 (N_43904,N_38893,N_32250);
xor U43905 (N_43905,N_35131,N_34861);
nor U43906 (N_43906,N_36482,N_32874);
or U43907 (N_43907,N_34435,N_36525);
or U43908 (N_43908,N_35787,N_38155);
and U43909 (N_43909,N_35135,N_39217);
xor U43910 (N_43910,N_34740,N_32993);
nor U43911 (N_43911,N_38970,N_33854);
and U43912 (N_43912,N_36780,N_33093);
nor U43913 (N_43913,N_33906,N_35626);
and U43914 (N_43914,N_30679,N_34426);
or U43915 (N_43915,N_33688,N_38779);
nand U43916 (N_43916,N_39025,N_31021);
or U43917 (N_43917,N_30079,N_38274);
xor U43918 (N_43918,N_35851,N_33365);
and U43919 (N_43919,N_30119,N_33862);
and U43920 (N_43920,N_39194,N_36044);
xor U43921 (N_43921,N_33708,N_31600);
or U43922 (N_43922,N_37283,N_32940);
or U43923 (N_43923,N_31373,N_32695);
nand U43924 (N_43924,N_34447,N_32187);
nor U43925 (N_43925,N_37786,N_31176);
nor U43926 (N_43926,N_37864,N_34622);
and U43927 (N_43927,N_38549,N_38718);
or U43928 (N_43928,N_37324,N_35794);
and U43929 (N_43929,N_35128,N_38082);
or U43930 (N_43930,N_32717,N_36603);
or U43931 (N_43931,N_37631,N_37117);
or U43932 (N_43932,N_39559,N_32664);
or U43933 (N_43933,N_31437,N_36950);
nor U43934 (N_43934,N_38483,N_35503);
nand U43935 (N_43935,N_38688,N_37230);
nand U43936 (N_43936,N_34045,N_32165);
nor U43937 (N_43937,N_33132,N_30876);
and U43938 (N_43938,N_36994,N_37666);
xnor U43939 (N_43939,N_36045,N_32230);
and U43940 (N_43940,N_37734,N_39976);
or U43941 (N_43941,N_33579,N_34702);
or U43942 (N_43942,N_38227,N_32726);
nand U43943 (N_43943,N_30557,N_35475);
and U43944 (N_43944,N_30518,N_38631);
and U43945 (N_43945,N_30861,N_30102);
and U43946 (N_43946,N_33317,N_37588);
and U43947 (N_43947,N_38600,N_31542);
xnor U43948 (N_43948,N_38283,N_35231);
nor U43949 (N_43949,N_30265,N_36453);
nand U43950 (N_43950,N_34769,N_34370);
and U43951 (N_43951,N_31727,N_38670);
nand U43952 (N_43952,N_35143,N_37475);
nand U43953 (N_43953,N_34394,N_39717);
and U43954 (N_43954,N_32354,N_34757);
and U43955 (N_43955,N_30927,N_37897);
nor U43956 (N_43956,N_35630,N_33277);
nand U43957 (N_43957,N_30216,N_37492);
and U43958 (N_43958,N_36217,N_38083);
xor U43959 (N_43959,N_39365,N_39679);
nor U43960 (N_43960,N_38120,N_30133);
xor U43961 (N_43961,N_30722,N_39595);
nor U43962 (N_43962,N_32616,N_37544);
nand U43963 (N_43963,N_34979,N_37155);
nor U43964 (N_43964,N_39610,N_33017);
xor U43965 (N_43965,N_35636,N_37814);
nand U43966 (N_43966,N_33159,N_34057);
and U43967 (N_43967,N_38366,N_39267);
nor U43968 (N_43968,N_34284,N_39355);
nor U43969 (N_43969,N_35436,N_38493);
and U43970 (N_43970,N_35575,N_34100);
nor U43971 (N_43971,N_38564,N_37361);
and U43972 (N_43972,N_33027,N_39297);
or U43973 (N_43973,N_34929,N_32793);
xor U43974 (N_43974,N_32505,N_30053);
nor U43975 (N_43975,N_37927,N_38563);
or U43976 (N_43976,N_33486,N_30288);
nand U43977 (N_43977,N_36216,N_34044);
and U43978 (N_43978,N_36111,N_33794);
nand U43979 (N_43979,N_38177,N_38256);
and U43980 (N_43980,N_32414,N_33650);
and U43981 (N_43981,N_38400,N_33099);
nand U43982 (N_43982,N_38377,N_34958);
or U43983 (N_43983,N_31634,N_31417);
nand U43984 (N_43984,N_37606,N_38024);
nand U43985 (N_43985,N_35379,N_37759);
nand U43986 (N_43986,N_39923,N_31713);
nor U43987 (N_43987,N_35522,N_39870);
nand U43988 (N_43988,N_39572,N_34927);
nand U43989 (N_43989,N_30170,N_38887);
nand U43990 (N_43990,N_36318,N_33144);
nand U43991 (N_43991,N_39918,N_32712);
xnor U43992 (N_43992,N_35587,N_37039);
nand U43993 (N_43993,N_39187,N_39432);
nand U43994 (N_43994,N_38048,N_32833);
xnor U43995 (N_43995,N_38110,N_37571);
and U43996 (N_43996,N_32820,N_33858);
and U43997 (N_43997,N_31468,N_33539);
xor U43998 (N_43998,N_33273,N_30653);
and U43999 (N_43999,N_32151,N_36835);
nand U44000 (N_44000,N_38742,N_37901);
xnor U44001 (N_44001,N_32404,N_33699);
nand U44002 (N_44002,N_35827,N_33066);
or U44003 (N_44003,N_38186,N_39454);
and U44004 (N_44004,N_37413,N_31957);
xor U44005 (N_44005,N_38648,N_30739);
nor U44006 (N_44006,N_39057,N_39795);
nand U44007 (N_44007,N_34836,N_30479);
xor U44008 (N_44008,N_39608,N_36334);
and U44009 (N_44009,N_33266,N_38557);
xor U44010 (N_44010,N_34619,N_39731);
and U44011 (N_44011,N_32844,N_39720);
nor U44012 (N_44012,N_36062,N_30808);
nor U44013 (N_44013,N_30137,N_33012);
xnor U44014 (N_44014,N_38281,N_30203);
or U44015 (N_44015,N_36567,N_32601);
nor U44016 (N_44016,N_33120,N_35961);
nand U44017 (N_44017,N_39936,N_32237);
xnor U44018 (N_44018,N_36636,N_31083);
or U44019 (N_44019,N_36680,N_30574);
nand U44020 (N_44020,N_37601,N_31447);
or U44021 (N_44021,N_38988,N_32142);
or U44022 (N_44022,N_30083,N_37956);
nand U44023 (N_44023,N_30461,N_34276);
or U44024 (N_44024,N_33665,N_38245);
xnor U44025 (N_44025,N_39196,N_30359);
nand U44026 (N_44026,N_36378,N_30035);
or U44027 (N_44027,N_32636,N_35488);
nand U44028 (N_44028,N_31744,N_30176);
and U44029 (N_44029,N_38453,N_35689);
and U44030 (N_44030,N_30920,N_32335);
and U44031 (N_44031,N_38834,N_30433);
xor U44032 (N_44032,N_32953,N_39251);
nand U44033 (N_44033,N_37583,N_37400);
and U44034 (N_44034,N_35119,N_35895);
or U44035 (N_44035,N_35415,N_30990);
nor U44036 (N_44036,N_33371,N_36646);
and U44037 (N_44037,N_37359,N_32443);
and U44038 (N_44038,N_31578,N_30273);
xor U44039 (N_44039,N_39791,N_39255);
and U44040 (N_44040,N_33566,N_34443);
nor U44041 (N_44041,N_31909,N_36596);
xnor U44042 (N_44042,N_35896,N_31950);
xnor U44043 (N_44043,N_32788,N_34218);
xor U44044 (N_44044,N_38933,N_34760);
or U44045 (N_44045,N_30269,N_33109);
nand U44046 (N_44046,N_37855,N_39861);
nor U44047 (N_44047,N_34314,N_32845);
nand U44048 (N_44048,N_36645,N_36096);
xor U44049 (N_44049,N_32750,N_36948);
or U44050 (N_44050,N_36492,N_35875);
or U44051 (N_44051,N_30305,N_30032);
nand U44052 (N_44052,N_38775,N_39435);
or U44053 (N_44053,N_34065,N_32731);
nand U44054 (N_44054,N_37644,N_34061);
nor U44055 (N_44055,N_39207,N_33983);
and U44056 (N_44056,N_36144,N_31493);
xnor U44057 (N_44057,N_31354,N_36988);
nand U44058 (N_44058,N_39370,N_38710);
xnor U44059 (N_44059,N_30202,N_34779);
or U44060 (N_44060,N_30702,N_35422);
nand U44061 (N_44061,N_33498,N_35654);
and U44062 (N_44062,N_31774,N_33551);
xor U44063 (N_44063,N_34318,N_38232);
nand U44064 (N_44064,N_36516,N_37528);
or U44065 (N_44065,N_38681,N_35000);
xor U44066 (N_44066,N_38497,N_38238);
or U44067 (N_44067,N_36749,N_33868);
and U44068 (N_44068,N_37843,N_33606);
nand U44069 (N_44069,N_30770,N_38408);
and U44070 (N_44070,N_30865,N_32283);
nand U44071 (N_44071,N_34521,N_37690);
or U44072 (N_44072,N_30803,N_33938);
and U44073 (N_44073,N_39170,N_30290);
nor U44074 (N_44074,N_31709,N_36821);
or U44075 (N_44075,N_35062,N_34470);
nand U44076 (N_44076,N_33507,N_39197);
nand U44077 (N_44077,N_37951,N_30640);
nand U44078 (N_44078,N_31847,N_33165);
xnor U44079 (N_44079,N_30012,N_37333);
or U44080 (N_44080,N_36442,N_30187);
or U44081 (N_44081,N_30443,N_34358);
or U44082 (N_44082,N_38249,N_34623);
nor U44083 (N_44083,N_35713,N_37477);
and U44084 (N_44084,N_38895,N_37279);
and U44085 (N_44085,N_34724,N_35933);
nand U44086 (N_44086,N_32390,N_32574);
nor U44087 (N_44087,N_37870,N_39204);
nor U44088 (N_44088,N_31954,N_31604);
and U44089 (N_44089,N_37723,N_33564);
nand U44090 (N_44090,N_34996,N_31376);
xnor U44091 (N_44091,N_30086,N_35972);
and U44092 (N_44092,N_34215,N_31382);
nor U44093 (N_44093,N_35405,N_31409);
nand U44094 (N_44094,N_39246,N_39044);
nand U44095 (N_44095,N_32950,N_36640);
and U44096 (N_44096,N_30194,N_30859);
xnor U44097 (N_44097,N_31764,N_36549);
and U44098 (N_44098,N_36643,N_37221);
nor U44099 (N_44099,N_33936,N_32519);
nor U44100 (N_44100,N_33710,N_32065);
and U44101 (N_44101,N_31776,N_31398);
and U44102 (N_44102,N_31652,N_34614);
nor U44103 (N_44103,N_32245,N_35908);
nand U44104 (N_44104,N_33919,N_30153);
and U44105 (N_44105,N_30907,N_37758);
and U44106 (N_44106,N_39593,N_30560);
or U44107 (N_44107,N_35214,N_35774);
xnor U44108 (N_44108,N_37813,N_38986);
nand U44109 (N_44109,N_35661,N_34977);
nand U44110 (N_44110,N_35857,N_37735);
nor U44111 (N_44111,N_39528,N_32930);
nand U44112 (N_44112,N_34684,N_30240);
xor U44113 (N_44113,N_34292,N_38490);
nor U44114 (N_44114,N_32363,N_35988);
xor U44115 (N_44115,N_39782,N_31548);
xnor U44116 (N_44116,N_37053,N_35550);
nor U44117 (N_44117,N_35595,N_31252);
or U44118 (N_44118,N_38127,N_37485);
nor U44119 (N_44119,N_37922,N_33997);
xnor U44120 (N_44120,N_36805,N_37947);
nand U44121 (N_44121,N_36896,N_30071);
xor U44122 (N_44122,N_30709,N_39565);
xnor U44123 (N_44123,N_31642,N_38492);
nor U44124 (N_44124,N_34734,N_31448);
xnor U44125 (N_44125,N_30111,N_33284);
nor U44126 (N_44126,N_34809,N_35365);
nand U44127 (N_44127,N_34679,N_32031);
and U44128 (N_44128,N_33918,N_38081);
xnor U44129 (N_44129,N_32987,N_35821);
and U44130 (N_44130,N_31922,N_37928);
xnor U44131 (N_44131,N_36581,N_36605);
nor U44132 (N_44132,N_38911,N_33818);
xnor U44133 (N_44133,N_39211,N_35600);
and U44134 (N_44134,N_38299,N_38533);
nand U44135 (N_44135,N_37575,N_37042);
nand U44136 (N_44136,N_34439,N_37858);
nor U44137 (N_44137,N_34077,N_30195);
nor U44138 (N_44138,N_35336,N_31700);
and U44139 (N_44139,N_33890,N_34530);
nor U44140 (N_44140,N_33203,N_34059);
nor U44141 (N_44141,N_35887,N_35390);
nand U44142 (N_44142,N_33955,N_33888);
nor U44143 (N_44143,N_34674,N_31719);
or U44144 (N_44144,N_32919,N_30939);
or U44145 (N_44145,N_39213,N_35900);
or U44146 (N_44146,N_30639,N_35705);
and U44147 (N_44147,N_30762,N_36527);
nand U44148 (N_44148,N_31633,N_39562);
xnor U44149 (N_44149,N_35492,N_34665);
xnor U44150 (N_44150,N_30316,N_31595);
and U44151 (N_44151,N_39278,N_35471);
nand U44152 (N_44152,N_31390,N_34870);
nor U44153 (N_44153,N_34835,N_39775);
xnor U44154 (N_44154,N_38856,N_32306);
nand U44155 (N_44155,N_37716,N_36104);
nand U44156 (N_44156,N_37911,N_35088);
xor U44157 (N_44157,N_30038,N_38042);
nand U44158 (N_44158,N_32631,N_36125);
nand U44159 (N_44159,N_39193,N_38207);
or U44160 (N_44160,N_33493,N_38028);
nor U44161 (N_44161,N_33496,N_36799);
or U44162 (N_44162,N_37976,N_34172);
xor U44163 (N_44163,N_32219,N_30767);
xnor U44164 (N_44164,N_32894,N_35880);
xnor U44165 (N_44165,N_35067,N_33661);
or U44166 (N_44166,N_35530,N_39941);
xor U44167 (N_44167,N_35103,N_34564);
nor U44168 (N_44168,N_37869,N_39443);
or U44169 (N_44169,N_37236,N_38569);
and U44170 (N_44170,N_39225,N_32420);
nand U44171 (N_44171,N_32957,N_36797);
nor U44172 (N_44172,N_31396,N_37183);
nand U44173 (N_44173,N_36281,N_36025);
nor U44174 (N_44174,N_37481,N_37863);
and U44175 (N_44175,N_39549,N_36077);
xnor U44176 (N_44176,N_31698,N_31118);
nor U44177 (N_44177,N_30831,N_32815);
nand U44178 (N_44178,N_30520,N_39414);
or U44179 (N_44179,N_37511,N_30329);
xnor U44180 (N_44180,N_34104,N_31415);
nand U44181 (N_44181,N_33596,N_31697);
xnor U44182 (N_44182,N_37486,N_31110);
and U44183 (N_44183,N_39300,N_39505);
nand U44184 (N_44184,N_36955,N_38159);
nor U44185 (N_44185,N_39468,N_37676);
and U44186 (N_44186,N_35954,N_32445);
or U44187 (N_44187,N_33667,N_37831);
and U44188 (N_44188,N_33216,N_34011);
and U44189 (N_44189,N_31748,N_37238);
or U44190 (N_44190,N_35174,N_35490);
xor U44191 (N_44191,N_30744,N_36794);
nand U44192 (N_44192,N_31223,N_38426);
nand U44193 (N_44193,N_34151,N_31862);
and U44194 (N_44194,N_36969,N_38596);
nand U44195 (N_44195,N_31859,N_32482);
xnor U44196 (N_44196,N_36162,N_35738);
and U44197 (N_44197,N_34932,N_31687);
xor U44198 (N_44198,N_33002,N_38720);
nand U44199 (N_44199,N_36986,N_32075);
nor U44200 (N_44200,N_30487,N_31940);
and U44201 (N_44201,N_38023,N_39890);
nor U44202 (N_44202,N_37574,N_39830);
and U44203 (N_44203,N_39320,N_35389);
and U44204 (N_44204,N_38236,N_31379);
xnor U44205 (N_44205,N_32126,N_35945);
or U44206 (N_44206,N_30661,N_39794);
nor U44207 (N_44207,N_33715,N_32853);
nand U44208 (N_44208,N_38163,N_30294);
nor U44209 (N_44209,N_36657,N_36771);
and U44210 (N_44210,N_39675,N_34683);
xnor U44211 (N_44211,N_34113,N_35421);
nand U44212 (N_44212,N_30896,N_30374);
xor U44213 (N_44213,N_31079,N_36319);
xor U44214 (N_44214,N_37988,N_37781);
or U44215 (N_44215,N_30445,N_36420);
or U44216 (N_44216,N_32262,N_33199);
or U44217 (N_44217,N_31100,N_32514);
nand U44218 (N_44218,N_30589,N_38612);
and U44219 (N_44219,N_35830,N_33885);
or U44220 (N_44220,N_33728,N_35468);
or U44221 (N_44221,N_30544,N_39174);
and U44222 (N_44222,N_39837,N_37094);
xnor U44223 (N_44223,N_32985,N_38347);
and U44224 (N_44224,N_32575,N_33702);
nor U44225 (N_44225,N_35145,N_36726);
or U44226 (N_44226,N_30155,N_31881);
or U44227 (N_44227,N_31545,N_31318);
nand U44228 (N_44228,N_37586,N_38478);
or U44229 (N_44229,N_34714,N_31377);
or U44230 (N_44230,N_36366,N_34153);
xnor U44231 (N_44231,N_32148,N_33383);
nand U44232 (N_44232,N_35715,N_37184);
nand U44233 (N_44233,N_39014,N_39668);
or U44234 (N_44234,N_35329,N_39759);
and U44235 (N_44235,N_35637,N_32797);
xnor U44236 (N_44236,N_39928,N_33628);
nor U44237 (N_44237,N_38597,N_31926);
or U44238 (N_44238,N_32118,N_37849);
or U44239 (N_44239,N_37126,N_36017);
xnor U44240 (N_44240,N_31166,N_39676);
nor U44241 (N_44241,N_35268,N_38618);
or U44242 (N_44242,N_33824,N_37918);
or U44243 (N_44243,N_35261,N_37205);
or U44244 (N_44244,N_38043,N_35110);
or U44245 (N_44245,N_36852,N_36908);
nand U44246 (N_44246,N_30816,N_37374);
nor U44247 (N_44247,N_34771,N_39698);
nor U44248 (N_44248,N_34584,N_31980);
xnor U44249 (N_44249,N_32480,N_38915);
or U44250 (N_44250,N_33877,N_38094);
nor U44251 (N_44251,N_36435,N_33602);
xnor U44252 (N_44252,N_32878,N_37199);
and U44253 (N_44253,N_35230,N_31564);
nor U44254 (N_44254,N_39451,N_36252);
or U44255 (N_44255,N_34825,N_39820);
or U44256 (N_44256,N_33117,N_38605);
or U44257 (N_44257,N_39550,N_36306);
xor U44258 (N_44258,N_34847,N_32920);
xnor U44259 (N_44259,N_35252,N_34028);
xnor U44260 (N_44260,N_34383,N_34948);
or U44261 (N_44261,N_33219,N_31924);
nor U44262 (N_44262,N_32039,N_33461);
and U44263 (N_44263,N_35339,N_33962);
or U44264 (N_44264,N_32057,N_33657);
xor U44265 (N_44265,N_30103,N_35776);
nand U44266 (N_44266,N_31227,N_39103);
or U44267 (N_44267,N_37862,N_39031);
and U44268 (N_44268,N_39109,N_34431);
and U44269 (N_44269,N_30011,N_33078);
and U44270 (N_44270,N_36696,N_32798);
nor U44271 (N_44271,N_32669,N_34403);
xor U44272 (N_44272,N_30304,N_37741);
and U44273 (N_44273,N_31923,N_33064);
and U44274 (N_44274,N_36195,N_37508);
nand U44275 (N_44275,N_30567,N_34853);
nand U44276 (N_44276,N_34391,N_30136);
xnor U44277 (N_44277,N_35870,N_37344);
and U44278 (N_44278,N_38424,N_34495);
and U44279 (N_44279,N_31470,N_31955);
and U44280 (N_44280,N_36807,N_30749);
nand U44281 (N_44281,N_32467,N_33615);
or U44282 (N_44282,N_31519,N_38980);
and U44283 (N_44283,N_39344,N_32918);
xor U44284 (N_44284,N_33553,N_32632);
xor U44285 (N_44285,N_38076,N_39094);
nor U44286 (N_44286,N_32139,N_39863);
xor U44287 (N_44287,N_30181,N_30784);
nand U44288 (N_44288,N_35182,N_34829);
and U44289 (N_44289,N_30549,N_33502);
and U44290 (N_44290,N_31821,N_35467);
nand U44291 (N_44291,N_33008,N_35132);
nand U44292 (N_44292,N_33337,N_32770);
and U44293 (N_44293,N_32640,N_36056);
and U44294 (N_44294,N_38927,N_39477);
nor U44295 (N_44295,N_32571,N_34127);
or U44296 (N_44296,N_32409,N_30300);
nand U44297 (N_44297,N_34017,N_34696);
or U44298 (N_44298,N_38987,N_35474);
and U44299 (N_44299,N_31850,N_30411);
and U44300 (N_44300,N_34353,N_39276);
and U44301 (N_44301,N_32900,N_32702);
nand U44302 (N_44302,N_30314,N_37437);
xor U44303 (N_44303,N_30506,N_33705);
nand U44304 (N_44304,N_32359,N_35378);
nand U44305 (N_44305,N_35646,N_31155);
xnor U44306 (N_44306,N_37380,N_34107);
and U44307 (N_44307,N_33326,N_37672);
or U44308 (N_44308,N_34271,N_37418);
nand U44309 (N_44309,N_31338,N_30682);
nor U44310 (N_44310,N_31148,N_35770);
xnor U44311 (N_44311,N_30672,N_31401);
nor U44312 (N_44312,N_33872,N_37409);
nand U44313 (N_44313,N_38124,N_32185);
or U44314 (N_44314,N_32272,N_32261);
nand U44315 (N_44315,N_31463,N_31613);
and U44316 (N_44316,N_31192,N_35668);
xor U44317 (N_44317,N_34362,N_34713);
or U44318 (N_44318,N_37627,N_30438);
xor U44319 (N_44319,N_34905,N_38824);
and U44320 (N_44320,N_33364,N_37525);
nand U44321 (N_44321,N_36877,N_32041);
nand U44322 (N_44322,N_32321,N_37564);
xor U44323 (N_44323,N_34618,N_30823);
and U44324 (N_44324,N_36296,N_38622);
and U44325 (N_44325,N_38441,N_31443);
xor U44326 (N_44326,N_33059,N_37694);
xor U44327 (N_44327,N_30998,N_33288);
and U44328 (N_44328,N_36855,N_30109);
and U44329 (N_44329,N_37752,N_36935);
nand U44330 (N_44330,N_39304,N_37130);
nand U44331 (N_44331,N_38442,N_34776);
xor U44332 (N_44332,N_31000,N_33091);
nor U44333 (N_44333,N_30708,N_33453);
xnor U44334 (N_44334,N_38216,N_37809);
or U44335 (N_44335,N_33560,N_36313);
xor U44336 (N_44336,N_37260,N_32952);
or U44337 (N_44337,N_35004,N_34307);
and U44338 (N_44338,N_32804,N_39306);
and U44339 (N_44339,N_36628,N_36766);
nand U44340 (N_44340,N_34768,N_33556);
or U44341 (N_44341,N_31543,N_33291);
nor U44342 (N_44342,N_37874,N_33205);
nand U44343 (N_44343,N_39539,N_38417);
and U44344 (N_44344,N_38992,N_32581);
xnor U44345 (N_44345,N_33767,N_39850);
xnor U44346 (N_44346,N_31747,N_35285);
and U44347 (N_44347,N_30019,N_39334);
nor U44348 (N_44348,N_33905,N_38705);
xnor U44349 (N_44349,N_39180,N_39664);
and U44350 (N_44350,N_35031,N_34255);
or U44351 (N_44351,N_32124,N_35457);
xnor U44352 (N_44352,N_36849,N_37594);
xor U44353 (N_44353,N_37299,N_39313);
nand U44354 (N_44354,N_39354,N_32275);
or U44355 (N_44355,N_39102,N_36412);
and U44356 (N_44356,N_35431,N_36764);
and U44357 (N_44357,N_32192,N_36770);
nand U44358 (N_44358,N_39852,N_32544);
xor U44359 (N_44359,N_38745,N_35243);
and U44360 (N_44360,N_37365,N_35536);
and U44361 (N_44361,N_34386,N_38089);
nor U44362 (N_44362,N_37745,N_36421);
xnor U44363 (N_44363,N_33923,N_34576);
xnor U44364 (N_44364,N_33331,N_33344);
nor U44365 (N_44365,N_36838,N_34995);
nand U44366 (N_44366,N_34103,N_37204);
nand U44367 (N_44367,N_34592,N_31818);
nand U44368 (N_44368,N_33074,N_36502);
or U44369 (N_44369,N_30363,N_36206);
and U44370 (N_44370,N_31590,N_34211);
or U44371 (N_44371,N_35886,N_38433);
nand U44372 (N_44372,N_32834,N_39473);
or U44373 (N_44373,N_31696,N_35499);
nand U44374 (N_44374,N_30668,N_34973);
xnor U44375 (N_44375,N_36505,N_36085);
xor U44376 (N_44376,N_33497,N_32827);
or U44377 (N_44377,N_37051,N_36788);
and U44378 (N_44378,N_39330,N_32835);
or U44379 (N_44379,N_37643,N_39800);
and U44380 (N_44380,N_34552,N_31728);
xnor U44381 (N_44381,N_38396,N_33255);
nor U44382 (N_44382,N_34938,N_36667);
xor U44383 (N_44383,N_39977,N_38381);
or U44384 (N_44384,N_37407,N_35829);
and U44385 (N_44385,N_33624,N_33261);
xor U44386 (N_44386,N_31968,N_32257);
or U44387 (N_44387,N_33167,N_32371);
xnor U44388 (N_44388,N_39844,N_30378);
and U44389 (N_44389,N_38552,N_37829);
nor U44390 (N_44390,N_35391,N_33209);
nand U44391 (N_44391,N_38623,N_36333);
xor U44392 (N_44392,N_33792,N_39958);
and U44393 (N_44393,N_32402,N_30504);
nand U44394 (N_44394,N_38717,N_30585);
nor U44395 (N_44395,N_39920,N_37314);
nor U44396 (N_44396,N_33642,N_36291);
nor U44397 (N_44397,N_32288,N_34140);
nor U44398 (N_44398,N_32029,N_37137);
xor U44399 (N_44399,N_31740,N_33129);
xor U44400 (N_44400,N_36769,N_31087);
nand U44401 (N_44401,N_33441,N_37325);
xor U44402 (N_44402,N_33154,N_39042);
nor U44403 (N_44403,N_35077,N_35533);
and U44404 (N_44404,N_36373,N_32251);
or U44405 (N_44405,N_30226,N_35432);
or U44406 (N_44406,N_35166,N_34968);
nor U44407 (N_44407,N_30353,N_34943);
or U44408 (N_44408,N_37711,N_33462);
nor U44409 (N_44409,N_35586,N_35920);
nor U44410 (N_44410,N_33352,N_31737);
and U44411 (N_44411,N_37837,N_38953);
nor U44412 (N_44412,N_36497,N_33574);
or U44413 (N_44413,N_39972,N_34031);
or U44414 (N_44414,N_30646,N_35152);
xnor U44415 (N_44415,N_33972,N_34712);
xor U44416 (N_44416,N_32975,N_39390);
and U44417 (N_44417,N_37749,N_39536);
nand U44418 (N_44418,N_35607,N_31839);
and U44419 (N_44419,N_34094,N_30792);
and U44420 (N_44420,N_30760,N_30569);
nand U44421 (N_44421,N_34626,N_32990);
and U44422 (N_44422,N_38545,N_38903);
xnor U44423 (N_44423,N_31843,N_32442);
nand U44424 (N_44424,N_39979,N_34590);
nor U44425 (N_44425,N_32130,N_39241);
nand U44426 (N_44426,N_34535,N_36033);
xor U44427 (N_44427,N_39074,N_35963);
and U44428 (N_44428,N_39115,N_36057);
and U44429 (N_44429,N_31572,N_38624);
and U44430 (N_44430,N_37600,N_32461);
nand U44431 (N_44431,N_35545,N_34166);
xnor U44432 (N_44432,N_31717,N_30961);
nand U44433 (N_44433,N_38014,N_38271);
nand U44434 (N_44434,N_38526,N_38954);
and U44435 (N_44435,N_37175,N_36397);
nor U44436 (N_44436,N_37742,N_31145);
nand U44437 (N_44437,N_36570,N_37072);
or U44438 (N_44438,N_39924,N_35165);
or U44439 (N_44439,N_38351,N_36945);
nand U44440 (N_44440,N_39479,N_38066);
and U44441 (N_44441,N_37297,N_34589);
nor U44442 (N_44442,N_39784,N_39178);
nand U44443 (N_44443,N_35169,N_37937);
or U44444 (N_44444,N_37171,N_39082);
nor U44445 (N_44445,N_36861,N_34417);
or U44446 (N_44446,N_39010,N_39421);
nor U44447 (N_44447,N_35398,N_30251);
nand U44448 (N_44448,N_38716,N_39582);
xnor U44449 (N_44449,N_31253,N_36170);
or U44450 (N_44450,N_36840,N_34283);
and U44451 (N_44451,N_39945,N_32168);
xor U44452 (N_44452,N_32898,N_36750);
and U44453 (N_44453,N_30968,N_34288);
xor U44454 (N_44454,N_34763,N_39500);
nand U44455 (N_44455,N_35330,N_38534);
or U44456 (N_44456,N_30158,N_32429);
xnor U44457 (N_44457,N_35281,N_39614);
or U44458 (N_44458,N_30785,N_30692);
nand U44459 (N_44459,N_37680,N_36913);
xor U44460 (N_44460,N_30875,N_31655);
or U44461 (N_44461,N_31400,N_38759);
xnor U44462 (N_44462,N_39436,N_30737);
nor U44463 (N_44463,N_33252,N_34723);
nor U44464 (N_44464,N_33776,N_34926);
or U44465 (N_44465,N_39865,N_38841);
xnor U44466 (N_44466,N_39864,N_39054);
xnor U44467 (N_44467,N_33305,N_32452);
or U44468 (N_44468,N_33569,N_38736);
xnor U44469 (N_44469,N_38945,N_35287);
xor U44470 (N_44470,N_37421,N_35149);
nor U44471 (N_44471,N_31385,N_30483);
nor U44472 (N_44472,N_39058,N_37016);
nor U44473 (N_44473,N_34499,N_30622);
or U44474 (N_44474,N_34070,N_36386);
nand U44475 (N_44475,N_38220,N_39404);
nor U44476 (N_44476,N_39853,N_35227);
nand U44477 (N_44477,N_30358,N_32137);
and U44478 (N_44478,N_36146,N_33005);
xnor U44479 (N_44479,N_36088,N_35280);
or U44480 (N_44480,N_32147,N_36579);
xnor U44481 (N_44481,N_39646,N_34917);
nor U44482 (N_44482,N_34682,N_36478);
or U44483 (N_44483,N_34415,N_31561);
or U44484 (N_44484,N_35259,N_32040);
xnor U44485 (N_44485,N_37603,N_39699);
nor U44486 (N_44486,N_37179,N_33108);
xnor U44487 (N_44487,N_38588,N_37765);
nor U44488 (N_44488,N_30262,N_38658);
or U44489 (N_44489,N_38484,N_34799);
nor U44490 (N_44490,N_31616,N_36931);
nand U44491 (N_44491,N_38358,N_36602);
nand U44492 (N_44492,N_33024,N_30696);
xor U44493 (N_44493,N_39515,N_33750);
nor U44494 (N_44494,N_32383,N_38525);
xnor U44495 (N_44495,N_37169,N_33153);
nand U44496 (N_44496,N_39585,N_34489);
nand U44497 (N_44497,N_31429,N_32562);
nand U44498 (N_44498,N_31113,N_33231);
or U44499 (N_44499,N_34743,N_38195);
nand U44500 (N_44500,N_37635,N_31979);
nor U44501 (N_44501,N_32617,N_35675);
nor U44502 (N_44502,N_39397,N_36467);
and U44503 (N_44503,N_31793,N_36585);
or U44504 (N_44504,N_35441,N_39933);
and U44505 (N_44505,N_37123,N_33143);
xnor U44506 (N_44506,N_39615,N_34819);
xor U44507 (N_44507,N_38335,N_36310);
xnor U44508 (N_44508,N_39659,N_38931);
xor U44509 (N_44509,N_35966,N_32511);
or U44510 (N_44510,N_35674,N_36556);
and U44511 (N_44511,N_33513,N_33038);
or U44512 (N_44512,N_31766,N_35325);
and U44513 (N_44513,N_33061,N_34058);
and U44514 (N_44514,N_35288,N_34290);
and U44515 (N_44515,N_38892,N_36201);
or U44516 (N_44516,N_36440,N_34837);
or U44517 (N_44517,N_34004,N_34690);
or U44518 (N_44518,N_30519,N_38686);
xnor U44519 (N_44519,N_30444,N_33401);
nand U44520 (N_44520,N_38693,N_39971);
or U44521 (N_44521,N_34272,N_30717);
xnor U44522 (N_44522,N_32078,N_37173);
xor U44523 (N_44523,N_34488,N_31948);
nor U44524 (N_44524,N_37193,N_36215);
or U44525 (N_44525,N_35608,N_36557);
and U44526 (N_44526,N_31093,N_36032);
and U44527 (N_44527,N_36051,N_38641);
nand U44528 (N_44528,N_32223,N_33748);
nor U44529 (N_44529,N_31074,N_36732);
and U44530 (N_44530,N_37659,N_30197);
nor U44531 (N_44531,N_38485,N_38201);
or U44532 (N_44532,N_30689,N_33976);
nand U44533 (N_44533,N_32877,N_31537);
nor U44534 (N_44534,N_35872,N_38311);
xnor U44535 (N_44535,N_37091,N_39035);
or U44536 (N_44536,N_31619,N_35979);
xor U44537 (N_44537,N_34546,N_33075);
xor U44538 (N_44538,N_35224,N_39444);
nor U44539 (N_44539,N_34747,N_37058);
xor U44540 (N_44540,N_33418,N_37585);
nor U44541 (N_44541,N_37391,N_34298);
xnor U44542 (N_44542,N_30340,N_39486);
or U44543 (N_44543,N_39917,N_30263);
and U44544 (N_44544,N_34216,N_36812);
nand U44545 (N_44545,N_30576,N_38384);
xnor U44546 (N_44546,N_34945,N_31181);
nor U44547 (N_44547,N_34795,N_35058);
and U44548 (N_44548,N_30897,N_32961);
or U44549 (N_44549,N_39095,N_32502);
xor U44550 (N_44550,N_33733,N_33166);
nand U44551 (N_44551,N_39915,N_39618);
xor U44552 (N_44552,N_30135,N_37251);
and U44553 (N_44553,N_38264,N_30527);
xor U44554 (N_44554,N_37298,N_32350);
nor U44555 (N_44555,N_38121,N_39856);
and U44556 (N_44556,N_39133,N_32806);
xor U44557 (N_44557,N_32191,N_38630);
or U44558 (N_44558,N_38239,N_33304);
or U44559 (N_44559,N_30244,N_34300);
xor U44560 (N_44560,N_30763,N_30375);
nand U44561 (N_44561,N_31803,N_33821);
nand U44562 (N_44562,N_32984,N_34568);
or U44563 (N_44563,N_37772,N_32560);
nor U44564 (N_44564,N_38075,N_35233);
nand U44565 (N_44565,N_39626,N_36604);
or U44566 (N_44566,N_38506,N_30586);
nand U44567 (N_44567,N_38153,N_38831);
nand U44568 (N_44568,N_31098,N_38721);
nor U44569 (N_44569,N_35617,N_31147);
xor U44570 (N_44570,N_34900,N_31589);
xor U44571 (N_44571,N_32912,N_31402);
xnor U44572 (N_44572,N_39088,N_39866);
or U44573 (N_44573,N_30074,N_34373);
nand U44574 (N_44574,N_31427,N_38680);
and U44575 (N_44575,N_38457,N_31210);
nand U44576 (N_44576,N_31034,N_34869);
and U44577 (N_44577,N_30588,N_36608);
or U44578 (N_44578,N_37685,N_38808);
and U44579 (N_44579,N_31514,N_30604);
nand U44580 (N_44580,N_39096,N_32141);
xnor U44581 (N_44581,N_31823,N_35272);
xor U44582 (N_44582,N_39891,N_39689);
xor U44583 (N_44583,N_36261,N_32576);
xor U44584 (N_44584,N_32753,N_34542);
and U44585 (N_44585,N_30028,N_37576);
nor U44586 (N_44586,N_32967,N_37034);
nand U44587 (N_44587,N_33062,N_33963);
nand U44588 (N_44588,N_30480,N_32252);
xor U44589 (N_44589,N_35046,N_33965);
nand U44590 (N_44590,N_37587,N_38134);
and U44591 (N_44591,N_35483,N_30883);
nand U44592 (N_44592,N_31011,N_32805);
nor U44593 (N_44593,N_33835,N_34722);
or U44594 (N_44594,N_39210,N_35563);
and U44595 (N_44595,N_30160,N_34754);
or U44596 (N_44596,N_33925,N_38225);
or U44597 (N_44597,N_37788,N_34728);
or U44598 (N_44598,N_33051,N_38919);
or U44599 (N_44599,N_39658,N_36233);
xor U44600 (N_44600,N_38386,N_35275);
nor U44601 (N_44601,N_30157,N_30725);
or U44602 (N_44602,N_35042,N_38055);
xor U44603 (N_44603,N_33021,N_36415);
or U44604 (N_44604,N_38765,N_34753);
and U44605 (N_44605,N_37425,N_36767);
nand U44606 (N_44606,N_35725,N_34349);
xor U44607 (N_44607,N_36364,N_31531);
nand U44608 (N_44608,N_31243,N_34297);
nand U44609 (N_44609,N_31241,N_31646);
xor U44610 (N_44610,N_33664,N_35164);
xnor U44611 (N_44611,N_30386,N_30908);
nand U44612 (N_44612,N_35775,N_31663);
nor U44613 (N_44613,N_38728,N_36197);
nor U44614 (N_44614,N_39540,N_34649);
nor U44615 (N_44615,N_32578,N_31566);
nand U44616 (N_44616,N_38896,N_36582);
xor U44617 (N_44617,N_33959,N_34145);
nor U44618 (N_44618,N_37244,N_39456);
and U44619 (N_44619,N_35981,N_31975);
and U44620 (N_44620,N_37147,N_38839);
nor U44621 (N_44621,N_34219,N_37267);
nand U44622 (N_44622,N_39564,N_35438);
nor U44623 (N_44623,N_34414,N_33618);
nor U44624 (N_44624,N_32434,N_31588);
and U44625 (N_44625,N_36140,N_30967);
nor U44626 (N_44626,N_30229,N_33427);
and U44627 (N_44627,N_39029,N_36244);
nand U44628 (N_44628,N_36015,N_30396);
nor U44629 (N_44629,N_39426,N_39269);
nand U44630 (N_44630,N_31334,N_38604);
nand U44631 (N_44631,N_39149,N_34055);
or U44632 (N_44632,N_36630,N_39434);
and U44633 (N_44633,N_39630,N_30101);
nor U44634 (N_44634,N_34540,N_31976);
nand U44635 (N_44635,N_36175,N_36564);
xnor U44636 (N_44636,N_32197,N_33428);
and U44637 (N_44637,N_30776,N_33110);
or U44638 (N_44638,N_38825,N_34301);
nor U44639 (N_44639,N_35708,N_31444);
nand U44640 (N_44640,N_37785,N_34844);
nor U44641 (N_44641,N_39968,N_36878);
nor U44642 (N_44642,N_36258,N_35463);
and U44643 (N_44643,N_39793,N_30901);
and U44644 (N_44644,N_35018,N_34909);
or U44645 (N_44645,N_39575,N_39257);
and U44646 (N_44646,N_39809,N_38243);
xor U44647 (N_44647,N_35066,N_38989);
and U44648 (N_44648,N_33753,N_30954);
xnor U44649 (N_44649,N_37131,N_36642);
nor U44650 (N_44650,N_31951,N_34596);
nor U44651 (N_44651,N_36713,N_32385);
nand U44652 (N_44652,N_31861,N_37435);
nand U44653 (N_44653,N_32100,N_31901);
nor U44654 (N_44654,N_32934,N_30844);
nand U44655 (N_44655,N_33466,N_35712);
xnor U44656 (N_44656,N_39123,N_34796);
nor U44657 (N_44657,N_33845,N_30837);
xnor U44658 (N_44658,N_39769,N_37793);
xnor U44659 (N_44659,N_32113,N_31149);
and U44660 (N_44660,N_33037,N_30891);
or U44661 (N_44661,N_35994,N_36169);
nor U44662 (N_44662,N_36110,N_33290);
and U44663 (N_44663,N_34486,N_30726);
or U44664 (N_44664,N_37224,N_37077);
and U44665 (N_44665,N_36857,N_39009);
xnor U44666 (N_44666,N_34655,N_33875);
nand U44667 (N_44667,N_33370,N_32678);
nand U44668 (N_44668,N_34248,N_37878);
nor U44669 (N_44669,N_35878,N_32196);
nand U44670 (N_44670,N_34303,N_37699);
nor U44671 (N_44671,N_33555,N_30944);
nand U44672 (N_44672,N_34473,N_34922);
xor U44673 (N_44673,N_33817,N_35109);
or U44674 (N_44674,N_32608,N_33457);
and U44675 (N_44675,N_30951,N_37543);
nor U44676 (N_44676,N_35298,N_39469);
and U44677 (N_44677,N_34516,N_34860);
xnor U44678 (N_44678,N_31488,N_34569);
or U44679 (N_44679,N_36982,N_37727);
or U44680 (N_44680,N_34672,N_36280);
nand U44681 (N_44681,N_34196,N_33651);
or U44682 (N_44682,N_37640,N_30493);
or U44683 (N_44683,N_36243,N_37355);
and U44684 (N_44684,N_32325,N_39705);
nor U44685 (N_44685,N_32503,N_36571);
xor U44686 (N_44686,N_33984,N_30159);
and U44687 (N_44687,N_36256,N_35894);
nor U44688 (N_44688,N_38284,N_34392);
or U44689 (N_44689,N_36394,N_35832);
and U44690 (N_44690,N_32379,N_31106);
nor U44691 (N_44691,N_36276,N_39842);
xnor U44692 (N_44692,N_39053,N_31782);
nor U44693 (N_44693,N_35101,N_33670);
xor U44694 (N_44694,N_35804,N_33289);
nand U44695 (N_44695,N_36241,N_39152);
nor U44696 (N_44696,N_38105,N_39826);
nor U44697 (N_44697,N_33999,N_31612);
nand U44698 (N_44698,N_30437,N_32110);
and U44699 (N_44699,N_37889,N_37015);
or U44700 (N_44700,N_33692,N_30768);
nor U44701 (N_44701,N_37743,N_32654);
nand U44702 (N_44702,N_30849,N_32723);
nand U44703 (N_44703,N_38866,N_31917);
nor U44704 (N_44704,N_30471,N_36692);
and U44705 (N_44705,N_38948,N_36521);
nor U44706 (N_44706,N_38737,N_37195);
nand U44707 (N_44707,N_39023,N_35038);
nand U44708 (N_44708,N_30248,N_37255);
and U44709 (N_44709,N_34812,N_32395);
nand U44710 (N_44710,N_39460,N_37102);
xor U44711 (N_44711,N_36255,N_38059);
nor U44712 (N_44712,N_31284,N_33782);
xnor U44713 (N_44713,N_34981,N_37542);
nor U44714 (N_44714,N_37835,N_31773);
nor U44715 (N_44715,N_34639,N_32832);
nand U44716 (N_44716,N_34232,N_37280);
and U44717 (N_44717,N_38182,N_31888);
and U44718 (N_44718,N_36430,N_37523);
nand U44719 (N_44719,N_37804,N_37998);
nor U44720 (N_44720,N_34450,N_37158);
and U44721 (N_44721,N_31609,N_33018);
nor U44722 (N_44722,N_37784,N_38885);
or U44723 (N_44723,N_38252,N_32406);
nand U44724 (N_44724,N_33545,N_36120);
or U44725 (N_44725,N_33101,N_33619);
and U44726 (N_44726,N_36848,N_37830);
nor U44727 (N_44727,N_35141,N_32396);
xnor U44728 (N_44728,N_30130,N_31523);
xor U44729 (N_44729,N_38202,N_36672);
or U44730 (N_44730,N_36629,N_35435);
nor U44731 (N_44731,N_36290,N_32828);
or U44732 (N_44732,N_33302,N_33790);
or U44733 (N_44733,N_30206,N_34481);
and U44734 (N_44734,N_38211,N_37483);
nand U44735 (N_44735,N_31878,N_30189);
nor U44736 (N_44736,N_36894,N_30070);
xor U44737 (N_44737,N_38941,N_34105);
nor U44738 (N_44738,N_35641,N_32446);
xnor U44739 (N_44739,N_35388,N_39166);
or U44740 (N_44740,N_39064,N_33156);
xnor U44741 (N_44741,N_37020,N_37026);
or U44742 (N_44742,N_33548,N_38984);
nor U44743 (N_44743,N_35235,N_33774);
nand U44744 (N_44744,N_38998,N_36315);
xor U44745 (N_44745,N_32850,N_31169);
or U44746 (N_44746,N_39874,N_30724);
xor U44747 (N_44747,N_38142,N_38580);
nand U44748 (N_44748,N_32541,N_36115);
nor U44749 (N_44749,N_30076,N_38877);
nand U44750 (N_44750,N_34667,N_38348);
nor U44751 (N_44751,N_30971,N_37828);
xor U44752 (N_44752,N_34332,N_36754);
nand U44753 (N_44753,N_33172,N_34518);
and U44754 (N_44754,N_30539,N_36972);
xor U44755 (N_44755,N_30602,N_31143);
and U44756 (N_44756,N_36231,N_37466);
and U44757 (N_44757,N_35697,N_39878);
and U44758 (N_44758,N_36300,N_30783);
or U44759 (N_44759,N_32455,N_32188);
and U44760 (N_44760,N_31767,N_38898);
and U44761 (N_44761,N_39989,N_32212);
or U44762 (N_44762,N_38212,N_39683);
nor U44763 (N_44763,N_35809,N_39681);
xor U44764 (N_44764,N_38852,N_39612);
nand U44765 (N_44765,N_38743,N_30087);
and U44766 (N_44766,N_34789,N_30637);
nand U44767 (N_44767,N_36528,N_34312);
nor U44768 (N_44768,N_32393,N_36381);
and U44769 (N_44769,N_36736,N_30541);
nand U44770 (N_44770,N_35864,N_39796);
nor U44771 (N_44771,N_31175,N_33477);
and U44772 (N_44772,N_35932,N_39016);
nor U44773 (N_44773,N_35568,N_33929);
or U44774 (N_44774,N_36671,N_35579);
or U44775 (N_44775,N_34600,N_32042);
xnor U44776 (N_44776,N_36164,N_31835);
or U44777 (N_44777,N_37530,N_34274);
or U44778 (N_44778,N_35771,N_36221);
xor U44779 (N_44779,N_30914,N_36561);
nand U44780 (N_44780,N_31019,N_38401);
xnor U44781 (N_44781,N_33666,N_36147);
and U44782 (N_44782,N_36791,N_30913);
or U44783 (N_44783,N_34912,N_32848);
nor U44784 (N_44784,N_37070,N_30747);
nand U44785 (N_44785,N_36389,N_37552);
nand U44786 (N_44786,N_39358,N_33054);
nor U44787 (N_44787,N_37410,N_35286);
nand U44788 (N_44788,N_36324,N_30382);
xnor U44789 (N_44789,N_39156,N_32881);
xor U44790 (N_44790,N_36719,N_33379);
or U44791 (N_44791,N_36929,N_37291);
xor U44792 (N_44792,N_39955,N_37028);
and U44793 (N_44793,N_38907,N_31375);
nand U44794 (N_44794,N_31010,N_31185);
nor U44795 (N_44795,N_31297,N_30395);
nand U44796 (N_44796,N_34852,N_39060);
and U44797 (N_44797,N_33384,N_32346);
xnor U44798 (N_44798,N_35375,N_35178);
and U44799 (N_44799,N_34160,N_37499);
or U44800 (N_44800,N_38802,N_35253);
nor U44801 (N_44801,N_32679,N_34188);
nor U44802 (N_44802,N_36340,N_30295);
nand U44803 (N_44803,N_33050,N_36176);
nand U44804 (N_44804,N_39571,N_38443);
nand U44805 (N_44805,N_31671,N_34265);
and U44806 (N_44806,N_30791,N_34021);
xor U44807 (N_44807,N_32706,N_32751);
nand U44808 (N_44808,N_37732,N_38962);
xor U44809 (N_44809,N_33632,N_37369);
or U44810 (N_44810,N_34342,N_38509);
or U44811 (N_44811,N_36647,N_39002);
nor U44812 (N_44812,N_35041,N_33373);
and U44813 (N_44813,N_31656,N_32809);
nor U44814 (N_44814,N_31779,N_33968);
and U44815 (N_44815,N_36495,N_34954);
or U44816 (N_44816,N_35810,N_38315);
and U44817 (N_44817,N_32852,N_34565);
nand U44818 (N_44818,N_30138,N_31568);
and U44819 (N_44819,N_35924,N_32675);
nand U44820 (N_44820,N_35142,N_31484);
and U44821 (N_44821,N_34496,N_38078);
and U44822 (N_44822,N_39701,N_30446);
or U44823 (N_44823,N_31177,N_30410);
or U44824 (N_44824,N_36037,N_33977);
xnor U44825 (N_44825,N_39558,N_35158);
xor U44826 (N_44826,N_31036,N_36803);
nor U44827 (N_44827,N_34647,N_39667);
nor U44828 (N_44828,N_33784,N_35476);
nand U44829 (N_44829,N_30060,N_35168);
nor U44830 (N_44830,N_37209,N_37623);
nand U44831 (N_44831,N_33995,N_32077);
and U44832 (N_44832,N_31689,N_36562);
nand U44833 (N_44833,N_38669,N_32448);
or U44834 (N_44834,N_33696,N_38538);
and U44835 (N_44835,N_36132,N_31278);
or U44836 (N_44836,N_35709,N_37363);
and U44837 (N_44837,N_33786,N_34256);
nor U44838 (N_44838,N_31403,N_34891);
nand U44839 (N_44839,N_39947,N_30734);
nand U44840 (N_44840,N_35151,N_31054);
nand U44841 (N_44841,N_34988,N_34076);
or U44842 (N_44842,N_33224,N_36678);
nand U44843 (N_44843,N_34411,N_30651);
and U44844 (N_44844,N_31775,N_32140);
and U44845 (N_44845,N_33901,N_39507);
nor U44846 (N_44846,N_31577,N_30107);
nor U44847 (N_44847,N_39579,N_34859);
or U44848 (N_44848,N_30994,N_32399);
xor U44849 (N_44849,N_38071,N_31863);
nand U44850 (N_44850,N_38991,N_32517);
nand U44851 (N_44851,N_31558,N_30088);
nor U44852 (N_44852,N_35927,N_31525);
nand U44853 (N_44853,N_34250,N_36673);
nand U44854 (N_44854,N_30743,N_34834);
nor U44855 (N_44855,N_35464,N_38031);
nand U44856 (N_44856,N_31817,N_33367);
nor U44857 (N_44857,N_31505,N_36632);
nand U44858 (N_44858,N_30105,N_39144);
nor U44859 (N_44859,N_38181,N_31020);
and U44860 (N_44860,N_36809,N_31749);
nor U44861 (N_44861,N_38857,N_34897);
nand U44862 (N_44862,N_34984,N_33402);
or U44863 (N_44863,N_37517,N_35323);
nor U44864 (N_44864,N_39312,N_36924);
nor U44865 (N_44865,N_39325,N_38521);
nor U44866 (N_44866,N_34640,N_35313);
nor U44867 (N_44867,N_33787,N_36029);
nand U44868 (N_44868,N_34176,N_36890);
nor U44869 (N_44869,N_36772,N_33998);
xor U44870 (N_44870,N_39489,N_35406);
xnor U44871 (N_44871,N_35576,N_30370);
and U44872 (N_44872,N_31544,N_32802);
xnor U44873 (N_44873,N_30077,N_32558);
nor U44874 (N_44874,N_38785,N_37747);
nand U44875 (N_44875,N_33575,N_39963);
nand U44876 (N_44876,N_38218,N_30801);
nand U44877 (N_44877,N_39774,N_39119);
nor U44878 (N_44878,N_30172,N_33121);
nor U44879 (N_44879,N_38244,N_30460);
nor U44880 (N_44880,N_39706,N_30649);
or U44881 (N_44881,N_37799,N_31295);
nand U44882 (N_44882,N_30393,N_32931);
xor U44883 (N_44883,N_31006,N_36317);
or U44884 (N_44884,N_34194,N_39424);
and U44885 (N_44885,N_39420,N_32719);
xor U44886 (N_44886,N_38837,N_30152);
nor U44887 (N_44887,N_31547,N_38126);
nor U44888 (N_44888,N_38154,N_33944);
xnor U44889 (N_44889,N_37602,N_39956);
nor U44890 (N_44890,N_33798,N_33586);
nor U44891 (N_44891,N_36874,N_34029);
nor U44892 (N_44892,N_30507,N_36682);
and U44893 (N_44893,N_38061,N_36897);
or U44894 (N_44894,N_30081,N_31875);
nand U44895 (N_44895,N_30733,N_33227);
or U44896 (N_44896,N_32083,N_34404);
and U44897 (N_44897,N_36473,N_30474);
or U44898 (N_44898,N_35137,N_33660);
or U44899 (N_44899,N_37932,N_35479);
nand U44900 (N_44900,N_30193,N_32481);
and U44901 (N_44901,N_38302,N_36859);
nand U44902 (N_44902,N_30530,N_33590);
nor U44903 (N_44903,N_36131,N_36725);
nand U44904 (N_44904,N_32225,N_37294);
or U44905 (N_44905,N_33210,N_35148);
or U44906 (N_44906,N_35105,N_35482);
and U44907 (N_44907,N_33739,N_37549);
nor U44908 (N_44908,N_33842,N_36302);
and U44909 (N_44909,N_38594,N_37235);
nand U44910 (N_44910,N_37853,N_39832);
nand U44911 (N_44911,N_36129,N_34630);
nor U44912 (N_44912,N_35238,N_34273);
and U44913 (N_44913,N_39472,N_35846);
nor U44914 (N_44914,N_33621,N_38322);
and U44915 (N_44915,N_35123,N_36130);
xor U44916 (N_44916,N_37296,N_39386);
nand U44917 (N_44917,N_36756,N_35613);
nand U44918 (N_44918,N_31194,N_38459);
or U44919 (N_44919,N_30605,N_33242);
or U44920 (N_44920,N_32381,N_32768);
or U44921 (N_44921,N_37520,N_33634);
nand U44922 (N_44922,N_30315,N_32776);
xor U44923 (N_44923,N_33973,N_35799);
and U44924 (N_44924,N_37695,N_36448);
or U44925 (N_44925,N_34206,N_38797);
or U44926 (N_44926,N_38266,N_33933);
nor U44927 (N_44927,N_37987,N_31915);
nor U44928 (N_44928,N_38147,N_31781);
or U44929 (N_44929,N_36488,N_37821);
nand U44930 (N_44930,N_33257,N_36995);
nor U44931 (N_44931,N_39510,N_36789);
xnor U44932 (N_44932,N_37986,N_39825);
xor U44933 (N_44933,N_35372,N_34816);
xnor U44934 (N_44934,N_35540,N_39164);
or U44935 (N_44935,N_39028,N_36178);
nand U44936 (N_44936,N_31235,N_31891);
nor U44937 (N_44937,N_30029,N_39901);
xor U44938 (N_44938,N_37222,N_35363);
nor U44939 (N_44939,N_35112,N_37043);
and U44940 (N_44940,N_33488,N_36081);
and U44941 (N_44941,N_36983,N_38584);
nand U44942 (N_44942,N_32388,N_38356);
and U44943 (N_44943,N_30050,N_39835);
nor U44944 (N_44944,N_38395,N_31784);
and U44945 (N_44945,N_33313,N_33605);
nand U44946 (N_44946,N_35321,N_31575);
xor U44947 (N_44947,N_37382,N_37740);
nand U44948 (N_44948,N_39952,N_33914);
nor U44949 (N_44949,N_33116,N_39997);
or U44950 (N_44950,N_30054,N_36271);
nor U44951 (N_44951,N_34164,N_38644);
and U44952 (N_44952,N_35507,N_34087);
xnor U44953 (N_44953,N_36984,N_34147);
and U44954 (N_44954,N_37902,N_36040);
nand U44955 (N_44955,N_30782,N_39959);
or U44956 (N_44956,N_37153,N_35410);
nor U44957 (N_44957,N_34883,N_31610);
or U44958 (N_44958,N_31161,N_36171);
nor U44959 (N_44959,N_38621,N_32462);
nand U44960 (N_44960,N_39845,N_33351);
or U44961 (N_44961,N_32374,N_33992);
and U44962 (N_44962,N_37379,N_32977);
or U44963 (N_44963,N_31983,N_34788);
nor U44964 (N_44964,N_32175,N_30697);
nand U44965 (N_44965,N_35304,N_35072);
xnor U44966 (N_44966,N_34811,N_38467);
and U44967 (N_44967,N_38924,N_38750);
nand U44968 (N_44968,N_36214,N_34503);
xnor U44969 (N_44969,N_35317,N_33994);
nor U44970 (N_44970,N_39684,N_36523);
nand U44971 (N_44971,N_34865,N_34942);
nand U44972 (N_44972,N_30684,N_34483);
and U44973 (N_44973,N_35546,N_33184);
nand U44974 (N_44974,N_32486,N_31660);
and U44975 (N_44975,N_37770,N_36107);
or U44976 (N_44976,N_38744,N_36889);
or U44977 (N_44977,N_30629,N_35026);
or U44978 (N_44978,N_37093,N_32935);
or U44979 (N_44979,N_36533,N_35818);
nand U44980 (N_44980,N_35634,N_39171);
nor U44981 (N_44981,N_38505,N_36275);
nor U44982 (N_44982,N_34899,N_30485);
or U44983 (N_44983,N_39818,N_35916);
nand U44984 (N_44984,N_39499,N_37120);
nor U44985 (N_44985,N_37229,N_33085);
xnor U44986 (N_44986,N_38205,N_32506);
nand U44987 (N_44987,N_39859,N_34035);
nand U44988 (N_44988,N_30241,N_35701);
and U44989 (N_44989,N_30550,N_37271);
and U44990 (N_44990,N_32226,N_33450);
xnor U44991 (N_44991,N_37933,N_37953);
nand U44992 (N_44992,N_30094,N_35248);
or U44993 (N_44993,N_38767,N_30650);
nor U44994 (N_44994,N_32496,N_33738);
xnor U44995 (N_44995,N_32740,N_34800);
xnor U44996 (N_44996,N_33140,N_30283);
or U44997 (N_44997,N_39633,N_30429);
and U44998 (N_44998,N_32071,N_31250);
and U44999 (N_44999,N_31853,N_36061);
xor U45000 (N_45000,N_35726,N_30292);
nor U45001 (N_45001,N_31400,N_30195);
nand U45002 (N_45002,N_36485,N_30878);
nor U45003 (N_45003,N_36151,N_31693);
xor U45004 (N_45004,N_33246,N_38556);
nand U45005 (N_45005,N_36590,N_32906);
nor U45006 (N_45006,N_37899,N_37819);
nand U45007 (N_45007,N_36178,N_33977);
nor U45008 (N_45008,N_32785,N_32339);
or U45009 (N_45009,N_39705,N_36526);
xnor U45010 (N_45010,N_33071,N_34319);
and U45011 (N_45011,N_37797,N_31186);
nor U45012 (N_45012,N_32240,N_31775);
nor U45013 (N_45013,N_37462,N_39429);
and U45014 (N_45014,N_38986,N_38542);
nor U45015 (N_45015,N_36014,N_38489);
and U45016 (N_45016,N_33553,N_36345);
xor U45017 (N_45017,N_34509,N_38807);
nand U45018 (N_45018,N_37134,N_34072);
xnor U45019 (N_45019,N_31328,N_36362);
nand U45020 (N_45020,N_31729,N_33652);
and U45021 (N_45021,N_35287,N_36715);
nand U45022 (N_45022,N_33614,N_38823);
or U45023 (N_45023,N_35256,N_37752);
xnor U45024 (N_45024,N_32632,N_30168);
xor U45025 (N_45025,N_35609,N_31077);
or U45026 (N_45026,N_37728,N_39658);
nor U45027 (N_45027,N_32205,N_38037);
xnor U45028 (N_45028,N_34084,N_35847);
nand U45029 (N_45029,N_34499,N_31404);
xor U45030 (N_45030,N_36025,N_35157);
and U45031 (N_45031,N_35548,N_39529);
nand U45032 (N_45032,N_33000,N_36145);
and U45033 (N_45033,N_37725,N_39717);
nor U45034 (N_45034,N_36932,N_31195);
nor U45035 (N_45035,N_33928,N_36182);
xnor U45036 (N_45036,N_33812,N_33142);
xor U45037 (N_45037,N_31282,N_38709);
nor U45038 (N_45038,N_39285,N_31523);
and U45039 (N_45039,N_35203,N_36527);
nor U45040 (N_45040,N_31226,N_37597);
nand U45041 (N_45041,N_34972,N_36715);
xnor U45042 (N_45042,N_34820,N_33501);
nor U45043 (N_45043,N_36619,N_32155);
nand U45044 (N_45044,N_31117,N_35610);
nand U45045 (N_45045,N_35141,N_32516);
xnor U45046 (N_45046,N_34120,N_32287);
nand U45047 (N_45047,N_30703,N_36952);
and U45048 (N_45048,N_39289,N_34089);
nor U45049 (N_45049,N_32931,N_35544);
xnor U45050 (N_45050,N_30570,N_34833);
or U45051 (N_45051,N_33012,N_38126);
xor U45052 (N_45052,N_36019,N_38169);
nor U45053 (N_45053,N_33698,N_31832);
nor U45054 (N_45054,N_33854,N_36287);
xnor U45055 (N_45055,N_37012,N_37171);
nand U45056 (N_45056,N_39037,N_31676);
nor U45057 (N_45057,N_39597,N_31996);
or U45058 (N_45058,N_33082,N_35645);
nor U45059 (N_45059,N_31984,N_35599);
or U45060 (N_45060,N_30796,N_34223);
nand U45061 (N_45061,N_39003,N_34930);
xor U45062 (N_45062,N_36873,N_30724);
xnor U45063 (N_45063,N_33242,N_31532);
or U45064 (N_45064,N_35133,N_30711);
nand U45065 (N_45065,N_34145,N_37411);
xnor U45066 (N_45066,N_35185,N_37772);
nand U45067 (N_45067,N_36788,N_36595);
nor U45068 (N_45068,N_38231,N_36847);
or U45069 (N_45069,N_33495,N_34923);
xnor U45070 (N_45070,N_37794,N_35780);
or U45071 (N_45071,N_33819,N_32971);
xnor U45072 (N_45072,N_33401,N_38325);
or U45073 (N_45073,N_34619,N_30434);
or U45074 (N_45074,N_32525,N_38161);
nor U45075 (N_45075,N_31375,N_31396);
or U45076 (N_45076,N_34071,N_34201);
xor U45077 (N_45077,N_32182,N_37154);
and U45078 (N_45078,N_37213,N_39887);
xnor U45079 (N_45079,N_32861,N_30211);
or U45080 (N_45080,N_31744,N_33807);
nor U45081 (N_45081,N_33970,N_34166);
xor U45082 (N_45082,N_36236,N_30960);
xnor U45083 (N_45083,N_34077,N_37964);
nor U45084 (N_45084,N_35950,N_32161);
nor U45085 (N_45085,N_34179,N_30419);
or U45086 (N_45086,N_35672,N_38707);
or U45087 (N_45087,N_31790,N_33662);
xor U45088 (N_45088,N_32400,N_36360);
nand U45089 (N_45089,N_34518,N_30308);
xnor U45090 (N_45090,N_38595,N_35388);
xor U45091 (N_45091,N_37115,N_38230);
nand U45092 (N_45092,N_38860,N_35201);
xnor U45093 (N_45093,N_33422,N_31201);
or U45094 (N_45094,N_30155,N_31515);
or U45095 (N_45095,N_34766,N_36011);
or U45096 (N_45096,N_39721,N_34873);
and U45097 (N_45097,N_32503,N_36629);
or U45098 (N_45098,N_34379,N_35934);
or U45099 (N_45099,N_38167,N_31814);
nor U45100 (N_45100,N_37247,N_34783);
nor U45101 (N_45101,N_38444,N_30368);
or U45102 (N_45102,N_35957,N_30923);
xor U45103 (N_45103,N_39981,N_30962);
nor U45104 (N_45104,N_36184,N_33786);
xnor U45105 (N_45105,N_31025,N_32575);
nand U45106 (N_45106,N_35314,N_36310);
or U45107 (N_45107,N_39651,N_37890);
and U45108 (N_45108,N_36101,N_30931);
nand U45109 (N_45109,N_32597,N_38617);
and U45110 (N_45110,N_36800,N_39369);
nor U45111 (N_45111,N_34749,N_34401);
or U45112 (N_45112,N_33155,N_37996);
xnor U45113 (N_45113,N_35341,N_39738);
nand U45114 (N_45114,N_35477,N_37804);
or U45115 (N_45115,N_33494,N_33749);
nand U45116 (N_45116,N_38860,N_32424);
nor U45117 (N_45117,N_30870,N_35145);
or U45118 (N_45118,N_32019,N_39243);
nand U45119 (N_45119,N_33814,N_30494);
or U45120 (N_45120,N_38971,N_33080);
or U45121 (N_45121,N_39120,N_30289);
nand U45122 (N_45122,N_38382,N_39786);
xnor U45123 (N_45123,N_33377,N_38131);
nor U45124 (N_45124,N_32324,N_35953);
or U45125 (N_45125,N_37500,N_33360);
and U45126 (N_45126,N_33584,N_33798);
and U45127 (N_45127,N_33032,N_39461);
and U45128 (N_45128,N_32027,N_35636);
xnor U45129 (N_45129,N_32605,N_37239);
or U45130 (N_45130,N_38645,N_35361);
xnor U45131 (N_45131,N_30304,N_39126);
nor U45132 (N_45132,N_30363,N_31294);
and U45133 (N_45133,N_38655,N_33486);
nor U45134 (N_45134,N_35923,N_37783);
nor U45135 (N_45135,N_36966,N_37343);
nor U45136 (N_45136,N_39200,N_36026);
nor U45137 (N_45137,N_31185,N_36270);
nand U45138 (N_45138,N_33083,N_30624);
or U45139 (N_45139,N_36577,N_34792);
nand U45140 (N_45140,N_36399,N_32755);
and U45141 (N_45141,N_39132,N_33280);
nor U45142 (N_45142,N_32016,N_32683);
or U45143 (N_45143,N_38866,N_37619);
nor U45144 (N_45144,N_34103,N_31981);
nand U45145 (N_45145,N_33035,N_36005);
nor U45146 (N_45146,N_38579,N_33273);
nor U45147 (N_45147,N_30520,N_38656);
and U45148 (N_45148,N_32408,N_32290);
or U45149 (N_45149,N_38543,N_34123);
and U45150 (N_45150,N_32001,N_37036);
nand U45151 (N_45151,N_34248,N_32014);
xor U45152 (N_45152,N_39825,N_39695);
or U45153 (N_45153,N_33296,N_36807);
nand U45154 (N_45154,N_35641,N_31260);
xnor U45155 (N_45155,N_30120,N_32777);
and U45156 (N_45156,N_39467,N_38882);
and U45157 (N_45157,N_33527,N_37355);
and U45158 (N_45158,N_31419,N_30661);
nand U45159 (N_45159,N_35707,N_35852);
nor U45160 (N_45160,N_34657,N_39150);
or U45161 (N_45161,N_34799,N_32234);
nand U45162 (N_45162,N_33120,N_34228);
or U45163 (N_45163,N_31072,N_37807);
and U45164 (N_45164,N_33320,N_30758);
and U45165 (N_45165,N_37058,N_39973);
nand U45166 (N_45166,N_36323,N_30735);
nor U45167 (N_45167,N_30455,N_32304);
or U45168 (N_45168,N_32617,N_38780);
xor U45169 (N_45169,N_34234,N_33200);
or U45170 (N_45170,N_30572,N_39494);
xnor U45171 (N_45171,N_30420,N_36512);
nand U45172 (N_45172,N_35167,N_30763);
xnor U45173 (N_45173,N_30887,N_32383);
nand U45174 (N_45174,N_31349,N_36570);
or U45175 (N_45175,N_35385,N_39984);
nor U45176 (N_45176,N_30108,N_38724);
nand U45177 (N_45177,N_38777,N_37837);
nand U45178 (N_45178,N_33415,N_33421);
nand U45179 (N_45179,N_32132,N_36896);
nor U45180 (N_45180,N_33979,N_36189);
xnor U45181 (N_45181,N_35843,N_32215);
nand U45182 (N_45182,N_32861,N_38012);
nand U45183 (N_45183,N_36685,N_30140);
xor U45184 (N_45184,N_37105,N_30248);
nand U45185 (N_45185,N_31176,N_35159);
nor U45186 (N_45186,N_37513,N_32248);
xnor U45187 (N_45187,N_30585,N_35025);
or U45188 (N_45188,N_32160,N_32985);
xnor U45189 (N_45189,N_32185,N_38367);
nand U45190 (N_45190,N_38169,N_36594);
xor U45191 (N_45191,N_32489,N_36599);
or U45192 (N_45192,N_38752,N_39754);
nand U45193 (N_45193,N_32378,N_33109);
xor U45194 (N_45194,N_34648,N_33163);
nor U45195 (N_45195,N_31097,N_35865);
or U45196 (N_45196,N_33043,N_31602);
nand U45197 (N_45197,N_38404,N_30010);
xnor U45198 (N_45198,N_37194,N_36005);
xnor U45199 (N_45199,N_33273,N_32693);
or U45200 (N_45200,N_32877,N_36828);
nor U45201 (N_45201,N_33256,N_33240);
or U45202 (N_45202,N_30218,N_33820);
nand U45203 (N_45203,N_37525,N_38958);
nand U45204 (N_45204,N_36607,N_31463);
and U45205 (N_45205,N_37598,N_36044);
nor U45206 (N_45206,N_37071,N_34043);
and U45207 (N_45207,N_34055,N_38278);
nand U45208 (N_45208,N_32309,N_37163);
nand U45209 (N_45209,N_32243,N_33018);
or U45210 (N_45210,N_34150,N_37890);
nor U45211 (N_45211,N_36860,N_33306);
or U45212 (N_45212,N_34859,N_38097);
xor U45213 (N_45213,N_37412,N_31540);
xor U45214 (N_45214,N_31311,N_31134);
nand U45215 (N_45215,N_35803,N_30680);
nor U45216 (N_45216,N_31463,N_32826);
xnor U45217 (N_45217,N_35592,N_30508);
nor U45218 (N_45218,N_33599,N_30315);
nand U45219 (N_45219,N_37036,N_33811);
nor U45220 (N_45220,N_36490,N_39618);
or U45221 (N_45221,N_36130,N_31163);
xor U45222 (N_45222,N_33868,N_33273);
nand U45223 (N_45223,N_31556,N_36054);
nand U45224 (N_45224,N_32768,N_37451);
or U45225 (N_45225,N_31226,N_35867);
nor U45226 (N_45226,N_34535,N_31669);
nor U45227 (N_45227,N_32535,N_33659);
xnor U45228 (N_45228,N_31158,N_32879);
nor U45229 (N_45229,N_31929,N_35199);
xor U45230 (N_45230,N_37052,N_36662);
nand U45231 (N_45231,N_39682,N_32283);
xnor U45232 (N_45232,N_37580,N_37438);
nand U45233 (N_45233,N_30292,N_34538);
or U45234 (N_45234,N_35081,N_32818);
or U45235 (N_45235,N_36257,N_33151);
nand U45236 (N_45236,N_32496,N_33917);
nand U45237 (N_45237,N_33176,N_38856);
or U45238 (N_45238,N_38407,N_32362);
or U45239 (N_45239,N_34052,N_36400);
nand U45240 (N_45240,N_38455,N_38296);
or U45241 (N_45241,N_31758,N_39062);
nor U45242 (N_45242,N_33919,N_31193);
xor U45243 (N_45243,N_30077,N_37617);
and U45244 (N_45244,N_31526,N_34873);
nor U45245 (N_45245,N_39217,N_30411);
nor U45246 (N_45246,N_31690,N_32296);
nand U45247 (N_45247,N_36759,N_37181);
xor U45248 (N_45248,N_30391,N_38666);
and U45249 (N_45249,N_39699,N_34117);
or U45250 (N_45250,N_35868,N_34696);
nor U45251 (N_45251,N_32852,N_30363);
or U45252 (N_45252,N_35654,N_30488);
nand U45253 (N_45253,N_39413,N_32262);
xnor U45254 (N_45254,N_38667,N_30755);
xnor U45255 (N_45255,N_37115,N_30534);
nand U45256 (N_45256,N_36954,N_38972);
or U45257 (N_45257,N_31080,N_33851);
and U45258 (N_45258,N_37663,N_33055);
and U45259 (N_45259,N_37337,N_33209);
nand U45260 (N_45260,N_35851,N_33796);
nand U45261 (N_45261,N_33537,N_33974);
nor U45262 (N_45262,N_32904,N_32663);
xnor U45263 (N_45263,N_31013,N_37821);
xor U45264 (N_45264,N_36696,N_35847);
or U45265 (N_45265,N_33743,N_34280);
nand U45266 (N_45266,N_38215,N_38468);
xor U45267 (N_45267,N_37350,N_31956);
and U45268 (N_45268,N_33339,N_37020);
or U45269 (N_45269,N_32473,N_32509);
and U45270 (N_45270,N_30747,N_35402);
or U45271 (N_45271,N_31337,N_32653);
xor U45272 (N_45272,N_31378,N_30272);
nand U45273 (N_45273,N_30629,N_38860);
or U45274 (N_45274,N_31623,N_35539);
or U45275 (N_45275,N_39535,N_36217);
or U45276 (N_45276,N_36320,N_39203);
or U45277 (N_45277,N_33450,N_33626);
xor U45278 (N_45278,N_37521,N_31880);
and U45279 (N_45279,N_35941,N_36405);
xnor U45280 (N_45280,N_30474,N_31906);
xor U45281 (N_45281,N_37859,N_34817);
nand U45282 (N_45282,N_34419,N_38738);
and U45283 (N_45283,N_37466,N_37148);
nand U45284 (N_45284,N_38744,N_35900);
or U45285 (N_45285,N_38172,N_35920);
xnor U45286 (N_45286,N_35211,N_30755);
xnor U45287 (N_45287,N_38772,N_39098);
xor U45288 (N_45288,N_33891,N_32435);
nor U45289 (N_45289,N_32107,N_37693);
and U45290 (N_45290,N_37074,N_36123);
xnor U45291 (N_45291,N_33395,N_39984);
or U45292 (N_45292,N_38082,N_39444);
nand U45293 (N_45293,N_31502,N_35231);
nor U45294 (N_45294,N_37432,N_39710);
nor U45295 (N_45295,N_34733,N_38164);
xnor U45296 (N_45296,N_35433,N_33098);
nand U45297 (N_45297,N_31503,N_33953);
and U45298 (N_45298,N_35702,N_33367);
nand U45299 (N_45299,N_34261,N_33146);
nand U45300 (N_45300,N_36537,N_31614);
or U45301 (N_45301,N_38770,N_36904);
xnor U45302 (N_45302,N_31458,N_33384);
and U45303 (N_45303,N_34022,N_30813);
nand U45304 (N_45304,N_30771,N_34705);
and U45305 (N_45305,N_38222,N_30043);
and U45306 (N_45306,N_32280,N_32307);
and U45307 (N_45307,N_32762,N_39189);
nor U45308 (N_45308,N_36702,N_32082);
or U45309 (N_45309,N_37467,N_32596);
xor U45310 (N_45310,N_31314,N_36710);
nand U45311 (N_45311,N_34495,N_37218);
xnor U45312 (N_45312,N_35839,N_36517);
xor U45313 (N_45313,N_34166,N_30932);
xor U45314 (N_45314,N_36004,N_37685);
xnor U45315 (N_45315,N_39125,N_30819);
nor U45316 (N_45316,N_30181,N_37485);
and U45317 (N_45317,N_31153,N_33542);
nor U45318 (N_45318,N_30271,N_39310);
nor U45319 (N_45319,N_30277,N_36518);
and U45320 (N_45320,N_38202,N_32241);
nor U45321 (N_45321,N_32305,N_38951);
and U45322 (N_45322,N_34226,N_38735);
or U45323 (N_45323,N_34316,N_32504);
and U45324 (N_45324,N_35570,N_31777);
nand U45325 (N_45325,N_37302,N_32754);
or U45326 (N_45326,N_35224,N_33255);
nand U45327 (N_45327,N_32417,N_38537);
nand U45328 (N_45328,N_38814,N_33228);
xor U45329 (N_45329,N_36051,N_32080);
and U45330 (N_45330,N_33382,N_37342);
nor U45331 (N_45331,N_38117,N_32963);
nor U45332 (N_45332,N_30636,N_38953);
or U45333 (N_45333,N_37067,N_31974);
xor U45334 (N_45334,N_35360,N_35976);
nor U45335 (N_45335,N_31452,N_32515);
xnor U45336 (N_45336,N_35708,N_35352);
and U45337 (N_45337,N_33658,N_31001);
nand U45338 (N_45338,N_37120,N_32662);
nand U45339 (N_45339,N_33904,N_31673);
or U45340 (N_45340,N_34076,N_31884);
nor U45341 (N_45341,N_30481,N_37438);
and U45342 (N_45342,N_39276,N_30335);
or U45343 (N_45343,N_33505,N_33903);
and U45344 (N_45344,N_34900,N_37664);
or U45345 (N_45345,N_39584,N_33374);
xnor U45346 (N_45346,N_36816,N_33542);
xor U45347 (N_45347,N_35872,N_35250);
and U45348 (N_45348,N_39426,N_36122);
or U45349 (N_45349,N_33700,N_31396);
xor U45350 (N_45350,N_33581,N_37578);
and U45351 (N_45351,N_34024,N_33565);
or U45352 (N_45352,N_32505,N_32263);
xnor U45353 (N_45353,N_30104,N_32838);
and U45354 (N_45354,N_35457,N_30534);
nor U45355 (N_45355,N_35722,N_32383);
nand U45356 (N_45356,N_35764,N_39904);
nor U45357 (N_45357,N_33015,N_39445);
and U45358 (N_45358,N_31880,N_38713);
xor U45359 (N_45359,N_32666,N_31078);
nor U45360 (N_45360,N_38912,N_38402);
xor U45361 (N_45361,N_38973,N_36342);
nor U45362 (N_45362,N_33095,N_38875);
nor U45363 (N_45363,N_38585,N_37616);
or U45364 (N_45364,N_36266,N_32602);
or U45365 (N_45365,N_35940,N_36668);
or U45366 (N_45366,N_35215,N_34381);
and U45367 (N_45367,N_35093,N_35241);
xnor U45368 (N_45368,N_31431,N_32413);
and U45369 (N_45369,N_36256,N_33791);
nand U45370 (N_45370,N_37601,N_38041);
xor U45371 (N_45371,N_31986,N_33490);
or U45372 (N_45372,N_30222,N_36288);
or U45373 (N_45373,N_32186,N_35751);
nand U45374 (N_45374,N_31836,N_38689);
nand U45375 (N_45375,N_35325,N_34015);
xor U45376 (N_45376,N_39323,N_36190);
and U45377 (N_45377,N_36217,N_31808);
xor U45378 (N_45378,N_33677,N_30248);
xor U45379 (N_45379,N_38323,N_33363);
or U45380 (N_45380,N_31175,N_36788);
xnor U45381 (N_45381,N_39247,N_39182);
nand U45382 (N_45382,N_32567,N_32830);
or U45383 (N_45383,N_35912,N_33389);
xor U45384 (N_45384,N_38822,N_33094);
and U45385 (N_45385,N_35651,N_30309);
or U45386 (N_45386,N_39519,N_34716);
or U45387 (N_45387,N_31915,N_36177);
and U45388 (N_45388,N_37847,N_32841);
nor U45389 (N_45389,N_38335,N_38862);
xnor U45390 (N_45390,N_39031,N_30845);
xor U45391 (N_45391,N_32450,N_32773);
nand U45392 (N_45392,N_39382,N_35300);
nand U45393 (N_45393,N_38715,N_38516);
nand U45394 (N_45394,N_35844,N_36911);
xor U45395 (N_45395,N_33005,N_37914);
or U45396 (N_45396,N_32331,N_32351);
xor U45397 (N_45397,N_37616,N_39411);
and U45398 (N_45398,N_33119,N_32239);
or U45399 (N_45399,N_32589,N_30607);
nand U45400 (N_45400,N_39280,N_37628);
xnor U45401 (N_45401,N_31827,N_32796);
and U45402 (N_45402,N_32173,N_37618);
or U45403 (N_45403,N_36221,N_33209);
nor U45404 (N_45404,N_38768,N_31209);
and U45405 (N_45405,N_36196,N_34568);
nand U45406 (N_45406,N_34356,N_33790);
or U45407 (N_45407,N_30399,N_31115);
nand U45408 (N_45408,N_30371,N_30824);
nand U45409 (N_45409,N_33353,N_32729);
xor U45410 (N_45410,N_39438,N_37833);
nand U45411 (N_45411,N_36407,N_32794);
xor U45412 (N_45412,N_38641,N_36679);
or U45413 (N_45413,N_36849,N_38532);
and U45414 (N_45414,N_37173,N_36950);
and U45415 (N_45415,N_32179,N_34810);
xor U45416 (N_45416,N_30617,N_30185);
or U45417 (N_45417,N_38817,N_34370);
nor U45418 (N_45418,N_35542,N_31369);
nor U45419 (N_45419,N_38783,N_38113);
and U45420 (N_45420,N_39301,N_38920);
and U45421 (N_45421,N_39613,N_38836);
xor U45422 (N_45422,N_31474,N_36959);
and U45423 (N_45423,N_35284,N_37525);
xor U45424 (N_45424,N_35553,N_38157);
xnor U45425 (N_45425,N_37924,N_38582);
nand U45426 (N_45426,N_31124,N_32142);
and U45427 (N_45427,N_35142,N_31588);
nand U45428 (N_45428,N_33786,N_39335);
or U45429 (N_45429,N_38019,N_32467);
xor U45430 (N_45430,N_30304,N_33912);
xor U45431 (N_45431,N_36163,N_38151);
nand U45432 (N_45432,N_30097,N_33529);
and U45433 (N_45433,N_37809,N_35324);
nor U45434 (N_45434,N_32240,N_38774);
nand U45435 (N_45435,N_34090,N_30951);
or U45436 (N_45436,N_36118,N_35222);
xor U45437 (N_45437,N_39145,N_30578);
nand U45438 (N_45438,N_38917,N_37495);
xor U45439 (N_45439,N_35707,N_39192);
nand U45440 (N_45440,N_31491,N_30295);
or U45441 (N_45441,N_31505,N_34390);
nand U45442 (N_45442,N_38282,N_33835);
nand U45443 (N_45443,N_37300,N_37188);
nand U45444 (N_45444,N_33431,N_32962);
and U45445 (N_45445,N_35845,N_36446);
or U45446 (N_45446,N_33506,N_30130);
nor U45447 (N_45447,N_39495,N_39106);
or U45448 (N_45448,N_38739,N_30504);
nand U45449 (N_45449,N_34180,N_35961);
nand U45450 (N_45450,N_30499,N_38349);
xor U45451 (N_45451,N_31800,N_35454);
nor U45452 (N_45452,N_34955,N_30230);
xnor U45453 (N_45453,N_31005,N_30563);
nor U45454 (N_45454,N_34830,N_38740);
nor U45455 (N_45455,N_31675,N_39471);
and U45456 (N_45456,N_31723,N_39600);
and U45457 (N_45457,N_38956,N_39033);
and U45458 (N_45458,N_30915,N_39301);
xnor U45459 (N_45459,N_34369,N_38810);
or U45460 (N_45460,N_38023,N_38226);
or U45461 (N_45461,N_36332,N_32962);
nand U45462 (N_45462,N_37852,N_31414);
or U45463 (N_45463,N_36311,N_34555);
or U45464 (N_45464,N_39883,N_36628);
nor U45465 (N_45465,N_34238,N_39668);
or U45466 (N_45466,N_36764,N_30660);
nor U45467 (N_45467,N_32532,N_38014);
xor U45468 (N_45468,N_34131,N_39243);
and U45469 (N_45469,N_33734,N_30564);
nand U45470 (N_45470,N_39835,N_30845);
xor U45471 (N_45471,N_39363,N_38120);
nor U45472 (N_45472,N_34456,N_38309);
nand U45473 (N_45473,N_36084,N_32765);
or U45474 (N_45474,N_36354,N_38688);
nor U45475 (N_45475,N_32771,N_34529);
nor U45476 (N_45476,N_36182,N_30831);
and U45477 (N_45477,N_35316,N_37866);
or U45478 (N_45478,N_38847,N_32761);
nand U45479 (N_45479,N_33713,N_37285);
or U45480 (N_45480,N_32748,N_30607);
or U45481 (N_45481,N_35767,N_37149);
or U45482 (N_45482,N_33228,N_35984);
nor U45483 (N_45483,N_31364,N_36753);
nor U45484 (N_45484,N_37139,N_32390);
nor U45485 (N_45485,N_30301,N_32036);
xor U45486 (N_45486,N_31251,N_35848);
xor U45487 (N_45487,N_31585,N_31450);
nor U45488 (N_45488,N_30070,N_30971);
nand U45489 (N_45489,N_34343,N_31127);
nand U45490 (N_45490,N_37139,N_38470);
nor U45491 (N_45491,N_32400,N_37686);
and U45492 (N_45492,N_33299,N_32162);
or U45493 (N_45493,N_30099,N_37327);
and U45494 (N_45494,N_36962,N_32709);
nor U45495 (N_45495,N_32790,N_33921);
or U45496 (N_45496,N_33306,N_33726);
nand U45497 (N_45497,N_38208,N_33570);
nand U45498 (N_45498,N_36884,N_30826);
or U45499 (N_45499,N_31423,N_32815);
or U45500 (N_45500,N_37722,N_36759);
nor U45501 (N_45501,N_31903,N_34196);
or U45502 (N_45502,N_38667,N_32463);
and U45503 (N_45503,N_31357,N_32120);
and U45504 (N_45504,N_35927,N_38992);
and U45505 (N_45505,N_35116,N_30404);
nand U45506 (N_45506,N_36821,N_38122);
nor U45507 (N_45507,N_36350,N_33419);
and U45508 (N_45508,N_31318,N_32909);
nor U45509 (N_45509,N_31344,N_30093);
nand U45510 (N_45510,N_38461,N_35633);
and U45511 (N_45511,N_31373,N_36815);
nand U45512 (N_45512,N_31298,N_39381);
nand U45513 (N_45513,N_36865,N_30117);
or U45514 (N_45514,N_39407,N_35396);
nor U45515 (N_45515,N_34443,N_30834);
nor U45516 (N_45516,N_35711,N_35868);
nand U45517 (N_45517,N_39439,N_39818);
and U45518 (N_45518,N_35377,N_33624);
nand U45519 (N_45519,N_39642,N_31210);
and U45520 (N_45520,N_35396,N_33841);
nand U45521 (N_45521,N_31809,N_30594);
nor U45522 (N_45522,N_38042,N_30056);
xnor U45523 (N_45523,N_38786,N_31381);
nand U45524 (N_45524,N_37596,N_30286);
nand U45525 (N_45525,N_37019,N_34670);
or U45526 (N_45526,N_33098,N_36978);
nor U45527 (N_45527,N_39976,N_35596);
nor U45528 (N_45528,N_33132,N_30467);
and U45529 (N_45529,N_32912,N_37832);
xnor U45530 (N_45530,N_39707,N_37735);
nand U45531 (N_45531,N_38571,N_39355);
nor U45532 (N_45532,N_37127,N_34932);
nand U45533 (N_45533,N_38815,N_38343);
nand U45534 (N_45534,N_38977,N_31367);
nor U45535 (N_45535,N_34598,N_36516);
nand U45536 (N_45536,N_39302,N_36224);
nor U45537 (N_45537,N_36020,N_36452);
and U45538 (N_45538,N_39261,N_37331);
nand U45539 (N_45539,N_30447,N_32842);
or U45540 (N_45540,N_36128,N_31574);
or U45541 (N_45541,N_32980,N_34737);
and U45542 (N_45542,N_35077,N_39816);
and U45543 (N_45543,N_38805,N_36250);
and U45544 (N_45544,N_35014,N_36332);
nand U45545 (N_45545,N_39083,N_33952);
nand U45546 (N_45546,N_35909,N_33540);
or U45547 (N_45547,N_33093,N_30706);
nand U45548 (N_45548,N_36115,N_37898);
and U45549 (N_45549,N_37616,N_34970);
nand U45550 (N_45550,N_39300,N_38445);
nor U45551 (N_45551,N_34904,N_39503);
nor U45552 (N_45552,N_31778,N_34614);
or U45553 (N_45553,N_38727,N_34163);
xnor U45554 (N_45554,N_33193,N_37129);
nor U45555 (N_45555,N_38413,N_31586);
nor U45556 (N_45556,N_34306,N_39385);
and U45557 (N_45557,N_33657,N_33282);
nor U45558 (N_45558,N_34250,N_31730);
xnor U45559 (N_45559,N_33003,N_34118);
or U45560 (N_45560,N_30834,N_36260);
and U45561 (N_45561,N_37657,N_33470);
nand U45562 (N_45562,N_32145,N_38875);
or U45563 (N_45563,N_39265,N_34688);
xor U45564 (N_45564,N_32971,N_36278);
or U45565 (N_45565,N_31101,N_38857);
xnor U45566 (N_45566,N_37041,N_33801);
and U45567 (N_45567,N_36429,N_34439);
nor U45568 (N_45568,N_39256,N_31827);
nor U45569 (N_45569,N_39409,N_37188);
or U45570 (N_45570,N_31554,N_33227);
xor U45571 (N_45571,N_35744,N_39106);
nand U45572 (N_45572,N_33248,N_32869);
xnor U45573 (N_45573,N_39791,N_30803);
nor U45574 (N_45574,N_34135,N_31597);
xor U45575 (N_45575,N_35215,N_30914);
or U45576 (N_45576,N_30829,N_38959);
nand U45577 (N_45577,N_38329,N_30948);
or U45578 (N_45578,N_35689,N_36162);
nand U45579 (N_45579,N_31696,N_34671);
or U45580 (N_45580,N_39078,N_37820);
nand U45581 (N_45581,N_35863,N_33309);
and U45582 (N_45582,N_32288,N_39323);
nor U45583 (N_45583,N_33398,N_36954);
nor U45584 (N_45584,N_32745,N_33635);
xnor U45585 (N_45585,N_38971,N_38848);
or U45586 (N_45586,N_37378,N_33109);
xnor U45587 (N_45587,N_32411,N_32275);
xnor U45588 (N_45588,N_39562,N_35558);
or U45589 (N_45589,N_38232,N_37665);
xnor U45590 (N_45590,N_39898,N_33340);
and U45591 (N_45591,N_37173,N_35600);
xnor U45592 (N_45592,N_38701,N_31415);
xor U45593 (N_45593,N_32482,N_37830);
nor U45594 (N_45594,N_34384,N_39122);
nand U45595 (N_45595,N_30295,N_37434);
nand U45596 (N_45596,N_36520,N_35503);
xnor U45597 (N_45597,N_39225,N_36228);
and U45598 (N_45598,N_38811,N_33470);
nand U45599 (N_45599,N_35588,N_32397);
xnor U45600 (N_45600,N_32661,N_30091);
and U45601 (N_45601,N_39028,N_31002);
nand U45602 (N_45602,N_37314,N_39940);
or U45603 (N_45603,N_35542,N_32050);
and U45604 (N_45604,N_32727,N_37969);
xor U45605 (N_45605,N_37633,N_33114);
nor U45606 (N_45606,N_31722,N_35959);
nor U45607 (N_45607,N_34538,N_30475);
nand U45608 (N_45608,N_39056,N_32243);
xor U45609 (N_45609,N_31434,N_37095);
nand U45610 (N_45610,N_31355,N_30562);
or U45611 (N_45611,N_38117,N_33728);
nor U45612 (N_45612,N_32757,N_39525);
xor U45613 (N_45613,N_35936,N_38034);
nor U45614 (N_45614,N_34204,N_35846);
nor U45615 (N_45615,N_32418,N_32955);
or U45616 (N_45616,N_30698,N_39229);
nor U45617 (N_45617,N_37633,N_31673);
xor U45618 (N_45618,N_31977,N_36400);
nor U45619 (N_45619,N_39073,N_32564);
and U45620 (N_45620,N_32631,N_32574);
xor U45621 (N_45621,N_37815,N_30105);
or U45622 (N_45622,N_36414,N_37329);
or U45623 (N_45623,N_34868,N_34770);
or U45624 (N_45624,N_33006,N_32227);
nor U45625 (N_45625,N_34045,N_39062);
and U45626 (N_45626,N_39125,N_35251);
or U45627 (N_45627,N_38684,N_33856);
xnor U45628 (N_45628,N_32140,N_34458);
and U45629 (N_45629,N_33392,N_35461);
nand U45630 (N_45630,N_33748,N_32947);
nand U45631 (N_45631,N_35017,N_38453);
nand U45632 (N_45632,N_30275,N_32637);
or U45633 (N_45633,N_38215,N_37421);
or U45634 (N_45634,N_37291,N_33899);
nor U45635 (N_45635,N_33108,N_34766);
or U45636 (N_45636,N_33703,N_30414);
and U45637 (N_45637,N_38473,N_38047);
nor U45638 (N_45638,N_32428,N_33548);
or U45639 (N_45639,N_34258,N_35261);
or U45640 (N_45640,N_37705,N_39122);
nor U45641 (N_45641,N_31455,N_33910);
and U45642 (N_45642,N_33373,N_36783);
nor U45643 (N_45643,N_39284,N_32797);
nor U45644 (N_45644,N_38019,N_39200);
xnor U45645 (N_45645,N_34785,N_37092);
nor U45646 (N_45646,N_34795,N_39106);
xor U45647 (N_45647,N_34303,N_37955);
and U45648 (N_45648,N_30321,N_30170);
xnor U45649 (N_45649,N_37703,N_38795);
nand U45650 (N_45650,N_31735,N_36690);
xnor U45651 (N_45651,N_34477,N_35927);
or U45652 (N_45652,N_34746,N_39148);
nand U45653 (N_45653,N_37254,N_32991);
and U45654 (N_45654,N_34244,N_38197);
xnor U45655 (N_45655,N_34939,N_39458);
xor U45656 (N_45656,N_35054,N_30391);
or U45657 (N_45657,N_39216,N_39226);
xor U45658 (N_45658,N_32689,N_30401);
xor U45659 (N_45659,N_39030,N_37571);
xor U45660 (N_45660,N_33721,N_30271);
and U45661 (N_45661,N_36451,N_33218);
and U45662 (N_45662,N_34119,N_35432);
or U45663 (N_45663,N_35358,N_32905);
xor U45664 (N_45664,N_37994,N_30024);
or U45665 (N_45665,N_31983,N_33865);
nor U45666 (N_45666,N_32234,N_32495);
or U45667 (N_45667,N_33154,N_32287);
nand U45668 (N_45668,N_30333,N_33950);
nor U45669 (N_45669,N_30501,N_33703);
xor U45670 (N_45670,N_38976,N_32282);
or U45671 (N_45671,N_33175,N_38509);
nor U45672 (N_45672,N_34702,N_36466);
or U45673 (N_45673,N_33113,N_39308);
nand U45674 (N_45674,N_37651,N_39679);
xnor U45675 (N_45675,N_34124,N_38807);
or U45676 (N_45676,N_34597,N_36751);
xor U45677 (N_45677,N_36131,N_31396);
nand U45678 (N_45678,N_36761,N_31057);
or U45679 (N_45679,N_33238,N_35774);
and U45680 (N_45680,N_38927,N_35448);
and U45681 (N_45681,N_31587,N_33332);
or U45682 (N_45682,N_33483,N_32678);
nand U45683 (N_45683,N_34961,N_35055);
xnor U45684 (N_45684,N_31789,N_30603);
xnor U45685 (N_45685,N_31396,N_34432);
nor U45686 (N_45686,N_32255,N_38517);
nand U45687 (N_45687,N_37076,N_38843);
and U45688 (N_45688,N_32838,N_36291);
or U45689 (N_45689,N_32226,N_39351);
xor U45690 (N_45690,N_37586,N_34475);
nor U45691 (N_45691,N_32892,N_36970);
or U45692 (N_45692,N_34184,N_33505);
nand U45693 (N_45693,N_30424,N_33205);
nor U45694 (N_45694,N_30793,N_34379);
nor U45695 (N_45695,N_37251,N_34855);
xor U45696 (N_45696,N_37049,N_37865);
nor U45697 (N_45697,N_36789,N_31518);
xor U45698 (N_45698,N_39177,N_34051);
xor U45699 (N_45699,N_30515,N_32472);
nor U45700 (N_45700,N_37750,N_35689);
or U45701 (N_45701,N_35404,N_35164);
or U45702 (N_45702,N_36124,N_37144);
xnor U45703 (N_45703,N_30090,N_30133);
and U45704 (N_45704,N_36756,N_31397);
or U45705 (N_45705,N_39539,N_35092);
nor U45706 (N_45706,N_31924,N_36772);
or U45707 (N_45707,N_30623,N_38027);
nand U45708 (N_45708,N_35210,N_39879);
and U45709 (N_45709,N_33481,N_33602);
or U45710 (N_45710,N_37303,N_36257);
and U45711 (N_45711,N_36623,N_34987);
nand U45712 (N_45712,N_39202,N_34212);
or U45713 (N_45713,N_33348,N_32514);
xnor U45714 (N_45714,N_34806,N_35004);
or U45715 (N_45715,N_30165,N_34370);
and U45716 (N_45716,N_32210,N_36197);
nand U45717 (N_45717,N_33929,N_33219);
or U45718 (N_45718,N_37734,N_36863);
nand U45719 (N_45719,N_32681,N_30477);
and U45720 (N_45720,N_35700,N_38756);
or U45721 (N_45721,N_32747,N_37641);
xnor U45722 (N_45722,N_32630,N_38238);
xor U45723 (N_45723,N_34866,N_39781);
nor U45724 (N_45724,N_36760,N_39616);
xnor U45725 (N_45725,N_36580,N_30133);
or U45726 (N_45726,N_30589,N_34106);
and U45727 (N_45727,N_39989,N_35774);
or U45728 (N_45728,N_33075,N_32002);
or U45729 (N_45729,N_35768,N_32362);
or U45730 (N_45730,N_37033,N_37438);
nand U45731 (N_45731,N_33651,N_37634);
and U45732 (N_45732,N_35385,N_35752);
and U45733 (N_45733,N_31758,N_36023);
or U45734 (N_45734,N_31867,N_37241);
nor U45735 (N_45735,N_35863,N_31861);
or U45736 (N_45736,N_38812,N_30832);
or U45737 (N_45737,N_35773,N_36000);
xnor U45738 (N_45738,N_32303,N_31314);
and U45739 (N_45739,N_31446,N_30661);
and U45740 (N_45740,N_37257,N_34277);
or U45741 (N_45741,N_37912,N_39755);
nand U45742 (N_45742,N_39462,N_37413);
nor U45743 (N_45743,N_32556,N_39043);
or U45744 (N_45744,N_38356,N_30790);
xor U45745 (N_45745,N_38265,N_38939);
or U45746 (N_45746,N_30454,N_39788);
nor U45747 (N_45747,N_37061,N_30810);
and U45748 (N_45748,N_38851,N_32800);
and U45749 (N_45749,N_30154,N_32294);
xnor U45750 (N_45750,N_37480,N_30942);
or U45751 (N_45751,N_30561,N_31313);
nand U45752 (N_45752,N_37420,N_38695);
nor U45753 (N_45753,N_38529,N_37244);
nor U45754 (N_45754,N_35427,N_39413);
nor U45755 (N_45755,N_30304,N_33850);
or U45756 (N_45756,N_30503,N_33392);
and U45757 (N_45757,N_39015,N_37392);
nand U45758 (N_45758,N_36193,N_39493);
and U45759 (N_45759,N_33965,N_37305);
and U45760 (N_45760,N_32980,N_31863);
nor U45761 (N_45761,N_33560,N_39768);
nand U45762 (N_45762,N_37533,N_37343);
xor U45763 (N_45763,N_30463,N_35997);
or U45764 (N_45764,N_30227,N_35353);
nor U45765 (N_45765,N_31061,N_31765);
nand U45766 (N_45766,N_31043,N_30882);
nor U45767 (N_45767,N_33737,N_38364);
or U45768 (N_45768,N_34696,N_30271);
or U45769 (N_45769,N_30952,N_32773);
and U45770 (N_45770,N_37487,N_30310);
and U45771 (N_45771,N_32639,N_38938);
nand U45772 (N_45772,N_31104,N_34574);
or U45773 (N_45773,N_39299,N_34791);
nor U45774 (N_45774,N_32653,N_39526);
nand U45775 (N_45775,N_39068,N_39728);
and U45776 (N_45776,N_36744,N_34832);
nand U45777 (N_45777,N_38178,N_34591);
and U45778 (N_45778,N_33614,N_33976);
nand U45779 (N_45779,N_36065,N_39215);
and U45780 (N_45780,N_36905,N_36884);
nor U45781 (N_45781,N_34118,N_33405);
xor U45782 (N_45782,N_35560,N_31522);
xor U45783 (N_45783,N_31691,N_35169);
or U45784 (N_45784,N_30454,N_36082);
or U45785 (N_45785,N_33465,N_35646);
and U45786 (N_45786,N_34386,N_33350);
nand U45787 (N_45787,N_38700,N_39303);
xnor U45788 (N_45788,N_38503,N_34025);
xor U45789 (N_45789,N_32094,N_30574);
xor U45790 (N_45790,N_36570,N_36106);
xor U45791 (N_45791,N_32167,N_38877);
or U45792 (N_45792,N_30473,N_31825);
nor U45793 (N_45793,N_35205,N_34406);
nand U45794 (N_45794,N_30045,N_39720);
nor U45795 (N_45795,N_36832,N_33641);
xor U45796 (N_45796,N_32154,N_35281);
nor U45797 (N_45797,N_36980,N_34278);
xnor U45798 (N_45798,N_31288,N_31825);
nand U45799 (N_45799,N_35133,N_36219);
xnor U45800 (N_45800,N_30111,N_36492);
and U45801 (N_45801,N_36219,N_37183);
and U45802 (N_45802,N_34822,N_32425);
nand U45803 (N_45803,N_36627,N_35209);
and U45804 (N_45804,N_31653,N_38295);
nor U45805 (N_45805,N_34220,N_34505);
xnor U45806 (N_45806,N_30555,N_30659);
and U45807 (N_45807,N_39394,N_39507);
or U45808 (N_45808,N_34190,N_39458);
nor U45809 (N_45809,N_35977,N_34817);
and U45810 (N_45810,N_30659,N_30460);
or U45811 (N_45811,N_31938,N_33421);
or U45812 (N_45812,N_35517,N_39341);
or U45813 (N_45813,N_32062,N_38176);
xor U45814 (N_45814,N_38920,N_31286);
nand U45815 (N_45815,N_30226,N_33366);
nor U45816 (N_45816,N_39913,N_36428);
nor U45817 (N_45817,N_37455,N_33746);
xor U45818 (N_45818,N_32529,N_32962);
nand U45819 (N_45819,N_32029,N_36662);
or U45820 (N_45820,N_31908,N_32461);
and U45821 (N_45821,N_36261,N_34010);
and U45822 (N_45822,N_36950,N_38666);
nor U45823 (N_45823,N_34932,N_38687);
nor U45824 (N_45824,N_30607,N_31345);
or U45825 (N_45825,N_32126,N_36769);
or U45826 (N_45826,N_31471,N_30354);
or U45827 (N_45827,N_39441,N_35591);
nor U45828 (N_45828,N_31956,N_36984);
or U45829 (N_45829,N_39860,N_36722);
xor U45830 (N_45830,N_34308,N_31412);
or U45831 (N_45831,N_37958,N_38799);
or U45832 (N_45832,N_30800,N_33783);
or U45833 (N_45833,N_31416,N_38600);
nand U45834 (N_45834,N_36640,N_32922);
and U45835 (N_45835,N_37866,N_33879);
and U45836 (N_45836,N_38484,N_37620);
nor U45837 (N_45837,N_31353,N_37966);
xor U45838 (N_45838,N_32403,N_33285);
nor U45839 (N_45839,N_35778,N_34682);
or U45840 (N_45840,N_32264,N_39823);
nand U45841 (N_45841,N_39133,N_32915);
nand U45842 (N_45842,N_34975,N_32390);
xor U45843 (N_45843,N_35047,N_39008);
nor U45844 (N_45844,N_33523,N_35053);
nor U45845 (N_45845,N_38048,N_38614);
nor U45846 (N_45846,N_36967,N_39296);
xnor U45847 (N_45847,N_37665,N_39197);
nand U45848 (N_45848,N_30413,N_33855);
and U45849 (N_45849,N_30107,N_37411);
or U45850 (N_45850,N_39901,N_32760);
and U45851 (N_45851,N_35526,N_38791);
or U45852 (N_45852,N_36125,N_32155);
xnor U45853 (N_45853,N_38213,N_34137);
nand U45854 (N_45854,N_39259,N_36618);
or U45855 (N_45855,N_38585,N_33425);
xnor U45856 (N_45856,N_32407,N_32656);
or U45857 (N_45857,N_39829,N_30358);
nand U45858 (N_45858,N_30272,N_36671);
nor U45859 (N_45859,N_37280,N_33876);
xor U45860 (N_45860,N_30045,N_36663);
nand U45861 (N_45861,N_36605,N_35763);
xnor U45862 (N_45862,N_39402,N_30132);
xnor U45863 (N_45863,N_39496,N_38340);
xnor U45864 (N_45864,N_33336,N_36219);
nor U45865 (N_45865,N_37581,N_33293);
nor U45866 (N_45866,N_38988,N_38785);
nand U45867 (N_45867,N_34446,N_37863);
or U45868 (N_45868,N_39309,N_33419);
or U45869 (N_45869,N_31291,N_34464);
or U45870 (N_45870,N_39400,N_35365);
nand U45871 (N_45871,N_37534,N_31337);
xor U45872 (N_45872,N_38869,N_37056);
nor U45873 (N_45873,N_39982,N_30899);
xor U45874 (N_45874,N_30095,N_38257);
xor U45875 (N_45875,N_36253,N_37123);
and U45876 (N_45876,N_31035,N_36510);
or U45877 (N_45877,N_37764,N_39158);
nand U45878 (N_45878,N_34877,N_34794);
or U45879 (N_45879,N_36133,N_37131);
xor U45880 (N_45880,N_39463,N_30738);
xnor U45881 (N_45881,N_38852,N_31833);
or U45882 (N_45882,N_31429,N_38918);
nand U45883 (N_45883,N_35306,N_37618);
and U45884 (N_45884,N_36750,N_34907);
nand U45885 (N_45885,N_38163,N_39620);
or U45886 (N_45886,N_35951,N_35872);
xor U45887 (N_45887,N_32514,N_37815);
nand U45888 (N_45888,N_32047,N_39578);
nand U45889 (N_45889,N_30322,N_31498);
and U45890 (N_45890,N_38135,N_31121);
xor U45891 (N_45891,N_32611,N_34444);
and U45892 (N_45892,N_33626,N_34864);
nor U45893 (N_45893,N_36025,N_35957);
nand U45894 (N_45894,N_30778,N_39141);
and U45895 (N_45895,N_30566,N_38413);
xor U45896 (N_45896,N_37581,N_38125);
or U45897 (N_45897,N_31020,N_36948);
nor U45898 (N_45898,N_31431,N_30902);
xnor U45899 (N_45899,N_34952,N_34550);
xnor U45900 (N_45900,N_33621,N_36142);
and U45901 (N_45901,N_36797,N_32141);
nor U45902 (N_45902,N_31649,N_35304);
nand U45903 (N_45903,N_39212,N_34610);
xor U45904 (N_45904,N_36400,N_36318);
nor U45905 (N_45905,N_37469,N_36980);
xnor U45906 (N_45906,N_34030,N_38615);
or U45907 (N_45907,N_36597,N_30814);
and U45908 (N_45908,N_33423,N_36964);
xnor U45909 (N_45909,N_36255,N_32787);
and U45910 (N_45910,N_36569,N_30116);
nand U45911 (N_45911,N_34458,N_33692);
or U45912 (N_45912,N_31318,N_37350);
and U45913 (N_45913,N_30468,N_36775);
and U45914 (N_45914,N_36372,N_38738);
nor U45915 (N_45915,N_31291,N_39674);
nand U45916 (N_45916,N_32764,N_34549);
nor U45917 (N_45917,N_32034,N_38716);
or U45918 (N_45918,N_39417,N_32516);
and U45919 (N_45919,N_37621,N_38280);
nand U45920 (N_45920,N_31932,N_39924);
or U45921 (N_45921,N_38492,N_30216);
and U45922 (N_45922,N_35272,N_33486);
nand U45923 (N_45923,N_38882,N_36116);
nor U45924 (N_45924,N_32051,N_31193);
nor U45925 (N_45925,N_31725,N_30671);
or U45926 (N_45926,N_37902,N_39751);
nor U45927 (N_45927,N_34484,N_33726);
or U45928 (N_45928,N_35176,N_35458);
nand U45929 (N_45929,N_39004,N_30723);
xnor U45930 (N_45930,N_37209,N_38962);
nor U45931 (N_45931,N_39403,N_33779);
xor U45932 (N_45932,N_33617,N_38527);
or U45933 (N_45933,N_35198,N_38480);
and U45934 (N_45934,N_35724,N_34599);
xnor U45935 (N_45935,N_35755,N_36088);
nor U45936 (N_45936,N_37354,N_38261);
or U45937 (N_45937,N_34143,N_31198);
and U45938 (N_45938,N_37155,N_30437);
or U45939 (N_45939,N_31431,N_37940);
nand U45940 (N_45940,N_33407,N_33521);
and U45941 (N_45941,N_33648,N_33383);
xor U45942 (N_45942,N_32695,N_39409);
nor U45943 (N_45943,N_35040,N_36410);
and U45944 (N_45944,N_38355,N_33234);
nand U45945 (N_45945,N_36119,N_31146);
xor U45946 (N_45946,N_30054,N_33534);
nor U45947 (N_45947,N_39208,N_38271);
or U45948 (N_45948,N_30040,N_32237);
and U45949 (N_45949,N_37814,N_34422);
nor U45950 (N_45950,N_33590,N_30648);
xnor U45951 (N_45951,N_37273,N_39194);
nand U45952 (N_45952,N_39168,N_35091);
and U45953 (N_45953,N_37088,N_39172);
and U45954 (N_45954,N_35301,N_36711);
nand U45955 (N_45955,N_37926,N_38475);
and U45956 (N_45956,N_38963,N_37313);
and U45957 (N_45957,N_30635,N_39422);
nand U45958 (N_45958,N_31323,N_33465);
xnor U45959 (N_45959,N_32131,N_36877);
and U45960 (N_45960,N_34454,N_35043);
nand U45961 (N_45961,N_38426,N_37853);
or U45962 (N_45962,N_33266,N_37247);
nand U45963 (N_45963,N_37221,N_35628);
nor U45964 (N_45964,N_30823,N_33642);
xnor U45965 (N_45965,N_38967,N_32507);
and U45966 (N_45966,N_39374,N_32399);
xnor U45967 (N_45967,N_31067,N_37054);
or U45968 (N_45968,N_37404,N_36993);
xnor U45969 (N_45969,N_35694,N_30507);
nand U45970 (N_45970,N_31925,N_31609);
or U45971 (N_45971,N_38247,N_33933);
xor U45972 (N_45972,N_39933,N_38996);
and U45973 (N_45973,N_30726,N_38221);
or U45974 (N_45974,N_34261,N_38884);
nor U45975 (N_45975,N_33099,N_33462);
nor U45976 (N_45976,N_31024,N_32293);
nand U45977 (N_45977,N_33246,N_32713);
xnor U45978 (N_45978,N_33254,N_35145);
or U45979 (N_45979,N_37576,N_39495);
or U45980 (N_45980,N_32325,N_37922);
nor U45981 (N_45981,N_33447,N_38634);
or U45982 (N_45982,N_32452,N_39704);
nor U45983 (N_45983,N_35216,N_34637);
xnor U45984 (N_45984,N_38576,N_39369);
and U45985 (N_45985,N_33789,N_35263);
or U45986 (N_45986,N_33256,N_39390);
nor U45987 (N_45987,N_33904,N_39252);
nand U45988 (N_45988,N_39732,N_36064);
nor U45989 (N_45989,N_37309,N_30020);
nand U45990 (N_45990,N_30719,N_33557);
nand U45991 (N_45991,N_38937,N_31079);
nand U45992 (N_45992,N_31098,N_30200);
nand U45993 (N_45993,N_34332,N_38429);
nand U45994 (N_45994,N_38160,N_31131);
nand U45995 (N_45995,N_37175,N_38695);
nor U45996 (N_45996,N_32863,N_34250);
xor U45997 (N_45997,N_36269,N_34163);
xor U45998 (N_45998,N_33495,N_34005);
or U45999 (N_45999,N_32097,N_34887);
xnor U46000 (N_46000,N_30565,N_37706);
nand U46001 (N_46001,N_31420,N_35689);
or U46002 (N_46002,N_38650,N_31734);
nand U46003 (N_46003,N_35718,N_32068);
nand U46004 (N_46004,N_31639,N_36302);
nand U46005 (N_46005,N_30364,N_33799);
xor U46006 (N_46006,N_30564,N_37424);
nand U46007 (N_46007,N_38547,N_37607);
xnor U46008 (N_46008,N_38144,N_36553);
nand U46009 (N_46009,N_33987,N_32082);
and U46010 (N_46010,N_36882,N_33017);
nor U46011 (N_46011,N_38618,N_39828);
and U46012 (N_46012,N_37645,N_33540);
nand U46013 (N_46013,N_30180,N_31437);
or U46014 (N_46014,N_34240,N_37005);
xnor U46015 (N_46015,N_30459,N_34786);
xnor U46016 (N_46016,N_34623,N_37504);
or U46017 (N_46017,N_34020,N_30738);
nand U46018 (N_46018,N_31263,N_33823);
or U46019 (N_46019,N_39501,N_36798);
and U46020 (N_46020,N_38342,N_36709);
or U46021 (N_46021,N_34524,N_37345);
and U46022 (N_46022,N_37098,N_30857);
or U46023 (N_46023,N_35200,N_38140);
xnor U46024 (N_46024,N_37549,N_33896);
nand U46025 (N_46025,N_30822,N_36020);
or U46026 (N_46026,N_34273,N_36049);
or U46027 (N_46027,N_33541,N_38614);
and U46028 (N_46028,N_33771,N_36446);
nor U46029 (N_46029,N_34358,N_36407);
nand U46030 (N_46030,N_36451,N_31011);
and U46031 (N_46031,N_33777,N_32310);
nor U46032 (N_46032,N_30842,N_33091);
xnor U46033 (N_46033,N_38774,N_35440);
and U46034 (N_46034,N_30401,N_31611);
xor U46035 (N_46035,N_38526,N_31250);
or U46036 (N_46036,N_30034,N_30027);
or U46037 (N_46037,N_32568,N_30539);
nand U46038 (N_46038,N_33320,N_34245);
or U46039 (N_46039,N_33836,N_35701);
nor U46040 (N_46040,N_34075,N_38887);
xnor U46041 (N_46041,N_37493,N_36932);
xor U46042 (N_46042,N_30464,N_30403);
xor U46043 (N_46043,N_34552,N_32831);
nand U46044 (N_46044,N_34082,N_39369);
nor U46045 (N_46045,N_34169,N_30337);
xor U46046 (N_46046,N_38272,N_33827);
and U46047 (N_46047,N_33967,N_39927);
nor U46048 (N_46048,N_39480,N_39398);
xnor U46049 (N_46049,N_39408,N_36757);
nand U46050 (N_46050,N_34662,N_30602);
nand U46051 (N_46051,N_37185,N_38499);
or U46052 (N_46052,N_39781,N_31814);
or U46053 (N_46053,N_39276,N_31873);
or U46054 (N_46054,N_33044,N_39472);
nand U46055 (N_46055,N_36712,N_34364);
or U46056 (N_46056,N_36274,N_38150);
nand U46057 (N_46057,N_35275,N_33050);
or U46058 (N_46058,N_37383,N_33485);
xnor U46059 (N_46059,N_37254,N_36977);
nand U46060 (N_46060,N_39340,N_32521);
nor U46061 (N_46061,N_37891,N_33376);
nand U46062 (N_46062,N_36399,N_34702);
nand U46063 (N_46063,N_30678,N_33799);
nor U46064 (N_46064,N_33657,N_37279);
xor U46065 (N_46065,N_31038,N_33969);
nor U46066 (N_46066,N_32510,N_38920);
nand U46067 (N_46067,N_35392,N_35353);
and U46068 (N_46068,N_30549,N_31270);
and U46069 (N_46069,N_34836,N_39826);
nor U46070 (N_46070,N_37020,N_34599);
nor U46071 (N_46071,N_36421,N_32750);
and U46072 (N_46072,N_39447,N_36284);
nor U46073 (N_46073,N_36590,N_33755);
or U46074 (N_46074,N_33689,N_33362);
nor U46075 (N_46075,N_30450,N_30704);
and U46076 (N_46076,N_36208,N_32903);
nor U46077 (N_46077,N_35190,N_37738);
nand U46078 (N_46078,N_31912,N_34340);
xnor U46079 (N_46079,N_32352,N_30068);
or U46080 (N_46080,N_36064,N_34270);
nand U46081 (N_46081,N_34558,N_34291);
nor U46082 (N_46082,N_30802,N_30566);
nor U46083 (N_46083,N_30415,N_38607);
and U46084 (N_46084,N_30061,N_32217);
nand U46085 (N_46085,N_33666,N_38373);
and U46086 (N_46086,N_34111,N_37469);
or U46087 (N_46087,N_38344,N_32892);
and U46088 (N_46088,N_31689,N_32729);
nor U46089 (N_46089,N_33159,N_34188);
nor U46090 (N_46090,N_30134,N_30602);
xor U46091 (N_46091,N_33219,N_32903);
or U46092 (N_46092,N_37753,N_36682);
and U46093 (N_46093,N_37383,N_32768);
xnor U46094 (N_46094,N_36939,N_37249);
nor U46095 (N_46095,N_33698,N_38613);
nand U46096 (N_46096,N_31336,N_38760);
xnor U46097 (N_46097,N_34170,N_34978);
xor U46098 (N_46098,N_38739,N_31514);
or U46099 (N_46099,N_32469,N_38643);
nand U46100 (N_46100,N_37301,N_33400);
nand U46101 (N_46101,N_37510,N_36791);
nor U46102 (N_46102,N_37393,N_33231);
and U46103 (N_46103,N_39578,N_39590);
nor U46104 (N_46104,N_33530,N_33151);
and U46105 (N_46105,N_36648,N_38862);
nor U46106 (N_46106,N_38836,N_31203);
nor U46107 (N_46107,N_35894,N_35406);
nor U46108 (N_46108,N_33060,N_32494);
or U46109 (N_46109,N_31277,N_33356);
or U46110 (N_46110,N_37014,N_33663);
nor U46111 (N_46111,N_34610,N_39458);
nand U46112 (N_46112,N_33584,N_36831);
and U46113 (N_46113,N_33211,N_39781);
xor U46114 (N_46114,N_39433,N_30443);
and U46115 (N_46115,N_38165,N_38911);
and U46116 (N_46116,N_37166,N_38633);
or U46117 (N_46117,N_32395,N_38572);
or U46118 (N_46118,N_36474,N_39758);
nand U46119 (N_46119,N_38711,N_34312);
nand U46120 (N_46120,N_39802,N_32651);
and U46121 (N_46121,N_30979,N_33420);
or U46122 (N_46122,N_37850,N_34015);
xor U46123 (N_46123,N_33738,N_34885);
nand U46124 (N_46124,N_30237,N_35148);
xor U46125 (N_46125,N_34983,N_33591);
nor U46126 (N_46126,N_36959,N_36360);
and U46127 (N_46127,N_30933,N_31378);
or U46128 (N_46128,N_30324,N_35728);
or U46129 (N_46129,N_33240,N_35420);
and U46130 (N_46130,N_38899,N_35460);
or U46131 (N_46131,N_39942,N_32038);
nand U46132 (N_46132,N_38697,N_33459);
nor U46133 (N_46133,N_38719,N_37759);
nor U46134 (N_46134,N_38565,N_32816);
or U46135 (N_46135,N_38038,N_31341);
xnor U46136 (N_46136,N_37799,N_32087);
nor U46137 (N_46137,N_36340,N_32551);
xor U46138 (N_46138,N_34004,N_36591);
or U46139 (N_46139,N_39371,N_39266);
xnor U46140 (N_46140,N_37979,N_32578);
or U46141 (N_46141,N_39567,N_30120);
and U46142 (N_46142,N_36332,N_36914);
and U46143 (N_46143,N_37630,N_39168);
nor U46144 (N_46144,N_39861,N_35182);
xor U46145 (N_46145,N_38289,N_31708);
xor U46146 (N_46146,N_39686,N_39830);
nand U46147 (N_46147,N_36229,N_38639);
nor U46148 (N_46148,N_39601,N_35945);
and U46149 (N_46149,N_32779,N_38678);
or U46150 (N_46150,N_32373,N_34516);
and U46151 (N_46151,N_30203,N_39603);
or U46152 (N_46152,N_32187,N_37056);
or U46153 (N_46153,N_36506,N_30165);
or U46154 (N_46154,N_31937,N_34321);
xnor U46155 (N_46155,N_31122,N_31753);
or U46156 (N_46156,N_35905,N_31368);
nand U46157 (N_46157,N_37888,N_35157);
xor U46158 (N_46158,N_39172,N_38703);
nand U46159 (N_46159,N_39716,N_34882);
or U46160 (N_46160,N_37258,N_34485);
and U46161 (N_46161,N_33359,N_35378);
and U46162 (N_46162,N_36298,N_35742);
nor U46163 (N_46163,N_36079,N_31646);
nand U46164 (N_46164,N_34144,N_34030);
nand U46165 (N_46165,N_32600,N_39877);
xnor U46166 (N_46166,N_32758,N_37361);
and U46167 (N_46167,N_34275,N_35188);
and U46168 (N_46168,N_35819,N_35829);
or U46169 (N_46169,N_37575,N_38115);
or U46170 (N_46170,N_39544,N_31990);
nor U46171 (N_46171,N_38880,N_39850);
nand U46172 (N_46172,N_35795,N_39051);
xor U46173 (N_46173,N_34186,N_31196);
and U46174 (N_46174,N_32663,N_37396);
xor U46175 (N_46175,N_36045,N_35644);
or U46176 (N_46176,N_33915,N_39143);
or U46177 (N_46177,N_37303,N_34711);
nor U46178 (N_46178,N_37833,N_31995);
nor U46179 (N_46179,N_32287,N_36709);
xor U46180 (N_46180,N_33372,N_32371);
nand U46181 (N_46181,N_31161,N_32343);
or U46182 (N_46182,N_39241,N_32876);
xnor U46183 (N_46183,N_31271,N_39066);
and U46184 (N_46184,N_33739,N_35062);
or U46185 (N_46185,N_31008,N_34250);
or U46186 (N_46186,N_37176,N_34366);
and U46187 (N_46187,N_34781,N_33500);
nor U46188 (N_46188,N_35041,N_33392);
nor U46189 (N_46189,N_33964,N_32474);
xor U46190 (N_46190,N_39480,N_35870);
or U46191 (N_46191,N_31615,N_37749);
and U46192 (N_46192,N_33824,N_35174);
nand U46193 (N_46193,N_32488,N_32129);
or U46194 (N_46194,N_31247,N_39923);
nand U46195 (N_46195,N_34571,N_34694);
nand U46196 (N_46196,N_35839,N_32713);
nand U46197 (N_46197,N_39712,N_37467);
and U46198 (N_46198,N_31850,N_38480);
nor U46199 (N_46199,N_35019,N_36682);
nand U46200 (N_46200,N_39943,N_36988);
or U46201 (N_46201,N_34040,N_31391);
and U46202 (N_46202,N_38789,N_39005);
nor U46203 (N_46203,N_33112,N_39952);
nand U46204 (N_46204,N_34866,N_31970);
nand U46205 (N_46205,N_33573,N_36506);
or U46206 (N_46206,N_39636,N_38545);
nor U46207 (N_46207,N_33458,N_33532);
xnor U46208 (N_46208,N_39453,N_39337);
nand U46209 (N_46209,N_31408,N_31732);
or U46210 (N_46210,N_35990,N_31933);
or U46211 (N_46211,N_36744,N_36741);
or U46212 (N_46212,N_35724,N_39619);
nand U46213 (N_46213,N_31413,N_32229);
nor U46214 (N_46214,N_37445,N_32148);
or U46215 (N_46215,N_32243,N_38080);
xor U46216 (N_46216,N_37841,N_35014);
nand U46217 (N_46217,N_38832,N_31530);
or U46218 (N_46218,N_35119,N_36052);
nand U46219 (N_46219,N_33626,N_32126);
nor U46220 (N_46220,N_30439,N_39776);
and U46221 (N_46221,N_38245,N_37223);
and U46222 (N_46222,N_35854,N_31169);
nand U46223 (N_46223,N_38990,N_34684);
and U46224 (N_46224,N_36853,N_39377);
xor U46225 (N_46225,N_34234,N_38601);
or U46226 (N_46226,N_31113,N_35705);
and U46227 (N_46227,N_36058,N_33817);
or U46228 (N_46228,N_39118,N_37217);
and U46229 (N_46229,N_30648,N_38965);
or U46230 (N_46230,N_31789,N_39405);
and U46231 (N_46231,N_38074,N_30244);
nor U46232 (N_46232,N_39720,N_32945);
nand U46233 (N_46233,N_38649,N_35027);
xor U46234 (N_46234,N_34664,N_31080);
or U46235 (N_46235,N_30014,N_31850);
nor U46236 (N_46236,N_33941,N_36798);
nand U46237 (N_46237,N_33777,N_38855);
nor U46238 (N_46238,N_34717,N_39878);
and U46239 (N_46239,N_33073,N_39381);
nor U46240 (N_46240,N_39046,N_30456);
nand U46241 (N_46241,N_35510,N_30342);
nor U46242 (N_46242,N_37629,N_39465);
nand U46243 (N_46243,N_33760,N_37301);
nor U46244 (N_46244,N_33727,N_39299);
or U46245 (N_46245,N_32943,N_30876);
or U46246 (N_46246,N_30916,N_30767);
nor U46247 (N_46247,N_33183,N_33310);
xor U46248 (N_46248,N_36368,N_37066);
and U46249 (N_46249,N_31070,N_35066);
xnor U46250 (N_46250,N_31262,N_39280);
nor U46251 (N_46251,N_32966,N_39149);
or U46252 (N_46252,N_34345,N_31227);
xnor U46253 (N_46253,N_32249,N_33570);
nor U46254 (N_46254,N_30281,N_39223);
xnor U46255 (N_46255,N_31973,N_36666);
or U46256 (N_46256,N_38852,N_39801);
nor U46257 (N_46257,N_39827,N_37484);
xor U46258 (N_46258,N_37396,N_38495);
nand U46259 (N_46259,N_37231,N_33053);
or U46260 (N_46260,N_38951,N_38256);
and U46261 (N_46261,N_31741,N_31825);
nor U46262 (N_46262,N_38942,N_38763);
and U46263 (N_46263,N_37390,N_32880);
and U46264 (N_46264,N_32544,N_34465);
nor U46265 (N_46265,N_30375,N_37570);
nor U46266 (N_46266,N_38526,N_35490);
or U46267 (N_46267,N_37818,N_31121);
xor U46268 (N_46268,N_34971,N_36416);
nor U46269 (N_46269,N_35283,N_34643);
nor U46270 (N_46270,N_31801,N_37940);
xnor U46271 (N_46271,N_37547,N_32937);
or U46272 (N_46272,N_35895,N_37448);
nand U46273 (N_46273,N_35364,N_39217);
or U46274 (N_46274,N_36447,N_39991);
nand U46275 (N_46275,N_34590,N_39604);
nor U46276 (N_46276,N_32538,N_32182);
xnor U46277 (N_46277,N_30022,N_37626);
nor U46278 (N_46278,N_32962,N_33347);
nor U46279 (N_46279,N_31414,N_33123);
nor U46280 (N_46280,N_39662,N_34045);
and U46281 (N_46281,N_39985,N_38059);
xor U46282 (N_46282,N_36407,N_31034);
xor U46283 (N_46283,N_39729,N_34590);
and U46284 (N_46284,N_34270,N_37871);
xor U46285 (N_46285,N_37814,N_30855);
or U46286 (N_46286,N_35224,N_32272);
and U46287 (N_46287,N_30522,N_32179);
and U46288 (N_46288,N_34672,N_34018);
xnor U46289 (N_46289,N_30276,N_36632);
or U46290 (N_46290,N_36869,N_35369);
nand U46291 (N_46291,N_33269,N_38733);
nand U46292 (N_46292,N_33731,N_31280);
xor U46293 (N_46293,N_30357,N_39076);
nor U46294 (N_46294,N_34636,N_39994);
xnor U46295 (N_46295,N_36505,N_36654);
xnor U46296 (N_46296,N_36266,N_30154);
and U46297 (N_46297,N_31004,N_39616);
and U46298 (N_46298,N_33341,N_32177);
nand U46299 (N_46299,N_34375,N_31310);
and U46300 (N_46300,N_37581,N_32638);
nor U46301 (N_46301,N_37793,N_38771);
and U46302 (N_46302,N_32797,N_32140);
nand U46303 (N_46303,N_33878,N_36307);
nand U46304 (N_46304,N_30739,N_32490);
and U46305 (N_46305,N_34130,N_33126);
nor U46306 (N_46306,N_37358,N_34026);
xor U46307 (N_46307,N_32701,N_34200);
nand U46308 (N_46308,N_38026,N_35121);
or U46309 (N_46309,N_35559,N_33362);
or U46310 (N_46310,N_32519,N_30772);
and U46311 (N_46311,N_38271,N_38933);
and U46312 (N_46312,N_31543,N_38183);
xor U46313 (N_46313,N_36500,N_39578);
nand U46314 (N_46314,N_37064,N_38582);
nor U46315 (N_46315,N_35045,N_30504);
and U46316 (N_46316,N_32572,N_36928);
xor U46317 (N_46317,N_36237,N_33591);
xor U46318 (N_46318,N_36162,N_37288);
nor U46319 (N_46319,N_32056,N_38782);
xnor U46320 (N_46320,N_38718,N_36005);
nand U46321 (N_46321,N_33181,N_31379);
xnor U46322 (N_46322,N_30682,N_32337);
or U46323 (N_46323,N_30867,N_32483);
nand U46324 (N_46324,N_38733,N_31198);
nor U46325 (N_46325,N_39472,N_37917);
or U46326 (N_46326,N_31432,N_32219);
nand U46327 (N_46327,N_35169,N_33732);
xor U46328 (N_46328,N_35087,N_34709);
nor U46329 (N_46329,N_39076,N_33448);
xnor U46330 (N_46330,N_31187,N_34435);
or U46331 (N_46331,N_30785,N_32554);
nor U46332 (N_46332,N_32348,N_39801);
nand U46333 (N_46333,N_33785,N_33986);
or U46334 (N_46334,N_30508,N_37729);
and U46335 (N_46335,N_39996,N_31028);
nand U46336 (N_46336,N_30406,N_38060);
nand U46337 (N_46337,N_39315,N_32805);
nand U46338 (N_46338,N_31726,N_31296);
xnor U46339 (N_46339,N_32283,N_30869);
xnor U46340 (N_46340,N_39312,N_36207);
and U46341 (N_46341,N_39164,N_38030);
nor U46342 (N_46342,N_32660,N_32987);
or U46343 (N_46343,N_36206,N_32364);
nand U46344 (N_46344,N_30615,N_36409);
or U46345 (N_46345,N_36791,N_31663);
nor U46346 (N_46346,N_36992,N_31850);
nand U46347 (N_46347,N_32594,N_33104);
nand U46348 (N_46348,N_35573,N_36856);
and U46349 (N_46349,N_30696,N_32785);
xnor U46350 (N_46350,N_37046,N_37692);
nor U46351 (N_46351,N_36986,N_33124);
nand U46352 (N_46352,N_30516,N_30490);
nor U46353 (N_46353,N_34215,N_37261);
nor U46354 (N_46354,N_39996,N_39656);
nand U46355 (N_46355,N_37025,N_33617);
nand U46356 (N_46356,N_32132,N_32350);
xor U46357 (N_46357,N_30188,N_32296);
nand U46358 (N_46358,N_39629,N_39980);
nand U46359 (N_46359,N_33247,N_33489);
and U46360 (N_46360,N_36357,N_33910);
nand U46361 (N_46361,N_32877,N_38885);
or U46362 (N_46362,N_31860,N_31595);
xor U46363 (N_46363,N_32336,N_38389);
and U46364 (N_46364,N_35317,N_36784);
nor U46365 (N_46365,N_38517,N_39828);
or U46366 (N_46366,N_33897,N_33678);
nor U46367 (N_46367,N_34604,N_37329);
nand U46368 (N_46368,N_30635,N_39827);
xnor U46369 (N_46369,N_38086,N_39996);
xor U46370 (N_46370,N_39922,N_33905);
xor U46371 (N_46371,N_30829,N_38585);
xor U46372 (N_46372,N_31038,N_34435);
xor U46373 (N_46373,N_38712,N_36059);
or U46374 (N_46374,N_37369,N_36271);
nor U46375 (N_46375,N_38792,N_37194);
nor U46376 (N_46376,N_36093,N_37342);
or U46377 (N_46377,N_32592,N_31093);
xnor U46378 (N_46378,N_35435,N_36349);
nor U46379 (N_46379,N_31804,N_39558);
and U46380 (N_46380,N_37444,N_31204);
xnor U46381 (N_46381,N_38308,N_35870);
and U46382 (N_46382,N_31851,N_35352);
nand U46383 (N_46383,N_32653,N_35115);
xnor U46384 (N_46384,N_36469,N_38819);
xnor U46385 (N_46385,N_34465,N_30092);
xor U46386 (N_46386,N_37454,N_32210);
or U46387 (N_46387,N_38345,N_32569);
nand U46388 (N_46388,N_31296,N_37302);
or U46389 (N_46389,N_32531,N_39639);
nand U46390 (N_46390,N_37228,N_35803);
nand U46391 (N_46391,N_34957,N_32380);
or U46392 (N_46392,N_38204,N_35811);
xnor U46393 (N_46393,N_32801,N_39216);
or U46394 (N_46394,N_33775,N_32334);
nand U46395 (N_46395,N_37831,N_30021);
xor U46396 (N_46396,N_37532,N_35800);
nor U46397 (N_46397,N_33927,N_34892);
nand U46398 (N_46398,N_33719,N_38047);
nor U46399 (N_46399,N_38748,N_31139);
and U46400 (N_46400,N_31124,N_32335);
xnor U46401 (N_46401,N_36671,N_33968);
nand U46402 (N_46402,N_34224,N_34302);
nand U46403 (N_46403,N_36463,N_36180);
or U46404 (N_46404,N_33762,N_39000);
nor U46405 (N_46405,N_38336,N_37534);
xnor U46406 (N_46406,N_31960,N_32295);
nand U46407 (N_46407,N_38979,N_33489);
nand U46408 (N_46408,N_36390,N_32897);
or U46409 (N_46409,N_35248,N_32725);
nand U46410 (N_46410,N_32579,N_32185);
nand U46411 (N_46411,N_35122,N_39387);
xor U46412 (N_46412,N_37945,N_39483);
xnor U46413 (N_46413,N_34157,N_32312);
nor U46414 (N_46414,N_36475,N_30939);
nor U46415 (N_46415,N_36828,N_33783);
nand U46416 (N_46416,N_32884,N_39742);
or U46417 (N_46417,N_31624,N_37751);
and U46418 (N_46418,N_37005,N_31580);
nand U46419 (N_46419,N_31384,N_38501);
nand U46420 (N_46420,N_38144,N_35155);
and U46421 (N_46421,N_32805,N_32452);
nor U46422 (N_46422,N_36512,N_39786);
nor U46423 (N_46423,N_34897,N_39998);
and U46424 (N_46424,N_37811,N_30918);
or U46425 (N_46425,N_39567,N_35282);
or U46426 (N_46426,N_36791,N_34537);
xnor U46427 (N_46427,N_37943,N_30899);
or U46428 (N_46428,N_33340,N_34258);
or U46429 (N_46429,N_31975,N_32430);
xor U46430 (N_46430,N_36426,N_32072);
and U46431 (N_46431,N_35367,N_35285);
nor U46432 (N_46432,N_37840,N_37268);
nand U46433 (N_46433,N_34042,N_30934);
nor U46434 (N_46434,N_36389,N_36883);
or U46435 (N_46435,N_32066,N_30392);
nor U46436 (N_46436,N_38108,N_33398);
nand U46437 (N_46437,N_39601,N_33638);
and U46438 (N_46438,N_36781,N_34579);
or U46439 (N_46439,N_35283,N_30239);
xnor U46440 (N_46440,N_31505,N_38284);
xor U46441 (N_46441,N_32311,N_34955);
nand U46442 (N_46442,N_35034,N_32946);
xor U46443 (N_46443,N_34159,N_35591);
nand U46444 (N_46444,N_32869,N_33792);
nand U46445 (N_46445,N_30364,N_31629);
nor U46446 (N_46446,N_34297,N_34463);
nor U46447 (N_46447,N_35258,N_36424);
xnor U46448 (N_46448,N_37663,N_38641);
nor U46449 (N_46449,N_31544,N_34163);
and U46450 (N_46450,N_38860,N_31760);
xnor U46451 (N_46451,N_37947,N_35985);
nand U46452 (N_46452,N_38353,N_39040);
or U46453 (N_46453,N_36644,N_37377);
nor U46454 (N_46454,N_35512,N_34364);
xor U46455 (N_46455,N_38439,N_39474);
and U46456 (N_46456,N_35152,N_39593);
nand U46457 (N_46457,N_31880,N_32566);
nor U46458 (N_46458,N_38481,N_36270);
nor U46459 (N_46459,N_32578,N_38939);
and U46460 (N_46460,N_34062,N_37478);
xnor U46461 (N_46461,N_30283,N_39570);
xnor U46462 (N_46462,N_34562,N_30090);
xnor U46463 (N_46463,N_38900,N_38963);
xnor U46464 (N_46464,N_35401,N_30020);
xor U46465 (N_46465,N_35191,N_34751);
or U46466 (N_46466,N_38041,N_35596);
or U46467 (N_46467,N_32367,N_32495);
xor U46468 (N_46468,N_35589,N_37737);
nand U46469 (N_46469,N_38840,N_34020);
or U46470 (N_46470,N_35199,N_36389);
or U46471 (N_46471,N_30816,N_36545);
and U46472 (N_46472,N_37927,N_31024);
and U46473 (N_46473,N_35074,N_39494);
and U46474 (N_46474,N_31646,N_30765);
or U46475 (N_46475,N_33059,N_39046);
and U46476 (N_46476,N_32470,N_32262);
xnor U46477 (N_46477,N_34987,N_30068);
or U46478 (N_46478,N_37587,N_34320);
nor U46479 (N_46479,N_36270,N_36625);
nand U46480 (N_46480,N_35023,N_36020);
nor U46481 (N_46481,N_35274,N_34233);
nor U46482 (N_46482,N_38736,N_31524);
xnor U46483 (N_46483,N_33505,N_30017);
or U46484 (N_46484,N_37919,N_39600);
xnor U46485 (N_46485,N_31079,N_39020);
and U46486 (N_46486,N_31827,N_38237);
and U46487 (N_46487,N_34383,N_33839);
and U46488 (N_46488,N_31278,N_35630);
nand U46489 (N_46489,N_39543,N_38597);
and U46490 (N_46490,N_30451,N_33466);
or U46491 (N_46491,N_38391,N_38458);
nand U46492 (N_46492,N_37812,N_37146);
nor U46493 (N_46493,N_37101,N_39235);
xnor U46494 (N_46494,N_38075,N_30727);
or U46495 (N_46495,N_32078,N_30121);
and U46496 (N_46496,N_37040,N_30058);
nor U46497 (N_46497,N_31018,N_37064);
and U46498 (N_46498,N_39651,N_30103);
or U46499 (N_46499,N_34542,N_31916);
nor U46500 (N_46500,N_31064,N_38520);
nor U46501 (N_46501,N_33260,N_31810);
and U46502 (N_46502,N_35945,N_31586);
xor U46503 (N_46503,N_34228,N_31949);
nor U46504 (N_46504,N_38991,N_33370);
xor U46505 (N_46505,N_30139,N_35222);
xor U46506 (N_46506,N_34786,N_33621);
xor U46507 (N_46507,N_34853,N_39120);
nor U46508 (N_46508,N_38295,N_37261);
or U46509 (N_46509,N_31508,N_32273);
nor U46510 (N_46510,N_36372,N_35797);
and U46511 (N_46511,N_36238,N_31026);
xnor U46512 (N_46512,N_38539,N_31606);
xor U46513 (N_46513,N_38631,N_32588);
nor U46514 (N_46514,N_37617,N_35343);
or U46515 (N_46515,N_35797,N_30045);
xnor U46516 (N_46516,N_30918,N_32226);
and U46517 (N_46517,N_35029,N_34039);
nor U46518 (N_46518,N_37017,N_30365);
or U46519 (N_46519,N_31427,N_31037);
and U46520 (N_46520,N_34231,N_37800);
xnor U46521 (N_46521,N_34007,N_31967);
or U46522 (N_46522,N_38611,N_31781);
or U46523 (N_46523,N_38911,N_38198);
nor U46524 (N_46524,N_34374,N_30042);
nand U46525 (N_46525,N_37608,N_37604);
or U46526 (N_46526,N_34012,N_35497);
or U46527 (N_46527,N_35025,N_32594);
or U46528 (N_46528,N_32723,N_38760);
and U46529 (N_46529,N_31559,N_37239);
xor U46530 (N_46530,N_39681,N_31742);
xor U46531 (N_46531,N_31619,N_38420);
or U46532 (N_46532,N_34308,N_36591);
nand U46533 (N_46533,N_31333,N_37788);
and U46534 (N_46534,N_38717,N_33330);
or U46535 (N_46535,N_30796,N_31151);
and U46536 (N_46536,N_35192,N_39553);
nand U46537 (N_46537,N_30138,N_38449);
nand U46538 (N_46538,N_30904,N_38534);
nor U46539 (N_46539,N_38789,N_35844);
nand U46540 (N_46540,N_32522,N_38586);
and U46541 (N_46541,N_34494,N_38353);
nor U46542 (N_46542,N_32080,N_32529);
nor U46543 (N_46543,N_36184,N_32399);
xor U46544 (N_46544,N_38266,N_33142);
xnor U46545 (N_46545,N_32700,N_37198);
xnor U46546 (N_46546,N_34497,N_31317);
and U46547 (N_46547,N_37069,N_33380);
xor U46548 (N_46548,N_33065,N_39088);
xnor U46549 (N_46549,N_34358,N_34626);
xnor U46550 (N_46550,N_30257,N_36518);
and U46551 (N_46551,N_36393,N_32465);
or U46552 (N_46552,N_33880,N_36038);
nor U46553 (N_46553,N_37825,N_30806);
nand U46554 (N_46554,N_35364,N_39159);
or U46555 (N_46555,N_38924,N_39270);
xnor U46556 (N_46556,N_38986,N_33946);
nor U46557 (N_46557,N_35958,N_30520);
nor U46558 (N_46558,N_37683,N_31044);
nor U46559 (N_46559,N_30171,N_35854);
and U46560 (N_46560,N_33570,N_30461);
or U46561 (N_46561,N_31946,N_37417);
nand U46562 (N_46562,N_33163,N_37474);
or U46563 (N_46563,N_36748,N_38930);
nor U46564 (N_46564,N_35209,N_34583);
and U46565 (N_46565,N_38985,N_36139);
xnor U46566 (N_46566,N_32441,N_36798);
and U46567 (N_46567,N_30615,N_31902);
or U46568 (N_46568,N_36052,N_38413);
and U46569 (N_46569,N_36292,N_35372);
nand U46570 (N_46570,N_31582,N_33964);
or U46571 (N_46571,N_33831,N_39177);
nor U46572 (N_46572,N_39798,N_31497);
nor U46573 (N_46573,N_32149,N_30817);
nand U46574 (N_46574,N_38972,N_37508);
nand U46575 (N_46575,N_39348,N_39890);
and U46576 (N_46576,N_39357,N_38837);
nand U46577 (N_46577,N_33137,N_36172);
and U46578 (N_46578,N_36053,N_37478);
xnor U46579 (N_46579,N_38801,N_33507);
xnor U46580 (N_46580,N_34054,N_32648);
and U46581 (N_46581,N_36625,N_36006);
xnor U46582 (N_46582,N_39947,N_38632);
nand U46583 (N_46583,N_38630,N_31070);
nor U46584 (N_46584,N_39156,N_30456);
and U46585 (N_46585,N_31989,N_31179);
or U46586 (N_46586,N_32203,N_38481);
xor U46587 (N_46587,N_32040,N_35903);
xor U46588 (N_46588,N_32163,N_33518);
nand U46589 (N_46589,N_38032,N_34388);
xnor U46590 (N_46590,N_37427,N_39745);
and U46591 (N_46591,N_35886,N_30594);
nor U46592 (N_46592,N_33261,N_30503);
nand U46593 (N_46593,N_32788,N_36135);
nand U46594 (N_46594,N_37536,N_39775);
nor U46595 (N_46595,N_32066,N_35704);
xnor U46596 (N_46596,N_30457,N_33232);
nand U46597 (N_46597,N_37607,N_38665);
or U46598 (N_46598,N_32537,N_30277);
xor U46599 (N_46599,N_37094,N_38613);
and U46600 (N_46600,N_37783,N_38215);
nand U46601 (N_46601,N_39505,N_37918);
and U46602 (N_46602,N_35555,N_33725);
nand U46603 (N_46603,N_39375,N_37287);
nand U46604 (N_46604,N_32512,N_38521);
nor U46605 (N_46605,N_33060,N_31076);
xnor U46606 (N_46606,N_38835,N_37655);
and U46607 (N_46607,N_36500,N_32138);
and U46608 (N_46608,N_39654,N_31356);
and U46609 (N_46609,N_32695,N_39406);
nand U46610 (N_46610,N_38440,N_36227);
xnor U46611 (N_46611,N_30869,N_35052);
and U46612 (N_46612,N_39443,N_37549);
and U46613 (N_46613,N_31074,N_38198);
xor U46614 (N_46614,N_35793,N_37815);
xor U46615 (N_46615,N_37887,N_31508);
nand U46616 (N_46616,N_30775,N_39642);
or U46617 (N_46617,N_30654,N_36380);
or U46618 (N_46618,N_33793,N_36281);
and U46619 (N_46619,N_31423,N_34608);
nand U46620 (N_46620,N_39038,N_35951);
and U46621 (N_46621,N_35744,N_39642);
xor U46622 (N_46622,N_32791,N_35185);
nor U46623 (N_46623,N_30605,N_39313);
or U46624 (N_46624,N_37700,N_35916);
xor U46625 (N_46625,N_34006,N_37104);
nand U46626 (N_46626,N_35114,N_31358);
and U46627 (N_46627,N_33671,N_38227);
xor U46628 (N_46628,N_39133,N_30463);
nand U46629 (N_46629,N_32443,N_36555);
xnor U46630 (N_46630,N_35752,N_34508);
nor U46631 (N_46631,N_39986,N_33734);
xnor U46632 (N_46632,N_33365,N_34029);
nor U46633 (N_46633,N_35936,N_38834);
or U46634 (N_46634,N_31279,N_32926);
nor U46635 (N_46635,N_39439,N_37041);
nor U46636 (N_46636,N_32600,N_34182);
nor U46637 (N_46637,N_34673,N_34604);
and U46638 (N_46638,N_38804,N_33626);
and U46639 (N_46639,N_30404,N_30616);
and U46640 (N_46640,N_34147,N_33053);
xor U46641 (N_46641,N_36964,N_37414);
xnor U46642 (N_46642,N_36463,N_35055);
or U46643 (N_46643,N_39158,N_36713);
or U46644 (N_46644,N_33545,N_32418);
and U46645 (N_46645,N_35274,N_35612);
nand U46646 (N_46646,N_36130,N_33077);
or U46647 (N_46647,N_33888,N_37194);
or U46648 (N_46648,N_38872,N_36738);
and U46649 (N_46649,N_37183,N_36302);
nor U46650 (N_46650,N_37194,N_35878);
nor U46651 (N_46651,N_34751,N_36773);
and U46652 (N_46652,N_36426,N_33872);
or U46653 (N_46653,N_33105,N_38217);
nor U46654 (N_46654,N_35676,N_36391);
or U46655 (N_46655,N_37061,N_39430);
or U46656 (N_46656,N_37191,N_32964);
xnor U46657 (N_46657,N_31988,N_39704);
and U46658 (N_46658,N_36924,N_36003);
xnor U46659 (N_46659,N_30312,N_38233);
nor U46660 (N_46660,N_36474,N_38106);
and U46661 (N_46661,N_32239,N_34141);
and U46662 (N_46662,N_36385,N_39331);
xnor U46663 (N_46663,N_35169,N_31193);
nor U46664 (N_46664,N_34669,N_34016);
nand U46665 (N_46665,N_36930,N_38573);
or U46666 (N_46666,N_33521,N_36395);
nand U46667 (N_46667,N_34315,N_37812);
nor U46668 (N_46668,N_33603,N_35017);
nand U46669 (N_46669,N_39703,N_34470);
xor U46670 (N_46670,N_31468,N_39505);
and U46671 (N_46671,N_36067,N_38583);
or U46672 (N_46672,N_33416,N_36243);
and U46673 (N_46673,N_36546,N_34246);
nor U46674 (N_46674,N_36534,N_37681);
and U46675 (N_46675,N_35668,N_32645);
or U46676 (N_46676,N_31168,N_38003);
xnor U46677 (N_46677,N_35663,N_39498);
or U46678 (N_46678,N_31501,N_38773);
and U46679 (N_46679,N_30645,N_33655);
xnor U46680 (N_46680,N_35506,N_30356);
xnor U46681 (N_46681,N_33393,N_30020);
nor U46682 (N_46682,N_33939,N_30160);
xor U46683 (N_46683,N_38556,N_31414);
nand U46684 (N_46684,N_37633,N_31134);
nand U46685 (N_46685,N_33008,N_34116);
xor U46686 (N_46686,N_30215,N_33777);
or U46687 (N_46687,N_33983,N_34258);
nor U46688 (N_46688,N_38921,N_33951);
nor U46689 (N_46689,N_36131,N_30273);
and U46690 (N_46690,N_36873,N_32784);
xor U46691 (N_46691,N_35974,N_37277);
nand U46692 (N_46692,N_39059,N_34046);
xnor U46693 (N_46693,N_32802,N_31415);
xor U46694 (N_46694,N_30187,N_34848);
nor U46695 (N_46695,N_35901,N_35777);
xor U46696 (N_46696,N_35982,N_37717);
or U46697 (N_46697,N_33024,N_38204);
nor U46698 (N_46698,N_30085,N_39989);
or U46699 (N_46699,N_35741,N_31009);
and U46700 (N_46700,N_34023,N_35310);
xor U46701 (N_46701,N_33799,N_38653);
nand U46702 (N_46702,N_37007,N_30876);
or U46703 (N_46703,N_38085,N_35601);
nor U46704 (N_46704,N_35960,N_36395);
or U46705 (N_46705,N_34927,N_37052);
or U46706 (N_46706,N_33926,N_32409);
and U46707 (N_46707,N_30636,N_35656);
nand U46708 (N_46708,N_38061,N_30818);
nand U46709 (N_46709,N_34160,N_39396);
and U46710 (N_46710,N_38414,N_32587);
xor U46711 (N_46711,N_32720,N_37442);
nor U46712 (N_46712,N_34987,N_36653);
or U46713 (N_46713,N_39680,N_31745);
nand U46714 (N_46714,N_35463,N_31437);
nand U46715 (N_46715,N_33059,N_33726);
xor U46716 (N_46716,N_34620,N_39567);
nand U46717 (N_46717,N_34394,N_34653);
xnor U46718 (N_46718,N_38994,N_30872);
nor U46719 (N_46719,N_38631,N_33383);
and U46720 (N_46720,N_31883,N_38370);
nor U46721 (N_46721,N_35829,N_36853);
or U46722 (N_46722,N_37125,N_33118);
or U46723 (N_46723,N_31048,N_38455);
or U46724 (N_46724,N_33719,N_36149);
nor U46725 (N_46725,N_39052,N_39632);
or U46726 (N_46726,N_39364,N_38021);
nand U46727 (N_46727,N_35479,N_35293);
nand U46728 (N_46728,N_34770,N_33891);
or U46729 (N_46729,N_30631,N_36260);
nor U46730 (N_46730,N_33389,N_32373);
nand U46731 (N_46731,N_30058,N_38181);
or U46732 (N_46732,N_38157,N_39509);
or U46733 (N_46733,N_35058,N_30798);
and U46734 (N_46734,N_38589,N_32497);
xor U46735 (N_46735,N_36107,N_30051);
xor U46736 (N_46736,N_35996,N_30709);
nand U46737 (N_46737,N_33576,N_36735);
xor U46738 (N_46738,N_35850,N_30379);
nor U46739 (N_46739,N_30518,N_32698);
nand U46740 (N_46740,N_33649,N_39717);
xor U46741 (N_46741,N_32277,N_35302);
and U46742 (N_46742,N_32605,N_37489);
and U46743 (N_46743,N_31091,N_39542);
or U46744 (N_46744,N_32737,N_34130);
xor U46745 (N_46745,N_34513,N_34002);
or U46746 (N_46746,N_39790,N_37526);
nor U46747 (N_46747,N_36052,N_38185);
or U46748 (N_46748,N_34767,N_33737);
nor U46749 (N_46749,N_31465,N_30795);
and U46750 (N_46750,N_30449,N_31073);
or U46751 (N_46751,N_31493,N_36913);
nand U46752 (N_46752,N_36781,N_32448);
or U46753 (N_46753,N_30054,N_32186);
and U46754 (N_46754,N_35702,N_34825);
nor U46755 (N_46755,N_38186,N_34849);
nor U46756 (N_46756,N_39042,N_31604);
xor U46757 (N_46757,N_31096,N_37750);
xor U46758 (N_46758,N_33602,N_31958);
nor U46759 (N_46759,N_35428,N_36204);
or U46760 (N_46760,N_36444,N_37157);
nor U46761 (N_46761,N_33311,N_31802);
xor U46762 (N_46762,N_38228,N_33434);
nor U46763 (N_46763,N_33239,N_30064);
xnor U46764 (N_46764,N_30811,N_37983);
and U46765 (N_46765,N_39376,N_33789);
xor U46766 (N_46766,N_38931,N_33925);
or U46767 (N_46767,N_36645,N_39787);
xor U46768 (N_46768,N_37445,N_30184);
nor U46769 (N_46769,N_37371,N_31389);
and U46770 (N_46770,N_36618,N_35940);
nand U46771 (N_46771,N_36900,N_39717);
xnor U46772 (N_46772,N_34555,N_35386);
xor U46773 (N_46773,N_37260,N_39826);
xor U46774 (N_46774,N_34036,N_30043);
nor U46775 (N_46775,N_38527,N_33667);
and U46776 (N_46776,N_35272,N_39337);
or U46777 (N_46777,N_32318,N_31576);
or U46778 (N_46778,N_31346,N_38492);
and U46779 (N_46779,N_39743,N_34249);
xnor U46780 (N_46780,N_34243,N_38890);
nor U46781 (N_46781,N_36000,N_36865);
xnor U46782 (N_46782,N_33529,N_31371);
nand U46783 (N_46783,N_32274,N_32001);
xnor U46784 (N_46784,N_36311,N_31309);
nor U46785 (N_46785,N_35982,N_33514);
nand U46786 (N_46786,N_32275,N_32741);
or U46787 (N_46787,N_35498,N_36551);
and U46788 (N_46788,N_39461,N_30615);
xor U46789 (N_46789,N_31061,N_33303);
nand U46790 (N_46790,N_36691,N_38645);
nand U46791 (N_46791,N_34535,N_39520);
nor U46792 (N_46792,N_30013,N_39974);
nand U46793 (N_46793,N_36158,N_35123);
xor U46794 (N_46794,N_39010,N_39149);
or U46795 (N_46795,N_30786,N_39186);
xnor U46796 (N_46796,N_30427,N_34403);
nand U46797 (N_46797,N_34450,N_36715);
nor U46798 (N_46798,N_35183,N_32367);
or U46799 (N_46799,N_35669,N_37748);
and U46800 (N_46800,N_30568,N_37362);
and U46801 (N_46801,N_36616,N_33796);
xor U46802 (N_46802,N_33734,N_37948);
nor U46803 (N_46803,N_36752,N_30055);
nand U46804 (N_46804,N_37823,N_32818);
nor U46805 (N_46805,N_34897,N_33994);
xor U46806 (N_46806,N_39564,N_34179);
nor U46807 (N_46807,N_36040,N_38406);
xor U46808 (N_46808,N_33385,N_31341);
nand U46809 (N_46809,N_34470,N_35905);
or U46810 (N_46810,N_38362,N_35835);
xor U46811 (N_46811,N_37543,N_30932);
or U46812 (N_46812,N_39045,N_32693);
xor U46813 (N_46813,N_32838,N_38218);
xor U46814 (N_46814,N_38691,N_30944);
and U46815 (N_46815,N_35340,N_32503);
xor U46816 (N_46816,N_30309,N_38705);
nand U46817 (N_46817,N_36972,N_32246);
xor U46818 (N_46818,N_31006,N_32826);
nand U46819 (N_46819,N_39331,N_33602);
xor U46820 (N_46820,N_36927,N_33832);
or U46821 (N_46821,N_35204,N_39070);
nor U46822 (N_46822,N_38116,N_30042);
nor U46823 (N_46823,N_39969,N_35320);
and U46824 (N_46824,N_37101,N_36712);
or U46825 (N_46825,N_35932,N_32419);
nand U46826 (N_46826,N_36774,N_33333);
and U46827 (N_46827,N_39883,N_36849);
nor U46828 (N_46828,N_33659,N_37459);
xnor U46829 (N_46829,N_35969,N_30126);
nand U46830 (N_46830,N_30767,N_33169);
or U46831 (N_46831,N_37804,N_33934);
or U46832 (N_46832,N_36350,N_37370);
or U46833 (N_46833,N_37493,N_37330);
or U46834 (N_46834,N_36685,N_32155);
nor U46835 (N_46835,N_37346,N_30097);
xnor U46836 (N_46836,N_34203,N_32870);
or U46837 (N_46837,N_39149,N_31262);
nor U46838 (N_46838,N_36671,N_36692);
or U46839 (N_46839,N_32276,N_38119);
nand U46840 (N_46840,N_36399,N_37638);
nand U46841 (N_46841,N_34869,N_33124);
xnor U46842 (N_46842,N_39840,N_34382);
nand U46843 (N_46843,N_38719,N_31064);
and U46844 (N_46844,N_39758,N_33544);
nand U46845 (N_46845,N_31444,N_35676);
nor U46846 (N_46846,N_32363,N_38456);
nor U46847 (N_46847,N_38808,N_30464);
nand U46848 (N_46848,N_38442,N_39405);
xnor U46849 (N_46849,N_32950,N_38910);
nor U46850 (N_46850,N_39631,N_30236);
nor U46851 (N_46851,N_39491,N_32056);
and U46852 (N_46852,N_35325,N_35059);
and U46853 (N_46853,N_32940,N_31369);
or U46854 (N_46854,N_32015,N_31236);
and U46855 (N_46855,N_31299,N_31237);
nor U46856 (N_46856,N_35016,N_38588);
xnor U46857 (N_46857,N_37476,N_34395);
and U46858 (N_46858,N_33521,N_31546);
xnor U46859 (N_46859,N_36472,N_38148);
xor U46860 (N_46860,N_30646,N_36616);
nor U46861 (N_46861,N_37212,N_32108);
xor U46862 (N_46862,N_30346,N_30751);
nor U46863 (N_46863,N_32304,N_38586);
or U46864 (N_46864,N_31106,N_33078);
xor U46865 (N_46865,N_36162,N_33239);
and U46866 (N_46866,N_35670,N_39746);
or U46867 (N_46867,N_31595,N_34105);
nand U46868 (N_46868,N_35989,N_30290);
xor U46869 (N_46869,N_31651,N_34248);
nor U46870 (N_46870,N_33548,N_33241);
or U46871 (N_46871,N_32317,N_33150);
or U46872 (N_46872,N_31659,N_39548);
nand U46873 (N_46873,N_33968,N_32842);
and U46874 (N_46874,N_39202,N_36817);
nor U46875 (N_46875,N_33543,N_30146);
or U46876 (N_46876,N_32295,N_30344);
and U46877 (N_46877,N_30849,N_30769);
nand U46878 (N_46878,N_38586,N_35020);
xor U46879 (N_46879,N_34457,N_31775);
or U46880 (N_46880,N_34868,N_37314);
or U46881 (N_46881,N_37190,N_34235);
xor U46882 (N_46882,N_34673,N_35105);
nor U46883 (N_46883,N_34321,N_33899);
nor U46884 (N_46884,N_31932,N_30381);
or U46885 (N_46885,N_37810,N_38440);
and U46886 (N_46886,N_39843,N_33418);
nand U46887 (N_46887,N_39611,N_30598);
nor U46888 (N_46888,N_33336,N_38771);
xor U46889 (N_46889,N_36779,N_30639);
xor U46890 (N_46890,N_35945,N_36400);
xor U46891 (N_46891,N_30820,N_33060);
nor U46892 (N_46892,N_30878,N_36988);
nor U46893 (N_46893,N_34703,N_32149);
nor U46894 (N_46894,N_35253,N_36470);
or U46895 (N_46895,N_37412,N_32773);
and U46896 (N_46896,N_37819,N_32451);
nand U46897 (N_46897,N_36788,N_35940);
nor U46898 (N_46898,N_32494,N_37917);
xor U46899 (N_46899,N_36077,N_36174);
nand U46900 (N_46900,N_32576,N_38540);
xor U46901 (N_46901,N_37968,N_31524);
and U46902 (N_46902,N_35479,N_31913);
nand U46903 (N_46903,N_36588,N_37016);
and U46904 (N_46904,N_34906,N_32339);
nand U46905 (N_46905,N_39172,N_37213);
and U46906 (N_46906,N_35911,N_35956);
nor U46907 (N_46907,N_32841,N_34498);
nor U46908 (N_46908,N_34044,N_39024);
nand U46909 (N_46909,N_37364,N_30718);
nor U46910 (N_46910,N_33880,N_32167);
nand U46911 (N_46911,N_34686,N_31143);
xnor U46912 (N_46912,N_38932,N_34279);
xor U46913 (N_46913,N_33295,N_37936);
nor U46914 (N_46914,N_31323,N_31279);
xnor U46915 (N_46915,N_32713,N_31868);
nand U46916 (N_46916,N_32957,N_39867);
or U46917 (N_46917,N_30206,N_33281);
xor U46918 (N_46918,N_36695,N_34195);
xor U46919 (N_46919,N_33822,N_38849);
xor U46920 (N_46920,N_35853,N_33511);
and U46921 (N_46921,N_31225,N_38176);
nand U46922 (N_46922,N_34051,N_37717);
nor U46923 (N_46923,N_30294,N_34507);
nor U46924 (N_46924,N_36776,N_31763);
xor U46925 (N_46925,N_31861,N_35259);
nand U46926 (N_46926,N_38348,N_33521);
and U46927 (N_46927,N_37563,N_33617);
nor U46928 (N_46928,N_30099,N_39720);
or U46929 (N_46929,N_34562,N_32717);
and U46930 (N_46930,N_39834,N_39817);
nand U46931 (N_46931,N_33994,N_35361);
xnor U46932 (N_46932,N_31722,N_37910);
nand U46933 (N_46933,N_32068,N_30621);
or U46934 (N_46934,N_37112,N_34880);
and U46935 (N_46935,N_35721,N_37946);
or U46936 (N_46936,N_32446,N_31235);
and U46937 (N_46937,N_34898,N_34492);
and U46938 (N_46938,N_36560,N_34470);
nand U46939 (N_46939,N_33592,N_38467);
nand U46940 (N_46940,N_30676,N_35278);
xnor U46941 (N_46941,N_36695,N_33952);
nand U46942 (N_46942,N_32542,N_34284);
nand U46943 (N_46943,N_33564,N_31063);
nor U46944 (N_46944,N_39078,N_32192);
or U46945 (N_46945,N_39853,N_39329);
nor U46946 (N_46946,N_32931,N_33595);
xnor U46947 (N_46947,N_32483,N_32522);
nand U46948 (N_46948,N_36912,N_31245);
nand U46949 (N_46949,N_36387,N_35018);
or U46950 (N_46950,N_32057,N_33985);
and U46951 (N_46951,N_36676,N_34760);
xor U46952 (N_46952,N_34299,N_36096);
xor U46953 (N_46953,N_38842,N_33676);
xnor U46954 (N_46954,N_36333,N_37179);
nor U46955 (N_46955,N_38027,N_37213);
nor U46956 (N_46956,N_34929,N_31703);
and U46957 (N_46957,N_37900,N_32756);
or U46958 (N_46958,N_35710,N_34169);
or U46959 (N_46959,N_36881,N_39424);
xnor U46960 (N_46960,N_34352,N_33369);
nor U46961 (N_46961,N_38489,N_37457);
or U46962 (N_46962,N_31325,N_32535);
nor U46963 (N_46963,N_33533,N_34132);
and U46964 (N_46964,N_33506,N_35543);
nand U46965 (N_46965,N_37976,N_36979);
nor U46966 (N_46966,N_38397,N_38544);
nand U46967 (N_46967,N_35277,N_32770);
nand U46968 (N_46968,N_36832,N_39407);
nor U46969 (N_46969,N_38017,N_35338);
or U46970 (N_46970,N_31875,N_32924);
nor U46971 (N_46971,N_39673,N_35350);
or U46972 (N_46972,N_30013,N_33849);
or U46973 (N_46973,N_37560,N_37834);
nand U46974 (N_46974,N_35708,N_34907);
or U46975 (N_46975,N_31767,N_34672);
or U46976 (N_46976,N_33607,N_38416);
nand U46977 (N_46977,N_34387,N_34871);
xnor U46978 (N_46978,N_38149,N_38155);
or U46979 (N_46979,N_32455,N_33622);
nand U46980 (N_46980,N_33575,N_30517);
or U46981 (N_46981,N_34322,N_33536);
xor U46982 (N_46982,N_34213,N_31956);
nand U46983 (N_46983,N_34893,N_30488);
xor U46984 (N_46984,N_34558,N_37331);
or U46985 (N_46985,N_31749,N_33846);
nand U46986 (N_46986,N_31538,N_32378);
xor U46987 (N_46987,N_30857,N_39369);
or U46988 (N_46988,N_38746,N_36451);
nand U46989 (N_46989,N_34752,N_39773);
nand U46990 (N_46990,N_34446,N_35136);
and U46991 (N_46991,N_30539,N_35461);
xor U46992 (N_46992,N_34053,N_36253);
or U46993 (N_46993,N_34905,N_37269);
nand U46994 (N_46994,N_32634,N_33645);
xnor U46995 (N_46995,N_33739,N_35452);
and U46996 (N_46996,N_38128,N_30412);
nand U46997 (N_46997,N_33446,N_30839);
or U46998 (N_46998,N_36073,N_35603);
nand U46999 (N_46999,N_30736,N_32677);
nor U47000 (N_47000,N_33535,N_36949);
or U47001 (N_47001,N_38970,N_39672);
nor U47002 (N_47002,N_35486,N_39298);
and U47003 (N_47003,N_32741,N_31428);
xnor U47004 (N_47004,N_36586,N_34551);
xor U47005 (N_47005,N_37349,N_38422);
nand U47006 (N_47006,N_36502,N_37233);
nand U47007 (N_47007,N_36459,N_32462);
nor U47008 (N_47008,N_30668,N_30149);
nor U47009 (N_47009,N_38736,N_30473);
or U47010 (N_47010,N_35491,N_37827);
nor U47011 (N_47011,N_31218,N_38373);
or U47012 (N_47012,N_35566,N_36182);
nor U47013 (N_47013,N_34030,N_35865);
xnor U47014 (N_47014,N_34843,N_36038);
or U47015 (N_47015,N_32154,N_38052);
xor U47016 (N_47016,N_32180,N_30864);
and U47017 (N_47017,N_38593,N_33915);
and U47018 (N_47018,N_32628,N_30834);
and U47019 (N_47019,N_32988,N_36783);
and U47020 (N_47020,N_32289,N_36401);
xor U47021 (N_47021,N_31744,N_35123);
nor U47022 (N_47022,N_38955,N_30808);
and U47023 (N_47023,N_34501,N_31362);
and U47024 (N_47024,N_32760,N_38429);
and U47025 (N_47025,N_33631,N_35448);
nor U47026 (N_47026,N_34925,N_32862);
nand U47027 (N_47027,N_35072,N_38791);
nor U47028 (N_47028,N_34587,N_32145);
nand U47029 (N_47029,N_38710,N_38097);
or U47030 (N_47030,N_39284,N_36524);
nand U47031 (N_47031,N_37362,N_32323);
nor U47032 (N_47032,N_38344,N_32237);
nand U47033 (N_47033,N_34476,N_39778);
xor U47034 (N_47034,N_38038,N_39846);
nor U47035 (N_47035,N_38399,N_32727);
nor U47036 (N_47036,N_30464,N_38057);
nor U47037 (N_47037,N_32795,N_32847);
or U47038 (N_47038,N_39712,N_37611);
and U47039 (N_47039,N_39469,N_32309);
nor U47040 (N_47040,N_33170,N_39317);
xor U47041 (N_47041,N_34977,N_30851);
nand U47042 (N_47042,N_37969,N_35255);
nor U47043 (N_47043,N_35164,N_36508);
xor U47044 (N_47044,N_32513,N_35138);
nand U47045 (N_47045,N_38369,N_37225);
and U47046 (N_47046,N_33739,N_35537);
and U47047 (N_47047,N_36225,N_31931);
nor U47048 (N_47048,N_37858,N_38407);
and U47049 (N_47049,N_34343,N_34686);
or U47050 (N_47050,N_31346,N_38201);
nor U47051 (N_47051,N_32115,N_36026);
nand U47052 (N_47052,N_36635,N_39903);
and U47053 (N_47053,N_32055,N_35775);
and U47054 (N_47054,N_39516,N_31313);
xor U47055 (N_47055,N_36118,N_32513);
or U47056 (N_47056,N_35737,N_37420);
and U47057 (N_47057,N_36720,N_34551);
nand U47058 (N_47058,N_36176,N_30859);
or U47059 (N_47059,N_30143,N_38980);
nand U47060 (N_47060,N_33822,N_37685);
or U47061 (N_47061,N_39244,N_38056);
or U47062 (N_47062,N_36429,N_38629);
or U47063 (N_47063,N_34459,N_35638);
and U47064 (N_47064,N_34899,N_37167);
nand U47065 (N_47065,N_36277,N_39802);
or U47066 (N_47066,N_33623,N_38014);
nor U47067 (N_47067,N_38948,N_36337);
and U47068 (N_47068,N_30858,N_37733);
and U47069 (N_47069,N_33547,N_37105);
nand U47070 (N_47070,N_37112,N_32517);
nand U47071 (N_47071,N_38495,N_30804);
nor U47072 (N_47072,N_32674,N_31909);
xor U47073 (N_47073,N_38037,N_38720);
nand U47074 (N_47074,N_31165,N_38044);
nand U47075 (N_47075,N_35725,N_39294);
nor U47076 (N_47076,N_33862,N_38270);
nor U47077 (N_47077,N_39401,N_31013);
xor U47078 (N_47078,N_35979,N_35067);
or U47079 (N_47079,N_33850,N_38981);
or U47080 (N_47080,N_39216,N_38566);
and U47081 (N_47081,N_32762,N_34339);
or U47082 (N_47082,N_31970,N_33967);
nor U47083 (N_47083,N_31879,N_36188);
nor U47084 (N_47084,N_32945,N_33397);
nor U47085 (N_47085,N_38774,N_37361);
or U47086 (N_47086,N_34309,N_37328);
nand U47087 (N_47087,N_30609,N_38739);
or U47088 (N_47088,N_31103,N_34255);
or U47089 (N_47089,N_38896,N_34293);
nand U47090 (N_47090,N_30770,N_35376);
or U47091 (N_47091,N_30809,N_30070);
and U47092 (N_47092,N_39018,N_31645);
and U47093 (N_47093,N_30819,N_39618);
xor U47094 (N_47094,N_35166,N_32140);
or U47095 (N_47095,N_38364,N_39254);
and U47096 (N_47096,N_30320,N_37035);
or U47097 (N_47097,N_38872,N_35920);
or U47098 (N_47098,N_39588,N_36778);
nor U47099 (N_47099,N_33902,N_37519);
xor U47100 (N_47100,N_39079,N_32399);
xnor U47101 (N_47101,N_38922,N_31762);
nor U47102 (N_47102,N_32443,N_37535);
or U47103 (N_47103,N_36142,N_39699);
nor U47104 (N_47104,N_36996,N_36768);
nor U47105 (N_47105,N_38653,N_31267);
or U47106 (N_47106,N_32012,N_36697);
and U47107 (N_47107,N_33721,N_34809);
nand U47108 (N_47108,N_37719,N_39712);
xor U47109 (N_47109,N_35917,N_37393);
nand U47110 (N_47110,N_32986,N_32106);
xor U47111 (N_47111,N_34751,N_39615);
nand U47112 (N_47112,N_36734,N_39066);
and U47113 (N_47113,N_35926,N_33115);
and U47114 (N_47114,N_36266,N_35411);
nor U47115 (N_47115,N_31119,N_35063);
or U47116 (N_47116,N_35238,N_35996);
and U47117 (N_47117,N_39576,N_31012);
and U47118 (N_47118,N_32490,N_33778);
and U47119 (N_47119,N_33778,N_30529);
xor U47120 (N_47120,N_35055,N_34781);
or U47121 (N_47121,N_39858,N_38389);
or U47122 (N_47122,N_37423,N_35090);
or U47123 (N_47123,N_32998,N_36832);
xor U47124 (N_47124,N_30606,N_37200);
nor U47125 (N_47125,N_30745,N_35176);
and U47126 (N_47126,N_35927,N_30160);
xnor U47127 (N_47127,N_30604,N_33323);
nand U47128 (N_47128,N_34659,N_30711);
nand U47129 (N_47129,N_37943,N_39701);
nand U47130 (N_47130,N_38538,N_39706);
and U47131 (N_47131,N_35848,N_34398);
nor U47132 (N_47132,N_38640,N_35252);
nor U47133 (N_47133,N_36029,N_31208);
nor U47134 (N_47134,N_30638,N_34296);
and U47135 (N_47135,N_31833,N_38319);
and U47136 (N_47136,N_38413,N_31617);
nor U47137 (N_47137,N_30596,N_34657);
or U47138 (N_47138,N_36461,N_36341);
or U47139 (N_47139,N_32103,N_35264);
nor U47140 (N_47140,N_37191,N_32945);
xnor U47141 (N_47141,N_36617,N_39069);
or U47142 (N_47142,N_35412,N_33644);
or U47143 (N_47143,N_38359,N_38382);
nor U47144 (N_47144,N_37877,N_39868);
xor U47145 (N_47145,N_32669,N_32468);
and U47146 (N_47146,N_38798,N_36789);
nand U47147 (N_47147,N_33563,N_32658);
or U47148 (N_47148,N_39945,N_38673);
or U47149 (N_47149,N_39390,N_36815);
or U47150 (N_47150,N_30399,N_35580);
nor U47151 (N_47151,N_38948,N_32593);
nor U47152 (N_47152,N_36463,N_35935);
and U47153 (N_47153,N_36868,N_32944);
and U47154 (N_47154,N_30481,N_34607);
nor U47155 (N_47155,N_34730,N_33611);
xor U47156 (N_47156,N_37764,N_37804);
or U47157 (N_47157,N_37287,N_36323);
and U47158 (N_47158,N_39905,N_37204);
xor U47159 (N_47159,N_33286,N_39828);
and U47160 (N_47160,N_34058,N_30198);
nand U47161 (N_47161,N_37110,N_33810);
and U47162 (N_47162,N_37026,N_37476);
nor U47163 (N_47163,N_39745,N_33740);
nand U47164 (N_47164,N_33039,N_30084);
or U47165 (N_47165,N_32376,N_36587);
nor U47166 (N_47166,N_39387,N_39262);
and U47167 (N_47167,N_38683,N_34372);
and U47168 (N_47168,N_31157,N_31138);
nor U47169 (N_47169,N_36243,N_30729);
and U47170 (N_47170,N_32436,N_31950);
nor U47171 (N_47171,N_32996,N_33389);
nand U47172 (N_47172,N_33894,N_34216);
or U47173 (N_47173,N_35023,N_30012);
nand U47174 (N_47174,N_39811,N_39123);
nand U47175 (N_47175,N_34574,N_39253);
nor U47176 (N_47176,N_33742,N_31137);
or U47177 (N_47177,N_34235,N_37508);
nor U47178 (N_47178,N_37022,N_36801);
nor U47179 (N_47179,N_32650,N_32404);
and U47180 (N_47180,N_30598,N_39222);
nand U47181 (N_47181,N_39862,N_36831);
and U47182 (N_47182,N_33270,N_31643);
nand U47183 (N_47183,N_30502,N_32730);
nand U47184 (N_47184,N_36677,N_39834);
and U47185 (N_47185,N_30878,N_33685);
nor U47186 (N_47186,N_30847,N_32340);
nor U47187 (N_47187,N_30981,N_37267);
and U47188 (N_47188,N_33088,N_31345);
nand U47189 (N_47189,N_36767,N_38854);
and U47190 (N_47190,N_37988,N_37187);
nor U47191 (N_47191,N_39538,N_38938);
and U47192 (N_47192,N_33051,N_38824);
nor U47193 (N_47193,N_30517,N_34723);
nand U47194 (N_47194,N_38981,N_36504);
and U47195 (N_47195,N_34721,N_38635);
nand U47196 (N_47196,N_36051,N_30177);
xnor U47197 (N_47197,N_33633,N_34095);
and U47198 (N_47198,N_35750,N_37450);
and U47199 (N_47199,N_37026,N_36659);
or U47200 (N_47200,N_34756,N_38696);
or U47201 (N_47201,N_30496,N_31772);
nand U47202 (N_47202,N_38767,N_39773);
nand U47203 (N_47203,N_33013,N_36056);
nand U47204 (N_47204,N_32865,N_32822);
and U47205 (N_47205,N_39424,N_30291);
nand U47206 (N_47206,N_35290,N_33104);
nand U47207 (N_47207,N_30681,N_36762);
nor U47208 (N_47208,N_31157,N_31662);
nor U47209 (N_47209,N_35317,N_37176);
and U47210 (N_47210,N_35996,N_36586);
nand U47211 (N_47211,N_30566,N_32123);
nand U47212 (N_47212,N_32232,N_31304);
or U47213 (N_47213,N_33245,N_37930);
nor U47214 (N_47214,N_39339,N_33721);
nor U47215 (N_47215,N_37714,N_38938);
xnor U47216 (N_47216,N_34908,N_30394);
nand U47217 (N_47217,N_35646,N_36064);
nor U47218 (N_47218,N_31832,N_35436);
xor U47219 (N_47219,N_39993,N_36735);
nand U47220 (N_47220,N_39230,N_30695);
xnor U47221 (N_47221,N_37147,N_34763);
xor U47222 (N_47222,N_31844,N_36834);
nand U47223 (N_47223,N_38526,N_36749);
or U47224 (N_47224,N_35218,N_37822);
xnor U47225 (N_47225,N_35369,N_34551);
nand U47226 (N_47226,N_30343,N_39357);
nor U47227 (N_47227,N_35919,N_31338);
or U47228 (N_47228,N_38548,N_34117);
xnor U47229 (N_47229,N_36339,N_32205);
or U47230 (N_47230,N_35142,N_38023);
or U47231 (N_47231,N_35570,N_31129);
xnor U47232 (N_47232,N_30455,N_38057);
nor U47233 (N_47233,N_32684,N_33706);
xnor U47234 (N_47234,N_39698,N_34113);
or U47235 (N_47235,N_32181,N_32545);
nor U47236 (N_47236,N_35273,N_32361);
nor U47237 (N_47237,N_38463,N_38353);
xnor U47238 (N_47238,N_39120,N_37782);
xor U47239 (N_47239,N_32177,N_34103);
nor U47240 (N_47240,N_34600,N_30307);
or U47241 (N_47241,N_36797,N_34079);
nand U47242 (N_47242,N_31481,N_31311);
and U47243 (N_47243,N_36804,N_38383);
nor U47244 (N_47244,N_31649,N_30478);
xnor U47245 (N_47245,N_31235,N_39215);
nor U47246 (N_47246,N_34730,N_34902);
nor U47247 (N_47247,N_37003,N_30148);
xnor U47248 (N_47248,N_38537,N_35591);
nor U47249 (N_47249,N_30370,N_35659);
nor U47250 (N_47250,N_30974,N_33226);
or U47251 (N_47251,N_37258,N_30399);
and U47252 (N_47252,N_39250,N_33011);
nor U47253 (N_47253,N_35324,N_30998);
nor U47254 (N_47254,N_32539,N_32114);
or U47255 (N_47255,N_35774,N_39383);
and U47256 (N_47256,N_32023,N_35785);
or U47257 (N_47257,N_34629,N_37941);
xnor U47258 (N_47258,N_31695,N_32263);
xor U47259 (N_47259,N_34134,N_35799);
and U47260 (N_47260,N_37754,N_36647);
xor U47261 (N_47261,N_36945,N_30082);
nor U47262 (N_47262,N_36251,N_35342);
nor U47263 (N_47263,N_30252,N_33472);
nand U47264 (N_47264,N_37599,N_33350);
xor U47265 (N_47265,N_39109,N_37685);
or U47266 (N_47266,N_33233,N_32573);
xor U47267 (N_47267,N_39124,N_37814);
nand U47268 (N_47268,N_37788,N_33709);
nor U47269 (N_47269,N_36576,N_36514);
xor U47270 (N_47270,N_36134,N_39104);
or U47271 (N_47271,N_38603,N_30667);
nor U47272 (N_47272,N_38063,N_30206);
nor U47273 (N_47273,N_30742,N_39258);
nor U47274 (N_47274,N_38629,N_38868);
or U47275 (N_47275,N_32902,N_37369);
or U47276 (N_47276,N_38797,N_32507);
xor U47277 (N_47277,N_34906,N_32335);
and U47278 (N_47278,N_36747,N_37346);
xnor U47279 (N_47279,N_39914,N_35599);
and U47280 (N_47280,N_35479,N_32733);
or U47281 (N_47281,N_36133,N_36511);
nor U47282 (N_47282,N_39686,N_31360);
nor U47283 (N_47283,N_36054,N_37247);
nor U47284 (N_47284,N_35882,N_32091);
nand U47285 (N_47285,N_36018,N_37994);
and U47286 (N_47286,N_34380,N_32219);
and U47287 (N_47287,N_34123,N_36531);
xor U47288 (N_47288,N_30614,N_31683);
nor U47289 (N_47289,N_38775,N_35552);
and U47290 (N_47290,N_36303,N_38169);
xor U47291 (N_47291,N_39869,N_31480);
nand U47292 (N_47292,N_32090,N_31219);
or U47293 (N_47293,N_39491,N_33214);
nor U47294 (N_47294,N_33013,N_39150);
nor U47295 (N_47295,N_31434,N_32725);
and U47296 (N_47296,N_38929,N_37247);
or U47297 (N_47297,N_30282,N_34693);
xor U47298 (N_47298,N_36174,N_38929);
xor U47299 (N_47299,N_35500,N_37762);
nand U47300 (N_47300,N_36097,N_35211);
xor U47301 (N_47301,N_32972,N_32551);
nor U47302 (N_47302,N_32063,N_37520);
nand U47303 (N_47303,N_36174,N_34684);
xnor U47304 (N_47304,N_32844,N_36270);
nor U47305 (N_47305,N_30442,N_33045);
xor U47306 (N_47306,N_38559,N_30736);
nand U47307 (N_47307,N_35145,N_33227);
nand U47308 (N_47308,N_39994,N_34967);
and U47309 (N_47309,N_39281,N_39378);
nand U47310 (N_47310,N_35148,N_38096);
nand U47311 (N_47311,N_34897,N_32670);
xnor U47312 (N_47312,N_36070,N_34697);
xnor U47313 (N_47313,N_34331,N_37782);
nand U47314 (N_47314,N_39271,N_36678);
or U47315 (N_47315,N_34558,N_32082);
xnor U47316 (N_47316,N_35996,N_32371);
xnor U47317 (N_47317,N_33969,N_38673);
or U47318 (N_47318,N_35591,N_34972);
and U47319 (N_47319,N_31456,N_36376);
nand U47320 (N_47320,N_34223,N_31168);
nand U47321 (N_47321,N_33195,N_35765);
xnor U47322 (N_47322,N_33579,N_37069);
nand U47323 (N_47323,N_37127,N_39622);
xnor U47324 (N_47324,N_35354,N_38318);
and U47325 (N_47325,N_38963,N_38261);
and U47326 (N_47326,N_39926,N_37830);
nand U47327 (N_47327,N_32950,N_39113);
xor U47328 (N_47328,N_34977,N_34146);
xor U47329 (N_47329,N_37717,N_34068);
and U47330 (N_47330,N_39114,N_37446);
or U47331 (N_47331,N_33740,N_31446);
and U47332 (N_47332,N_38670,N_34622);
xnor U47333 (N_47333,N_32762,N_35467);
xor U47334 (N_47334,N_31968,N_34222);
and U47335 (N_47335,N_38402,N_39566);
nand U47336 (N_47336,N_36224,N_34583);
nand U47337 (N_47337,N_34137,N_33804);
and U47338 (N_47338,N_39146,N_37219);
and U47339 (N_47339,N_37213,N_33761);
xnor U47340 (N_47340,N_37317,N_36683);
nand U47341 (N_47341,N_35880,N_37518);
nand U47342 (N_47342,N_31230,N_33492);
or U47343 (N_47343,N_36966,N_39454);
xnor U47344 (N_47344,N_31275,N_35401);
nand U47345 (N_47345,N_30453,N_31302);
nor U47346 (N_47346,N_35178,N_33758);
and U47347 (N_47347,N_32290,N_39111);
xor U47348 (N_47348,N_32431,N_35628);
nor U47349 (N_47349,N_35665,N_35567);
nor U47350 (N_47350,N_31235,N_35148);
nor U47351 (N_47351,N_38040,N_34329);
nor U47352 (N_47352,N_33844,N_31139);
nand U47353 (N_47353,N_34957,N_39237);
xnor U47354 (N_47354,N_36768,N_30151);
xnor U47355 (N_47355,N_34154,N_35989);
nand U47356 (N_47356,N_34307,N_33213);
xor U47357 (N_47357,N_30385,N_31481);
nor U47358 (N_47358,N_32196,N_38097);
xor U47359 (N_47359,N_35569,N_37284);
nand U47360 (N_47360,N_30434,N_33294);
and U47361 (N_47361,N_34917,N_37218);
xnor U47362 (N_47362,N_34283,N_33725);
and U47363 (N_47363,N_37015,N_31193);
nor U47364 (N_47364,N_39659,N_33775);
and U47365 (N_47365,N_34750,N_39939);
nor U47366 (N_47366,N_31439,N_36134);
or U47367 (N_47367,N_35816,N_31839);
and U47368 (N_47368,N_33499,N_32327);
nor U47369 (N_47369,N_39395,N_36648);
nor U47370 (N_47370,N_34584,N_32912);
nand U47371 (N_47371,N_34803,N_36644);
or U47372 (N_47372,N_32435,N_30382);
and U47373 (N_47373,N_36301,N_37989);
or U47374 (N_47374,N_31396,N_30145);
and U47375 (N_47375,N_31641,N_35198);
nand U47376 (N_47376,N_34979,N_37652);
nor U47377 (N_47377,N_36905,N_32254);
nor U47378 (N_47378,N_31610,N_32801);
or U47379 (N_47379,N_38319,N_37515);
or U47380 (N_47380,N_39993,N_30187);
xor U47381 (N_47381,N_39812,N_30760);
xnor U47382 (N_47382,N_39100,N_36925);
nor U47383 (N_47383,N_35210,N_32649);
xor U47384 (N_47384,N_36277,N_38134);
nand U47385 (N_47385,N_35652,N_37601);
or U47386 (N_47386,N_38562,N_30318);
nor U47387 (N_47387,N_37104,N_35058);
or U47388 (N_47388,N_36757,N_37224);
nand U47389 (N_47389,N_36899,N_33541);
or U47390 (N_47390,N_32895,N_32466);
and U47391 (N_47391,N_32012,N_36032);
xor U47392 (N_47392,N_37145,N_39863);
nor U47393 (N_47393,N_39074,N_39188);
xor U47394 (N_47394,N_37534,N_32938);
and U47395 (N_47395,N_30399,N_38402);
or U47396 (N_47396,N_34165,N_32364);
xnor U47397 (N_47397,N_31777,N_31397);
or U47398 (N_47398,N_30459,N_33194);
xnor U47399 (N_47399,N_36191,N_38751);
and U47400 (N_47400,N_31269,N_34651);
nand U47401 (N_47401,N_36028,N_38098);
nor U47402 (N_47402,N_38428,N_31367);
and U47403 (N_47403,N_35523,N_31996);
and U47404 (N_47404,N_36588,N_38047);
nand U47405 (N_47405,N_31903,N_37908);
nor U47406 (N_47406,N_37146,N_36754);
or U47407 (N_47407,N_35494,N_39893);
and U47408 (N_47408,N_34095,N_37643);
or U47409 (N_47409,N_36233,N_38800);
xnor U47410 (N_47410,N_38583,N_38375);
and U47411 (N_47411,N_33595,N_36487);
nand U47412 (N_47412,N_35923,N_34774);
nand U47413 (N_47413,N_38469,N_33706);
nand U47414 (N_47414,N_35264,N_31259);
and U47415 (N_47415,N_32768,N_36921);
nor U47416 (N_47416,N_36744,N_37292);
nand U47417 (N_47417,N_39865,N_39132);
nand U47418 (N_47418,N_36866,N_39382);
nand U47419 (N_47419,N_32722,N_31097);
and U47420 (N_47420,N_36475,N_39693);
xor U47421 (N_47421,N_30721,N_38922);
and U47422 (N_47422,N_38301,N_39577);
xor U47423 (N_47423,N_34664,N_38013);
or U47424 (N_47424,N_39585,N_36343);
and U47425 (N_47425,N_37108,N_37179);
and U47426 (N_47426,N_30695,N_38633);
and U47427 (N_47427,N_34182,N_36963);
nor U47428 (N_47428,N_30350,N_30270);
or U47429 (N_47429,N_32017,N_37158);
and U47430 (N_47430,N_30736,N_36934);
and U47431 (N_47431,N_32237,N_32552);
or U47432 (N_47432,N_30817,N_36069);
and U47433 (N_47433,N_34141,N_30333);
xnor U47434 (N_47434,N_35426,N_33227);
xor U47435 (N_47435,N_37135,N_36105);
and U47436 (N_47436,N_36994,N_35853);
nor U47437 (N_47437,N_30125,N_30767);
or U47438 (N_47438,N_37457,N_33217);
or U47439 (N_47439,N_36550,N_36332);
nor U47440 (N_47440,N_34377,N_31767);
or U47441 (N_47441,N_38907,N_31922);
or U47442 (N_47442,N_37839,N_30635);
nor U47443 (N_47443,N_37841,N_30408);
xnor U47444 (N_47444,N_30491,N_33130);
xnor U47445 (N_47445,N_37268,N_38862);
or U47446 (N_47446,N_37435,N_31323);
or U47447 (N_47447,N_35905,N_31437);
or U47448 (N_47448,N_38884,N_30342);
and U47449 (N_47449,N_34952,N_33698);
xor U47450 (N_47450,N_33572,N_31610);
xor U47451 (N_47451,N_30595,N_39856);
nor U47452 (N_47452,N_38699,N_30559);
or U47453 (N_47453,N_32156,N_35933);
or U47454 (N_47454,N_36436,N_31491);
or U47455 (N_47455,N_38037,N_33524);
or U47456 (N_47456,N_39566,N_39563);
nand U47457 (N_47457,N_36537,N_32810);
xor U47458 (N_47458,N_31925,N_31840);
nand U47459 (N_47459,N_30552,N_38516);
nor U47460 (N_47460,N_36613,N_31840);
nor U47461 (N_47461,N_38950,N_30358);
and U47462 (N_47462,N_36370,N_35343);
and U47463 (N_47463,N_33043,N_30366);
xnor U47464 (N_47464,N_30689,N_31262);
and U47465 (N_47465,N_30402,N_33509);
nor U47466 (N_47466,N_38796,N_33074);
nor U47467 (N_47467,N_35404,N_36715);
nand U47468 (N_47468,N_32338,N_30944);
or U47469 (N_47469,N_32040,N_34138);
nor U47470 (N_47470,N_38732,N_31863);
nand U47471 (N_47471,N_31991,N_35986);
and U47472 (N_47472,N_37399,N_36336);
or U47473 (N_47473,N_32901,N_35671);
nand U47474 (N_47474,N_38898,N_39385);
xnor U47475 (N_47475,N_37218,N_34824);
nand U47476 (N_47476,N_39515,N_33164);
or U47477 (N_47477,N_32981,N_31522);
and U47478 (N_47478,N_36883,N_39438);
and U47479 (N_47479,N_31882,N_35620);
and U47480 (N_47480,N_31802,N_39808);
or U47481 (N_47481,N_35635,N_34160);
nand U47482 (N_47482,N_35483,N_34059);
xnor U47483 (N_47483,N_39183,N_34262);
xnor U47484 (N_47484,N_30829,N_38690);
nand U47485 (N_47485,N_38695,N_35412);
and U47486 (N_47486,N_39483,N_30108);
and U47487 (N_47487,N_35443,N_39897);
xor U47488 (N_47488,N_31857,N_31855);
nand U47489 (N_47489,N_30582,N_31588);
and U47490 (N_47490,N_36201,N_37820);
nor U47491 (N_47491,N_36822,N_36403);
nor U47492 (N_47492,N_37604,N_32982);
and U47493 (N_47493,N_37719,N_30625);
and U47494 (N_47494,N_37029,N_31760);
and U47495 (N_47495,N_32651,N_39713);
or U47496 (N_47496,N_36837,N_30122);
or U47497 (N_47497,N_38614,N_39307);
xor U47498 (N_47498,N_31944,N_36040);
nor U47499 (N_47499,N_31891,N_36364);
or U47500 (N_47500,N_37288,N_33167);
xor U47501 (N_47501,N_38879,N_39367);
xor U47502 (N_47502,N_30262,N_37464);
nand U47503 (N_47503,N_36619,N_36984);
and U47504 (N_47504,N_32768,N_36618);
nand U47505 (N_47505,N_31863,N_33776);
and U47506 (N_47506,N_31248,N_34406);
xnor U47507 (N_47507,N_38193,N_32215);
and U47508 (N_47508,N_30727,N_30694);
nand U47509 (N_47509,N_31687,N_31546);
xnor U47510 (N_47510,N_35265,N_39548);
and U47511 (N_47511,N_33681,N_38824);
xnor U47512 (N_47512,N_37864,N_30712);
xnor U47513 (N_47513,N_35071,N_35201);
and U47514 (N_47514,N_32570,N_35065);
or U47515 (N_47515,N_38479,N_38916);
and U47516 (N_47516,N_34059,N_38243);
and U47517 (N_47517,N_31657,N_32181);
nand U47518 (N_47518,N_34651,N_37399);
nand U47519 (N_47519,N_38525,N_34942);
xor U47520 (N_47520,N_37489,N_35868);
nor U47521 (N_47521,N_36455,N_33485);
nand U47522 (N_47522,N_38138,N_31653);
or U47523 (N_47523,N_36613,N_31763);
nor U47524 (N_47524,N_31182,N_31391);
nand U47525 (N_47525,N_32626,N_31894);
or U47526 (N_47526,N_37845,N_37279);
xnor U47527 (N_47527,N_30965,N_30032);
and U47528 (N_47528,N_31881,N_34876);
nor U47529 (N_47529,N_35568,N_32110);
or U47530 (N_47530,N_35147,N_38961);
nand U47531 (N_47531,N_30850,N_37017);
and U47532 (N_47532,N_38601,N_38306);
nand U47533 (N_47533,N_31537,N_36454);
nand U47534 (N_47534,N_34633,N_31230);
nor U47535 (N_47535,N_39525,N_31392);
nand U47536 (N_47536,N_39234,N_38050);
and U47537 (N_47537,N_35981,N_38524);
nand U47538 (N_47538,N_31763,N_37246);
nand U47539 (N_47539,N_32615,N_32112);
or U47540 (N_47540,N_37997,N_33596);
and U47541 (N_47541,N_39127,N_36054);
nand U47542 (N_47542,N_36486,N_37424);
or U47543 (N_47543,N_33625,N_39383);
nor U47544 (N_47544,N_33548,N_37345);
nor U47545 (N_47545,N_39672,N_38648);
or U47546 (N_47546,N_34779,N_37130);
xnor U47547 (N_47547,N_37247,N_32693);
xor U47548 (N_47548,N_34201,N_34374);
or U47549 (N_47549,N_39869,N_33401);
nor U47550 (N_47550,N_36085,N_33296);
and U47551 (N_47551,N_39357,N_31048);
nand U47552 (N_47552,N_38716,N_34067);
nor U47553 (N_47553,N_32686,N_31921);
nor U47554 (N_47554,N_35754,N_34092);
or U47555 (N_47555,N_35441,N_37292);
nand U47556 (N_47556,N_34405,N_39280);
or U47557 (N_47557,N_36759,N_34826);
nand U47558 (N_47558,N_35085,N_31690);
and U47559 (N_47559,N_39118,N_33709);
nand U47560 (N_47560,N_31151,N_36665);
and U47561 (N_47561,N_30545,N_36144);
xor U47562 (N_47562,N_35968,N_31335);
xnor U47563 (N_47563,N_30263,N_33392);
xnor U47564 (N_47564,N_38025,N_30098);
or U47565 (N_47565,N_38490,N_34973);
xor U47566 (N_47566,N_33048,N_39652);
nor U47567 (N_47567,N_33249,N_35204);
xnor U47568 (N_47568,N_33369,N_34304);
nand U47569 (N_47569,N_37484,N_38958);
xor U47570 (N_47570,N_30957,N_39086);
xnor U47571 (N_47571,N_30068,N_33916);
and U47572 (N_47572,N_39103,N_34227);
and U47573 (N_47573,N_38134,N_33214);
or U47574 (N_47574,N_30580,N_39934);
and U47575 (N_47575,N_31887,N_30475);
nor U47576 (N_47576,N_33845,N_34008);
nor U47577 (N_47577,N_39621,N_30724);
xor U47578 (N_47578,N_31173,N_30339);
nor U47579 (N_47579,N_31447,N_37047);
nand U47580 (N_47580,N_38750,N_30204);
or U47581 (N_47581,N_31790,N_33034);
nand U47582 (N_47582,N_38434,N_33244);
xor U47583 (N_47583,N_34508,N_32491);
and U47584 (N_47584,N_31825,N_39343);
nor U47585 (N_47585,N_34993,N_34647);
nor U47586 (N_47586,N_34853,N_35722);
nor U47587 (N_47587,N_37888,N_36764);
nand U47588 (N_47588,N_39543,N_39391);
nor U47589 (N_47589,N_32977,N_38374);
or U47590 (N_47590,N_30760,N_39328);
nor U47591 (N_47591,N_38162,N_30696);
xor U47592 (N_47592,N_39994,N_30896);
xnor U47593 (N_47593,N_38090,N_36615);
or U47594 (N_47594,N_34929,N_36499);
nor U47595 (N_47595,N_34561,N_38200);
nor U47596 (N_47596,N_34274,N_36850);
nand U47597 (N_47597,N_32402,N_35885);
or U47598 (N_47598,N_38989,N_33821);
or U47599 (N_47599,N_38789,N_34601);
nor U47600 (N_47600,N_34127,N_30348);
and U47601 (N_47601,N_31352,N_39868);
nor U47602 (N_47602,N_32672,N_33126);
or U47603 (N_47603,N_32392,N_31969);
nor U47604 (N_47604,N_33578,N_32549);
xor U47605 (N_47605,N_30432,N_39075);
or U47606 (N_47606,N_38821,N_34565);
and U47607 (N_47607,N_30561,N_35722);
nor U47608 (N_47608,N_39050,N_34707);
and U47609 (N_47609,N_36289,N_39229);
nand U47610 (N_47610,N_38269,N_35087);
and U47611 (N_47611,N_36696,N_38479);
and U47612 (N_47612,N_36318,N_36281);
and U47613 (N_47613,N_35089,N_30844);
nand U47614 (N_47614,N_32316,N_35086);
nand U47615 (N_47615,N_39504,N_31866);
xnor U47616 (N_47616,N_36139,N_32614);
or U47617 (N_47617,N_35501,N_37036);
and U47618 (N_47618,N_31982,N_34988);
and U47619 (N_47619,N_33949,N_30217);
or U47620 (N_47620,N_35258,N_36603);
and U47621 (N_47621,N_32427,N_39764);
xnor U47622 (N_47622,N_30020,N_35690);
or U47623 (N_47623,N_32605,N_39299);
nor U47624 (N_47624,N_38420,N_35914);
xor U47625 (N_47625,N_39334,N_38741);
nand U47626 (N_47626,N_38114,N_31372);
nand U47627 (N_47627,N_38320,N_35960);
nor U47628 (N_47628,N_34234,N_34642);
xnor U47629 (N_47629,N_35855,N_32483);
or U47630 (N_47630,N_36277,N_34304);
or U47631 (N_47631,N_34551,N_37274);
nor U47632 (N_47632,N_36247,N_39816);
nand U47633 (N_47633,N_32542,N_39749);
nor U47634 (N_47634,N_32445,N_37669);
and U47635 (N_47635,N_37438,N_36056);
and U47636 (N_47636,N_37849,N_36407);
or U47637 (N_47637,N_35100,N_33203);
and U47638 (N_47638,N_35323,N_35105);
or U47639 (N_47639,N_32362,N_37547);
nand U47640 (N_47640,N_37936,N_39551);
nand U47641 (N_47641,N_35708,N_35573);
or U47642 (N_47642,N_36375,N_38901);
xnor U47643 (N_47643,N_36316,N_32110);
or U47644 (N_47644,N_30352,N_32834);
nor U47645 (N_47645,N_32372,N_32861);
xnor U47646 (N_47646,N_35495,N_34849);
xor U47647 (N_47647,N_32642,N_36413);
nand U47648 (N_47648,N_31790,N_38601);
and U47649 (N_47649,N_31903,N_34940);
nor U47650 (N_47650,N_38600,N_38890);
nand U47651 (N_47651,N_39293,N_34375);
or U47652 (N_47652,N_31728,N_34331);
and U47653 (N_47653,N_34186,N_35724);
nand U47654 (N_47654,N_35488,N_30956);
or U47655 (N_47655,N_32232,N_34746);
xor U47656 (N_47656,N_32087,N_39149);
nor U47657 (N_47657,N_30466,N_30651);
nand U47658 (N_47658,N_39013,N_32741);
and U47659 (N_47659,N_32972,N_32341);
or U47660 (N_47660,N_39650,N_39671);
xor U47661 (N_47661,N_30784,N_38900);
or U47662 (N_47662,N_38937,N_38023);
xnor U47663 (N_47663,N_39710,N_32421);
and U47664 (N_47664,N_35246,N_30472);
and U47665 (N_47665,N_38402,N_35477);
nand U47666 (N_47666,N_38972,N_33831);
xor U47667 (N_47667,N_31006,N_33855);
nand U47668 (N_47668,N_33521,N_39687);
nand U47669 (N_47669,N_37249,N_39466);
xor U47670 (N_47670,N_32517,N_32142);
xor U47671 (N_47671,N_37526,N_34210);
and U47672 (N_47672,N_37233,N_31312);
nand U47673 (N_47673,N_32597,N_30391);
and U47674 (N_47674,N_34775,N_30386);
and U47675 (N_47675,N_30523,N_33238);
nor U47676 (N_47676,N_35130,N_30747);
nor U47677 (N_47677,N_36586,N_32393);
nand U47678 (N_47678,N_31407,N_30964);
xnor U47679 (N_47679,N_37728,N_39568);
nor U47680 (N_47680,N_30050,N_39940);
and U47681 (N_47681,N_31880,N_35701);
or U47682 (N_47682,N_33469,N_34230);
nor U47683 (N_47683,N_39912,N_39446);
and U47684 (N_47684,N_30080,N_35708);
and U47685 (N_47685,N_35511,N_35505);
xnor U47686 (N_47686,N_35398,N_30811);
nor U47687 (N_47687,N_30181,N_30013);
xnor U47688 (N_47688,N_39053,N_33544);
nor U47689 (N_47689,N_33838,N_30994);
nand U47690 (N_47690,N_35497,N_39746);
and U47691 (N_47691,N_37372,N_38779);
and U47692 (N_47692,N_37427,N_39693);
nor U47693 (N_47693,N_34594,N_36284);
xnor U47694 (N_47694,N_35045,N_37652);
nor U47695 (N_47695,N_35436,N_35223);
xnor U47696 (N_47696,N_30271,N_39133);
xnor U47697 (N_47697,N_39628,N_33039);
nand U47698 (N_47698,N_34772,N_39767);
nand U47699 (N_47699,N_36822,N_31114);
xnor U47700 (N_47700,N_33113,N_32365);
or U47701 (N_47701,N_34206,N_35437);
nand U47702 (N_47702,N_35007,N_39250);
and U47703 (N_47703,N_32415,N_37583);
xor U47704 (N_47704,N_35666,N_32652);
or U47705 (N_47705,N_39414,N_39406);
or U47706 (N_47706,N_36582,N_31968);
and U47707 (N_47707,N_35490,N_30045);
or U47708 (N_47708,N_34121,N_31084);
xor U47709 (N_47709,N_33419,N_33212);
nand U47710 (N_47710,N_34561,N_33425);
nor U47711 (N_47711,N_36186,N_39120);
nor U47712 (N_47712,N_31785,N_38229);
xnor U47713 (N_47713,N_39294,N_37960);
or U47714 (N_47714,N_30830,N_38589);
nand U47715 (N_47715,N_38216,N_38411);
or U47716 (N_47716,N_30497,N_39642);
nor U47717 (N_47717,N_36673,N_35517);
or U47718 (N_47718,N_32792,N_33814);
or U47719 (N_47719,N_31613,N_38494);
xnor U47720 (N_47720,N_30594,N_30856);
xor U47721 (N_47721,N_37619,N_33585);
nor U47722 (N_47722,N_39525,N_39460);
or U47723 (N_47723,N_37647,N_38176);
nor U47724 (N_47724,N_35986,N_34986);
and U47725 (N_47725,N_34364,N_30253);
or U47726 (N_47726,N_37656,N_30920);
and U47727 (N_47727,N_39765,N_35383);
nor U47728 (N_47728,N_36849,N_36596);
nand U47729 (N_47729,N_37139,N_31314);
xor U47730 (N_47730,N_33364,N_36974);
nor U47731 (N_47731,N_33434,N_31374);
xnor U47732 (N_47732,N_35493,N_34199);
nand U47733 (N_47733,N_32168,N_30464);
xnor U47734 (N_47734,N_30781,N_30505);
or U47735 (N_47735,N_37505,N_35735);
and U47736 (N_47736,N_39616,N_38229);
and U47737 (N_47737,N_31325,N_39745);
xor U47738 (N_47738,N_34392,N_35606);
nor U47739 (N_47739,N_33232,N_32526);
or U47740 (N_47740,N_32821,N_31116);
xor U47741 (N_47741,N_38830,N_34550);
and U47742 (N_47742,N_32125,N_39584);
or U47743 (N_47743,N_34066,N_31937);
xor U47744 (N_47744,N_31471,N_39560);
xnor U47745 (N_47745,N_39419,N_39545);
or U47746 (N_47746,N_36282,N_30956);
xor U47747 (N_47747,N_32459,N_37477);
nand U47748 (N_47748,N_33522,N_34884);
nand U47749 (N_47749,N_39878,N_37926);
xor U47750 (N_47750,N_31461,N_38825);
and U47751 (N_47751,N_38569,N_37768);
or U47752 (N_47752,N_37173,N_30229);
nand U47753 (N_47753,N_32652,N_34481);
nor U47754 (N_47754,N_33715,N_35127);
nand U47755 (N_47755,N_35522,N_36176);
nand U47756 (N_47756,N_32535,N_32144);
nand U47757 (N_47757,N_38884,N_33839);
or U47758 (N_47758,N_37607,N_31535);
or U47759 (N_47759,N_35079,N_30845);
nand U47760 (N_47760,N_32723,N_38541);
xnor U47761 (N_47761,N_37613,N_34488);
nand U47762 (N_47762,N_31866,N_33043);
or U47763 (N_47763,N_34393,N_36872);
nand U47764 (N_47764,N_35611,N_34580);
nand U47765 (N_47765,N_33419,N_33768);
and U47766 (N_47766,N_38776,N_31051);
xor U47767 (N_47767,N_33838,N_35750);
or U47768 (N_47768,N_30292,N_36122);
and U47769 (N_47769,N_39379,N_31779);
nor U47770 (N_47770,N_38222,N_31915);
nand U47771 (N_47771,N_31200,N_30062);
nand U47772 (N_47772,N_34272,N_38989);
nand U47773 (N_47773,N_35272,N_32746);
nand U47774 (N_47774,N_34516,N_32640);
or U47775 (N_47775,N_37265,N_32038);
nor U47776 (N_47776,N_34565,N_36184);
xor U47777 (N_47777,N_33149,N_35873);
nand U47778 (N_47778,N_30602,N_35261);
nor U47779 (N_47779,N_37983,N_37559);
nor U47780 (N_47780,N_35390,N_31540);
xnor U47781 (N_47781,N_39792,N_35814);
xor U47782 (N_47782,N_38255,N_34017);
and U47783 (N_47783,N_31643,N_32133);
or U47784 (N_47784,N_31833,N_36437);
xor U47785 (N_47785,N_30444,N_31053);
nor U47786 (N_47786,N_39085,N_38837);
xor U47787 (N_47787,N_36846,N_35944);
nand U47788 (N_47788,N_34466,N_39759);
nor U47789 (N_47789,N_38891,N_31888);
or U47790 (N_47790,N_33677,N_33657);
or U47791 (N_47791,N_30688,N_39864);
and U47792 (N_47792,N_30364,N_36926);
xnor U47793 (N_47793,N_37712,N_36242);
xor U47794 (N_47794,N_37027,N_39522);
nand U47795 (N_47795,N_33162,N_35187);
nand U47796 (N_47796,N_33706,N_36709);
nor U47797 (N_47797,N_34276,N_31529);
xnor U47798 (N_47798,N_38511,N_30761);
or U47799 (N_47799,N_32857,N_38819);
nand U47800 (N_47800,N_36794,N_38273);
nand U47801 (N_47801,N_35288,N_36651);
xor U47802 (N_47802,N_39791,N_37943);
and U47803 (N_47803,N_32393,N_31244);
nor U47804 (N_47804,N_34255,N_39691);
xnor U47805 (N_47805,N_36717,N_38922);
xor U47806 (N_47806,N_32530,N_33806);
or U47807 (N_47807,N_31432,N_31394);
xnor U47808 (N_47808,N_39916,N_31190);
and U47809 (N_47809,N_31644,N_30074);
xnor U47810 (N_47810,N_34887,N_34096);
xnor U47811 (N_47811,N_30052,N_34921);
and U47812 (N_47812,N_33345,N_31500);
or U47813 (N_47813,N_38903,N_30520);
xor U47814 (N_47814,N_30863,N_37931);
nand U47815 (N_47815,N_37085,N_39402);
and U47816 (N_47816,N_38452,N_34439);
xor U47817 (N_47817,N_32945,N_33074);
xnor U47818 (N_47818,N_39525,N_37296);
nor U47819 (N_47819,N_35409,N_32015);
or U47820 (N_47820,N_31355,N_36395);
or U47821 (N_47821,N_30394,N_36653);
xnor U47822 (N_47822,N_30645,N_38715);
or U47823 (N_47823,N_36885,N_32624);
or U47824 (N_47824,N_30153,N_34789);
xor U47825 (N_47825,N_35783,N_34532);
nand U47826 (N_47826,N_39821,N_37189);
or U47827 (N_47827,N_35451,N_34477);
nor U47828 (N_47828,N_30815,N_33363);
and U47829 (N_47829,N_31107,N_35467);
xnor U47830 (N_47830,N_35005,N_33645);
nand U47831 (N_47831,N_30549,N_31023);
nor U47832 (N_47832,N_32855,N_30955);
nand U47833 (N_47833,N_38003,N_30650);
and U47834 (N_47834,N_37205,N_38339);
nand U47835 (N_47835,N_32959,N_35679);
nor U47836 (N_47836,N_34148,N_31271);
and U47837 (N_47837,N_34978,N_35389);
and U47838 (N_47838,N_30392,N_34081);
nand U47839 (N_47839,N_38412,N_31743);
nor U47840 (N_47840,N_31216,N_31073);
xnor U47841 (N_47841,N_33870,N_34706);
or U47842 (N_47842,N_35764,N_37673);
or U47843 (N_47843,N_34306,N_35868);
nand U47844 (N_47844,N_32206,N_37996);
xor U47845 (N_47845,N_38280,N_36623);
nand U47846 (N_47846,N_32124,N_33033);
nor U47847 (N_47847,N_37794,N_30414);
nand U47848 (N_47848,N_30241,N_39003);
nand U47849 (N_47849,N_38758,N_30849);
and U47850 (N_47850,N_33447,N_38311);
xnor U47851 (N_47851,N_35897,N_34480);
and U47852 (N_47852,N_38164,N_33362);
and U47853 (N_47853,N_39093,N_37818);
nor U47854 (N_47854,N_32638,N_30093);
or U47855 (N_47855,N_37560,N_39914);
or U47856 (N_47856,N_33382,N_34688);
xnor U47857 (N_47857,N_34054,N_38271);
nor U47858 (N_47858,N_31773,N_39265);
or U47859 (N_47859,N_39233,N_36723);
and U47860 (N_47860,N_35208,N_39976);
xor U47861 (N_47861,N_31802,N_32158);
and U47862 (N_47862,N_39593,N_34734);
xor U47863 (N_47863,N_36787,N_35848);
and U47864 (N_47864,N_36533,N_39335);
nor U47865 (N_47865,N_39334,N_32890);
and U47866 (N_47866,N_33751,N_32587);
and U47867 (N_47867,N_33053,N_30045);
and U47868 (N_47868,N_31501,N_39369);
or U47869 (N_47869,N_35343,N_35659);
nor U47870 (N_47870,N_39581,N_33101);
xnor U47871 (N_47871,N_31720,N_33724);
nand U47872 (N_47872,N_35196,N_37956);
or U47873 (N_47873,N_31865,N_33046);
or U47874 (N_47874,N_38593,N_35150);
or U47875 (N_47875,N_33120,N_34170);
xor U47876 (N_47876,N_36987,N_33754);
or U47877 (N_47877,N_37781,N_35933);
or U47878 (N_47878,N_32616,N_34478);
or U47879 (N_47879,N_38611,N_32360);
nor U47880 (N_47880,N_32179,N_34233);
and U47881 (N_47881,N_30710,N_33024);
xor U47882 (N_47882,N_33800,N_30152);
and U47883 (N_47883,N_33019,N_39503);
nand U47884 (N_47884,N_32802,N_34623);
and U47885 (N_47885,N_34507,N_35428);
xor U47886 (N_47886,N_38827,N_33888);
or U47887 (N_47887,N_33849,N_36107);
nand U47888 (N_47888,N_34759,N_30903);
and U47889 (N_47889,N_37101,N_32207);
or U47890 (N_47890,N_33947,N_31272);
nor U47891 (N_47891,N_36236,N_39497);
nand U47892 (N_47892,N_39306,N_34554);
xor U47893 (N_47893,N_38582,N_39878);
xnor U47894 (N_47894,N_30200,N_33632);
or U47895 (N_47895,N_30251,N_39591);
or U47896 (N_47896,N_33012,N_39885);
xor U47897 (N_47897,N_34992,N_32595);
and U47898 (N_47898,N_38057,N_31325);
or U47899 (N_47899,N_36647,N_30399);
or U47900 (N_47900,N_33825,N_31787);
or U47901 (N_47901,N_33108,N_39742);
nand U47902 (N_47902,N_32259,N_32734);
nor U47903 (N_47903,N_35151,N_37714);
nand U47904 (N_47904,N_34369,N_36074);
and U47905 (N_47905,N_36256,N_32418);
nand U47906 (N_47906,N_34100,N_37826);
xor U47907 (N_47907,N_39493,N_38162);
nor U47908 (N_47908,N_36195,N_38533);
nand U47909 (N_47909,N_32978,N_30138);
xnor U47910 (N_47910,N_38739,N_31685);
or U47911 (N_47911,N_39304,N_36238);
xor U47912 (N_47912,N_30309,N_30639);
xor U47913 (N_47913,N_34935,N_38008);
xor U47914 (N_47914,N_39346,N_32342);
and U47915 (N_47915,N_35672,N_37833);
and U47916 (N_47916,N_38077,N_31318);
nor U47917 (N_47917,N_31439,N_31697);
nor U47918 (N_47918,N_31107,N_32472);
or U47919 (N_47919,N_39642,N_30548);
or U47920 (N_47920,N_32411,N_34483);
nand U47921 (N_47921,N_39307,N_37133);
and U47922 (N_47922,N_31891,N_34550);
xor U47923 (N_47923,N_31086,N_33526);
xnor U47924 (N_47924,N_30531,N_36929);
nand U47925 (N_47925,N_34279,N_33614);
or U47926 (N_47926,N_32280,N_34678);
and U47927 (N_47927,N_35768,N_32265);
xnor U47928 (N_47928,N_33665,N_30287);
nor U47929 (N_47929,N_34081,N_36116);
or U47930 (N_47930,N_37661,N_32970);
or U47931 (N_47931,N_36878,N_37541);
nor U47932 (N_47932,N_37544,N_31722);
or U47933 (N_47933,N_39047,N_32316);
and U47934 (N_47934,N_33214,N_34606);
or U47935 (N_47935,N_31683,N_36803);
nand U47936 (N_47936,N_33424,N_30330);
and U47937 (N_47937,N_31397,N_38257);
nor U47938 (N_47938,N_31023,N_39060);
and U47939 (N_47939,N_32343,N_34866);
or U47940 (N_47940,N_30447,N_35777);
nand U47941 (N_47941,N_39928,N_39565);
xnor U47942 (N_47942,N_34086,N_39380);
nand U47943 (N_47943,N_31027,N_38054);
nand U47944 (N_47944,N_33251,N_38959);
nand U47945 (N_47945,N_39091,N_39782);
nand U47946 (N_47946,N_31863,N_32128);
xnor U47947 (N_47947,N_38338,N_35956);
or U47948 (N_47948,N_39638,N_39287);
and U47949 (N_47949,N_35865,N_38028);
nor U47950 (N_47950,N_36875,N_39310);
nand U47951 (N_47951,N_37045,N_37266);
or U47952 (N_47952,N_37540,N_34100);
and U47953 (N_47953,N_34868,N_32904);
nor U47954 (N_47954,N_35116,N_34790);
nand U47955 (N_47955,N_32268,N_33562);
nor U47956 (N_47956,N_38559,N_31265);
nand U47957 (N_47957,N_37484,N_39949);
or U47958 (N_47958,N_37482,N_32631);
nor U47959 (N_47959,N_39741,N_39418);
nand U47960 (N_47960,N_35761,N_31057);
or U47961 (N_47961,N_33516,N_30575);
nand U47962 (N_47962,N_37565,N_36820);
nand U47963 (N_47963,N_35094,N_31117);
or U47964 (N_47964,N_39099,N_31337);
and U47965 (N_47965,N_39943,N_34530);
or U47966 (N_47966,N_37454,N_39870);
and U47967 (N_47967,N_34285,N_39677);
nor U47968 (N_47968,N_35950,N_30677);
or U47969 (N_47969,N_30382,N_35013);
or U47970 (N_47970,N_30959,N_39036);
nand U47971 (N_47971,N_37168,N_31173);
nor U47972 (N_47972,N_32378,N_38508);
nand U47973 (N_47973,N_33062,N_32922);
xnor U47974 (N_47974,N_35472,N_30287);
or U47975 (N_47975,N_31609,N_37842);
xnor U47976 (N_47976,N_35454,N_37550);
xor U47977 (N_47977,N_30927,N_34713);
nand U47978 (N_47978,N_38421,N_35994);
nor U47979 (N_47979,N_32407,N_38973);
and U47980 (N_47980,N_37636,N_37311);
and U47981 (N_47981,N_32132,N_37075);
xor U47982 (N_47982,N_33443,N_35743);
nor U47983 (N_47983,N_33240,N_31068);
and U47984 (N_47984,N_33378,N_30875);
nor U47985 (N_47985,N_31674,N_32326);
xnor U47986 (N_47986,N_38998,N_35782);
or U47987 (N_47987,N_37570,N_39332);
nand U47988 (N_47988,N_39149,N_37436);
or U47989 (N_47989,N_30348,N_36848);
nand U47990 (N_47990,N_38474,N_38101);
nand U47991 (N_47991,N_31589,N_35497);
nand U47992 (N_47992,N_36586,N_38864);
nand U47993 (N_47993,N_37380,N_37843);
nor U47994 (N_47994,N_33669,N_35204);
and U47995 (N_47995,N_33886,N_30932);
nand U47996 (N_47996,N_31896,N_31439);
and U47997 (N_47997,N_31796,N_35819);
nand U47998 (N_47998,N_37968,N_32039);
nand U47999 (N_47999,N_31392,N_37326);
and U48000 (N_48000,N_32501,N_39542);
nand U48001 (N_48001,N_39820,N_37161);
nor U48002 (N_48002,N_32920,N_33304);
xor U48003 (N_48003,N_31649,N_30524);
nand U48004 (N_48004,N_39590,N_30392);
nor U48005 (N_48005,N_30812,N_33390);
and U48006 (N_48006,N_30086,N_30918);
xor U48007 (N_48007,N_30574,N_30343);
and U48008 (N_48008,N_33648,N_34811);
xor U48009 (N_48009,N_33668,N_38285);
or U48010 (N_48010,N_37079,N_32444);
nand U48011 (N_48011,N_32416,N_38350);
xor U48012 (N_48012,N_32461,N_30930);
nor U48013 (N_48013,N_30921,N_38723);
nor U48014 (N_48014,N_31850,N_38360);
or U48015 (N_48015,N_37582,N_30377);
and U48016 (N_48016,N_32570,N_30888);
nand U48017 (N_48017,N_37396,N_38123);
or U48018 (N_48018,N_34669,N_33914);
or U48019 (N_48019,N_38457,N_31338);
nand U48020 (N_48020,N_35679,N_30524);
nand U48021 (N_48021,N_38918,N_37434);
xor U48022 (N_48022,N_39860,N_35370);
or U48023 (N_48023,N_35429,N_31438);
nor U48024 (N_48024,N_30702,N_35095);
nor U48025 (N_48025,N_31510,N_32515);
nand U48026 (N_48026,N_38998,N_38839);
nand U48027 (N_48027,N_37190,N_38956);
and U48028 (N_48028,N_35137,N_37080);
nor U48029 (N_48029,N_34596,N_35945);
and U48030 (N_48030,N_38365,N_30367);
and U48031 (N_48031,N_34785,N_31867);
nand U48032 (N_48032,N_33678,N_30466);
or U48033 (N_48033,N_30434,N_32229);
xnor U48034 (N_48034,N_38414,N_39343);
xnor U48035 (N_48035,N_37991,N_33591);
nand U48036 (N_48036,N_39181,N_36240);
or U48037 (N_48037,N_39937,N_35673);
xor U48038 (N_48038,N_37609,N_30652);
nand U48039 (N_48039,N_36261,N_33020);
nor U48040 (N_48040,N_35872,N_34921);
xor U48041 (N_48041,N_36169,N_38562);
and U48042 (N_48042,N_34168,N_34601);
nand U48043 (N_48043,N_34220,N_38067);
or U48044 (N_48044,N_31394,N_39922);
nand U48045 (N_48045,N_35999,N_39048);
nand U48046 (N_48046,N_36949,N_37779);
nor U48047 (N_48047,N_39747,N_34431);
nand U48048 (N_48048,N_36127,N_30710);
xor U48049 (N_48049,N_37153,N_32900);
and U48050 (N_48050,N_33054,N_31953);
and U48051 (N_48051,N_35293,N_37833);
nand U48052 (N_48052,N_34345,N_35565);
nand U48053 (N_48053,N_33279,N_30459);
nand U48054 (N_48054,N_32688,N_33990);
or U48055 (N_48055,N_34033,N_31893);
nand U48056 (N_48056,N_30740,N_32521);
nand U48057 (N_48057,N_33835,N_37778);
nor U48058 (N_48058,N_38287,N_38872);
and U48059 (N_48059,N_37269,N_35023);
nand U48060 (N_48060,N_35761,N_32101);
xor U48061 (N_48061,N_36705,N_32812);
xor U48062 (N_48062,N_39327,N_34096);
or U48063 (N_48063,N_34815,N_34645);
and U48064 (N_48064,N_32276,N_31892);
nor U48065 (N_48065,N_30561,N_38208);
and U48066 (N_48066,N_36591,N_31241);
nand U48067 (N_48067,N_35986,N_34338);
or U48068 (N_48068,N_31176,N_30855);
or U48069 (N_48069,N_33303,N_37113);
xor U48070 (N_48070,N_38320,N_35463);
xor U48071 (N_48071,N_39533,N_38876);
or U48072 (N_48072,N_39554,N_38611);
xor U48073 (N_48073,N_35207,N_33215);
xnor U48074 (N_48074,N_38192,N_37547);
and U48075 (N_48075,N_33004,N_34683);
or U48076 (N_48076,N_30553,N_39997);
xnor U48077 (N_48077,N_36062,N_32532);
xnor U48078 (N_48078,N_33920,N_33432);
xnor U48079 (N_48079,N_32905,N_31487);
or U48080 (N_48080,N_37606,N_31838);
xor U48081 (N_48081,N_35376,N_35861);
nor U48082 (N_48082,N_37223,N_33739);
nor U48083 (N_48083,N_31901,N_37730);
or U48084 (N_48084,N_39302,N_34318);
xnor U48085 (N_48085,N_38938,N_34290);
and U48086 (N_48086,N_37578,N_36087);
and U48087 (N_48087,N_38388,N_31887);
or U48088 (N_48088,N_33042,N_30078);
or U48089 (N_48089,N_34315,N_38544);
xnor U48090 (N_48090,N_30783,N_36242);
and U48091 (N_48091,N_37974,N_35053);
and U48092 (N_48092,N_34057,N_33613);
and U48093 (N_48093,N_32418,N_30365);
or U48094 (N_48094,N_37668,N_37909);
nor U48095 (N_48095,N_33802,N_38267);
nor U48096 (N_48096,N_38752,N_39736);
and U48097 (N_48097,N_31499,N_32183);
or U48098 (N_48098,N_37556,N_32522);
nand U48099 (N_48099,N_31939,N_31693);
or U48100 (N_48100,N_31278,N_39666);
and U48101 (N_48101,N_38583,N_37540);
and U48102 (N_48102,N_35157,N_31806);
or U48103 (N_48103,N_35745,N_31299);
xor U48104 (N_48104,N_39040,N_36695);
nor U48105 (N_48105,N_32646,N_35292);
nor U48106 (N_48106,N_35461,N_30890);
or U48107 (N_48107,N_37290,N_30180);
nor U48108 (N_48108,N_34978,N_35385);
nor U48109 (N_48109,N_30183,N_30487);
nand U48110 (N_48110,N_32413,N_31984);
and U48111 (N_48111,N_32038,N_38969);
and U48112 (N_48112,N_34133,N_39872);
nand U48113 (N_48113,N_33176,N_38202);
xnor U48114 (N_48114,N_32928,N_33330);
nand U48115 (N_48115,N_36937,N_31859);
and U48116 (N_48116,N_36189,N_34340);
and U48117 (N_48117,N_36290,N_31416);
nor U48118 (N_48118,N_36190,N_36822);
and U48119 (N_48119,N_36317,N_34935);
and U48120 (N_48120,N_35196,N_35193);
xnor U48121 (N_48121,N_34942,N_33340);
nor U48122 (N_48122,N_34950,N_32848);
nor U48123 (N_48123,N_32493,N_32863);
nor U48124 (N_48124,N_31279,N_33782);
nand U48125 (N_48125,N_36268,N_34615);
nor U48126 (N_48126,N_32595,N_30081);
nand U48127 (N_48127,N_32573,N_31936);
and U48128 (N_48128,N_37358,N_31891);
and U48129 (N_48129,N_38673,N_30999);
nand U48130 (N_48130,N_35720,N_34658);
xnor U48131 (N_48131,N_37336,N_30043);
or U48132 (N_48132,N_39210,N_32958);
xnor U48133 (N_48133,N_31635,N_32489);
nand U48134 (N_48134,N_33267,N_31623);
nand U48135 (N_48135,N_33276,N_37651);
xor U48136 (N_48136,N_35666,N_36906);
nand U48137 (N_48137,N_33677,N_38661);
and U48138 (N_48138,N_39943,N_36226);
and U48139 (N_48139,N_36004,N_30084);
or U48140 (N_48140,N_36358,N_32535);
or U48141 (N_48141,N_30450,N_33576);
and U48142 (N_48142,N_32145,N_37313);
or U48143 (N_48143,N_38561,N_34396);
nor U48144 (N_48144,N_34172,N_36441);
and U48145 (N_48145,N_31679,N_37553);
or U48146 (N_48146,N_38771,N_34991);
xor U48147 (N_48147,N_35472,N_36666);
or U48148 (N_48148,N_36380,N_36851);
and U48149 (N_48149,N_38370,N_38599);
or U48150 (N_48150,N_39885,N_34650);
nand U48151 (N_48151,N_31730,N_38091);
or U48152 (N_48152,N_32039,N_34402);
and U48153 (N_48153,N_31535,N_34890);
xnor U48154 (N_48154,N_36880,N_31616);
and U48155 (N_48155,N_36760,N_32433);
nand U48156 (N_48156,N_31470,N_35623);
nand U48157 (N_48157,N_32189,N_35570);
xor U48158 (N_48158,N_32844,N_37734);
and U48159 (N_48159,N_38348,N_39719);
nand U48160 (N_48160,N_34338,N_36240);
and U48161 (N_48161,N_37228,N_37611);
xor U48162 (N_48162,N_37763,N_35049);
nor U48163 (N_48163,N_31760,N_31380);
nand U48164 (N_48164,N_39733,N_36445);
and U48165 (N_48165,N_38611,N_33623);
and U48166 (N_48166,N_33582,N_31254);
nand U48167 (N_48167,N_31272,N_31516);
nand U48168 (N_48168,N_34209,N_35068);
and U48169 (N_48169,N_34487,N_32717);
xor U48170 (N_48170,N_30053,N_34202);
nor U48171 (N_48171,N_32039,N_30864);
nand U48172 (N_48172,N_35303,N_37638);
nor U48173 (N_48173,N_35357,N_39920);
xnor U48174 (N_48174,N_39553,N_31185);
xnor U48175 (N_48175,N_33479,N_35699);
xor U48176 (N_48176,N_38883,N_38542);
nand U48177 (N_48177,N_32301,N_33667);
xnor U48178 (N_48178,N_30732,N_36001);
and U48179 (N_48179,N_35128,N_30973);
xnor U48180 (N_48180,N_31392,N_36898);
and U48181 (N_48181,N_34696,N_37130);
xnor U48182 (N_48182,N_32117,N_38581);
or U48183 (N_48183,N_36151,N_33015);
and U48184 (N_48184,N_36454,N_32680);
or U48185 (N_48185,N_38833,N_33452);
or U48186 (N_48186,N_32062,N_30069);
nand U48187 (N_48187,N_38960,N_31612);
and U48188 (N_48188,N_35850,N_31322);
nor U48189 (N_48189,N_34817,N_35786);
xnor U48190 (N_48190,N_31765,N_39659);
nor U48191 (N_48191,N_39571,N_32601);
or U48192 (N_48192,N_36513,N_36708);
and U48193 (N_48193,N_31174,N_32827);
nand U48194 (N_48194,N_34113,N_32747);
nor U48195 (N_48195,N_33773,N_32828);
nor U48196 (N_48196,N_31416,N_38739);
and U48197 (N_48197,N_35075,N_38985);
and U48198 (N_48198,N_38617,N_30340);
nand U48199 (N_48199,N_36401,N_32910);
or U48200 (N_48200,N_30725,N_39896);
or U48201 (N_48201,N_37693,N_39104);
xor U48202 (N_48202,N_30117,N_34835);
nand U48203 (N_48203,N_33266,N_33158);
nand U48204 (N_48204,N_33198,N_31650);
xnor U48205 (N_48205,N_39252,N_31491);
nor U48206 (N_48206,N_30785,N_34557);
and U48207 (N_48207,N_30632,N_35598);
nor U48208 (N_48208,N_32478,N_36587);
or U48209 (N_48209,N_38873,N_36777);
or U48210 (N_48210,N_36824,N_37191);
or U48211 (N_48211,N_34624,N_36757);
nand U48212 (N_48212,N_36701,N_38005);
xor U48213 (N_48213,N_33073,N_38169);
or U48214 (N_48214,N_34067,N_35547);
or U48215 (N_48215,N_37786,N_39250);
xor U48216 (N_48216,N_33318,N_33953);
nand U48217 (N_48217,N_39431,N_30073);
and U48218 (N_48218,N_35169,N_33752);
and U48219 (N_48219,N_30584,N_35420);
nor U48220 (N_48220,N_35148,N_39192);
nand U48221 (N_48221,N_35952,N_35949);
or U48222 (N_48222,N_38069,N_38107);
and U48223 (N_48223,N_31652,N_34894);
and U48224 (N_48224,N_31781,N_38090);
nor U48225 (N_48225,N_37049,N_39235);
and U48226 (N_48226,N_37504,N_38307);
nand U48227 (N_48227,N_30237,N_34110);
and U48228 (N_48228,N_33566,N_33068);
or U48229 (N_48229,N_38947,N_31409);
nand U48230 (N_48230,N_30055,N_30837);
or U48231 (N_48231,N_38244,N_37047);
xor U48232 (N_48232,N_38929,N_32876);
xor U48233 (N_48233,N_38660,N_38742);
nor U48234 (N_48234,N_30074,N_35260);
or U48235 (N_48235,N_37661,N_30353);
nand U48236 (N_48236,N_32413,N_38104);
nor U48237 (N_48237,N_37574,N_30871);
or U48238 (N_48238,N_39172,N_38973);
and U48239 (N_48239,N_36958,N_30990);
and U48240 (N_48240,N_34352,N_31512);
xnor U48241 (N_48241,N_39051,N_38214);
nor U48242 (N_48242,N_34277,N_35552);
nor U48243 (N_48243,N_37078,N_32928);
xor U48244 (N_48244,N_35923,N_31437);
nor U48245 (N_48245,N_36421,N_31359);
nor U48246 (N_48246,N_37266,N_31071);
nor U48247 (N_48247,N_34340,N_34938);
xor U48248 (N_48248,N_36564,N_31449);
nand U48249 (N_48249,N_38973,N_32655);
xor U48250 (N_48250,N_32910,N_35988);
and U48251 (N_48251,N_39231,N_35486);
nor U48252 (N_48252,N_34472,N_35328);
nand U48253 (N_48253,N_31211,N_31200);
and U48254 (N_48254,N_35477,N_33496);
xnor U48255 (N_48255,N_36026,N_38754);
and U48256 (N_48256,N_34461,N_35859);
nand U48257 (N_48257,N_35328,N_39363);
or U48258 (N_48258,N_35655,N_36347);
nor U48259 (N_48259,N_39352,N_31190);
nand U48260 (N_48260,N_34937,N_37353);
nand U48261 (N_48261,N_33445,N_33956);
or U48262 (N_48262,N_34425,N_36228);
xnor U48263 (N_48263,N_30904,N_38864);
nand U48264 (N_48264,N_35690,N_39128);
or U48265 (N_48265,N_33898,N_32803);
xor U48266 (N_48266,N_39365,N_33291);
nand U48267 (N_48267,N_30772,N_32252);
xnor U48268 (N_48268,N_32622,N_36420);
or U48269 (N_48269,N_35716,N_30534);
nor U48270 (N_48270,N_31695,N_37176);
nor U48271 (N_48271,N_33249,N_30321);
and U48272 (N_48272,N_36528,N_34933);
xor U48273 (N_48273,N_34921,N_34379);
or U48274 (N_48274,N_36158,N_33651);
or U48275 (N_48275,N_36894,N_37957);
xor U48276 (N_48276,N_36201,N_36202);
or U48277 (N_48277,N_35404,N_31829);
nand U48278 (N_48278,N_39234,N_33674);
nand U48279 (N_48279,N_36536,N_32464);
nand U48280 (N_48280,N_39272,N_37344);
or U48281 (N_48281,N_38921,N_38602);
and U48282 (N_48282,N_38650,N_30403);
xor U48283 (N_48283,N_31144,N_34455);
xnor U48284 (N_48284,N_32579,N_35136);
or U48285 (N_48285,N_33299,N_36990);
nand U48286 (N_48286,N_39935,N_33697);
nor U48287 (N_48287,N_32435,N_36971);
nor U48288 (N_48288,N_30612,N_38991);
and U48289 (N_48289,N_34614,N_38057);
or U48290 (N_48290,N_31822,N_35065);
nor U48291 (N_48291,N_39643,N_30155);
nor U48292 (N_48292,N_32397,N_39178);
and U48293 (N_48293,N_38364,N_35205);
xor U48294 (N_48294,N_37878,N_36899);
and U48295 (N_48295,N_31706,N_39090);
or U48296 (N_48296,N_30495,N_35328);
nor U48297 (N_48297,N_33062,N_37949);
or U48298 (N_48298,N_35403,N_32969);
or U48299 (N_48299,N_34929,N_32568);
nand U48300 (N_48300,N_31311,N_36244);
nor U48301 (N_48301,N_39063,N_39971);
or U48302 (N_48302,N_35552,N_30446);
nand U48303 (N_48303,N_31286,N_33112);
and U48304 (N_48304,N_39348,N_39968);
nand U48305 (N_48305,N_33654,N_31323);
nor U48306 (N_48306,N_30832,N_35490);
and U48307 (N_48307,N_32574,N_39989);
and U48308 (N_48308,N_34830,N_35901);
nand U48309 (N_48309,N_37444,N_37901);
nand U48310 (N_48310,N_32419,N_36849);
xnor U48311 (N_48311,N_34829,N_37503);
nand U48312 (N_48312,N_30357,N_30325);
nor U48313 (N_48313,N_34626,N_32549);
and U48314 (N_48314,N_39599,N_31648);
and U48315 (N_48315,N_34672,N_36955);
nor U48316 (N_48316,N_31818,N_30798);
or U48317 (N_48317,N_37065,N_35270);
and U48318 (N_48318,N_31817,N_33745);
nand U48319 (N_48319,N_32861,N_32072);
and U48320 (N_48320,N_30728,N_39663);
xor U48321 (N_48321,N_37926,N_38678);
xnor U48322 (N_48322,N_34441,N_34098);
nor U48323 (N_48323,N_38143,N_36682);
or U48324 (N_48324,N_32106,N_38969);
xor U48325 (N_48325,N_36234,N_33372);
nand U48326 (N_48326,N_38854,N_39448);
or U48327 (N_48327,N_37661,N_31091);
xnor U48328 (N_48328,N_33402,N_35438);
nand U48329 (N_48329,N_32811,N_32015);
and U48330 (N_48330,N_30197,N_35765);
nand U48331 (N_48331,N_36720,N_36357);
xor U48332 (N_48332,N_32700,N_37030);
nand U48333 (N_48333,N_36719,N_31576);
or U48334 (N_48334,N_35271,N_38181);
and U48335 (N_48335,N_30983,N_34855);
xor U48336 (N_48336,N_35126,N_34166);
nand U48337 (N_48337,N_33471,N_39704);
xor U48338 (N_48338,N_30628,N_39063);
and U48339 (N_48339,N_39979,N_39585);
nor U48340 (N_48340,N_30274,N_37403);
or U48341 (N_48341,N_38632,N_33034);
xnor U48342 (N_48342,N_39956,N_35000);
nor U48343 (N_48343,N_32001,N_31023);
nand U48344 (N_48344,N_38524,N_37033);
or U48345 (N_48345,N_32107,N_36961);
nor U48346 (N_48346,N_33181,N_39219);
nor U48347 (N_48347,N_39220,N_36041);
xor U48348 (N_48348,N_32885,N_32826);
xor U48349 (N_48349,N_33913,N_37565);
nand U48350 (N_48350,N_36398,N_30434);
nor U48351 (N_48351,N_33678,N_39726);
nor U48352 (N_48352,N_33972,N_33603);
xnor U48353 (N_48353,N_35112,N_37908);
xor U48354 (N_48354,N_39864,N_31461);
xnor U48355 (N_48355,N_37689,N_33705);
and U48356 (N_48356,N_32681,N_38456);
nor U48357 (N_48357,N_35458,N_30901);
and U48358 (N_48358,N_32896,N_35117);
nand U48359 (N_48359,N_39610,N_38361);
nand U48360 (N_48360,N_37311,N_37662);
nand U48361 (N_48361,N_37545,N_33609);
and U48362 (N_48362,N_32983,N_32594);
and U48363 (N_48363,N_38255,N_31888);
or U48364 (N_48364,N_36862,N_30699);
nor U48365 (N_48365,N_35916,N_38919);
nor U48366 (N_48366,N_39472,N_30862);
xor U48367 (N_48367,N_35737,N_33571);
nand U48368 (N_48368,N_34078,N_32276);
or U48369 (N_48369,N_32226,N_32804);
or U48370 (N_48370,N_36672,N_38584);
or U48371 (N_48371,N_39122,N_32650);
xnor U48372 (N_48372,N_33659,N_32091);
or U48373 (N_48373,N_36966,N_36280);
and U48374 (N_48374,N_32358,N_33285);
or U48375 (N_48375,N_35790,N_31372);
nand U48376 (N_48376,N_32381,N_30896);
or U48377 (N_48377,N_33777,N_33911);
nand U48378 (N_48378,N_32879,N_39110);
nor U48379 (N_48379,N_38199,N_38162);
or U48380 (N_48380,N_31454,N_39148);
nor U48381 (N_48381,N_39412,N_37360);
nor U48382 (N_48382,N_38495,N_32308);
nand U48383 (N_48383,N_37568,N_31341);
nor U48384 (N_48384,N_34259,N_33941);
nand U48385 (N_48385,N_33415,N_30172);
or U48386 (N_48386,N_34472,N_30561);
xor U48387 (N_48387,N_34454,N_38431);
and U48388 (N_48388,N_35783,N_34757);
nor U48389 (N_48389,N_35491,N_34442);
nor U48390 (N_48390,N_31210,N_32731);
nor U48391 (N_48391,N_35165,N_38836);
xnor U48392 (N_48392,N_38509,N_30427);
and U48393 (N_48393,N_38278,N_38257);
nand U48394 (N_48394,N_31360,N_34264);
or U48395 (N_48395,N_31247,N_38669);
nand U48396 (N_48396,N_36158,N_36035);
nand U48397 (N_48397,N_33333,N_30502);
xnor U48398 (N_48398,N_38110,N_38254);
nand U48399 (N_48399,N_34698,N_39161);
and U48400 (N_48400,N_35203,N_33095);
nor U48401 (N_48401,N_31855,N_34476);
or U48402 (N_48402,N_32604,N_37639);
nand U48403 (N_48403,N_35800,N_34580);
nand U48404 (N_48404,N_36095,N_33002);
nand U48405 (N_48405,N_31730,N_32910);
nand U48406 (N_48406,N_32120,N_30143);
or U48407 (N_48407,N_39860,N_38808);
nand U48408 (N_48408,N_33439,N_31553);
xor U48409 (N_48409,N_31672,N_37414);
and U48410 (N_48410,N_31741,N_37779);
nand U48411 (N_48411,N_32821,N_37346);
nor U48412 (N_48412,N_35632,N_31771);
nor U48413 (N_48413,N_31090,N_35707);
xor U48414 (N_48414,N_31981,N_32498);
nor U48415 (N_48415,N_34143,N_38042);
xnor U48416 (N_48416,N_36755,N_38354);
or U48417 (N_48417,N_39918,N_39731);
and U48418 (N_48418,N_38027,N_33630);
and U48419 (N_48419,N_39856,N_36254);
and U48420 (N_48420,N_34801,N_36438);
xor U48421 (N_48421,N_39094,N_31740);
nor U48422 (N_48422,N_34315,N_35407);
nand U48423 (N_48423,N_36530,N_38862);
nand U48424 (N_48424,N_33131,N_31443);
or U48425 (N_48425,N_33949,N_39287);
and U48426 (N_48426,N_32665,N_38773);
nor U48427 (N_48427,N_36055,N_30997);
nor U48428 (N_48428,N_32945,N_32961);
xor U48429 (N_48429,N_35807,N_37962);
nand U48430 (N_48430,N_32391,N_35228);
nand U48431 (N_48431,N_34256,N_37159);
nand U48432 (N_48432,N_39482,N_38396);
and U48433 (N_48433,N_36403,N_30977);
nor U48434 (N_48434,N_35182,N_33050);
or U48435 (N_48435,N_33470,N_34291);
xnor U48436 (N_48436,N_34948,N_32889);
nor U48437 (N_48437,N_35425,N_39290);
and U48438 (N_48438,N_37558,N_37978);
nand U48439 (N_48439,N_36290,N_34805);
nand U48440 (N_48440,N_30195,N_37377);
xor U48441 (N_48441,N_39932,N_34137);
or U48442 (N_48442,N_32596,N_31097);
or U48443 (N_48443,N_32156,N_34727);
and U48444 (N_48444,N_39821,N_31204);
and U48445 (N_48445,N_39515,N_35079);
or U48446 (N_48446,N_38105,N_36686);
nor U48447 (N_48447,N_35515,N_32315);
xnor U48448 (N_48448,N_31934,N_30570);
nor U48449 (N_48449,N_39397,N_30117);
nor U48450 (N_48450,N_36778,N_32164);
nand U48451 (N_48451,N_34122,N_33617);
nor U48452 (N_48452,N_30949,N_36530);
and U48453 (N_48453,N_39744,N_31288);
and U48454 (N_48454,N_32829,N_32598);
xor U48455 (N_48455,N_34914,N_35859);
nand U48456 (N_48456,N_35643,N_31023);
nand U48457 (N_48457,N_34601,N_38217);
nor U48458 (N_48458,N_35681,N_30793);
xnor U48459 (N_48459,N_38520,N_36624);
and U48460 (N_48460,N_38785,N_34205);
and U48461 (N_48461,N_39777,N_31360);
or U48462 (N_48462,N_38196,N_36867);
nand U48463 (N_48463,N_37375,N_37452);
or U48464 (N_48464,N_34233,N_35058);
xnor U48465 (N_48465,N_37605,N_30924);
nand U48466 (N_48466,N_36718,N_31155);
nor U48467 (N_48467,N_38137,N_33351);
nor U48468 (N_48468,N_35488,N_33985);
nor U48469 (N_48469,N_30889,N_37255);
nor U48470 (N_48470,N_34631,N_30719);
nor U48471 (N_48471,N_37287,N_35322);
nor U48472 (N_48472,N_37057,N_32310);
nor U48473 (N_48473,N_32977,N_32443);
nand U48474 (N_48474,N_31387,N_38599);
and U48475 (N_48475,N_39955,N_30098);
xor U48476 (N_48476,N_34307,N_37907);
nand U48477 (N_48477,N_32402,N_39850);
or U48478 (N_48478,N_39996,N_39774);
nand U48479 (N_48479,N_36635,N_34760);
nor U48480 (N_48480,N_36743,N_36297);
xor U48481 (N_48481,N_31928,N_32336);
and U48482 (N_48482,N_34075,N_33280);
or U48483 (N_48483,N_33524,N_36751);
xnor U48484 (N_48484,N_39612,N_35823);
or U48485 (N_48485,N_33389,N_33863);
nand U48486 (N_48486,N_33612,N_34041);
nand U48487 (N_48487,N_31315,N_34341);
nor U48488 (N_48488,N_36517,N_31858);
nor U48489 (N_48489,N_35107,N_31810);
and U48490 (N_48490,N_36569,N_35567);
or U48491 (N_48491,N_32627,N_31449);
nor U48492 (N_48492,N_35936,N_39593);
nand U48493 (N_48493,N_31950,N_39208);
or U48494 (N_48494,N_37904,N_38452);
xor U48495 (N_48495,N_30563,N_39670);
and U48496 (N_48496,N_34513,N_32046);
nor U48497 (N_48497,N_31568,N_35890);
xnor U48498 (N_48498,N_37983,N_31508);
xnor U48499 (N_48499,N_34433,N_31387);
and U48500 (N_48500,N_32328,N_35439);
xor U48501 (N_48501,N_35756,N_31492);
nor U48502 (N_48502,N_34376,N_30558);
nor U48503 (N_48503,N_35130,N_31326);
or U48504 (N_48504,N_39657,N_38067);
nand U48505 (N_48505,N_33653,N_39042);
nor U48506 (N_48506,N_32919,N_38088);
or U48507 (N_48507,N_39153,N_38031);
nand U48508 (N_48508,N_35518,N_32019);
xor U48509 (N_48509,N_36500,N_31907);
xor U48510 (N_48510,N_37728,N_34605);
or U48511 (N_48511,N_39260,N_39634);
or U48512 (N_48512,N_30733,N_35072);
and U48513 (N_48513,N_32210,N_39196);
nor U48514 (N_48514,N_30504,N_37578);
and U48515 (N_48515,N_38300,N_32372);
xnor U48516 (N_48516,N_35185,N_30688);
xor U48517 (N_48517,N_36593,N_38793);
and U48518 (N_48518,N_32605,N_35643);
nand U48519 (N_48519,N_39485,N_32006);
and U48520 (N_48520,N_38487,N_36150);
and U48521 (N_48521,N_37392,N_34095);
nor U48522 (N_48522,N_36193,N_37216);
or U48523 (N_48523,N_31163,N_31803);
nor U48524 (N_48524,N_38596,N_38519);
or U48525 (N_48525,N_39843,N_37144);
nand U48526 (N_48526,N_31559,N_34351);
nand U48527 (N_48527,N_33679,N_35018);
nand U48528 (N_48528,N_34986,N_36879);
nor U48529 (N_48529,N_35209,N_34249);
nor U48530 (N_48530,N_35999,N_38707);
nand U48531 (N_48531,N_30658,N_32794);
nor U48532 (N_48532,N_35794,N_32875);
nand U48533 (N_48533,N_39119,N_37122);
and U48534 (N_48534,N_32321,N_37511);
xnor U48535 (N_48535,N_36012,N_36479);
nor U48536 (N_48536,N_38386,N_38280);
xnor U48537 (N_48537,N_30113,N_32663);
and U48538 (N_48538,N_34897,N_32156);
or U48539 (N_48539,N_35853,N_35198);
nand U48540 (N_48540,N_31763,N_32578);
nor U48541 (N_48541,N_35279,N_36321);
and U48542 (N_48542,N_37386,N_37302);
and U48543 (N_48543,N_38943,N_31021);
nand U48544 (N_48544,N_36346,N_31379);
nor U48545 (N_48545,N_34604,N_35049);
and U48546 (N_48546,N_36961,N_30494);
and U48547 (N_48547,N_31556,N_30616);
xor U48548 (N_48548,N_39450,N_36097);
nand U48549 (N_48549,N_31117,N_34893);
nor U48550 (N_48550,N_33973,N_38305);
or U48551 (N_48551,N_36102,N_32478);
and U48552 (N_48552,N_38472,N_38192);
or U48553 (N_48553,N_39357,N_30485);
or U48554 (N_48554,N_30496,N_37027);
nand U48555 (N_48555,N_31754,N_30014);
or U48556 (N_48556,N_34868,N_36815);
or U48557 (N_48557,N_38075,N_39931);
xor U48558 (N_48558,N_34901,N_39445);
nand U48559 (N_48559,N_36115,N_37252);
xnor U48560 (N_48560,N_34100,N_38772);
nand U48561 (N_48561,N_37486,N_32720);
nor U48562 (N_48562,N_35920,N_33136);
and U48563 (N_48563,N_37648,N_30303);
nor U48564 (N_48564,N_32235,N_38900);
nand U48565 (N_48565,N_35505,N_39118);
xor U48566 (N_48566,N_37013,N_39000);
or U48567 (N_48567,N_33689,N_32402);
nor U48568 (N_48568,N_36711,N_35150);
or U48569 (N_48569,N_38371,N_30939);
nand U48570 (N_48570,N_38139,N_34263);
nand U48571 (N_48571,N_36211,N_33956);
nand U48572 (N_48572,N_39669,N_35044);
nor U48573 (N_48573,N_33254,N_38944);
or U48574 (N_48574,N_39801,N_35513);
nand U48575 (N_48575,N_35900,N_31908);
xor U48576 (N_48576,N_39962,N_38029);
nor U48577 (N_48577,N_36561,N_39920);
xnor U48578 (N_48578,N_30056,N_36188);
nor U48579 (N_48579,N_35898,N_39595);
and U48580 (N_48580,N_32848,N_32370);
or U48581 (N_48581,N_31223,N_34661);
or U48582 (N_48582,N_39550,N_37410);
nor U48583 (N_48583,N_32254,N_32162);
or U48584 (N_48584,N_39500,N_36164);
nor U48585 (N_48585,N_32262,N_39547);
nand U48586 (N_48586,N_30120,N_34191);
xnor U48587 (N_48587,N_37872,N_36530);
or U48588 (N_48588,N_38722,N_32282);
and U48589 (N_48589,N_30498,N_33253);
nand U48590 (N_48590,N_36391,N_35845);
xnor U48591 (N_48591,N_36904,N_37183);
nor U48592 (N_48592,N_34116,N_36086);
nor U48593 (N_48593,N_32801,N_34253);
nand U48594 (N_48594,N_35495,N_39111);
nor U48595 (N_48595,N_35625,N_39648);
nor U48596 (N_48596,N_34102,N_34326);
xnor U48597 (N_48597,N_33796,N_39232);
xnor U48598 (N_48598,N_30087,N_36681);
or U48599 (N_48599,N_35725,N_32502);
nor U48600 (N_48600,N_32460,N_33812);
and U48601 (N_48601,N_35633,N_32987);
nor U48602 (N_48602,N_37613,N_31040);
nor U48603 (N_48603,N_32652,N_36235);
xnor U48604 (N_48604,N_39871,N_30714);
nor U48605 (N_48605,N_30003,N_37276);
or U48606 (N_48606,N_35089,N_38782);
nand U48607 (N_48607,N_37536,N_38119);
nor U48608 (N_48608,N_33329,N_38721);
xnor U48609 (N_48609,N_38747,N_33164);
or U48610 (N_48610,N_33155,N_34139);
or U48611 (N_48611,N_32662,N_32233);
and U48612 (N_48612,N_30529,N_36945);
nand U48613 (N_48613,N_33880,N_32190);
xor U48614 (N_48614,N_31361,N_37966);
nor U48615 (N_48615,N_34200,N_30449);
nor U48616 (N_48616,N_34365,N_35948);
or U48617 (N_48617,N_37488,N_34072);
xor U48618 (N_48618,N_35707,N_34593);
nand U48619 (N_48619,N_33085,N_30090);
xnor U48620 (N_48620,N_33427,N_34047);
and U48621 (N_48621,N_35685,N_38961);
nor U48622 (N_48622,N_34231,N_37907);
nand U48623 (N_48623,N_39204,N_35794);
xnor U48624 (N_48624,N_31868,N_37346);
and U48625 (N_48625,N_31378,N_37242);
and U48626 (N_48626,N_30259,N_30469);
or U48627 (N_48627,N_36501,N_32178);
or U48628 (N_48628,N_35706,N_35428);
nor U48629 (N_48629,N_32158,N_34922);
nand U48630 (N_48630,N_38596,N_33954);
nand U48631 (N_48631,N_35408,N_34731);
nand U48632 (N_48632,N_35384,N_37959);
or U48633 (N_48633,N_30892,N_39090);
xor U48634 (N_48634,N_35085,N_36046);
nor U48635 (N_48635,N_31551,N_35650);
nor U48636 (N_48636,N_36466,N_32068);
and U48637 (N_48637,N_35726,N_39689);
nand U48638 (N_48638,N_32112,N_30588);
nand U48639 (N_48639,N_38627,N_39390);
nor U48640 (N_48640,N_32485,N_33666);
nor U48641 (N_48641,N_33390,N_36617);
nor U48642 (N_48642,N_39219,N_39638);
and U48643 (N_48643,N_34945,N_39423);
xor U48644 (N_48644,N_30778,N_38627);
xor U48645 (N_48645,N_34471,N_32103);
or U48646 (N_48646,N_39391,N_38031);
nor U48647 (N_48647,N_39197,N_30706);
or U48648 (N_48648,N_30814,N_30444);
nand U48649 (N_48649,N_32860,N_31026);
nand U48650 (N_48650,N_34104,N_38555);
nor U48651 (N_48651,N_32108,N_31385);
or U48652 (N_48652,N_33118,N_30312);
xor U48653 (N_48653,N_32580,N_37658);
nor U48654 (N_48654,N_30886,N_31366);
nor U48655 (N_48655,N_32655,N_32419);
nor U48656 (N_48656,N_34108,N_38980);
or U48657 (N_48657,N_35334,N_33303);
nor U48658 (N_48658,N_31193,N_34727);
nor U48659 (N_48659,N_30626,N_39186);
nand U48660 (N_48660,N_31636,N_34473);
nand U48661 (N_48661,N_37006,N_31729);
nor U48662 (N_48662,N_39018,N_39921);
nor U48663 (N_48663,N_36005,N_33254);
or U48664 (N_48664,N_38404,N_36014);
nand U48665 (N_48665,N_36586,N_30163);
xor U48666 (N_48666,N_30763,N_36105);
nand U48667 (N_48667,N_37767,N_33789);
nand U48668 (N_48668,N_36810,N_35891);
xor U48669 (N_48669,N_30439,N_34462);
and U48670 (N_48670,N_34482,N_38260);
and U48671 (N_48671,N_37628,N_35202);
nand U48672 (N_48672,N_36955,N_35445);
nand U48673 (N_48673,N_37316,N_31382);
nor U48674 (N_48674,N_36420,N_39801);
nor U48675 (N_48675,N_30712,N_32989);
nor U48676 (N_48676,N_33524,N_33858);
nand U48677 (N_48677,N_37418,N_35844);
nor U48678 (N_48678,N_36306,N_33738);
xnor U48679 (N_48679,N_35877,N_37548);
xnor U48680 (N_48680,N_31734,N_36263);
and U48681 (N_48681,N_31350,N_33497);
nor U48682 (N_48682,N_31074,N_34978);
or U48683 (N_48683,N_30031,N_30096);
nor U48684 (N_48684,N_35113,N_32158);
nor U48685 (N_48685,N_38333,N_34736);
and U48686 (N_48686,N_30674,N_35155);
and U48687 (N_48687,N_37303,N_36334);
or U48688 (N_48688,N_37567,N_39736);
nand U48689 (N_48689,N_35137,N_32049);
nand U48690 (N_48690,N_31219,N_36889);
and U48691 (N_48691,N_31919,N_37260);
nand U48692 (N_48692,N_32686,N_31256);
or U48693 (N_48693,N_30174,N_37197);
xor U48694 (N_48694,N_35192,N_30364);
xnor U48695 (N_48695,N_31320,N_34011);
nand U48696 (N_48696,N_37640,N_34979);
nand U48697 (N_48697,N_32707,N_32086);
and U48698 (N_48698,N_39146,N_32230);
nand U48699 (N_48699,N_33214,N_39859);
nor U48700 (N_48700,N_31810,N_32092);
nand U48701 (N_48701,N_31542,N_36542);
nand U48702 (N_48702,N_31393,N_37131);
or U48703 (N_48703,N_32766,N_32099);
xnor U48704 (N_48704,N_32420,N_32741);
xnor U48705 (N_48705,N_37307,N_38021);
or U48706 (N_48706,N_34138,N_39506);
or U48707 (N_48707,N_37438,N_30524);
nand U48708 (N_48708,N_35701,N_32124);
nand U48709 (N_48709,N_30283,N_35243);
xnor U48710 (N_48710,N_31504,N_35749);
nand U48711 (N_48711,N_33462,N_30140);
nand U48712 (N_48712,N_32543,N_32599);
and U48713 (N_48713,N_39908,N_34716);
xnor U48714 (N_48714,N_37761,N_31725);
and U48715 (N_48715,N_32050,N_36540);
nor U48716 (N_48716,N_36336,N_35932);
nand U48717 (N_48717,N_33786,N_35287);
nor U48718 (N_48718,N_38308,N_37163);
or U48719 (N_48719,N_38114,N_35035);
nand U48720 (N_48720,N_39144,N_36092);
or U48721 (N_48721,N_39923,N_38872);
xnor U48722 (N_48722,N_38545,N_33605);
nor U48723 (N_48723,N_38270,N_33699);
nand U48724 (N_48724,N_32509,N_36794);
or U48725 (N_48725,N_30003,N_32160);
xor U48726 (N_48726,N_35907,N_35822);
or U48727 (N_48727,N_30437,N_39387);
nand U48728 (N_48728,N_34502,N_30103);
xor U48729 (N_48729,N_33790,N_35375);
or U48730 (N_48730,N_34336,N_35849);
nor U48731 (N_48731,N_39314,N_31919);
nand U48732 (N_48732,N_30293,N_30769);
nor U48733 (N_48733,N_39807,N_30113);
nand U48734 (N_48734,N_37739,N_31147);
nand U48735 (N_48735,N_31317,N_33723);
and U48736 (N_48736,N_34517,N_31078);
and U48737 (N_48737,N_32854,N_30078);
and U48738 (N_48738,N_32770,N_33774);
nand U48739 (N_48739,N_34496,N_38113);
xnor U48740 (N_48740,N_32202,N_35207);
xor U48741 (N_48741,N_35974,N_38445);
nand U48742 (N_48742,N_34705,N_33619);
nand U48743 (N_48743,N_35452,N_33619);
and U48744 (N_48744,N_34991,N_32441);
and U48745 (N_48745,N_38752,N_32443);
and U48746 (N_48746,N_30193,N_37606);
xor U48747 (N_48747,N_32581,N_30138);
xor U48748 (N_48748,N_30296,N_30842);
nand U48749 (N_48749,N_31641,N_36337);
xor U48750 (N_48750,N_37814,N_36470);
and U48751 (N_48751,N_31978,N_36730);
xor U48752 (N_48752,N_36715,N_34563);
nor U48753 (N_48753,N_30243,N_37502);
nand U48754 (N_48754,N_31111,N_33171);
nor U48755 (N_48755,N_37588,N_38310);
nand U48756 (N_48756,N_35010,N_36366);
and U48757 (N_48757,N_38597,N_37593);
and U48758 (N_48758,N_39122,N_33168);
and U48759 (N_48759,N_30325,N_31252);
or U48760 (N_48760,N_36825,N_39244);
or U48761 (N_48761,N_34121,N_38433);
xnor U48762 (N_48762,N_31289,N_30223);
and U48763 (N_48763,N_35872,N_32209);
nand U48764 (N_48764,N_33390,N_34799);
xor U48765 (N_48765,N_39038,N_31266);
nand U48766 (N_48766,N_36473,N_34793);
nand U48767 (N_48767,N_31746,N_38984);
nand U48768 (N_48768,N_39123,N_31058);
xnor U48769 (N_48769,N_30074,N_30572);
nand U48770 (N_48770,N_31930,N_33109);
or U48771 (N_48771,N_31499,N_31943);
nand U48772 (N_48772,N_32565,N_39687);
nand U48773 (N_48773,N_31044,N_30668);
xor U48774 (N_48774,N_35696,N_38651);
xnor U48775 (N_48775,N_37425,N_38811);
nand U48776 (N_48776,N_38415,N_32140);
xnor U48777 (N_48777,N_36160,N_34824);
nand U48778 (N_48778,N_39364,N_39634);
and U48779 (N_48779,N_38031,N_36634);
nor U48780 (N_48780,N_30920,N_39736);
nand U48781 (N_48781,N_35314,N_35189);
or U48782 (N_48782,N_37733,N_32540);
and U48783 (N_48783,N_33290,N_30633);
and U48784 (N_48784,N_30618,N_30826);
or U48785 (N_48785,N_36276,N_36536);
and U48786 (N_48786,N_37969,N_34954);
nor U48787 (N_48787,N_38335,N_39414);
and U48788 (N_48788,N_39136,N_38346);
or U48789 (N_48789,N_32475,N_33275);
or U48790 (N_48790,N_30258,N_31107);
xnor U48791 (N_48791,N_36684,N_37154);
xor U48792 (N_48792,N_36986,N_38771);
nor U48793 (N_48793,N_30088,N_30807);
or U48794 (N_48794,N_35617,N_30727);
nand U48795 (N_48795,N_39236,N_34299);
nand U48796 (N_48796,N_37536,N_31729);
or U48797 (N_48797,N_31858,N_34318);
nor U48798 (N_48798,N_38769,N_32780);
and U48799 (N_48799,N_39434,N_31061);
nor U48800 (N_48800,N_39994,N_32962);
and U48801 (N_48801,N_35906,N_33907);
and U48802 (N_48802,N_31381,N_34697);
and U48803 (N_48803,N_32293,N_32780);
xor U48804 (N_48804,N_34054,N_35033);
nand U48805 (N_48805,N_33769,N_37124);
xnor U48806 (N_48806,N_30468,N_36931);
xnor U48807 (N_48807,N_38365,N_33396);
or U48808 (N_48808,N_33988,N_39379);
and U48809 (N_48809,N_35560,N_36119);
and U48810 (N_48810,N_37507,N_34989);
and U48811 (N_48811,N_31561,N_33188);
or U48812 (N_48812,N_31968,N_39329);
or U48813 (N_48813,N_33006,N_31556);
and U48814 (N_48814,N_38919,N_37561);
xor U48815 (N_48815,N_36220,N_35161);
nand U48816 (N_48816,N_36917,N_34787);
and U48817 (N_48817,N_36353,N_38194);
xor U48818 (N_48818,N_31441,N_35357);
xnor U48819 (N_48819,N_30909,N_37880);
and U48820 (N_48820,N_35285,N_30063);
and U48821 (N_48821,N_32987,N_33443);
xnor U48822 (N_48822,N_33812,N_37078);
nand U48823 (N_48823,N_30050,N_34238);
and U48824 (N_48824,N_38971,N_32046);
xnor U48825 (N_48825,N_39350,N_31508);
and U48826 (N_48826,N_35995,N_32194);
nor U48827 (N_48827,N_37452,N_33503);
nor U48828 (N_48828,N_36926,N_32938);
nand U48829 (N_48829,N_37917,N_38599);
or U48830 (N_48830,N_36680,N_32970);
xnor U48831 (N_48831,N_38375,N_37031);
xor U48832 (N_48832,N_32313,N_34068);
nor U48833 (N_48833,N_37822,N_34827);
nand U48834 (N_48834,N_38377,N_30824);
and U48835 (N_48835,N_36865,N_30395);
nor U48836 (N_48836,N_35717,N_33901);
xnor U48837 (N_48837,N_32601,N_34130);
xor U48838 (N_48838,N_34854,N_37237);
or U48839 (N_48839,N_34705,N_38476);
xnor U48840 (N_48840,N_31088,N_39542);
nor U48841 (N_48841,N_36857,N_31859);
xnor U48842 (N_48842,N_37381,N_38276);
xnor U48843 (N_48843,N_32716,N_38948);
xor U48844 (N_48844,N_37402,N_38726);
and U48845 (N_48845,N_37194,N_35077);
and U48846 (N_48846,N_33100,N_36416);
nand U48847 (N_48847,N_34697,N_30029);
and U48848 (N_48848,N_38532,N_31991);
nand U48849 (N_48849,N_39566,N_34223);
xor U48850 (N_48850,N_32466,N_37231);
nand U48851 (N_48851,N_33587,N_36196);
xnor U48852 (N_48852,N_34990,N_35131);
nor U48853 (N_48853,N_37050,N_34705);
nor U48854 (N_48854,N_30106,N_37621);
xor U48855 (N_48855,N_30225,N_34938);
and U48856 (N_48856,N_34653,N_36526);
xor U48857 (N_48857,N_35130,N_30490);
xor U48858 (N_48858,N_39378,N_37846);
or U48859 (N_48859,N_34053,N_35398);
and U48860 (N_48860,N_38605,N_34160);
nand U48861 (N_48861,N_30896,N_38680);
nor U48862 (N_48862,N_38422,N_36428);
nand U48863 (N_48863,N_33188,N_33930);
or U48864 (N_48864,N_37323,N_37457);
and U48865 (N_48865,N_34057,N_30077);
nor U48866 (N_48866,N_33989,N_35675);
or U48867 (N_48867,N_39530,N_33323);
nor U48868 (N_48868,N_33582,N_39015);
or U48869 (N_48869,N_37646,N_39338);
nor U48870 (N_48870,N_32905,N_35060);
nand U48871 (N_48871,N_38604,N_38684);
nand U48872 (N_48872,N_34232,N_33009);
or U48873 (N_48873,N_30936,N_32126);
or U48874 (N_48874,N_31246,N_34267);
or U48875 (N_48875,N_35321,N_38467);
xor U48876 (N_48876,N_34925,N_39387);
nor U48877 (N_48877,N_37527,N_34524);
or U48878 (N_48878,N_36550,N_38170);
xnor U48879 (N_48879,N_34467,N_34673);
or U48880 (N_48880,N_33044,N_37899);
nor U48881 (N_48881,N_39562,N_31759);
and U48882 (N_48882,N_37719,N_32036);
nand U48883 (N_48883,N_34856,N_32610);
nand U48884 (N_48884,N_33852,N_39565);
xor U48885 (N_48885,N_30972,N_39292);
nand U48886 (N_48886,N_33581,N_38728);
nor U48887 (N_48887,N_38302,N_32401);
xor U48888 (N_48888,N_38217,N_39165);
xnor U48889 (N_48889,N_34862,N_37415);
or U48890 (N_48890,N_30822,N_39218);
xor U48891 (N_48891,N_39339,N_37077);
xor U48892 (N_48892,N_34612,N_31150);
xnor U48893 (N_48893,N_33629,N_35859);
xnor U48894 (N_48894,N_37770,N_34925);
nor U48895 (N_48895,N_31538,N_31601);
xnor U48896 (N_48896,N_34832,N_35399);
or U48897 (N_48897,N_30934,N_31028);
nor U48898 (N_48898,N_31851,N_32966);
and U48899 (N_48899,N_37287,N_33334);
and U48900 (N_48900,N_31583,N_39295);
xnor U48901 (N_48901,N_34503,N_32214);
or U48902 (N_48902,N_37978,N_36991);
and U48903 (N_48903,N_39130,N_39630);
xnor U48904 (N_48904,N_33204,N_33635);
nand U48905 (N_48905,N_36074,N_34583);
nand U48906 (N_48906,N_35556,N_36608);
nor U48907 (N_48907,N_30387,N_39595);
xnor U48908 (N_48908,N_38070,N_32441);
nand U48909 (N_48909,N_32113,N_30496);
and U48910 (N_48910,N_37443,N_35851);
nand U48911 (N_48911,N_32765,N_39179);
nand U48912 (N_48912,N_30649,N_32815);
nand U48913 (N_48913,N_36273,N_31959);
and U48914 (N_48914,N_35274,N_31442);
and U48915 (N_48915,N_37338,N_36796);
xnor U48916 (N_48916,N_39363,N_37754);
xor U48917 (N_48917,N_36272,N_37366);
xor U48918 (N_48918,N_39434,N_39053);
nand U48919 (N_48919,N_38325,N_36721);
or U48920 (N_48920,N_33737,N_31201);
nand U48921 (N_48921,N_37998,N_39245);
nand U48922 (N_48922,N_32294,N_37898);
xnor U48923 (N_48923,N_34856,N_39470);
xnor U48924 (N_48924,N_33910,N_30734);
and U48925 (N_48925,N_32695,N_33251);
and U48926 (N_48926,N_33360,N_39436);
or U48927 (N_48927,N_37490,N_32632);
and U48928 (N_48928,N_38590,N_36532);
xnor U48929 (N_48929,N_30434,N_36235);
nor U48930 (N_48930,N_36029,N_38785);
xnor U48931 (N_48931,N_39624,N_30718);
nand U48932 (N_48932,N_36150,N_31340);
nor U48933 (N_48933,N_33727,N_34746);
nor U48934 (N_48934,N_33582,N_31990);
and U48935 (N_48935,N_32945,N_37250);
or U48936 (N_48936,N_38694,N_34083);
xor U48937 (N_48937,N_39195,N_39070);
and U48938 (N_48938,N_31166,N_33920);
or U48939 (N_48939,N_33257,N_35148);
or U48940 (N_48940,N_39568,N_37716);
or U48941 (N_48941,N_33640,N_39346);
xor U48942 (N_48942,N_33256,N_32827);
and U48943 (N_48943,N_39968,N_36307);
or U48944 (N_48944,N_39427,N_39110);
or U48945 (N_48945,N_38347,N_34679);
nor U48946 (N_48946,N_32728,N_39635);
xor U48947 (N_48947,N_33945,N_35175);
nand U48948 (N_48948,N_31504,N_32329);
nor U48949 (N_48949,N_32094,N_31664);
and U48950 (N_48950,N_36919,N_39718);
and U48951 (N_48951,N_35716,N_30424);
nor U48952 (N_48952,N_33366,N_30930);
and U48953 (N_48953,N_35863,N_35240);
xnor U48954 (N_48954,N_35377,N_31988);
nand U48955 (N_48955,N_31526,N_31251);
or U48956 (N_48956,N_33413,N_38722);
xor U48957 (N_48957,N_34144,N_36485);
xor U48958 (N_48958,N_34675,N_30850);
xor U48959 (N_48959,N_37466,N_38231);
nand U48960 (N_48960,N_39086,N_30677);
and U48961 (N_48961,N_38727,N_37085);
or U48962 (N_48962,N_37116,N_36646);
and U48963 (N_48963,N_34914,N_31636);
nor U48964 (N_48964,N_34892,N_30502);
nand U48965 (N_48965,N_39731,N_39404);
nor U48966 (N_48966,N_35788,N_37143);
nor U48967 (N_48967,N_36516,N_38449);
nor U48968 (N_48968,N_35811,N_33070);
xor U48969 (N_48969,N_30887,N_34208);
nand U48970 (N_48970,N_30549,N_35121);
or U48971 (N_48971,N_32989,N_35226);
or U48972 (N_48972,N_33348,N_36878);
or U48973 (N_48973,N_34063,N_37106);
and U48974 (N_48974,N_31933,N_39991);
nor U48975 (N_48975,N_39798,N_31143);
xor U48976 (N_48976,N_32142,N_38262);
and U48977 (N_48977,N_36992,N_33935);
xnor U48978 (N_48978,N_37015,N_31267);
nor U48979 (N_48979,N_36398,N_39878);
nand U48980 (N_48980,N_32099,N_34938);
or U48981 (N_48981,N_30517,N_32787);
and U48982 (N_48982,N_34777,N_39062);
or U48983 (N_48983,N_38412,N_34366);
or U48984 (N_48984,N_30995,N_30845);
nand U48985 (N_48985,N_35386,N_35332);
nand U48986 (N_48986,N_35172,N_30323);
nand U48987 (N_48987,N_32116,N_30586);
or U48988 (N_48988,N_35817,N_37221);
and U48989 (N_48989,N_34579,N_30586);
nand U48990 (N_48990,N_36777,N_31603);
and U48991 (N_48991,N_37127,N_33164);
nand U48992 (N_48992,N_38517,N_36359);
nand U48993 (N_48993,N_33611,N_31565);
nor U48994 (N_48994,N_38231,N_34009);
nand U48995 (N_48995,N_34819,N_30804);
nand U48996 (N_48996,N_33865,N_32234);
and U48997 (N_48997,N_31413,N_38756);
or U48998 (N_48998,N_36397,N_34059);
nand U48999 (N_48999,N_31948,N_33851);
nand U49000 (N_49000,N_37253,N_37511);
or U49001 (N_49001,N_35661,N_39935);
and U49002 (N_49002,N_31815,N_31545);
or U49003 (N_49003,N_34584,N_37488);
or U49004 (N_49004,N_31992,N_32992);
and U49005 (N_49005,N_34398,N_31366);
or U49006 (N_49006,N_31519,N_39664);
nand U49007 (N_49007,N_33976,N_36644);
nand U49008 (N_49008,N_39365,N_39915);
nand U49009 (N_49009,N_34456,N_31870);
nor U49010 (N_49010,N_35337,N_34714);
nand U49011 (N_49011,N_38659,N_38606);
nor U49012 (N_49012,N_30742,N_39858);
or U49013 (N_49013,N_37410,N_39193);
xnor U49014 (N_49014,N_35677,N_38769);
nand U49015 (N_49015,N_32763,N_32528);
xor U49016 (N_49016,N_34046,N_34791);
nand U49017 (N_49017,N_32081,N_33431);
and U49018 (N_49018,N_35105,N_30026);
xor U49019 (N_49019,N_32243,N_39312);
nand U49020 (N_49020,N_33822,N_38295);
or U49021 (N_49021,N_32831,N_37921);
nand U49022 (N_49022,N_38087,N_33381);
and U49023 (N_49023,N_32440,N_30879);
xnor U49024 (N_49024,N_35817,N_31942);
xnor U49025 (N_49025,N_34652,N_34819);
and U49026 (N_49026,N_36588,N_37331);
and U49027 (N_49027,N_32956,N_30571);
or U49028 (N_49028,N_34844,N_37965);
nand U49029 (N_49029,N_36740,N_32971);
nand U49030 (N_49030,N_35095,N_31607);
nand U49031 (N_49031,N_31849,N_35972);
nand U49032 (N_49032,N_33873,N_39526);
nor U49033 (N_49033,N_39815,N_37272);
nand U49034 (N_49034,N_39364,N_33580);
xnor U49035 (N_49035,N_35873,N_37614);
and U49036 (N_49036,N_37363,N_39172);
xnor U49037 (N_49037,N_39409,N_39883);
xor U49038 (N_49038,N_30403,N_33940);
xor U49039 (N_49039,N_35536,N_30185);
xnor U49040 (N_49040,N_31546,N_31403);
xor U49041 (N_49041,N_34231,N_32026);
xnor U49042 (N_49042,N_31016,N_39584);
xnor U49043 (N_49043,N_35316,N_38602);
xnor U49044 (N_49044,N_34159,N_34904);
nand U49045 (N_49045,N_31566,N_39091);
and U49046 (N_49046,N_38674,N_30034);
xnor U49047 (N_49047,N_32364,N_32319);
xor U49048 (N_49048,N_31768,N_38144);
or U49049 (N_49049,N_31098,N_30265);
or U49050 (N_49050,N_33781,N_30350);
xnor U49051 (N_49051,N_33896,N_34407);
xor U49052 (N_49052,N_33531,N_37081);
nor U49053 (N_49053,N_30502,N_31876);
and U49054 (N_49054,N_37225,N_35913);
nand U49055 (N_49055,N_38816,N_37875);
and U49056 (N_49056,N_38114,N_37905);
nand U49057 (N_49057,N_31338,N_33806);
nor U49058 (N_49058,N_30874,N_32161);
and U49059 (N_49059,N_35054,N_36164);
nor U49060 (N_49060,N_36310,N_34117);
xor U49061 (N_49061,N_35799,N_35610);
nand U49062 (N_49062,N_31310,N_34943);
and U49063 (N_49063,N_35333,N_33565);
nand U49064 (N_49064,N_36623,N_35440);
xor U49065 (N_49065,N_37195,N_30009);
or U49066 (N_49066,N_37143,N_33029);
or U49067 (N_49067,N_37205,N_34428);
nand U49068 (N_49068,N_35431,N_39086);
and U49069 (N_49069,N_38291,N_38391);
nor U49070 (N_49070,N_38071,N_31048);
and U49071 (N_49071,N_35362,N_35492);
nand U49072 (N_49072,N_33354,N_32071);
nor U49073 (N_49073,N_34179,N_36091);
xnor U49074 (N_49074,N_36449,N_31530);
nor U49075 (N_49075,N_33449,N_39032);
or U49076 (N_49076,N_34720,N_32524);
and U49077 (N_49077,N_31901,N_32738);
and U49078 (N_49078,N_30219,N_38960);
xor U49079 (N_49079,N_34196,N_36861);
nand U49080 (N_49080,N_32045,N_30439);
nor U49081 (N_49081,N_35039,N_39282);
nand U49082 (N_49082,N_33859,N_36595);
nor U49083 (N_49083,N_33117,N_31441);
or U49084 (N_49084,N_34726,N_37513);
and U49085 (N_49085,N_32201,N_38644);
and U49086 (N_49086,N_34923,N_35656);
nand U49087 (N_49087,N_34042,N_36120);
nor U49088 (N_49088,N_37754,N_36053);
or U49089 (N_49089,N_31964,N_39838);
xnor U49090 (N_49090,N_37634,N_38949);
and U49091 (N_49091,N_30223,N_30484);
or U49092 (N_49092,N_38136,N_37986);
nor U49093 (N_49093,N_36247,N_35689);
nand U49094 (N_49094,N_39806,N_30521);
or U49095 (N_49095,N_33211,N_34043);
or U49096 (N_49096,N_30291,N_32624);
nand U49097 (N_49097,N_32464,N_33393);
xor U49098 (N_49098,N_36754,N_35165);
and U49099 (N_49099,N_31728,N_39214);
nor U49100 (N_49100,N_30726,N_35144);
or U49101 (N_49101,N_32290,N_32298);
and U49102 (N_49102,N_33919,N_36136);
nand U49103 (N_49103,N_34053,N_33888);
xor U49104 (N_49104,N_37934,N_32146);
xnor U49105 (N_49105,N_32785,N_32562);
nand U49106 (N_49106,N_34875,N_30529);
nand U49107 (N_49107,N_31528,N_31556);
or U49108 (N_49108,N_34366,N_30777);
nand U49109 (N_49109,N_38769,N_37172);
and U49110 (N_49110,N_38884,N_36340);
xnor U49111 (N_49111,N_38371,N_32471);
and U49112 (N_49112,N_31427,N_32521);
and U49113 (N_49113,N_33193,N_38399);
nor U49114 (N_49114,N_38250,N_34911);
or U49115 (N_49115,N_37749,N_39548);
and U49116 (N_49116,N_31493,N_35699);
and U49117 (N_49117,N_32940,N_38430);
nand U49118 (N_49118,N_30616,N_30165);
and U49119 (N_49119,N_36375,N_33624);
and U49120 (N_49120,N_34830,N_32952);
xor U49121 (N_49121,N_33631,N_37507);
and U49122 (N_49122,N_39824,N_38225);
or U49123 (N_49123,N_36551,N_38631);
and U49124 (N_49124,N_31728,N_32128);
or U49125 (N_49125,N_38565,N_39059);
nand U49126 (N_49126,N_34322,N_35059);
nor U49127 (N_49127,N_30053,N_34891);
or U49128 (N_49128,N_34543,N_39134);
xnor U49129 (N_49129,N_38000,N_33400);
nand U49130 (N_49130,N_34721,N_30941);
or U49131 (N_49131,N_31990,N_30839);
or U49132 (N_49132,N_33770,N_33260);
and U49133 (N_49133,N_33841,N_30540);
nand U49134 (N_49134,N_37770,N_35133);
and U49135 (N_49135,N_33815,N_34857);
and U49136 (N_49136,N_35665,N_30527);
and U49137 (N_49137,N_33521,N_38379);
and U49138 (N_49138,N_35923,N_36044);
nand U49139 (N_49139,N_39091,N_39115);
or U49140 (N_49140,N_37179,N_32137);
and U49141 (N_49141,N_39677,N_30743);
nand U49142 (N_49142,N_36011,N_34419);
nor U49143 (N_49143,N_38507,N_37701);
nor U49144 (N_49144,N_31534,N_37816);
nand U49145 (N_49145,N_35603,N_36413);
or U49146 (N_49146,N_31327,N_39609);
nor U49147 (N_49147,N_31883,N_30768);
nor U49148 (N_49148,N_33149,N_31069);
or U49149 (N_49149,N_35828,N_37037);
xor U49150 (N_49150,N_30764,N_31961);
nand U49151 (N_49151,N_30189,N_31610);
nor U49152 (N_49152,N_31199,N_32281);
xor U49153 (N_49153,N_38283,N_34386);
and U49154 (N_49154,N_33419,N_30409);
nand U49155 (N_49155,N_36133,N_39359);
xor U49156 (N_49156,N_36113,N_39293);
nor U49157 (N_49157,N_35910,N_30369);
nor U49158 (N_49158,N_37574,N_35957);
or U49159 (N_49159,N_30244,N_32459);
xnor U49160 (N_49160,N_35312,N_32870);
and U49161 (N_49161,N_33593,N_35447);
and U49162 (N_49162,N_37647,N_38581);
xnor U49163 (N_49163,N_30923,N_39834);
xnor U49164 (N_49164,N_35675,N_35144);
nand U49165 (N_49165,N_38994,N_31714);
xnor U49166 (N_49166,N_34276,N_36992);
and U49167 (N_49167,N_31635,N_34327);
xor U49168 (N_49168,N_39431,N_36784);
nand U49169 (N_49169,N_31171,N_39073);
or U49170 (N_49170,N_36207,N_37944);
xor U49171 (N_49171,N_32412,N_34158);
and U49172 (N_49172,N_36225,N_30114);
nand U49173 (N_49173,N_39747,N_32411);
and U49174 (N_49174,N_30060,N_36479);
nand U49175 (N_49175,N_35838,N_38207);
and U49176 (N_49176,N_38999,N_38690);
nand U49177 (N_49177,N_32946,N_33426);
and U49178 (N_49178,N_30982,N_37959);
nand U49179 (N_49179,N_30849,N_31514);
nor U49180 (N_49180,N_36266,N_35359);
nor U49181 (N_49181,N_30002,N_39225);
nor U49182 (N_49182,N_37537,N_32173);
or U49183 (N_49183,N_30648,N_34523);
or U49184 (N_49184,N_37574,N_31656);
nand U49185 (N_49185,N_38467,N_33121);
nor U49186 (N_49186,N_34742,N_33487);
or U49187 (N_49187,N_32600,N_37236);
xnor U49188 (N_49188,N_39381,N_35780);
or U49189 (N_49189,N_38819,N_39717);
nor U49190 (N_49190,N_31448,N_33086);
and U49191 (N_49191,N_31460,N_37102);
nand U49192 (N_49192,N_32338,N_31280);
nand U49193 (N_49193,N_37391,N_32237);
and U49194 (N_49194,N_34183,N_36133);
and U49195 (N_49195,N_33338,N_34496);
nor U49196 (N_49196,N_37162,N_32344);
nand U49197 (N_49197,N_33188,N_30161);
nand U49198 (N_49198,N_31311,N_39401);
nand U49199 (N_49199,N_31413,N_38110);
or U49200 (N_49200,N_36552,N_39053);
nor U49201 (N_49201,N_38895,N_35549);
xor U49202 (N_49202,N_34899,N_30324);
or U49203 (N_49203,N_32529,N_38150);
nand U49204 (N_49204,N_31903,N_30824);
xnor U49205 (N_49205,N_30844,N_34066);
xnor U49206 (N_49206,N_36803,N_31756);
nor U49207 (N_49207,N_31956,N_32376);
nand U49208 (N_49208,N_32042,N_38608);
and U49209 (N_49209,N_39255,N_39926);
and U49210 (N_49210,N_31630,N_30383);
nor U49211 (N_49211,N_31460,N_32760);
and U49212 (N_49212,N_34543,N_33172);
xor U49213 (N_49213,N_33744,N_34908);
nand U49214 (N_49214,N_38470,N_35803);
nor U49215 (N_49215,N_38737,N_30081);
and U49216 (N_49216,N_35152,N_32488);
and U49217 (N_49217,N_31222,N_31825);
nand U49218 (N_49218,N_32450,N_32292);
xor U49219 (N_49219,N_36523,N_38664);
xor U49220 (N_49220,N_36086,N_37224);
nand U49221 (N_49221,N_32000,N_37440);
xnor U49222 (N_49222,N_38287,N_30884);
nand U49223 (N_49223,N_35519,N_38681);
and U49224 (N_49224,N_36535,N_39326);
or U49225 (N_49225,N_38331,N_37904);
nand U49226 (N_49226,N_31237,N_32694);
or U49227 (N_49227,N_39826,N_37755);
nand U49228 (N_49228,N_33829,N_31851);
or U49229 (N_49229,N_33718,N_37011);
and U49230 (N_49230,N_39398,N_34165);
nand U49231 (N_49231,N_39240,N_36593);
nand U49232 (N_49232,N_31769,N_35958);
or U49233 (N_49233,N_35202,N_30763);
and U49234 (N_49234,N_33104,N_30863);
xnor U49235 (N_49235,N_39934,N_34221);
and U49236 (N_49236,N_31156,N_39961);
and U49237 (N_49237,N_33744,N_33288);
nand U49238 (N_49238,N_37066,N_30427);
nor U49239 (N_49239,N_33730,N_35741);
nand U49240 (N_49240,N_36090,N_38475);
or U49241 (N_49241,N_33425,N_39536);
nor U49242 (N_49242,N_31887,N_34424);
nand U49243 (N_49243,N_31776,N_30663);
and U49244 (N_49244,N_32900,N_33512);
or U49245 (N_49245,N_37302,N_37165);
nor U49246 (N_49246,N_36634,N_31793);
and U49247 (N_49247,N_35416,N_35059);
and U49248 (N_49248,N_30328,N_35478);
or U49249 (N_49249,N_30417,N_34396);
nor U49250 (N_49250,N_32942,N_33786);
and U49251 (N_49251,N_39890,N_38096);
or U49252 (N_49252,N_39745,N_33264);
nand U49253 (N_49253,N_31006,N_34973);
or U49254 (N_49254,N_32241,N_39474);
nand U49255 (N_49255,N_36002,N_36318);
nand U49256 (N_49256,N_30551,N_38600);
nor U49257 (N_49257,N_31542,N_30889);
nand U49258 (N_49258,N_39572,N_35322);
xnor U49259 (N_49259,N_38838,N_37169);
and U49260 (N_49260,N_39482,N_38060);
nand U49261 (N_49261,N_35712,N_31729);
xnor U49262 (N_49262,N_30245,N_39067);
nor U49263 (N_49263,N_32268,N_39239);
nor U49264 (N_49264,N_32024,N_37920);
or U49265 (N_49265,N_34029,N_38123);
nand U49266 (N_49266,N_38190,N_35596);
and U49267 (N_49267,N_37019,N_35778);
xor U49268 (N_49268,N_38056,N_35419);
nor U49269 (N_49269,N_30286,N_36540);
and U49270 (N_49270,N_39607,N_39642);
or U49271 (N_49271,N_31049,N_39265);
nand U49272 (N_49272,N_37403,N_39233);
and U49273 (N_49273,N_35101,N_38035);
xnor U49274 (N_49274,N_35449,N_33387);
xnor U49275 (N_49275,N_35173,N_30305);
and U49276 (N_49276,N_37755,N_36846);
nor U49277 (N_49277,N_32775,N_33095);
nor U49278 (N_49278,N_30039,N_36739);
or U49279 (N_49279,N_36996,N_32174);
xor U49280 (N_49280,N_35021,N_34175);
or U49281 (N_49281,N_33214,N_30460);
xor U49282 (N_49282,N_38171,N_31372);
xnor U49283 (N_49283,N_38753,N_38217);
nor U49284 (N_49284,N_36239,N_34015);
xor U49285 (N_49285,N_38673,N_31484);
and U49286 (N_49286,N_31577,N_34817);
or U49287 (N_49287,N_34998,N_32387);
xor U49288 (N_49288,N_33648,N_37115);
or U49289 (N_49289,N_31881,N_34214);
nor U49290 (N_49290,N_38178,N_33495);
xor U49291 (N_49291,N_33970,N_36687);
or U49292 (N_49292,N_31805,N_31139);
or U49293 (N_49293,N_38656,N_30834);
xnor U49294 (N_49294,N_30407,N_37391);
or U49295 (N_49295,N_30768,N_39136);
nor U49296 (N_49296,N_31713,N_35504);
nand U49297 (N_49297,N_38781,N_34941);
nand U49298 (N_49298,N_33373,N_31579);
or U49299 (N_49299,N_38256,N_32700);
nand U49300 (N_49300,N_31122,N_38591);
xnor U49301 (N_49301,N_35811,N_33173);
or U49302 (N_49302,N_37184,N_32282);
nand U49303 (N_49303,N_38979,N_37491);
xor U49304 (N_49304,N_34187,N_32849);
or U49305 (N_49305,N_35531,N_33719);
nor U49306 (N_49306,N_33673,N_39694);
and U49307 (N_49307,N_33391,N_32301);
nor U49308 (N_49308,N_36319,N_39277);
nand U49309 (N_49309,N_36146,N_36974);
or U49310 (N_49310,N_36152,N_39700);
xor U49311 (N_49311,N_37513,N_39005);
or U49312 (N_49312,N_39080,N_39116);
xnor U49313 (N_49313,N_36845,N_36775);
nand U49314 (N_49314,N_35450,N_34095);
and U49315 (N_49315,N_38948,N_39507);
or U49316 (N_49316,N_38260,N_38552);
nand U49317 (N_49317,N_39647,N_30114);
nand U49318 (N_49318,N_33676,N_33322);
xor U49319 (N_49319,N_34771,N_32002);
nor U49320 (N_49320,N_32762,N_31955);
nand U49321 (N_49321,N_38168,N_39066);
nand U49322 (N_49322,N_30651,N_39029);
and U49323 (N_49323,N_33035,N_35827);
xnor U49324 (N_49324,N_31039,N_36241);
and U49325 (N_49325,N_37853,N_30375);
nand U49326 (N_49326,N_38005,N_30167);
or U49327 (N_49327,N_36866,N_33610);
nor U49328 (N_49328,N_38663,N_37333);
nand U49329 (N_49329,N_39047,N_39443);
or U49330 (N_49330,N_31993,N_30418);
nand U49331 (N_49331,N_37586,N_39922);
and U49332 (N_49332,N_32431,N_39527);
nor U49333 (N_49333,N_34669,N_39305);
or U49334 (N_49334,N_31760,N_35545);
xor U49335 (N_49335,N_32574,N_30661);
and U49336 (N_49336,N_36602,N_35428);
nor U49337 (N_49337,N_35027,N_34999);
xor U49338 (N_49338,N_37016,N_33109);
nor U49339 (N_49339,N_38045,N_30053);
nand U49340 (N_49340,N_30228,N_39050);
nor U49341 (N_49341,N_37598,N_33839);
nor U49342 (N_49342,N_32535,N_35528);
xnor U49343 (N_49343,N_36606,N_31615);
nand U49344 (N_49344,N_38974,N_31923);
and U49345 (N_49345,N_32070,N_30881);
or U49346 (N_49346,N_31779,N_32549);
or U49347 (N_49347,N_30443,N_36191);
or U49348 (N_49348,N_37992,N_34568);
nand U49349 (N_49349,N_31716,N_31372);
nor U49350 (N_49350,N_38109,N_32183);
nand U49351 (N_49351,N_33740,N_35322);
or U49352 (N_49352,N_31970,N_37523);
nor U49353 (N_49353,N_39070,N_31846);
nand U49354 (N_49354,N_35556,N_34189);
or U49355 (N_49355,N_38802,N_31635);
nor U49356 (N_49356,N_36758,N_30658);
nand U49357 (N_49357,N_35321,N_31406);
nand U49358 (N_49358,N_33210,N_31518);
xnor U49359 (N_49359,N_36568,N_33043);
or U49360 (N_49360,N_30033,N_30731);
nor U49361 (N_49361,N_32131,N_33503);
nand U49362 (N_49362,N_33943,N_32284);
or U49363 (N_49363,N_32709,N_34527);
xnor U49364 (N_49364,N_35620,N_31111);
xor U49365 (N_49365,N_33149,N_37331);
or U49366 (N_49366,N_33361,N_35307);
nand U49367 (N_49367,N_30933,N_38226);
or U49368 (N_49368,N_38957,N_38099);
and U49369 (N_49369,N_37867,N_30600);
xnor U49370 (N_49370,N_38262,N_36773);
xnor U49371 (N_49371,N_30940,N_35231);
xor U49372 (N_49372,N_37347,N_38136);
nand U49373 (N_49373,N_31869,N_31635);
xnor U49374 (N_49374,N_30051,N_32208);
xor U49375 (N_49375,N_31273,N_33498);
and U49376 (N_49376,N_34558,N_38691);
xnor U49377 (N_49377,N_32329,N_39164);
or U49378 (N_49378,N_36086,N_33792);
or U49379 (N_49379,N_34500,N_37735);
and U49380 (N_49380,N_30127,N_33449);
nor U49381 (N_49381,N_38947,N_37531);
nand U49382 (N_49382,N_36791,N_30637);
or U49383 (N_49383,N_36717,N_34451);
nor U49384 (N_49384,N_38306,N_37461);
and U49385 (N_49385,N_39476,N_38706);
nand U49386 (N_49386,N_31573,N_35848);
xor U49387 (N_49387,N_31803,N_36092);
nor U49388 (N_49388,N_38304,N_36545);
or U49389 (N_49389,N_37654,N_30609);
xor U49390 (N_49390,N_38228,N_30417);
and U49391 (N_49391,N_37513,N_38599);
nand U49392 (N_49392,N_30682,N_30421);
or U49393 (N_49393,N_31511,N_33363);
xnor U49394 (N_49394,N_35477,N_32089);
and U49395 (N_49395,N_34487,N_33035);
and U49396 (N_49396,N_37159,N_35205);
nand U49397 (N_49397,N_38609,N_39825);
nor U49398 (N_49398,N_30015,N_34861);
and U49399 (N_49399,N_36011,N_32561);
nand U49400 (N_49400,N_36270,N_35629);
nand U49401 (N_49401,N_39846,N_38585);
nor U49402 (N_49402,N_32472,N_31184);
nor U49403 (N_49403,N_35396,N_39677);
xnor U49404 (N_49404,N_38637,N_32957);
and U49405 (N_49405,N_31849,N_37526);
and U49406 (N_49406,N_34191,N_32855);
nand U49407 (N_49407,N_35894,N_36977);
nand U49408 (N_49408,N_31372,N_35537);
and U49409 (N_49409,N_35023,N_32209);
nor U49410 (N_49410,N_36098,N_37718);
nor U49411 (N_49411,N_38363,N_33925);
and U49412 (N_49412,N_37952,N_30334);
nand U49413 (N_49413,N_31771,N_30238);
xor U49414 (N_49414,N_31270,N_35451);
nand U49415 (N_49415,N_38601,N_37454);
and U49416 (N_49416,N_35083,N_38677);
xor U49417 (N_49417,N_39079,N_31064);
nand U49418 (N_49418,N_37018,N_32340);
nand U49419 (N_49419,N_35943,N_32668);
xnor U49420 (N_49420,N_31467,N_33400);
or U49421 (N_49421,N_37982,N_35887);
nand U49422 (N_49422,N_39418,N_35127);
xor U49423 (N_49423,N_31365,N_36031);
xor U49424 (N_49424,N_32158,N_35937);
and U49425 (N_49425,N_34798,N_35497);
nor U49426 (N_49426,N_39510,N_33056);
nand U49427 (N_49427,N_31375,N_31909);
and U49428 (N_49428,N_39196,N_32786);
and U49429 (N_49429,N_36591,N_31782);
and U49430 (N_49430,N_33484,N_32889);
or U49431 (N_49431,N_38656,N_38759);
nand U49432 (N_49432,N_30734,N_30856);
nor U49433 (N_49433,N_38208,N_34232);
and U49434 (N_49434,N_32036,N_38689);
nand U49435 (N_49435,N_35909,N_30411);
nor U49436 (N_49436,N_31482,N_39334);
nand U49437 (N_49437,N_33899,N_37813);
xnor U49438 (N_49438,N_37428,N_35493);
xnor U49439 (N_49439,N_39269,N_33816);
nand U49440 (N_49440,N_32453,N_37088);
nand U49441 (N_49441,N_39947,N_34038);
or U49442 (N_49442,N_34274,N_30665);
and U49443 (N_49443,N_35665,N_35291);
nor U49444 (N_49444,N_39196,N_39364);
nor U49445 (N_49445,N_33564,N_33340);
or U49446 (N_49446,N_33645,N_34351);
or U49447 (N_49447,N_37368,N_38941);
or U49448 (N_49448,N_31044,N_32429);
nor U49449 (N_49449,N_32390,N_37177);
xnor U49450 (N_49450,N_36284,N_37851);
xor U49451 (N_49451,N_30300,N_39499);
nand U49452 (N_49452,N_38275,N_39898);
and U49453 (N_49453,N_31362,N_30741);
xnor U49454 (N_49454,N_35897,N_30215);
nor U49455 (N_49455,N_30959,N_34733);
and U49456 (N_49456,N_30441,N_33292);
nor U49457 (N_49457,N_36367,N_39775);
or U49458 (N_49458,N_32126,N_38885);
or U49459 (N_49459,N_33470,N_32723);
and U49460 (N_49460,N_35137,N_39838);
and U49461 (N_49461,N_36644,N_37628);
xnor U49462 (N_49462,N_34920,N_31878);
xnor U49463 (N_49463,N_33983,N_37845);
or U49464 (N_49464,N_34341,N_34687);
xor U49465 (N_49465,N_34257,N_38231);
nand U49466 (N_49466,N_39805,N_30946);
xor U49467 (N_49467,N_37400,N_33763);
or U49468 (N_49468,N_38357,N_33281);
nor U49469 (N_49469,N_39465,N_35834);
and U49470 (N_49470,N_36074,N_34184);
or U49471 (N_49471,N_32501,N_36611);
or U49472 (N_49472,N_33438,N_38826);
or U49473 (N_49473,N_36976,N_33707);
or U49474 (N_49474,N_30592,N_35340);
nor U49475 (N_49475,N_35287,N_35741);
nor U49476 (N_49476,N_30496,N_32731);
xor U49477 (N_49477,N_38221,N_39082);
nor U49478 (N_49478,N_35425,N_33997);
nor U49479 (N_49479,N_39828,N_32536);
nor U49480 (N_49480,N_37457,N_37573);
and U49481 (N_49481,N_34585,N_31630);
and U49482 (N_49482,N_34005,N_39182);
or U49483 (N_49483,N_35298,N_32449);
nand U49484 (N_49484,N_33133,N_37548);
and U49485 (N_49485,N_30528,N_35128);
nand U49486 (N_49486,N_37747,N_31677);
xor U49487 (N_49487,N_33703,N_33828);
nand U49488 (N_49488,N_35018,N_36532);
xor U49489 (N_49489,N_36438,N_36851);
nand U49490 (N_49490,N_39858,N_35887);
nor U49491 (N_49491,N_31710,N_38597);
and U49492 (N_49492,N_31273,N_31084);
nand U49493 (N_49493,N_37491,N_33828);
nand U49494 (N_49494,N_35531,N_39197);
nor U49495 (N_49495,N_35588,N_35030);
xnor U49496 (N_49496,N_32376,N_39773);
nor U49497 (N_49497,N_37320,N_38792);
and U49498 (N_49498,N_37746,N_34747);
and U49499 (N_49499,N_32669,N_32474);
nand U49500 (N_49500,N_39892,N_33931);
nor U49501 (N_49501,N_30277,N_30390);
and U49502 (N_49502,N_35535,N_39183);
or U49503 (N_49503,N_36143,N_30649);
and U49504 (N_49504,N_32888,N_32027);
and U49505 (N_49505,N_30437,N_33063);
nand U49506 (N_49506,N_33545,N_30834);
or U49507 (N_49507,N_33646,N_39509);
nor U49508 (N_49508,N_30605,N_30969);
or U49509 (N_49509,N_31682,N_37508);
and U49510 (N_49510,N_33905,N_33835);
and U49511 (N_49511,N_36798,N_32447);
nand U49512 (N_49512,N_30711,N_30063);
xnor U49513 (N_49513,N_35338,N_37390);
xnor U49514 (N_49514,N_36633,N_35457);
and U49515 (N_49515,N_37709,N_39619);
nand U49516 (N_49516,N_39620,N_30959);
xor U49517 (N_49517,N_34663,N_30198);
or U49518 (N_49518,N_35242,N_37858);
nor U49519 (N_49519,N_35278,N_39793);
nand U49520 (N_49520,N_30737,N_35047);
or U49521 (N_49521,N_36086,N_38073);
nor U49522 (N_49522,N_30009,N_37249);
or U49523 (N_49523,N_30746,N_31329);
nand U49524 (N_49524,N_39383,N_33349);
xnor U49525 (N_49525,N_38799,N_39522);
xnor U49526 (N_49526,N_33489,N_37585);
and U49527 (N_49527,N_36611,N_39376);
or U49528 (N_49528,N_37683,N_36924);
nand U49529 (N_49529,N_38322,N_34878);
xor U49530 (N_49530,N_37441,N_39059);
nand U49531 (N_49531,N_35067,N_34124);
xor U49532 (N_49532,N_39168,N_34852);
or U49533 (N_49533,N_32547,N_35281);
xor U49534 (N_49534,N_38815,N_36466);
and U49535 (N_49535,N_39727,N_32297);
nand U49536 (N_49536,N_34686,N_37136);
or U49537 (N_49537,N_34519,N_39178);
xor U49538 (N_49538,N_32961,N_33463);
and U49539 (N_49539,N_30753,N_30349);
and U49540 (N_49540,N_39475,N_36911);
xnor U49541 (N_49541,N_33264,N_35902);
and U49542 (N_49542,N_35133,N_36482);
and U49543 (N_49543,N_30355,N_39987);
nand U49544 (N_49544,N_30113,N_34787);
nor U49545 (N_49545,N_36704,N_35109);
and U49546 (N_49546,N_32822,N_31213);
nor U49547 (N_49547,N_39785,N_38990);
or U49548 (N_49548,N_37905,N_32730);
nor U49549 (N_49549,N_34500,N_37691);
nor U49550 (N_49550,N_38642,N_32063);
nand U49551 (N_49551,N_38293,N_31183);
nor U49552 (N_49552,N_37824,N_34815);
nor U49553 (N_49553,N_34545,N_37701);
xor U49554 (N_49554,N_39050,N_36373);
xnor U49555 (N_49555,N_39571,N_39426);
xnor U49556 (N_49556,N_38370,N_32970);
xor U49557 (N_49557,N_35881,N_38762);
nor U49558 (N_49558,N_30008,N_31991);
xnor U49559 (N_49559,N_39645,N_34286);
nand U49560 (N_49560,N_38870,N_36468);
xnor U49561 (N_49561,N_36108,N_38893);
nand U49562 (N_49562,N_36917,N_39088);
nand U49563 (N_49563,N_33862,N_32871);
nor U49564 (N_49564,N_32259,N_39370);
and U49565 (N_49565,N_34329,N_34410);
xnor U49566 (N_49566,N_38490,N_36471);
nor U49567 (N_49567,N_39206,N_39652);
and U49568 (N_49568,N_38685,N_36394);
or U49569 (N_49569,N_31690,N_31600);
or U49570 (N_49570,N_38242,N_35512);
xnor U49571 (N_49571,N_33174,N_32422);
and U49572 (N_49572,N_36322,N_38460);
and U49573 (N_49573,N_36230,N_31940);
and U49574 (N_49574,N_39476,N_36857);
and U49575 (N_49575,N_35319,N_36574);
nor U49576 (N_49576,N_30386,N_31659);
nor U49577 (N_49577,N_37716,N_38458);
and U49578 (N_49578,N_34007,N_38038);
nor U49579 (N_49579,N_33144,N_38176);
nor U49580 (N_49580,N_39071,N_33213);
nand U49581 (N_49581,N_31838,N_37720);
nor U49582 (N_49582,N_31345,N_37026);
or U49583 (N_49583,N_35274,N_32966);
or U49584 (N_49584,N_35606,N_32279);
xor U49585 (N_49585,N_35673,N_35008);
nor U49586 (N_49586,N_31168,N_32519);
and U49587 (N_49587,N_30673,N_39776);
and U49588 (N_49588,N_31675,N_32275);
xnor U49589 (N_49589,N_34962,N_38829);
xor U49590 (N_49590,N_35046,N_37603);
or U49591 (N_49591,N_36830,N_32806);
nor U49592 (N_49592,N_31514,N_30875);
nor U49593 (N_49593,N_32908,N_33211);
and U49594 (N_49594,N_34165,N_36821);
nor U49595 (N_49595,N_31644,N_31824);
xor U49596 (N_49596,N_38230,N_31078);
and U49597 (N_49597,N_39824,N_39187);
or U49598 (N_49598,N_38976,N_30861);
xor U49599 (N_49599,N_36070,N_37223);
xor U49600 (N_49600,N_35287,N_30239);
nor U49601 (N_49601,N_32422,N_37753);
or U49602 (N_49602,N_32039,N_33976);
or U49603 (N_49603,N_31610,N_31896);
nand U49604 (N_49604,N_39342,N_38431);
or U49605 (N_49605,N_39591,N_36955);
nor U49606 (N_49606,N_30856,N_37756);
xor U49607 (N_49607,N_30063,N_38491);
and U49608 (N_49608,N_34010,N_35660);
nand U49609 (N_49609,N_34016,N_33376);
and U49610 (N_49610,N_31477,N_38581);
nand U49611 (N_49611,N_33702,N_37398);
and U49612 (N_49612,N_30948,N_38318);
and U49613 (N_49613,N_34679,N_34134);
nor U49614 (N_49614,N_39685,N_34596);
or U49615 (N_49615,N_35847,N_39682);
xnor U49616 (N_49616,N_33151,N_33073);
or U49617 (N_49617,N_38979,N_36595);
or U49618 (N_49618,N_30310,N_31294);
and U49619 (N_49619,N_35169,N_34469);
and U49620 (N_49620,N_35764,N_30820);
xor U49621 (N_49621,N_31179,N_38732);
xnor U49622 (N_49622,N_36931,N_36063);
xor U49623 (N_49623,N_37804,N_31881);
and U49624 (N_49624,N_31240,N_35192);
nor U49625 (N_49625,N_36048,N_31246);
nor U49626 (N_49626,N_30576,N_30604);
nor U49627 (N_49627,N_34245,N_35076);
nor U49628 (N_49628,N_35326,N_33977);
or U49629 (N_49629,N_37817,N_32785);
or U49630 (N_49630,N_31902,N_39238);
or U49631 (N_49631,N_34014,N_36120);
or U49632 (N_49632,N_30905,N_35383);
nand U49633 (N_49633,N_35033,N_30830);
nor U49634 (N_49634,N_32957,N_33242);
or U49635 (N_49635,N_31242,N_38411);
nor U49636 (N_49636,N_36420,N_30907);
or U49637 (N_49637,N_32220,N_31391);
and U49638 (N_49638,N_34582,N_37792);
xor U49639 (N_49639,N_35718,N_35133);
xor U49640 (N_49640,N_32746,N_39817);
nor U49641 (N_49641,N_34485,N_31434);
nor U49642 (N_49642,N_36930,N_36401);
and U49643 (N_49643,N_33040,N_34651);
and U49644 (N_49644,N_30357,N_31078);
and U49645 (N_49645,N_30096,N_34238);
nand U49646 (N_49646,N_39118,N_31563);
nor U49647 (N_49647,N_34007,N_36268);
nand U49648 (N_49648,N_33011,N_38358);
or U49649 (N_49649,N_38196,N_30782);
and U49650 (N_49650,N_33654,N_39612);
or U49651 (N_49651,N_31205,N_37423);
nand U49652 (N_49652,N_30093,N_31767);
xnor U49653 (N_49653,N_37931,N_32408);
xnor U49654 (N_49654,N_39366,N_38218);
nand U49655 (N_49655,N_37516,N_33836);
nand U49656 (N_49656,N_30294,N_35058);
nand U49657 (N_49657,N_33811,N_36626);
xnor U49658 (N_49658,N_33238,N_30356);
or U49659 (N_49659,N_31224,N_39302);
nand U49660 (N_49660,N_35684,N_36427);
and U49661 (N_49661,N_34432,N_37707);
xor U49662 (N_49662,N_33861,N_33851);
xnor U49663 (N_49663,N_36727,N_31689);
nor U49664 (N_49664,N_38566,N_38252);
xor U49665 (N_49665,N_30531,N_32300);
and U49666 (N_49666,N_39076,N_33091);
xnor U49667 (N_49667,N_36592,N_38633);
nor U49668 (N_49668,N_38252,N_33127);
and U49669 (N_49669,N_30042,N_38804);
nor U49670 (N_49670,N_30298,N_32073);
nand U49671 (N_49671,N_38561,N_33462);
xor U49672 (N_49672,N_38391,N_39909);
nor U49673 (N_49673,N_34975,N_34449);
and U49674 (N_49674,N_35069,N_39948);
nor U49675 (N_49675,N_34190,N_34797);
or U49676 (N_49676,N_30227,N_34017);
xor U49677 (N_49677,N_34724,N_31320);
nand U49678 (N_49678,N_35852,N_32269);
nand U49679 (N_49679,N_37855,N_36173);
nand U49680 (N_49680,N_39376,N_32012);
nor U49681 (N_49681,N_32379,N_32647);
nand U49682 (N_49682,N_35874,N_34026);
nand U49683 (N_49683,N_31179,N_36252);
nor U49684 (N_49684,N_39729,N_31203);
nor U49685 (N_49685,N_30576,N_38516);
or U49686 (N_49686,N_30402,N_37828);
and U49687 (N_49687,N_35626,N_36609);
and U49688 (N_49688,N_33192,N_37385);
or U49689 (N_49689,N_37904,N_32542);
and U49690 (N_49690,N_39189,N_32472);
nand U49691 (N_49691,N_39072,N_38168);
nand U49692 (N_49692,N_31792,N_36325);
nor U49693 (N_49693,N_35420,N_37883);
xnor U49694 (N_49694,N_39143,N_37906);
nor U49695 (N_49695,N_34531,N_31377);
and U49696 (N_49696,N_35770,N_30553);
nand U49697 (N_49697,N_32695,N_38455);
or U49698 (N_49698,N_33074,N_30608);
xor U49699 (N_49699,N_35978,N_38609);
nand U49700 (N_49700,N_37735,N_38299);
nand U49701 (N_49701,N_30849,N_33637);
xnor U49702 (N_49702,N_39548,N_37708);
nand U49703 (N_49703,N_35294,N_34767);
nand U49704 (N_49704,N_30855,N_37069);
nor U49705 (N_49705,N_38415,N_38427);
nand U49706 (N_49706,N_39180,N_38654);
or U49707 (N_49707,N_35927,N_32184);
or U49708 (N_49708,N_39297,N_37888);
nand U49709 (N_49709,N_31987,N_31986);
xor U49710 (N_49710,N_30638,N_32989);
xnor U49711 (N_49711,N_34138,N_35224);
or U49712 (N_49712,N_37145,N_36934);
and U49713 (N_49713,N_34637,N_32235);
xnor U49714 (N_49714,N_36217,N_38343);
or U49715 (N_49715,N_39295,N_30952);
nand U49716 (N_49716,N_31905,N_36350);
and U49717 (N_49717,N_30501,N_35791);
or U49718 (N_49718,N_30813,N_33272);
xor U49719 (N_49719,N_34523,N_34225);
nand U49720 (N_49720,N_32192,N_34283);
xnor U49721 (N_49721,N_37623,N_38276);
and U49722 (N_49722,N_33908,N_38831);
and U49723 (N_49723,N_30149,N_34249);
nand U49724 (N_49724,N_35867,N_32337);
or U49725 (N_49725,N_37472,N_33233);
nand U49726 (N_49726,N_31124,N_37120);
or U49727 (N_49727,N_31877,N_31283);
nand U49728 (N_49728,N_31274,N_36112);
nor U49729 (N_49729,N_33106,N_33968);
nor U49730 (N_49730,N_33971,N_38783);
xor U49731 (N_49731,N_38263,N_38247);
xor U49732 (N_49732,N_30360,N_30952);
nor U49733 (N_49733,N_30801,N_32001);
and U49734 (N_49734,N_32544,N_33251);
nand U49735 (N_49735,N_35546,N_33936);
xor U49736 (N_49736,N_33498,N_32731);
and U49737 (N_49737,N_39995,N_35783);
nand U49738 (N_49738,N_32288,N_37934);
nor U49739 (N_49739,N_34218,N_38146);
nand U49740 (N_49740,N_35344,N_36129);
nor U49741 (N_49741,N_33370,N_31052);
or U49742 (N_49742,N_31186,N_33079);
or U49743 (N_49743,N_34869,N_31473);
xnor U49744 (N_49744,N_36257,N_39988);
nand U49745 (N_49745,N_38195,N_38488);
or U49746 (N_49746,N_35713,N_36537);
or U49747 (N_49747,N_36063,N_37557);
or U49748 (N_49748,N_31787,N_32097);
nor U49749 (N_49749,N_36774,N_34041);
or U49750 (N_49750,N_35644,N_39462);
or U49751 (N_49751,N_39120,N_37531);
and U49752 (N_49752,N_32164,N_37866);
nor U49753 (N_49753,N_37295,N_39328);
and U49754 (N_49754,N_33500,N_36632);
and U49755 (N_49755,N_39771,N_35672);
nor U49756 (N_49756,N_30133,N_31504);
and U49757 (N_49757,N_36482,N_30169);
nor U49758 (N_49758,N_37397,N_38360);
nor U49759 (N_49759,N_32254,N_30170);
xnor U49760 (N_49760,N_34070,N_35355);
and U49761 (N_49761,N_37834,N_33828);
and U49762 (N_49762,N_36488,N_33815);
nand U49763 (N_49763,N_33963,N_37669);
and U49764 (N_49764,N_33006,N_35368);
xnor U49765 (N_49765,N_39904,N_37879);
nor U49766 (N_49766,N_37765,N_32518);
and U49767 (N_49767,N_35856,N_38569);
xnor U49768 (N_49768,N_33729,N_34839);
nand U49769 (N_49769,N_35783,N_37771);
or U49770 (N_49770,N_34256,N_38537);
or U49771 (N_49771,N_32302,N_39390);
or U49772 (N_49772,N_38620,N_31240);
xor U49773 (N_49773,N_37852,N_34145);
and U49774 (N_49774,N_31804,N_39824);
and U49775 (N_49775,N_36221,N_32574);
or U49776 (N_49776,N_38184,N_30459);
and U49777 (N_49777,N_34180,N_30527);
and U49778 (N_49778,N_37106,N_34078);
nor U49779 (N_49779,N_32799,N_30255);
nor U49780 (N_49780,N_34899,N_39531);
or U49781 (N_49781,N_36474,N_30336);
and U49782 (N_49782,N_36138,N_37423);
nand U49783 (N_49783,N_38730,N_38804);
nand U49784 (N_49784,N_31648,N_31294);
nor U49785 (N_49785,N_30407,N_39647);
nand U49786 (N_49786,N_33143,N_31505);
nor U49787 (N_49787,N_38790,N_30447);
nor U49788 (N_49788,N_30144,N_30838);
nor U49789 (N_49789,N_34644,N_36473);
or U49790 (N_49790,N_37565,N_34554);
nand U49791 (N_49791,N_35694,N_34695);
nor U49792 (N_49792,N_31440,N_32476);
nand U49793 (N_49793,N_36308,N_32719);
and U49794 (N_49794,N_37994,N_31311);
nand U49795 (N_49795,N_39667,N_35059);
or U49796 (N_49796,N_36196,N_35229);
nand U49797 (N_49797,N_36946,N_31716);
xor U49798 (N_49798,N_34808,N_39818);
nand U49799 (N_49799,N_34218,N_32389);
or U49800 (N_49800,N_31324,N_35883);
nand U49801 (N_49801,N_30900,N_30432);
and U49802 (N_49802,N_34725,N_32940);
or U49803 (N_49803,N_33808,N_34867);
nand U49804 (N_49804,N_34738,N_34532);
and U49805 (N_49805,N_39710,N_31351);
xor U49806 (N_49806,N_36327,N_38802);
nor U49807 (N_49807,N_32233,N_32231);
and U49808 (N_49808,N_37549,N_34778);
xnor U49809 (N_49809,N_34313,N_32679);
and U49810 (N_49810,N_35680,N_35143);
xnor U49811 (N_49811,N_31463,N_36001);
xnor U49812 (N_49812,N_30863,N_31636);
nand U49813 (N_49813,N_30067,N_38065);
or U49814 (N_49814,N_31363,N_37974);
and U49815 (N_49815,N_32292,N_31452);
nand U49816 (N_49816,N_35211,N_39730);
or U49817 (N_49817,N_30135,N_32774);
xor U49818 (N_49818,N_39787,N_30706);
nor U49819 (N_49819,N_39519,N_30328);
nand U49820 (N_49820,N_38477,N_36190);
nor U49821 (N_49821,N_34536,N_39851);
and U49822 (N_49822,N_35591,N_32863);
nand U49823 (N_49823,N_31524,N_37777);
nor U49824 (N_49824,N_39317,N_37546);
and U49825 (N_49825,N_35570,N_35967);
or U49826 (N_49826,N_31880,N_38329);
nor U49827 (N_49827,N_30964,N_37904);
xnor U49828 (N_49828,N_32199,N_34137);
or U49829 (N_49829,N_30798,N_37878);
and U49830 (N_49830,N_32910,N_31659);
and U49831 (N_49831,N_39471,N_36812);
nand U49832 (N_49832,N_35786,N_33079);
xnor U49833 (N_49833,N_36284,N_37432);
and U49834 (N_49834,N_33027,N_38843);
nor U49835 (N_49835,N_34982,N_37147);
and U49836 (N_49836,N_38260,N_35423);
or U49837 (N_49837,N_37604,N_36724);
or U49838 (N_49838,N_31988,N_33298);
or U49839 (N_49839,N_37311,N_34738);
and U49840 (N_49840,N_34264,N_36149);
and U49841 (N_49841,N_39464,N_31961);
nand U49842 (N_49842,N_38648,N_37843);
or U49843 (N_49843,N_38420,N_33388);
nand U49844 (N_49844,N_37836,N_34385);
or U49845 (N_49845,N_38789,N_30199);
nor U49846 (N_49846,N_38548,N_30213);
xor U49847 (N_49847,N_31309,N_39259);
and U49848 (N_49848,N_33244,N_39439);
nor U49849 (N_49849,N_38073,N_35217);
nand U49850 (N_49850,N_37895,N_37293);
and U49851 (N_49851,N_32396,N_39259);
or U49852 (N_49852,N_39420,N_33016);
nor U49853 (N_49853,N_30511,N_38130);
xnor U49854 (N_49854,N_37235,N_33145);
xnor U49855 (N_49855,N_32887,N_33131);
nor U49856 (N_49856,N_30794,N_32183);
and U49857 (N_49857,N_36253,N_39699);
or U49858 (N_49858,N_31891,N_31758);
or U49859 (N_49859,N_32909,N_32658);
nand U49860 (N_49860,N_38808,N_39712);
or U49861 (N_49861,N_39606,N_39288);
xor U49862 (N_49862,N_38264,N_35395);
nand U49863 (N_49863,N_34336,N_39218);
and U49864 (N_49864,N_33385,N_38683);
xnor U49865 (N_49865,N_30045,N_35700);
xnor U49866 (N_49866,N_38996,N_33835);
and U49867 (N_49867,N_38443,N_33190);
xnor U49868 (N_49868,N_30882,N_30935);
xor U49869 (N_49869,N_35850,N_39814);
nor U49870 (N_49870,N_32722,N_33845);
nand U49871 (N_49871,N_35083,N_35742);
nor U49872 (N_49872,N_32368,N_38031);
nand U49873 (N_49873,N_32640,N_39800);
nand U49874 (N_49874,N_33261,N_35306);
nor U49875 (N_49875,N_39646,N_30966);
and U49876 (N_49876,N_33350,N_32430);
or U49877 (N_49877,N_30034,N_39987);
or U49878 (N_49878,N_31204,N_38744);
nor U49879 (N_49879,N_33105,N_35713);
and U49880 (N_49880,N_37308,N_39379);
xnor U49881 (N_49881,N_38921,N_31806);
nand U49882 (N_49882,N_31617,N_38799);
nand U49883 (N_49883,N_39143,N_36148);
nor U49884 (N_49884,N_33309,N_34016);
and U49885 (N_49885,N_32344,N_36675);
xor U49886 (N_49886,N_33287,N_37481);
and U49887 (N_49887,N_35899,N_31326);
nor U49888 (N_49888,N_36768,N_38993);
nand U49889 (N_49889,N_35664,N_31547);
xor U49890 (N_49890,N_33634,N_33305);
xor U49891 (N_49891,N_37565,N_33904);
or U49892 (N_49892,N_30648,N_38349);
xor U49893 (N_49893,N_35507,N_34396);
xor U49894 (N_49894,N_34209,N_36957);
xor U49895 (N_49895,N_33325,N_33182);
nand U49896 (N_49896,N_36195,N_37261);
and U49897 (N_49897,N_34262,N_33419);
or U49898 (N_49898,N_37765,N_30927);
nand U49899 (N_49899,N_33888,N_30477);
nor U49900 (N_49900,N_30597,N_36201);
and U49901 (N_49901,N_34451,N_30445);
nand U49902 (N_49902,N_36060,N_36208);
and U49903 (N_49903,N_34787,N_39972);
or U49904 (N_49904,N_38116,N_30016);
or U49905 (N_49905,N_36896,N_35793);
nand U49906 (N_49906,N_31959,N_31749);
nor U49907 (N_49907,N_33703,N_36856);
nor U49908 (N_49908,N_39462,N_35000);
and U49909 (N_49909,N_34938,N_34591);
and U49910 (N_49910,N_30230,N_34156);
or U49911 (N_49911,N_39156,N_37648);
xnor U49912 (N_49912,N_33739,N_34908);
or U49913 (N_49913,N_34902,N_32717);
and U49914 (N_49914,N_33681,N_38641);
nor U49915 (N_49915,N_36293,N_32561);
xor U49916 (N_49916,N_37528,N_38913);
nor U49917 (N_49917,N_38983,N_31503);
nand U49918 (N_49918,N_31275,N_31780);
xnor U49919 (N_49919,N_32167,N_38986);
nor U49920 (N_49920,N_34723,N_31963);
nand U49921 (N_49921,N_36355,N_37344);
or U49922 (N_49922,N_35299,N_31037);
nand U49923 (N_49923,N_34034,N_33040);
or U49924 (N_49924,N_39463,N_39197);
nor U49925 (N_49925,N_35727,N_37915);
or U49926 (N_49926,N_38304,N_36732);
nor U49927 (N_49927,N_37217,N_33355);
and U49928 (N_49928,N_34900,N_39985);
nand U49929 (N_49929,N_38363,N_38603);
nand U49930 (N_49930,N_36797,N_35131);
nor U49931 (N_49931,N_30647,N_38720);
nor U49932 (N_49932,N_30448,N_33710);
or U49933 (N_49933,N_39671,N_39098);
or U49934 (N_49934,N_33528,N_39783);
nand U49935 (N_49935,N_38889,N_36283);
xnor U49936 (N_49936,N_37377,N_37566);
xor U49937 (N_49937,N_31985,N_39255);
nor U49938 (N_49938,N_38627,N_33183);
nor U49939 (N_49939,N_30142,N_37183);
nand U49940 (N_49940,N_32622,N_36984);
nor U49941 (N_49941,N_35980,N_38230);
nor U49942 (N_49942,N_33001,N_39461);
or U49943 (N_49943,N_31986,N_37766);
xnor U49944 (N_49944,N_34735,N_38117);
or U49945 (N_49945,N_32551,N_34248);
or U49946 (N_49946,N_31834,N_30410);
or U49947 (N_49947,N_30307,N_38244);
nor U49948 (N_49948,N_38505,N_35649);
and U49949 (N_49949,N_38659,N_36452);
nor U49950 (N_49950,N_34379,N_36625);
and U49951 (N_49951,N_38010,N_32297);
nand U49952 (N_49952,N_34472,N_34695);
nor U49953 (N_49953,N_34049,N_34987);
and U49954 (N_49954,N_38511,N_38621);
xor U49955 (N_49955,N_33012,N_32990);
nand U49956 (N_49956,N_30952,N_35834);
and U49957 (N_49957,N_30986,N_34314);
and U49958 (N_49958,N_36671,N_35590);
nor U49959 (N_49959,N_34796,N_38312);
xor U49960 (N_49960,N_32167,N_32796);
and U49961 (N_49961,N_38531,N_35667);
and U49962 (N_49962,N_39578,N_35123);
nand U49963 (N_49963,N_38002,N_38245);
xnor U49964 (N_49964,N_32651,N_36929);
nor U49965 (N_49965,N_34806,N_36160);
nand U49966 (N_49966,N_34684,N_34531);
xnor U49967 (N_49967,N_34112,N_36013);
xor U49968 (N_49968,N_32880,N_33260);
or U49969 (N_49969,N_35274,N_36540);
nand U49970 (N_49970,N_31209,N_38686);
nand U49971 (N_49971,N_38611,N_35501);
or U49972 (N_49972,N_32863,N_31843);
nand U49973 (N_49973,N_34364,N_34165);
nor U49974 (N_49974,N_37517,N_39967);
and U49975 (N_49975,N_31373,N_39661);
or U49976 (N_49976,N_30959,N_33142);
nand U49977 (N_49977,N_39811,N_31819);
nor U49978 (N_49978,N_33882,N_35720);
xor U49979 (N_49979,N_39069,N_31254);
xnor U49980 (N_49980,N_35255,N_34929);
and U49981 (N_49981,N_30747,N_32299);
and U49982 (N_49982,N_36341,N_34564);
nor U49983 (N_49983,N_33246,N_36955);
or U49984 (N_49984,N_37818,N_36082);
and U49985 (N_49985,N_31780,N_39802);
or U49986 (N_49986,N_34325,N_39344);
nor U49987 (N_49987,N_35671,N_34024);
nor U49988 (N_49988,N_36473,N_39610);
nand U49989 (N_49989,N_35405,N_35170);
or U49990 (N_49990,N_34687,N_30447);
and U49991 (N_49991,N_31515,N_34434);
or U49992 (N_49992,N_39716,N_35265);
or U49993 (N_49993,N_34175,N_35531);
or U49994 (N_49994,N_31387,N_34566);
nand U49995 (N_49995,N_37517,N_31952);
or U49996 (N_49996,N_34133,N_35121);
and U49997 (N_49997,N_30599,N_30309);
xnor U49998 (N_49998,N_38123,N_32599);
or U49999 (N_49999,N_37350,N_33125);
and UO_0 (O_0,N_42185,N_44829);
nand UO_1 (O_1,N_45108,N_45200);
nand UO_2 (O_2,N_49555,N_44265);
nor UO_3 (O_3,N_45677,N_44160);
nor UO_4 (O_4,N_42201,N_41137);
and UO_5 (O_5,N_47856,N_45403);
or UO_6 (O_6,N_41818,N_49273);
nand UO_7 (O_7,N_45850,N_41432);
and UO_8 (O_8,N_45229,N_41391);
nor UO_9 (O_9,N_47202,N_43707);
nor UO_10 (O_10,N_41332,N_40010);
and UO_11 (O_11,N_49300,N_42147);
nor UO_12 (O_12,N_45139,N_47878);
nand UO_13 (O_13,N_46543,N_48140);
xor UO_14 (O_14,N_48161,N_48154);
or UO_15 (O_15,N_44225,N_42047);
nor UO_16 (O_16,N_48131,N_40274);
xor UO_17 (O_17,N_40147,N_49079);
nor UO_18 (O_18,N_46961,N_40177);
nand UO_19 (O_19,N_41773,N_40815);
nand UO_20 (O_20,N_46880,N_49285);
or UO_21 (O_21,N_46762,N_45664);
xnor UO_22 (O_22,N_45797,N_44579);
or UO_23 (O_23,N_43923,N_40121);
xnor UO_24 (O_24,N_43389,N_47982);
nand UO_25 (O_25,N_42847,N_46559);
nor UO_26 (O_26,N_40375,N_40912);
nand UO_27 (O_27,N_48319,N_43507);
xnor UO_28 (O_28,N_45806,N_49157);
nor UO_29 (O_29,N_49679,N_46286);
nor UO_30 (O_30,N_46500,N_48500);
nor UO_31 (O_31,N_47454,N_42187);
nand UO_32 (O_32,N_44589,N_45918);
and UO_33 (O_33,N_48861,N_46003);
nand UO_34 (O_34,N_44112,N_41995);
nor UO_35 (O_35,N_45774,N_42693);
xor UO_36 (O_36,N_41881,N_49419);
or UO_37 (O_37,N_47865,N_48942);
and UO_38 (O_38,N_47297,N_41823);
nor UO_39 (O_39,N_45451,N_46677);
nand UO_40 (O_40,N_41839,N_44753);
or UO_41 (O_41,N_47668,N_47497);
and UO_42 (O_42,N_42261,N_40405);
nand UO_43 (O_43,N_42453,N_45932);
nand UO_44 (O_44,N_42610,N_49210);
or UO_45 (O_45,N_41403,N_49714);
nand UO_46 (O_46,N_45743,N_42461);
nand UO_47 (O_47,N_43444,N_44202);
xnor UO_48 (O_48,N_43855,N_44405);
or UO_49 (O_49,N_41087,N_43877);
nor UO_50 (O_50,N_44518,N_42068);
nor UO_51 (O_51,N_43416,N_46467);
nor UO_52 (O_52,N_44000,N_44923);
xor UO_53 (O_53,N_49667,N_48599);
and UO_54 (O_54,N_47830,N_47937);
nand UO_55 (O_55,N_49970,N_44971);
xor UO_56 (O_56,N_47310,N_44972);
nor UO_57 (O_57,N_40792,N_44892);
and UO_58 (O_58,N_42036,N_47406);
nand UO_59 (O_59,N_44625,N_44844);
and UO_60 (O_60,N_49546,N_47492);
and UO_61 (O_61,N_43465,N_49299);
xnor UO_62 (O_62,N_48177,N_41015);
nand UO_63 (O_63,N_48116,N_42286);
and UO_64 (O_64,N_49003,N_43794);
nand UO_65 (O_65,N_46679,N_46618);
nand UO_66 (O_66,N_43652,N_43278);
nand UO_67 (O_67,N_44904,N_48582);
nand UO_68 (O_68,N_42938,N_46183);
and UO_69 (O_69,N_40066,N_41366);
nor UO_70 (O_70,N_49090,N_44024);
and UO_71 (O_71,N_47203,N_48504);
and UO_72 (O_72,N_43271,N_43384);
xnor UO_73 (O_73,N_41780,N_46774);
or UO_74 (O_74,N_48538,N_49486);
or UO_75 (O_75,N_45911,N_41861);
or UO_76 (O_76,N_46941,N_42942);
or UO_77 (O_77,N_48743,N_45304);
xor UO_78 (O_78,N_46840,N_47796);
nor UO_79 (O_79,N_45579,N_41052);
nor UO_80 (O_80,N_46477,N_42849);
or UO_81 (O_81,N_43590,N_49183);
or UO_82 (O_82,N_45776,N_48361);
and UO_83 (O_83,N_41478,N_41836);
or UO_84 (O_84,N_45129,N_44268);
and UO_85 (O_85,N_45880,N_42781);
or UO_86 (O_86,N_45433,N_41518);
xnor UO_87 (O_87,N_49883,N_42476);
or UO_88 (O_88,N_41098,N_49496);
xnor UO_89 (O_89,N_44436,N_49902);
xor UO_90 (O_90,N_43928,N_44184);
nor UO_91 (O_91,N_48239,N_48844);
nand UO_92 (O_92,N_45699,N_45436);
nor UO_93 (O_93,N_49089,N_42298);
and UO_94 (O_94,N_49246,N_44033);
and UO_95 (O_95,N_48093,N_44280);
nand UO_96 (O_96,N_47321,N_42128);
or UO_97 (O_97,N_45900,N_45808);
nor UO_98 (O_98,N_44164,N_43025);
or UO_99 (O_99,N_41146,N_44679);
or UO_100 (O_100,N_46140,N_46891);
nor UO_101 (O_101,N_44963,N_43312);
and UO_102 (O_102,N_46918,N_40252);
nor UO_103 (O_103,N_44951,N_42957);
nor UO_104 (O_104,N_46560,N_40917);
nor UO_105 (O_105,N_45987,N_49729);
or UO_106 (O_106,N_43948,N_47393);
nand UO_107 (O_107,N_42734,N_45870);
or UO_108 (O_108,N_48581,N_47994);
or UO_109 (O_109,N_45319,N_46201);
and UO_110 (O_110,N_41447,N_48685);
and UO_111 (O_111,N_42940,N_46624);
xnor UO_112 (O_112,N_49848,N_43508);
xnor UO_113 (O_113,N_47315,N_40080);
nor UO_114 (O_114,N_46521,N_41126);
nand UO_115 (O_115,N_44135,N_42794);
nand UO_116 (O_116,N_45629,N_41103);
nor UO_117 (O_117,N_49207,N_43138);
xor UO_118 (O_118,N_47400,N_46110);
nand UO_119 (O_119,N_48781,N_46928);
and UO_120 (O_120,N_41690,N_41916);
nor UO_121 (O_121,N_42835,N_41212);
and UO_122 (O_122,N_43662,N_43127);
nor UO_123 (O_123,N_41525,N_49776);
and UO_124 (O_124,N_48086,N_46851);
and UO_125 (O_125,N_43920,N_42104);
nand UO_126 (O_126,N_42926,N_40836);
or UO_127 (O_127,N_43400,N_45786);
and UO_128 (O_128,N_45829,N_48021);
or UO_129 (O_129,N_43167,N_45038);
xor UO_130 (O_130,N_47291,N_49825);
or UO_131 (O_131,N_49125,N_47008);
or UO_132 (O_132,N_45135,N_45177);
nand UO_133 (O_133,N_43449,N_43204);
nor UO_134 (O_134,N_43496,N_40773);
xnor UO_135 (O_135,N_48334,N_49915);
nor UO_136 (O_136,N_44221,N_49863);
nor UO_137 (O_137,N_46220,N_49209);
xnor UO_138 (O_138,N_47598,N_40366);
nor UO_139 (O_139,N_47739,N_42810);
xnor UO_140 (O_140,N_40119,N_48918);
and UO_141 (O_141,N_42801,N_47069);
xor UO_142 (O_142,N_45744,N_42554);
nor UO_143 (O_143,N_41461,N_44715);
and UO_144 (O_144,N_44794,N_43348);
nor UO_145 (O_145,N_45551,N_41265);
and UO_146 (O_146,N_43876,N_48986);
or UO_147 (O_147,N_45198,N_44684);
nand UO_148 (O_148,N_48237,N_44100);
nor UO_149 (O_149,N_46645,N_43874);
xnor UO_150 (O_150,N_48422,N_42115);
or UO_151 (O_151,N_48243,N_48812);
nor UO_152 (O_152,N_42339,N_48231);
nor UO_153 (O_153,N_46044,N_48993);
or UO_154 (O_154,N_40873,N_45312);
nor UO_155 (O_155,N_41236,N_42851);
nand UO_156 (O_156,N_49898,N_49931);
nand UO_157 (O_157,N_46612,N_44620);
nand UO_158 (O_158,N_42325,N_47430);
nor UO_159 (O_159,N_46969,N_44352);
or UO_160 (O_160,N_47952,N_42609);
nor UO_161 (O_161,N_42795,N_49531);
nand UO_162 (O_162,N_49893,N_44658);
xnor UO_163 (O_163,N_44647,N_48998);
xor UO_164 (O_164,N_48805,N_44549);
xor UO_165 (O_165,N_43749,N_48146);
or UO_166 (O_166,N_42925,N_49618);
or UO_167 (O_167,N_45514,N_43474);
nor UO_168 (O_168,N_49591,N_49073);
and UO_169 (O_169,N_47740,N_48145);
nor UO_170 (O_170,N_40886,N_46086);
or UO_171 (O_171,N_41941,N_41563);
xor UO_172 (O_172,N_48734,N_42401);
xnor UO_173 (O_173,N_45573,N_49118);
nor UO_174 (O_174,N_43976,N_46253);
and UO_175 (O_175,N_48497,N_49055);
xnor UO_176 (O_176,N_45442,N_46692);
nor UO_177 (O_177,N_49117,N_45054);
and UO_178 (O_178,N_40860,N_44609);
nand UO_179 (O_179,N_43060,N_46799);
and UO_180 (O_180,N_40790,N_42805);
nor UO_181 (O_181,N_44199,N_43762);
nor UO_182 (O_182,N_47450,N_41040);
and UO_183 (O_183,N_44596,N_43269);
nor UO_184 (O_184,N_42907,N_41049);
or UO_185 (O_185,N_40441,N_41777);
and UO_186 (O_186,N_42216,N_47344);
xor UO_187 (O_187,N_49065,N_42330);
nand UO_188 (O_188,N_41646,N_45990);
and UO_189 (O_189,N_44755,N_47829);
nor UO_190 (O_190,N_40734,N_48573);
nand UO_191 (O_191,N_48910,N_42802);
and UO_192 (O_192,N_42143,N_43746);
xor UO_193 (O_193,N_48190,N_43189);
xnor UO_194 (O_194,N_43265,N_44997);
and UO_195 (O_195,N_47775,N_47418);
nand UO_196 (O_196,N_43973,N_45447);
and UO_197 (O_197,N_40193,N_49286);
nand UO_198 (O_198,N_45331,N_41549);
xor UO_199 (O_199,N_46486,N_47754);
xnor UO_200 (O_200,N_40862,N_48933);
or UO_201 (O_201,N_44292,N_43797);
xnor UO_202 (O_202,N_40782,N_42276);
xor UO_203 (O_203,N_45263,N_46042);
nand UO_204 (O_204,N_42522,N_46650);
and UO_205 (O_205,N_41567,N_47704);
nor UO_206 (O_206,N_49109,N_49313);
xor UO_207 (O_207,N_44431,N_46155);
and UO_208 (O_208,N_45396,N_46218);
nor UO_209 (O_209,N_45578,N_48107);
or UO_210 (O_210,N_43101,N_47350);
nand UO_211 (O_211,N_49004,N_46327);
or UO_212 (O_212,N_48954,N_49258);
or UO_213 (O_213,N_48283,N_49650);
or UO_214 (O_214,N_45714,N_48523);
nor UO_215 (O_215,N_41868,N_48279);
xnor UO_216 (O_216,N_45341,N_41529);
or UO_217 (O_217,N_42384,N_41960);
or UO_218 (O_218,N_45212,N_45720);
and UO_219 (O_219,N_48212,N_41885);
nand UO_220 (O_220,N_47281,N_44328);
xor UO_221 (O_221,N_48090,N_41550);
and UO_222 (O_222,N_43667,N_42236);
xnor UO_223 (O_223,N_44492,N_41134);
nor UO_224 (O_224,N_47874,N_47312);
and UO_225 (O_225,N_46797,N_43203);
and UO_226 (O_226,N_45328,N_46430);
nand UO_227 (O_227,N_46784,N_48758);
nand UO_228 (O_228,N_43814,N_49469);
xor UO_229 (O_229,N_47957,N_43547);
nor UO_230 (O_230,N_41004,N_46636);
nand UO_231 (O_231,N_41257,N_42645);
and UO_232 (O_232,N_41085,N_47958);
or UO_233 (O_233,N_40443,N_44355);
or UO_234 (O_234,N_46468,N_47162);
nand UO_235 (O_235,N_47885,N_45916);
nor UO_236 (O_236,N_40187,N_45449);
xnor UO_237 (O_237,N_47804,N_46248);
nand UO_238 (O_238,N_42714,N_49520);
and UO_239 (O_239,N_43770,N_48095);
nand UO_240 (O_240,N_42960,N_49678);
and UO_241 (O_241,N_49656,N_44051);
xnor UO_242 (O_242,N_43977,N_41614);
and UO_243 (O_243,N_43267,N_41063);
nor UO_244 (O_244,N_48578,N_48747);
and UO_245 (O_245,N_40472,N_43723);
and UO_246 (O_246,N_48701,N_41656);
nor UO_247 (O_247,N_49060,N_42534);
and UO_248 (O_248,N_46591,N_44953);
or UO_249 (O_249,N_44856,N_47005);
xnor UO_250 (O_250,N_41315,N_40754);
or UO_251 (O_251,N_45611,N_44373);
nor UO_252 (O_252,N_44418,N_47520);
nand UO_253 (O_253,N_45721,N_47811);
and UO_254 (O_254,N_40277,N_49025);
xnor UO_255 (O_255,N_40138,N_40584);
or UO_256 (O_256,N_48440,N_48318);
xor UO_257 (O_257,N_42371,N_40381);
nor UO_258 (O_258,N_44612,N_45818);
nor UO_259 (O_259,N_40331,N_40447);
or UO_260 (O_260,N_48443,N_46871);
xor UO_261 (O_261,N_40001,N_44660);
xnor UO_262 (O_262,N_47228,N_49375);
nand UO_263 (O_263,N_42025,N_47169);
and UO_264 (O_264,N_46388,N_45209);
nor UO_265 (O_265,N_49621,N_45379);
or UO_266 (O_266,N_40194,N_41491);
xor UO_267 (O_267,N_40148,N_49525);
or UO_268 (O_268,N_46292,N_41001);
nor UO_269 (O_269,N_45013,N_43134);
nor UO_270 (O_270,N_45995,N_41443);
and UO_271 (O_271,N_44214,N_43035);
and UO_272 (O_272,N_43671,N_48262);
nor UO_273 (O_273,N_44009,N_48493);
or UO_274 (O_274,N_45560,N_40871);
and UO_275 (O_275,N_43032,N_43222);
xor UO_276 (O_276,N_44310,N_42962);
nor UO_277 (O_277,N_47265,N_43106);
nand UO_278 (O_278,N_43155,N_48425);
and UO_279 (O_279,N_45004,N_48201);
and UO_280 (O_280,N_49024,N_47688);
nor UO_281 (O_281,N_49627,N_41230);
xnor UO_282 (O_282,N_40677,N_49865);
and UO_283 (O_283,N_44060,N_41934);
nand UO_284 (O_284,N_47530,N_49563);
nand UO_285 (O_285,N_41019,N_40823);
xnor UO_286 (O_286,N_48785,N_41292);
or UO_287 (O_287,N_40913,N_49264);
or UO_288 (O_288,N_47611,N_42126);
nand UO_289 (O_289,N_45032,N_41634);
or UO_290 (O_290,N_41974,N_43630);
nor UO_291 (O_291,N_49455,N_41523);
nor UO_292 (O_292,N_42485,N_44504);
and UO_293 (O_293,N_49453,N_46014);
or UO_294 (O_294,N_49078,N_43372);
and UO_295 (O_295,N_41947,N_45896);
xnor UO_296 (O_296,N_41588,N_48191);
and UO_297 (O_297,N_45087,N_42178);
nor UO_298 (O_298,N_49252,N_47593);
nand UO_299 (O_299,N_43309,N_47566);
or UO_300 (O_300,N_42658,N_40481);
and UO_301 (O_301,N_47037,N_49763);
xnor UO_302 (O_302,N_49899,N_41029);
nand UO_303 (O_303,N_46368,N_41185);
or UO_304 (O_304,N_40619,N_49099);
nor UO_305 (O_305,N_40021,N_41912);
or UO_306 (O_306,N_46384,N_44717);
nand UO_307 (O_307,N_40803,N_47780);
nand UO_308 (O_308,N_47339,N_46572);
and UO_309 (O_309,N_45411,N_40589);
xnor UO_310 (O_310,N_49401,N_41080);
nand UO_311 (O_311,N_46848,N_42282);
or UO_312 (O_312,N_43461,N_46027);
nor UO_313 (O_313,N_46204,N_46258);
nor UO_314 (O_314,N_43363,N_42396);
nand UO_315 (O_315,N_44366,N_44582);
or UO_316 (O_316,N_42394,N_41414);
nand UO_317 (O_317,N_49516,N_42297);
nor UO_318 (O_318,N_49501,N_44026);
or UO_319 (O_319,N_43589,N_41510);
nor UO_320 (O_320,N_45353,N_46493);
xor UO_321 (O_321,N_43042,N_43256);
and UO_322 (O_322,N_46390,N_47123);
xnor UO_323 (O_323,N_43756,N_45419);
and UO_324 (O_324,N_49858,N_43390);
or UO_325 (O_325,N_42843,N_47539);
or UO_326 (O_326,N_43443,N_48557);
xor UO_327 (O_327,N_45475,N_44547);
nor UO_328 (O_328,N_41232,N_43343);
nand UO_329 (O_329,N_41632,N_48087);
nor UO_330 (O_330,N_47822,N_49597);
nand UO_331 (O_331,N_41195,N_44970);
nand UO_332 (O_332,N_42160,N_48903);
and UO_333 (O_333,N_48587,N_43629);
nand UO_334 (O_334,N_44180,N_43113);
nor UO_335 (O_335,N_47546,N_48188);
nor UO_336 (O_336,N_47873,N_42981);
xor UO_337 (O_337,N_40538,N_40821);
and UO_338 (O_338,N_47806,N_44798);
nand UO_339 (O_339,N_42120,N_45051);
xnor UO_340 (O_340,N_43074,N_47717);
and UO_341 (O_341,N_46723,N_44627);
and UO_342 (O_342,N_49296,N_40454);
nor UO_343 (O_343,N_40135,N_49105);
and UO_344 (O_344,N_46828,N_49731);
xor UO_345 (O_345,N_44573,N_42706);
nor UO_346 (O_346,N_49617,N_48516);
xnor UO_347 (O_347,N_42613,N_45636);
and UO_348 (O_348,N_46551,N_42604);
nor UO_349 (O_349,N_48732,N_47442);
and UO_350 (O_350,N_42964,N_45042);
xnor UO_351 (O_351,N_46479,N_42991);
nand UO_352 (O_352,N_42430,N_40249);
nor UO_353 (O_353,N_41889,N_46525);
xor UO_354 (O_354,N_49672,N_40387);
xor UO_355 (O_355,N_49795,N_41058);
xor UO_356 (O_356,N_49572,N_43011);
or UO_357 (O_357,N_41824,N_44134);
or UO_358 (O_358,N_40920,N_46660);
nor UO_359 (O_359,N_47685,N_47572);
xor UO_360 (O_360,N_45950,N_43484);
and UO_361 (O_361,N_47670,N_41162);
nand UO_362 (O_362,N_44118,N_46785);
or UO_363 (O_363,N_46209,N_49693);
or UO_364 (O_364,N_40571,N_48865);
nand UO_365 (O_365,N_46347,N_42204);
xnor UO_366 (O_366,N_40012,N_47104);
and UO_367 (O_367,N_44098,N_43118);
xnor UO_368 (O_368,N_40494,N_40445);
nor UO_369 (O_369,N_49341,N_44412);
nor UO_370 (O_370,N_46605,N_48829);
xor UO_371 (O_371,N_47642,N_47789);
or UO_372 (O_372,N_43294,N_43862);
or UO_373 (O_373,N_47388,N_44457);
nor UO_374 (O_374,N_44042,N_40961);
xnor UO_375 (O_375,N_45409,N_42555);
xor UO_376 (O_376,N_49480,N_42248);
nand UO_377 (O_377,N_44630,N_44124);
nand UO_378 (O_378,N_40670,N_43806);
and UO_379 (O_379,N_45697,N_40614);
nand UO_380 (O_380,N_45878,N_40036);
xor UO_381 (O_381,N_46549,N_48471);
xor UO_382 (O_382,N_40367,N_47727);
xor UO_383 (O_383,N_48967,N_41283);
nor UO_384 (O_384,N_49796,N_41675);
xor UO_385 (O_385,N_49981,N_42245);
or UO_386 (O_386,N_48803,N_48399);
or UO_387 (O_387,N_47560,N_44023);
or UO_388 (O_388,N_44713,N_48024);
xnor UO_389 (O_389,N_40546,N_47769);
and UO_390 (O_390,N_44003,N_45694);
xnor UO_391 (O_391,N_42121,N_46245);
nand UO_392 (O_392,N_48871,N_41853);
nand UO_393 (O_393,N_41397,N_44653);
and UO_394 (O_394,N_47614,N_43292);
nand UO_395 (O_395,N_44057,N_48569);
xor UO_396 (O_396,N_43608,N_42351);
nand UO_397 (O_397,N_40426,N_43865);
nor UO_398 (O_398,N_47462,N_42521);
xnor UO_399 (O_399,N_45690,N_40767);
nor UO_400 (O_400,N_47185,N_41289);
and UO_401 (O_401,N_48476,N_48548);
nor UO_402 (O_402,N_42319,N_49732);
and UO_403 (O_403,N_48220,N_41383);
nand UO_404 (O_404,N_46070,N_48077);
or UO_405 (O_405,N_42516,N_49822);
nor UO_406 (O_406,N_44610,N_40428);
nand UO_407 (O_407,N_47965,N_40174);
nor UO_408 (O_408,N_49785,N_43836);
nor UO_409 (O_409,N_45431,N_45503);
nor UO_410 (O_410,N_42308,N_47129);
xnor UO_411 (O_411,N_40763,N_43592);
xnor UO_412 (O_412,N_40764,N_44411);
xor UO_413 (O_413,N_47047,N_47276);
nor UO_414 (O_414,N_44986,N_44583);
or UO_415 (O_415,N_43700,N_43638);
and UO_416 (O_416,N_40113,N_46869);
and UO_417 (O_417,N_43344,N_45446);
or UO_418 (O_418,N_40753,N_42786);
nand UO_419 (O_419,N_45577,N_49519);
nand UO_420 (O_420,N_45441,N_40977);
or UO_421 (O_421,N_48091,N_40240);
nor UO_422 (O_422,N_45622,N_47338);
nand UO_423 (O_423,N_42884,N_43049);
or UO_424 (O_424,N_49014,N_46598);
nand UO_425 (O_425,N_48519,N_45607);
nor UO_426 (O_426,N_44629,N_41784);
nor UO_427 (O_427,N_46104,N_44803);
xor UO_428 (O_428,N_45305,N_48136);
xnor UO_429 (O_429,N_43214,N_48850);
nor UO_430 (O_430,N_48505,N_48184);
nand UO_431 (O_431,N_46967,N_44452);
nor UO_432 (O_432,N_44807,N_43225);
or UO_433 (O_433,N_40988,N_40201);
or UO_434 (O_434,N_43937,N_43644);
and UO_435 (O_435,N_47999,N_40768);
and UO_436 (O_436,N_44503,N_48634);
or UO_437 (O_437,N_43907,N_47213);
or UO_438 (O_438,N_46008,N_43459);
nor UO_439 (O_439,N_41144,N_48526);
xnor UO_440 (O_440,N_49059,N_45080);
and UO_441 (O_441,N_42977,N_43968);
xnor UO_442 (O_442,N_44099,N_45060);
xor UO_443 (O_443,N_45912,N_44251);
and UO_444 (O_444,N_47062,N_41356);
nor UO_445 (O_445,N_49409,N_47337);
nor UO_446 (O_446,N_42355,N_40478);
nand UO_447 (O_447,N_41404,N_40935);
nand UO_448 (O_448,N_47777,N_44561);
nor UO_449 (O_449,N_49165,N_45898);
or UO_450 (O_450,N_41090,N_46073);
nand UO_451 (O_451,N_43181,N_43854);
xor UO_452 (O_452,N_45588,N_42638);
nor UO_453 (O_453,N_42808,N_45370);
xor UO_454 (O_454,N_48754,N_49721);
xor UO_455 (O_455,N_42595,N_40607);
xnor UO_456 (O_456,N_46632,N_43607);
or UO_457 (O_457,N_45239,N_49013);
nor UO_458 (O_458,N_49945,N_41262);
nor UO_459 (O_459,N_42797,N_47122);
and UO_460 (O_460,N_45726,N_42196);
xor UO_461 (O_461,N_40798,N_40479);
nand UO_462 (O_462,N_42184,N_44937);
or UO_463 (O_463,N_47666,N_48366);
nand UO_464 (O_464,N_48432,N_45375);
nand UO_465 (O_465,N_44190,N_44701);
nor UO_466 (O_466,N_44071,N_41537);
nand UO_467 (O_467,N_42885,N_48514);
or UO_468 (O_468,N_48677,N_44740);
and UO_469 (O_469,N_41931,N_49388);
nor UO_470 (O_470,N_41507,N_49613);
xnor UO_471 (O_471,N_47272,N_47888);
nand UO_472 (O_472,N_49768,N_47141);
nand UO_473 (O_473,N_47918,N_47986);
or UO_474 (O_474,N_43172,N_43767);
nor UO_475 (O_475,N_43984,N_40772);
or UO_476 (O_476,N_49927,N_45834);
nor UO_477 (O_477,N_43000,N_43664);
or UO_478 (O_478,N_42290,N_45923);
nand UO_479 (O_479,N_48576,N_45891);
and UO_480 (O_480,N_49799,N_43005);
nand UO_481 (O_481,N_48470,N_47855);
nand UO_482 (O_482,N_44534,N_45556);
nor UO_483 (O_483,N_43533,N_44390);
nand UO_484 (O_484,N_45106,N_48724);
nand UO_485 (O_485,N_45471,N_49770);
nor UO_486 (O_486,N_48828,N_42041);
nor UO_487 (O_487,N_46100,N_45856);
or UO_488 (O_488,N_47271,N_46074);
or UO_489 (O_489,N_49686,N_47112);
nand UO_490 (O_490,N_47961,N_49051);
xnor UO_491 (O_491,N_45805,N_43743);
and UO_492 (O_492,N_42498,N_42924);
nor UO_493 (O_493,N_42736,N_48234);
nor UO_494 (O_494,N_44137,N_46064);
xnor UO_495 (O_495,N_47814,N_47000);
or UO_496 (O_496,N_47783,N_46257);
or UO_497 (O_497,N_46580,N_42566);
or UO_498 (O_498,N_45023,N_46089);
nand UO_499 (O_499,N_49689,N_48592);
nand UO_500 (O_500,N_41705,N_49075);
xnor UO_501 (O_501,N_40225,N_44489);
nor UO_502 (O_502,N_45865,N_47026);
and UO_503 (O_503,N_42983,N_47851);
nor UO_504 (O_504,N_47419,N_45874);
and UO_505 (O_505,N_43478,N_43196);
and UO_506 (O_506,N_42746,N_47189);
and UO_507 (O_507,N_48678,N_47429);
nor UO_508 (O_508,N_46936,N_49733);
and UO_509 (O_509,N_40243,N_48182);
and UO_510 (O_510,N_49394,N_47819);
or UO_511 (O_511,N_40672,N_41269);
nor UO_512 (O_512,N_44260,N_48480);
nand UO_513 (O_513,N_45421,N_45654);
or UO_514 (O_514,N_41112,N_43540);
and UO_515 (O_515,N_48101,N_47768);
and UO_516 (O_516,N_45059,N_40323);
and UO_517 (O_517,N_43497,N_49601);
nor UO_518 (O_518,N_43503,N_47273);
or UO_519 (O_519,N_49211,N_40509);
xor UO_520 (O_520,N_40127,N_48199);
xnor UO_521 (O_521,N_43143,N_44159);
xor UO_522 (O_522,N_46039,N_44224);
nor UO_523 (O_523,N_43481,N_43579);
and UO_524 (O_524,N_47908,N_48294);
xnor UO_525 (O_525,N_41071,N_45068);
xnor UO_526 (O_526,N_44078,N_43549);
nand UO_527 (O_527,N_45663,N_45235);
or UO_528 (O_528,N_49787,N_47734);
nor UO_529 (O_529,N_47807,N_44013);
nor UO_530 (O_530,N_40828,N_40743);
xnor UO_531 (O_531,N_47127,N_44148);
nand UO_532 (O_532,N_40878,N_40911);
nand UO_533 (O_533,N_49047,N_45644);
nand UO_534 (O_534,N_44559,N_41891);
and UO_535 (O_535,N_47175,N_40981);
nand UO_536 (O_536,N_41980,N_41437);
and UO_537 (O_537,N_45222,N_42902);
and UO_538 (O_538,N_49359,N_49132);
and UO_539 (O_539,N_44893,N_44036);
xor UO_540 (O_540,N_43987,N_45460);
nand UO_541 (O_541,N_49747,N_48583);
and UO_542 (O_542,N_41658,N_48662);
xor UO_543 (O_543,N_41374,N_42507);
and UO_544 (O_544,N_44465,N_41505);
and UO_545 (O_545,N_44061,N_44285);
or UO_546 (O_546,N_48004,N_43788);
and UO_547 (O_547,N_44181,N_40498);
or UO_548 (O_548,N_43744,N_45075);
xnor UO_549 (O_549,N_46831,N_42989);
nand UO_550 (O_550,N_43212,N_44246);
or UO_551 (O_551,N_42570,N_42525);
nor UO_552 (O_552,N_47637,N_40662);
nand UO_553 (O_553,N_48621,N_47868);
xnor UO_554 (O_554,N_48506,N_43486);
or UO_555 (O_555,N_46030,N_40110);
nand UO_556 (O_556,N_43908,N_41707);
nand UO_557 (O_557,N_45488,N_47416);
and UO_558 (O_558,N_44389,N_41714);
and UO_559 (O_559,N_42215,N_46050);
and UO_560 (O_560,N_48687,N_47905);
nor UO_561 (O_561,N_41669,N_41766);
nand UO_562 (O_562,N_42207,N_44363);
xor UO_563 (O_563,N_44991,N_46850);
nand UO_564 (O_564,N_42776,N_40344);
or UO_565 (O_565,N_48033,N_42186);
nor UO_566 (O_566,N_41944,N_41351);
nand UO_567 (O_567,N_44096,N_49538);
nand UO_568 (O_568,N_44510,N_49467);
or UO_569 (O_569,N_49262,N_45094);
xor UO_570 (O_570,N_48670,N_44001);
nor UO_571 (O_571,N_44847,N_42634);
or UO_572 (O_572,N_47238,N_44948);
or UO_573 (O_573,N_49941,N_49527);
nor UO_574 (O_574,N_42491,N_47673);
nand UO_575 (O_575,N_49160,N_48068);
nor UO_576 (O_576,N_45746,N_40802);
or UO_577 (O_577,N_40731,N_46952);
or UO_578 (O_578,N_43253,N_43537);
and UO_579 (O_579,N_45147,N_41738);
xnor UO_580 (O_580,N_45555,N_46326);
nor UO_581 (O_581,N_48765,N_45067);
nand UO_582 (O_582,N_41748,N_46617);
or UO_583 (O_583,N_41698,N_49544);
xnor UO_584 (O_584,N_49378,N_47060);
nand UO_585 (O_585,N_44782,N_40835);
nor UO_586 (O_586,N_49489,N_46835);
or UO_587 (O_587,N_44325,N_47266);
or UO_588 (O_588,N_49873,N_47901);
nor UO_589 (O_589,N_44779,N_44074);
nor UO_590 (O_590,N_48860,N_45113);
nand UO_591 (O_591,N_45747,N_46191);
and UO_592 (O_592,N_42422,N_44183);
xnor UO_593 (O_593,N_40991,N_49696);
nand UO_594 (O_594,N_40293,N_44065);
and UO_595 (O_595,N_46031,N_43954);
and UO_596 (O_596,N_48949,N_43230);
xor UO_597 (O_597,N_48028,N_46681);
nor UO_598 (O_598,N_42179,N_41079);
or UO_599 (O_599,N_48588,N_49340);
or UO_600 (O_600,N_42974,N_43135);
nand UO_601 (O_601,N_47882,N_44037);
or UO_602 (O_602,N_49052,N_42244);
xor UO_603 (O_603,N_42790,N_44537);
nor UO_604 (O_604,N_45364,N_43213);
nor UO_605 (O_605,N_44608,N_42527);
nand UO_606 (O_606,N_43401,N_40796);
nand UO_607 (O_607,N_48051,N_46233);
and UO_608 (O_608,N_47723,N_47974);
or UO_609 (O_609,N_46538,N_48742);
nor UO_610 (O_610,N_42803,N_40000);
nand UO_611 (O_611,N_49404,N_42747);
nand UO_612 (O_612,N_49989,N_40947);
xor UO_613 (O_613,N_43102,N_40003);
nand UO_614 (O_614,N_41164,N_49800);
and UO_615 (O_615,N_44535,N_46372);
and UO_616 (O_616,N_46547,N_49251);
xnor UO_617 (O_617,N_45425,N_45942);
xnor UO_618 (O_618,N_46288,N_42858);
nand UO_619 (O_619,N_49122,N_49061);
and UO_620 (O_620,N_42304,N_49310);
or UO_621 (O_621,N_40505,N_44505);
or UO_622 (O_622,N_41102,N_46765);
nor UO_623 (O_623,N_43015,N_40616);
and UO_624 (O_624,N_47833,N_45443);
xnor UO_625 (O_625,N_49463,N_45978);
and UO_626 (O_626,N_43368,N_44817);
and UO_627 (O_627,N_41915,N_42617);
and UO_628 (O_628,N_47394,N_46392);
nor UO_629 (O_629,N_47778,N_45324);
nand UO_630 (O_630,N_42163,N_44705);
nand UO_631 (O_631,N_49630,N_44988);
and UO_632 (O_632,N_44901,N_40719);
xor UO_633 (O_633,N_44106,N_48920);
and UO_634 (O_634,N_46808,N_43921);
nand UO_635 (O_635,N_44513,N_49529);
and UO_636 (O_636,N_47166,N_42105);
nand UO_637 (O_637,N_46365,N_49478);
xnor UO_638 (O_638,N_40918,N_42113);
nor UO_639 (O_639,N_41908,N_44879);
and UO_640 (O_640,N_41533,N_42413);
nand UO_641 (O_641,N_40362,N_43588);
nor UO_642 (O_642,N_47398,N_43594);
xnor UO_643 (O_643,N_41093,N_47533);
nand UO_644 (O_644,N_41739,N_45241);
xor UO_645 (O_645,N_41155,N_41992);
nor UO_646 (O_646,N_42511,N_40533);
nor UO_647 (O_647,N_45592,N_41068);
or UO_648 (O_648,N_45030,N_47006);
or UO_649 (O_649,N_48722,N_44243);
or UO_650 (O_650,N_48749,N_43398);
xnor UO_651 (O_651,N_45486,N_40691);
xor UO_652 (O_652,N_46361,N_48276);
and UO_653 (O_653,N_40171,N_41602);
or UO_654 (O_654,N_47096,N_48338);
xor UO_655 (O_655,N_42098,N_47658);
or UO_656 (O_656,N_48671,N_44708);
xor UO_657 (O_657,N_42280,N_43215);
nand UO_658 (O_658,N_48833,N_46349);
or UO_659 (O_659,N_41109,N_49921);
and UO_660 (O_660,N_44356,N_47118);
nand UO_661 (O_661,N_42920,N_41305);
xnor UO_662 (O_662,N_40655,N_47070);
xor UO_663 (O_663,N_40537,N_41812);
and UO_664 (O_664,N_49345,N_48789);
nor UO_665 (O_665,N_44750,N_43017);
xnor UO_666 (O_666,N_44462,N_42123);
nand UO_667 (O_667,N_49035,N_45128);
nor UO_668 (O_668,N_48235,N_40256);
nor UO_669 (O_669,N_49610,N_45778);
or UO_670 (O_670,N_47969,N_44838);
xnor UO_671 (O_671,N_48948,N_41847);
and UO_672 (O_672,N_43124,N_47784);
or UO_673 (O_673,N_48236,N_46775);
nor UO_674 (O_674,N_43380,N_41204);
xnor UO_675 (O_675,N_45399,N_48979);
xnor UO_676 (O_676,N_47978,N_44121);
and UO_677 (O_677,N_43006,N_46766);
nand UO_678 (O_678,N_42644,N_40015);
or UO_679 (O_679,N_40483,N_47601);
and UO_680 (O_680,N_47165,N_42615);
and UO_681 (O_681,N_47226,N_45798);
nor UO_682 (O_682,N_47087,N_48770);
nor UO_683 (O_683,N_49552,N_43824);
xnor UO_684 (O_684,N_45155,N_48931);
nor UO_685 (O_685,N_40879,N_42859);
xor UO_686 (O_686,N_40969,N_45736);
nand UO_687 (O_687,N_46726,N_43902);
nand UO_688 (O_688,N_43885,N_45759);
and UO_689 (O_689,N_47328,N_47995);
nand UO_690 (O_690,N_40970,N_43621);
nor UO_691 (O_691,N_43084,N_49471);
nor UO_692 (O_692,N_40915,N_40311);
nand UO_693 (O_693,N_47206,N_45922);
nor UO_694 (O_694,N_44619,N_48094);
and UO_695 (O_695,N_47680,N_49654);
nand UO_696 (O_696,N_47613,N_46892);
xor UO_697 (O_697,N_46157,N_44357);
nand UO_698 (O_698,N_41603,N_49201);
or UO_699 (O_699,N_44327,N_46773);
nor UO_700 (O_700,N_46870,N_41095);
xor UO_701 (O_701,N_41619,N_49369);
or UO_702 (O_702,N_47242,N_45945);
nand UO_703 (O_703,N_42605,N_42806);
nor UO_704 (O_704,N_47080,N_40396);
nor UO_705 (O_705,N_44162,N_49748);
and UO_706 (O_706,N_49297,N_40203);
nor UO_707 (O_707,N_43957,N_49674);
xor UO_708 (O_708,N_43764,N_47200);
nor UO_709 (O_709,N_42827,N_42557);
nand UO_710 (O_710,N_43433,N_47157);
or UO_711 (O_711,N_42811,N_44200);
or UO_712 (O_712,N_48762,N_42165);
and UO_713 (O_713,N_41294,N_49062);
xor UO_714 (O_714,N_48215,N_41554);
or UO_715 (O_715,N_42543,N_43873);
or UO_716 (O_716,N_48802,N_43293);
nand UO_717 (O_717,N_49232,N_43631);
and UO_718 (O_718,N_49974,N_49923);
and UO_719 (O_719,N_48719,N_42151);
xnor UO_720 (O_720,N_44132,N_47632);
nand UO_721 (O_721,N_42440,N_46237);
nand UO_722 (O_722,N_41830,N_49964);
nand UO_723 (O_723,N_43705,N_44053);
or UO_724 (O_724,N_48543,N_49911);
nand UO_725 (O_725,N_44604,N_46370);
nor UO_726 (O_726,N_49615,N_43725);
nand UO_727 (O_727,N_48030,N_40668);
nor UO_728 (O_728,N_44641,N_44785);
or UO_729 (O_729,N_41898,N_49975);
nor UO_730 (O_730,N_48650,N_42340);
and UO_731 (O_731,N_42370,N_43479);
xnor UO_732 (O_732,N_49938,N_42967);
xor UO_733 (O_733,N_42946,N_49798);
nor UO_734 (O_734,N_41241,N_42824);
nor UO_735 (O_735,N_49386,N_42086);
nand UO_736 (O_736,N_43317,N_47446);
and UO_737 (O_737,N_41598,N_44038);
nor UO_738 (O_738,N_40156,N_41746);
and UO_739 (O_739,N_44256,N_44211);
and UO_740 (O_740,N_47221,N_46893);
nand UO_741 (O_741,N_41928,N_44015);
xor UO_742 (O_742,N_49603,N_47795);
and UO_743 (O_743,N_45596,N_40017);
nand UO_744 (O_744,N_47176,N_46400);
or UO_745 (O_745,N_48128,N_41636);
xnor UO_746 (O_746,N_46407,N_42229);
and UO_747 (O_747,N_42684,N_43051);
or UO_748 (O_748,N_41893,N_46552);
nor UO_749 (O_749,N_49427,N_49971);
nand UO_750 (O_750,N_49389,N_40793);
and UO_751 (O_751,N_45050,N_41778);
xor UO_752 (O_752,N_42449,N_48601);
and UO_753 (O_753,N_41111,N_45107);
or UO_754 (O_754,N_49930,N_46354);
and UO_755 (O_755,N_48488,N_41176);
or UO_756 (O_756,N_48607,N_49728);
nor UO_757 (O_757,N_45552,N_45053);
and UO_758 (O_758,N_46858,N_47973);
nand UO_759 (O_759,N_41797,N_41271);
xnor UO_760 (O_760,N_46606,N_46029);
nor UO_761 (O_761,N_45689,N_45434);
nor UO_762 (O_762,N_45788,N_46461);
or UO_763 (O_763,N_46956,N_44792);
nor UO_764 (O_764,N_43090,N_46105);
or UO_765 (O_765,N_44564,N_44525);
xor UO_766 (O_766,N_46807,N_48016);
or UO_767 (O_767,N_46962,N_44767);
xnor UO_768 (O_768,N_49707,N_40583);
nand UO_769 (O_769,N_41640,N_46634);
nand UO_770 (O_770,N_44206,N_42984);
xnor UO_771 (O_771,N_46474,N_45879);
and UO_772 (O_772,N_44637,N_45943);
and UO_773 (O_773,N_46478,N_48771);
nor UO_774 (O_774,N_41829,N_49237);
and UO_775 (O_775,N_49571,N_45581);
xnor UO_776 (O_776,N_43438,N_45024);
xnor UO_777 (O_777,N_45568,N_48729);
nor UO_778 (O_778,N_44031,N_43755);
xnor UO_779 (O_779,N_43254,N_45323);
nor UO_780 (O_780,N_46825,N_47990);
or UO_781 (O_781,N_43397,N_47191);
or UO_782 (O_782,N_41583,N_41955);
nor UO_783 (O_783,N_45415,N_46426);
and UO_784 (O_784,N_43748,N_48363);
nand UO_785 (O_785,N_42375,N_42054);
nand UO_786 (O_786,N_41643,N_48078);
nand UO_787 (O_787,N_45076,N_46860);
xor UO_788 (O_788,N_40899,N_42274);
or UO_789 (O_789,N_47282,N_46371);
or UO_790 (O_790,N_46036,N_42836);
nand UO_791 (O_791,N_47967,N_42758);
and UO_792 (O_792,N_47787,N_47919);
nand UO_793 (O_793,N_49637,N_45658);
nand UO_794 (O_794,N_43288,N_42437);
nor UO_795 (O_795,N_41886,N_44027);
nor UO_796 (O_796,N_46926,N_46463);
xnor UO_797 (O_797,N_46561,N_43442);
nor UO_798 (O_798,N_42825,N_49253);
nand UO_799 (O_799,N_48285,N_46193);
and UO_800 (O_800,N_48520,N_40199);
nand UO_801 (O_801,N_46098,N_46047);
nand UO_802 (O_802,N_44780,N_45044);
nand UO_803 (O_803,N_49924,N_44110);
xor UO_804 (O_804,N_47945,N_41737);
xor UO_805 (O_805,N_46635,N_47864);
and UO_806 (O_806,N_49708,N_40490);
nor UO_807 (O_807,N_43096,N_49022);
or UO_808 (O_808,N_41415,N_41022);
nand UO_809 (O_809,N_48241,N_47816);
or UO_810 (O_810,N_48980,N_43969);
xnor UO_811 (O_811,N_46758,N_46091);
and UO_812 (O_812,N_43546,N_41736);
or UO_813 (O_813,N_42921,N_45453);
and UO_814 (O_814,N_44403,N_43218);
nand UO_815 (O_815,N_49639,N_40224);
and UO_816 (O_816,N_44869,N_46285);
nand UO_817 (O_817,N_45927,N_40843);
and UO_818 (O_818,N_48222,N_49354);
xnor UO_819 (O_819,N_45570,N_48123);
nor UO_820 (O_820,N_40335,N_49541);
nand UO_821 (O_821,N_43881,N_41148);
or UO_822 (O_822,N_47131,N_44595);
nor UO_823 (O_823,N_42980,N_42494);
or UO_824 (O_824,N_43958,N_48535);
xor UO_825 (O_825,N_47009,N_43494);
xor UO_826 (O_826,N_48079,N_48159);
nand UO_827 (O_827,N_47217,N_49756);
xor UO_828 (O_828,N_49936,N_48898);
and UO_829 (O_829,N_44726,N_49900);
nand UO_830 (O_830,N_47627,N_47349);
nand UO_831 (O_831,N_40316,N_45114);
nor UO_832 (O_832,N_42266,N_41413);
xor UO_833 (O_833,N_47378,N_46977);
and UO_834 (O_834,N_49994,N_46906);
nand UO_835 (O_835,N_42970,N_45467);
nor UO_836 (O_836,N_42897,N_41490);
nor UO_837 (O_837,N_49036,N_47375);
nor UO_838 (O_838,N_44092,N_41783);
xor UO_839 (O_839,N_45144,N_47913);
nand UO_840 (O_840,N_40818,N_45974);
nand UO_841 (O_841,N_42944,N_41384);
nand UO_842 (O_842,N_42250,N_41128);
nor UO_843 (O_843,N_48495,N_46750);
nand UO_844 (O_844,N_42360,N_42834);
or UO_845 (O_845,N_46639,N_44695);
and UO_846 (O_846,N_47588,N_49995);
or UO_847 (O_847,N_40044,N_40880);
and UO_848 (O_848,N_44673,N_48180);
nor UO_849 (O_849,N_41431,N_41703);
nand UO_850 (O_850,N_43934,N_41599);
or UO_851 (O_851,N_42329,N_45186);
and UO_852 (O_852,N_49920,N_42976);
nor UO_853 (O_853,N_41156,N_45010);
or UO_854 (O_854,N_47548,N_44337);
or UO_855 (O_855,N_47887,N_42529);
nand UO_856 (O_856,N_40626,N_47099);
xnor UO_857 (O_857,N_43200,N_49304);
and UO_858 (O_858,N_44095,N_48304);
and UO_859 (O_859,N_40732,N_40319);
nand UO_860 (O_860,N_41907,N_40591);
xnor UO_861 (O_861,N_40322,N_43763);
nor UO_862 (O_862,N_44133,N_43765);
nand UO_863 (O_863,N_46777,N_41530);
nand UO_864 (O_864,N_47147,N_40442);
xor UO_865 (O_865,N_44633,N_49102);
and UO_866 (O_866,N_42588,N_44063);
nor UO_867 (O_867,N_41512,N_41903);
nand UO_868 (O_868,N_41037,N_42475);
and UO_869 (O_869,N_42695,N_48748);
or UO_870 (O_870,N_47879,N_40721);
and UO_871 (O_871,N_44725,N_46208);
or UO_872 (O_872,N_49884,N_41759);
or UO_873 (O_873,N_49275,N_47606);
nor UO_874 (O_874,N_43115,N_40776);
or UO_875 (O_875,N_41641,N_49476);
xnor UO_876 (O_876,N_48194,N_41852);
nor UO_877 (O_877,N_49569,N_43999);
nand UO_878 (O_878,N_42337,N_44279);
and UO_879 (O_879,N_48885,N_47972);
nor UO_880 (O_880,N_45890,N_42556);
nand UO_881 (O_881,N_40294,N_41187);
and UO_882 (O_882,N_47834,N_46410);
or UO_883 (O_883,N_40658,N_47153);
nor UO_884 (O_884,N_48836,N_42314);
or UO_885 (O_885,N_42101,N_47396);
xnor UO_886 (O_886,N_40501,N_41485);
nand UO_887 (O_887,N_40833,N_44188);
nand UO_888 (O_888,N_48278,N_42757);
nor UO_889 (O_889,N_40022,N_47599);
nor UO_890 (O_890,N_42155,N_42295);
xnor UO_891 (O_891,N_40402,N_42012);
nand UO_892 (O_892,N_47925,N_49918);
xnor UO_893 (O_893,N_49254,N_48189);
nor UO_894 (O_894,N_49724,N_48987);
or UO_895 (O_895,N_47170,N_47316);
or UO_896 (O_896,N_42444,N_45162);
nand UO_897 (O_897,N_44108,N_41196);
or UO_898 (O_898,N_44622,N_49191);
nor UO_899 (O_899,N_43364,N_46826);
xnor UO_900 (O_900,N_44994,N_43847);
xnor UO_901 (O_901,N_44613,N_49346);
or UO_902 (O_902,N_44002,N_47705);
nor UO_903 (O_903,N_48779,N_48579);
or UO_904 (O_904,N_45764,N_49937);
and UO_905 (O_905,N_41972,N_45532);
xnor UO_906 (O_906,N_48108,N_47730);
xor UO_907 (O_907,N_42793,N_40482);
or UO_908 (O_908,N_49765,N_45905);
nor UO_909 (O_909,N_46658,N_41831);
xor UO_910 (O_910,N_46102,N_46992);
nor UO_911 (O_911,N_42569,N_45546);
xor UO_912 (O_912,N_40650,N_44599);
nand UO_913 (O_913,N_48081,N_48302);
xor UO_914 (O_914,N_45633,N_40324);
nand UO_915 (O_915,N_44544,N_44895);
or UO_916 (O_916,N_46712,N_41061);
nor UO_917 (O_917,N_41246,N_44094);
or UO_918 (O_918,N_48127,N_44498);
nor UO_919 (O_919,N_47928,N_43674);
and UO_920 (O_920,N_48089,N_46999);
nor UO_921 (O_921,N_47551,N_44548);
nand UO_922 (O_922,N_43614,N_43568);
xnor UO_923 (O_923,N_41387,N_43314);
or UO_924 (O_924,N_47915,N_48173);
and UO_925 (O_925,N_40649,N_48259);
nand UO_926 (O_926,N_49806,N_44899);
or UO_927 (O_927,N_40265,N_43030);
and UO_928 (O_928,N_49499,N_45261);
and UO_929 (O_929,N_47317,N_48309);
xor UO_930 (O_930,N_45174,N_45360);
xor UO_931 (O_931,N_40245,N_49145);
xnor UO_932 (O_932,N_41611,N_44039);
and UO_933 (O_933,N_47645,N_40453);
nor UO_934 (O_934,N_44295,N_43679);
nor UO_935 (O_935,N_43582,N_42766);
nand UO_936 (O_936,N_44668,N_44707);
xnor UO_937 (O_937,N_44174,N_43800);
xnor UO_938 (O_938,N_42545,N_44929);
xnor UO_939 (O_939,N_43327,N_44274);
xnor UO_940 (O_940,N_44577,N_49352);
xor UO_941 (O_941,N_43161,N_40185);
xnor UO_942 (O_942,N_41925,N_49046);
xor UO_943 (O_943,N_42701,N_49164);
nor UO_944 (O_944,N_44400,N_48787);
or UO_945 (O_945,N_49575,N_42336);
nand UO_946 (O_946,N_45093,N_43597);
nor UO_947 (O_947,N_45232,N_40728);
nor UO_948 (O_948,N_46845,N_44888);
nand UO_949 (O_949,N_41701,N_45823);
or UO_950 (O_950,N_40104,N_41321);
xor UO_951 (O_951,N_44563,N_44958);
and UO_952 (O_952,N_41369,N_45124);
xor UO_953 (O_953,N_47146,N_46579);
nand UO_954 (O_954,N_47285,N_42089);
xnor UO_955 (O_955,N_48031,N_43081);
xor UO_956 (O_956,N_41017,N_44232);
xnor UO_957 (O_957,N_42531,N_45687);
xnor UO_958 (O_958,N_49385,N_43429);
xnor UO_959 (O_959,N_40757,N_44305);
nor UO_960 (O_960,N_45594,N_49907);
nor UO_961 (O_961,N_49488,N_40418);
nor UO_962 (O_962,N_42095,N_49856);
nor UO_963 (O_963,N_46129,N_47110);
nor UO_964 (O_964,N_41067,N_48469);
xnor UO_965 (O_965,N_47840,N_43146);
and UO_966 (O_966,N_43116,N_42415);
and UO_967 (O_967,N_44655,N_45296);
and UO_968 (O_968,N_49712,N_45490);
xor UO_969 (O_969,N_49616,N_49871);
xor UO_970 (O_970,N_41201,N_45386);
xnor UO_971 (O_971,N_48835,N_42958);
nand UO_972 (O_972,N_41419,N_43832);
or UO_973 (O_973,N_42048,N_47149);
and UO_974 (O_974,N_46380,N_45031);
or UO_975 (O_975,N_44866,N_49431);
xnor UO_976 (O_976,N_44771,N_41425);
nor UO_977 (O_977,N_40500,N_47371);
or UO_978 (O_978,N_45779,N_47979);
nor UO_979 (O_979,N_45566,N_47148);
nand UO_980 (O_980,N_42436,N_49851);
or UO_981 (O_981,N_43297,N_40994);
nor UO_982 (O_982,N_48367,N_43575);
nand UO_983 (O_983,N_45722,N_41666);
xnor UO_984 (O_984,N_42683,N_44916);
nor UO_985 (O_985,N_44444,N_42167);
nor UO_986 (O_986,N_45478,N_44995);
or UO_987 (O_987,N_47628,N_47066);
nor UO_988 (O_988,N_48692,N_45363);
or UO_989 (O_989,N_48697,N_47320);
or UO_990 (O_990,N_43149,N_41732);
xnor UO_991 (O_991,N_41920,N_46680);
nor UO_992 (O_992,N_47397,N_46702);
nor UO_993 (O_993,N_43132,N_48393);
xor UO_994 (O_994,N_47983,N_46200);
xor UO_995 (O_995,N_42131,N_42462);
or UO_996 (O_996,N_45371,N_41850);
nand UO_997 (O_997,N_49828,N_49245);
nand UO_998 (O_998,N_42685,N_45755);
nor UO_999 (O_999,N_46083,N_42672);
nor UO_1000 (O_1000,N_49284,N_44123);
nor UO_1001 (O_1001,N_49133,N_45868);
or UO_1002 (O_1002,N_43287,N_41213);
or UO_1003 (O_1003,N_44385,N_43538);
nor UO_1004 (O_1004,N_45610,N_49468);
nor UO_1005 (O_1005,N_47381,N_41874);
nand UO_1006 (O_1006,N_42930,N_42717);
and UO_1007 (O_1007,N_48282,N_49096);
nand UO_1008 (O_1008,N_40115,N_44430);
nor UO_1009 (O_1009,N_41526,N_45660);
and UO_1010 (O_1010,N_48329,N_44998);
nand UO_1011 (O_1011,N_49985,N_40413);
xor UO_1012 (O_1012,N_42134,N_48401);
and UO_1013 (O_1013,N_45815,N_40712);
nand UO_1014 (O_1014,N_47633,N_48437);
xor UO_1015 (O_1015,N_46743,N_49864);
nand UO_1016 (O_1016,N_40725,N_42421);
and UO_1017 (O_1017,N_48217,N_43353);
or UO_1018 (O_1018,N_45104,N_46494);
nor UO_1019 (O_1019,N_47030,N_49559);
nand UO_1020 (O_1020,N_41851,N_43321);
nor UO_1021 (O_1021,N_42996,N_42000);
nand UO_1022 (O_1022,N_45192,N_46043);
nand UO_1023 (O_1023,N_45484,N_42928);
nand UO_1024 (O_1024,N_44718,N_46131);
nand UO_1025 (O_1025,N_40780,N_40643);
and UO_1026 (O_1026,N_48169,N_47653);
and UO_1027 (O_1027,N_49523,N_42799);
xnor UO_1028 (O_1028,N_40320,N_47498);
or UO_1029 (O_1029,N_40378,N_40938);
xnor UO_1030 (O_1030,N_42823,N_40457);
xor UO_1031 (O_1031,N_43757,N_40376);
or UO_1032 (O_1032,N_49342,N_47687);
xnor UO_1033 (O_1033,N_47697,N_47032);
nor UO_1034 (O_1034,N_42538,N_49919);
and UO_1035 (O_1035,N_42221,N_42666);
and UO_1036 (O_1036,N_45649,N_44101);
and UO_1037 (O_1037,N_49371,N_43485);
nor UO_1038 (O_1038,N_49085,N_45752);
nand UO_1039 (O_1039,N_47359,N_40685);
xor UO_1040 (O_1040,N_44161,N_40283);
and UO_1041 (O_1041,N_44196,N_46298);
or UO_1042 (O_1042,N_49599,N_47250);
nand UO_1043 (O_1043,N_44519,N_41065);
and UO_1044 (O_1044,N_49655,N_44990);
nand UO_1045 (O_1045,N_48817,N_43861);
and UO_1046 (O_1046,N_44379,N_45071);
xnor UO_1047 (O_1047,N_45440,N_46754);
or UO_1048 (O_1048,N_48156,N_41538);
xor UO_1049 (O_1049,N_49521,N_41873);
nor UO_1050 (O_1050,N_41242,N_47883);
nand UO_1051 (O_1051,N_45420,N_46088);
or UO_1052 (O_1052,N_48550,N_44789);
nand UO_1053 (O_1053,N_45913,N_45065);
nor UO_1054 (O_1054,N_42963,N_48921);
or UO_1055 (O_1055,N_40218,N_46160);
nand UO_1056 (O_1056,N_48970,N_40748);
nor UO_1057 (O_1057,N_43620,N_40909);
xor UO_1058 (O_1058,N_46925,N_47582);
nand UO_1059 (O_1059,N_43117,N_43918);
or UO_1060 (O_1060,N_49593,N_43385);
and UO_1061 (O_1061,N_48296,N_43733);
or UO_1062 (O_1062,N_49680,N_49764);
nand UO_1063 (O_1063,N_44146,N_46798);
and UO_1064 (O_1064,N_40209,N_40422);
and UO_1065 (O_1065,N_46603,N_45435);
nand UO_1066 (O_1066,N_48672,N_42641);
nor UO_1067 (O_1067,N_46108,N_49175);
nand UO_1068 (O_1068,N_48472,N_46133);
xnor UO_1069 (O_1069,N_47045,N_42457);
and UO_1070 (O_1070,N_46462,N_46881);
nand UO_1071 (O_1071,N_46955,N_45320);
nand UO_1072 (O_1072,N_45016,N_40380);
or UO_1073 (O_1073,N_44521,N_40134);
nor UO_1074 (O_1074,N_45536,N_49514);
xnor UO_1075 (O_1075,N_44788,N_40296);
xnor UO_1076 (O_1076,N_45811,N_42321);
nor UO_1077 (O_1077,N_40715,N_49753);
and UO_1078 (O_1078,N_45944,N_48006);
nand UO_1079 (O_1079,N_41994,N_41051);
xor UO_1080 (O_1080,N_42466,N_40239);
or UO_1081 (O_1081,N_49508,N_44618);
or UO_1082 (O_1082,N_41219,N_42119);
and UO_1083 (O_1083,N_49097,N_49098);
or UO_1084 (O_1084,N_41681,N_47136);
nand UO_1085 (O_1085,N_44103,N_40207);
nand UO_1086 (O_1086,N_41000,N_41256);
nor UO_1087 (O_1087,N_43520,N_40368);
xor UO_1088 (O_1088,N_44870,N_46005);
or UO_1089 (O_1089,N_40968,N_49384);
or UO_1090 (O_1090,N_43340,N_47657);
or UO_1091 (O_1091,N_44361,N_49368);
nor UO_1092 (O_1092,N_44488,N_49854);
and UO_1093 (O_1093,N_49406,N_41513);
and UO_1094 (O_1094,N_45272,N_44539);
nor UO_1095 (O_1095,N_44857,N_46640);
nor UO_1096 (O_1096,N_48813,N_40694);
nand UO_1097 (O_1097,N_44102,N_44638);
nand UO_1098 (O_1098,N_41869,N_49643);
nor UO_1099 (O_1099,N_40054,N_44182);
nor UO_1100 (O_1100,N_44115,N_45273);
xor UO_1101 (O_1101,N_44796,N_40577);
nor UO_1102 (O_1102,N_49429,N_45921);
nand UO_1103 (O_1103,N_46391,N_41964);
nand UO_1104 (O_1104,N_47289,N_42060);
and UO_1105 (O_1105,N_40228,N_42189);
nand UO_1106 (O_1106,N_49759,N_46495);
nand UO_1107 (O_1107,N_42819,N_47478);
nand UO_1108 (O_1108,N_44511,N_47311);
or UO_1109 (O_1109,N_44172,N_45197);
nor UO_1110 (O_1110,N_41650,N_45423);
nand UO_1111 (O_1111,N_41358,N_41376);
and UO_1112 (O_1112,N_48784,N_49845);
xor UO_1113 (O_1113,N_49644,N_48632);
xor UO_1114 (O_1114,N_40459,N_40856);
or UO_1115 (O_1115,N_45961,N_47626);
nor UO_1116 (O_1116,N_46259,N_42813);
and UO_1117 (O_1117,N_43139,N_40159);
nand UO_1118 (O_1118,N_48788,N_40964);
nand UO_1119 (O_1119,N_49757,N_44657);
or UO_1120 (O_1120,N_48013,N_48580);
and UO_1121 (O_1121,N_42489,N_43054);
nand UO_1122 (O_1122,N_47557,N_48610);
and UO_1123 (O_1123,N_44634,N_49344);
or UO_1124 (O_1124,N_49723,N_43998);
nand UO_1125 (O_1125,N_46498,N_49786);
nor UO_1126 (O_1126,N_44566,N_41798);
xnor UO_1127 (O_1127,N_42265,N_47507);
xor UO_1128 (O_1128,N_44578,N_45529);
or UO_1129 (O_1129,N_43945,N_47116);
nand UO_1130 (O_1130,N_45640,N_46883);
and UO_1131 (O_1131,N_43406,N_43734);
or UO_1132 (O_1132,N_40671,N_48143);
xnor UO_1133 (O_1133,N_49112,N_47555);
nor UO_1134 (O_1134,N_40963,N_49294);
nand UO_1135 (O_1135,N_40410,N_40937);
nand UO_1136 (O_1136,N_42161,N_46277);
nor UO_1137 (O_1137,N_46528,N_40212);
nor UO_1138 (O_1138,N_41466,N_48320);
and UO_1139 (O_1139,N_45250,N_41322);
and UO_1140 (O_1140,N_42597,N_47435);
xnor UO_1141 (O_1141,N_49792,N_43683);
xor UO_1142 (O_1142,N_42148,N_40379);
nand UO_1143 (O_1143,N_46672,N_46563);
or UO_1144 (O_1144,N_41457,N_41653);
or UO_1145 (O_1145,N_40388,N_46934);
or UO_1146 (O_1146,N_41092,N_43606);
xor UO_1147 (O_1147,N_48005,N_42263);
and UO_1148 (O_1148,N_48874,N_41438);
or UO_1149 (O_1149,N_46471,N_47631);
nor UO_1150 (O_1150,N_41275,N_43460);
and UO_1151 (O_1151,N_44097,N_41670);
or UO_1152 (O_1152,N_40026,N_49592);
nor UO_1153 (O_1153,N_44059,N_40996);
xnor UO_1154 (O_1154,N_47433,N_41657);
or UO_1155 (O_1155,N_41036,N_46697);
or UO_1156 (O_1156,N_44334,N_42191);
nand UO_1157 (O_1157,N_41430,N_45334);
or UO_1158 (O_1158,N_42034,N_40688);
xnor UO_1159 (O_1159,N_42354,N_47485);
and UO_1160 (O_1160,N_41138,N_40944);
and UO_1161 (O_1161,N_48240,N_47825);
nand UO_1162 (O_1162,N_45343,N_47055);
and UO_1163 (O_1163,N_40002,N_47749);
nand UO_1164 (O_1164,N_45948,N_48630);
or UO_1165 (O_1165,N_40078,N_42032);
or UO_1166 (O_1166,N_43120,N_45039);
and UO_1167 (O_1167,N_42528,N_49505);
xnor UO_1168 (O_1168,N_40812,N_45853);
or UO_1169 (O_1169,N_45999,N_46202);
xor UO_1170 (O_1170,N_49405,N_40824);
nand UO_1171 (O_1171,N_41635,N_44946);
and UO_1172 (O_1172,N_42343,N_43352);
nand UO_1173 (O_1173,N_41273,N_49982);
xnor UO_1174 (O_1174,N_48380,N_46838);
nand UO_1175 (O_1175,N_43548,N_46328);
or UO_1176 (O_1176,N_48597,N_45407);
nand UO_1177 (O_1177,N_44365,N_42192);
xor UO_1178 (O_1178,N_46015,N_48883);
nand UO_1179 (O_1179,N_49684,N_43053);
or UO_1180 (O_1180,N_45957,N_48667);
or UO_1181 (O_1181,N_49543,N_45525);
and UO_1182 (O_1182,N_47092,N_47609);
nand UO_1183 (O_1183,N_40480,N_40612);
or UO_1184 (O_1184,N_45333,N_42603);
xor UO_1185 (O_1185,N_41184,N_41147);
nand UO_1186 (O_1186,N_40433,N_41375);
nor UO_1187 (O_1187,N_47340,N_43077);
and UO_1188 (O_1188,N_41601,N_41744);
nor UO_1189 (O_1189,N_44333,N_48384);
nor UO_1190 (O_1190,N_49156,N_47452);
nor UO_1191 (O_1191,N_42624,N_41064);
and UO_1192 (O_1192,N_48657,N_44607);
xnor UO_1193 (O_1193,N_44008,N_45372);
nand UO_1194 (O_1194,N_43511,N_41034);
nand UO_1195 (O_1195,N_41626,N_45709);
and UO_1196 (O_1196,N_47183,N_45993);
xor UO_1197 (O_1197,N_42596,N_43018);
nand UO_1198 (O_1198,N_47709,N_41753);
nand UO_1199 (O_1199,N_47001,N_46558);
xnor UO_1200 (O_1200,N_41540,N_45279);
xnor UO_1201 (O_1201,N_42373,N_43941);
or UO_1202 (O_1202,N_48839,N_46676);
nand UO_1203 (O_1203,N_41720,N_46427);
nor UO_1204 (O_1204,N_40837,N_49411);
or UO_1205 (O_1205,N_40553,N_40259);
nand UO_1206 (O_1206,N_43509,N_45196);
or UO_1207 (O_1207,N_45003,N_41515);
nor UO_1208 (O_1208,N_42922,N_40253);
and UO_1209 (O_1209,N_47917,N_40087);
nor UO_1210 (O_1210,N_46130,N_47034);
or UO_1211 (O_1211,N_48541,N_48531);
xor UO_1212 (O_1212,N_47902,N_49914);
nand UO_1213 (O_1213,N_45875,N_46511);
nor UO_1214 (O_1214,N_43052,N_48392);
xnor UO_1215 (O_1215,N_40945,N_46115);
nand UO_1216 (O_1216,N_46644,N_40700);
xnor UO_1217 (O_1217,N_45603,N_44429);
nor UO_1218 (O_1218,N_47295,N_45416);
or UO_1219 (O_1219,N_47924,N_43634);
xor UO_1220 (O_1220,N_40749,N_42551);
nand UO_1221 (O_1221,N_49793,N_47235);
nor UO_1222 (O_1222,N_49200,N_42602);
xnor UO_1223 (O_1223,N_42526,N_48893);
or UO_1224 (O_1224,N_45456,N_48229);
and UO_1225 (O_1225,N_48428,N_44809);
xor UO_1226 (O_1226,N_48418,N_47135);
and UO_1227 (O_1227,N_44427,N_49551);
nand UO_1228 (O_1228,N_42868,N_43981);
xor UO_1229 (O_1229,N_40622,N_45455);
or UO_1230 (O_1230,N_40328,N_40784);
nor UO_1231 (O_1231,N_47875,N_47290);
xor UO_1232 (O_1232,N_45780,N_40726);
and UO_1233 (O_1233,N_45833,N_45740);
and UO_1234 (O_1234,N_43842,N_40312);
or UO_1235 (O_1235,N_42501,N_44044);
nor UO_1236 (O_1236,N_47861,N_45153);
xnor UO_1237 (O_1237,N_49741,N_49638);
nand UO_1238 (O_1238,N_48700,N_46541);
nand UO_1239 (O_1239,N_46429,N_43165);
xor UO_1240 (O_1240,N_42792,N_47224);
and UO_1241 (O_1241,N_41021,N_42203);
nor UO_1242 (O_1242,N_49347,N_48084);
xnor UO_1243 (O_1243,N_47839,N_45368);
and UO_1244 (O_1244,N_48738,N_42788);
nor UO_1245 (O_1245,N_49947,N_44332);
xnor UO_1246 (O_1246,N_46281,N_40709);
xor UO_1247 (O_1247,N_47247,N_41178);
and UO_1248 (O_1248,N_47385,N_45735);
nor UO_1249 (O_1249,N_48978,N_48129);
or UO_1250 (O_1250,N_46984,N_45839);
nand UO_1251 (O_1251,N_49511,N_43716);
nand UO_1252 (O_1252,N_48308,N_45599);
nand UO_1253 (O_1253,N_40760,N_48553);
xnor UO_1254 (O_1254,N_49367,N_42423);
xnor UO_1255 (O_1255,N_40846,N_43448);
and UO_1256 (O_1256,N_46302,N_48513);
xor UO_1257 (O_1257,N_49094,N_47710);
and UO_1258 (O_1258,N_42975,N_45373);
nand UO_1259 (O_1259,N_46369,N_46872);
nand UO_1260 (O_1260,N_41418,N_46865);
xnor UO_1261 (O_1261,N_46562,N_48059);
xnor UO_1262 (O_1262,N_47652,N_46336);
nand UO_1263 (O_1263,N_46661,N_47964);
or UO_1264 (O_1264,N_42426,N_49996);
xnor UO_1265 (O_1265,N_48638,N_47284);
or UO_1266 (O_1266,N_41450,N_41770);
nand UO_1267 (O_1267,N_47679,N_48622);
and UO_1268 (O_1268,N_46760,N_41905);
nand UO_1269 (O_1269,N_46207,N_49633);
and UO_1270 (O_1270,N_48546,N_42045);
nor UO_1271 (O_1271,N_42839,N_42572);
and UO_1272 (O_1272,N_40746,N_41218);
and UO_1273 (O_1273,N_45617,N_47441);
xnor UO_1274 (O_1274,N_44437,N_40893);
nor UO_1275 (O_1275,N_44956,N_41172);
nor UO_1276 (O_1276,N_40189,N_49648);
xor UO_1277 (O_1277,N_42347,N_45543);
and UO_1278 (O_1278,N_40302,N_47443);
and UO_1279 (O_1279,N_47939,N_46585);
nand UO_1280 (O_1280,N_47190,N_43626);
nand UO_1281 (O_1281,N_49230,N_46497);
nor UO_1282 (O_1282,N_48646,N_46340);
nor UO_1283 (O_1283,N_41651,N_47656);
or UO_1284 (O_1284,N_43075,N_45586);
or UO_1285 (O_1285,N_44298,N_41927);
nor UO_1286 (O_1286,N_48944,N_43545);
and UO_1287 (O_1287,N_42697,N_44632);
nand UO_1288 (O_1288,N_43875,N_42934);
and UO_1289 (O_1289,N_40984,N_42483);
and UO_1290 (O_1290,N_49151,N_44208);
nand UO_1291 (O_1291,N_41066,N_44667);
nand UO_1292 (O_1292,N_44032,N_42174);
nand UO_1293 (O_1293,N_42283,N_42911);
nand UO_1294 (O_1294,N_41655,N_43624);
nor UO_1295 (O_1295,N_47793,N_44831);
nor UO_1296 (O_1296,N_49482,N_43373);
or UO_1297 (O_1297,N_45223,N_48888);
nor UO_1298 (O_1298,N_49801,N_43675);
xor UO_1299 (O_1299,N_47411,N_40151);
xnor UO_1300 (O_1300,N_43289,N_43777);
and UO_1301 (O_1301,N_46986,N_46165);
xnor UO_1302 (O_1302,N_43358,N_48620);
nand UO_1303 (O_1303,N_40096,N_48092);
nand UO_1304 (O_1304,N_45828,N_49221);
xor UO_1305 (O_1305,N_42443,N_41247);
nand UO_1306 (O_1306,N_47573,N_45047);
nand UO_1307 (O_1307,N_46449,N_42589);
nor UO_1308 (O_1308,N_46902,N_40737);
xnor UO_1309 (O_1309,N_48820,N_45099);
or UO_1310 (O_1310,N_46907,N_41553);
and UO_1311 (O_1311,N_42816,N_49549);
nand UO_1312 (O_1312,N_43462,N_47647);
nand UO_1313 (O_1313,N_47726,N_47695);
nor UO_1314 (O_1314,N_41459,N_47623);
and UO_1315 (O_1315,N_43882,N_45194);
nand UO_1316 (O_1316,N_41334,N_49301);
nor UO_1317 (O_1317,N_43952,N_48641);
or UO_1318 (O_1318,N_46067,N_42109);
and UO_1319 (O_1319,N_41743,N_42400);
or UO_1320 (O_1320,N_45625,N_42635);
nor UO_1321 (O_1321,N_42646,N_42710);
or UO_1322 (O_1322,N_46203,N_41410);
and UO_1323 (O_1323,N_48999,N_41901);
or UO_1324 (O_1324,N_43692,N_48837);
nand UO_1325 (O_1325,N_44635,N_42590);
nand UO_1326 (O_1326,N_48890,N_44747);
nor UO_1327 (O_1327,N_49334,N_47423);
nand UO_1328 (O_1328,N_44127,N_41191);
or UO_1329 (O_1329,N_45621,N_44204);
nor UO_1330 (O_1330,N_46124,N_44043);
nor UO_1331 (O_1331,N_40286,N_49890);
xor UO_1332 (O_1332,N_47702,N_45958);
xnor UO_1333 (O_1333,N_47331,N_49769);
and UO_1334 (O_1334,N_42721,N_47354);
and UO_1335 (O_1335,N_42775,N_40512);
nor UO_1336 (O_1336,N_44974,N_46403);
xor UO_1337 (O_1337,N_43374,N_44523);
xnor UO_1338 (O_1338,N_48056,N_47852);
xnor UO_1339 (O_1339,N_41760,N_41751);
nor UO_1340 (O_1340,N_48435,N_43224);
nor UO_1341 (O_1341,N_48395,N_49576);
and UO_1342 (O_1342,N_45637,N_46472);
xor UO_1343 (O_1343,N_47547,N_42749);
nor UO_1344 (O_1344,N_48750,N_46454);
nand UO_1345 (O_1345,N_48752,N_48260);
and UO_1346 (O_1346,N_47538,N_42842);
and UO_1347 (O_1347,N_44816,N_47477);
nand UO_1348 (O_1348,N_42326,N_42657);
nand UO_1349 (O_1349,N_48307,N_48727);
xnor UO_1350 (O_1350,N_41475,N_40559);
and UO_1351 (O_1351,N_41362,N_42692);
nor UO_1352 (O_1352,N_43194,N_42601);
nor UO_1353 (O_1353,N_43583,N_48406);
nor UO_1354 (O_1354,N_45002,N_41896);
nand UO_1355 (O_1355,N_43898,N_47167);
or UO_1356 (O_1356,N_45602,N_42091);
xor UO_1357 (O_1357,N_47750,N_47422);
nand UO_1358 (O_1358,N_46629,N_46973);
xor UO_1359 (O_1359,N_46945,N_42982);
and UO_1360 (O_1360,N_47061,N_45770);
xnor UO_1361 (O_1361,N_48605,N_43825);
and UO_1362 (O_1362,N_49142,N_48467);
xnor UO_1363 (O_1363,N_45626,N_48098);
nor UO_1364 (O_1364,N_40091,N_47160);
xor UO_1365 (O_1365,N_42260,N_43068);
and UO_1366 (O_1366,N_46151,N_46190);
and UO_1367 (O_1367,N_48412,N_42087);
nand UO_1368 (O_1368,N_42270,N_42335);
and UO_1369 (O_1369,N_40101,N_42632);
nand UO_1370 (O_1370,N_43094,N_49817);
xnor UO_1371 (O_1371,N_47534,N_47966);
nor UO_1372 (O_1372,N_44416,N_41268);
xnor UO_1373 (O_1373,N_45872,N_47130);
xor UO_1374 (O_1374,N_42509,N_48939);
nor UO_1375 (O_1375,N_41449,N_45218);
and UO_1376 (O_1376,N_49676,N_49660);
xnor UO_1377 (O_1377,N_48015,N_40439);
xor UO_1378 (O_1378,N_40075,N_45315);
xor UO_1379 (O_1379,N_45836,N_49400);
and UO_1380 (O_1380,N_47230,N_40627);
xnor UO_1381 (O_1381,N_44387,N_43950);
and UO_1382 (O_1382,N_49350,N_45507);
nor UO_1383 (O_1383,N_47417,N_46386);
xor UO_1384 (O_1384,N_40341,N_44909);
xnor UO_1385 (O_1385,N_42452,N_43335);
or UO_1386 (O_1386,N_40855,N_49446);
nand UO_1387 (O_1387,N_44278,N_47042);
and UO_1388 (O_1388,N_47771,N_42019);
and UO_1389 (O_1389,N_43956,N_44853);
and UO_1390 (O_1390,N_43695,N_46227);
nor UO_1391 (O_1391,N_43754,N_46291);
and UO_1392 (O_1392,N_43962,N_41826);
and UO_1393 (O_1393,N_43126,N_48268);
and UO_1394 (O_1394,N_40456,N_44475);
or UO_1395 (O_1395,N_42222,N_47984);
nand UO_1396 (O_1396,N_44439,N_44372);
nor UO_1397 (O_1397,N_48524,N_44491);
or UO_1398 (O_1398,N_48627,N_43301);
xnor UO_1399 (O_1399,N_47929,N_48267);
xnor UO_1400 (O_1400,N_49223,N_48997);
nor UO_1401 (O_1401,N_41434,N_46844);
xor UO_1402 (O_1402,N_41800,N_40747);
nor UO_1403 (O_1403,N_41976,N_46343);
nand UO_1404 (O_1404,N_43078,N_48991);
nor UO_1405 (O_1405,N_47845,N_47355);
xnor UO_1406 (O_1406,N_46145,N_48312);
nand UO_1407 (O_1407,N_42620,N_48884);
or UO_1408 (O_1408,N_44083,N_47583);
or UO_1409 (O_1409,N_40072,N_46418);
nand UO_1410 (O_1410,N_43512,N_42357);
or UO_1411 (O_1411,N_45187,N_45558);
and UO_1412 (O_1412,N_44047,N_43492);
and UO_1413 (O_1413,N_43911,N_47625);
xnor UO_1414 (O_1414,N_42815,N_46841);
nor UO_1415 (O_1415,N_47365,N_41712);
or UO_1416 (O_1416,N_49155,N_47421);
nand UO_1417 (O_1417,N_42583,N_40609);
nor UO_1418 (O_1418,N_46856,N_40637);
nand UO_1419 (O_1419,N_48449,N_45213);
nor UO_1420 (O_1420,N_40931,N_47343);
nor UO_1421 (O_1421,N_48755,N_46506);
nand UO_1422 (O_1422,N_41462,N_47858);
nor UO_1423 (O_1423,N_42743,N_48053);
or UO_1424 (O_1424,N_44272,N_46318);
and UO_1425 (O_1425,N_42987,N_40051);
and UO_1426 (O_1426,N_46522,N_47301);
xor UO_1427 (O_1427,N_44832,N_42385);
and UO_1428 (O_1428,N_40924,N_46749);
or UO_1429 (O_1429,N_49671,N_45703);
nor UO_1430 (O_1430,N_45125,N_46109);
nand UO_1431 (O_1431,N_40130,N_41629);
nor UO_1432 (O_1432,N_49460,N_40550);
nand UO_1433 (O_1433,N_45025,N_42063);
nor UO_1434 (O_1434,N_45462,N_47306);
or UO_1435 (O_1435,N_45342,N_44840);
or UO_1436 (O_1436,N_43445,N_44683);
nand UO_1437 (O_1437,N_48711,N_44223);
and UO_1438 (O_1438,N_43089,N_49289);
and UO_1439 (O_1439,N_41806,N_46473);
nor UO_1440 (O_1440,N_45101,N_44370);
nand UO_1441 (O_1441,N_48873,N_47002);
or UO_1442 (O_1442,N_48273,N_41113);
xor UO_1443 (O_1443,N_49779,N_45873);
nor UO_1444 (O_1444,N_41159,N_46719);
and UO_1445 (O_1445,N_48940,N_43758);
and UO_1446 (O_1446,N_45367,N_49271);
nor UO_1447 (O_1447,N_47872,N_48761);
or UO_1448 (O_1448,N_46839,N_48185);
nand UO_1449 (O_1449,N_46357,N_47143);
nand UO_1450 (O_1450,N_45078,N_41962);
or UO_1451 (O_1451,N_45754,N_46951);
and UO_1452 (O_1452,N_44245,N_46767);
or UO_1453 (O_1453,N_42731,N_45227);
xor UO_1454 (O_1454,N_42459,N_43403);
nor UO_1455 (O_1455,N_44848,N_48266);
nor UO_1456 (O_1456,N_43091,N_48880);
nor UO_1457 (O_1457,N_48479,N_49000);
nor UO_1458 (O_1458,N_48445,N_47108);
or UO_1459 (O_1459,N_42333,N_45777);
or UO_1460 (O_1460,N_41799,N_42789);
nand UO_1461 (O_1461,N_40766,N_43324);
and UO_1462 (O_1462,N_40371,N_44757);
nand UO_1463 (O_1463,N_49434,N_49138);
nor UO_1464 (O_1464,N_47481,N_42090);
and UO_1465 (O_1465,N_48352,N_48049);
nand UO_1466 (O_1466,N_45612,N_49661);
nor UO_1467 (O_1467,N_49234,N_43360);
nand UO_1468 (O_1468,N_49754,N_42419);
xor UO_1469 (O_1469,N_42022,N_49844);
xnor UO_1470 (O_1470,N_48668,N_45897);
nand UO_1471 (O_1471,N_40170,N_40181);
or UO_1472 (O_1472,N_45459,N_43523);
or UO_1473 (O_1473,N_44587,N_41547);
nand UO_1474 (O_1474,N_47399,N_49217);
and UO_1475 (O_1475,N_47713,N_46593);
or UO_1476 (O_1476,N_41882,N_41959);
or UO_1477 (O_1477,N_48359,N_45616);
xnor UO_1478 (O_1478,N_45949,N_49247);
nor UO_1479 (O_1479,N_48721,N_45141);
and UO_1480 (O_1480,N_46305,N_49435);
or UO_1481 (O_1481,N_45204,N_46117);
and UO_1482 (O_1482,N_49017,N_43148);
xor UO_1483 (O_1483,N_41813,N_46198);
xor UO_1484 (O_1484,N_49180,N_41497);
nand UO_1485 (O_1485,N_47587,N_45018);
or UO_1486 (O_1486,N_45647,N_40995);
nand UO_1487 (O_1487,N_45846,N_45970);
xor UO_1488 (O_1488,N_40222,N_49236);
xor UO_1489 (O_1489,N_40708,N_42009);
xnor UO_1490 (O_1490,N_47720,N_43665);
nand UO_1491 (O_1491,N_42103,N_47159);
xnor UO_1492 (O_1492,N_43927,N_49278);
nand UO_1493 (O_1493,N_45112,N_48542);
and UO_1494 (O_1494,N_41244,N_48426);
nand UO_1495 (O_1495,N_44054,N_44093);
or UO_1496 (O_1496,N_44981,N_46114);
xnor UO_1497 (O_1497,N_45849,N_44714);
xnor UO_1498 (O_1498,N_48492,N_46101);
xnor UO_1499 (O_1499,N_49392,N_44979);
nand UO_1500 (O_1500,N_47940,N_48796);
or UO_1501 (O_1501,N_45741,N_48521);
or UO_1502 (O_1502,N_44811,N_46460);
xnor UO_1503 (O_1503,N_48608,N_44868);
nand UO_1504 (O_1504,N_44827,N_44470);
nand UO_1505 (O_1505,N_41354,N_48810);
nand UO_1506 (O_1506,N_40952,N_45983);
or UO_1507 (O_1507,N_42499,N_44450);
nor UO_1508 (O_1508,N_48210,N_47013);
nand UO_1509 (O_1509,N_42269,N_44712);
or UO_1510 (O_1510,N_40703,N_43110);
xor UO_1511 (O_1511,N_47038,N_44616);
nor UO_1512 (O_1512,N_42618,N_40641);
or UO_1513 (O_1513,N_46782,N_40385);
and UO_1514 (O_1514,N_49361,N_48152);
and UO_1515 (O_1515,N_41198,N_46621);
nor UO_1516 (O_1516,N_40965,N_43323);
nor UO_1517 (O_1517,N_44473,N_45313);
or UO_1518 (O_1518,N_44818,N_46701);
or UO_1519 (O_1519,N_41259,N_41062);
or UO_1520 (O_1520,N_49509,N_46422);
nor UO_1521 (O_1521,N_41879,N_41310);
nor UO_1522 (O_1522,N_41248,N_41300);
nor UO_1523 (O_1523,N_42367,N_41565);
nor UO_1524 (O_1524,N_44744,N_40651);
or UO_1525 (O_1525,N_49568,N_47472);
nor UO_1526 (O_1526,N_43772,N_45515);
and UO_1527 (O_1527,N_42729,N_47667);
nor UO_1528 (O_1528,N_42202,N_42378);
or UO_1529 (O_1529,N_43349,N_46923);
or UO_1530 (O_1530,N_46887,N_46740);
nand UO_1531 (O_1531,N_41592,N_42709);
nand UO_1532 (O_1532,N_44401,N_40569);
nand UO_1533 (O_1533,N_42629,N_49006);
nor UO_1534 (O_1534,N_42224,N_43048);
nand UO_1535 (O_1535,N_48992,N_41078);
and UO_1536 (O_1536,N_45086,N_41007);
or UO_1537 (O_1537,N_46375,N_46531);
xor UO_1538 (O_1538,N_44874,N_43069);
nand UO_1539 (O_1539,N_48288,N_47565);
nor UO_1540 (O_1540,N_40979,N_43164);
or UO_1541 (O_1541,N_46540,N_49239);
xnor UO_1542 (O_1542,N_47357,N_40408);
nor UO_1543 (O_1543,N_43044,N_40382);
xnor UO_1544 (O_1544,N_44329,N_45166);
nor UO_1545 (O_1545,N_41320,N_41352);
nand UO_1546 (O_1546,N_41864,N_40572);
xnor UO_1547 (O_1547,N_41235,N_48574);
xnor UO_1548 (O_1548,N_40082,N_40544);
or UO_1549 (O_1549,N_48941,N_44358);
nand UO_1550 (O_1550,N_40625,N_49735);
nand UO_1551 (O_1551,N_42312,N_49809);
xor UO_1552 (O_1552,N_45739,N_47204);
nand UO_1553 (O_1553,N_45814,N_46657);
nor UO_1554 (O_1554,N_43848,N_47244);
and UO_1555 (O_1555,N_42647,N_45306);
nor UO_1556 (O_1556,N_45157,N_46307);
xor UO_1557 (O_1557,N_47461,N_48551);
nor UO_1558 (O_1558,N_45133,N_49363);
nor UO_1559 (O_1559,N_49162,N_40364);
xnor UO_1560 (O_1560,N_49773,N_49136);
or UO_1561 (O_1561,N_47278,N_44845);
and UO_1562 (O_1562,N_44189,N_49106);
nor UO_1563 (O_1563,N_47299,N_41239);
or UO_1564 (O_1564,N_46779,N_47179);
nand UO_1565 (O_1565,N_48726,N_49283);
nand UO_1566 (O_1566,N_45487,N_49874);
nand UO_1567 (O_1567,N_44993,N_45052);
nand UO_1568 (O_1568,N_49740,N_49550);
or UO_1569 (O_1569,N_49373,N_45807);
nor UO_1570 (O_1570,N_44558,N_45077);
and UO_1571 (O_1571,N_43647,N_47738);
and UO_1572 (O_1572,N_41135,N_47641);
xor UO_1573 (O_1573,N_44734,N_45955);
xor UO_1574 (O_1574,N_43565,N_49978);
or UO_1575 (O_1575,N_42159,N_45095);
and UO_1576 (O_1576,N_46499,N_44524);
and UO_1577 (O_1577,N_43759,N_49144);
or UO_1578 (O_1578,N_40508,N_46519);
nor UO_1579 (O_1579,N_41900,N_45221);
or UO_1580 (O_1580,N_44380,N_42237);
nor UO_1581 (O_1581,N_40019,N_42652);
or UO_1582 (O_1582,N_48698,N_48847);
xnor UO_1583 (O_1583,N_47363,N_43544);
nor UO_1584 (O_1584,N_41940,N_43332);
xor UO_1585 (O_1585,N_45877,N_48048);
xnor UO_1586 (O_1586,N_41516,N_48664);
xor UO_1587 (O_1587,N_44485,N_42448);
nand UO_1588 (O_1588,N_41522,N_40432);
and UO_1589 (O_1589,N_44149,N_48554);
nor UO_1590 (O_1590,N_41649,N_49248);
or UO_1591 (O_1591,N_41688,N_47988);
xor UO_1592 (O_1592,N_44277,N_40642);
and UO_1593 (O_1593,N_43543,N_45063);
nand UO_1594 (O_1594,N_47847,N_48737);
and UO_1595 (O_1595,N_47892,N_42310);
and UO_1596 (O_1596,N_45559,N_45827);
nand UO_1597 (O_1597,N_44567,N_49064);
nor UO_1598 (O_1598,N_49461,N_42231);
and UO_1599 (O_1599,N_45300,N_46953);
xnor UO_1600 (O_1600,N_41956,N_49477);
or UO_1601 (O_1601,N_46235,N_41856);
or UO_1602 (O_1602,N_48057,N_47700);
xor UO_1603 (O_1603,N_41749,N_48929);
nand UO_1604 (O_1604,N_46345,N_45686);
nor UO_1605 (O_1605,N_44480,N_42857);
xor UO_1606 (O_1606,N_41966,N_45606);
and UO_1607 (O_1607,N_47491,N_45518);
nor UO_1608 (O_1608,N_40160,N_49202);
nand UO_1609 (O_1609,N_46214,N_49485);
nor UO_1610 (O_1610,N_43686,N_40848);
and UO_1611 (O_1611,N_41237,N_47490);
nand UO_1612 (O_1612,N_44307,N_43541);
nor UO_1613 (O_1613,N_45657,N_45257);
nand UO_1614 (O_1614,N_45500,N_41225);
xor UO_1615 (O_1615,N_43480,N_46168);
nor UO_1616 (O_1616,N_45998,N_49925);
nand UO_1617 (O_1617,N_45685,N_43904);
nor UO_1618 (O_1618,N_41979,N_41416);
xnor UO_1619 (O_1619,N_40827,N_41880);
or UO_1620 (O_1620,N_47802,N_42212);
xor UO_1621 (O_1621,N_44294,N_49697);
or UO_1622 (O_1622,N_49980,N_43645);
nand UO_1623 (O_1623,N_47119,N_43598);
or UO_1624 (O_1624,N_40155,N_43574);
and UO_1625 (O_1625,N_45782,N_48830);
xnor UO_1626 (O_1626,N_40462,N_44222);
or UO_1627 (O_1627,N_42515,N_44364);
nor UO_1628 (O_1628,N_46053,N_40663);
or UO_1629 (O_1629,N_42565,N_43639);
nor UO_1630 (O_1630,N_48733,N_46914);
nor UO_1631 (O_1631,N_40421,N_48540);
and UO_1632 (O_1632,N_40730,N_46197);
xor UO_1633 (O_1633,N_48114,N_42180);
and UO_1634 (O_1634,N_48821,N_46033);
and UO_1635 (O_1635,N_43405,N_44359);
nand UO_1636 (O_1636,N_41595,N_43837);
nor UO_1637 (O_1637,N_42621,N_49953);
xnor UO_1638 (O_1638,N_41771,N_49224);
xnor UO_1639 (O_1639,N_46002,N_41243);
xnor UO_1640 (O_1640,N_41661,N_47377);
and UO_1641 (O_1641,N_40980,N_43551);
and UO_1642 (O_1642,N_40114,N_48705);
nand UO_1643 (O_1643,N_49607,N_49530);
xnor UO_1644 (O_1644,N_46264,N_43910);
xnor UO_1645 (O_1645,N_46315,N_46024);
nor UO_1646 (O_1646,N_47402,N_47927);
nor UO_1647 (O_1647,N_45567,N_40123);
xor UO_1648 (O_1648,N_47439,N_47889);
and UO_1649 (O_1649,N_42904,N_48478);
xnor UO_1650 (O_1650,N_40613,N_49781);
or UO_1651 (O_1651,N_46035,N_43693);
or UO_1652 (O_1652,N_49343,N_43940);
nand UO_1653 (O_1653,N_48555,N_49108);
nor UO_1654 (O_1654,N_44756,N_48658);
or UO_1655 (O_1655,N_42947,N_45854);
or UO_1656 (O_1656,N_42125,N_41919);
nor UO_1657 (O_1657,N_44593,N_44466);
or UO_1658 (O_1658,N_42990,N_48047);
nand UO_1659 (O_1659,N_43566,N_46309);
and UO_1660 (O_1660,N_44897,N_44252);
nand UO_1661 (O_1661,N_46037,N_48339);
and UO_1662 (O_1662,N_46855,N_49412);
or UO_1663 (O_1663,N_47302,N_46379);
nand UO_1664 (O_1664,N_40427,N_44453);
or UO_1665 (O_1665,N_44600,N_44864);
or UO_1666 (O_1666,N_40702,N_46447);
or UO_1667 (O_1667,N_49454,N_49005);
and UO_1668 (O_1668,N_45268,N_44455);
nor UO_1669 (O_1669,N_42033,N_49946);
and UO_1670 (O_1670,N_49131,N_45426);
nor UO_1671 (O_1671,N_44468,N_48846);
and UO_1672 (O_1672,N_46356,N_40167);
and UO_1673 (O_1673,N_44226,N_44396);
and UO_1674 (O_1674,N_44905,N_41463);
xnor UO_1675 (O_1675,N_42680,N_45397);
xor UO_1676 (O_1676,N_49072,N_47761);
and UO_1677 (O_1677,N_48009,N_49843);
xor UO_1678 (O_1678,N_43337,N_44271);
xor UO_1679 (O_1679,N_41586,N_46394);
nor UO_1680 (O_1680,N_41678,N_46787);
nand UO_1681 (O_1681,N_47683,N_47595);
nor UO_1682 (O_1682,N_42720,N_48533);
or UO_1683 (O_1683,N_42445,N_43387);
nand UO_1684 (O_1684,N_40291,N_49823);
or UO_1685 (O_1685,N_48675,N_45176);
or UO_1686 (O_1686,N_42580,N_43211);
and UO_1687 (O_1687,N_43277,N_45238);
and UO_1688 (O_1688,N_44598,N_41045);
nor UO_1689 (O_1689,N_48438,N_42676);
or UO_1690 (O_1690,N_40474,N_43336);
nor UO_1691 (O_1691,N_41454,N_42020);
nor UO_1692 (O_1692,N_47920,N_43055);
nand UO_1693 (O_1693,N_40386,N_43542);
or UO_1694 (O_1694,N_49266,N_47531);
or UO_1695 (O_1695,N_40004,N_49877);
nand UO_1696 (O_1696,N_40305,N_46459);
nor UO_1697 (O_1697,N_46975,N_49991);
or UO_1698 (O_1698,N_45215,N_46226);
nor UO_1699 (O_1699,N_42735,N_42441);
xnor UO_1700 (O_1700,N_49250,N_41123);
or UO_1701 (O_1701,N_40551,N_46965);
xnor UO_1702 (O_1702,N_43086,N_44859);
nand UO_1703 (O_1703,N_49268,N_43810);
xor UO_1704 (O_1704,N_40434,N_42467);
or UO_1705 (O_1705,N_46267,N_48254);
and UO_1706 (O_1706,N_48624,N_47464);
nand UO_1707 (O_1707,N_46550,N_43711);
xnor UO_1708 (O_1708,N_41909,N_42866);
nand UO_1709 (O_1709,N_43868,N_40861);
and UO_1710 (O_1710,N_41492,N_40306);
nor UO_1711 (O_1711,N_46107,N_42616);
and UO_1712 (O_1712,N_48947,N_43266);
xnor UO_1713 (O_1713,N_43615,N_48074);
nand UO_1714 (O_1714,N_40959,N_45928);
nand UO_1715 (O_1715,N_41929,N_45069);
or UO_1716 (O_1716,N_41313,N_47168);
nor UO_1717 (O_1717,N_46875,N_46348);
or UO_1718 (O_1718,N_42936,N_49702);
nand UO_1719 (O_1719,N_43864,N_44006);
and UO_1720 (O_1720,N_45929,N_40639);
and UO_1721 (O_1721,N_48594,N_48115);
or UO_1722 (O_1722,N_42540,N_48315);
nor UO_1723 (O_1723,N_40424,N_42916);
nor UO_1724 (O_1724,N_45680,N_49683);
nand UO_1725 (O_1725,N_42542,N_47960);
xnor UO_1726 (O_1726,N_47516,N_49322);
xor UO_1727 (O_1727,N_42268,N_47081);
xor UO_1728 (O_1728,N_47073,N_45860);
or UO_1729 (O_1729,N_43193,N_45163);
and UO_1730 (O_1730,N_47029,N_49897);
xor UO_1731 (O_1731,N_43296,N_48872);
nand UO_1732 (O_1732,N_46397,N_48455);
xor UO_1733 (O_1733,N_47559,N_41584);
nand UO_1734 (O_1734,N_41756,N_42256);
or UO_1735 (O_1735,N_48297,N_49657);
nand UO_1736 (O_1736,N_47946,N_41511);
or UO_1737 (O_1737,N_45329,N_45220);
nand UO_1738 (O_1738,N_42303,N_43562);
and UO_1739 (O_1739,N_49940,N_45199);
xor UO_1740 (O_1740,N_46553,N_45005);
or UO_1741 (O_1741,N_40854,N_47156);
xnor UO_1742 (O_1742,N_41541,N_46162);
and UO_1743 (O_1743,N_42663,N_40047);
nor UO_1744 (O_1744,N_43174,N_40949);
and UO_1745 (O_1745,N_42840,N_43012);
and UO_1746 (O_1746,N_43899,N_47773);
and UO_1747 (O_1747,N_48027,N_43206);
and UO_1748 (O_1748,N_43715,N_48138);
and UO_1749 (O_1749,N_47746,N_44975);
xor UO_1750 (O_1750,N_42077,N_40971);
nor UO_1751 (O_1751,N_43701,N_47805);
or UO_1752 (O_1752,N_47590,N_48485);
nand UO_1753 (O_1753,N_47214,N_40389);
and UO_1754 (O_1754,N_40751,N_40473);
and UO_1755 (O_1755,N_42059,N_41790);
nand UO_1756 (O_1756,N_46161,N_41033);
xnor UO_1757 (O_1757,N_42767,N_43158);
nand UO_1758 (O_1758,N_41131,N_45432);
or UO_1759 (O_1759,N_48552,N_43473);
nand UO_1760 (O_1760,N_40273,N_47494);
nor UO_1761 (O_1761,N_40412,N_46485);
nor UO_1762 (O_1762,N_47899,N_48457);
or UO_1763 (O_1763,N_48699,N_41179);
nand UO_1764 (O_1764,N_48295,N_44056);
nand UO_1765 (O_1765,N_46150,N_45848);
xnor UO_1766 (O_1766,N_48629,N_40632);
or UO_1767 (O_1767,N_45914,N_43182);
or UO_1768 (O_1768,N_42567,N_43354);
nand UO_1769 (O_1769,N_40863,N_41668);
nor UO_1770 (O_1770,N_41194,N_48142);
nor UO_1771 (O_1771,N_40333,N_45219);
and UO_1772 (O_1772,N_47553,N_41188);
xnor UO_1773 (O_1773,N_40050,N_49811);
xor UO_1774 (O_1774,N_45613,N_41923);
and UO_1775 (O_1775,N_47781,N_45253);
xnor UO_1776 (O_1776,N_45553,N_40762);
and UO_1777 (O_1777,N_41296,N_40196);
nand UO_1778 (O_1778,N_41993,N_49356);
and UO_1779 (O_1779,N_41220,N_44474);
or UO_1780 (O_1780,N_41386,N_40587);
and UO_1781 (O_1781,N_47074,N_40258);
xor UO_1782 (O_1782,N_42454,N_46308);
nor UO_1783 (O_1783,N_46916,N_44079);
xor UO_1784 (O_1784,N_45598,N_48549);
and UO_1785 (O_1785,N_42864,N_44264);
nand UO_1786 (O_1786,N_43887,N_45021);
xor UO_1787 (O_1787,N_40536,N_45266);
and UO_1788 (O_1788,N_42254,N_49573);
and UO_1789 (O_1789,N_43414,N_43955);
nand UO_1790 (O_1790,N_41715,N_46894);
nand UO_1791 (O_1791,N_47078,N_47996);
xnor UO_1792 (O_1792,N_48099,N_40722);
nor UO_1793 (O_1793,N_49158,N_48055);
and UO_1794 (O_1794,N_41023,N_47722);
xor UO_1795 (O_1795,N_40543,N_40510);
and UO_1796 (O_1796,N_41371,N_47841);
xor UO_1797 (O_1797,N_49442,N_46861);
nand UO_1798 (O_1798,N_40365,N_41904);
nand UO_1799 (O_1799,N_41842,N_44943);
or UO_1800 (O_1800,N_42188,N_40133);
xnor UO_1801 (O_1801,N_45696,N_41664);
or UO_1802 (O_1802,N_49420,N_44050);
xor UO_1803 (O_1803,N_46113,N_40310);
or UO_1804 (O_1804,N_47755,N_40877);
nor UO_1805 (O_1805,N_49992,N_47053);
xor UO_1806 (O_1806,N_44703,N_46075);
and UO_1807 (O_1807,N_40885,N_42345);
and UO_1808 (O_1808,N_47848,N_48859);
or UO_1809 (O_1809,N_47854,N_46590);
nor UO_1810 (O_1810,N_45563,N_43618);
or UO_1811 (O_1811,N_44402,N_45259);
nand UO_1812 (O_1812,N_44109,N_45683);
nor UO_1813 (O_1813,N_46827,N_43179);
and UO_1814 (O_1814,N_44787,N_42150);
nor UO_1815 (O_1815,N_45027,N_41820);
nand UO_1816 (O_1816,N_47264,N_45048);
xor UO_1817 (O_1817,N_44075,N_44116);
nor UO_1818 (O_1818,N_42278,N_44205);
nor UO_1819 (O_1819,N_40714,N_44791);
and UO_1820 (O_1820,N_49054,N_43425);
nor UO_1821 (O_1821,N_42935,N_43783);
xnor UO_1822 (O_1822,N_42183,N_41787);
nand UO_1823 (O_1823,N_46959,N_47703);
and UO_1824 (O_1824,N_44908,N_48490);
and UO_1825 (O_1825,N_46420,N_49185);
nand UO_1826 (O_1826,N_44681,N_41805);
or UO_1827 (O_1827,N_43622,N_44546);
or UO_1828 (O_1828,N_42198,N_40644);
nand UO_1829 (O_1829,N_43248,N_46981);
nor UO_1830 (O_1830,N_40695,N_47051);
nand UO_1831 (O_1831,N_46711,N_45996);
or UO_1832 (O_1832,N_42723,N_48305);
and UO_1833 (O_1833,N_47144,N_40241);
and UO_1834 (O_1834,N_48870,N_46602);
nor UO_1835 (O_1835,N_42688,N_40237);
and UO_1836 (O_1836,N_45760,N_45585);
and UO_1837 (O_1837,N_42251,N_49973);
xor UO_1838 (O_1838,N_43154,N_43008);
and UO_1839 (O_1839,N_43404,N_48311);
and UO_1840 (O_1840,N_45154,N_46275);
xnor UO_1841 (O_1841,N_49129,N_44072);
nor UO_1842 (O_1842,N_46863,N_46338);
xor UO_1843 (O_1843,N_47714,N_43727);
nand UO_1844 (O_1844,N_47198,N_42220);
and UO_1845 (O_1845,N_48831,N_47448);
nor UO_1846 (O_1846,N_43627,N_48228);
or UO_1847 (O_1847,N_47571,N_49645);
nand UO_1848 (O_1848,N_47951,N_45338);
nand UO_1849 (O_1849,N_40338,N_42703);
or UO_1850 (O_1850,N_41899,N_43599);
and UO_1851 (O_1851,N_42062,N_49647);
xor UO_1852 (O_1852,N_45193,N_40779);
and UO_1853 (O_1853,N_45707,N_44442);
xnor UO_1854 (O_1854,N_49390,N_48205);
or UO_1855 (O_1855,N_47241,N_41003);
nor UO_1856 (O_1856,N_45429,N_49335);
xnor UO_1857 (O_1857,N_42127,N_46249);
or UO_1858 (O_1858,N_41479,N_40595);
nor UO_1859 (O_1859,N_43257,N_47663);
nand UO_1860 (O_1860,N_40982,N_48905);
xor UO_1861 (O_1861,N_42910,N_42600);
or UO_1862 (O_1862,N_40788,N_46724);
xor UO_1863 (O_1863,N_42759,N_44735);
or UO_1864 (O_1864,N_45597,N_42397);
or UO_1865 (O_1865,N_41221,N_43217);
nor UO_1866 (O_1866,N_44270,N_40007);
nand UO_1867 (O_1867,N_44741,N_47333);
or UO_1868 (O_1868,N_42145,N_49850);
nor UO_1869 (O_1869,N_41367,N_43307);
nor UO_1870 (O_1870,N_46299,N_49839);
or UO_1871 (O_1871,N_49256,N_41394);
nand UO_1872 (O_1872,N_42486,N_47537);
xor UO_1873 (O_1873,N_41645,N_40358);
xor UO_1874 (O_1874,N_46877,N_44376);
xnor UO_1875 (O_1875,N_47579,N_42172);
xnor UO_1876 (O_1876,N_40902,N_40985);
and UO_1877 (O_1877,N_44960,N_45022);
xor UO_1878 (O_1878,N_46698,N_48611);
or UO_1879 (O_1879,N_40210,N_40578);
nor UO_1880 (O_1880,N_44777,N_47280);
nor UO_1881 (O_1881,N_46032,N_44592);
and UO_1882 (O_1882,N_45140,N_49771);
and UO_1883 (O_1883,N_47383,N_49882);
or UO_1884 (O_1884,N_43002,N_44157);
or UO_1885 (O_1885,N_46121,N_43061);
nand UO_1886 (O_1886,N_49695,N_45274);
xor UO_1887 (O_1887,N_41817,N_40089);
nor UO_1888 (O_1888,N_44812,N_40806);
nand UO_1889 (O_1889,N_48420,N_48815);
and UO_1890 (O_1890,N_46709,N_48786);
nand UO_1891 (O_1891,N_48659,N_45496);
nand UO_1892 (O_1892,N_45794,N_41933);
or UO_1893 (O_1893,N_45859,N_46671);
and UO_1894 (O_1894,N_41487,N_44490);
xor UO_1895 (O_1895,N_49119,N_40870);
or UO_1896 (O_1896,N_41348,N_46062);
xnor UO_1897 (O_1897,N_46649,N_47484);
nand UO_1898 (O_1898,N_49457,N_46889);
and UO_1899 (O_1899,N_48598,N_41573);
xor UO_1900 (O_1900,N_43815,N_40112);
nor UO_1901 (O_1901,N_45587,N_41038);
and UO_1902 (O_1902,N_41030,N_43046);
nand UO_1903 (O_1903,N_48149,N_49364);
and UO_1904 (O_1904,N_46832,N_40765);
and UO_1905 (O_1905,N_46238,N_44949);
and UO_1906 (O_1906,N_48002,N_46052);
nand UO_1907 (O_1907,N_48450,N_45941);
xnor UO_1908 (O_1908,N_40936,N_40552);
xnor UO_1909 (O_1909,N_45126,N_46180);
or UO_1910 (O_1910,N_42643,N_41186);
nor UO_1911 (O_1911,N_44309,N_42655);
nand UO_1912 (O_1912,N_45591,N_46395);
and UO_1913 (O_1913,N_40420,N_41536);
or UO_1914 (O_1914,N_46770,N_46019);
nand UO_1915 (O_1915,N_43170,N_47785);
nand UO_1916 (O_1916,N_46597,N_42728);
or UO_1917 (O_1917,N_43205,N_48643);
xnor UO_1918 (O_1918,N_41932,N_40921);
nand UO_1919 (O_1919,N_48452,N_45391);
nor UO_1920 (O_1920,N_49274,N_46402);
xnor UO_1921 (O_1921,N_44739,N_49019);
nand UO_1922 (O_1922,N_45748,N_42037);
or UO_1923 (O_1923,N_45482,N_45881);
or UO_1924 (O_1924,N_45565,N_44085);
nor UO_1925 (O_1925,N_46678,N_49497);
or UO_1926 (O_1926,N_44560,N_40906);
xor UO_1927 (O_1927,N_48332,N_43095);
nand UO_1928 (O_1928,N_41938,N_43680);
and UO_1929 (O_1929,N_48238,N_47745);
nor UO_1930 (O_1930,N_47090,N_40027);
nand UO_1931 (O_1931,N_49892,N_43632);
nor UO_1932 (O_1932,N_43381,N_49827);
nand UO_1933 (O_1933,N_46628,N_43640);
nand UO_1934 (O_1934,N_48913,N_49807);
or UO_1935 (O_1935,N_46589,N_45105);
nand UO_1936 (O_1936,N_44062,N_48187);
nor UO_1937 (O_1937,N_44982,N_40900);
nand UO_1938 (O_1938,N_45960,N_42208);
nand UO_1939 (O_1939,N_49846,N_49438);
nor UO_1940 (O_1940,N_48151,N_44469);
xor UO_1941 (O_1941,N_43216,N_49778);
nand UO_1942 (O_1942,N_42668,N_47049);
nor UO_1943 (O_1943,N_44728,N_44154);
and UO_1944 (O_1944,N_42473,N_48510);
nor UO_1945 (O_1945,N_48858,N_49726);
nor UO_1946 (O_1946,N_45414,N_47968);
nand UO_1947 (O_1947,N_43024,N_48926);
nor UO_1948 (O_1948,N_49381,N_43625);
or UO_1949 (O_1949,N_43818,N_48527);
xnor UO_1950 (O_1950,N_42285,N_44287);
nand UO_1951 (O_1951,N_41593,N_46985);
xnor UO_1952 (O_1952,N_41859,N_42878);
nand UO_1953 (O_1953,N_48419,N_40041);
xnor UO_1954 (O_1954,N_49829,N_49762);
nor UO_1955 (O_1955,N_48628,N_45926);
nand UO_1956 (O_1956,N_49001,N_40350);
xnor UO_1957 (O_1957,N_46940,N_43932);
and UO_1958 (O_1958,N_41168,N_48603);
and UO_1959 (O_1959,N_43482,N_44890);
or UO_1960 (O_1960,N_44145,N_40250);
xor UO_1961 (O_1961,N_48845,N_41009);
and UO_1962 (O_1962,N_49761,N_44035);
xnor UO_1963 (O_1963,N_46212,N_45646);
and UO_1964 (O_1964,N_45340,N_41988);
xor UO_1965 (O_1965,N_48216,N_43303);
or UO_1966 (O_1966,N_47218,N_42999);
nand UO_1967 (O_1967,N_42021,N_47661);
nor UO_1968 (O_1968,N_47655,N_44259);
nand UO_1969 (O_1969,N_41075,N_44477);
nor UO_1970 (O_1970,N_42053,N_48403);
and UO_1971 (O_1971,N_40292,N_42901);
or UO_1972 (O_1972,N_47173,N_41337);
xor UO_1973 (O_1973,N_47708,N_42293);
and UO_1974 (O_1974,N_49203,N_42738);
nand UO_1975 (O_1975,N_48163,N_49417);
nand UO_1976 (O_1976,N_45802,N_47318);
nand UO_1977 (O_1977,N_44020,N_45670);
nand UO_1978 (O_1978,N_40690,N_46405);
xor UO_1979 (O_1979,N_45513,N_41060);
and UO_1980 (O_1980,N_43559,N_41151);
or UO_1981 (O_1981,N_41936,N_49580);
nor UO_1982 (O_1982,N_43412,N_41918);
and UO_1983 (O_1983,N_43260,N_40231);
and UO_1984 (O_1984,N_47480,N_47205);
nor UO_1985 (O_1985,N_49261,N_47742);
nand UO_1986 (O_1986,N_47254,N_48879);
nand UO_1987 (O_1987,N_46993,N_41291);
and UO_1988 (O_1988,N_45867,N_42639);
and UO_1989 (O_1989,N_44965,N_44650);
nand UO_1990 (O_1990,N_44362,N_47922);
xnor UO_1991 (O_1991,N_43883,N_44481);
nand UO_1992 (O_1992,N_49107,N_41725);
xor UO_1993 (O_1993,N_45376,N_42661);
xnor UO_1994 (O_1994,N_48388,N_48763);
or UO_1995 (O_1995,N_48043,N_43038);
xnor UO_1996 (O_1996,N_49808,N_49954);
nand UO_1997 (O_1997,N_43004,N_45791);
nor UO_1998 (O_1998,N_40774,N_47977);
nand UO_1999 (O_1999,N_49259,N_43376);
or UO_2000 (O_2000,N_45028,N_49329);
and UO_2001 (O_2001,N_46126,N_49605);
and UO_2002 (O_2002,N_42742,N_42853);
xor UO_2003 (O_2003,N_49687,N_43853);
and UO_2004 (O_2004,N_43539,N_46476);
nor UO_2005 (O_2005,N_46972,N_43290);
nand UO_2006 (O_2006,N_46176,N_41924);
nand UO_2007 (O_2007,N_45547,N_40489);
xnor UO_2008 (O_2008,N_46310,N_48386);
and UO_2009 (O_2009,N_44872,N_49545);
xnor UO_2010 (O_2010,N_44925,N_48974);
nand UO_2011 (O_2011,N_47208,N_43532);
nand UO_2012 (O_2012,N_44090,N_47083);
or UO_2013 (O_2013,N_40204,N_44621);
nand UO_2014 (O_2014,N_42753,N_43166);
or UO_2015 (O_2015,N_43866,N_42309);
or UO_2016 (O_2016,N_46284,N_45962);
xnor UO_2017 (O_2017,N_41578,N_40448);
or UO_2018 (O_2018,N_45084,N_47292);
xor UO_2019 (O_2019,N_45965,N_40137);
nor UO_2020 (O_2020,N_48407,N_47850);
nand UO_2021 (O_2021,N_48112,N_42364);
and UO_2022 (O_2022,N_43085,N_42755);
nor UO_2023 (O_2023,N_43995,N_41677);
xnor UO_2024 (O_2024,N_45725,N_49706);
nand UO_2025 (O_2025,N_42577,N_48811);
or UO_2026 (O_2026,N_48961,N_42455);
nor UO_2027 (O_2027,N_42535,N_46505);
nor UO_2028 (O_2028,N_46817,N_45454);
xnor UO_2029 (O_2029,N_46295,N_48373);
xnor UO_2030 (O_2030,N_42071,N_45007);
xnor UO_2031 (O_2031,N_40867,N_47639);
or UO_2032 (O_2032,N_49554,N_45575);
and UO_2033 (O_2033,N_43550,N_42182);
and UO_2034 (O_2034,N_43912,N_48710);
and UO_2035 (O_2035,N_42973,N_45548);
or UO_2036 (O_2036,N_46263,N_45322);
nor UO_2037 (O_2037,N_46093,N_42227);
xor UO_2038 (O_2038,N_44234,N_41551);
xor UO_2039 (O_2039,N_49705,N_41420);
or UO_2040 (O_2040,N_41327,N_47827);
or UO_2041 (O_2041,N_46172,N_45762);
and UO_2042 (O_2042,N_41943,N_45468);
and UO_2043 (O_2043,N_43493,N_41258);
nand UO_2044 (O_2044,N_41948,N_40526);
xnor UO_2045 (O_2045,N_43375,N_49320);
or UO_2046 (O_2046,N_42517,N_45641);
nor UO_2047 (O_2047,N_42678,N_47549);
nand UO_2048 (O_2048,N_40014,N_40820);
and UO_2049 (O_2049,N_47188,N_45991);
nor UO_2050 (O_2050,N_40565,N_41667);
nand UO_2051 (O_2051,N_44399,N_44824);
nor UO_2052 (O_2052,N_45175,N_45907);
xor UO_2053 (O_2053,N_40811,N_43424);
nand UO_2054 (O_2054,N_44497,N_42046);
nor UO_2055 (O_2055,N_40326,N_45671);
nand UO_2056 (O_2056,N_48501,N_40465);
nor UO_2057 (O_2057,N_42149,N_43555);
and UO_2058 (O_2058,N_46496,N_42798);
xor UO_2059 (O_2059,N_43241,N_40557);
or UO_2060 (O_2060,N_45448,N_42503);
and UO_2061 (O_2061,N_43795,N_43728);
nor UO_2062 (O_2062,N_41312,N_47615);
and UO_2063 (O_2063,N_47669,N_43207);
nand UO_2064 (O_2064,N_44494,N_40620);
and UO_2065 (O_2065,N_46659,N_46582);
nor UO_2066 (O_2066,N_46451,N_48825);
xnor UO_2067 (O_2067,N_43557,N_48679);
xor UO_2068 (O_2068,N_41991,N_46010);
and UO_2069 (O_2069,N_41717,N_42530);
and UO_2070 (O_2070,N_47953,N_46763);
or UO_2071 (O_2071,N_47815,N_46335);
xnor UO_2072 (O_2072,N_45058,N_46581);
xor UO_2073 (O_2073,N_43238,N_41249);
or UO_2074 (O_2074,N_44045,N_42064);
and UO_2075 (O_2075,N_45008,N_40495);
nand UO_2076 (O_2076,N_40596,N_45037);
or UO_2077 (O_2077,N_41039,N_47801);
and UO_2078 (O_2078,N_46139,N_48271);
nand UO_2079 (O_2079,N_44931,N_46138);
xor UO_2080 (O_2080,N_41887,N_47102);
and UO_2081 (O_2081,N_41769,N_48368);
or UO_2082 (O_2082,N_40729,N_47881);
nor UO_2083 (O_2083,N_48911,N_42199);
nand UO_2084 (O_2084,N_49049,N_45642);
nor UO_2085 (O_2085,N_48258,N_49220);
nand UO_2086 (O_2086,N_47392,N_41165);
nand UO_2087 (O_2087,N_43697,N_47063);
xnor UO_2088 (O_2088,N_40679,N_43915);
nand UO_2089 (O_2089,N_41427,N_48464);
nor UO_2090 (O_2090,N_42408,N_40930);
nand UO_2091 (O_2091,N_45234,N_45600);
xor UO_2092 (O_2092,N_46385,N_45400);
and UO_2093 (O_2093,N_49011,N_43280);
and UO_2094 (O_2094,N_40698,N_48613);
nor UO_2095 (O_2095,N_40681,N_49852);
nand UO_2096 (O_2096,N_41706,N_42581);
and UO_2097 (O_2097,N_48411,N_42856);
nor UO_2098 (O_2098,N_46518,N_45701);
xor UO_2099 (O_2099,N_48150,N_46282);
or UO_2100 (O_2100,N_47330,N_46700);
or UO_2101 (O_2101,N_44528,N_41299);
or UO_2102 (O_2102,N_40629,N_41500);
or UO_2103 (O_2103,N_46303,N_47342);
nor UO_2104 (O_2104,N_49095,N_49777);
xnor UO_2105 (O_2105,N_42377,N_48387);
and UO_2106 (O_2106,N_46886,N_45783);
or UO_2107 (O_2107,N_44846,N_41145);
nand UO_2108 (O_2108,N_42463,N_49081);
or UO_2109 (O_2109,N_44678,N_47731);
and UO_2110 (O_2110,N_45763,N_42052);
nand UO_2111 (O_2111,N_45590,N_45290);
nand UO_2112 (O_2112,N_41260,N_44512);
or UO_2113 (O_2113,N_44674,N_49281);
nor UO_2114 (O_2114,N_46970,N_41150);
and UO_2115 (O_2115,N_42642,N_47348);
nor UO_2116 (O_2116,N_45382,N_41568);
xor UO_2117 (O_2117,N_48394,N_46714);
nand UO_2118 (O_2118,N_41171,N_43964);
nor UO_2119 (O_2119,N_42230,N_43872);
and UO_2120 (O_2120,N_41961,N_45264);
or UO_2121 (O_2121,N_43088,N_45014);
and UO_2122 (O_2122,N_47103,N_46539);
nor UO_2123 (O_2123,N_46888,N_40661);
and UO_2124 (O_2124,N_49518,N_49104);
xor UO_2125 (O_2125,N_44257,N_48822);
or UO_2126 (O_2126,N_47900,N_42972);
nand UO_2127 (O_2127,N_42633,N_45917);
nor UO_2128 (O_2128,N_40183,N_43516);
nand UO_2129 (O_2129,N_48769,N_48306);
nand UO_2130 (O_2130,N_49790,N_43988);
nand UO_2131 (O_2131,N_49287,N_41460);
xnor UO_2132 (O_2132,N_44942,N_43379);
or UO_2133 (O_2133,N_47517,N_44055);
or UO_2134 (O_2134,N_49474,N_48255);
nand UO_2135 (O_2135,N_42112,N_49393);
or UO_2136 (O_2136,N_47401,N_41564);
xnor UO_2137 (O_2137,N_43506,N_42582);
xnor UO_2138 (O_2138,N_41471,N_47434);
or UO_2139 (O_2139,N_40400,N_46246);
nand UO_2140 (O_2140,N_47117,N_49847);
and UO_2141 (O_2141,N_44004,N_41319);
nor UO_2142 (O_2142,N_41699,N_46715);
nand UO_2143 (O_2143,N_42739,N_45816);
or UO_2144 (O_2144,N_40298,N_41205);
nor UO_2145 (O_2145,N_46147,N_47142);
xnor UO_2146 (O_2146,N_45480,N_49619);
xnor UO_2147 (O_2147,N_41199,N_41807);
nor UO_2148 (O_2148,N_40966,N_49174);
or UO_2149 (O_2149,N_47976,N_40070);
nor UO_2150 (O_2150,N_41054,N_42405);
xor UO_2151 (O_2151,N_48481,N_47031);
nand UO_2152 (O_2152,N_44576,N_42490);
xor UO_2153 (O_2153,N_46364,N_46300);
nand UO_2154 (O_2154,N_41399,N_48673);
nor UO_2155 (O_2155,N_40615,N_41837);
nor UO_2156 (O_2156,N_40461,N_44386);
and UO_2157 (O_2157,N_41166,N_42379);
nand UO_2158 (O_2158,N_40169,N_44944);
xor UO_2159 (O_2159,N_44932,N_44340);
or UO_2160 (O_2160,N_42882,N_49596);
xnor UO_2161 (O_2161,N_41702,N_41193);
or UO_2162 (O_2162,N_41484,N_42005);
nand UO_2163 (O_2163,N_44565,N_46578);
xnor UO_2164 (O_2164,N_41983,N_43377);
or UO_2165 (O_2165,N_43001,N_47201);
xor UO_2166 (O_2166,N_47744,N_46830);
xnor UO_2167 (O_2167,N_48924,N_41326);
xor UO_2168 (O_2168,N_48378,N_44530);
and UO_2169 (O_2169,N_40435,N_46329);
and UO_2170 (O_2170,N_49128,N_45561);
or UO_2171 (O_2171,N_49784,N_42677);
nor UO_2172 (O_2172,N_40786,N_43345);
nor UO_2173 (O_2173,N_48409,N_45631);
xor UO_2174 (O_2174,N_41930,N_45675);
nand UO_2175 (O_2175,N_41028,N_46241);
nor UO_2176 (O_2176,N_48489,N_45530);
and UO_2177 (O_2177,N_43273,N_44795);
nand UO_2178 (O_2178,N_45302,N_47586);
and UO_2179 (O_2179,N_47361,N_40664);
nand UO_2180 (O_2180,N_43672,N_41272);
nor UO_2181 (O_2181,N_42003,N_42768);
or UO_2182 (O_2182,N_45216,N_48768);
xnor UO_2183 (O_2183,N_49987,N_42740);
nor UO_2184 (O_2184,N_45810,N_46567);
xnor UO_2185 (O_2185,N_49170,N_40636);
and UO_2186 (O_2186,N_47630,N_46415);
and UO_2187 (O_2187,N_40242,N_44694);
xnor UO_2188 (O_2188,N_47138,N_46170);
nor UO_2189 (O_2189,N_49416,N_45043);
xor UO_2190 (O_2190,N_46555,N_48875);
and UO_2191 (O_2191,N_44406,N_43177);
nor UO_2192 (O_2192,N_43946,N_43676);
nand UO_2193 (O_2193,N_40519,N_46919);
nor UO_2194 (O_2194,N_43228,N_49121);
and UO_2195 (O_2195,N_47075,N_46548);
and UO_2196 (O_2196,N_48965,N_41846);
and UO_2197 (O_2197,N_49606,N_46457);
or UO_2198 (O_2198,N_49184,N_45301);
nor UO_2199 (O_2199,N_44536,N_43534);
and UO_2200 (O_2200,N_42674,N_48507);
nand UO_2201 (O_2201,N_46912,N_41096);
nor UO_2202 (O_2202,N_47287,N_47023);
nand UO_2203 (O_2203,N_44554,N_46189);
xnor UO_2204 (O_2204,N_41363,N_43131);
nand UO_2205 (O_2205,N_48827,N_42152);
nand UO_2206 (O_2206,N_44506,N_48461);
and UO_2207 (O_2207,N_46231,N_46230);
and UO_2208 (O_2208,N_48756,N_46696);
nand UO_2209 (O_2209,N_40710,N_48415);
nor UO_2210 (O_2210,N_45977,N_40876);
and UO_2211 (O_2211,N_45601,N_44865);
xnor UO_2212 (O_2212,N_41441,N_41704);
xor UO_2213 (O_2213,N_40592,N_47425);
nand UO_2214 (O_2214,N_41848,N_40513);
nand UO_2215 (O_2215,N_42349,N_49027);
xor UO_2216 (O_2216,N_41922,N_40052);
and UO_2217 (O_2217,N_49608,N_49087);
or UO_2218 (O_2218,N_40401,N_44347);
nand UO_2219 (O_2219,N_44903,N_49682);
or UO_2220 (O_2220,N_48562,N_49737);
xor UO_2221 (O_2221,N_48496,N_43359);
and UO_2222 (O_2222,N_46611,N_44167);
nand UO_2223 (O_2223,N_48792,N_41012);
or UO_2224 (O_2224,N_41795,N_49942);
xor UO_2225 (O_2225,N_47493,N_43311);
or UO_2226 (O_2226,N_47358,N_41341);
and UO_2227 (O_2227,N_44834,N_46819);
nor UO_2228 (O_2228,N_42023,N_49249);
nor UO_2229 (O_2229,N_40720,N_48119);
nor UO_2230 (O_2230,N_42505,N_43884);
and UO_2231 (O_2231,N_46320,N_48010);
nand UO_2232 (O_2232,N_43961,N_44286);
and UO_2233 (O_2233,N_42030,N_44151);
xnor UO_2234 (O_2234,N_41721,N_41532);
and UO_2235 (O_2235,N_42243,N_41104);
and UO_2236 (O_2236,N_46991,N_41872);
xnor UO_2237 (O_2237,N_48990,N_47438);
xnor UO_2238 (O_2238,N_42715,N_48703);
and UO_2239 (O_2239,N_41888,N_45994);
nand UO_2240 (O_2240,N_44711,N_46695);
xor UO_2241 (O_2241,N_47303,N_42193);
or UO_2242 (O_2242,N_42951,N_45408);
nor UO_2243 (O_2243,N_46018,N_48323);
or UO_2244 (O_2244,N_40125,N_42968);
nand UO_2245 (O_2245,N_47428,N_49451);
or UO_2246 (O_2246,N_44736,N_48720);
or UO_2247 (O_2247,N_42301,N_40939);
or UO_2248 (O_2248,N_43123,N_48120);
or UO_2249 (O_2249,N_43773,N_46544);
nand UO_2250 (O_2250,N_48851,N_40107);
nand UO_2251 (O_2251,N_48537,N_48764);
nand UO_2252 (O_2252,N_48778,N_48887);
or UO_2253 (O_2253,N_42061,N_45593);
and UO_2254 (O_2254,N_48430,N_46849);
xor UO_2255 (O_2255,N_43330,N_45499);
xnor UO_2256 (O_2256,N_42284,N_47636);
and UO_2257 (O_2257,N_45134,N_49956);
or UO_2258 (O_2258,N_44969,N_47518);
and UO_2259 (O_2259,N_40588,N_48937);
nor UO_2260 (O_2260,N_44353,N_48060);
nor UO_2261 (O_2261,N_48381,N_42206);
xor UO_2262 (O_2262,N_44419,N_41694);
or UO_2263 (O_2263,N_41597,N_48517);
nor UO_2264 (O_2264,N_48617,N_40705);
or UO_2265 (O_2265,N_43188,N_41562);
xnor UO_2266 (O_2266,N_47071,N_49751);
xnor UO_2267 (O_2267,N_41967,N_46604);
and UO_2268 (O_2268,N_42998,N_44721);
xor UO_2269 (O_2269,N_42623,N_46938);
and UO_2270 (O_2270,N_48096,N_49577);
nor UO_2271 (O_2271,N_43107,N_45909);
or UO_2272 (O_2272,N_41228,N_46566);
or UO_2273 (O_2273,N_40597,N_45713);
xor UO_2274 (O_2274,N_42016,N_47125);
and UO_2275 (O_2275,N_48876,N_49456);
or UO_2276 (O_2276,N_49838,N_42429);
nand UO_2277 (O_2277,N_42561,N_40180);
and UO_2278 (O_2278,N_45325,N_47088);
nand UO_2279 (O_2279,N_49114,N_42931);
xnor UO_2280 (O_2280,N_49556,N_40586);
nand UO_2281 (O_2281,N_48453,N_43322);
and UO_2282 (O_2282,N_44509,N_46971);
xnor UO_2283 (O_2283,N_46795,N_46446);
and UO_2284 (O_2284,N_42754,N_48623);
nand UO_2285 (O_2285,N_48735,N_49387);
xnor UO_2286 (O_2286,N_48148,N_42255);
nand UO_2287 (O_2287,N_40173,N_43010);
xor UO_2288 (O_2288,N_45214,N_44752);
xor UO_2289 (O_2289,N_44913,N_48179);
nand UO_2290 (O_2290,N_45724,N_46631);
and UO_2291 (O_2291,N_46722,N_45968);
nand UO_2292 (O_2292,N_49718,N_44672);
or UO_2293 (O_2293,N_42264,N_43603);
or UO_2294 (O_2294,N_45495,N_40423);
and UO_2295 (O_2295,N_49976,N_49780);
or UO_2296 (O_2296,N_41303,N_41582);
nor UO_2297 (O_2297,N_42506,N_47403);
and UO_2298 (O_2298,N_42049,N_47675);
nand UO_2299 (O_2299,N_41379,N_43399);
nand UO_2300 (O_2300,N_45252,N_49513);
nor UO_2301 (O_2301,N_49837,N_42744);
nor UO_2302 (O_2302,N_44688,N_45692);
or UO_2303 (O_2303,N_43070,N_42170);
or UO_2304 (O_2304,N_46842,N_40163);
or UO_2305 (O_2305,N_46051,N_44410);
and UO_2306 (O_2306,N_43371,N_40392);
and UO_2307 (O_2307,N_45491,N_46173);
and UO_2308 (O_2308,N_47936,N_44935);
xnor UO_2309 (O_2309,N_45015,N_49634);
or UO_2310 (O_2310,N_47824,N_40914);
xor UO_2311 (O_2311,N_45820,N_44017);
nand UO_2312 (O_2312,N_41659,N_46721);
nor UO_2313 (O_2313,N_41170,N_47207);
and UO_2314 (O_2314,N_48515,N_46224);
xor UO_2315 (O_2315,N_43965,N_46236);
and UO_2316 (O_2316,N_46788,N_46732);
nor UO_2317 (O_2317,N_45893,N_41996);
or UO_2318 (O_2318,N_44808,N_44166);
and UO_2319 (O_2319,N_44284,N_44575);
xnor UO_2320 (O_2320,N_49842,N_46069);
and UO_2321 (O_2321,N_44768,N_44863);
or UO_2322 (O_2322,N_46225,N_40795);
or UO_2323 (O_2323,N_41439,N_40278);
nand UO_2324 (O_2324,N_43691,N_40373);
and UO_2325 (O_2325,N_46983,N_45285);
and UO_2326 (O_2326,N_48848,N_43774);
xnor UO_2327 (O_2327,N_45847,N_41747);
nor UO_2328 (O_2328,N_40997,N_45691);
and UO_2329 (O_2329,N_47095,N_41295);
nand UO_2330 (O_2330,N_41978,N_49736);
nand UO_2331 (O_2331,N_49272,N_43463);
nand UO_2332 (O_2332,N_42579,N_47649);
or UO_2333 (O_2333,N_45524,N_47648);
nand UO_2334 (O_2334,N_49713,N_46056);
xor UO_2335 (O_2335,N_46363,N_49418);
nand UO_2336 (O_2336,N_46673,N_41498);
nor UO_2337 (O_2337,N_45265,N_43726);
xnor UO_2338 (O_2338,N_43925,N_43974);
or UO_2339 (O_2339,N_46759,N_42362);
and UO_2340 (O_2340,N_42510,N_47113);
xnor UO_2341 (O_2341,N_45650,N_41742);
nor UO_2342 (O_2342,N_49216,N_46821);
nor UO_2343 (O_2343,N_41671,N_44322);
or UO_2344 (O_2344,N_43529,N_45967);
and UO_2345 (O_2345,N_44724,N_43781);
nor UO_2346 (O_2346,N_48124,N_41476);
and UO_2347 (O_2347,N_47506,N_49548);
xnor UO_2348 (O_2348,N_42118,N_42173);
and UO_2349 (O_2349,N_46864,N_48483);
nor UO_2350 (O_2350,N_42997,N_44242);
nand UO_2351 (O_2351,N_49862,N_42751);
nand UO_2352 (O_2352,N_48730,N_46352);
nand UO_2353 (O_2353,N_46475,N_40028);
nand UO_2354 (O_2354,N_43426,N_42100);
xor UO_2355 (O_2355,N_43576,N_47640);
and UO_2356 (O_2356,N_45184,N_46854);
and UO_2357 (O_2357,N_43760,N_47813);
and UO_2358 (O_2358,N_49859,N_47239);
or UO_2359 (O_2359,N_40407,N_42809);
nor UO_2360 (O_2360,N_44984,N_45885);
nor UO_2361 (O_2361,N_42281,N_48097);
nand UO_2362 (O_2362,N_42598,N_44686);
nand UO_2363 (O_2363,N_46818,N_48790);
and UO_2364 (O_2364,N_43786,N_41035);
nor UO_2365 (O_2365,N_44269,N_45073);
and UO_2366 (O_2366,N_49338,N_46592);
nor UO_2367 (O_2367,N_40598,N_48275);
nand UO_2368 (O_2368,N_48322,N_47897);
nor UO_2369 (O_2369,N_40251,N_46199);
nor UO_2370 (O_2370,N_46484,N_44338);
and UO_2371 (O_2371,N_44482,N_49789);
nor UO_2372 (O_2372,N_43396,N_45768);
or UO_2373 (O_2373,N_45337,N_43895);
nor UO_2374 (O_2374,N_40953,N_49587);
nor UO_2375 (O_2375,N_40383,N_41683);
xor UO_2376 (O_2376,N_45643,N_41192);
nand UO_2377 (O_2377,N_40517,N_40020);
and UO_2378 (O_2378,N_40706,N_41855);
xor UO_2379 (O_2379,N_40318,N_49351);
or UO_2380 (O_2380,N_48454,N_40229);
or UO_2381 (O_2381,N_46908,N_43413);
or UO_2382 (O_2382,N_49872,N_46586);
and UO_2383 (O_2383,N_40343,N_42067);
nand UO_2384 (O_2384,N_47043,N_42862);
or UO_2385 (O_2385,N_48689,N_44299);
or UO_2386 (O_2386,N_44770,N_40943);
nand UO_2387 (O_2387,N_46927,N_44733);
nand UO_2388 (O_2388,N_44178,N_48807);
nand UO_2389 (O_2389,N_44354,N_44424);
nand UO_2390 (O_2390,N_40676,N_45097);
or UO_2391 (O_2391,N_48355,N_46963);
and UO_2392 (O_2392,N_44878,N_44318);
or UO_2393 (O_2393,N_43717,N_48530);
or UO_2394 (O_2394,N_47876,N_43434);
xnor UO_2395 (O_2395,N_40845,N_47570);
nand UO_2396 (O_2396,N_45981,N_49752);
nor UO_2397 (O_2397,N_45498,N_45424);
nor UO_2398 (O_2398,N_47786,N_49493);
nor UO_2399 (O_2399,N_43176,N_46899);
xor UO_2400 (O_2400,N_48350,N_47947);
nand UO_2401 (O_2401,N_41827,N_42412);
and UO_2402 (O_2402,N_41267,N_47541);
nand UO_2403 (O_2403,N_44331,N_41274);
xnor UO_2404 (O_2404,N_47741,N_42533);
and UO_2405 (O_2405,N_45233,N_42481);
nor UO_2406 (O_2406,N_46187,N_42670);
xnor UO_2407 (O_2407,N_46333,N_45908);
or UO_2408 (O_2408,N_41207,N_41423);
xnor UO_2409 (O_2409,N_43668,N_49604);
or UO_2410 (O_2410,N_42804,N_47307);
nor UO_2411 (O_2411,N_44927,N_49830);
and UO_2412 (O_2412,N_41574,N_45572);
xnor UO_2413 (O_2413,N_40669,N_40978);
and UO_2414 (O_2414,N_49168,N_48265);
nor UO_2415 (O_2415,N_43250,N_40347);
or UO_2416 (O_2416,N_40055,N_43721);
nand UO_2417 (O_2417,N_41089,N_40315);
or UO_2418 (O_2418,N_48840,N_41048);
nor UO_2419 (O_2419,N_41451,N_40266);
nand UO_2420 (O_2420,N_46090,N_46713);
nand UO_2421 (O_2421,N_43704,N_40006);
or UO_2422 (O_2422,N_40922,N_46196);
xnor UO_2423 (O_2423,N_42586,N_47524);
xnor UO_2424 (O_2424,N_43967,N_44773);
nand UO_2425 (O_2425,N_45492,N_47415);
and UO_2426 (O_2426,N_42386,N_40284);
nand UO_2427 (O_2427,N_45352,N_42253);
or UO_2428 (O_2428,N_48923,N_40660);
or UO_2429 (O_2429,N_45668,N_40605);
xnor UO_2430 (O_2430,N_49091,N_49917);
nand UO_2431 (O_2431,N_49328,N_40024);
and UO_2432 (O_2432,N_46924,N_44543);
nor UO_2433 (O_2433,N_40983,N_41382);
nand UO_2434 (O_2434,N_46382,N_44978);
nor UO_2435 (O_2435,N_44320,N_46653);
nand UO_2436 (O_2436,N_42872,N_47046);
nand UO_2437 (O_2437,N_42690,N_49860);
nand UO_2438 (O_2438,N_42102,N_46152);
or UO_2439 (O_2439,N_46570,N_44461);
nand UO_2440 (O_2440,N_45576,N_47690);
or UO_2441 (O_2441,N_47993,N_47369);
and UO_2442 (O_2442,N_41508,N_40451);
xor UO_2443 (O_2443,N_46909,N_48982);
nand UO_2444 (O_2444,N_49624,N_40263);
and UO_2445 (O_2445,N_45033,N_47155);
xnor UO_2446 (O_2446,N_48303,N_48486);
or UO_2447 (O_2447,N_49124,N_40951);
nand UO_2448 (O_2448,N_46929,N_46438);
xor UO_2449 (O_2449,N_45049,N_44894);
and UO_2450 (O_2450,N_46058,N_40724);
and UO_2451 (O_2451,N_46378,N_46442);
nor UO_2452 (O_2452,N_46699,N_48196);
and UO_2453 (O_2453,N_47126,N_45217);
xnor UO_2454 (O_2454,N_44645,N_47455);
or UO_2455 (O_2455,N_43178,N_43226);
nor UO_2456 (O_2456,N_41119,N_44732);
xnor UO_2457 (O_2457,N_40499,N_43419);
nor UO_2458 (O_2458,N_45761,N_49758);
nand UO_2459 (O_2459,N_48663,N_41311);
and UO_2460 (O_2460,N_46455,N_43737);
nor UO_2461 (O_2461,N_49958,N_48907);
nand UO_2462 (O_2462,N_48448,N_40260);
and UO_2463 (O_2463,N_45378,N_40393);
or UO_2464 (O_2464,N_40172,N_45623);
xnor UO_2465 (O_2465,N_43435,N_44407);
nand UO_2466 (O_2466,N_44315,N_44185);
or UO_2467 (O_2467,N_43114,N_49225);
and UO_2468 (O_2468,N_40297,N_44250);
or UO_2469 (O_2469,N_46185,N_45299);
nor UO_2470 (O_2470,N_41774,N_41426);
and UO_2471 (O_2471,N_45362,N_46244);
xnor UO_2472 (O_2472,N_43677,N_42226);
xnor UO_2473 (O_2473,N_44572,N_43903);
xnor UO_2474 (O_2474,N_42886,N_43919);
nand UO_2475 (O_2475,N_47482,N_49539);
or UO_2476 (O_2476,N_43183,N_43996);
or UO_2477 (O_2477,N_45822,N_46175);
and UO_2478 (O_2478,N_45469,N_43283);
xnor UO_2479 (O_2479,N_42169,N_46268);
xnor UO_2480 (O_2480,N_40987,N_45317);
nand UO_2481 (O_2481,N_47124,N_42099);
nor UO_2482 (O_2482,N_45516,N_46771);
and UO_2483 (O_2483,N_46276,N_44142);
xnor UO_2484 (O_2484,N_45336,N_43471);
or UO_2485 (O_2485,N_40549,N_49629);
and UO_2486 (O_2486,N_45539,N_49651);
nor UO_2487 (O_2487,N_42713,N_43033);
nor UO_2488 (O_2488,N_41841,N_48413);
or UO_2489 (O_2489,N_47689,N_44153);
xor UO_2490 (O_2490,N_42389,N_44590);
or UO_2491 (O_2491,N_41607,N_49652);
nor UO_2492 (O_2492,N_48571,N_40576);
xor UO_2493 (O_2493,N_49255,N_49564);
xnor UO_2494 (O_2494,N_44520,N_47269);
nand UO_2495 (O_2495,N_43808,N_42140);
xnor UO_2496 (O_2496,N_42356,N_42088);
or UO_2497 (O_2497,N_41844,N_42770);
or UO_2498 (O_2498,N_47067,N_40289);
or UO_2499 (O_2499,N_41280,N_40804);
nand UO_2500 (O_2500,N_41950,N_49181);
xor UO_2501 (O_2501,N_42427,N_46710);
xor UO_2502 (O_2502,N_45785,N_40370);
and UO_2503 (O_2503,N_41576,N_45284);
or UO_2504 (O_2504,N_46057,N_41910);
xor UO_2505 (O_2505,N_48900,N_42627);
xnor UO_2506 (O_2506,N_43792,N_43274);
or UO_2507 (O_2507,N_42358,N_47181);
xnor UO_2508 (O_2508,N_42553,N_42614);
xor UO_2509 (O_2509,N_42874,N_43057);
and UO_2510 (O_2510,N_43971,N_48565);
and UO_2511 (O_2511,N_40404,N_43302);
nand UO_2512 (O_2512,N_47152,N_41140);
and UO_2513 (O_2513,N_47511,N_45619);
and UO_2514 (O_2514,N_43100,N_48365);
nand UO_2515 (O_2515,N_44957,N_40857);
nand UO_2516 (O_2516,N_40262,N_46915);
nand UO_2517 (O_2517,N_48686,N_42042);
nor UO_2518 (O_2518,N_43157,N_46094);
or UO_2519 (O_2519,N_47767,N_45659);
and UO_2520 (O_2520,N_48709,N_44830);
and UO_2521 (O_2521,N_47137,N_46996);
or UO_2522 (O_2522,N_40468,N_49263);
or UO_2523 (O_2523,N_45182,N_41408);
nor UO_2524 (O_2524,N_44300,N_40067);
nand UO_2525 (O_2525,N_48041,N_42026);
nor UO_2526 (O_2526,N_48606,N_41581);
xnor UO_2527 (O_2527,N_45226,N_42769);
nand UO_2528 (O_2528,N_41990,N_44454);
or UO_2529 (O_2529,N_49670,N_40822);
xor UO_2530 (O_2530,N_44193,N_44114);
and UO_2531 (O_2531,N_47056,N_42388);
nor UO_2532 (O_2532,N_43850,N_42458);
nand UO_2533 (O_2533,N_41615,N_47543);
or UO_2534 (O_2534,N_45208,N_42376);
or UO_2535 (O_2535,N_45915,N_48263);
nand UO_2536 (O_2536,N_43308,N_48360);
nor UO_2537 (O_2537,N_41973,N_46078);
xor UO_2538 (O_2538,N_45438,N_49189);
xnor UO_2539 (O_2539,N_47178,N_46106);
and UO_2540 (O_2540,N_43003,N_40281);
nor UO_2541 (O_2541,N_49084,N_42418);
nand UO_2542 (O_2542,N_46125,N_45925);
nand UO_2543 (O_2543,N_45959,N_47326);
nor UO_2544 (O_2544,N_48032,N_41470);
nor UO_2545 (O_2545,N_42626,N_47453);
nor UO_2546 (O_2546,N_43197,N_49152);
and UO_2547 (O_2547,N_44392,N_43852);
xnor UO_2548 (O_2548,N_46283,N_44291);
or UO_2549 (O_2549,N_42432,N_48996);
or UO_2550 (O_2550,N_48336,N_45862);
nand UO_2551 (O_2551,N_45711,N_40604);
nor UO_2552 (O_2552,N_46017,N_48818);
or UO_2553 (O_2553,N_45939,N_40659);
or UO_2554 (O_2554,N_41261,N_49484);
and UO_2555 (O_2555,N_43678,N_48372);
and UO_2556 (O_2556,N_46251,N_44395);
and UO_2557 (O_2557,N_40727,N_48775);
nor UO_2558 (O_2558,N_49522,N_43264);
or UO_2559 (O_2559,N_40234,N_47803);
nand UO_2560 (O_2560,N_45604,N_41304);
nor UO_2561 (O_2561,N_40908,N_43041);
nor UO_2562 (O_2562,N_41378,N_44440);
xnor UO_2563 (O_2563,N_42075,N_45189);
and UO_2564 (O_2564,N_43488,N_40106);
xor UO_2565 (O_2565,N_45533,N_49007);
or UO_2566 (O_2566,N_47474,N_44203);
nand UO_2567 (O_2567,N_47194,N_45066);
or UO_2568 (O_2568,N_42783,N_48525);
and UO_2569 (O_2569,N_43605,N_45972);
nand UO_2570 (O_2570,N_41018,N_47884);
nor UO_2571 (O_2571,N_45549,N_40515);
xnor UO_2572 (O_2572,N_40794,N_49810);
xor UO_2573 (O_2573,N_43080,N_42435);
nand UO_2574 (O_2574,N_46080,N_40111);
and UO_2575 (O_2575,N_47921,N_48741);
or UO_2576 (O_2576,N_49126,N_49260);
or UO_2577 (O_2577,N_44945,N_47894);
and UO_2578 (O_2578,N_44574,N_46922);
xnor UO_2579 (O_2579,N_49668,N_42438);
or UO_2580 (O_2580,N_43886,N_40431);
xor UO_2581 (O_2581,N_42232,N_47810);
and UO_2582 (O_2582,N_44709,N_46879);
nor UO_2583 (O_2583,N_46166,N_49557);
or UO_2584 (O_2584,N_46174,N_42289);
and UO_2585 (O_2585,N_40568,N_48684);
xnor UO_2586 (O_2586,N_46141,N_43180);
xnor UO_2587 (O_2587,N_45858,N_44985);
nor UO_2588 (O_2588,N_42961,N_40956);
nor UO_2589 (O_2589,N_41347,N_44308);
nand UO_2590 (O_2590,N_48560,N_45380);
xnor UO_2591 (O_2591,N_43991,N_48852);
xnor UO_2592 (O_2592,N_49179,N_48680);
nand UO_2593 (O_2593,N_45412,N_40416);
xor UO_2594 (O_2594,N_48473,N_49302);
nor UO_2595 (O_2595,N_44194,N_42612);
nand UO_2596 (O_2596,N_41585,N_44570);
nor UO_2597 (O_2597,N_45920,N_41815);
and UO_2598 (O_2598,N_47368,N_41163);
and UO_2599 (O_2599,N_41402,N_45930);
nor UO_2600 (O_2600,N_49437,N_42978);
and UO_2601 (O_2601,N_40777,N_49290);
and UO_2602 (O_2602,N_41731,N_40244);
xor UO_2603 (O_2603,N_41210,N_41412);
nand UO_2604 (O_2604,N_45528,N_44603);
or UO_2605 (O_2605,N_43554,N_44261);
nand UO_2606 (O_2606,N_49727,N_44198);
or UO_2607 (O_2607,N_41016,N_47508);
nand UO_2608 (O_2608,N_48776,N_49699);
nor UO_2609 (O_2609,N_40144,N_40403);
xnor UO_2610 (O_2610,N_47617,N_48375);
nand UO_2611 (O_2611,N_47832,N_47577);
nor UO_2612 (O_2612,N_40858,N_42240);
and UO_2613 (O_2613,N_40723,N_44666);
xnor UO_2614 (O_2614,N_40950,N_47580);
and UO_2615 (O_2615,N_42774,N_42699);
xnor UO_2616 (O_2616,N_48934,N_43719);
nor UO_2617 (O_2617,N_43650,N_48000);
or UO_2618 (O_2618,N_47629,N_44339);
xor UO_2619 (O_2619,N_42732,N_48270);
or UO_2620 (O_2620,N_42890,N_46616);
nand UO_2621 (O_2621,N_45389,N_42069);
xnor UO_2622 (O_2622,N_48814,N_45270);
or UO_2623 (O_2623,N_49399,N_46958);
xnor UO_2624 (O_2624,N_47380,N_49063);
xnor UO_2625 (O_2625,N_45494,N_43452);
nand UO_2626 (O_2626,N_49588,N_49066);
xor UO_2627 (O_2627,N_42675,N_41344);
nand UO_2628 (O_2628,N_44989,N_46583);
xnor UO_2629 (O_2629,N_49475,N_45635);
nor UO_2630 (O_2630,N_43428,N_47529);
and UO_2631 (O_2631,N_47779,N_47916);
xnor UO_2632 (O_2632,N_46802,N_45085);
or UO_2633 (O_2633,N_42807,N_43688);
or UO_2634 (O_2634,N_41734,N_41963);
nand UO_2635 (O_2635,N_44704,N_43653);
or UO_2636 (O_2636,N_42008,N_48693);
nor UO_2637 (O_2637,N_45729,N_43510);
nand UO_2638 (O_2638,N_45136,N_46571);
nand UO_2639 (O_2639,N_49583,N_46853);
xor UO_2640 (O_2640,N_43658,N_40139);
nor UO_2641 (O_2641,N_41452,N_42460);
or UO_2642 (O_2642,N_42072,N_49472);
xor UO_2643 (O_2643,N_48269,N_41227);
and UO_2644 (O_2644,N_49349,N_45639);
or UO_2645 (O_2645,N_43059,N_41849);
xor UO_2646 (O_2646,N_41407,N_46502);
nand UO_2647 (O_2647,N_44382,N_42410);
and UO_2648 (O_2648,N_40334,N_49242);
xnor UO_2649 (O_2649,N_40150,N_46717);
or UO_2650 (O_2650,N_41654,N_48539);
nor UO_2651 (O_2651,N_46537,N_48462);
nand UO_2652 (O_2652,N_49675,N_44636);
xor UO_2653 (O_2653,N_47510,N_40713);
and UO_2654 (O_2654,N_42238,N_43150);
nand UO_2655 (O_2655,N_46009,N_42492);
xnor UO_2656 (O_2656,N_42727,N_40034);
nor UO_2657 (O_2657,N_42854,N_46667);
nand UO_2658 (O_2658,N_41857,N_44508);
or UO_2659 (O_2659,N_47602,N_43552);
xnor UO_2660 (O_2660,N_40759,N_44052);
nor UO_2661 (O_2661,N_47678,N_40610);
and UO_2662 (O_2662,N_46065,N_46082);
nand UO_2663 (O_2663,N_47693,N_42002);
or UO_2664 (O_2664,N_47721,N_49957);
xnor UO_2665 (O_2665,N_46401,N_42888);
nand UO_2666 (O_2666,N_42176,N_42562);
and UO_2667 (O_2667,N_45185,N_45956);
nand UO_2668 (O_2668,N_42417,N_48040);
and UO_2669 (O_2669,N_46049,N_44784);
and UO_2670 (O_2670,N_43843,N_43892);
and UO_2671 (O_2671,N_48292,N_43585);
or UO_2672 (O_2672,N_42841,N_46443);
xor UO_2673 (O_2673,N_43867,N_48466);
and UO_2674 (O_2674,N_47014,N_40184);
nor UO_2675 (O_2675,N_49803,N_44918);
and UO_2676 (O_2676,N_46055,N_45282);
or UO_2677 (O_2677,N_45509,N_44947);
nand UO_2678 (O_2678,N_44662,N_48272);
or UO_2679 (O_2679,N_40807,N_46515);
or UO_2680 (O_2680,N_46608,N_47556);
xor UO_2681 (O_2681,N_42578,N_44980);
nor UO_2682 (O_2682,N_47503,N_42887);
and UO_2683 (O_2683,N_47258,N_46769);
xnor UO_2684 (O_2684,N_42585,N_45564);
nand UO_2685 (O_2685,N_46159,N_46366);
nand UO_2686 (O_2686,N_49323,N_48063);
xor UO_2687 (O_2687,N_43906,N_40359);
nand UO_2688 (O_2688,N_43513,N_44420);
nor UO_2689 (O_2689,N_43232,N_46794);
xor UO_2690 (O_2690,N_49023,N_46149);
or UO_2691 (O_2691,N_47019,N_41287);
nand UO_2692 (O_2692,N_45645,N_45574);
xor UO_2693 (O_2693,N_43300,N_40437);
nand UO_2694 (O_2694,N_48441,N_43499);
xor UO_2695 (O_2695,N_45886,N_40016);
xor UO_2696 (O_2696,N_48953,N_42544);
nor UO_2697 (O_2697,N_45098,N_43990);
or UO_2698 (O_2698,N_44283,N_44397);
and UO_2699 (O_2699,N_49963,N_44855);
nand UO_2700 (O_2700,N_45466,N_44996);
xnor UO_2701 (O_2701,N_40496,N_42006);
and UO_2702 (O_2702,N_47216,N_43637);
nor UO_2703 (O_2703,N_47077,N_42752);
nand UO_2704 (O_2704,N_46481,N_49231);
and UO_2705 (O_2705,N_47886,N_46707);
nand UO_2706 (O_2706,N_41401,N_48799);
nor UO_2707 (O_2707,N_42106,N_42719);
and UO_2708 (O_2708,N_43587,N_46950);
nand UO_2709 (O_2709,N_40208,N_49880);
or UO_2710 (O_2710,N_43616,N_43518);
nor UO_2711 (O_2711,N_47523,N_44216);
and UO_2712 (O_2712,N_40314,N_43058);
or UO_2713 (O_2713,N_44191,N_48046);
xor UO_2714 (O_2714,N_41353,N_41788);
nand UO_2715 (O_2715,N_45648,N_47105);
and UO_2716 (O_2716,N_49891,N_45728);
or UO_2717 (O_2717,N_44661,N_47223);
and UO_2718 (O_2718,N_41984,N_41965);
and UO_2719 (O_2719,N_49355,N_47174);
and UO_2720 (O_2720,N_43959,N_46730);
or UO_2721 (O_2721,N_41728,N_44915);
nand UO_2722 (O_2722,N_47391,N_41796);
nor UO_2723 (O_2723,N_40081,N_40832);
and UO_2724 (O_2724,N_48951,N_47954);
and UO_2725 (O_2725,N_40506,N_41733);
nor UO_2726 (O_2726,N_44914,N_40755);
nor UO_2727 (O_2727,N_45316,N_49031);
and UO_2728 (O_2728,N_47909,N_44150);
or UO_2729 (O_2729,N_42322,N_41240);
or UO_2730 (O_2730,N_49948,N_43341);
nor UO_2731 (O_2731,N_43789,N_46252);
xor UO_2732 (O_2732,N_48316,N_46337);
nand UO_2733 (O_2733,N_43251,N_41307);
and UO_2734 (O_2734,N_40143,N_40257);
xor UO_2735 (O_2735,N_42791,N_48935);
nand UO_2736 (O_2736,N_41791,N_47992);
nand UO_2737 (O_2737,N_46939,N_43804);
xor UO_2738 (O_2738,N_45738,N_47797);
and UO_2739 (O_2739,N_45934,N_40999);
nand UO_2740 (O_2740,N_48503,N_40539);
nor UO_2741 (O_2741,N_41406,N_46822);
or UO_2742 (O_2742,N_40165,N_43365);
and UO_2743 (O_2743,N_48458,N_41647);
nand UO_2744 (O_2744,N_43105,N_40527);
xnor UO_2745 (O_2745,N_44551,N_48665);
or UO_2746 (O_2746,N_45179,N_47335);
nor UO_2747 (O_2747,N_48139,N_48225);
nor UO_2748 (O_2748,N_44648,N_40716);
nand UO_2749 (O_2749,N_49365,N_48780);
or UO_2750 (O_2750,N_49212,N_42361);
xnor UO_2751 (O_2751,N_40285,N_48975);
xor UO_2752 (O_2752,N_48122,N_40859);
nor UO_2753 (O_2753,N_47792,N_46213);
and UO_2754 (O_2754,N_41124,N_44391);
and UO_2755 (O_2755,N_46708,N_49360);
nor UO_2756 (O_2756,N_43698,N_46279);
nor UO_2757 (O_2757,N_40621,N_43483);
nand UO_2758 (O_2758,N_40449,N_44218);
nor UO_2759 (O_2759,N_49649,N_40916);
nand UO_2760 (O_2760,N_44516,N_46112);
nor UO_2761 (O_2761,N_40295,N_43328);
nand UO_2762 (O_2762,N_41074,N_47237);
nor UO_2763 (O_2763,N_41776,N_48153);
nand UO_2764 (O_2764,N_40458,N_42066);
nor UO_2765 (O_2765,N_44471,N_40455);
nand UO_2766 (O_2766,N_41997,N_43320);
xnor UO_2767 (O_2767,N_43468,N_47838);
and UO_2768 (O_2768,N_40817,N_45508);
or UO_2769 (O_2769,N_47294,N_49566);
nand UO_2770 (O_2770,N_41099,N_43476);
or UO_2771 (O_2771,N_45205,N_45248);
nand UO_2772 (O_2772,N_45723,N_49972);
or UO_2773 (O_2773,N_49532,N_48600);
and UO_2774 (O_2774,N_44884,N_47616);
and UO_2775 (O_2775,N_48429,N_42313);
or UO_2776 (O_2776,N_47270,N_44231);
and UO_2777 (O_2777,N_46167,N_41288);
xor UO_2778 (O_2778,N_43202,N_43252);
or UO_2779 (O_2779,N_41723,N_46630);
and UO_2780 (O_2780,N_43152,N_43661);
or UO_2781 (O_2781,N_47751,N_49041);
nor UO_2782 (O_2782,N_48333,N_46976);
and UO_2783 (O_2783,N_46737,N_45335);
and UO_2784 (O_2784,N_44067,N_43286);
nor UO_2785 (O_2785,N_48899,N_46688);
and UO_2786 (O_2786,N_47684,N_41323);
or UO_2787 (O_2787,N_47163,N_44445);
or UO_2788 (O_2788,N_48017,N_44141);
nand UO_2789 (O_2789,N_49612,N_44624);
or UO_2790 (O_2790,N_48038,N_45667);
xnor UO_2791 (O_2791,N_45545,N_45244);
or UO_2792 (O_2792,N_47109,N_41676);
nand UO_2793 (O_2793,N_45117,N_48757);
xor UO_2794 (O_2794,N_40640,N_40353);
nand UO_2795 (O_2795,N_47253,N_40197);
nor UO_2796 (O_2796,N_42190,N_46304);
or UO_2797 (O_2797,N_47487,N_44105);
nand UO_2798 (O_2798,N_47251,N_45813);
and UO_2799 (O_2799,N_47956,N_46885);
and UO_2800 (O_2800,N_48635,N_49888);
and UO_2801 (O_2801,N_43156,N_41772);
and UO_2802 (O_2802,N_44447,N_48952);
nand UO_2803 (O_2803,N_47225,N_44276);
nor UO_2804 (O_2804,N_40040,N_49198);
nand UO_2805 (O_2805,N_46905,N_43636);
nor UO_2806 (O_2806,N_46421,N_40692);
xnor UO_2807 (O_2807,N_40398,N_42628);
xor UO_2808 (O_2808,N_43315,N_47935);
or UO_2809 (O_2809,N_40554,N_41010);
nor UO_2810 (O_2810,N_46843,N_40369);
and UO_2811 (O_2811,N_46642,N_47234);
xnor UO_2812 (O_2812,N_40736,N_46776);
nand UO_2813 (O_2813,N_45803,N_42691);
nor UO_2814 (O_2814,N_43407,N_42447);
nand UO_2815 (O_2815,N_42380,N_44288);
nor UO_2816 (O_2816,N_43972,N_43466);
or UO_2817 (O_2817,N_41069,N_49056);
nand UO_2818 (O_2818,N_40874,N_44542);
xor UO_2819 (O_2819,N_40141,N_41233);
or UO_2820 (O_2820,N_44522,N_45291);
or UO_2821 (O_2821,N_42622,N_42246);
and UO_2822 (O_2822,N_47620,N_43142);
nand UO_2823 (O_2823,N_47252,N_44793);
xor UO_2824 (O_2824,N_44014,N_42259);
xnor UO_2825 (O_2825,N_46882,N_43082);
nor UO_2826 (O_2826,N_46556,N_46355);
and UO_2827 (O_2827,N_46823,N_43752);
nand UO_2828 (O_2828,N_47345,N_48653);
or UO_2829 (O_2829,N_46813,N_48424);
xnor UO_2830 (O_2830,N_47842,N_49620);
or UO_2831 (O_2831,N_48901,N_47107);
or UO_2832 (O_2832,N_45061,N_40992);
nand UO_2833 (O_2833,N_43905,N_40217);
xnor UO_2834 (O_2834,N_48547,N_42252);
xnor UO_2835 (O_2835,N_49909,N_43393);
xnor UO_2836 (O_2836,N_43738,N_40102);
nand UO_2837 (O_2837,N_47644,N_41999);
and UO_2838 (O_2838,N_48170,N_43504);
xor UO_2839 (O_2839,N_44138,N_44344);
or UO_2840 (O_2840,N_44699,N_45544);
and UO_2841 (O_2841,N_45710,N_41105);
nand UO_2842 (O_2842,N_49560,N_48528);
nand UO_2843 (O_2843,N_43893,N_41616);
and UO_2844 (O_2844,N_43231,N_43949);
or UO_2845 (O_2845,N_47384,N_47500);
and UO_2846 (O_2846,N_48529,N_44665);
or UO_2847 (O_2847,N_41467,N_43720);
and UO_2848 (O_2848,N_43785,N_48602);
or UO_2849 (O_2849,N_43655,N_48335);
nand UO_2850 (O_2850,N_45989,N_44837);
and UO_2851 (O_2851,N_40673,N_44458);
or UO_2852 (O_2852,N_45463,N_42575);
xnor UO_2853 (O_2853,N_45838,N_40192);
nor UO_2854 (O_2854,N_43535,N_45969);
nor UO_2855 (O_2855,N_41346,N_43782);
nor UO_2856 (O_2856,N_40654,N_44961);
or UO_2857 (O_2857,N_44941,N_48575);
and UO_2858 (O_2858,N_45240,N_49950);
nand UO_2859 (O_2859,N_41448,N_44375);
or UO_2860 (O_2860,N_47930,N_43931);
nor UO_2861 (O_2861,N_49316,N_47211);
or UO_2862 (O_2862,N_49362,N_46060);
or UO_2863 (O_2863,N_40477,N_49700);
and UO_2864 (O_2864,N_46059,N_46297);
and UO_2865 (O_2865,N_40100,N_45700);
nor UO_2866 (O_2866,N_42915,N_47820);
or UO_2867 (O_2867,N_48396,N_45618);
xor UO_2868 (O_2868,N_45799,N_42242);
or UO_2869 (O_2869,N_49912,N_44769);
xor UO_2870 (O_2870,N_41528,N_46706);
and UO_2871 (O_2871,N_44487,N_46061);
xnor UO_2872 (O_2872,N_45688,N_41867);
or UO_2873 (O_2873,N_43243,N_45864);
and UO_2874 (O_2874,N_41302,N_42649);
and UO_2875 (O_2875,N_48242,N_41234);
nor UO_2876 (O_2876,N_49704,N_43063);
or UO_2877 (O_2877,N_47322,N_49282);
xor UO_2878 (O_2878,N_43975,N_44195);
or UO_2879 (O_2879,N_41211,N_49410);
or UO_2880 (O_2880,N_48369,N_47341);
or UO_2881 (O_2881,N_40570,N_42954);
and UO_2882 (O_2882,N_46154,N_41405);
xor UO_2883 (O_2883,N_43617,N_46685);
or UO_2884 (O_2884,N_43431,N_40198);
nor UO_2885 (O_2885,N_48637,N_44173);
nand UO_2886 (O_2886,N_44849,N_48321);
or UO_2887 (O_2887,N_46529,N_40602);
or UO_2888 (O_2888,N_47427,N_47449);
xor UO_2889 (O_2889,N_47692,N_46633);
nand UO_2890 (O_2890,N_41364,N_44896);
nand UO_2891 (O_2891,N_49433,N_43712);
nand UO_2892 (O_2892,N_43787,N_45294);
and UO_2893 (O_2893,N_45652,N_45772);
xor UO_2894 (O_2894,N_43657,N_44168);
nor UO_2895 (O_2895,N_47535,N_40898);
and UO_2896 (O_2896,N_45502,N_40735);
xnor UO_2897 (O_2897,N_44394,N_46873);
xor UO_2898 (O_2898,N_44217,N_44654);
nor UO_2899 (O_2899,N_41127,N_47456);
and UO_2900 (O_2900,N_42708,N_48647);
nor UO_2901 (O_2901,N_42162,N_40372);
or UO_2902 (O_2902,N_43793,N_47387);
and UO_2903 (O_2903,N_45669,N_49421);
or UO_2904 (O_2904,N_44289,N_46007);
or UO_2905 (O_2905,N_45132,N_44084);
nand UO_2906 (O_2906,N_49422,N_49745);
xor UO_2907 (O_2907,N_40348,N_49835);
xnor UO_2908 (O_2908,N_49534,N_41026);
or UO_2909 (O_2909,N_40890,N_40340);
or UO_2910 (O_2910,N_47231,N_41214);
xnor UO_2911 (O_2911,N_41385,N_42985);
or UO_2912 (O_2912,N_45831,N_47762);
nand UO_2913 (O_2913,N_48105,N_41684);
nand UO_2914 (O_2914,N_42074,N_44876);
and UO_2915 (O_2915,N_43871,N_43500);
or UO_2916 (O_2916,N_49590,N_43316);
nand UO_2917 (O_2917,N_43062,N_43034);
nand UO_2918 (O_2918,N_47701,N_47719);
xor UO_2919 (O_2919,N_47558,N_41025);
or UO_2920 (O_2920,N_42873,N_46048);
and UO_2921 (O_2921,N_47089,N_47576);
nor UO_2922 (O_2922,N_43013,N_48773);
or UO_2923 (O_2923,N_42696,N_45790);
and UO_2924 (O_2924,N_47585,N_47467);
xor UO_2925 (O_2925,N_41101,N_47724);
xor UO_2926 (O_2926,N_46781,N_40491);
and UO_2927 (O_2927,N_41785,N_42763);
or UO_2928 (O_2928,N_41428,N_48645);
xor UO_2929 (O_2929,N_40108,N_48324);
xor UO_2930 (O_2930,N_43313,N_42209);
and UO_2931 (O_2931,N_44639,N_45742);
or UO_2932 (O_2932,N_43515,N_42017);
xor UO_2933 (O_2933,N_42988,N_49692);
xnor UO_2934 (O_2934,N_43285,N_42277);
xor UO_2935 (O_2935,N_40190,N_47676);
nor UO_2936 (O_2936,N_43747,N_42451);
or UO_2937 (O_2937,N_48233,N_46096);
or UO_2938 (O_2938,N_49008,N_44586);
nand UO_2939 (O_2939,N_41472,N_40593);
xor UO_2940 (O_2940,N_43362,N_49547);
xnor UO_2941 (O_2941,N_43043,N_44463);
nor UO_2942 (O_2942,N_43979,N_47100);
nand UO_2943 (O_2943,N_48289,N_43423);
and UO_2944 (O_2944,N_44460,N_48795);
xnor UO_2945 (O_2945,N_41935,N_44117);
nor UO_2946 (O_2946,N_44882,N_44324);
nor UO_2947 (O_2947,N_42821,N_42541);
and UO_2948 (O_2948,N_43249,N_40154);
and UO_2949 (O_2949,N_48008,N_43901);
nand UO_2950 (O_2950,N_44070,N_44762);
nand UO_2951 (O_2951,N_45883,N_42029);
xor UO_2952 (O_2952,N_45402,N_46768);
xor UO_2953 (O_2953,N_43803,N_44451);
and UO_2954 (O_2954,N_43122,N_47718);
nor UO_2955 (O_2955,N_49291,N_41097);
or UO_2956 (O_2956,N_48317,N_49665);
and UO_2957 (O_2957,N_45249,N_49849);
xnor UO_2958 (O_2958,N_48287,N_45895);
nand UO_2959 (O_2959,N_42539,N_44019);
xnor UO_2960 (O_2960,N_41757,N_41436);
nand UO_2961 (O_2961,N_41309,N_46066);
and UO_2962 (O_2962,N_44501,N_41373);
or UO_2963 (O_2963,N_42393,N_46313);
nor UO_2964 (O_2964,N_49479,N_46428);
nor UO_2965 (O_2965,N_45673,N_43087);
nand UO_2966 (O_2966,N_44515,N_48383);
nor UO_2967 (O_2967,N_45381,N_44751);
and UO_2968 (O_2968,N_43357,N_40464);
xor UO_2969 (O_2969,N_41197,N_45938);
xor UO_2970 (O_2970,N_45988,N_45497);
or UO_2971 (O_2971,N_48026,N_43339);
xnor UO_2972 (O_2972,N_44819,N_46837);
xor UO_2973 (O_2973,N_40255,N_48966);
and UO_2974 (O_2974,N_42671,N_47091);
nor UO_2975 (O_2975,N_48137,N_46012);
and UO_2976 (O_2976,N_47512,N_46683);
and UO_2977 (O_2977,N_43229,N_47085);
or UO_2978 (O_2978,N_47809,N_42979);
and UO_2979 (O_2979,N_49462,N_45775);
xnor UO_2980 (O_2980,N_48052,N_49314);
nor UO_2981 (O_2981,N_44852,N_41623);
nand UO_2982 (O_2982,N_48615,N_42213);
nor UO_2983 (O_2983,N_45542,N_40247);
and UO_2984 (O_2984,N_40955,N_45111);
nor UO_2985 (O_2985,N_40809,N_40638);
and UO_2986 (O_2986,N_42855,N_43261);
nand UO_2987 (O_2987,N_41572,N_42195);
nand UO_2988 (O_2988,N_44540,N_44950);
nor UO_2989 (O_2989,N_49470,N_49214);
or UO_2990 (O_2990,N_40752,N_43410);
nor UO_2991 (O_2991,N_48534,N_49178);
xnor UO_2992 (O_2992,N_45242,N_46184);
and UO_2993 (O_2993,N_42478,N_45789);
and UO_2994 (O_2994,N_40617,N_40826);
nor UO_2995 (O_2995,N_41157,N_47791);
xnor UO_2996 (O_2996,N_43439,N_46988);
or UO_2997 (O_2997,N_42306,N_48208);
and UO_2998 (O_2998,N_45889,N_45035);
nand UO_2999 (O_2999,N_40600,N_41884);
or UO_3000 (O_3000,N_46904,N_47376);
nand UO_3001 (O_3001,N_45869,N_43894);
xnor UO_3002 (O_3002,N_48740,N_47835);
and UO_3003 (O_3003,N_48777,N_48640);
or UO_3004 (O_3004,N_44761,N_47261);
xor UO_3005 (O_3005,N_47828,N_45258);
nand UO_3006 (O_3006,N_47084,N_48868);
and UO_3007 (O_3007,N_48299,N_48751);
nand UO_3008 (O_3008,N_49465,N_49965);
nor UO_3009 (O_3009,N_46994,N_47327);
nor UO_3010 (O_3010,N_49783,N_42296);
nor UO_3011 (O_3011,N_48011,N_43185);
xor UO_3012 (O_3012,N_48644,N_45519);
and UO_3013 (O_3013,N_47975,N_45183);
xor UO_3014 (O_3014,N_48227,N_40770);
nor UO_3015 (O_3015,N_46577,N_41672);
xor UO_3016 (O_3016,N_46596,N_45130);
and UO_3017 (O_3017,N_41433,N_42108);
or UO_3018 (O_3018,N_45251,N_49279);
nand UO_3019 (O_3019,N_40905,N_48468);
nor UO_3020 (O_3020,N_49959,N_40560);
xnor UO_3021 (O_3021,N_40084,N_40666);
nor UO_3022 (O_3022,N_41845,N_44086);
nor UO_3023 (O_3023,N_42718,N_44745);
nand UO_3024 (O_3024,N_48676,N_44028);
nor UO_3025 (O_3025,N_40563,N_43519);
nand UO_3026 (O_3026,N_47329,N_48181);
and UO_3027 (O_3027,N_48681,N_40805);
nor UO_3028 (O_3028,N_45843,N_45458);
xor UO_3029 (O_3029,N_44871,N_49372);
and UO_3030 (O_3030,N_43983,N_48340);
xor UO_3031 (O_3031,N_41730,N_46038);
and UO_3032 (O_3032,N_42891,N_45474);
nand UO_3033 (O_3033,N_40009,N_40475);
xor UO_3034 (O_3034,N_45288,N_49439);
or UO_3035 (O_3035,N_42350,N_47279);
xnor UO_3036 (O_3036,N_49020,N_44977);
and UO_3037 (O_3037,N_47184,N_48691);
nor UO_3038 (O_3038,N_46445,N_49270);
nor UO_3039 (O_3039,N_40497,N_43109);
nand UO_3040 (O_3040,N_45571,N_45237);
and UO_3041 (O_3041,N_45072,N_40656);
xor UO_3042 (O_3042,N_48618,N_48969);
xor UO_3043 (O_3043,N_44156,N_41819);
or UO_3044 (O_3044,N_41226,N_41481);
xnor UO_3045 (O_3045,N_43284,N_47706);
nor UO_3046 (O_3046,N_40363,N_40791);
nor UO_3047 (O_3047,N_46085,N_40090);
nand UO_3048 (O_3048,N_48908,N_48162);
xor UO_3049 (O_3049,N_42992,N_42737);
xnor UO_3050 (O_3050,N_45236,N_46425);
and UO_3051 (O_3051,N_48891,N_46568);
or UO_3052 (O_3052,N_47436,N_46317);
or UO_3053 (O_3053,N_44716,N_45452);
xor UO_3054 (O_3054,N_48113,N_44021);
and UO_3055 (O_3055,N_40157,N_41539);
and UO_3056 (O_3056,N_44077,N_47985);
nand UO_3057 (O_3057,N_44007,N_40840);
or UO_3058 (O_3058,N_47458,N_42406);
xnor UO_3059 (O_3059,N_48085,N_44483);
or UO_3060 (O_3060,N_42107,N_48326);
or UO_3061 (O_3061,N_40095,N_40929);
nor UO_3062 (O_3062,N_42640,N_42470);
and UO_3063 (O_3063,N_47132,N_43833);
and UO_3064 (O_3064,N_47798,N_47473);
or UO_3065 (O_3065,N_49926,N_40271);
xor UO_3066 (O_3066,N_46123,N_45116);
xor UO_3067 (O_3067,N_43926,N_42210);
or UO_3068 (O_3068,N_46534,N_46651);
and UO_3069 (O_3069,N_41953,N_43020);
nand UO_3070 (O_3070,N_47229,N_42966);
nor UO_3071 (O_3071,N_44775,N_46524);
and UO_3072 (O_3072,N_48073,N_41982);
and UO_3073 (O_3073,N_42943,N_47756);
xnor UO_3074 (O_3074,N_42879,N_46542);
nor UO_3075 (O_3075,N_43527,N_48290);
nor UO_3076 (O_3076,N_46954,N_46716);
xor UO_3077 (O_3077,N_45832,N_43567);
and UO_3078 (O_3078,N_49424,N_45009);
or UO_3079 (O_3079,N_41998,N_43310);
xnor UO_3080 (O_3080,N_46686,N_49315);
or UO_3081 (O_3081,N_48558,N_41298);
nor UO_3082 (O_3082,N_41190,N_47563);
or UO_3083 (O_3083,N_45830,N_49653);
nand UO_3084 (O_3084,N_42782,N_43809);
or UO_3085 (O_3085,N_41862,N_40888);
and UO_3086 (O_3086,N_45171,N_47459);
nand UO_3087 (O_3087,N_42262,N_40093);
and UO_3088 (O_3088,N_49458,N_46655);
or UO_3089 (O_3089,N_42764,N_49853);
nor UO_3090 (O_3090,N_47495,N_47846);
and UO_3091 (O_3091,N_48421,N_48356);
nand UO_3092 (O_3092,N_43835,N_49348);
nand UO_3093 (O_3093,N_47475,N_44611);
xnor UO_3094 (O_3094,N_42903,N_48328);
xnor UO_3095 (O_3095,N_41398,N_49397);
nor UO_3096 (O_3096,N_42497,N_41175);
nand UO_3097 (O_3097,N_43656,N_45583);
and UO_3098 (O_3098,N_43944,N_45842);
nor UO_3099 (O_3099,N_40339,N_45000);
xor UO_3100 (O_3100,N_43536,N_47407);
or UO_3101 (O_3101,N_48310,N_42341);
or UO_3102 (O_3102,N_41116,N_41110);
nor UO_3103 (O_3103,N_48707,N_48166);
nor UO_3104 (O_3104,N_40230,N_47021);
xnor UO_3105 (O_3105,N_45019,N_49012);
nor UO_3106 (O_3106,N_40750,N_44992);
nand UO_3107 (O_3107,N_45377,N_42785);
and UO_3108 (O_3108,N_46419,N_42403);
nand UO_3109 (O_3109,N_45931,N_41804);
or UO_3110 (O_3110,N_46290,N_41182);
nand UO_3111 (O_3111,N_41114,N_43351);
nor UO_3112 (O_3112,N_44316,N_41142);
nor UO_3113 (O_3113,N_46803,N_47332);
nand UO_3114 (O_3114,N_47732,N_43609);
nand UO_3115 (O_3115,N_48132,N_47862);
xor UO_3116 (O_3116,N_43953,N_45119);
nand UO_3117 (O_3117,N_47386,N_42407);
xnor UO_3118 (O_3118,N_45512,N_48202);
nand UO_3119 (O_3119,N_40993,N_45569);
and UO_3120 (O_3120,N_47664,N_48930);
nand UO_3121 (O_3121,N_41713,N_45012);
nand UO_3122 (O_3122,N_46796,N_42712);
nand UO_3123 (O_3123,N_48772,N_46247);
and UO_3124 (O_3124,N_48042,N_47437);
nor UO_3125 (O_3125,N_42611,N_45510);
nand UO_3126 (O_3126,N_47171,N_47757);
nand UO_3127 (O_3127,N_45540,N_46995);
nor UO_3128 (O_3128,N_43635,N_44434);
xor UO_3129 (O_3129,N_49725,N_45347);
xor UO_3130 (O_3130,N_43646,N_43714);
or UO_3131 (O_3131,N_49585,N_45169);
xor UO_3132 (O_3132,N_41027,N_45110);
xor UO_3133 (O_3133,N_44883,N_40395);
nand UO_3134 (O_3134,N_41561,N_43451);
and UO_3135 (O_3135,N_43813,N_45580);
xnor UO_3136 (O_3136,N_43820,N_44675);
nand UO_3137 (O_3137,N_48864,N_49870);
xor UO_3138 (O_3138,N_48614,N_40696);
nor UO_3139 (O_3139,N_48034,N_44215);
xor UO_3140 (O_3140,N_45428,N_46016);
nor UO_3141 (O_3141,N_47955,N_45665);
xnor UO_3142 (O_3142,N_47654,N_47262);
nand UO_3143 (O_3143,N_44484,N_44089);
xnor UO_3144 (O_3144,N_45882,N_45283);
and UO_3145 (O_3145,N_48716,N_41579);
xnor UO_3146 (O_3146,N_43502,N_48325);
nor UO_3147 (O_3147,N_40575,N_40409);
nor UO_3148 (O_3148,N_43151,N_48736);
nor UO_3149 (O_3149,N_48402,N_41548);
or UO_3150 (O_3150,N_43740,N_46341);
or UO_3151 (O_3151,N_46229,N_42773);
nand UO_3152 (O_3152,N_42353,N_40098);
nor UO_3153 (O_3153,N_47098,N_41514);
and UO_3154 (O_3154,N_45679,N_49103);
and UO_3155 (O_3155,N_48364,N_47154);
nor UO_3156 (O_3156,N_48398,N_48717);
nor UO_3157 (O_3157,N_40085,N_45143);
xnor UO_3158 (O_3158,N_44939,N_43455);
and UO_3159 (O_3159,N_45971,N_42217);
nor UO_3160 (O_3160,N_48160,N_42197);
or UO_3161 (O_3161,N_44029,N_40646);
xor UO_3162 (O_3162,N_46431,N_42387);
nor UO_3163 (O_3163,N_48007,N_49288);
xnor UO_3164 (O_3164,N_49150,N_47800);
or UO_3165 (O_3165,N_49832,N_45040);
nor UO_3166 (O_3166,N_43246,N_46262);
nor UO_3167 (O_3167,N_49009,N_46466);
nor UO_3168 (O_3168,N_49703,N_45715);
and UO_3169 (O_3169,N_41892,N_49358);
and UO_3170 (O_3170,N_49984,N_43816);
xnor UO_3171 (O_3171,N_46211,N_44128);
nand UO_3172 (O_3172,N_46982,N_45303);
and UO_3173 (O_3173,N_41775,N_40657);
xor UO_3174 (O_3174,N_45314,N_45485);
nand UO_3175 (O_3175,N_49473,N_41985);
nand UO_3176 (O_3176,N_49116,N_41464);
nand UO_3177 (O_3177,N_42571,N_45947);
xnor UO_3178 (O_3178,N_46600,N_45100);
or UO_3179 (O_3179,N_42110,N_49537);
or UO_3180 (O_3180,N_48460,N_40866);
and UO_3181 (O_3181,N_43819,N_49632);
nand UO_3182 (O_3182,N_45627,N_44049);
or UO_3183 (O_3183,N_49600,N_46144);
and UO_3184 (O_3184,N_45121,N_42031);
or UO_3185 (O_3185,N_43441,N_44776);
and UO_3186 (O_3186,N_42219,N_49602);
xor UO_3187 (O_3187,N_46806,N_48498);
or UO_3188 (O_3188,N_42136,N_44058);
or UO_3189 (O_3189,N_44212,N_47914);
or UO_3190 (O_3190,N_49819,N_49309);
or UO_3191 (O_3191,N_44175,N_41613);
xor UO_3192 (O_3192,N_46669,N_43242);
nand UO_3193 (O_3193,N_40083,N_48206);
nand UO_3194 (O_3194,N_47027,N_43236);
nand UO_3195 (O_3195,N_41130,N_48567);
xnor UO_3196 (O_3196,N_45309,N_41808);
and UO_3197 (O_3197,N_44122,N_48745);
and UO_3198 (O_3198,N_43834,N_42665);
or UO_3199 (O_3199,N_47694,N_44472);
or UO_3200 (O_3200,N_41008,N_44448);
xor UO_3201 (O_3201,N_49922,N_47522);
nor UO_3202 (O_3202,N_41117,N_45006);
nand UO_3203 (O_3203,N_44502,N_45427);
xor UO_3204 (O_3204,N_40645,N_47440);
or UO_3205 (O_3205,N_46736,N_41222);
nor UO_3206 (O_3206,N_43924,N_47460);
or UO_3207 (O_3207,N_41552,N_44553);
nand UO_3208 (O_3208,N_47942,N_42667);
and UO_3209 (O_3209,N_40775,N_45792);
nand UO_3210 (O_3210,N_41811,N_46169);
nor UO_3211 (O_3211,N_46072,N_41002);
nor UO_3212 (O_3212,N_46077,N_46900);
nor UO_3213 (O_3213,N_45982,N_43275);
nand UO_3214 (O_3214,N_49929,N_46408);
or UO_3215 (O_3215,N_47686,N_43896);
or UO_3216 (O_3216,N_49028,N_41149);
or UO_3217 (O_3217,N_40849,N_46087);
or UO_3218 (O_3218,N_41316,N_43306);
nand UO_3219 (O_3219,N_47050,N_42863);
and UO_3220 (O_3220,N_44835,N_40872);
nand UO_3221 (O_3221,N_49415,N_47003);
xnor UO_3222 (O_3222,N_49324,N_49403);
nand UO_3223 (O_3223,N_42941,N_40092);
or UO_3224 (O_3224,N_44936,N_45318);
xnor UO_3225 (O_3225,N_42344,N_45717);
or UO_3226 (O_3226,N_44938,N_48556);
or UO_3227 (O_3227,N_43951,N_40701);
xnor UO_3228 (O_3228,N_46487,N_41325);
nor UO_3229 (O_3229,N_49896,N_46119);
or UO_3230 (O_3230,N_40060,N_42233);
xnor UO_3231 (O_3231,N_41697,N_43561);
or UO_3232 (O_3232,N_49167,N_49398);
and UO_3233 (O_3233,N_46974,N_44171);
or UO_3234 (O_3234,N_48408,N_41206);
nand UO_3235 (O_3235,N_42318,N_43857);
nand UO_3236 (O_3236,N_42194,N_43856);
and UO_3237 (O_3237,N_43023,N_49208);
xnor UO_3238 (O_3238,N_48349,N_42130);
and UO_3239 (O_3239,N_46748,N_42625);
or UO_3240 (O_3240,N_47010,N_44514);
or UO_3241 (O_3241,N_46512,N_47682);
or UO_3242 (O_3242,N_42327,N_46316);
nand UO_3243 (O_3243,N_45892,N_46417);
nand UO_3244 (O_3244,N_41914,N_42532);
xor UO_3245 (O_3245,N_45260,N_46514);
or UO_3246 (O_3246,N_42917,N_40406);
nor UO_3247 (O_3247,N_44220,N_44532);
or UO_3248 (O_3248,N_41968,N_48226);
xnor UO_3249 (O_3249,N_43739,N_45286);
and UO_3250 (O_3250,N_43031,N_48616);
or UO_3251 (O_3251,N_45681,N_48843);
and UO_3252 (O_3252,N_44659,N_49589);
nor UO_3253 (O_3253,N_47196,N_49952);
nand UO_3254 (O_3254,N_45766,N_43247);
or UO_3255 (O_3255,N_40246,N_44233);
xor UO_3256 (O_3256,N_44642,N_45522);
and UO_3257 (O_3257,N_44858,N_44507);
nand UO_3258 (O_3258,N_41006,N_40097);
or UO_3259 (O_3259,N_41129,N_41047);
and UO_3260 (O_3260,N_48853,N_40884);
or UO_3261 (O_3261,N_43556,N_41660);
nor UO_3262 (O_3262,N_42894,N_46266);
and UO_3263 (O_3263,N_41254,N_46801);
nand UO_3264 (O_3264,N_41685,N_46081);
and UO_3265 (O_3265,N_41724,N_40062);
or UO_3266 (O_3266,N_41763,N_43356);
and UO_3267 (O_3267,N_46250,N_48896);
or UO_3268 (O_3268,N_47255,N_43913);
nor UO_3269 (O_3269,N_42493,N_40330);
xor UO_3270 (O_3270,N_43186,N_46933);
xor UO_3271 (O_3271,N_49662,N_40742);
nand UO_3272 (O_3272,N_40045,N_43613);
xnor UO_3273 (O_3273,N_45178,N_44786);
xnor UO_3274 (O_3274,N_49916,N_49413);
nand UO_3275 (O_3275,N_40556,N_48251);
nor UO_3276 (O_3276,N_49353,N_46682);
and UO_3277 (O_3277,N_43526,N_43703);
or UO_3278 (O_3278,N_49395,N_49339);
nand UO_3279 (O_3279,N_47209,N_44614);
nand UO_3280 (O_3280,N_49908,N_43978);
nor UO_3281 (O_3281,N_43079,N_44526);
xnor UO_3282 (O_3282,N_44281,N_43849);
xnor UO_3283 (O_3283,N_42275,N_48559);
nand UO_3284 (O_3284,N_45036,N_47263);
nand UO_3285 (O_3285,N_44730,N_49734);
nor UO_3286 (O_3286,N_46346,N_40524);
nand UO_3287 (O_3287,N_45505,N_40761);
or UO_3288 (O_3288,N_42826,N_48568);
and UO_3289 (O_3289,N_44187,N_42914);
nand UO_3290 (O_3290,N_44813,N_42606);
xor UO_3291 (O_3291,N_40079,N_40528);
nand UO_3292 (O_3292,N_44346,N_47028);
xnor UO_3293 (O_3293,N_48382,N_47600);
and UO_3294 (O_3294,N_43184,N_40484);
nor UO_3295 (O_3295,N_43572,N_43722);
nand UO_3296 (O_3296,N_40865,N_44804);
nand UO_3297 (O_3297,N_43391,N_49311);
nand UO_3298 (O_3298,N_41917,N_47923);
or UO_3299 (O_3299,N_48104,N_46132);
xor UO_3300 (O_3300,N_41544,N_43696);
xor UO_3301 (O_3301,N_46666,N_49659);
nand UO_3302 (O_3302,N_47766,N_48994);
or UO_3303 (O_3303,N_49739,N_46325);
and UO_3304 (O_3304,N_44011,N_48103);
xor UO_3305 (O_3305,N_45127,N_43475);
and UO_3306 (O_3306,N_44842,N_49166);
nor UO_3307 (O_3307,N_43596,N_43258);
or UO_3308 (O_3308,N_48400,N_42607);
xor UO_3309 (O_3309,N_46434,N_47943);
nand UO_3310 (O_3310,N_48385,N_47277);
or UO_3311 (O_3311,N_45131,N_41945);
nor UO_3312 (O_3312,N_48050,N_42949);
or UO_3313 (O_3313,N_46240,N_45719);
or UO_3314 (O_3314,N_42702,N_40216);
nor UO_3315 (O_3315,N_43643,N_49074);
or UO_3316 (O_3316,N_45706,N_43028);
and UO_3317 (O_3317,N_46205,N_48512);
nor UO_3318 (O_3318,N_42659,N_42480);
or UO_3319 (O_3319,N_42166,N_45361);
nand UO_3320 (O_3320,N_41639,N_49173);
nor UO_3321 (O_3321,N_49332,N_49715);
nand UO_3322 (O_3322,N_48728,N_40153);
and UO_3323 (O_3323,N_44727,N_41203);
and UO_3324 (O_3324,N_46332,N_47267);
nand UO_3325 (O_3325,N_40948,N_43112);
xor UO_3326 (O_3326,N_44640,N_42830);
nor UO_3327 (O_3327,N_45812,N_40444);
or UO_3328 (O_3328,N_47612,N_44584);
nor UO_3329 (O_3329,N_47758,N_44833);
nand UO_3330 (O_3330,N_40471,N_49494);
or UO_3331 (O_3331,N_45584,N_49504);
and UO_3332 (O_3332,N_44131,N_48012);
nand UO_3333 (O_3333,N_41764,N_45538);
nor UO_3334 (O_3334,N_43411,N_47743);
nor UO_3335 (O_3335,N_42402,N_49010);
nor UO_3336 (O_3336,N_40547,N_44441);
xor UO_3337 (O_3337,N_44862,N_42442);
nor UO_3338 (O_3338,N_49716,N_43611);
or UO_3339 (O_3339,N_42956,N_48938);
or UO_3340 (O_3340,N_41282,N_49034);
and UO_3341 (O_3341,N_47681,N_48404);
and UO_3342 (O_3342,N_47128,N_46022);
and UO_3343 (O_3343,N_48117,N_45470);
or UO_3344 (O_3344,N_43456,N_43083);
nand UO_3345 (O_3345,N_42334,N_42307);
nand UO_3346 (O_3346,N_49425,N_49535);
or UO_3347 (O_3347,N_44034,N_42524);
or UO_3348 (O_3348,N_43573,N_49466);
and UO_3349 (O_3349,N_43771,N_48186);
nor UO_3350 (O_3350,N_47959,N_46809);
xor UO_3351 (O_3351,N_42933,N_40063);
and UO_3352 (O_3352,N_46099,N_44700);
or UO_3353 (O_3353,N_40304,N_42142);
nor UO_3354 (O_3354,N_44080,N_43420);
nor UO_3355 (O_3355,N_43826,N_45146);
and UO_3356 (O_3356,N_49943,N_49204);
and UO_3357 (O_3357,N_44854,N_45678);
nand UO_3358 (O_3358,N_47463,N_47643);
nand UO_3359 (O_3359,N_47408,N_49794);
nor UO_3360 (O_3360,N_49824,N_40514);
or UO_3361 (O_3361,N_46374,N_45081);
or UO_3362 (O_3362,N_43528,N_44760);
or UO_3363 (O_3363,N_40687,N_44304);
nor UO_3364 (O_3364,N_48936,N_43829);
or UO_3365 (O_3365,N_49934,N_48167);
and UO_3366 (O_3366,N_45088,N_41231);
nor UO_3367 (O_3367,N_45345,N_42817);
and UO_3368 (O_3368,N_48487,N_48661);
or UO_3369 (O_3369,N_41989,N_43731);
xnor UO_3370 (O_3370,N_48342,N_48972);
xnor UO_3371 (O_3371,N_45844,N_44531);
nor UO_3372 (O_3372,N_48649,N_45390);
nor UO_3373 (O_3373,N_46607,N_40436);
nor UO_3374 (O_3374,N_40008,N_44825);
nand UO_3375 (O_3375,N_44676,N_41120);
or UO_3376 (O_3376,N_46287,N_47934);
nor UO_3377 (O_3377,N_45045,N_40852);
nand UO_3378 (O_3378,N_43477,N_47981);
and UO_3379 (O_3379,N_46690,N_49528);
xnor UO_3380 (O_3380,N_42986,N_48856);
nand UO_3381 (O_3381,N_49816,N_48045);
nand UO_3382 (O_3382,N_44165,N_46846);
nand UO_3383 (O_3383,N_42324,N_46412);
nand UO_3384 (O_3384,N_49961,N_49968);
xnor UO_3385 (O_3385,N_43272,N_49717);
nand UO_3386 (O_3386,N_46040,N_42392);
and UO_3387 (O_3387,N_46545,N_44697);
nand UO_3388 (O_3388,N_42833,N_45225);
nand UO_3389 (O_3389,N_47818,N_47065);
nand UO_3390 (O_3390,N_40005,N_48927);
nand UO_3391 (O_3391,N_47076,N_41263);
xor UO_3392 (O_3392,N_42660,N_49492);
xnor UO_3393 (O_3393,N_40254,N_46725);
nor UO_3394 (O_3394,N_42560,N_45628);
xor UO_3395 (O_3395,N_40518,N_42456);
and UO_3396 (O_3396,N_46652,N_43173);
nand UO_3397 (O_3397,N_40783,N_46930);
nand UO_3398 (O_3398,N_40717,N_41580);
and UO_3399 (O_3399,N_46439,N_47592);
or UO_3400 (O_3400,N_49791,N_43014);
nor UO_3401 (O_3401,N_40345,N_40276);
nand UO_3402 (O_3402,N_47420,N_48633);
nor UO_3403 (O_3403,N_46946,N_47948);
or UO_3404 (O_3404,N_41453,N_42316);
nor UO_3405 (O_3405,N_49445,N_49498);
xnor UO_3406 (O_3406,N_45271,N_42299);
and UO_3407 (O_3407,N_45029,N_43525);
nand UO_3408 (O_3408,N_48277,N_44968);
xor UO_3409 (O_3409,N_46944,N_42546);
or UO_3410 (O_3410,N_48044,N_47353);
xnor UO_3411 (O_3411,N_47665,N_46693);
or UO_3412 (O_3412,N_47759,N_45472);
nand UO_3413 (O_3413,N_47893,N_49861);
or UO_3414 (O_3414,N_46041,N_48376);
or UO_3415 (O_3415,N_44841,N_41084);
or UO_3416 (O_3416,N_44643,N_46444);
nor UO_3417 (O_3417,N_43673,N_40683);
and UO_3418 (O_3418,N_47870,N_45410);
nand UO_3419 (O_3419,N_48596,N_48482);
xor UO_3420 (O_3420,N_42778,N_44486);
nand UO_3421 (O_3421,N_42076,N_48696);
nand UO_3422 (O_3422,N_48192,N_48639);
nand UO_3423 (O_3423,N_41951,N_45256);
nor UO_3424 (O_3424,N_41343,N_45287);
nand UO_3425 (O_3425,N_44693,N_46957);
or UO_3426 (O_3426,N_40161,N_44236);
xor UO_3427 (O_3427,N_43994,N_40932);
xor UO_3428 (O_3428,N_44230,N_44891);
xor UO_3429 (O_3429,N_43845,N_48595);
or UO_3430 (O_3430,N_44646,N_41825);
and UO_3431 (O_3431,N_44258,N_48682);
xnor UO_3432 (O_3432,N_46480,N_46273);
nand UO_3433 (O_3433,N_42395,N_47772);
or UO_3434 (O_3434,N_47298,N_45138);
xnor UO_3435 (O_3435,N_49887,N_42431);
or UO_3436 (O_3436,N_44748,N_40485);
and UO_3437 (O_3437,N_40853,N_40158);
xnor UO_3438 (O_3438,N_49820,N_48585);
nor UO_3439 (O_3439,N_42305,N_47323);
and UO_3440 (O_3440,N_48702,N_43235);
and UO_3441 (O_3441,N_43595,N_45195);
and UO_3442 (O_3442,N_42945,N_40077);
nand UO_3443 (O_3443,N_43709,N_46569);
and UO_3444 (O_3444,N_46670,N_47187);
and UO_3445 (O_3445,N_41388,N_44873);
or UO_3446 (O_3446,N_46613,N_48203);
xnor UO_3447 (O_3447,N_46921,N_40186);
or UO_3448 (O_3448,N_44235,N_44615);
or UO_3449 (O_3449,N_42241,N_44571);
and UO_3450 (O_3450,N_44248,N_41503);
or UO_3451 (O_3451,N_44012,N_43586);
nor UO_3452 (O_3452,N_43129,N_44016);
nand UO_3453 (O_3453,N_43610,N_44025);
or UO_3454 (O_3454,N_41534,N_40665);
or UO_3455 (O_3455,N_47545,N_40086);
nand UO_3456 (O_3456,N_41663,N_41345);
xor UO_3457 (O_3457,N_49432,N_42716);
nor UO_3458 (O_3458,N_43936,N_42908);
or UO_3459 (O_3459,N_41594,N_49330);
nand UO_3460 (O_3460,N_49866,N_47794);
nand UO_3461 (O_3461,N_47094,N_49694);
and UO_3462 (O_3462,N_48656,N_41600);
xor UO_3463 (O_3463,N_45465,N_41400);
nand UO_3464 (O_3464,N_43830,N_44341);
and UO_3465 (O_3465,N_40707,N_46409);
nand UO_3466 (O_3466,N_49134,N_48357);
nor UO_3467 (O_3467,N_48370,N_45405);
nor UO_3468 (O_3468,N_44421,N_47812);
xor UO_3469 (O_3469,N_47015,N_44104);
nand UO_3470 (O_3470,N_45888,N_46398);
xor UO_3471 (O_3471,N_47890,N_42040);
xnor UO_3472 (O_3472,N_47971,N_41482);
nand UO_3473 (O_3473,N_47826,N_46897);
or UO_3474 (O_3474,N_45609,N_47910);
or UO_3475 (O_3475,N_44605,N_47944);
or UO_3476 (O_3476,N_49195,N_43418);
or UO_3477 (O_3477,N_49414,N_48767);
xnor UO_3478 (O_3478,N_40076,N_49038);
xor UO_3479 (O_3479,N_45461,N_47527);
xnor UO_3480 (O_3480,N_46898,N_40841);
nand UO_3481 (O_3481,N_47172,N_44048);
xor UO_3482 (O_3482,N_40300,N_45358);
nand UO_3483 (O_3483,N_46523,N_41665);
xnor UO_3484 (O_3484,N_46573,N_48957);
or UO_3485 (O_3485,N_48439,N_44046);
xnor UO_3486 (O_3486,N_48405,N_45698);
nor UO_3487 (O_3487,N_49050,N_48410);
nor UO_3488 (O_3488,N_45899,N_47451);
nand UO_3489 (O_3489,N_40680,N_47877);
xnor UO_3490 (O_3490,N_43329,N_40103);
or UO_3491 (O_3491,N_46280,N_41913);
xor UO_3492 (O_3492,N_41499,N_47597);
xor UO_3493 (O_3493,N_45011,N_44139);
and UO_3494 (O_3494,N_47544,N_40411);
xnor UO_3495 (O_3495,N_41200,N_46811);
nor UO_3496 (O_3496,N_43125,N_46464);
nor UO_3497 (O_3497,N_41883,N_47949);
or UO_3498 (O_3498,N_41264,N_42390);
and UO_3499 (O_3499,N_49760,N_42549);
nand UO_3500 (O_3500,N_45937,N_49677);
or UO_3501 (O_3501,N_41877,N_46492);
and UO_3502 (O_3502,N_42168,N_49093);
and UO_3503 (O_3503,N_46239,N_43190);
xnor UO_3504 (O_3504,N_44302,N_47004);
or UO_3505 (O_3505,N_47186,N_41556);
nand UO_3506 (O_3506,N_45289,N_44467);
nand UO_3507 (O_3507,N_42765,N_40269);
or UO_3508 (O_3508,N_46321,N_45102);
nand UO_3509 (O_3509,N_48463,N_44426);
nor UO_3510 (O_3510,N_49382,N_43602);
nor UO_3511 (O_3511,N_46509,N_45489);
nand UO_3512 (O_3512,N_47578,N_42994);
or UO_3513 (O_3513,N_44550,N_49502);
nor UO_3514 (O_3514,N_46448,N_43221);
or UO_3515 (O_3515,N_46243,N_44999);
or UO_3516 (O_3516,N_45450,N_48959);
nand UO_3517 (O_3517,N_49691,N_47568);
or UO_3518 (O_3518,N_44737,N_44702);
xnor UO_3519 (O_3519,N_46960,N_41474);
xnor UO_3520 (O_3520,N_40558,N_42409);
nor UO_3521 (O_3521,N_49969,N_40926);
or UO_3522 (O_3522,N_49738,N_47057);
xor UO_3523 (O_3523,N_43019,N_47604);
or UO_3524 (O_3524,N_45137,N_41118);
nor UO_3525 (O_3525,N_49058,N_47733);
nand UO_3526 (O_3526,N_49526,N_41365);
nor UO_3527 (O_3527,N_44843,N_42328);
nor UO_3528 (O_3528,N_43036,N_41489);
or UO_3529 (O_3529,N_43208,N_47817);
and UO_3530 (O_3530,N_48590,N_48945);
nand UO_3531 (O_3531,N_41053,N_42496);
xnor UO_3532 (O_3532,N_42896,N_49663);
nand UO_3533 (O_3533,N_49448,N_45444);
nand UO_3534 (O_3534,N_41637,N_47509);
and UO_3535 (O_3535,N_47823,N_43633);
nor UO_3536 (O_3536,N_41153,N_45339);
or UO_3537 (O_3537,N_47621,N_46753);
nand UO_3538 (O_3538,N_48158,N_49515);
xnor UO_3539 (O_3539,N_40814,N_47895);
and UO_3540 (O_3540,N_40342,N_41360);
or UO_3541 (O_3541,N_41229,N_41627);
xor UO_3542 (O_3542,N_47079,N_43593);
xnor UO_3543 (O_3543,N_47101,N_45704);
nor UO_3544 (O_3544,N_46720,N_40068);
nor UO_3545 (O_3545,N_42205,N_49960);
nor UO_3546 (O_3546,N_46071,N_41372);
nor UO_3547 (O_3547,N_48475,N_46805);
nor UO_3548 (O_3548,N_40360,N_49540);
or UO_3549 (O_3549,N_49990,N_44282);
nor UO_3550 (O_3550,N_45034,N_40962);
and UO_3551 (O_3551,N_46120,N_41189);
or UO_3552 (O_3552,N_43651,N_40739);
and UO_3553 (O_3553,N_44696,N_41251);
nand UO_3554 (O_3554,N_40901,N_41417);
nand UO_3555 (O_3555,N_43570,N_44275);
nor UO_3556 (O_3556,N_49190,N_47907);
or UO_3557 (O_3557,N_47716,N_47699);
xor UO_3558 (O_3558,N_43840,N_40580);
nor UO_3559 (O_3559,N_47871,N_40206);
or UO_3560 (O_3560,N_49293,N_40503);
nand UO_3561 (O_3561,N_43133,N_48232);
nor UO_3562 (O_3562,N_42035,N_43076);
xnor UO_3563 (O_3563,N_41816,N_43766);
and UO_3564 (O_3564,N_49070,N_46859);
xor UO_3565 (O_3565,N_41863,N_45535);
or UO_3566 (O_3566,N_44323,N_42512);
xnor UO_3567 (O_3567,N_40582,N_44664);
and UO_3568 (O_3568,N_48688,N_43163);
xor UO_3569 (O_3569,N_46219,N_44690);
nand UO_3570 (O_3570,N_48712,N_49265);
or UO_3571 (O_3571,N_43581,N_43369);
nor UO_3572 (O_3572,N_48983,N_43071);
and UO_3573 (O_3573,N_46116,N_45142);
or UO_3574 (O_3574,N_41286,N_42796);
nand UO_3575 (O_3575,N_44158,N_44343);
xor UO_3576 (O_3576,N_42038,N_46968);
nand UO_3577 (O_3577,N_42724,N_46311);
or UO_3578 (O_3578,N_40611,N_43210);
nor UO_3579 (O_3579,N_46565,N_47268);
and UO_3580 (O_3580,N_49238,N_49979);
and UO_3581 (O_3581,N_48695,N_41494);
xnor UO_3582 (O_3582,N_46620,N_46122);
xnor UO_3583 (O_3583,N_47635,N_41393);
and UO_3584 (O_3584,N_41981,N_42272);
xor UO_3585 (O_3585,N_40013,N_41208);
nand UO_3586 (O_3586,N_43796,N_42122);
xor UO_3587 (O_3587,N_46406,N_48925);
xor UO_3588 (O_3588,N_46000,N_48642);
and UO_3589 (O_3589,N_45017,N_43888);
or UO_3590 (O_3590,N_49197,N_41059);
nor UO_3591 (O_3591,N_45884,N_49685);
or UO_3592 (O_3592,N_42154,N_44435);
and UO_3593 (O_3593,N_46383,N_45651);
xnor UO_3594 (O_3594,N_47248,N_44774);
nor UO_3595 (O_3595,N_41809,N_40601);
or UO_3596 (O_3596,N_44163,N_47245);
nand UO_3597 (O_3597,N_45866,N_42730);
nor UO_3598 (O_3598,N_49894,N_46389);
nor UO_3599 (O_3599,N_41524,N_46741);
xor UO_3600 (O_3600,N_42508,N_48175);
or UO_3601 (O_3601,N_45608,N_40032);
nor UO_3602 (O_3602,N_45795,N_49100);
nor UO_3603 (O_3603,N_49512,N_49562);
nand UO_3604 (O_3604,N_49750,N_47536);
or UO_3605 (O_3605,N_40042,N_40634);
nor UO_3606 (O_3606,N_44140,N_48849);
xor UO_3607 (O_3607,N_44821,N_41173);
xnor UO_3608 (O_3608,N_41389,N_44602);
xnor UO_3609 (O_3609,N_49910,N_40903);
and UO_3610 (O_3610,N_40162,N_42831);
nor UO_3611 (O_3611,N_42513,N_40561);
or UO_3612 (O_3612,N_48760,N_40329);
or UO_3613 (O_3613,N_48914,N_41606);
nand UO_3614 (O_3614,N_47379,N_42383);
and UO_3615 (O_3615,N_42869,N_46998);
and UO_3616 (O_3616,N_42346,N_43929);
nor UO_3617 (O_3617,N_42800,N_42007);
xnor UO_3618 (O_3618,N_40693,N_43259);
xor UO_3619 (O_3619,N_47471,N_45554);
and UO_3620 (O_3620,N_40415,N_46755);
and UO_3621 (O_3621,N_40118,N_41786);
nor UO_3622 (O_3622,N_41952,N_44263);
nand UO_3623 (O_3623,N_45855,N_41355);
xor UO_3624 (O_3624,N_46615,N_45070);
nor UO_3625 (O_3625,N_49376,N_43966);
nor UO_3626 (O_3626,N_46026,N_41350);
xor UO_3627 (O_3627,N_48250,N_43298);
nand UO_3628 (O_3628,N_42558,N_44556);
xor UO_3629 (O_3629,N_42477,N_43191);
or UO_3630 (O_3630,N_47469,N_48655);
nand UO_3631 (O_3631,N_46742,N_45145);
nand UO_3632 (O_3632,N_47362,N_45758);
nand UO_3633 (O_3633,N_41729,N_49143);
and UO_3634 (O_3634,N_42157,N_46260);
nand UO_3635 (O_3635,N_49402,N_45417);
nand UO_3636 (O_3636,N_49581,N_43879);
nand UO_3637 (O_3637,N_45401,N_46727);
nand UO_3638 (O_3638,N_48286,N_49269);
or UO_3639 (O_3639,N_49999,N_43822);
xnor UO_3640 (O_3640,N_40844,N_42520);
nor UO_3641 (O_3641,N_45115,N_48080);
xor UO_3642 (O_3642,N_44413,N_47404);
nand UO_3643 (O_3643,N_41152,N_42028);
and UO_3644 (O_3644,N_46654,N_47309);
xnor UO_3645 (O_3645,N_40213,N_48102);
nand UO_3646 (O_3646,N_46373,N_41577);
nor UO_3647 (O_3647,N_45979,N_40507);
nor UO_3648 (O_3648,N_43654,N_44966);
nand UO_3649 (O_3649,N_44723,N_47017);
nand UO_3650 (O_3650,N_41520,N_44155);
nand UO_3651 (O_3651,N_45550,N_44213);
nand UO_3652 (O_3652,N_45887,N_40094);
or UO_3653 (O_3653,N_43601,N_41082);
nor UO_3654 (O_3654,N_42323,N_41057);
nand UO_3655 (O_3655,N_43802,N_43938);
nor UO_3656 (O_3656,N_47610,N_47227);
xor UO_3657 (O_3657,N_40149,N_45243);
or UO_3658 (O_3658,N_41686,N_49307);
xor UO_3659 (O_3659,N_42057,N_47257);
or UO_3660 (O_3660,N_47505,N_45693);
and UO_3661 (O_3661,N_48061,N_46643);
or UO_3662 (O_3662,N_47025,N_43262);
or UO_3663 (O_3663,N_40417,N_42832);
nand UO_3664 (O_3664,N_47574,N_48950);
xnor UO_3665 (O_3665,N_43039,N_48474);
nor UO_3666 (O_3666,N_48955,N_40523);
nand UO_3667 (O_3667,N_45784,N_49383);
and UO_3668 (O_3668,N_45731,N_45310);
and UO_3669 (O_3669,N_42900,N_42001);
xnor UO_3670 (O_3670,N_47989,N_45262);
or UO_3671 (O_3671,N_49626,N_41860);
xnor UO_3672 (O_3672,N_49430,N_47903);
xor UO_3673 (O_3673,N_44219,N_41687);
nand UO_3674 (O_3674,N_41070,N_45837);
xnor UO_3675 (O_3675,N_44197,N_48390);
or UO_3676 (O_3676,N_47215,N_45122);
or UO_3677 (O_3677,N_49536,N_41445);
nor UO_3678 (O_3678,N_46367,N_41832);
nor UO_3679 (O_3679,N_49030,N_44907);
nor UO_3680 (O_3680,N_40223,N_48570);
nor UO_3681 (O_3681,N_44790,N_42116);
and UO_3682 (O_3682,N_48922,N_49939);
and UO_3683 (O_3683,N_40248,N_44293);
nor UO_3684 (O_3684,N_44983,N_45181);
nor UO_3685 (O_3685,N_41477,N_46358);
xor UO_3686 (O_3686,N_44349,N_43050);
nand UO_3687 (O_3687,N_43145,N_40309);
nand UO_3688 (O_3688,N_46293,N_42865);
xnor UO_3689 (O_3689,N_49579,N_44381);
nor UO_3690 (O_3690,N_40221,N_49169);
xnor UO_3691 (O_3691,N_44682,N_42070);
xor UO_3692 (O_3692,N_49071,N_40511);
nand UO_3693 (O_3693,N_44764,N_45164);
or UO_3694 (O_3694,N_43577,N_43325);
nand UO_3695 (O_3695,N_40307,N_48532);
or UO_3696 (O_3696,N_47869,N_49292);
and UO_3697 (O_3697,N_48774,N_44241);
xnor UO_3698 (O_3698,N_42082,N_41975);
xor UO_3699 (O_3699,N_49280,N_47390);
and UO_3700 (O_3700,N_40618,N_40686);
nand UO_3701 (O_3701,N_48819,N_44301);
nor UO_3702 (O_3702,N_42784,N_46404);
nand UO_3703 (O_3703,N_44922,N_46034);
nand UO_3704 (O_3704,N_40430,N_48863);
nand UO_3705 (O_3705,N_48806,N_41741);
nand UO_3706 (O_3706,N_47195,N_47210);
nor UO_3707 (O_3707,N_40355,N_43821);
xor UO_3708 (O_3708,N_46647,N_47072);
nor UO_3709 (O_3709,N_45201,N_49821);
nand UO_3710 (O_3710,N_42247,N_45092);
or UO_3711 (O_3711,N_46814,N_47618);
xnor UO_3712 (O_3712,N_49213,N_48211);
and UO_3713 (O_3713,N_47698,N_46836);
or UO_3714 (O_3714,N_44606,N_46619);
xor UO_3715 (O_3715,N_44738,N_41517);
nor UO_3716 (O_3716,N_40534,N_46917);
and UO_3717 (O_3717,N_45919,N_43338);
nand UO_3718 (O_3718,N_45732,N_48915);
xor UO_3719 (O_3719,N_46118,N_45388);
or UO_3720 (O_3720,N_42484,N_41501);
and UO_3721 (O_3721,N_48347,N_45326);
nand UO_3722 (O_3722,N_40191,N_46989);
or UO_3723 (O_3723,N_40268,N_40574);
xnor UO_3724 (O_3724,N_49235,N_40889);
xor UO_3725 (O_3725,N_47370,N_42550);
nor UO_3726 (O_3726,N_41290,N_40919);
xor UO_3727 (O_3727,N_47799,N_49635);
and UO_3728 (O_3728,N_42673,N_47844);
or UO_3729 (O_3729,N_44758,N_42479);
nor UO_3730 (O_3730,N_45170,N_47177);
nor UO_3731 (O_3731,N_42844,N_43982);
and UO_3732 (O_3732,N_49370,N_43319);
nand UO_3733 (O_3733,N_47314,N_43436);
nand UO_3734 (O_3734,N_44900,N_44692);
nand UO_3735 (O_3735,N_43040,N_40771);
nand UO_3736 (O_3736,N_42906,N_43960);
and UO_3737 (O_3737,N_49226,N_48522);
nor UO_3738 (O_3738,N_49452,N_45674);
and UO_3739 (O_3739,N_45656,N_41711);
nor UO_3740 (O_3740,N_42135,N_42368);
nor UO_3741 (O_3741,N_40219,N_42689);
nand UO_3742 (O_3742,N_43270,N_47575);
nand UO_3743 (O_3743,N_40797,N_45966);
nor UO_3744 (O_3744,N_40630,N_49080);
nand UO_3745 (O_3745,N_40842,N_45211);
nand UO_3746 (O_3746,N_44040,N_47853);
nand UO_3747 (O_3747,N_46314,N_46664);
and UO_3748 (O_3748,N_41217,N_48648);
or UO_3749 (O_3749,N_44147,N_40440);
nand UO_3750 (O_3750,N_43402,N_43745);
or UO_3751 (O_3751,N_41340,N_48808);
and UO_3752 (O_3752,N_48198,N_48111);
xor UO_3753 (O_3753,N_49594,N_49709);
nand UO_3754 (O_3754,N_46134,N_48917);
xor UO_3755 (O_3755,N_46436,N_42726);
xor UO_3756 (O_3756,N_46937,N_42787);
xor UO_3757 (O_3757,N_40179,N_49032);
and UO_3758 (O_3758,N_46756,N_47896);
xor UO_3759 (O_3759,N_41284,N_44933);
nor UO_3760 (O_3760,N_42971,N_42955);
or UO_3761 (O_3761,N_47691,N_42748);
nand UO_3762 (O_3762,N_41161,N_43997);
nor UO_3763 (O_3763,N_42881,N_43098);
xnor UO_3764 (O_3764,N_49664,N_48135);
xnor UO_3765 (O_3765,N_46684,N_43009);
nand UO_3766 (O_3766,N_44066,N_40946);
or UO_3767 (O_3767,N_44330,N_45445);
or UO_3768 (O_3768,N_45562,N_49673);
and UO_3769 (O_3769,N_47024,N_44321);
or UO_3770 (O_3770,N_47660,N_45501);
nand UO_3771 (O_3771,N_44244,N_47274);
xor UO_3772 (O_3772,N_45655,N_47931);
nand UO_3773 (O_3773,N_40967,N_43776);
xor UO_3774 (O_3774,N_47728,N_46812);
nand UO_3775 (O_3775,N_44143,N_45861);
or UO_3776 (O_3776,N_43223,N_40038);
xnor UO_3777 (O_3777,N_42200,N_45280);
nand UO_3778 (O_3778,N_49977,N_41628);
xor UO_3779 (O_3779,N_45298,N_47526);
or UO_3780 (O_3780,N_47199,N_49141);
or UO_3781 (O_3781,N_45090,N_44422);
nand UO_3782 (O_3782,N_42504,N_41710);
and UO_3783 (O_3783,N_43027,N_40778);
nor UO_3784 (O_3784,N_40327,N_43130);
nand UO_3785 (O_3785,N_48069,N_44689);
or UO_3786 (O_3786,N_47093,N_42959);
nor UO_3787 (O_3787,N_41076,N_40799);
and UO_3788 (O_3788,N_41380,N_43889);
and UO_3789 (O_3789,N_47011,N_47765);
or UO_3790 (O_3790,N_41050,N_40910);
nor UO_3791 (O_3791,N_47672,N_43753);
nor UO_3792 (O_3792,N_49187,N_40061);
nand UO_3793 (O_3793,N_49053,N_49831);
and UO_3794 (O_3794,N_46574,N_47891);
nand UO_3795 (O_3795,N_48353,N_40785);
or UO_3796 (O_3796,N_42682,N_44663);
and UO_3797 (O_3797,N_48984,N_43281);
and UO_3798 (O_3798,N_47022,N_48586);
nand UO_3799 (O_3799,N_49998,N_44799);
nor UO_3800 (O_3800,N_40516,N_46735);
and UO_3801 (O_3801,N_42352,N_48134);
nor UO_3802 (O_3802,N_43490,N_44911);
or UO_3803 (O_3803,N_41121,N_47048);
xor UO_3804 (O_3804,N_48536,N_48171);
or UO_3805 (O_3805,N_43282,N_49380);
xor UO_3806 (O_3806,N_48022,N_45082);
xnor UO_3807 (O_3807,N_44569,N_47987);
xnor UO_3808 (O_3808,N_45630,N_42414);
and UO_3809 (O_3809,N_49295,N_46470);
xnor UO_3810 (O_3810,N_46739,N_46342);
and UO_3811 (O_3811,N_43160,N_46312);
nand UO_3812 (O_3812,N_42439,N_49904);
xor UO_3813 (O_3813,N_45727,N_43742);
and UO_3814 (O_3814,N_43741,N_47790);
xnor UO_3815 (O_3815,N_45676,N_44954);
nor UO_3816 (O_3816,N_47372,N_42700);
xnor UO_3817 (O_3817,N_45817,N_41308);
and UO_3818 (O_3818,N_47646,N_40023);
and UO_3819 (O_3819,N_40287,N_41559);
nor UO_3820 (O_3820,N_40892,N_44433);
nand UO_3821 (O_3821,N_47360,N_48300);
nor UO_3822 (O_3822,N_45954,N_45275);
or UO_3823 (O_3823,N_42175,N_48877);
or UO_3824 (O_3824,N_47502,N_46503);
xor UO_3825 (O_3825,N_48126,N_40566);
xor UO_3826 (O_3826,N_44119,N_47776);
nand UO_3827 (O_3827,N_43970,N_48631);
xnor UO_3828 (O_3828,N_45819,N_46910);
nand UO_3829 (O_3829,N_44912,N_40053);
and UO_3830 (O_3830,N_44594,N_41591);
and UO_3831 (O_3831,N_41782,N_44850);
or UO_3832 (O_3832,N_47821,N_44887);
and UO_3833 (O_3833,N_48834,N_48718);
or UO_3834 (O_3834,N_43553,N_42434);
or UO_3835 (O_3835,N_48912,N_43514);
and UO_3836 (O_3836,N_42608,N_47753);
or UO_3837 (O_3837,N_43791,N_48869);
nor UO_3838 (O_3838,N_48744,N_44192);
nand UO_3839 (O_3839,N_44839,N_40467);
nand UO_3840 (O_3840,N_44861,N_40188);
or UO_3841 (O_3841,N_44314,N_48804);
nor UO_3842 (O_3842,N_49746,N_49578);
and UO_3843 (O_3843,N_43056,N_49408);
or UO_3844 (O_3844,N_47941,N_44746);
and UO_3845 (O_3845,N_48147,N_40025);
nor UO_3846 (O_3846,N_49730,N_45906);
and UO_3847 (O_3847,N_40830,N_42899);
or UO_3848 (O_3848,N_41279,N_47468);
xor UO_3849 (O_3849,N_47904,N_46738);
or UO_3850 (O_3850,N_40740,N_42146);
and UO_3851 (O_3851,N_47550,N_41605);
nand UO_3852 (O_3852,N_42574,N_40469);
nor UO_3853 (O_3853,N_42929,N_44240);
or UO_3854 (O_3854,N_43386,N_49215);
or UO_3855 (O_3855,N_42909,N_40282);
nor UO_3856 (O_3856,N_44408,N_42257);
nand UO_3857 (O_3857,N_44631,N_46997);
xor UO_3858 (O_3858,N_47514,N_48932);
nor UO_3859 (O_3859,N_41357,N_44273);
or UO_3860 (O_3860,N_48066,N_49441);
or UO_3861 (O_3861,N_42948,N_48224);
nand UO_3862 (O_3862,N_48014,N_44926);
nand UO_3863 (O_3863,N_44229,N_40998);
nand UO_3864 (O_3864,N_45020,N_42300);
nand UO_3865 (O_3865,N_47659,N_45292);
nand UO_3866 (O_3866,N_42548,N_47619);
nand UO_3867 (O_3867,N_49154,N_44591);
nor UO_3868 (O_3868,N_49149,N_48715);
nor UO_3869 (O_3869,N_48070,N_42085);
xnor UO_3870 (O_3870,N_41679,N_41865);
nand UO_3871 (O_3871,N_43447,N_44345);
and UO_3872 (O_3872,N_46423,N_41527);
and UO_3873 (O_3873,N_40018,N_40974);
or UO_3874 (O_3874,N_47374,N_47808);
nor UO_3875 (O_3875,N_46331,N_48165);
xor UO_3876 (O_3876,N_40126,N_42653);
nand UO_3877 (O_3877,N_46001,N_46648);
nor UO_3878 (O_3878,N_43136,N_48866);
xor UO_3879 (O_3879,N_45712,N_42342);
nor UO_3880 (O_3880,N_41521,N_42177);
nand UO_3881 (O_3881,N_44669,N_41543);
nor UO_3882 (O_3882,N_47634,N_49641);
xnor UO_3883 (O_3883,N_48314,N_47735);
nor UO_3884 (O_3884,N_43985,N_48816);
and UO_3885 (O_3885,N_47465,N_41700);
or UO_3886 (O_3886,N_44306,N_42648);
or UO_3887 (O_3887,N_40532,N_44144);
or UO_3888 (O_3888,N_47561,N_44541);
nand UO_3889 (O_3889,N_45756,N_45046);
and UO_3890 (O_3890,N_45695,N_45902);
xor UO_3891 (O_3891,N_42117,N_46868);
nor UO_3892 (O_3892,N_41046,N_44064);
nor UO_3893 (O_3893,N_49205,N_46360);
nand UO_3894 (O_3894,N_43798,N_44374);
nand UO_3895 (O_3895,N_44820,N_41897);
or UO_3896 (O_3896,N_49834,N_48035);
and UO_3897 (O_3897,N_48110,N_48025);
nor UO_3898 (O_3898,N_47259,N_42760);
and UO_3899 (O_3899,N_40238,N_45346);
and UO_3900 (O_3900,N_47405,N_43227);
nor UO_3901 (O_3901,N_43600,N_49804);
or UO_3902 (O_3902,N_48130,N_46816);
or UO_3903 (O_3903,N_46949,N_40117);
nor UO_3904 (O_3904,N_41238,N_46535);
and UO_3905 (O_3905,N_48477,N_49092);
and UO_3906 (O_3906,N_48962,N_49658);
and UO_3907 (O_3907,N_47033,N_47233);
nor UO_3908 (O_3908,N_49336,N_46790);
nor UO_3909 (O_3909,N_47866,N_46195);
or UO_3910 (O_3910,N_44253,N_48491);
or UO_3911 (O_3911,N_43304,N_47466);
nor UO_3912 (O_3912,N_42650,N_46004);
nor UO_3913 (O_3913,N_45267,N_45531);
nand UO_3914 (O_3914,N_47351,N_42871);
nor UO_3915 (O_3915,N_41361,N_40142);
or UO_3916 (O_3916,N_46789,N_45387);
or UO_3917 (O_3917,N_42137,N_49196);
nand UO_3918 (O_3918,N_47521,N_44125);
xor UO_3919 (O_3919,N_41143,N_46234);
nor UO_3920 (O_3920,N_44415,N_41810);
nand UO_3921 (O_3921,N_42225,N_47650);
nand UO_3922 (O_3922,N_49868,N_46228);
xnor UO_3923 (O_3923,N_44759,N_43333);
and UO_3924 (O_3924,N_40152,N_43137);
and UO_3925 (O_3925,N_40573,N_40756);
or UO_3926 (O_3926,N_45661,N_40545);
or UO_3927 (O_3927,N_40819,N_41557);
xor UO_3928 (O_3928,N_40460,N_41854);
xor UO_3929 (O_3929,N_46274,N_40270);
nor UO_3930 (O_3930,N_48427,N_49306);
or UO_3931 (O_3931,N_46440,N_45662);
or UO_3932 (O_3932,N_42124,N_47140);
or UO_3933 (O_3933,N_49742,N_47134);
and UO_3934 (O_3934,N_41696,N_41266);
nand UO_3935 (O_3935,N_46068,N_48626);
and UO_3936 (O_3936,N_45247,N_42969);
nand UO_3937 (O_3937,N_42923,N_46215);
and UO_3938 (O_3938,N_44018,N_44885);
and UO_3939 (O_3939,N_49710,N_42828);
and UO_3940 (O_3940,N_40990,N_49407);
nand UO_3941 (O_3941,N_43943,N_40046);
nor UO_3942 (O_3942,N_44797,N_44449);
nor UO_3943 (O_3943,N_42133,N_48075);
nor UO_3944 (O_3944,N_40925,N_43388);
and UO_3945 (O_3945,N_49826,N_40608);
xnor UO_3946 (O_3946,N_49932,N_42488);
xnor UO_3947 (O_3947,N_48209,N_47926);
nand UO_3948 (O_3948,N_44877,N_47158);
nand UO_3949 (O_3949,N_45156,N_49139);
xnor UO_3950 (O_3950,N_43947,N_40299);
nand UO_3951 (O_3951,N_45074,N_41803);
nand UO_3952 (O_3952,N_44425,N_43878);
xor UO_3953 (O_3953,N_45793,N_46482);
nor UO_3954 (O_3954,N_40211,N_47180);
and UO_3955 (O_3955,N_44783,N_46747);
nor UO_3956 (O_3956,N_49317,N_48174);
or UO_3957 (O_3957,N_44934,N_42065);
nand UO_3958 (O_3958,N_49241,N_46913);
nand UO_3959 (O_3959,N_45161,N_41648);
xnor UO_3960 (O_3960,N_49161,N_49767);
nand UO_3961 (O_3961,N_48247,N_42518);
xnor UO_3962 (O_3962,N_49813,N_46278);
or UO_3963 (O_3963,N_49720,N_41789);
or UO_3964 (O_3964,N_48838,N_43065);
or UO_3965 (O_3965,N_42762,N_42722);
xnor UO_3966 (O_3966,N_47912,N_48584);
or UO_3967 (O_3967,N_49895,N_44207);
nor UO_3968 (O_3968,N_49933,N_48782);
or UO_3969 (O_3969,N_48301,N_41792);
nand UO_3970 (O_3970,N_41281,N_41011);
nor UO_3971 (O_3971,N_44976,N_40504);
and UO_3972 (O_3972,N_40745,N_41317);
and UO_3973 (O_3973,N_45476,N_41395);
xor UO_3974 (O_3974,N_45393,N_43844);
xnor UO_3975 (O_3975,N_45464,N_40264);
and UO_3976 (O_3976,N_45457,N_48141);
and UO_3977 (O_3977,N_41761,N_42381);
nand UO_3978 (O_3978,N_48878,N_41878);
or UO_3979 (O_3979,N_41270,N_42892);
or UO_3980 (O_3980,N_46296,N_42382);
xnor UO_3981 (O_3981,N_46387,N_47662);
or UO_3982 (O_3982,N_47651,N_43780);
or UO_3983 (O_3983,N_44388,N_42771);
and UO_3984 (O_3984,N_41285,N_44706);
and UO_3985 (O_3985,N_48725,N_49646);
nand UO_3986 (O_3986,N_48882,N_48389);
xor UO_3987 (O_3987,N_45997,N_48168);
xnor UO_3988 (O_3988,N_45159,N_44628);
xnor UO_3989 (O_3989,N_42576,N_42111);
or UO_3990 (O_3990,N_41875,N_43890);
or UO_3991 (O_3991,N_46353,N_47145);
nor UO_3992 (O_3992,N_40957,N_43201);
and UO_3993 (O_3993,N_42084,N_44152);
nor UO_3994 (O_3994,N_43584,N_46516);
or UO_3995 (O_3995,N_42094,N_47457);
xor UO_3996 (O_3996,N_49636,N_49305);
or UO_3997 (O_3997,N_49267,N_45228);
and UO_3998 (O_3998,N_42024,N_47007);
nand UO_3999 (O_3999,N_42636,N_47240);
and UO_4000 (O_4000,N_49743,N_41621);
or UO_4001 (O_4001,N_46435,N_40623);
xor UO_4002 (O_4002,N_44342,N_47352);
nor UO_4003 (O_4003,N_46867,N_45026);
and UO_4004 (O_4004,N_49044,N_41755);
nand UO_4005 (O_4005,N_43498,N_40520);
or UO_4006 (O_4006,N_40438,N_48377);
nor UO_4007 (O_4007,N_41545,N_46217);
or UO_4008 (O_4008,N_46520,N_45359);
nor UO_4009 (O_4009,N_47413,N_45165);
nand UO_4010 (O_4010,N_41086,N_43914);
nand UO_4011 (O_4011,N_41396,N_48434);
xor UO_4012 (O_4012,N_42918,N_40301);
xor UO_4013 (O_4013,N_49188,N_49443);
and UO_4014 (O_4014,N_49622,N_48446);
nor UO_4015 (O_4015,N_48801,N_41278);
or UO_4016 (O_4016,N_45055,N_44967);
or UO_4017 (O_4017,N_48223,N_49698);
nor UO_4018 (O_4018,N_45876,N_45946);
and UO_4019 (O_4019,N_45001,N_46815);
and UO_4020 (O_4020,N_42433,N_44130);
xor UO_4021 (O_4021,N_43724,N_41324);
nor UO_4022 (O_4022,N_40689,N_49327);
or UO_4023 (O_4023,N_45737,N_41662);
xnor UO_4024 (O_4024,N_43342,N_47041);
nand UO_4025 (O_4025,N_43299,N_45041);
and UO_4026 (O_4026,N_47389,N_41014);
and UO_4027 (O_4027,N_42662,N_40308);
xnor UO_4028 (O_4028,N_42860,N_44802);
and UO_4029 (O_4029,N_41329,N_41136);
and UO_4030 (O_4030,N_40131,N_42547);
or UO_4031 (O_4031,N_46674,N_45120);
nand UO_4032 (O_4032,N_41377,N_43491);
or UO_4033 (O_4033,N_48065,N_46964);
and UO_4034 (O_4034,N_49113,N_47880);
and UO_4035 (O_4035,N_42139,N_46458);
nor UO_4036 (O_4036,N_40399,N_49722);
nor UO_4037 (O_4037,N_47594,N_47324);
xnor UO_4038 (O_4038,N_43382,N_49490);
xor UO_4039 (O_4039,N_44378,N_45276);
nand UO_4040 (O_4040,N_46783,N_43501);
nor UO_4041 (O_4041,N_41177,N_43916);
and UO_4042 (O_4042,N_42500,N_42450);
and UO_4043 (O_4043,N_40039,N_45851);
nand UO_4044 (O_4044,N_42593,N_46791);
nand UO_4045 (O_4045,N_49015,N_44742);
nand UO_4046 (O_4046,N_40232,N_45767);
nand UO_4047 (O_4047,N_43846,N_44495);
nand UO_4048 (O_4048,N_49308,N_49193);
nor UO_4049 (O_4049,N_42374,N_49423);
nor UO_4050 (O_4050,N_46221,N_49962);
and UO_4051 (O_4051,N_45083,N_41624);
nand UO_4052 (O_4052,N_42425,N_40699);
or UO_4053 (O_4053,N_44311,N_44262);
xnor UO_4054 (O_4054,N_44924,N_43751);
nor UO_4055 (O_4055,N_45091,N_45901);
xor UO_4056 (O_4056,N_43628,N_43805);
nand UO_4057 (O_4057,N_46028,N_48298);
and UO_4058 (O_4058,N_46046,N_42079);
nand UO_4059 (O_4059,N_43175,N_49303);
nand UO_4060 (O_4060,N_49901,N_45422);
or UO_4061 (O_4061,N_43690,N_48109);
or UO_4062 (O_4062,N_43470,N_48577);
xor UO_4063 (O_4063,N_49886,N_46306);
xnor UO_4064 (O_4064,N_44930,N_41587);
and UO_4065 (O_4065,N_44698,N_48798);
nand UO_4066 (O_4066,N_49574,N_42829);
or UO_4067 (O_4067,N_46948,N_45527);
xor UO_4068 (O_4068,N_44557,N_46978);
xnor UO_4069 (O_4069,N_41132,N_40825);
nand UO_4070 (O_4070,N_40470,N_44348);
or UO_4071 (O_4071,N_48841,N_49881);
xor UO_4072 (O_4072,N_48666,N_42563);
nor UO_4073 (O_4073,N_42239,N_43992);
xnor UO_4074 (O_4074,N_41631,N_47018);
nor UO_4075 (O_4075,N_49321,N_45951);
or UO_4076 (O_4076,N_40933,N_40801);
xnor UO_4077 (O_4077,N_46156,N_46206);
nor UO_4078 (O_4078,N_41937,N_46595);
or UO_4079 (O_4079,N_46980,N_49021);
or UO_4080 (O_4080,N_46178,N_46614);
and UO_4081 (O_4081,N_41115,N_43446);
and UO_4082 (O_4082,N_49967,N_45605);
or UO_4083 (O_4083,N_49867,N_46874);
xor UO_4084 (O_4084,N_47581,N_48253);
nand UO_4085 (O_4085,N_41987,N_42927);
xor UO_4086 (O_4086,N_44120,N_47106);
nor UO_4087 (O_4087,N_49719,N_47603);
nand UO_4088 (O_4088,N_40233,N_45787);
xor UO_4089 (O_4089,N_41411,N_48442);
and UO_4090 (O_4090,N_43730,N_47605);
nand UO_4091 (O_4091,N_40074,N_46269);
xor UO_4092 (O_4092,N_40521,N_46656);
and UO_4093 (O_4093,N_46270,N_44851);
xor UO_4094 (O_4094,N_43531,N_41504);
xor UO_4095 (O_4095,N_43347,N_42050);
xnor UO_4096 (O_4096,N_47347,N_49669);
and UO_4097 (O_4097,N_49944,N_43169);
nor UO_4098 (O_4098,N_45255,N_48164);
nand UO_4099 (O_4099,N_46181,N_47212);
or UO_4100 (O_4100,N_41509,N_41032);
or UO_4101 (O_4101,N_45537,N_46942);
nand UO_4102 (O_4102,N_47725,N_45190);
or UO_4103 (O_4103,N_49016,N_48037);
xnor UO_4104 (O_4104,N_49233,N_49836);
or UO_4105 (O_4105,N_43370,N_40120);
nand UO_4106 (O_4106,N_49244,N_48067);
nor UO_4107 (O_4107,N_41446,N_48946);
nor UO_4108 (O_4108,N_42093,N_49503);
nand UO_4109 (O_4109,N_47504,N_43522);
nor UO_4110 (O_4110,N_44367,N_43838);
nor UO_4111 (O_4111,N_45964,N_45894);
xnor UO_4112 (O_4112,N_45582,N_46351);
nor UO_4113 (O_4113,N_44111,N_45781);
nand UO_4114 (O_4114,N_49040,N_44186);
and UO_4115 (O_4115,N_49146,N_42271);
nand UO_4116 (O_4116,N_44351,N_41833);
and UO_4117 (O_4117,N_49628,N_47489);
nor UO_4118 (O_4118,N_40030,N_41692);
xor UO_4119 (O_4119,N_44875,N_45149);
and UO_4120 (O_4120,N_41535,N_47622);
nand UO_4121 (O_4121,N_46862,N_43073);
xnor UO_4122 (O_4122,N_43718,N_46488);
xor UO_4123 (O_4123,N_48783,N_46393);
xnor UO_4124 (O_4124,N_44729,N_40594);
nor UO_4125 (O_4125,N_48609,N_48572);
nor UO_4126 (O_4126,N_42078,N_49039);
or UO_4127 (O_4127,N_41160,N_41630);
or UO_4128 (O_4128,N_48337,N_45980);
and UO_4129 (O_4129,N_41618,N_41181);
or UO_4130 (O_4130,N_48019,N_46136);
nand UO_4131 (O_4131,N_48897,N_48020);
nor UO_4132 (O_4132,N_40361,N_40058);
or UO_4133 (O_4133,N_47325,N_47426);
nand UO_4134 (O_4134,N_43641,N_47395);
or UO_4135 (O_4135,N_41954,N_42599);
or UO_4136 (O_4136,N_43713,N_42939);
nand UO_4137 (O_4137,N_46947,N_47097);
and UO_4138 (O_4138,N_45765,N_48862);
and UO_4139 (O_4139,N_45439,N_49312);
xor UO_4140 (O_4140,N_43942,N_40332);
and UO_4141 (O_4141,N_42004,N_41409);
nor UO_4142 (O_4142,N_41822,N_49123);
nand UO_4143 (O_4143,N_48636,N_48456);
and UO_4144 (O_4144,N_41139,N_46943);
nor UO_4145 (O_4145,N_46054,N_46507);
xor UO_4146 (O_4146,N_46396,N_44810);
or UO_4147 (O_4147,N_49077,N_46433);
xnor UO_4148 (O_4148,N_44350,N_41768);
nand UO_4149 (O_4149,N_49276,N_41958);
or UO_4150 (O_4150,N_41612,N_46256);
and UO_4151 (O_4151,N_43318,N_46734);
nor UO_4152 (O_4152,N_40599,N_47584);
nand UO_4153 (O_4153,N_40875,N_43863);
nand UO_4154 (O_4154,N_48354,N_48447);
nand UO_4155 (O_4155,N_42867,N_48791);
or UO_4156 (O_4156,N_44805,N_42158);
xor UO_4157 (O_4157,N_46728,N_49570);
nor UO_4158 (O_4158,N_41141,N_41468);
or UO_4159 (O_4159,N_43409,N_47760);
or UO_4160 (O_4160,N_40530,N_41250);
and UO_4161 (O_4161,N_46192,N_41245);
nor UO_4162 (O_4162,N_45804,N_42559);
xor UO_4163 (O_4163,N_49459,N_48218);
or UO_4164 (O_4164,N_43037,N_46179);
nand UO_4165 (O_4165,N_46148,N_43521);
nand UO_4166 (O_4166,N_49076,N_41301);
xor UO_4167 (O_4167,N_41570,N_41745);
and UO_4168 (O_4168,N_43989,N_48423);
xnor UO_4169 (O_4169,N_40011,N_42993);
and UO_4170 (O_4170,N_43649,N_48261);
or UO_4171 (O_4171,N_42898,N_40847);
nor UO_4172 (O_4172,N_46966,N_44384);
nor UO_4173 (O_4173,N_40989,N_40037);
xnor UO_4174 (O_4174,N_49993,N_46932);
or UO_4175 (O_4175,N_46216,N_49243);
xnor UO_4176 (O_4176,N_48544,N_46627);
nor UO_4177 (O_4177,N_44496,N_40904);
or UO_4178 (O_4178,N_46857,N_40073);
and UO_4179 (O_4179,N_41608,N_47120);
or UO_4180 (O_4180,N_42893,N_42141);
or UO_4181 (O_4181,N_41642,N_44917);
nor UO_4182 (O_4182,N_43199,N_40280);
and UO_4183 (O_4183,N_40813,N_40336);
or UO_4184 (O_4184,N_48824,N_40941);
xnor UO_4185 (O_4185,N_43263,N_41620);
nand UO_4186 (O_4186,N_44597,N_47161);
and UO_4187 (O_4187,N_45682,N_44290);
nand UO_4188 (O_4188,N_42681,N_44476);
and UO_4189 (O_4189,N_41044,N_45824);
nor UO_4190 (O_4190,N_41765,N_47831);
nor UO_4191 (O_4191,N_47608,N_44296);
nand UO_4192 (O_4192,N_41215,N_46142);
and UO_4193 (O_4193,N_41318,N_45904);
nor UO_4194 (O_4194,N_40261,N_43437);
and UO_4195 (O_4195,N_42273,N_44580);
or UO_4196 (O_4196,N_40883,N_47016);
or UO_4197 (O_4197,N_49186,N_48589);
nor UO_4198 (O_4198,N_47569,N_47409);
xor UO_4199 (O_4199,N_41255,N_45733);
xnor UO_4200 (O_4200,N_42138,N_40585);
nand UO_4201 (O_4201,N_46641,N_46847);
or UO_4202 (O_4202,N_47488,N_46294);
or UO_4203 (O_4203,N_46575,N_40555);
or UO_4204 (O_4204,N_46890,N_46527);
and UO_4205 (O_4205,N_48362,N_43108);
nand UO_4206 (O_4206,N_45521,N_45705);
nor UO_4207 (O_4207,N_43415,N_47837);
or UO_4208 (O_4208,N_40317,N_41339);
or UO_4209 (O_4209,N_49487,N_48264);
xor UO_4210 (O_4210,N_42587,N_44517);
or UO_4211 (O_4211,N_45430,N_48230);
and UO_4212 (O_4212,N_40647,N_45344);
or UO_4213 (O_4213,N_41622,N_42818);
nand UO_4214 (O_4214,N_48759,N_40303);
xor UO_4215 (O_4215,N_41083,N_40384);
nor UO_4216 (O_4216,N_43159,N_45821);
or UO_4217 (O_4217,N_43939,N_43558);
nor UO_4218 (O_4218,N_42056,N_44677);
and UO_4219 (O_4219,N_43897,N_46990);
xnor UO_4220 (O_4220,N_46896,N_42619);
nand UO_4221 (O_4221,N_41381,N_40450);
nand UO_4222 (O_4222,N_41726,N_49447);
nand UO_4223 (O_4223,N_47712,N_45103);
or UO_4224 (O_4224,N_42044,N_42267);
nand UO_4225 (O_4225,N_47424,N_48106);
nor UO_4226 (O_4226,N_41835,N_43326);
and UO_4227 (O_4227,N_41359,N_44902);
and UO_4228 (O_4228,N_41020,N_44955);
nand UO_4229 (O_4229,N_41767,N_43933);
or UO_4230 (O_4230,N_45392,N_47197);
or UO_4231 (O_4231,N_49788,N_41814);
nor UO_4232 (O_4232,N_44091,N_40816);
and UO_4233 (O_4233,N_48076,N_43417);
or UO_4234 (O_4234,N_49631,N_45148);
xor UO_4235 (O_4235,N_47554,N_48058);
nor UO_4236 (O_4236,N_40116,N_42704);
xnor UO_4237 (O_4237,N_48281,N_48713);
xnor UO_4238 (O_4238,N_41590,N_43831);
and UO_4239 (O_4239,N_40487,N_43395);
xor UO_4240 (O_4240,N_40146,N_43761);
nor UO_4241 (O_4241,N_47486,N_40831);
and UO_4242 (O_4242,N_43560,N_49491);
nor UO_4243 (O_4243,N_42171,N_46694);
and UO_4244 (O_4244,N_43450,N_48563);
nand UO_4245 (O_4245,N_44227,N_48794);
and UO_4246 (O_4246,N_48155,N_49331);
nor UO_4247 (O_4247,N_40942,N_47532);
nand UO_4248 (O_4248,N_42073,N_49782);
and UO_4249 (O_4249,N_41571,N_48593);
nor UO_4250 (O_4250,N_46637,N_40738);
xor UO_4251 (O_4251,N_45245,N_47366);
and UO_4252 (O_4252,N_42363,N_44499);
and UO_4253 (O_4253,N_41055,N_44886);
nand UO_4254 (O_4254,N_48723,N_46979);
or UO_4255 (O_4255,N_40635,N_42080);
nor UO_4256 (O_4256,N_42880,N_43140);
or UO_4257 (O_4257,N_42883,N_40182);
nor UO_4258 (O_4258,N_44438,N_49171);
nor UO_4259 (O_4259,N_43571,N_45173);
nand UO_4260 (O_4260,N_46646,N_41122);
nand UO_4261 (O_4261,N_46441,N_41977);
nand UO_4262 (O_4262,N_48484,N_44479);
nor UO_4263 (O_4263,N_40653,N_46557);
and UO_4264 (O_4264,N_49483,N_46513);
and UO_4265 (O_4265,N_49997,N_43239);
xnor UO_4266 (O_4266,N_44826,N_41531);
or UO_4267 (O_4267,N_48502,N_44910);
nor UO_4268 (O_4268,N_46127,N_40048);
nor UO_4269 (O_4269,N_48341,N_41821);
nand UO_4270 (O_4270,N_48894,N_46546);
nor UO_4271 (O_4271,N_49147,N_48943);
and UO_4272 (O_4272,N_42366,N_41708);
xor UO_4273 (O_4273,N_42331,N_44126);
nor UO_4274 (O_4274,N_42837,N_42469);
or UO_4275 (O_4275,N_40648,N_41392);
nor UO_4276 (O_4276,N_43245,N_46689);
nand UO_4277 (O_4277,N_45295,N_40352);
or UO_4278 (O_4278,N_43801,N_40829);
xnor UO_4279 (O_4279,N_41843,N_46416);
nor UO_4280 (O_4280,N_44959,N_46097);
nand UO_4281 (O_4281,N_43660,N_41793);
nand UO_4282 (O_4282,N_45349,N_41024);
xor UO_4283 (O_4283,N_43147,N_49840);
xnor UO_4284 (O_4284,N_42875,N_41674);
nand UO_4285 (O_4285,N_48857,N_45473);
nor UO_4286 (O_4286,N_41442,N_44801);
or UO_4287 (O_4287,N_48842,N_44581);
and UO_4288 (O_4288,N_45152,N_44881);
nor UO_4289 (O_4289,N_43045,N_47334);
and UO_4290 (O_4290,N_40882,N_42654);
and UO_4291 (O_4291,N_48274,N_48330);
nor UO_4292 (O_4292,N_43663,N_41328);
nand UO_4293 (O_4293,N_43729,N_44326);
nor UO_4294 (O_4294,N_41638,N_41689);
and UO_4295 (O_4295,N_40476,N_44317);
or UO_4296 (O_4296,N_41183,N_45413);
nor UO_4297 (O_4297,N_45254,N_40325);
or UO_4298 (O_4298,N_41081,N_40226);
and UO_4299 (O_4299,N_48291,N_46751);
nand UO_4300 (O_4300,N_48358,N_47540);
xnor UO_4301 (O_4301,N_49623,N_48797);
xnor UO_4302 (O_4302,N_48964,N_46876);
or UO_4303 (O_4303,N_43421,N_40769);
xor UO_4304 (O_4304,N_41926,N_47232);
and UO_4305 (O_4305,N_40346,N_44209);
and UO_4306 (O_4306,N_40056,N_41911);
nor UO_4307 (O_4307,N_40869,N_48881);
or UO_4308 (O_4308,N_45330,N_44247);
or UO_4309 (O_4309,N_48023,N_47962);
and UO_4310 (O_4310,N_41125,N_48766);
xor UO_4311 (O_4311,N_44822,N_47513);
nor UO_4312 (O_4312,N_40166,N_45933);
and UO_4313 (O_4313,N_41458,N_47589);
and UO_4314 (O_4314,N_40175,N_43276);
nand UO_4315 (O_4315,N_42568,N_40349);
and UO_4316 (O_4316,N_44781,N_47275);
and UO_4317 (O_4317,N_48499,N_40928);
nand UO_4318 (O_4318,N_42772,N_46450);
xnor UO_4319 (O_4319,N_49192,N_46271);
xnor UO_4320 (O_4320,N_48690,N_42745);
and UO_4321 (O_4321,N_44423,N_44228);
or UO_4322 (O_4322,N_40781,N_41558);
or UO_4323 (O_4323,N_41043,N_49325);
or UO_4324 (O_4324,N_41154,N_49111);
nor UO_4325 (O_4325,N_48674,N_44459);
or UO_4326 (O_4326,N_49227,N_47412);
xor UO_4327 (O_4327,N_44201,N_41750);
xnor UO_4328 (O_4328,N_44249,N_46829);
or UO_4329 (O_4329,N_42820,N_46143);
and UO_4330 (O_4330,N_46834,N_41342);
or UO_4331 (O_4331,N_49083,N_47933);
nor UO_4332 (O_4332,N_41942,N_49436);
nand UO_4333 (O_4333,N_40033,N_45638);
nor UO_4334 (O_4334,N_45718,N_40390);
or UO_4335 (O_4335,N_45595,N_48436);
nor UO_4336 (O_4336,N_43295,N_48973);
nor UO_4337 (O_4337,N_43790,N_45871);
xnor UO_4338 (O_4338,N_49586,N_45986);
and UO_4339 (O_4339,N_49018,N_45278);
xor UO_4340 (O_4340,N_48204,N_48195);
or UO_4341 (O_4341,N_46079,N_48459);
nand UO_4342 (O_4342,N_40227,N_40682);
or UO_4343 (O_4343,N_41758,N_42114);
xnor UO_4344 (O_4344,N_42519,N_43909);
xor UO_4345 (O_4345,N_40425,N_44081);
nor UO_4346 (O_4346,N_46265,N_44928);
nor UO_4347 (O_4347,N_40535,N_40934);
nor UO_4348 (O_4348,N_46903,N_45840);
nand UO_4349 (O_4349,N_44626,N_48968);
nand UO_4350 (O_4350,N_47296,N_46704);
xnor UO_4351 (O_4351,N_47040,N_47991);
or UO_4352 (O_4352,N_46599,N_49229);
nand UO_4353 (O_4353,N_41333,N_47748);
and UO_4354 (O_4354,N_44687,N_45384);
or UO_4355 (O_4355,N_47133,N_40675);
xor UO_4356 (O_4356,N_42687,N_40357);
nor UO_4357 (O_4357,N_41444,N_47035);
nor UO_4358 (O_4358,N_45751,N_48683);
nor UO_4359 (O_4359,N_48604,N_49159);
nand UO_4360 (O_4360,N_49558,N_48909);
or UO_4361 (O_4361,N_47036,N_46662);
and UO_4362 (O_4362,N_43930,N_41465);
and UO_4363 (O_4363,N_42214,N_47788);
nand UO_4364 (O_4364,N_48345,N_47139);
and UO_4365 (O_4365,N_47782,N_45224);
and UO_4366 (O_4366,N_44763,N_41502);
nor UO_4367 (O_4367,N_49495,N_46013);
or UO_4368 (O_4368,N_44177,N_48886);
or UO_4369 (O_4369,N_46469,N_44538);
or UO_4370 (O_4370,N_42591,N_40960);
or UO_4371 (O_4371,N_43623,N_49444);
nand UO_4372 (O_4372,N_40035,N_49042);
or UO_4373 (O_4373,N_44432,N_45297);
nor UO_4374 (O_4374,N_44710,N_43464);
xnor UO_4375 (O_4375,N_40839,N_44670);
nand UO_4376 (O_4376,N_44360,N_48348);
or UO_4377 (O_4377,N_45398,N_40164);
xnor UO_4378 (O_4378,N_46255,N_46792);
and UO_4379 (O_4379,N_49701,N_44823);
and UO_4380 (O_4380,N_47859,N_44464);
or UO_4381 (O_4381,N_41493,N_41560);
nand UO_4382 (O_4382,N_49120,N_47150);
nor UO_4383 (O_4383,N_43268,N_47860);
nand UO_4384 (O_4384,N_49377,N_42372);
or UO_4385 (O_4385,N_47260,N_45845);
xor UO_4386 (O_4386,N_45975,N_48118);
xor UO_4387 (O_4387,N_43383,N_40463);
nor UO_4388 (O_4388,N_48433,N_48176);
or UO_4389 (O_4389,N_45517,N_45481);
xor UO_4390 (O_4390,N_47249,N_43694);
nor UO_4391 (O_4391,N_48257,N_45277);
nor UO_4392 (O_4392,N_42058,N_47963);
nand UO_4393 (O_4393,N_40374,N_48200);
nor UO_4394 (O_4394,N_43708,N_48889);
nor UO_4395 (O_4395,N_49857,N_43458);
and UO_4396 (O_4396,N_41754,N_46526);
and UO_4397 (O_4397,N_42876,N_45348);
nor UO_4398 (O_4398,N_46103,N_40492);
nor UO_4399 (O_4399,N_41625,N_42750);
xor UO_4400 (O_4400,N_49949,N_48708);
xor UO_4401 (O_4401,N_45180,N_48121);
or UO_4402 (O_4402,N_44443,N_45350);
nor UO_4403 (O_4403,N_44562,N_45541);
and UO_4404 (O_4404,N_46344,N_49955);
or UO_4405 (O_4405,N_46733,N_45311);
nor UO_4406 (O_4406,N_40132,N_41330);
xor UO_4407 (O_4407,N_46006,N_46359);
nand UO_4408 (O_4408,N_42814,N_42514);
and UO_4409 (O_4409,N_43072,N_44169);
and UO_4410 (O_4410,N_49642,N_48625);
xor UO_4411 (O_4411,N_44691,N_46020);
nand UO_4412 (O_4412,N_43047,N_46691);
nand UO_4413 (O_4413,N_49426,N_42905);
or UO_4414 (O_4414,N_47911,N_48995);
and UO_4415 (O_4415,N_41106,N_48989);
or UO_4416 (O_4416,N_46703,N_41838);
nand UO_4417 (O_4417,N_47151,N_42845);
xor UO_4418 (O_4418,N_48371,N_48245);
or UO_4419 (O_4419,N_45624,N_45479);
or UO_4420 (O_4420,N_42592,N_49983);
and UO_4421 (O_4421,N_41596,N_48248);
and UO_4422 (O_4422,N_43255,N_46623);
nand UO_4423 (O_4423,N_41986,N_41174);
or UO_4424 (O_4424,N_46045,N_49057);
and UO_4425 (O_4425,N_45632,N_43685);
xnor UO_4426 (O_4426,N_44749,N_41652);
and UO_4427 (O_4427,N_45800,N_42761);
nand UO_4428 (O_4428,N_40136,N_47525);
xnor UO_4429 (O_4429,N_46536,N_41589);
or UO_4430 (O_4430,N_47950,N_41617);
nor UO_4431 (O_4431,N_46146,N_41091);
and UO_4432 (O_4432,N_42294,N_42391);
and UO_4433 (O_4433,N_42698,N_48652);
or UO_4434 (O_4434,N_44493,N_43732);
nand UO_4435 (O_4435,N_40522,N_45383);
or UO_4436 (O_4436,N_44555,N_44022);
and UO_4437 (O_4437,N_43851,N_47121);
xnor UO_4438 (O_4438,N_40704,N_48157);
xnor UO_4439 (O_4439,N_41224,N_42010);
and UO_4440 (O_4440,N_46324,N_40603);
and UO_4441 (O_4441,N_46824,N_44889);
and UO_4442 (O_4442,N_46483,N_40321);
and UO_4443 (O_4443,N_46588,N_48100);
or UO_4444 (O_4444,N_42097,N_43736);
xnor UO_4445 (O_4445,N_42495,N_42631);
nor UO_4446 (O_4446,N_42211,N_44176);
nand UO_4447 (O_4447,N_49812,N_41779);
nand UO_4448 (O_4448,N_47479,N_47236);
xor UO_4449 (O_4449,N_42092,N_42428);
or UO_4450 (O_4450,N_46584,N_47364);
nand UO_4451 (O_4451,N_44319,N_45369);
nor UO_4452 (O_4452,N_47836,N_48960);
xnor UO_4453 (O_4453,N_44371,N_47980);
or UO_4454 (O_4454,N_46901,N_40178);
or UO_4455 (O_4455,N_48249,N_43093);
xor UO_4456 (O_4456,N_48036,N_43563);
and UO_4457 (O_4457,N_43517,N_49043);
nor UO_4458 (O_4458,N_46322,N_49318);
and UO_4459 (O_4459,N_43104,N_43021);
xnor UO_4460 (O_4460,N_45973,N_41828);
xnor UO_4461 (O_4461,N_42705,N_40502);
xor UO_4462 (O_4462,N_46786,N_40176);
and UO_4463 (O_4463,N_44129,N_45123);
and UO_4464 (O_4464,N_43710,N_49045);
or UO_4465 (O_4465,N_44076,N_43870);
or UO_4466 (O_4466,N_49681,N_44254);
xnor UO_4467 (O_4467,N_44898,N_43361);
nand UO_4468 (O_4468,N_45750,N_49609);
or UO_4469 (O_4469,N_45483,N_47542);
xnor UO_4470 (O_4470,N_49815,N_45903);
or UO_4471 (O_4471,N_41335,N_49086);
nand UO_4472 (O_4472,N_48207,N_42472);
or UO_4473 (O_4473,N_41858,N_40529);
or UO_4474 (O_4474,N_40105,N_42679);
or UO_4475 (O_4475,N_40633,N_44754);
xor UO_4476 (O_4476,N_45826,N_43141);
nor UO_4477 (O_4477,N_40129,N_46063);
nor UO_4478 (O_4478,N_47863,N_47382);
nand UO_4479 (O_4479,N_48183,N_47562);
and UO_4480 (O_4480,N_45293,N_45852);
or UO_4481 (O_4481,N_44041,N_49935);
or UO_4482 (O_4482,N_40429,N_48144);
nor UO_4483 (O_4483,N_43578,N_41781);
nor UO_4484 (O_4484,N_44836,N_40606);
and UO_4485 (O_4485,N_43366,N_43472);
and UO_4486 (O_4486,N_46023,N_47012);
nor UO_4487 (O_4487,N_45230,N_40548);
and UO_4488 (O_4488,N_46752,N_45620);
xnor UO_4489 (O_4489,N_42468,N_45769);
nand UO_4490 (O_4490,N_47843,N_49082);
nand UO_4491 (O_4491,N_49068,N_46210);
nor UO_4492 (O_4492,N_40834,N_46745);
nor UO_4493 (O_4493,N_40674,N_47849);
and UO_4494 (O_4494,N_41077,N_41871);
and UO_4495 (O_4495,N_41180,N_40976);
and UO_4496 (O_4496,N_46025,N_43922);
nand UO_4497 (O_4497,N_45953,N_47677);
or UO_4498 (O_4498,N_46095,N_41486);
xnor UO_4499 (O_4499,N_43564,N_43119);
nand UO_4500 (O_4500,N_40065,N_45356);
or UO_4501 (O_4501,N_49688,N_40562);
and UO_4502 (O_4502,N_40414,N_40419);
xnor UO_4503 (O_4503,N_48654,N_49841);
or UO_4504 (O_4504,N_47638,N_47288);
or UO_4505 (O_4505,N_41005,N_44860);
or UO_4506 (O_4506,N_49500,N_40031);
and UO_4507 (O_4507,N_47596,N_43121);
xnor UO_4508 (O_4508,N_47770,N_41483);
or UO_4509 (O_4509,N_47501,N_45702);
nor UO_4510 (O_4510,N_40567,N_48904);
or UO_4511 (O_4511,N_42711,N_48746);
xnor UO_4512 (O_4512,N_43489,N_46432);
xnor UO_4513 (O_4513,N_41390,N_48219);
and UO_4514 (O_4514,N_47998,N_48981);
nand UO_4515 (O_4515,N_41368,N_41216);
and UO_4516 (O_4516,N_48706,N_47938);
or UO_4517 (O_4517,N_46564,N_46533);
nor UO_4518 (O_4518,N_44588,N_42664);
nand UO_4519 (O_4519,N_49002,N_48344);
or UO_4520 (O_4520,N_48977,N_41722);
nor UO_4521 (O_4521,N_46705,N_42537);
nor UO_4522 (O_4522,N_44545,N_49755);
or UO_4523 (O_4523,N_40140,N_46490);
and UO_4524 (O_4524,N_43495,N_41895);
and UO_4525 (O_4525,N_40540,N_44623);
and UO_4526 (O_4526,N_40531,N_46884);
and UO_4527 (O_4527,N_47256,N_40202);
nor UO_4528 (O_4528,N_43187,N_49218);
and UO_4529 (O_4529,N_47764,N_45167);
nor UO_4530 (O_4530,N_40356,N_45188);
or UO_4531 (O_4531,N_40124,N_49885);
nand UO_4532 (O_4532,N_44069,N_43769);
and UO_4533 (O_4533,N_42234,N_46137);
nor UO_4534 (O_4534,N_45589,N_46530);
nor UO_4535 (O_4535,N_41169,N_49802);
nor UO_4536 (O_4536,N_47020,N_40488);
and UO_4537 (O_4537,N_43807,N_43706);
nor UO_4538 (O_4538,N_44335,N_44940);
or UO_4539 (O_4539,N_43067,N_49257);
nand UO_4540 (O_4540,N_43350,N_41094);
xor UO_4541 (O_4541,N_46800,N_49326);
nor UO_4542 (O_4542,N_43234,N_42852);
and UO_4543 (O_4543,N_42014,N_45757);
xnor UO_4544 (O_4544,N_43859,N_45506);
or UO_4545 (O_4545,N_46414,N_46744);
and UO_4546 (O_4546,N_45841,N_46761);
and UO_4547 (O_4547,N_45203,N_41566);
or UO_4548 (O_4548,N_46456,N_46188);
nand UO_4549 (O_4549,N_46668,N_42953);
xnor UO_4550 (O_4550,N_47293,N_43612);
nand UO_4551 (O_4551,N_46576,N_42950);
xor UO_4552 (O_4552,N_43219,N_42249);
nand UO_4553 (O_4553,N_43505,N_46319);
nor UO_4554 (O_4554,N_44313,N_48660);
and UO_4555 (O_4555,N_48902,N_43869);
or UO_4556 (O_4556,N_45614,N_40986);
nor UO_4557 (O_4557,N_47432,N_44617);
xor UO_4558 (O_4558,N_40652,N_40667);
nor UO_4559 (O_4559,N_45771,N_44527);
xnor UO_4560 (O_4560,N_41336,N_43430);
nor UO_4561 (O_4561,N_45745,N_40337);
and UO_4562 (O_4562,N_47164,N_43097);
and UO_4563 (O_4563,N_49298,N_43334);
xnor UO_4564 (O_4564,N_44393,N_47219);
or UO_4565 (O_4565,N_48867,N_48854);
nor UO_4566 (O_4566,N_43891,N_45825);
xor UO_4567 (O_4567,N_47729,N_46289);
nor UO_4568 (O_4568,N_49775,N_41802);
xor UO_4569 (O_4569,N_44651,N_42181);
xnor UO_4570 (O_4570,N_45493,N_44336);
nor UO_4571 (O_4571,N_45523,N_42051);
nor UO_4572 (O_4572,N_47283,N_48062);
nand UO_4573 (O_4573,N_43378,N_49037);
nand UO_4574 (O_4574,N_44680,N_48731);
nand UO_4575 (O_4575,N_43305,N_42861);
nor UO_4576 (O_4576,N_48246,N_42332);
or UO_4577 (O_4577,N_47737,N_40275);
and UO_4578 (O_4578,N_44765,N_43026);
xor UO_4579 (O_4579,N_44962,N_40907);
nor UO_4580 (O_4580,N_44720,N_40927);
xnor UO_4581 (O_4581,N_46491,N_49614);
nand UO_4582 (O_4582,N_49889,N_49640);
xnor UO_4583 (O_4583,N_46532,N_41349);
xor UO_4584 (O_4584,N_42317,N_49524);
and UO_4585 (O_4585,N_45281,N_41277);
or UO_4586 (O_4586,N_43408,N_42725);
or UO_4587 (O_4587,N_41695,N_47222);
nand UO_4588 (O_4588,N_48284,N_43768);
nand UO_4589 (O_4589,N_40394,N_42637);
nand UO_4590 (O_4590,N_44255,N_44239);
nor UO_4591 (O_4591,N_43669,N_47674);
and UO_4592 (O_4592,N_45418,N_40864);
nand UO_4593 (O_4593,N_40088,N_40800);
and UO_4594 (O_4594,N_43682,N_48545);
or UO_4595 (O_4595,N_46437,N_46587);
and UO_4596 (O_4596,N_46920,N_44068);
nand UO_4597 (O_4597,N_40377,N_44867);
and UO_4598 (O_4598,N_44398,N_40891);
xor UO_4599 (O_4599,N_48221,N_48694);
xor UO_4600 (O_4600,N_40145,N_42235);
nor UO_4601 (O_4601,N_43670,N_47476);
nor UO_4602 (O_4602,N_41870,N_44719);
and UO_4603 (O_4603,N_49033,N_44170);
nand UO_4604 (O_4604,N_41969,N_41314);
nor UO_4605 (O_4605,N_44685,N_44010);
and UO_4606 (O_4606,N_41902,N_47058);
xor UO_4607 (O_4607,N_46675,N_42913);
xor UO_4608 (O_4608,N_48172,N_46186);
or UO_4609 (O_4609,N_48916,N_45327);
or UO_4610 (O_4610,N_47300,N_42015);
xnor UO_4611 (O_4611,N_49913,N_46111);
or UO_4612 (O_4612,N_41480,N_43986);
nand UO_4613 (O_4613,N_43935,N_44585);
nand UO_4614 (O_4614,N_48178,N_48214);
or UO_4615 (O_4615,N_49869,N_40486);
nor UO_4616 (O_4616,N_43858,N_40628);
xor UO_4617 (O_4617,N_43022,N_42707);
and UO_4618 (O_4618,N_48906,N_46764);
nor UO_4619 (O_4619,N_40099,N_42777);
and UO_4620 (O_4620,N_43993,N_43684);
xnor UO_4621 (O_4621,N_43799,N_47763);
and UO_4622 (O_4622,N_49374,N_49510);
or UO_4623 (O_4623,N_45936,N_48855);
xor UO_4624 (O_4624,N_48566,N_45160);
nor UO_4625 (O_4625,N_44656,N_49026);
nand UO_4626 (O_4626,N_47499,N_44082);
nor UO_4627 (O_4627,N_41440,N_41957);
or UO_4628 (O_4628,N_46377,N_45395);
xor UO_4629 (O_4629,N_43735,N_46323);
xor UO_4630 (O_4630,N_47059,N_46625);
or UO_4631 (O_4631,N_44377,N_41762);
xor UO_4632 (O_4632,N_47736,N_41740);
nand UO_4633 (O_4633,N_49584,N_49199);
and UO_4634 (O_4634,N_42223,N_42694);
nand UO_4635 (O_4635,N_42812,N_48029);
xor UO_4636 (O_4636,N_48256,N_43604);
or UO_4637 (O_4637,N_49988,N_49876);
xor UO_4638 (O_4638,N_42018,N_47111);
nor UO_4639 (O_4639,N_49140,N_43162);
nand UO_4640 (O_4640,N_42218,N_44815);
nand UO_4641 (O_4641,N_45910,N_43291);
nor UO_4642 (O_4642,N_46501,N_40718);
xnor UO_4643 (O_4643,N_49148,N_43827);
nor UO_4644 (O_4644,N_48619,N_48451);
and UO_4645 (O_4645,N_40838,N_46609);
nor UO_4646 (O_4646,N_48083,N_47068);
and UO_4647 (O_4647,N_48397,N_45672);
nor UO_4648 (O_4648,N_45809,N_44568);
xnor UO_4649 (O_4649,N_43775,N_45985);
nand UO_4650 (O_4650,N_40446,N_48892);
nand UO_4651 (O_4651,N_43784,N_49240);
and UO_4652 (O_4652,N_44814,N_49814);
xnor UO_4653 (O_4653,N_41306,N_48327);
and UO_4654 (O_4654,N_40205,N_41542);
nand UO_4655 (O_4655,N_43689,N_42156);
and UO_4656 (O_4656,N_48213,N_47483);
nor UO_4657 (O_4657,N_45332,N_44552);
xor UO_4658 (O_4658,N_49366,N_49533);
xnor UO_4659 (O_4659,N_44267,N_47774);
xor UO_4660 (O_4660,N_48714,N_49966);
and UO_4661 (O_4661,N_41293,N_42338);
and UO_4662 (O_4662,N_41041,N_47752);
xor UO_4663 (O_4663,N_49951,N_48976);
or UO_4664 (O_4664,N_47707,N_41555);
nand UO_4665 (O_4665,N_42822,N_46381);
and UO_4666 (O_4666,N_43860,N_42594);
or UO_4667 (O_4667,N_41693,N_42932);
nand UO_4668 (O_4668,N_46931,N_42416);
nor UO_4669 (O_4669,N_40868,N_49906);
nor UO_4670 (O_4670,N_49153,N_46350);
nand UO_4671 (O_4671,N_47624,N_40043);
nor UO_4672 (O_4672,N_45202,N_40881);
or UO_4673 (O_4673,N_42398,N_47591);
and UO_4674 (O_4674,N_41610,N_47246);
nor UO_4675 (O_4675,N_41876,N_47747);
nor UO_4676 (O_4676,N_40397,N_43007);
nand UO_4677 (O_4677,N_48612,N_49903);
and UO_4678 (O_4678,N_47898,N_42404);
or UO_4679 (O_4679,N_46731,N_44073);
nand UO_4680 (O_4680,N_47336,N_47515);
or UO_4681 (O_4681,N_44964,N_49088);
and UO_4682 (O_4682,N_46399,N_49337);
nand UO_4683 (O_4683,N_47857,N_48958);
nand UO_4684 (O_4684,N_49194,N_41496);
xnor UO_4685 (O_4685,N_40733,N_49625);
nand UO_4686 (O_4686,N_43687,N_44731);
xnor UO_4687 (O_4687,N_43841,N_48414);
nand UO_4688 (O_4688,N_49875,N_46757);
nand UO_4689 (O_4689,N_48018,N_49582);
nor UO_4690 (O_4690,N_46153,N_46804);
nor UO_4691 (O_4691,N_48509,N_42129);
nor UO_4692 (O_4692,N_43237,N_48826);
and UO_4693 (O_4693,N_43648,N_47305);
nand UO_4694 (O_4694,N_42895,N_42919);
nand UO_4695 (O_4695,N_46665,N_47220);
or UO_4696 (O_4696,N_45940,N_40758);
or UO_4697 (O_4697,N_47114,N_47607);
nor UO_4698 (O_4698,N_43099,N_44414);
nand UO_4699 (O_4699,N_44478,N_48252);
and UO_4700 (O_4700,N_47044,N_45366);
nand UO_4701 (O_4701,N_46987,N_48088);
xor UO_4702 (O_4702,N_42013,N_40789);
xor UO_4703 (O_4703,N_43699,N_40214);
xnor UO_4704 (O_4704,N_48331,N_48793);
or UO_4705 (O_4705,N_46413,N_46330);
xor UO_4706 (O_4706,N_41421,N_41716);
xnor UO_4707 (O_4707,N_48465,N_42288);
nor UO_4708 (O_4708,N_40850,N_45191);
nor UO_4709 (O_4709,N_46772,N_42889);
and UO_4710 (O_4710,N_40195,N_43240);
and UO_4711 (O_4711,N_46171,N_46718);
and UO_4712 (O_4712,N_48919,N_46362);
xor UO_4713 (O_4713,N_49222,N_49177);
or UO_4714 (O_4714,N_49172,N_48591);
nor UO_4715 (O_4715,N_46301,N_41031);
or UO_4716 (O_4716,N_44383,N_40678);
or UO_4717 (O_4717,N_40896,N_42464);
nand UO_4718 (O_4718,N_44087,N_40590);
nor UO_4719 (O_4719,N_43917,N_41133);
and UO_4720 (O_4720,N_46163,N_48988);
and UO_4721 (O_4721,N_49879,N_49115);
and UO_4722 (O_4722,N_44529,N_46194);
or UO_4723 (O_4723,N_46376,N_49666);
nor UO_4724 (O_4724,N_42465,N_45062);
nand UO_4725 (O_4725,N_49517,N_48313);
nand UO_4726 (O_4726,N_41680,N_47447);
xnor UO_4727 (O_4727,N_42315,N_45734);
and UO_4728 (O_4728,N_42311,N_40810);
nand UO_4729 (O_4729,N_44500,N_41519);
nor UO_4730 (O_4730,N_42081,N_46222);
or UO_4731 (O_4731,N_40200,N_46729);
nor UO_4732 (O_4732,N_42164,N_41056);
or UO_4733 (O_4733,N_44238,N_48985);
or UO_4734 (O_4734,N_45365,N_47519);
nand UO_4735 (O_4735,N_46878,N_45935);
nand UO_4736 (O_4736,N_41435,N_49219);
nand UO_4737 (O_4737,N_43619,N_44906);
and UO_4738 (O_4738,N_49182,N_49986);
nand UO_4739 (O_4739,N_40466,N_45526);
and UO_4740 (O_4740,N_45118,N_45684);
nand UO_4741 (O_4741,N_40069,N_47193);
xnor UO_4742 (O_4742,N_45207,N_48417);
xnor UO_4743 (O_4743,N_40057,N_42411);
or UO_4744 (O_4744,N_49029,N_47410);
xor UO_4745 (O_4745,N_49611,N_49391);
xor UO_4746 (O_4746,N_41456,N_46182);
and UO_4747 (O_4747,N_41088,N_44778);
or UO_4748 (O_4748,N_43168,N_49595);
nand UO_4749 (O_4749,N_46489,N_44921);
nor UO_4750 (O_4750,N_46334,N_46092);
nor UO_4751 (O_4751,N_40541,N_48739);
nor UO_4752 (O_4752,N_46254,N_43066);
or UO_4753 (O_4753,N_45634,N_41338);
and UO_4754 (O_4754,N_41107,N_46852);
and UO_4755 (O_4755,N_42027,N_41890);
nor UO_4756 (O_4756,N_46935,N_45653);
xnor UO_4757 (O_4757,N_46601,N_41297);
or UO_4758 (O_4758,N_41709,N_43750);
or UO_4759 (O_4759,N_40542,N_42848);
xor UO_4760 (O_4760,N_47445,N_42424);
xnor UO_4761 (O_4761,N_45150,N_45992);
or UO_4762 (O_4762,N_47867,N_40697);
xor UO_4763 (O_4763,N_46076,N_47567);
or UO_4764 (O_4764,N_45308,N_40631);
xnor UO_4765 (O_4765,N_40215,N_48072);
xnor UO_4766 (O_4766,N_46626,N_44179);
nand UO_4767 (O_4767,N_41794,N_42096);
and UO_4768 (O_4768,N_40940,N_46833);
nor UO_4769 (O_4769,N_44237,N_49772);
and UO_4770 (O_4770,N_41013,N_46638);
or UO_4771 (O_4771,N_47319,N_45534);
nor UO_4772 (O_4772,N_46810,N_49067);
or UO_4773 (O_4773,N_41718,N_45730);
xor UO_4774 (O_4774,N_40808,N_45269);
nor UO_4775 (O_4775,N_47313,N_47444);
xnor UO_4776 (O_4776,N_42846,N_41167);
nand UO_4777 (O_4777,N_49130,N_41834);
nor UO_4778 (O_4778,N_46158,N_43453);
nor UO_4779 (O_4779,N_45079,N_46424);
or UO_4780 (O_4780,N_40493,N_49565);
nand UO_4781 (O_4781,N_43487,N_41673);
nor UO_4782 (O_4782,N_46011,N_41488);
and UO_4783 (O_4783,N_43817,N_44722);
xnor UO_4784 (O_4784,N_48508,N_41158);
nand UO_4785 (O_4785,N_42779,N_41575);
xor UO_4786 (O_4786,N_47431,N_43367);
nor UO_4787 (O_4787,N_49805,N_40741);
and UO_4788 (O_4788,N_43811,N_41546);
or UO_4789 (O_4789,N_40564,N_47054);
or UO_4790 (O_4790,N_40973,N_49110);
nor UO_4791 (O_4791,N_43591,N_48416);
or UO_4792 (O_4792,N_46164,N_43198);
nand UO_4793 (O_4793,N_48832,N_48197);
or UO_4794 (O_4794,N_48956,N_45504);
and UO_4795 (O_4795,N_45924,N_45394);
nor UO_4796 (O_4796,N_41422,N_41735);
and UO_4797 (O_4797,N_48704,N_46508);
or UO_4798 (O_4798,N_49928,N_45056);
xnor UO_4799 (O_4799,N_43422,N_47192);
nor UO_4800 (O_4800,N_49542,N_49101);
xnor UO_4801 (O_4801,N_41253,N_40288);
or UO_4802 (O_4802,N_47308,N_44952);
and UO_4803 (O_4803,N_48054,N_47715);
or UO_4804 (O_4804,N_40049,N_49567);
or UO_4805 (O_4805,N_46911,N_41569);
or UO_4806 (O_4806,N_46866,N_47052);
xnor UO_4807 (O_4807,N_47711,N_45557);
nand UO_4808 (O_4808,N_40029,N_49440);
or UO_4809 (O_4809,N_46272,N_43880);
xnor UO_4810 (O_4810,N_45952,N_42780);
or UO_4811 (O_4811,N_43192,N_48374);
or UO_4812 (O_4812,N_40895,N_48071);
or UO_4813 (O_4813,N_47496,N_44671);
or UO_4814 (O_4814,N_42055,N_49428);
nand UO_4815 (O_4815,N_43779,N_41906);
nor UO_4816 (O_4816,N_47970,N_48651);
nor UO_4817 (O_4817,N_41691,N_44312);
or UO_4818 (O_4818,N_45057,N_42995);
and UO_4819 (O_4819,N_45749,N_41727);
or UO_4820 (O_4820,N_48809,N_44919);
and UO_4821 (O_4821,N_46261,N_49766);
or UO_4822 (O_4822,N_48928,N_45231);
and UO_4823 (O_4823,N_42228,N_41752);
nand UO_4824 (O_4824,N_46820,N_47286);
or UO_4825 (O_4825,N_45246,N_42937);
nor UO_4826 (O_4826,N_41801,N_41506);
and UO_4827 (O_4827,N_40744,N_49163);
and UO_4828 (O_4828,N_49561,N_46453);
xnor UO_4829 (O_4829,N_42756,N_40122);
xor UO_4830 (O_4830,N_45716,N_45109);
xor UO_4831 (O_4831,N_47552,N_42850);
nor UO_4832 (O_4832,N_41495,N_42471);
or UO_4833 (O_4833,N_44652,N_45168);
xor UO_4834 (O_4834,N_40071,N_42669);
nand UO_4835 (O_4835,N_43195,N_44987);
and UO_4836 (O_4836,N_42474,N_43440);
xnor UO_4837 (O_4837,N_42952,N_43569);
and UO_4838 (O_4838,N_40220,N_44404);
nor UO_4839 (O_4839,N_48125,N_47671);
nor UO_4840 (O_4840,N_41946,N_40624);
or UO_4841 (O_4841,N_45406,N_45357);
xnor UO_4842 (O_4842,N_49333,N_40059);
and UO_4843 (O_4843,N_44644,N_47367);
nor UO_4844 (O_4844,N_44368,N_46223);
nor UO_4845 (O_4845,N_48800,N_42573);
and UO_4846 (O_4846,N_49818,N_46021);
and UO_4847 (O_4847,N_49127,N_48351);
and UO_4848 (O_4848,N_41633,N_44369);
or UO_4849 (O_4849,N_43642,N_48064);
or UO_4850 (O_4850,N_40391,N_44743);
or UO_4851 (O_4851,N_40894,N_43103);
nand UO_4852 (O_4852,N_43812,N_45064);
nor UO_4853 (O_4853,N_41455,N_44303);
or UO_4854 (O_4854,N_46663,N_42446);
nand UO_4855 (O_4855,N_48518,N_45355);
and UO_4856 (O_4856,N_43209,N_41331);
nor UO_4857 (O_4857,N_42912,N_43029);
xnor UO_4858 (O_4858,N_41894,N_46232);
nand UO_4859 (O_4859,N_45835,N_44417);
xnor UO_4860 (O_4860,N_48280,N_43153);
xnor UO_4861 (O_4861,N_48669,N_47082);
and UO_4862 (O_4862,N_45158,N_46135);
or UO_4863 (O_4863,N_43279,N_40267);
xor UO_4864 (O_4864,N_43128,N_45773);
nand UO_4865 (O_4865,N_40313,N_44920);
nor UO_4866 (O_4866,N_48963,N_42536);
nor UO_4867 (O_4867,N_45857,N_42651);
nor UO_4868 (O_4868,N_43666,N_44210);
or UO_4869 (O_4869,N_45206,N_47564);
nand UO_4870 (O_4870,N_47086,N_44446);
nand UO_4871 (O_4871,N_49507,N_45385);
or UO_4872 (O_4872,N_42258,N_40354);
or UO_4873 (O_4873,N_49449,N_42359);
or UO_4874 (O_4874,N_42365,N_48343);
and UO_4875 (O_4875,N_41971,N_45089);
nand UO_4876 (O_4876,N_43355,N_45801);
and UO_4877 (O_4877,N_46895,N_43524);
nor UO_4878 (O_4878,N_42083,N_47696);
or UO_4879 (O_4879,N_43244,N_44088);
xor UO_4880 (O_4880,N_43394,N_43331);
or UO_4881 (O_4881,N_42153,N_49048);
xnor UO_4882 (O_4882,N_43432,N_48753);
xor UO_4883 (O_4883,N_42838,N_40972);
nand UO_4884 (O_4884,N_47304,N_49855);
nor UO_4885 (O_4885,N_46504,N_49450);
nor UO_4886 (O_4886,N_49797,N_40064);
nand UO_4887 (O_4887,N_46517,N_43064);
and UO_4888 (O_4888,N_42552,N_47182);
nor UO_4889 (O_4889,N_40109,N_42043);
xnor UO_4890 (O_4890,N_46465,N_41424);
and UO_4891 (O_4891,N_49905,N_48293);
and UO_4892 (O_4892,N_40236,N_43392);
or UO_4893 (O_4893,N_45404,N_42686);
or UO_4894 (O_4894,N_44297,N_44806);
and UO_4895 (O_4895,N_40975,N_42399);
xor UO_4896 (O_4896,N_42348,N_42733);
nor UO_4897 (O_4897,N_42279,N_43963);
or UO_4898 (O_4898,N_40923,N_47346);
nor UO_4899 (O_4899,N_49774,N_49357);
and UO_4900 (O_4900,N_42369,N_41921);
and UO_4901 (O_4901,N_41949,N_49878);
or UO_4902 (O_4902,N_45351,N_42877);
and UO_4903 (O_4903,N_47932,N_40168);
and UO_4904 (O_4904,N_40279,N_46554);
nor UO_4905 (O_4905,N_46128,N_43681);
xor UO_4906 (O_4906,N_49069,N_47243);
and UO_4907 (O_4907,N_46339,N_41429);
xor UO_4908 (O_4908,N_43778,N_49711);
or UO_4909 (O_4909,N_42630,N_42584);
nor UO_4910 (O_4910,N_48444,N_45753);
nand UO_4911 (O_4911,N_45796,N_48561);
nor UO_4912 (O_4912,N_49277,N_41202);
nand UO_4913 (O_4913,N_48431,N_45321);
nand UO_4914 (O_4914,N_47414,N_44409);
nand UO_4915 (O_4915,N_40235,N_46778);
xor UO_4916 (O_4916,N_44601,N_42287);
xor UO_4917 (O_4917,N_48379,N_48039);
nor UO_4918 (O_4918,N_48391,N_43111);
nor UO_4919 (O_4919,N_47528,N_46177);
and UO_4920 (O_4920,N_42741,N_46510);
nor UO_4921 (O_4921,N_48193,N_41719);
and UO_4922 (O_4922,N_41223,N_49228);
nand UO_4923 (O_4923,N_43016,N_48494);
nor UO_4924 (O_4924,N_43469,N_44828);
and UO_4925 (O_4925,N_44772,N_44030);
xor UO_4926 (O_4926,N_48003,N_43702);
or UO_4927 (O_4927,N_45210,N_44113);
xor UO_4928 (O_4928,N_42420,N_44880);
nor UO_4929 (O_4929,N_45151,N_40290);
nand UO_4930 (O_4930,N_42011,N_48564);
nand UO_4931 (O_4931,N_46622,N_43220);
or UO_4932 (O_4932,N_48971,N_40581);
or UO_4933 (O_4933,N_47906,N_40851);
and UO_4934 (O_4934,N_44136,N_49506);
xor UO_4935 (O_4935,N_41866,N_45708);
and UO_4936 (O_4936,N_49137,N_49749);
or UO_4937 (O_4937,N_41370,N_49833);
xnor UO_4938 (O_4938,N_40525,N_41840);
and UO_4939 (O_4939,N_41644,N_41108);
nand UO_4940 (O_4940,N_40128,N_49135);
or UO_4941 (O_4941,N_49379,N_45437);
or UO_4942 (O_4942,N_47064,N_41100);
or UO_4943 (O_4943,N_49464,N_41276);
nand UO_4944 (O_4944,N_43457,N_47373);
or UO_4945 (O_4945,N_43171,N_40887);
and UO_4946 (O_4946,N_41604,N_49744);
nor UO_4947 (O_4947,N_46687,N_45615);
nor UO_4948 (O_4948,N_42292,N_41609);
and UO_4949 (O_4949,N_47356,N_42320);
nand UO_4950 (O_4950,N_45520,N_43467);
and UO_4951 (O_4951,N_44800,N_40351);
xor UO_4952 (O_4952,N_42870,N_44005);
and UO_4953 (O_4953,N_45666,N_44266);
and UO_4954 (O_4954,N_44107,N_45477);
and UO_4955 (O_4955,N_46411,N_49553);
or UO_4956 (O_4956,N_40711,N_44428);
xnor UO_4957 (O_4957,N_41252,N_47470);
nor UO_4958 (O_4958,N_48244,N_47997);
nor UO_4959 (O_4959,N_41473,N_42564);
and UO_4960 (O_4960,N_42144,N_41072);
nor UO_4961 (O_4961,N_46610,N_46452);
xor UO_4962 (O_4962,N_45863,N_40684);
and UO_4963 (O_4963,N_40579,N_48001);
xnor UO_4964 (O_4964,N_45984,N_46793);
and UO_4965 (O_4965,N_44766,N_49598);
or UO_4966 (O_4966,N_45374,N_46594);
and UO_4967 (O_4967,N_40452,N_47115);
or UO_4968 (O_4968,N_44533,N_40958);
and UO_4969 (O_4969,N_45096,N_41682);
nand UO_4970 (O_4970,N_43092,N_43900);
nand UO_4971 (O_4971,N_41939,N_42039);
or UO_4972 (O_4972,N_48082,N_49690);
or UO_4973 (O_4973,N_41469,N_48346);
nor UO_4974 (O_4974,N_45511,N_42291);
nor UO_4975 (O_4975,N_43839,N_40272);
xnor UO_4976 (O_4976,N_41042,N_43980);
nand UO_4977 (O_4977,N_45354,N_40787);
nor UO_4978 (O_4978,N_42502,N_42132);
xnor UO_4979 (O_4979,N_46780,N_43346);
nand UO_4980 (O_4980,N_49206,N_49481);
and UO_4981 (O_4981,N_42487,N_43144);
and UO_4982 (O_4982,N_46746,N_42482);
or UO_4983 (O_4983,N_48823,N_43823);
or UO_4984 (O_4984,N_45976,N_43233);
and UO_4985 (O_4985,N_41073,N_42302);
and UO_4986 (O_4986,N_45307,N_49176);
or UO_4987 (O_4987,N_44973,N_44649);
nand UO_4988 (O_4988,N_43580,N_42965);
and UO_4989 (O_4989,N_41209,N_46242);
nand UO_4990 (O_4990,N_45172,N_46084);
xnor UO_4991 (O_4991,N_42656,N_43454);
xor UO_4992 (O_4992,N_43530,N_40897);
nand UO_4993 (O_4993,N_43659,N_42523);
xnor UO_4994 (O_4994,N_40954,N_44456);
or UO_4995 (O_4995,N_41970,N_45963);
and UO_4996 (O_4996,N_43427,N_48133);
and UO_4997 (O_4997,N_49319,N_48511);
xnor UO_4998 (O_4998,N_49396,N_43828);
nor UO_4999 (O_4999,N_48895,N_47039);
endmodule