module basic_1500_15000_2000_5_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_1301,In_573);
nand U1 (N_1,In_1171,In_663);
or U2 (N_2,In_1123,In_238);
nor U3 (N_3,In_630,In_893);
nand U4 (N_4,In_683,In_75);
nand U5 (N_5,In_1398,In_1302);
and U6 (N_6,In_140,In_1349);
xnor U7 (N_7,In_143,In_876);
nand U8 (N_8,In_1245,In_1083);
nor U9 (N_9,In_789,In_1283);
xor U10 (N_10,In_1189,In_72);
xnor U11 (N_11,In_1493,In_91);
xor U12 (N_12,In_1394,In_791);
and U13 (N_13,In_1144,In_491);
xor U14 (N_14,In_1403,In_361);
xor U15 (N_15,In_1456,In_196);
and U16 (N_16,In_1321,In_103);
nor U17 (N_17,In_468,In_183);
or U18 (N_18,In_656,In_287);
and U19 (N_19,In_526,In_706);
xnor U20 (N_20,In_705,In_785);
nor U21 (N_21,In_744,In_1054);
nor U22 (N_22,In_12,In_169);
or U23 (N_23,In_1066,In_1401);
xnor U24 (N_24,In_1478,In_21);
and U25 (N_25,In_1085,In_1204);
nor U26 (N_26,In_174,In_884);
or U27 (N_27,In_1001,In_1467);
or U28 (N_28,In_1265,In_478);
and U29 (N_29,In_356,In_1327);
nand U30 (N_30,In_1396,In_1243);
nor U31 (N_31,In_144,In_606);
nor U32 (N_32,In_610,In_992);
or U33 (N_33,In_1412,In_503);
or U34 (N_34,In_989,In_1450);
xnor U35 (N_35,In_569,In_245);
and U36 (N_36,In_1109,In_1421);
or U37 (N_37,In_123,In_321);
nor U38 (N_38,In_899,In_94);
xor U39 (N_39,In_659,In_901);
nand U40 (N_40,In_1309,In_1135);
and U41 (N_41,In_801,In_378);
and U42 (N_42,In_182,In_518);
and U43 (N_43,In_166,In_519);
and U44 (N_44,In_187,In_1288);
or U45 (N_45,In_684,In_743);
xor U46 (N_46,In_1365,In_550);
nand U47 (N_47,In_682,In_413);
and U48 (N_48,In_1381,In_1356);
nand U49 (N_49,In_1022,In_296);
nand U50 (N_50,In_52,In_1025);
nor U51 (N_51,In_6,In_699);
and U52 (N_52,In_930,In_243);
or U53 (N_53,In_765,In_620);
nand U54 (N_54,In_1073,In_186);
nor U55 (N_55,In_119,In_685);
and U56 (N_56,In_353,In_1407);
nand U57 (N_57,In_104,In_538);
xor U58 (N_58,In_763,In_1387);
or U59 (N_59,In_708,In_397);
and U60 (N_60,In_940,In_365);
or U61 (N_61,In_329,In_881);
nand U62 (N_62,In_475,In_253);
nor U63 (N_63,In_107,In_136);
xor U64 (N_64,In_770,In_464);
and U65 (N_65,In_1206,In_1297);
and U66 (N_66,In_1417,In_386);
or U67 (N_67,In_208,In_1136);
or U68 (N_68,In_761,In_390);
nand U69 (N_69,In_295,In_157);
nor U70 (N_70,In_480,In_835);
xnor U71 (N_71,In_1148,In_1378);
or U72 (N_72,In_1416,In_270);
nand U73 (N_73,In_634,In_534);
nand U74 (N_74,In_37,In_1488);
and U75 (N_75,In_758,In_1413);
nor U76 (N_76,In_1331,In_665);
xor U77 (N_77,In_316,In_1395);
nand U78 (N_78,In_1353,In_147);
and U79 (N_79,In_1350,In_318);
nor U80 (N_80,In_1479,In_1352);
and U81 (N_81,In_448,In_330);
nand U82 (N_82,In_1277,In_237);
nor U83 (N_83,In_1452,In_1196);
and U84 (N_84,In_1386,In_953);
or U85 (N_85,In_363,In_1260);
and U86 (N_86,In_830,In_1354);
nor U87 (N_87,In_324,In_589);
and U88 (N_88,In_779,In_585);
and U89 (N_89,In_343,In_1141);
nand U90 (N_90,In_996,In_939);
or U91 (N_91,In_1047,In_675);
nor U92 (N_92,In_1053,In_209);
nand U93 (N_93,In_1190,In_148);
and U94 (N_94,In_1465,In_1094);
nand U95 (N_95,In_1179,In_1017);
nor U96 (N_96,In_780,In_516);
or U97 (N_97,In_331,In_1463);
or U98 (N_98,In_439,In_979);
xnor U99 (N_99,In_161,In_34);
xnor U100 (N_100,In_1498,In_1182);
xnor U101 (N_101,In_220,In_1439);
nor U102 (N_102,In_179,In_333);
or U103 (N_103,In_470,In_1003);
nor U104 (N_104,In_215,In_1108);
and U105 (N_105,In_1121,In_142);
and U106 (N_106,In_15,In_1132);
xor U107 (N_107,In_738,In_697);
xor U108 (N_108,In_1226,In_1170);
or U109 (N_109,In_995,In_877);
xnor U110 (N_110,In_1449,In_1486);
nand U111 (N_111,In_1028,In_251);
nand U112 (N_112,In_751,In_558);
nand U113 (N_113,In_1207,In_312);
and U114 (N_114,In_1448,In_1459);
or U115 (N_115,In_1419,In_615);
nand U116 (N_116,In_134,In_872);
xor U117 (N_117,In_384,In_1031);
xor U118 (N_118,In_1317,In_497);
nand U119 (N_119,In_87,In_1186);
or U120 (N_120,In_1293,In_1058);
xnor U121 (N_121,In_855,In_734);
and U122 (N_122,In_1296,In_978);
nand U123 (N_123,In_1104,In_756);
nand U124 (N_124,In_667,In_1219);
nor U125 (N_125,In_1029,In_96);
and U126 (N_126,In_84,In_1015);
nor U127 (N_127,In_944,In_520);
xor U128 (N_128,In_152,In_1092);
or U129 (N_129,In_614,In_947);
and U130 (N_130,In_1429,In_1198);
xor U131 (N_131,In_976,In_809);
nor U132 (N_132,In_45,In_172);
xnor U133 (N_133,In_210,In_1079);
xnor U134 (N_134,In_406,In_882);
or U135 (N_135,In_1369,In_1099);
and U136 (N_136,In_403,In_1295);
nand U137 (N_137,In_0,In_693);
and U138 (N_138,In_78,In_733);
and U139 (N_139,In_803,In_1462);
xor U140 (N_140,In_849,In_1342);
xor U141 (N_141,In_900,In_1347);
nor U142 (N_142,In_1075,In_198);
nor U143 (N_143,In_185,In_891);
xnor U144 (N_144,In_974,In_422);
or U145 (N_145,In_1337,In_1322);
or U146 (N_146,In_871,In_1300);
and U147 (N_147,In_609,In_1193);
nor U148 (N_148,In_279,In_857);
and U149 (N_149,In_931,In_396);
and U150 (N_150,In_1051,In_13);
and U151 (N_151,In_374,In_44);
nor U152 (N_152,In_1238,In_820);
and U153 (N_153,In_1161,In_1359);
xor U154 (N_154,In_507,In_1495);
xor U155 (N_155,In_284,In_798);
and U156 (N_156,In_224,In_1246);
nand U157 (N_157,In_1038,In_115);
nand U158 (N_158,In_1059,In_263);
nand U159 (N_159,In_824,In_1101);
xnor U160 (N_160,In_8,In_1158);
nor U161 (N_161,In_175,In_178);
and U162 (N_162,In_83,In_309);
or U163 (N_163,In_963,In_275);
xnor U164 (N_164,In_1304,In_100);
or U165 (N_165,In_752,In_637);
nand U166 (N_166,In_278,In_582);
nor U167 (N_167,In_1026,In_1131);
nand U168 (N_168,In_1250,In_1223);
or U169 (N_169,In_1409,In_441);
nor U170 (N_170,In_1060,In_1270);
nor U171 (N_171,In_97,In_1251);
nand U172 (N_172,In_299,In_1320);
nand U173 (N_173,In_965,In_50);
nand U174 (N_174,In_677,In_866);
xor U175 (N_175,In_1384,In_1389);
xnor U176 (N_176,In_966,In_66);
nand U177 (N_177,In_796,In_367);
nand U178 (N_178,In_133,In_490);
nand U179 (N_179,In_845,In_1112);
or U180 (N_180,In_810,In_335);
nand U181 (N_181,In_393,In_354);
and U182 (N_182,In_1232,In_282);
and U183 (N_183,In_1166,In_1247);
or U184 (N_184,In_39,In_207);
xnor U185 (N_185,In_631,In_1007);
nand U186 (N_186,In_570,In_346);
nand U187 (N_187,In_760,In_303);
or U188 (N_188,In_306,In_276);
nor U189 (N_189,In_1391,In_364);
nand U190 (N_190,In_1485,In_280);
or U191 (N_191,In_1457,In_273);
nand U192 (N_192,In_586,In_509);
and U193 (N_193,In_466,In_216);
or U194 (N_194,In_1306,In_1267);
nor U195 (N_195,In_991,In_73);
nand U196 (N_196,In_943,In_1040);
and U197 (N_197,In_76,In_1216);
or U198 (N_198,In_19,In_577);
xnor U199 (N_199,In_1291,In_1063);
nor U200 (N_200,In_1415,In_56);
and U201 (N_201,In_1211,In_409);
xnor U202 (N_202,In_485,In_594);
xnor U203 (N_203,In_452,In_1185);
and U204 (N_204,In_696,In_671);
or U205 (N_205,In_177,In_20);
xnor U206 (N_206,In_494,In_607);
xnor U207 (N_207,In_351,In_1392);
nor U208 (N_208,In_408,In_1192);
and U209 (N_209,In_532,In_1023);
nand U210 (N_210,In_920,In_587);
or U211 (N_211,In_269,In_840);
nand U212 (N_212,In_493,In_896);
nand U213 (N_213,In_1009,In_151);
xnor U214 (N_214,In_1146,In_392);
xor U215 (N_215,In_806,In_1200);
xor U216 (N_216,In_687,In_540);
nand U217 (N_217,In_79,In_1050);
nor U218 (N_218,In_105,In_1366);
nand U219 (N_219,In_993,In_58);
nor U220 (N_220,In_852,In_811);
nand U221 (N_221,In_626,In_720);
xor U222 (N_222,In_542,In_1011);
nor U223 (N_223,In_247,In_1049);
and U224 (N_224,In_1290,In_563);
or U225 (N_225,In_874,In_323);
nand U226 (N_226,In_1126,In_604);
nor U227 (N_227,In_851,In_1425);
xor U228 (N_228,In_48,In_1002);
and U229 (N_229,In_7,In_795);
nor U230 (N_230,In_447,In_605);
or U231 (N_231,In_1351,In_244);
or U232 (N_232,In_1253,In_1379);
nand U233 (N_233,In_1315,In_1134);
nand U234 (N_234,In_618,In_360);
nor U235 (N_235,In_814,In_870);
nor U236 (N_236,In_660,In_514);
and U237 (N_237,In_646,In_1205);
xor U238 (N_238,In_918,In_1110);
or U239 (N_239,In_1080,In_1338);
or U240 (N_240,In_479,In_205);
and U241 (N_241,In_1242,In_1008);
or U242 (N_242,In_1077,In_1323);
nor U243 (N_243,In_93,In_528);
or U244 (N_244,In_1249,In_1256);
nor U245 (N_245,In_666,In_90);
nand U246 (N_246,In_1318,In_301);
or U247 (N_247,In_815,In_595);
xor U248 (N_248,In_669,In_249);
xor U249 (N_249,In_1362,In_990);
or U250 (N_250,In_1325,In_1018);
and U251 (N_251,In_1328,In_1129);
nor U252 (N_252,In_293,In_593);
xnor U253 (N_253,In_305,In_846);
and U254 (N_254,In_914,In_822);
nand U255 (N_255,In_977,In_1163);
nor U256 (N_256,In_612,In_640);
or U257 (N_257,In_496,In_372);
or U258 (N_258,In_718,In_1105);
or U259 (N_259,In_433,In_1484);
or U260 (N_260,In_1220,In_1169);
and U261 (N_261,In_1422,In_499);
xnor U262 (N_262,In_895,In_43);
xnor U263 (N_263,In_1371,In_1167);
xnor U264 (N_264,In_204,In_116);
xnor U265 (N_265,In_1043,In_171);
and U266 (N_266,In_150,In_1102);
nor U267 (N_267,In_1497,In_121);
nand U268 (N_268,In_1175,In_689);
nor U269 (N_269,In_435,In_544);
or U270 (N_270,In_1284,In_304);
or U271 (N_271,In_442,In_674);
xor U272 (N_272,In_1461,In_401);
xnor U273 (N_273,In_16,In_596);
nor U274 (N_274,In_1294,In_704);
xor U275 (N_275,In_928,In_691);
xnor U276 (N_276,In_938,In_42);
and U277 (N_277,In_77,In_213);
xor U278 (N_278,In_985,In_658);
and U279 (N_279,In_1287,In_1202);
xnor U280 (N_280,In_1036,In_265);
or U281 (N_281,In_581,In_1024);
xor U282 (N_282,In_1239,In_664);
or U283 (N_283,In_1305,In_1181);
and U284 (N_284,In_601,In_359);
xnor U285 (N_285,In_232,In_239);
xor U286 (N_286,In_410,In_381);
nand U287 (N_287,In_1312,In_235);
nor U288 (N_288,In_565,In_1272);
nand U289 (N_289,In_285,In_854);
nor U290 (N_290,In_1255,In_842);
nor U291 (N_291,In_522,In_561);
nand U292 (N_292,In_212,In_1042);
nor U293 (N_293,In_680,In_54);
or U294 (N_294,In_418,In_935);
xor U295 (N_295,In_1069,In_613);
nand U296 (N_296,In_986,In_1234);
nor U297 (N_297,In_767,In_181);
nand U298 (N_298,In_564,In_737);
and U299 (N_299,In_512,In_1435);
or U300 (N_300,In_787,In_110);
or U301 (N_301,In_81,In_1237);
nor U302 (N_302,In_252,In_1339);
xor U303 (N_303,In_1057,In_288);
or U304 (N_304,In_1269,In_964);
or U305 (N_305,In_527,In_719);
or U306 (N_306,In_913,In_414);
xnor U307 (N_307,In_619,In_860);
xor U308 (N_308,In_444,In_1274);
and U309 (N_309,In_4,In_217);
nor U310 (N_310,In_379,In_112);
xor U311 (N_311,In_428,In_813);
and U312 (N_312,In_531,In_59);
nand U313 (N_313,In_729,In_546);
nand U314 (N_314,In_853,In_598);
and U315 (N_315,In_289,In_25);
xnor U316 (N_316,In_1152,In_632);
or U317 (N_317,In_1364,In_1373);
and U318 (N_318,In_1056,In_398);
or U319 (N_319,In_957,In_1032);
and U320 (N_320,In_535,In_1363);
xor U321 (N_321,In_457,In_508);
and U322 (N_322,In_1428,In_591);
or U323 (N_323,In_347,In_1162);
and U324 (N_324,In_382,In_1133);
or U325 (N_325,In_562,In_924);
nand U326 (N_326,In_1156,In_225);
and U327 (N_327,In_972,In_625);
nor U328 (N_328,In_68,In_721);
nor U329 (N_329,In_825,In_1341);
or U330 (N_330,In_818,In_628);
nor U331 (N_331,In_462,In_1262);
xor U332 (N_332,In_17,In_755);
or U333 (N_333,In_388,In_994);
and U334 (N_334,In_29,In_24);
and U335 (N_335,In_879,In_1344);
xnor U336 (N_336,In_566,In_211);
or U337 (N_337,In_2,In_762);
nor U338 (N_338,In_1116,In_1377);
nand U339 (N_339,In_55,In_547);
and U340 (N_340,In_234,In_1380);
xnor U341 (N_341,In_513,In_1091);
and U342 (N_342,In_1374,In_549);
nand U343 (N_343,In_481,In_847);
and U344 (N_344,In_740,In_1184);
or U345 (N_345,In_707,In_156);
xnor U346 (N_346,In_644,In_1178);
or U347 (N_347,In_1367,In_500);
nand U348 (N_348,In_1346,In_983);
xnor U349 (N_349,In_848,In_838);
or U350 (N_350,In_650,In_1142);
xnor U351 (N_351,In_892,In_23);
nor U352 (N_352,In_641,In_426);
and U353 (N_353,In_695,In_255);
xnor U354 (N_354,In_400,In_63);
nor U355 (N_355,In_837,In_711);
nand U356 (N_356,In_341,In_937);
and U357 (N_357,In_1067,In_128);
nand U358 (N_358,In_768,In_970);
nor U359 (N_359,In_1229,In_274);
nor U360 (N_360,In_1114,In_1061);
nor U361 (N_361,In_567,In_902);
nand U362 (N_362,In_673,In_1411);
and U363 (N_363,In_1443,In_1183);
nand U364 (N_364,In_592,In_717);
xnor U365 (N_365,In_328,In_653);
or U366 (N_366,In_748,In_536);
nand U367 (N_367,In_1271,In_159);
or U368 (N_368,In_1180,In_741);
nor U369 (N_369,In_449,In_117);
nand U370 (N_370,In_1454,In_300);
and U371 (N_371,In_662,In_958);
nor U372 (N_372,In_35,In_191);
or U373 (N_373,In_1473,In_362);
or U374 (N_374,In_192,In_1263);
nor U375 (N_375,In_1402,In_971);
nand U376 (N_376,In_101,In_1188);
xor U377 (N_377,In_917,In_812);
and U378 (N_378,In_424,In_627);
or U379 (N_379,In_1149,In_1221);
nand U380 (N_380,In_89,In_1383);
xor U381 (N_381,In_754,In_1313);
nor U382 (N_382,In_639,In_222);
xnor U383 (N_383,In_1280,In_167);
or U384 (N_384,In_61,In_730);
or U385 (N_385,In_189,In_1281);
and U386 (N_386,In_556,In_445);
or U387 (N_387,In_859,In_1345);
nand U388 (N_388,In_484,In_450);
nand U389 (N_389,In_1336,In_336);
or U390 (N_390,In_771,In_190);
nor U391 (N_391,In_197,In_942);
xor U392 (N_392,In_1433,In_1410);
xnor U393 (N_393,In_469,In_311);
and U394 (N_394,In_1490,In_897);
and U395 (N_395,In_922,In_476);
nor U396 (N_396,In_261,In_772);
nor U397 (N_397,In_477,In_1434);
or U398 (N_398,In_260,In_799);
xor U399 (N_399,In_998,In_694);
nand U400 (N_400,In_130,In_385);
or U401 (N_401,In_1037,In_773);
nor U402 (N_402,In_141,In_616);
and U403 (N_403,In_702,In_858);
nor U404 (N_404,In_784,In_875);
xor U405 (N_405,In_817,In_1261);
or U406 (N_406,In_471,In_907);
nor U407 (N_407,In_723,In_350);
or U408 (N_408,In_473,In_1160);
nor U409 (N_409,In_1275,In_339);
nor U410 (N_410,In_1326,In_1308);
nor U411 (N_411,In_878,In_173);
nand U412 (N_412,In_1016,In_368);
xor U413 (N_413,In_1168,In_358);
or U414 (N_414,In_624,In_11);
or U415 (N_415,In_162,In_1203);
nor U416 (N_416,In_750,In_1375);
xor U417 (N_417,In_1404,In_1406);
nand U418 (N_418,In_1447,In_1471);
or U419 (N_419,In_1476,In_575);
nand U420 (N_420,In_1191,In_774);
and U421 (N_421,In_861,In_1150);
or U422 (N_422,In_108,In_1125);
nand U423 (N_423,In_890,In_1228);
nand U424 (N_424,In_543,In_766);
nand U425 (N_425,In_487,In_537);
xor U426 (N_426,In_1000,In_1187);
or U427 (N_427,In_927,In_394);
nor U428 (N_428,In_1086,In_572);
and U429 (N_429,In_1252,In_1487);
and U430 (N_430,In_686,In_1201);
nand U431 (N_431,In_1469,In_1393);
nand U432 (N_432,In_788,In_149);
nor U433 (N_433,In_1147,In_431);
xor U434 (N_434,In_256,In_1143);
nor U435 (N_435,In_629,In_975);
and U436 (N_436,In_1494,In_10);
xnor U437 (N_437,In_1195,In_488);
xnor U438 (N_438,In_1113,In_839);
or U439 (N_439,In_36,In_961);
nor U440 (N_440,In_501,In_395);
nor U441 (N_441,In_574,In_1235);
nand U442 (N_442,In_781,In_804);
nand U443 (N_443,In_1222,In_1090);
nand U444 (N_444,In_1070,In_389);
and U445 (N_445,In_794,In_375);
nand U446 (N_446,In_894,In_1355);
or U447 (N_447,In_676,In_405);
xor U448 (N_448,In_505,In_1213);
and U449 (N_449,In_831,In_124);
nor U450 (N_450,In_1432,In_672);
nand U451 (N_451,In_298,In_1084);
or U452 (N_452,In_492,In_511);
nor U453 (N_453,In_776,In_692);
and U454 (N_454,In_700,In_357);
xor U455 (N_455,In_1475,In_1072);
and U456 (N_456,In_557,In_1064);
nand U457 (N_457,In_636,In_862);
or U458 (N_458,In_125,In_28);
nand U459 (N_459,In_458,In_1414);
and U460 (N_460,In_26,In_272);
or U461 (N_461,In_373,In_661);
or U462 (N_462,In_419,In_923);
nand U463 (N_463,In_753,In_1004);
and U464 (N_464,In_973,In_1332);
or U465 (N_465,In_1451,In_1324);
and U466 (N_466,In_850,In_502);
and U467 (N_467,In_1157,In_308);
nor U468 (N_468,In_747,In_434);
xor U469 (N_469,In_310,In_40);
nand U470 (N_470,In_915,In_1021);
nand U471 (N_471,In_525,In_1240);
nand U472 (N_472,In_1074,In_713);
or U473 (N_473,In_340,In_1117);
nor U474 (N_474,In_246,In_194);
xor U475 (N_475,In_455,In_51);
nand U476 (N_476,In_764,In_99);
or U477 (N_477,In_982,In_908);
or U478 (N_478,In_1357,In_955);
or U479 (N_479,In_863,In_599);
and U480 (N_480,In_294,In_1289);
or U481 (N_481,In_1173,In_421);
and U482 (N_482,In_1436,In_1358);
nand U483 (N_483,In_523,In_1078);
nor U484 (N_484,In_446,In_1333);
and U485 (N_485,In_1119,In_38);
and U486 (N_486,In_1128,In_603);
and U487 (N_487,In_219,In_250);
nor U488 (N_488,In_1065,In_436);
xor U489 (N_489,In_529,In_127);
or U490 (N_490,In_281,In_1405);
xor U491 (N_491,In_1199,In_834);
xor U492 (N_492,In_377,In_214);
nor U493 (N_493,In_611,In_498);
nor U494 (N_494,In_617,In_1426);
or U495 (N_495,In_797,In_221);
nor U496 (N_496,In_1254,In_633);
nand U497 (N_497,In_1124,In_49);
nand U498 (N_498,In_137,In_1212);
xnor U499 (N_499,In_1013,In_726);
xnor U500 (N_500,In_325,In_657);
and U501 (N_501,In_1438,In_460);
and U502 (N_502,In_524,In_170);
or U503 (N_503,In_342,In_1388);
or U504 (N_504,In_555,In_1329);
xnor U505 (N_505,In_126,In_724);
nor U506 (N_506,In_521,In_887);
or U507 (N_507,In_856,In_1303);
and U508 (N_508,In_559,In_932);
nor U509 (N_509,In_1385,In_885);
nor U510 (N_510,In_459,In_1164);
nor U511 (N_511,In_402,In_652);
xor U512 (N_512,In_416,In_728);
and U513 (N_513,In_826,In_898);
nand U514 (N_514,In_1225,In_313);
xor U515 (N_515,In_554,In_146);
and U516 (N_516,In_1176,In_1044);
or U517 (N_517,In_909,In_936);
nor U518 (N_518,In_47,In_1012);
nand U519 (N_519,In_315,In_649);
and U520 (N_520,In_257,In_113);
nor U521 (N_521,In_1468,In_597);
and U522 (N_522,In_843,In_635);
and U523 (N_523,In_70,In_131);
nor U524 (N_524,In_732,In_230);
nor U525 (N_525,In_886,In_109);
and U526 (N_526,In_865,In_168);
xor U527 (N_527,In_33,In_701);
nor U528 (N_528,In_1311,In_64);
or U529 (N_529,In_1499,In_1020);
xnor U530 (N_530,In_155,In_106);
or U531 (N_531,In_541,In_816);
xnor U532 (N_532,In_841,In_948);
or U533 (N_533,In_407,In_945);
or U534 (N_534,In_1466,In_1285);
nor U535 (N_535,In_844,In_823);
xnor U536 (N_536,In_80,In_1441);
nor U537 (N_537,In_749,In_1041);
and U538 (N_538,In_602,In_725);
xnor U539 (N_539,In_1418,In_579);
nand U540 (N_540,In_1279,In_1455);
xor U541 (N_541,In_911,In_1153);
nand U542 (N_542,In_688,In_1241);
and U543 (N_543,In_946,In_474);
xor U544 (N_544,In_60,In_1081);
or U545 (N_545,In_576,In_320);
nor U546 (N_546,In_201,In_380);
and U547 (N_547,In_786,In_420);
nor U548 (N_548,In_266,In_775);
or U549 (N_549,In_651,In_712);
and U550 (N_550,In_355,In_1481);
nand U551 (N_551,In_1151,In_1382);
nor U552 (N_552,In_404,In_451);
nor U553 (N_553,In_836,In_1033);
xnor U554 (N_554,In_888,In_792);
and U555 (N_555,In_268,In_344);
and U556 (N_556,In_57,In_921);
nor U557 (N_557,In_352,In_709);
xnor U558 (N_558,In_46,In_95);
nand U559 (N_559,In_1420,In_132);
nand U560 (N_560,In_1089,In_370);
nand U561 (N_561,In_1052,In_427);
and U562 (N_562,In_1098,In_731);
and U563 (N_563,In_967,In_1445);
xnor U564 (N_564,In_1197,In_1400);
nor U565 (N_565,In_271,In_307);
nand U566 (N_566,In_348,In_1310);
or U567 (N_567,In_440,In_456);
nand U568 (N_568,In_1427,In_240);
and U569 (N_569,In_621,In_742);
xnor U570 (N_570,In_267,In_129);
or U571 (N_571,In_968,In_638);
and U572 (N_572,In_710,In_1483);
or U573 (N_573,In_1019,In_929);
or U574 (N_574,In_1082,In_997);
and U575 (N_575,In_1268,In_231);
xnor U576 (N_576,In_1068,In_1138);
or U577 (N_577,In_580,In_1477);
nand U578 (N_578,In_85,In_1442);
or U579 (N_579,In_551,In_437);
xor U580 (N_580,In_345,In_1444);
nor U581 (N_581,In_1276,In_1437);
xor U582 (N_582,In_461,In_869);
xor U583 (N_583,In_716,In_1224);
nand U584 (N_584,In_1368,In_432);
and U585 (N_585,In_1088,In_262);
nand U586 (N_586,In_757,In_678);
and U587 (N_587,In_1006,In_1076);
and U588 (N_588,In_905,In_415);
nor U589 (N_589,In_1278,In_1408);
nand U590 (N_590,In_1316,In_9);
and U591 (N_591,In_438,In_1424);
nand U592 (N_592,In_553,In_184);
or U593 (N_593,In_645,In_832);
and U594 (N_594,In_1460,In_1319);
nor U595 (N_595,In_1100,In_583);
xnor U596 (N_596,In_3,In_1039);
nand U597 (N_597,In_1370,In_486);
nand U598 (N_598,In_833,In_783);
nor U599 (N_599,In_1282,In_584);
nand U600 (N_600,In_111,In_1440);
xnor U601 (N_601,In_819,In_782);
or U602 (N_602,In_933,In_1430);
nor U603 (N_603,In_314,In_1115);
nand U604 (N_604,In_1340,In_291);
or U605 (N_605,In_643,In_655);
or U606 (N_606,In_199,In_163);
nand U607 (N_607,In_453,In_139);
nand U608 (N_608,In_912,In_302);
nor U609 (N_609,In_425,In_736);
nor U610 (N_610,In_1172,In_545);
and U611 (N_611,In_411,In_980);
nor U612 (N_612,In_988,In_956);
nand U613 (N_613,In_32,In_1399);
nor U614 (N_614,In_868,In_226);
xor U615 (N_615,In_67,In_925);
nor U616 (N_616,In_30,In_489);
and U617 (N_617,In_1472,In_1292);
and U618 (N_618,In_264,In_745);
and U619 (N_619,In_292,In_515);
or U620 (N_620,In_158,In_1120);
xnor U621 (N_621,In_322,In_102);
and U622 (N_622,In_338,In_277);
or U623 (N_623,In_319,In_188);
and U624 (N_624,In_417,In_118);
xnor U625 (N_625,In_1071,In_954);
and U626 (N_626,In_138,In_1087);
or U627 (N_627,In_1248,In_539);
or U628 (N_628,In_176,In_821);
nand U629 (N_629,In_366,In_254);
and U630 (N_630,In_828,In_950);
and U631 (N_631,In_376,In_1470);
and U632 (N_632,In_517,In_92);
nand U633 (N_633,In_1217,In_778);
nand U634 (N_634,In_248,In_1446);
or U635 (N_635,In_443,In_1127);
nor U636 (N_636,In_334,In_578);
or U637 (N_637,In_1453,In_1257);
nor U638 (N_638,In_777,In_873);
xor U639 (N_639,In_889,In_793);
and U640 (N_640,In_919,In_530);
nand U641 (N_641,In_999,In_74);
xnor U642 (N_642,In_1035,In_164);
xnor U643 (N_643,In_69,In_1264);
or U644 (N_644,In_349,In_883);
nand U645 (N_645,In_1107,In_1062);
and U646 (N_646,In_332,In_1231);
and U647 (N_647,In_71,In_467);
xnor U648 (N_648,In_227,In_337);
or U649 (N_649,In_283,In_1489);
xnor U650 (N_650,In_910,In_98);
or U651 (N_651,In_1055,In_1045);
or U652 (N_652,In_297,In_495);
nor U653 (N_653,In_369,In_654);
and U654 (N_654,In_317,In_802);
xor U655 (N_655,In_800,In_135);
or U656 (N_656,In_916,In_681);
nand U657 (N_657,In_981,In_1214);
nand U658 (N_658,In_259,In_951);
nand U659 (N_659,In_1139,In_1390);
xor U660 (N_660,In_1376,In_962);
or U661 (N_661,In_1314,In_829);
nand U662 (N_662,In_827,In_608);
or U663 (N_663,In_679,In_193);
nor U664 (N_664,In_642,In_1155);
and U665 (N_665,In_1140,In_22);
nand U666 (N_666,In_1027,In_504);
xnor U667 (N_667,In_1259,In_286);
nand U668 (N_668,In_31,In_1103);
or U669 (N_669,In_904,In_223);
or U670 (N_670,In_714,In_1111);
nor U671 (N_671,In_122,In_1096);
nor U672 (N_672,In_1492,In_202);
nand U673 (N_673,In_1154,In_241);
or U674 (N_674,In_560,In_568);
nand U675 (N_675,In_1244,In_114);
and U676 (N_676,In_622,In_1177);
xor U677 (N_677,In_926,In_383);
or U678 (N_678,In_1480,In_1048);
or U679 (N_679,In_952,In_1343);
xnor U680 (N_680,In_82,In_1194);
nand U681 (N_681,In_5,In_1118);
or U682 (N_682,In_1482,In_715);
and U683 (N_683,In_1236,In_588);
xnor U684 (N_684,In_1458,In_423);
nand U685 (N_685,In_1046,In_371);
or U686 (N_686,In_1106,In_1298);
or U687 (N_687,In_1208,In_941);
or U688 (N_688,In_1474,In_1266);
nor U689 (N_689,In_391,In_1137);
and U690 (N_690,In_1210,In_698);
nand U691 (N_691,In_258,In_430);
xnor U692 (N_692,In_1423,In_1233);
or U693 (N_693,In_229,In_759);
or U694 (N_694,In_290,In_808);
or U695 (N_695,In_722,In_154);
nand U696 (N_696,In_703,In_623);
or U697 (N_697,In_203,In_533);
xor U698 (N_698,In_1334,In_200);
xor U699 (N_699,In_1230,In_195);
nand U700 (N_700,In_1361,In_1286);
or U701 (N_701,In_1209,In_1227);
nor U702 (N_702,In_548,In_1130);
xnor U703 (N_703,In_1010,In_242);
nand U704 (N_704,In_670,In_153);
xor U705 (N_705,In_1095,In_571);
nor U706 (N_706,In_1097,In_145);
or U707 (N_707,In_552,In_1174);
nand U708 (N_708,In_960,In_807);
or U709 (N_709,In_1491,In_53);
xnor U710 (N_710,In_454,In_984);
xor U711 (N_711,In_668,In_1360);
xor U712 (N_712,In_735,In_1464);
xnor U713 (N_713,In_987,In_429);
or U714 (N_714,In_880,In_1307);
nor U715 (N_715,In_1014,In_1348);
nand U716 (N_716,In_483,In_236);
nand U717 (N_717,In_65,In_233);
xor U718 (N_718,In_1372,In_1159);
or U719 (N_719,In_14,In_1397);
nand U720 (N_720,In_590,In_790);
xor U721 (N_721,In_18,In_1005);
or U722 (N_722,In_465,In_1330);
xor U723 (N_723,In_463,In_1299);
nand U724 (N_724,In_88,In_1335);
and U725 (N_725,In_387,In_647);
nor U726 (N_726,In_1496,In_1034);
or U727 (N_727,In_120,In_1273);
nand U728 (N_728,In_805,In_165);
xor U729 (N_729,In_934,In_769);
xnor U730 (N_730,In_506,In_412);
and U731 (N_731,In_510,In_949);
nor U732 (N_732,In_41,In_327);
xor U733 (N_733,In_1,In_206);
and U734 (N_734,In_218,In_1145);
nor U735 (N_735,In_959,In_482);
and U736 (N_736,In_1122,In_690);
nand U737 (N_737,In_1165,In_160);
xor U738 (N_738,In_62,In_472);
xnor U739 (N_739,In_969,In_326);
nor U740 (N_740,In_903,In_1215);
xnor U741 (N_741,In_600,In_727);
nand U742 (N_742,In_867,In_86);
nand U743 (N_743,In_1258,In_399);
or U744 (N_744,In_27,In_739);
xor U745 (N_745,In_1431,In_648);
and U746 (N_746,In_228,In_864);
xor U747 (N_747,In_746,In_906);
nand U748 (N_748,In_1218,In_1093);
or U749 (N_749,In_180,In_1030);
nand U750 (N_750,In_1491,In_546);
nand U751 (N_751,In_1009,In_58);
nor U752 (N_752,In_106,In_262);
and U753 (N_753,In_533,In_450);
and U754 (N_754,In_1128,In_582);
nor U755 (N_755,In_123,In_597);
xnor U756 (N_756,In_571,In_1288);
or U757 (N_757,In_723,In_1160);
xnor U758 (N_758,In_590,In_3);
nor U759 (N_759,In_826,In_1310);
and U760 (N_760,In_752,In_224);
and U761 (N_761,In_517,In_655);
nand U762 (N_762,In_684,In_1063);
or U763 (N_763,In_1472,In_107);
and U764 (N_764,In_1382,In_314);
nor U765 (N_765,In_265,In_1408);
xnor U766 (N_766,In_1164,In_102);
nand U767 (N_767,In_421,In_1347);
and U768 (N_768,In_1208,In_1289);
and U769 (N_769,In_1163,In_251);
or U770 (N_770,In_833,In_1085);
xor U771 (N_771,In_1270,In_1110);
nor U772 (N_772,In_787,In_296);
and U773 (N_773,In_450,In_607);
or U774 (N_774,In_617,In_492);
xor U775 (N_775,In_1390,In_1343);
xnor U776 (N_776,In_171,In_951);
nand U777 (N_777,In_1268,In_893);
or U778 (N_778,In_296,In_149);
nand U779 (N_779,In_902,In_391);
xor U780 (N_780,In_277,In_992);
xor U781 (N_781,In_1029,In_2);
or U782 (N_782,In_799,In_102);
xor U783 (N_783,In_555,In_177);
nor U784 (N_784,In_146,In_0);
nor U785 (N_785,In_1205,In_735);
nand U786 (N_786,In_1239,In_96);
nand U787 (N_787,In_442,In_1239);
xor U788 (N_788,In_1160,In_478);
nor U789 (N_789,In_411,In_1445);
xnor U790 (N_790,In_502,In_1397);
xnor U791 (N_791,In_917,In_1256);
nor U792 (N_792,In_1355,In_200);
nand U793 (N_793,In_136,In_381);
or U794 (N_794,In_803,In_817);
nand U795 (N_795,In_357,In_983);
nand U796 (N_796,In_175,In_1211);
xor U797 (N_797,In_532,In_330);
xnor U798 (N_798,In_1119,In_620);
xor U799 (N_799,In_74,In_833);
nand U800 (N_800,In_1100,In_898);
nand U801 (N_801,In_510,In_1086);
nor U802 (N_802,In_940,In_1241);
and U803 (N_803,In_874,In_867);
and U804 (N_804,In_419,In_881);
nor U805 (N_805,In_1265,In_1060);
and U806 (N_806,In_226,In_61);
xnor U807 (N_807,In_1357,In_232);
or U808 (N_808,In_331,In_702);
nor U809 (N_809,In_773,In_154);
nand U810 (N_810,In_505,In_817);
xor U811 (N_811,In_1300,In_1112);
or U812 (N_812,In_988,In_9);
and U813 (N_813,In_99,In_1358);
xnor U814 (N_814,In_443,In_64);
xnor U815 (N_815,In_506,In_123);
xor U816 (N_816,In_1124,In_767);
or U817 (N_817,In_186,In_597);
and U818 (N_818,In_1137,In_449);
nor U819 (N_819,In_1152,In_1030);
and U820 (N_820,In_1185,In_396);
xnor U821 (N_821,In_296,In_832);
or U822 (N_822,In_431,In_296);
xnor U823 (N_823,In_1012,In_1429);
or U824 (N_824,In_1065,In_340);
xor U825 (N_825,In_251,In_351);
nor U826 (N_826,In_928,In_326);
and U827 (N_827,In_812,In_416);
nor U828 (N_828,In_1220,In_529);
and U829 (N_829,In_1408,In_614);
nor U830 (N_830,In_363,In_435);
nor U831 (N_831,In_822,In_1390);
nand U832 (N_832,In_216,In_59);
or U833 (N_833,In_1021,In_959);
nand U834 (N_834,In_1268,In_852);
and U835 (N_835,In_281,In_282);
xor U836 (N_836,In_1354,In_614);
or U837 (N_837,In_790,In_1034);
xor U838 (N_838,In_1277,In_1293);
and U839 (N_839,In_1450,In_839);
and U840 (N_840,In_695,In_1447);
or U841 (N_841,In_1482,In_67);
xnor U842 (N_842,In_1061,In_431);
and U843 (N_843,In_744,In_1286);
or U844 (N_844,In_987,In_547);
and U845 (N_845,In_266,In_1222);
nand U846 (N_846,In_793,In_829);
nand U847 (N_847,In_1393,In_731);
nand U848 (N_848,In_280,In_41);
xor U849 (N_849,In_1498,In_1441);
nor U850 (N_850,In_1365,In_1370);
or U851 (N_851,In_1055,In_806);
or U852 (N_852,In_501,In_1093);
nor U853 (N_853,In_679,In_1210);
xor U854 (N_854,In_686,In_266);
nand U855 (N_855,In_921,In_462);
nand U856 (N_856,In_726,In_1411);
nor U857 (N_857,In_309,In_565);
nor U858 (N_858,In_1391,In_351);
nor U859 (N_859,In_1446,In_1134);
or U860 (N_860,In_254,In_1100);
nand U861 (N_861,In_1305,In_703);
or U862 (N_862,In_1351,In_204);
xnor U863 (N_863,In_233,In_547);
or U864 (N_864,In_636,In_642);
or U865 (N_865,In_1109,In_964);
xnor U866 (N_866,In_1088,In_151);
or U867 (N_867,In_15,In_449);
or U868 (N_868,In_429,In_818);
nand U869 (N_869,In_1477,In_928);
nand U870 (N_870,In_1117,In_293);
nand U871 (N_871,In_327,In_914);
nand U872 (N_872,In_292,In_613);
xnor U873 (N_873,In_121,In_1437);
and U874 (N_874,In_1262,In_1255);
nor U875 (N_875,In_1065,In_991);
and U876 (N_876,In_602,In_1429);
nor U877 (N_877,In_1347,In_1278);
nor U878 (N_878,In_852,In_276);
or U879 (N_879,In_385,In_189);
nor U880 (N_880,In_1108,In_1063);
nor U881 (N_881,In_1206,In_243);
nand U882 (N_882,In_1426,In_762);
nand U883 (N_883,In_994,In_870);
nor U884 (N_884,In_1312,In_783);
xnor U885 (N_885,In_452,In_493);
or U886 (N_886,In_859,In_711);
nand U887 (N_887,In_1331,In_1414);
nand U888 (N_888,In_956,In_327);
nand U889 (N_889,In_933,In_1111);
and U890 (N_890,In_135,In_756);
and U891 (N_891,In_1321,In_1087);
and U892 (N_892,In_854,In_1230);
or U893 (N_893,In_1172,In_1421);
nor U894 (N_894,In_1188,In_475);
and U895 (N_895,In_686,In_812);
nand U896 (N_896,In_475,In_167);
or U897 (N_897,In_154,In_768);
xnor U898 (N_898,In_1326,In_1045);
nand U899 (N_899,In_1348,In_1239);
and U900 (N_900,In_66,In_1031);
nor U901 (N_901,In_1457,In_587);
nor U902 (N_902,In_273,In_711);
and U903 (N_903,In_890,In_882);
or U904 (N_904,In_163,In_462);
or U905 (N_905,In_850,In_1090);
xor U906 (N_906,In_624,In_1399);
and U907 (N_907,In_790,In_826);
xor U908 (N_908,In_1023,In_44);
and U909 (N_909,In_219,In_407);
nor U910 (N_910,In_34,In_1310);
and U911 (N_911,In_967,In_200);
nand U912 (N_912,In_50,In_152);
nor U913 (N_913,In_92,In_852);
xnor U914 (N_914,In_1142,In_552);
or U915 (N_915,In_1251,In_865);
or U916 (N_916,In_1197,In_573);
or U917 (N_917,In_1209,In_304);
and U918 (N_918,In_138,In_894);
xor U919 (N_919,In_247,In_48);
or U920 (N_920,In_382,In_808);
nand U921 (N_921,In_1310,In_53);
xor U922 (N_922,In_424,In_0);
nand U923 (N_923,In_667,In_1361);
or U924 (N_924,In_938,In_733);
or U925 (N_925,In_1155,In_427);
or U926 (N_926,In_138,In_55);
or U927 (N_927,In_796,In_1131);
nand U928 (N_928,In_1217,In_1294);
xor U929 (N_929,In_270,In_461);
xnor U930 (N_930,In_531,In_318);
nor U931 (N_931,In_380,In_748);
and U932 (N_932,In_1022,In_127);
and U933 (N_933,In_651,In_1414);
nand U934 (N_934,In_455,In_865);
nand U935 (N_935,In_1460,In_17);
and U936 (N_936,In_259,In_68);
and U937 (N_937,In_736,In_341);
xnor U938 (N_938,In_537,In_727);
and U939 (N_939,In_196,In_436);
or U940 (N_940,In_737,In_300);
nand U941 (N_941,In_180,In_1369);
or U942 (N_942,In_1140,In_1264);
nand U943 (N_943,In_927,In_786);
nand U944 (N_944,In_790,In_58);
or U945 (N_945,In_758,In_186);
nand U946 (N_946,In_354,In_87);
xor U947 (N_947,In_672,In_437);
nor U948 (N_948,In_187,In_1417);
nor U949 (N_949,In_735,In_408);
or U950 (N_950,In_1426,In_1310);
xnor U951 (N_951,In_514,In_742);
nor U952 (N_952,In_346,In_1035);
nor U953 (N_953,In_280,In_163);
nand U954 (N_954,In_157,In_1478);
and U955 (N_955,In_389,In_1275);
and U956 (N_956,In_1425,In_787);
or U957 (N_957,In_87,In_883);
and U958 (N_958,In_35,In_452);
and U959 (N_959,In_331,In_240);
nor U960 (N_960,In_198,In_583);
nor U961 (N_961,In_546,In_251);
or U962 (N_962,In_196,In_117);
or U963 (N_963,In_755,In_914);
nand U964 (N_964,In_1454,In_364);
nor U965 (N_965,In_279,In_672);
and U966 (N_966,In_1370,In_520);
nor U967 (N_967,In_1109,In_1461);
and U968 (N_968,In_613,In_354);
xnor U969 (N_969,In_1411,In_683);
and U970 (N_970,In_354,In_1086);
xnor U971 (N_971,In_358,In_452);
nor U972 (N_972,In_784,In_428);
and U973 (N_973,In_471,In_34);
nand U974 (N_974,In_24,In_650);
nor U975 (N_975,In_48,In_330);
xor U976 (N_976,In_1481,In_390);
and U977 (N_977,In_1038,In_144);
or U978 (N_978,In_1300,In_996);
or U979 (N_979,In_1417,In_1179);
or U980 (N_980,In_450,In_130);
xor U981 (N_981,In_1035,In_892);
and U982 (N_982,In_913,In_493);
or U983 (N_983,In_374,In_1079);
nor U984 (N_984,In_335,In_297);
xor U985 (N_985,In_1133,In_461);
xor U986 (N_986,In_1313,In_15);
xnor U987 (N_987,In_1169,In_428);
or U988 (N_988,In_854,In_42);
xor U989 (N_989,In_297,In_15);
or U990 (N_990,In_1164,In_763);
or U991 (N_991,In_1383,In_710);
and U992 (N_992,In_1240,In_509);
or U993 (N_993,In_1456,In_433);
nand U994 (N_994,In_1130,In_1355);
and U995 (N_995,In_205,In_1271);
nand U996 (N_996,In_149,In_53);
xnor U997 (N_997,In_750,In_478);
and U998 (N_998,In_582,In_818);
xor U999 (N_999,In_1424,In_203);
or U1000 (N_1000,In_381,In_1231);
nor U1001 (N_1001,In_1490,In_658);
nand U1002 (N_1002,In_960,In_1373);
and U1003 (N_1003,In_1317,In_1163);
or U1004 (N_1004,In_292,In_332);
nand U1005 (N_1005,In_552,In_825);
or U1006 (N_1006,In_208,In_1028);
nand U1007 (N_1007,In_302,In_1011);
and U1008 (N_1008,In_254,In_1218);
and U1009 (N_1009,In_776,In_86);
nand U1010 (N_1010,In_549,In_403);
nor U1011 (N_1011,In_1489,In_170);
xor U1012 (N_1012,In_1138,In_1071);
and U1013 (N_1013,In_748,In_189);
nand U1014 (N_1014,In_1339,In_1085);
xnor U1015 (N_1015,In_346,In_1457);
or U1016 (N_1016,In_1039,In_1377);
xor U1017 (N_1017,In_1180,In_303);
xnor U1018 (N_1018,In_1251,In_1409);
and U1019 (N_1019,In_953,In_1486);
xor U1020 (N_1020,In_1355,In_1140);
xor U1021 (N_1021,In_1169,In_947);
or U1022 (N_1022,In_1356,In_1264);
xnor U1023 (N_1023,In_781,In_255);
or U1024 (N_1024,In_1054,In_937);
or U1025 (N_1025,In_303,In_1244);
or U1026 (N_1026,In_355,In_1316);
or U1027 (N_1027,In_677,In_1264);
nor U1028 (N_1028,In_285,In_642);
and U1029 (N_1029,In_611,In_1491);
or U1030 (N_1030,In_230,In_771);
xor U1031 (N_1031,In_330,In_1128);
and U1032 (N_1032,In_1248,In_1003);
nor U1033 (N_1033,In_1256,In_111);
and U1034 (N_1034,In_330,In_1022);
xor U1035 (N_1035,In_1106,In_588);
or U1036 (N_1036,In_473,In_502);
nor U1037 (N_1037,In_117,In_765);
xnor U1038 (N_1038,In_928,In_159);
nor U1039 (N_1039,In_1327,In_438);
nand U1040 (N_1040,In_1402,In_1177);
and U1041 (N_1041,In_178,In_1089);
nand U1042 (N_1042,In_1194,In_648);
or U1043 (N_1043,In_373,In_1482);
nor U1044 (N_1044,In_1318,In_1433);
xor U1045 (N_1045,In_782,In_915);
or U1046 (N_1046,In_1403,In_436);
xor U1047 (N_1047,In_674,In_800);
nand U1048 (N_1048,In_1365,In_1187);
nand U1049 (N_1049,In_1273,In_1406);
or U1050 (N_1050,In_794,In_1224);
nand U1051 (N_1051,In_35,In_313);
or U1052 (N_1052,In_975,In_1452);
or U1053 (N_1053,In_538,In_563);
nand U1054 (N_1054,In_608,In_768);
nand U1055 (N_1055,In_1370,In_526);
or U1056 (N_1056,In_743,In_1250);
nor U1057 (N_1057,In_1097,In_453);
xnor U1058 (N_1058,In_294,In_1259);
and U1059 (N_1059,In_172,In_487);
nand U1060 (N_1060,In_1431,In_1397);
nor U1061 (N_1061,In_157,In_1367);
and U1062 (N_1062,In_1492,In_70);
and U1063 (N_1063,In_616,In_1213);
xnor U1064 (N_1064,In_1194,In_50);
nor U1065 (N_1065,In_989,In_181);
nor U1066 (N_1066,In_738,In_1050);
or U1067 (N_1067,In_54,In_1052);
xor U1068 (N_1068,In_1212,In_1277);
or U1069 (N_1069,In_1354,In_91);
xnor U1070 (N_1070,In_618,In_978);
xnor U1071 (N_1071,In_138,In_356);
or U1072 (N_1072,In_462,In_312);
xor U1073 (N_1073,In_161,In_1039);
nand U1074 (N_1074,In_1114,In_954);
nand U1075 (N_1075,In_662,In_63);
nand U1076 (N_1076,In_1466,In_214);
nand U1077 (N_1077,In_1221,In_573);
nor U1078 (N_1078,In_187,In_392);
or U1079 (N_1079,In_1075,In_449);
xnor U1080 (N_1080,In_876,In_438);
or U1081 (N_1081,In_886,In_1478);
nor U1082 (N_1082,In_948,In_1071);
nand U1083 (N_1083,In_82,In_788);
nand U1084 (N_1084,In_216,In_813);
nor U1085 (N_1085,In_649,In_173);
nor U1086 (N_1086,In_818,In_434);
or U1087 (N_1087,In_204,In_1249);
nor U1088 (N_1088,In_45,In_1457);
nand U1089 (N_1089,In_754,In_948);
xor U1090 (N_1090,In_658,In_1319);
or U1091 (N_1091,In_576,In_1326);
nand U1092 (N_1092,In_537,In_791);
nand U1093 (N_1093,In_40,In_901);
nand U1094 (N_1094,In_790,In_645);
nand U1095 (N_1095,In_7,In_328);
xnor U1096 (N_1096,In_472,In_1285);
xnor U1097 (N_1097,In_275,In_355);
nand U1098 (N_1098,In_260,In_592);
xnor U1099 (N_1099,In_1335,In_389);
nand U1100 (N_1100,In_884,In_1341);
nand U1101 (N_1101,In_698,In_735);
nand U1102 (N_1102,In_67,In_900);
or U1103 (N_1103,In_1424,In_814);
and U1104 (N_1104,In_943,In_263);
or U1105 (N_1105,In_178,In_256);
xnor U1106 (N_1106,In_575,In_1057);
nor U1107 (N_1107,In_1170,In_314);
xor U1108 (N_1108,In_12,In_1389);
nor U1109 (N_1109,In_1044,In_930);
xor U1110 (N_1110,In_59,In_505);
and U1111 (N_1111,In_1245,In_23);
or U1112 (N_1112,In_296,In_546);
xor U1113 (N_1113,In_1255,In_139);
xnor U1114 (N_1114,In_1421,In_503);
and U1115 (N_1115,In_733,In_815);
and U1116 (N_1116,In_880,In_1367);
or U1117 (N_1117,In_840,In_1029);
and U1118 (N_1118,In_1179,In_1434);
and U1119 (N_1119,In_1163,In_994);
or U1120 (N_1120,In_330,In_193);
nand U1121 (N_1121,In_810,In_1497);
nor U1122 (N_1122,In_562,In_82);
and U1123 (N_1123,In_745,In_112);
or U1124 (N_1124,In_1477,In_1180);
xor U1125 (N_1125,In_178,In_883);
nor U1126 (N_1126,In_639,In_903);
nor U1127 (N_1127,In_695,In_796);
xor U1128 (N_1128,In_69,In_922);
and U1129 (N_1129,In_895,In_728);
nor U1130 (N_1130,In_726,In_1410);
xnor U1131 (N_1131,In_174,In_391);
and U1132 (N_1132,In_594,In_126);
xnor U1133 (N_1133,In_363,In_490);
and U1134 (N_1134,In_1096,In_1088);
and U1135 (N_1135,In_385,In_207);
and U1136 (N_1136,In_746,In_1278);
or U1137 (N_1137,In_1351,In_621);
nor U1138 (N_1138,In_161,In_1071);
xnor U1139 (N_1139,In_1137,In_507);
nand U1140 (N_1140,In_1041,In_1474);
and U1141 (N_1141,In_192,In_34);
nand U1142 (N_1142,In_1427,In_1038);
or U1143 (N_1143,In_1380,In_1158);
xor U1144 (N_1144,In_900,In_961);
and U1145 (N_1145,In_748,In_1221);
xnor U1146 (N_1146,In_650,In_1275);
or U1147 (N_1147,In_759,In_747);
xnor U1148 (N_1148,In_1096,In_198);
nand U1149 (N_1149,In_262,In_380);
nand U1150 (N_1150,In_1360,In_1061);
or U1151 (N_1151,In_517,In_1146);
xnor U1152 (N_1152,In_39,In_830);
and U1153 (N_1153,In_80,In_492);
and U1154 (N_1154,In_215,In_1119);
or U1155 (N_1155,In_98,In_633);
nor U1156 (N_1156,In_167,In_943);
and U1157 (N_1157,In_1239,In_256);
nand U1158 (N_1158,In_773,In_1248);
nand U1159 (N_1159,In_123,In_210);
xor U1160 (N_1160,In_411,In_1408);
xnor U1161 (N_1161,In_709,In_1277);
and U1162 (N_1162,In_1095,In_1283);
or U1163 (N_1163,In_959,In_1497);
or U1164 (N_1164,In_993,In_1123);
nor U1165 (N_1165,In_1109,In_1462);
nand U1166 (N_1166,In_548,In_1210);
xor U1167 (N_1167,In_814,In_892);
nor U1168 (N_1168,In_1371,In_1477);
xor U1169 (N_1169,In_126,In_561);
and U1170 (N_1170,In_850,In_621);
nor U1171 (N_1171,In_1258,In_807);
and U1172 (N_1172,In_697,In_1405);
xnor U1173 (N_1173,In_599,In_1405);
xor U1174 (N_1174,In_549,In_195);
or U1175 (N_1175,In_323,In_813);
or U1176 (N_1176,In_291,In_512);
nor U1177 (N_1177,In_285,In_508);
or U1178 (N_1178,In_929,In_1079);
nand U1179 (N_1179,In_915,In_1092);
nand U1180 (N_1180,In_151,In_104);
xnor U1181 (N_1181,In_82,In_659);
nor U1182 (N_1182,In_776,In_771);
or U1183 (N_1183,In_1190,In_686);
xnor U1184 (N_1184,In_513,In_46);
nor U1185 (N_1185,In_323,In_1393);
xnor U1186 (N_1186,In_372,In_1005);
nand U1187 (N_1187,In_226,In_1153);
xnor U1188 (N_1188,In_42,In_823);
or U1189 (N_1189,In_200,In_620);
or U1190 (N_1190,In_90,In_908);
xor U1191 (N_1191,In_347,In_1143);
nand U1192 (N_1192,In_1109,In_667);
or U1193 (N_1193,In_201,In_300);
nor U1194 (N_1194,In_864,In_530);
xor U1195 (N_1195,In_314,In_205);
nand U1196 (N_1196,In_1300,In_1118);
and U1197 (N_1197,In_197,In_345);
and U1198 (N_1198,In_1247,In_948);
or U1199 (N_1199,In_1040,In_1239);
nand U1200 (N_1200,In_796,In_80);
and U1201 (N_1201,In_248,In_74);
and U1202 (N_1202,In_613,In_1290);
or U1203 (N_1203,In_1474,In_1140);
xnor U1204 (N_1204,In_125,In_86);
and U1205 (N_1205,In_618,In_579);
xor U1206 (N_1206,In_620,In_158);
nand U1207 (N_1207,In_731,In_1183);
and U1208 (N_1208,In_727,In_1034);
xor U1209 (N_1209,In_1405,In_679);
xor U1210 (N_1210,In_883,In_1394);
nand U1211 (N_1211,In_342,In_428);
and U1212 (N_1212,In_919,In_128);
nor U1213 (N_1213,In_954,In_1311);
nor U1214 (N_1214,In_118,In_1182);
nand U1215 (N_1215,In_1444,In_1269);
or U1216 (N_1216,In_1080,In_964);
nor U1217 (N_1217,In_374,In_548);
nor U1218 (N_1218,In_1403,In_319);
nand U1219 (N_1219,In_1416,In_1075);
or U1220 (N_1220,In_263,In_649);
and U1221 (N_1221,In_1484,In_280);
xnor U1222 (N_1222,In_781,In_1189);
xnor U1223 (N_1223,In_881,In_138);
or U1224 (N_1224,In_689,In_1494);
xor U1225 (N_1225,In_874,In_1186);
or U1226 (N_1226,In_1258,In_1001);
nand U1227 (N_1227,In_383,In_564);
or U1228 (N_1228,In_755,In_728);
nor U1229 (N_1229,In_837,In_130);
xor U1230 (N_1230,In_315,In_667);
nand U1231 (N_1231,In_465,In_672);
or U1232 (N_1232,In_529,In_1044);
xnor U1233 (N_1233,In_227,In_553);
and U1234 (N_1234,In_117,In_994);
nand U1235 (N_1235,In_279,In_839);
nor U1236 (N_1236,In_1336,In_1282);
xor U1237 (N_1237,In_1012,In_881);
nand U1238 (N_1238,In_358,In_1392);
and U1239 (N_1239,In_490,In_522);
nand U1240 (N_1240,In_1430,In_1161);
and U1241 (N_1241,In_708,In_1153);
nand U1242 (N_1242,In_1041,In_649);
nand U1243 (N_1243,In_1175,In_1128);
xor U1244 (N_1244,In_10,In_526);
nor U1245 (N_1245,In_408,In_1035);
and U1246 (N_1246,In_375,In_752);
nor U1247 (N_1247,In_118,In_1483);
or U1248 (N_1248,In_880,In_102);
or U1249 (N_1249,In_681,In_1469);
xor U1250 (N_1250,In_746,In_824);
nand U1251 (N_1251,In_1200,In_755);
nand U1252 (N_1252,In_851,In_1242);
nand U1253 (N_1253,In_1296,In_361);
xnor U1254 (N_1254,In_989,In_346);
nor U1255 (N_1255,In_272,In_224);
nor U1256 (N_1256,In_848,In_1047);
or U1257 (N_1257,In_142,In_798);
nor U1258 (N_1258,In_864,In_375);
and U1259 (N_1259,In_1109,In_1267);
nor U1260 (N_1260,In_400,In_836);
nor U1261 (N_1261,In_1439,In_19);
or U1262 (N_1262,In_895,In_1410);
nor U1263 (N_1263,In_691,In_265);
and U1264 (N_1264,In_1076,In_50);
nand U1265 (N_1265,In_408,In_1326);
or U1266 (N_1266,In_1114,In_1359);
nor U1267 (N_1267,In_747,In_141);
or U1268 (N_1268,In_1001,In_1264);
and U1269 (N_1269,In_1114,In_1381);
or U1270 (N_1270,In_275,In_916);
xnor U1271 (N_1271,In_844,In_112);
nand U1272 (N_1272,In_635,In_298);
or U1273 (N_1273,In_618,In_797);
and U1274 (N_1274,In_1062,In_1346);
xnor U1275 (N_1275,In_1300,In_808);
nand U1276 (N_1276,In_1255,In_477);
nand U1277 (N_1277,In_1306,In_1029);
or U1278 (N_1278,In_683,In_700);
nand U1279 (N_1279,In_1197,In_472);
nor U1280 (N_1280,In_803,In_4);
nor U1281 (N_1281,In_243,In_1461);
nand U1282 (N_1282,In_630,In_639);
or U1283 (N_1283,In_1439,In_672);
nor U1284 (N_1284,In_86,In_950);
xor U1285 (N_1285,In_1408,In_1126);
nand U1286 (N_1286,In_425,In_1009);
or U1287 (N_1287,In_1374,In_714);
nand U1288 (N_1288,In_318,In_485);
xor U1289 (N_1289,In_189,In_109);
nand U1290 (N_1290,In_1100,In_103);
and U1291 (N_1291,In_628,In_760);
or U1292 (N_1292,In_404,In_377);
nor U1293 (N_1293,In_904,In_836);
or U1294 (N_1294,In_662,In_405);
xnor U1295 (N_1295,In_903,In_219);
or U1296 (N_1296,In_542,In_1478);
xnor U1297 (N_1297,In_200,In_1008);
and U1298 (N_1298,In_802,In_1035);
nand U1299 (N_1299,In_758,In_335);
nor U1300 (N_1300,In_618,In_182);
nor U1301 (N_1301,In_765,In_222);
or U1302 (N_1302,In_956,In_678);
nor U1303 (N_1303,In_1379,In_708);
xnor U1304 (N_1304,In_58,In_1316);
or U1305 (N_1305,In_1244,In_688);
nand U1306 (N_1306,In_1185,In_453);
or U1307 (N_1307,In_381,In_1110);
xnor U1308 (N_1308,In_647,In_728);
or U1309 (N_1309,In_525,In_1104);
or U1310 (N_1310,In_408,In_1422);
nor U1311 (N_1311,In_512,In_339);
xnor U1312 (N_1312,In_339,In_1005);
nand U1313 (N_1313,In_339,In_112);
or U1314 (N_1314,In_1376,In_1068);
nor U1315 (N_1315,In_47,In_109);
nor U1316 (N_1316,In_761,In_45);
nor U1317 (N_1317,In_539,In_1394);
nand U1318 (N_1318,In_508,In_288);
and U1319 (N_1319,In_394,In_611);
and U1320 (N_1320,In_1064,In_921);
xor U1321 (N_1321,In_253,In_590);
nand U1322 (N_1322,In_725,In_179);
and U1323 (N_1323,In_311,In_1299);
nand U1324 (N_1324,In_534,In_1008);
nand U1325 (N_1325,In_1093,In_390);
and U1326 (N_1326,In_190,In_1471);
or U1327 (N_1327,In_826,In_4);
or U1328 (N_1328,In_483,In_886);
or U1329 (N_1329,In_650,In_263);
or U1330 (N_1330,In_651,In_1093);
or U1331 (N_1331,In_726,In_100);
and U1332 (N_1332,In_148,In_865);
nand U1333 (N_1333,In_1148,In_400);
and U1334 (N_1334,In_170,In_270);
or U1335 (N_1335,In_580,In_265);
nor U1336 (N_1336,In_883,In_717);
nand U1337 (N_1337,In_77,In_1031);
or U1338 (N_1338,In_1062,In_406);
nand U1339 (N_1339,In_343,In_1231);
and U1340 (N_1340,In_933,In_1140);
nand U1341 (N_1341,In_1053,In_1482);
nand U1342 (N_1342,In_481,In_796);
nor U1343 (N_1343,In_935,In_1334);
and U1344 (N_1344,In_107,In_1039);
or U1345 (N_1345,In_314,In_1066);
nor U1346 (N_1346,In_1400,In_701);
nand U1347 (N_1347,In_160,In_1219);
xnor U1348 (N_1348,In_1008,In_392);
or U1349 (N_1349,In_1078,In_704);
xnor U1350 (N_1350,In_592,In_736);
nor U1351 (N_1351,In_707,In_1159);
xnor U1352 (N_1352,In_343,In_1377);
nor U1353 (N_1353,In_482,In_1229);
or U1354 (N_1354,In_940,In_977);
or U1355 (N_1355,In_998,In_96);
or U1356 (N_1356,In_1089,In_368);
nor U1357 (N_1357,In_166,In_784);
and U1358 (N_1358,In_1462,In_1079);
or U1359 (N_1359,In_1,In_471);
or U1360 (N_1360,In_753,In_195);
and U1361 (N_1361,In_794,In_858);
xnor U1362 (N_1362,In_760,In_1265);
or U1363 (N_1363,In_158,In_1496);
xnor U1364 (N_1364,In_979,In_26);
and U1365 (N_1365,In_920,In_1304);
or U1366 (N_1366,In_842,In_1290);
nor U1367 (N_1367,In_1019,In_1375);
or U1368 (N_1368,In_937,In_1269);
or U1369 (N_1369,In_1344,In_1361);
xor U1370 (N_1370,In_608,In_1251);
or U1371 (N_1371,In_59,In_919);
and U1372 (N_1372,In_1318,In_1341);
and U1373 (N_1373,In_96,In_477);
nor U1374 (N_1374,In_776,In_1066);
xnor U1375 (N_1375,In_327,In_1085);
nand U1376 (N_1376,In_1110,In_1445);
xnor U1377 (N_1377,In_890,In_1209);
nand U1378 (N_1378,In_643,In_1474);
xor U1379 (N_1379,In_960,In_137);
xnor U1380 (N_1380,In_830,In_1333);
xnor U1381 (N_1381,In_323,In_1288);
nor U1382 (N_1382,In_279,In_1079);
xnor U1383 (N_1383,In_1494,In_691);
xor U1384 (N_1384,In_1476,In_1117);
or U1385 (N_1385,In_878,In_542);
and U1386 (N_1386,In_51,In_1319);
or U1387 (N_1387,In_1059,In_379);
and U1388 (N_1388,In_569,In_122);
and U1389 (N_1389,In_1179,In_1400);
or U1390 (N_1390,In_1062,In_1231);
or U1391 (N_1391,In_629,In_1038);
and U1392 (N_1392,In_1382,In_699);
nand U1393 (N_1393,In_1330,In_89);
xor U1394 (N_1394,In_1187,In_943);
nor U1395 (N_1395,In_639,In_473);
or U1396 (N_1396,In_13,In_1256);
nor U1397 (N_1397,In_1204,In_595);
or U1398 (N_1398,In_621,In_286);
xor U1399 (N_1399,In_417,In_687);
and U1400 (N_1400,In_1380,In_413);
or U1401 (N_1401,In_1127,In_865);
nor U1402 (N_1402,In_1254,In_368);
nor U1403 (N_1403,In_955,In_1167);
or U1404 (N_1404,In_121,In_1133);
and U1405 (N_1405,In_216,In_1475);
or U1406 (N_1406,In_1092,In_779);
xor U1407 (N_1407,In_453,In_1138);
nor U1408 (N_1408,In_688,In_1156);
xnor U1409 (N_1409,In_522,In_828);
nor U1410 (N_1410,In_220,In_509);
nand U1411 (N_1411,In_308,In_141);
nor U1412 (N_1412,In_681,In_558);
nor U1413 (N_1413,In_928,In_313);
nor U1414 (N_1414,In_23,In_131);
and U1415 (N_1415,In_288,In_603);
xor U1416 (N_1416,In_374,In_451);
nor U1417 (N_1417,In_1154,In_404);
or U1418 (N_1418,In_1073,In_1448);
xnor U1419 (N_1419,In_1166,In_628);
nor U1420 (N_1420,In_579,In_1493);
and U1421 (N_1421,In_502,In_207);
nor U1422 (N_1422,In_682,In_447);
or U1423 (N_1423,In_1283,In_820);
xnor U1424 (N_1424,In_990,In_311);
xor U1425 (N_1425,In_777,In_1311);
and U1426 (N_1426,In_1089,In_1212);
nor U1427 (N_1427,In_1244,In_921);
or U1428 (N_1428,In_1472,In_1039);
nand U1429 (N_1429,In_287,In_540);
xor U1430 (N_1430,In_1412,In_1043);
or U1431 (N_1431,In_299,In_134);
xnor U1432 (N_1432,In_1286,In_632);
xor U1433 (N_1433,In_271,In_1357);
nand U1434 (N_1434,In_11,In_501);
xor U1435 (N_1435,In_1221,In_28);
nand U1436 (N_1436,In_1359,In_978);
nor U1437 (N_1437,In_771,In_503);
xnor U1438 (N_1438,In_1419,In_852);
and U1439 (N_1439,In_971,In_825);
nand U1440 (N_1440,In_807,In_236);
or U1441 (N_1441,In_441,In_623);
and U1442 (N_1442,In_832,In_581);
and U1443 (N_1443,In_1223,In_364);
nor U1444 (N_1444,In_1055,In_737);
nor U1445 (N_1445,In_745,In_949);
xnor U1446 (N_1446,In_3,In_412);
nand U1447 (N_1447,In_176,In_856);
xnor U1448 (N_1448,In_430,In_558);
nand U1449 (N_1449,In_365,In_314);
nor U1450 (N_1450,In_312,In_956);
nand U1451 (N_1451,In_1143,In_274);
nand U1452 (N_1452,In_1019,In_1420);
and U1453 (N_1453,In_252,In_903);
and U1454 (N_1454,In_1111,In_1183);
or U1455 (N_1455,In_1117,In_228);
nand U1456 (N_1456,In_562,In_1489);
nor U1457 (N_1457,In_1336,In_79);
and U1458 (N_1458,In_1098,In_13);
nor U1459 (N_1459,In_76,In_972);
and U1460 (N_1460,In_1356,In_752);
xnor U1461 (N_1461,In_965,In_1210);
and U1462 (N_1462,In_430,In_1195);
and U1463 (N_1463,In_1382,In_311);
nor U1464 (N_1464,In_939,In_1129);
nand U1465 (N_1465,In_1094,In_98);
nand U1466 (N_1466,In_637,In_606);
xor U1467 (N_1467,In_1175,In_1123);
nor U1468 (N_1468,In_717,In_1428);
xor U1469 (N_1469,In_1348,In_751);
and U1470 (N_1470,In_208,In_458);
nand U1471 (N_1471,In_1487,In_448);
and U1472 (N_1472,In_7,In_1246);
nand U1473 (N_1473,In_1451,In_49);
nand U1474 (N_1474,In_1360,In_1342);
nor U1475 (N_1475,In_12,In_41);
nand U1476 (N_1476,In_1164,In_1320);
nor U1477 (N_1477,In_224,In_1140);
and U1478 (N_1478,In_719,In_966);
or U1479 (N_1479,In_1169,In_30);
nor U1480 (N_1480,In_1070,In_1145);
nand U1481 (N_1481,In_792,In_439);
and U1482 (N_1482,In_764,In_1039);
nand U1483 (N_1483,In_237,In_656);
or U1484 (N_1484,In_910,In_1152);
xnor U1485 (N_1485,In_692,In_181);
nor U1486 (N_1486,In_184,In_479);
nand U1487 (N_1487,In_1216,In_921);
or U1488 (N_1488,In_1220,In_359);
or U1489 (N_1489,In_1139,In_861);
or U1490 (N_1490,In_652,In_1162);
nor U1491 (N_1491,In_1110,In_1278);
and U1492 (N_1492,In_1031,In_1027);
nand U1493 (N_1493,In_1254,In_190);
xnor U1494 (N_1494,In_1188,In_1038);
nand U1495 (N_1495,In_942,In_1404);
xnor U1496 (N_1496,In_1252,In_826);
nor U1497 (N_1497,In_596,In_1436);
and U1498 (N_1498,In_556,In_1432);
and U1499 (N_1499,In_1027,In_345);
xnor U1500 (N_1500,In_14,In_147);
nor U1501 (N_1501,In_1388,In_116);
xor U1502 (N_1502,In_658,In_1204);
xnor U1503 (N_1503,In_1257,In_114);
nor U1504 (N_1504,In_744,In_316);
nor U1505 (N_1505,In_927,In_505);
nand U1506 (N_1506,In_878,In_928);
xnor U1507 (N_1507,In_1115,In_1396);
nand U1508 (N_1508,In_1170,In_1308);
nand U1509 (N_1509,In_1446,In_977);
xor U1510 (N_1510,In_801,In_825);
nor U1511 (N_1511,In_66,In_1105);
and U1512 (N_1512,In_1148,In_494);
nor U1513 (N_1513,In_974,In_443);
and U1514 (N_1514,In_316,In_1252);
and U1515 (N_1515,In_438,In_1034);
or U1516 (N_1516,In_1281,In_637);
nor U1517 (N_1517,In_961,In_997);
nor U1518 (N_1518,In_1168,In_190);
nor U1519 (N_1519,In_637,In_119);
nand U1520 (N_1520,In_352,In_880);
or U1521 (N_1521,In_1419,In_1442);
xor U1522 (N_1522,In_897,In_1108);
nand U1523 (N_1523,In_53,In_509);
and U1524 (N_1524,In_989,In_439);
or U1525 (N_1525,In_144,In_1309);
and U1526 (N_1526,In_96,In_1352);
and U1527 (N_1527,In_645,In_1426);
or U1528 (N_1528,In_1029,In_32);
nand U1529 (N_1529,In_307,In_1231);
xnor U1530 (N_1530,In_580,In_851);
xnor U1531 (N_1531,In_703,In_624);
and U1532 (N_1532,In_494,In_1089);
nor U1533 (N_1533,In_1480,In_15);
nor U1534 (N_1534,In_329,In_281);
and U1535 (N_1535,In_651,In_334);
or U1536 (N_1536,In_1201,In_799);
xnor U1537 (N_1537,In_649,In_236);
nand U1538 (N_1538,In_987,In_1296);
and U1539 (N_1539,In_1219,In_637);
and U1540 (N_1540,In_1106,In_322);
nor U1541 (N_1541,In_92,In_1065);
or U1542 (N_1542,In_1217,In_1020);
or U1543 (N_1543,In_94,In_685);
nor U1544 (N_1544,In_657,In_567);
nand U1545 (N_1545,In_1266,In_616);
xor U1546 (N_1546,In_203,In_1234);
and U1547 (N_1547,In_64,In_317);
nor U1548 (N_1548,In_632,In_723);
xor U1549 (N_1549,In_120,In_338);
or U1550 (N_1550,In_1446,In_675);
or U1551 (N_1551,In_1262,In_619);
xor U1552 (N_1552,In_544,In_328);
or U1553 (N_1553,In_604,In_1045);
nand U1554 (N_1554,In_339,In_474);
and U1555 (N_1555,In_1417,In_156);
nor U1556 (N_1556,In_632,In_519);
or U1557 (N_1557,In_660,In_681);
xor U1558 (N_1558,In_1345,In_376);
or U1559 (N_1559,In_512,In_35);
xor U1560 (N_1560,In_1271,In_624);
or U1561 (N_1561,In_1249,In_445);
and U1562 (N_1562,In_1463,In_101);
xor U1563 (N_1563,In_1124,In_553);
or U1564 (N_1564,In_1046,In_1197);
nand U1565 (N_1565,In_573,In_1103);
xor U1566 (N_1566,In_785,In_1101);
or U1567 (N_1567,In_1297,In_534);
and U1568 (N_1568,In_342,In_338);
xor U1569 (N_1569,In_819,In_523);
and U1570 (N_1570,In_807,In_973);
nand U1571 (N_1571,In_174,In_477);
and U1572 (N_1572,In_23,In_936);
or U1573 (N_1573,In_890,In_183);
and U1574 (N_1574,In_99,In_409);
or U1575 (N_1575,In_998,In_539);
and U1576 (N_1576,In_197,In_1027);
xnor U1577 (N_1577,In_579,In_672);
nand U1578 (N_1578,In_83,In_1320);
and U1579 (N_1579,In_753,In_1287);
nand U1580 (N_1580,In_388,In_246);
nor U1581 (N_1581,In_422,In_138);
or U1582 (N_1582,In_1427,In_646);
nor U1583 (N_1583,In_1495,In_277);
xnor U1584 (N_1584,In_922,In_1329);
xnor U1585 (N_1585,In_275,In_259);
or U1586 (N_1586,In_1455,In_549);
nor U1587 (N_1587,In_1443,In_577);
nor U1588 (N_1588,In_929,In_230);
nor U1589 (N_1589,In_367,In_943);
nand U1590 (N_1590,In_40,In_255);
xor U1591 (N_1591,In_1207,In_755);
or U1592 (N_1592,In_1242,In_584);
or U1593 (N_1593,In_1341,In_872);
and U1594 (N_1594,In_758,In_1372);
xor U1595 (N_1595,In_272,In_260);
or U1596 (N_1596,In_1078,In_17);
nor U1597 (N_1597,In_948,In_434);
and U1598 (N_1598,In_1363,In_531);
nor U1599 (N_1599,In_606,In_1033);
and U1600 (N_1600,In_331,In_770);
nand U1601 (N_1601,In_1376,In_158);
or U1602 (N_1602,In_73,In_759);
and U1603 (N_1603,In_1211,In_1094);
xnor U1604 (N_1604,In_334,In_144);
xor U1605 (N_1605,In_658,In_802);
nand U1606 (N_1606,In_670,In_1079);
nor U1607 (N_1607,In_684,In_83);
nor U1608 (N_1608,In_673,In_518);
nand U1609 (N_1609,In_57,In_1240);
nor U1610 (N_1610,In_1120,In_1143);
or U1611 (N_1611,In_485,In_301);
or U1612 (N_1612,In_1298,In_970);
nor U1613 (N_1613,In_1062,In_1359);
or U1614 (N_1614,In_412,In_33);
or U1615 (N_1615,In_1148,In_685);
and U1616 (N_1616,In_1130,In_105);
or U1617 (N_1617,In_869,In_983);
and U1618 (N_1618,In_260,In_1381);
nor U1619 (N_1619,In_235,In_88);
and U1620 (N_1620,In_789,In_1417);
nand U1621 (N_1621,In_14,In_530);
xnor U1622 (N_1622,In_1433,In_1476);
nor U1623 (N_1623,In_1090,In_958);
nor U1624 (N_1624,In_904,In_163);
xor U1625 (N_1625,In_20,In_287);
and U1626 (N_1626,In_97,In_905);
nor U1627 (N_1627,In_303,In_1273);
nand U1628 (N_1628,In_993,In_559);
nand U1629 (N_1629,In_757,In_595);
nand U1630 (N_1630,In_1117,In_75);
nor U1631 (N_1631,In_957,In_740);
and U1632 (N_1632,In_1075,In_37);
nand U1633 (N_1633,In_1362,In_949);
nor U1634 (N_1634,In_776,In_456);
nor U1635 (N_1635,In_73,In_1014);
xnor U1636 (N_1636,In_268,In_616);
or U1637 (N_1637,In_528,In_1078);
nand U1638 (N_1638,In_1102,In_298);
and U1639 (N_1639,In_268,In_157);
nor U1640 (N_1640,In_476,In_1121);
or U1641 (N_1641,In_1019,In_102);
xor U1642 (N_1642,In_1223,In_1087);
nor U1643 (N_1643,In_1009,In_1322);
nor U1644 (N_1644,In_1123,In_199);
or U1645 (N_1645,In_829,In_1409);
or U1646 (N_1646,In_378,In_1043);
or U1647 (N_1647,In_889,In_1333);
or U1648 (N_1648,In_835,In_1091);
and U1649 (N_1649,In_578,In_1160);
xor U1650 (N_1650,In_1182,In_319);
xor U1651 (N_1651,In_592,In_598);
nand U1652 (N_1652,In_426,In_873);
nor U1653 (N_1653,In_232,In_785);
nand U1654 (N_1654,In_1408,In_1073);
nand U1655 (N_1655,In_1120,In_1124);
nand U1656 (N_1656,In_913,In_981);
xor U1657 (N_1657,In_1362,In_1375);
and U1658 (N_1658,In_979,In_1057);
nor U1659 (N_1659,In_139,In_1347);
or U1660 (N_1660,In_1005,In_379);
or U1661 (N_1661,In_237,In_184);
or U1662 (N_1662,In_670,In_511);
nor U1663 (N_1663,In_585,In_385);
and U1664 (N_1664,In_188,In_1249);
nand U1665 (N_1665,In_1362,In_581);
nand U1666 (N_1666,In_1074,In_749);
xor U1667 (N_1667,In_427,In_902);
xor U1668 (N_1668,In_1402,In_1421);
nand U1669 (N_1669,In_1183,In_861);
nand U1670 (N_1670,In_296,In_594);
or U1671 (N_1671,In_1257,In_1477);
and U1672 (N_1672,In_1368,In_485);
and U1673 (N_1673,In_486,In_162);
nand U1674 (N_1674,In_1026,In_1325);
xnor U1675 (N_1675,In_775,In_333);
nor U1676 (N_1676,In_426,In_182);
and U1677 (N_1677,In_1261,In_1450);
or U1678 (N_1678,In_822,In_825);
or U1679 (N_1679,In_1045,In_203);
or U1680 (N_1680,In_158,In_256);
nand U1681 (N_1681,In_432,In_1392);
nand U1682 (N_1682,In_505,In_1284);
and U1683 (N_1683,In_914,In_535);
nand U1684 (N_1684,In_738,In_1124);
nor U1685 (N_1685,In_565,In_876);
nor U1686 (N_1686,In_1064,In_1200);
nor U1687 (N_1687,In_921,In_1189);
or U1688 (N_1688,In_868,In_1474);
nand U1689 (N_1689,In_1161,In_176);
xnor U1690 (N_1690,In_457,In_1369);
nand U1691 (N_1691,In_478,In_838);
xor U1692 (N_1692,In_1463,In_338);
nor U1693 (N_1693,In_564,In_276);
xor U1694 (N_1694,In_185,In_127);
nand U1695 (N_1695,In_138,In_603);
or U1696 (N_1696,In_1298,In_55);
xnor U1697 (N_1697,In_311,In_793);
nand U1698 (N_1698,In_450,In_764);
and U1699 (N_1699,In_94,In_295);
and U1700 (N_1700,In_206,In_890);
nand U1701 (N_1701,In_428,In_656);
nand U1702 (N_1702,In_953,In_1201);
nand U1703 (N_1703,In_733,In_551);
or U1704 (N_1704,In_1425,In_525);
nand U1705 (N_1705,In_682,In_115);
nand U1706 (N_1706,In_71,In_97);
xnor U1707 (N_1707,In_1235,In_412);
nand U1708 (N_1708,In_416,In_1257);
xor U1709 (N_1709,In_794,In_675);
nor U1710 (N_1710,In_1254,In_356);
xnor U1711 (N_1711,In_750,In_484);
nor U1712 (N_1712,In_554,In_1159);
xnor U1713 (N_1713,In_603,In_1483);
or U1714 (N_1714,In_528,In_1105);
and U1715 (N_1715,In_916,In_1420);
xor U1716 (N_1716,In_987,In_17);
or U1717 (N_1717,In_1312,In_83);
or U1718 (N_1718,In_802,In_213);
and U1719 (N_1719,In_686,In_1312);
xnor U1720 (N_1720,In_1168,In_1128);
nor U1721 (N_1721,In_1380,In_977);
or U1722 (N_1722,In_196,In_1142);
and U1723 (N_1723,In_726,In_1276);
nand U1724 (N_1724,In_641,In_89);
nand U1725 (N_1725,In_761,In_800);
nor U1726 (N_1726,In_97,In_182);
nand U1727 (N_1727,In_144,In_1061);
or U1728 (N_1728,In_1135,In_664);
and U1729 (N_1729,In_837,In_836);
or U1730 (N_1730,In_642,In_63);
or U1731 (N_1731,In_1261,In_1156);
and U1732 (N_1732,In_23,In_400);
or U1733 (N_1733,In_291,In_1200);
xor U1734 (N_1734,In_1063,In_1135);
or U1735 (N_1735,In_273,In_1441);
nand U1736 (N_1736,In_753,In_1108);
nor U1737 (N_1737,In_161,In_368);
nor U1738 (N_1738,In_935,In_272);
and U1739 (N_1739,In_1042,In_69);
nor U1740 (N_1740,In_45,In_1478);
nand U1741 (N_1741,In_878,In_255);
nor U1742 (N_1742,In_23,In_683);
and U1743 (N_1743,In_1061,In_810);
xnor U1744 (N_1744,In_1096,In_507);
or U1745 (N_1745,In_1498,In_521);
nand U1746 (N_1746,In_779,In_459);
nor U1747 (N_1747,In_1208,In_205);
nand U1748 (N_1748,In_933,In_1285);
or U1749 (N_1749,In_937,In_370);
nand U1750 (N_1750,In_165,In_106);
and U1751 (N_1751,In_1071,In_1463);
nor U1752 (N_1752,In_1174,In_191);
nor U1753 (N_1753,In_946,In_1309);
nand U1754 (N_1754,In_1154,In_625);
or U1755 (N_1755,In_501,In_65);
and U1756 (N_1756,In_396,In_36);
nand U1757 (N_1757,In_450,In_265);
or U1758 (N_1758,In_454,In_199);
nor U1759 (N_1759,In_684,In_63);
nand U1760 (N_1760,In_248,In_307);
xor U1761 (N_1761,In_214,In_1015);
or U1762 (N_1762,In_1143,In_267);
xnor U1763 (N_1763,In_660,In_800);
nor U1764 (N_1764,In_477,In_1081);
and U1765 (N_1765,In_1098,In_795);
or U1766 (N_1766,In_528,In_370);
or U1767 (N_1767,In_986,In_228);
nand U1768 (N_1768,In_1170,In_55);
and U1769 (N_1769,In_458,In_528);
or U1770 (N_1770,In_705,In_300);
or U1771 (N_1771,In_469,In_1439);
or U1772 (N_1772,In_468,In_1159);
nor U1773 (N_1773,In_777,In_282);
nor U1774 (N_1774,In_1287,In_18);
xnor U1775 (N_1775,In_412,In_1024);
xnor U1776 (N_1776,In_834,In_612);
nand U1777 (N_1777,In_139,In_154);
nand U1778 (N_1778,In_1386,In_176);
and U1779 (N_1779,In_43,In_1366);
or U1780 (N_1780,In_333,In_1234);
nor U1781 (N_1781,In_982,In_1419);
nor U1782 (N_1782,In_1297,In_975);
and U1783 (N_1783,In_300,In_118);
or U1784 (N_1784,In_558,In_1441);
xnor U1785 (N_1785,In_201,In_1299);
and U1786 (N_1786,In_1250,In_628);
nand U1787 (N_1787,In_1322,In_1191);
or U1788 (N_1788,In_716,In_1361);
and U1789 (N_1789,In_1016,In_565);
and U1790 (N_1790,In_1342,In_202);
nand U1791 (N_1791,In_1458,In_266);
or U1792 (N_1792,In_939,In_681);
or U1793 (N_1793,In_1277,In_730);
xnor U1794 (N_1794,In_296,In_1070);
nand U1795 (N_1795,In_366,In_1455);
xor U1796 (N_1796,In_14,In_1395);
or U1797 (N_1797,In_1245,In_1047);
nor U1798 (N_1798,In_114,In_1154);
or U1799 (N_1799,In_550,In_545);
xnor U1800 (N_1800,In_1378,In_1152);
and U1801 (N_1801,In_1359,In_863);
nor U1802 (N_1802,In_1349,In_1317);
or U1803 (N_1803,In_1074,In_677);
and U1804 (N_1804,In_829,In_1141);
or U1805 (N_1805,In_121,In_1455);
xor U1806 (N_1806,In_393,In_1303);
or U1807 (N_1807,In_1165,In_1429);
and U1808 (N_1808,In_692,In_1307);
nor U1809 (N_1809,In_577,In_155);
nand U1810 (N_1810,In_64,In_583);
or U1811 (N_1811,In_219,In_235);
and U1812 (N_1812,In_730,In_1008);
nor U1813 (N_1813,In_1012,In_1332);
nor U1814 (N_1814,In_568,In_1222);
and U1815 (N_1815,In_359,In_720);
or U1816 (N_1816,In_447,In_169);
or U1817 (N_1817,In_508,In_1356);
nor U1818 (N_1818,In_268,In_478);
xor U1819 (N_1819,In_295,In_522);
or U1820 (N_1820,In_1316,In_1256);
and U1821 (N_1821,In_191,In_1435);
nor U1822 (N_1822,In_76,In_1422);
xor U1823 (N_1823,In_350,In_629);
or U1824 (N_1824,In_877,In_389);
nand U1825 (N_1825,In_891,In_453);
nand U1826 (N_1826,In_76,In_561);
and U1827 (N_1827,In_119,In_360);
nor U1828 (N_1828,In_718,In_944);
xnor U1829 (N_1829,In_335,In_962);
nand U1830 (N_1830,In_716,In_576);
xnor U1831 (N_1831,In_624,In_93);
nand U1832 (N_1832,In_574,In_152);
nor U1833 (N_1833,In_1179,In_439);
nor U1834 (N_1834,In_786,In_937);
nor U1835 (N_1835,In_928,In_1287);
or U1836 (N_1836,In_589,In_1111);
and U1837 (N_1837,In_436,In_202);
or U1838 (N_1838,In_1135,In_758);
or U1839 (N_1839,In_311,In_1245);
nand U1840 (N_1840,In_502,In_587);
or U1841 (N_1841,In_1484,In_628);
nand U1842 (N_1842,In_1075,In_1335);
xnor U1843 (N_1843,In_1212,In_51);
xor U1844 (N_1844,In_1204,In_1448);
nor U1845 (N_1845,In_183,In_1423);
or U1846 (N_1846,In_1249,In_921);
nor U1847 (N_1847,In_42,In_825);
nand U1848 (N_1848,In_578,In_1043);
xor U1849 (N_1849,In_62,In_1443);
nand U1850 (N_1850,In_616,In_71);
and U1851 (N_1851,In_294,In_633);
and U1852 (N_1852,In_249,In_1010);
nor U1853 (N_1853,In_9,In_787);
nor U1854 (N_1854,In_1163,In_1383);
nand U1855 (N_1855,In_278,In_1410);
or U1856 (N_1856,In_1195,In_529);
nor U1857 (N_1857,In_111,In_53);
nand U1858 (N_1858,In_381,In_370);
nand U1859 (N_1859,In_1237,In_730);
and U1860 (N_1860,In_733,In_870);
or U1861 (N_1861,In_740,In_1034);
xnor U1862 (N_1862,In_119,In_1136);
or U1863 (N_1863,In_1427,In_598);
nand U1864 (N_1864,In_735,In_832);
or U1865 (N_1865,In_1414,In_685);
or U1866 (N_1866,In_704,In_125);
nand U1867 (N_1867,In_1438,In_219);
or U1868 (N_1868,In_1040,In_696);
nand U1869 (N_1869,In_933,In_350);
and U1870 (N_1870,In_1367,In_1430);
nor U1871 (N_1871,In_740,In_787);
nand U1872 (N_1872,In_277,In_898);
nand U1873 (N_1873,In_454,In_1133);
nand U1874 (N_1874,In_185,In_979);
and U1875 (N_1875,In_487,In_817);
xor U1876 (N_1876,In_1460,In_1222);
and U1877 (N_1877,In_1396,In_267);
nor U1878 (N_1878,In_586,In_1001);
xor U1879 (N_1879,In_890,In_1454);
xor U1880 (N_1880,In_1109,In_208);
nor U1881 (N_1881,In_192,In_1224);
nand U1882 (N_1882,In_199,In_143);
xor U1883 (N_1883,In_1482,In_519);
xnor U1884 (N_1884,In_923,In_1245);
or U1885 (N_1885,In_186,In_1221);
nand U1886 (N_1886,In_550,In_1406);
xnor U1887 (N_1887,In_724,In_999);
or U1888 (N_1888,In_183,In_328);
and U1889 (N_1889,In_1344,In_489);
nor U1890 (N_1890,In_966,In_872);
nor U1891 (N_1891,In_472,In_1291);
nor U1892 (N_1892,In_86,In_1257);
xor U1893 (N_1893,In_1387,In_1112);
and U1894 (N_1894,In_169,In_839);
and U1895 (N_1895,In_1244,In_1371);
nand U1896 (N_1896,In_142,In_1230);
or U1897 (N_1897,In_1387,In_1408);
nand U1898 (N_1898,In_1110,In_542);
and U1899 (N_1899,In_1122,In_256);
nand U1900 (N_1900,In_1074,In_1343);
nor U1901 (N_1901,In_524,In_808);
nor U1902 (N_1902,In_973,In_862);
xnor U1903 (N_1903,In_1378,In_1040);
nand U1904 (N_1904,In_846,In_110);
or U1905 (N_1905,In_663,In_967);
or U1906 (N_1906,In_1103,In_1151);
nand U1907 (N_1907,In_501,In_165);
nor U1908 (N_1908,In_688,In_485);
nand U1909 (N_1909,In_691,In_125);
and U1910 (N_1910,In_347,In_388);
xor U1911 (N_1911,In_899,In_169);
or U1912 (N_1912,In_560,In_1451);
nand U1913 (N_1913,In_1309,In_160);
xor U1914 (N_1914,In_1198,In_1181);
nand U1915 (N_1915,In_1379,In_987);
nor U1916 (N_1916,In_313,In_122);
nand U1917 (N_1917,In_1286,In_1391);
nor U1918 (N_1918,In_1476,In_567);
or U1919 (N_1919,In_91,In_232);
nand U1920 (N_1920,In_741,In_228);
and U1921 (N_1921,In_46,In_910);
or U1922 (N_1922,In_1169,In_774);
and U1923 (N_1923,In_281,In_140);
or U1924 (N_1924,In_233,In_259);
nor U1925 (N_1925,In_437,In_756);
xor U1926 (N_1926,In_20,In_64);
xnor U1927 (N_1927,In_624,In_923);
nor U1928 (N_1928,In_976,In_1377);
nor U1929 (N_1929,In_986,In_254);
xor U1930 (N_1930,In_1091,In_448);
or U1931 (N_1931,In_592,In_1262);
and U1932 (N_1932,In_718,In_729);
and U1933 (N_1933,In_602,In_989);
nor U1934 (N_1934,In_416,In_301);
or U1935 (N_1935,In_1285,In_155);
nor U1936 (N_1936,In_635,In_964);
and U1937 (N_1937,In_330,In_1490);
or U1938 (N_1938,In_212,In_773);
xor U1939 (N_1939,In_500,In_345);
nor U1940 (N_1940,In_828,In_930);
and U1941 (N_1941,In_421,In_79);
nand U1942 (N_1942,In_340,In_44);
nand U1943 (N_1943,In_256,In_1124);
xor U1944 (N_1944,In_522,In_427);
and U1945 (N_1945,In_869,In_98);
xnor U1946 (N_1946,In_1329,In_360);
and U1947 (N_1947,In_1111,In_1001);
nand U1948 (N_1948,In_349,In_398);
nand U1949 (N_1949,In_1193,In_533);
nor U1950 (N_1950,In_701,In_466);
and U1951 (N_1951,In_538,In_424);
and U1952 (N_1952,In_152,In_1457);
nor U1953 (N_1953,In_245,In_90);
nand U1954 (N_1954,In_318,In_426);
xor U1955 (N_1955,In_256,In_1155);
nor U1956 (N_1956,In_1410,In_723);
nor U1957 (N_1957,In_347,In_896);
nor U1958 (N_1958,In_1462,In_1168);
xor U1959 (N_1959,In_881,In_989);
nor U1960 (N_1960,In_1173,In_395);
or U1961 (N_1961,In_1358,In_1424);
nor U1962 (N_1962,In_0,In_1385);
and U1963 (N_1963,In_1474,In_1068);
nand U1964 (N_1964,In_1156,In_60);
xor U1965 (N_1965,In_1336,In_739);
or U1966 (N_1966,In_442,In_1040);
nand U1967 (N_1967,In_467,In_522);
nor U1968 (N_1968,In_929,In_1039);
nand U1969 (N_1969,In_9,In_562);
nand U1970 (N_1970,In_1469,In_364);
nand U1971 (N_1971,In_1199,In_388);
nor U1972 (N_1972,In_427,In_28);
xor U1973 (N_1973,In_470,In_582);
xor U1974 (N_1974,In_1061,In_1412);
nand U1975 (N_1975,In_1225,In_945);
nand U1976 (N_1976,In_756,In_783);
or U1977 (N_1977,In_302,In_347);
xnor U1978 (N_1978,In_742,In_1317);
or U1979 (N_1979,In_1264,In_778);
nand U1980 (N_1980,In_681,In_514);
and U1981 (N_1981,In_429,In_833);
xor U1982 (N_1982,In_944,In_1145);
and U1983 (N_1983,In_1469,In_881);
or U1984 (N_1984,In_61,In_907);
or U1985 (N_1985,In_476,In_172);
nor U1986 (N_1986,In_1421,In_122);
nor U1987 (N_1987,In_1023,In_511);
xnor U1988 (N_1988,In_807,In_1282);
nand U1989 (N_1989,In_229,In_193);
or U1990 (N_1990,In_91,In_43);
xnor U1991 (N_1991,In_945,In_330);
or U1992 (N_1992,In_1001,In_591);
xor U1993 (N_1993,In_677,In_1421);
or U1994 (N_1994,In_925,In_367);
and U1995 (N_1995,In_116,In_565);
or U1996 (N_1996,In_372,In_967);
and U1997 (N_1997,In_372,In_601);
and U1998 (N_1998,In_285,In_1304);
or U1999 (N_1999,In_27,In_439);
and U2000 (N_2000,In_464,In_510);
and U2001 (N_2001,In_1058,In_1305);
nand U2002 (N_2002,In_1453,In_809);
and U2003 (N_2003,In_1076,In_1197);
nand U2004 (N_2004,In_1385,In_60);
or U2005 (N_2005,In_1321,In_294);
xor U2006 (N_2006,In_751,In_790);
nor U2007 (N_2007,In_1383,In_1187);
xor U2008 (N_2008,In_1401,In_498);
nor U2009 (N_2009,In_1440,In_190);
or U2010 (N_2010,In_436,In_701);
xor U2011 (N_2011,In_104,In_1227);
nand U2012 (N_2012,In_1088,In_753);
nand U2013 (N_2013,In_1004,In_29);
nand U2014 (N_2014,In_879,In_353);
nor U2015 (N_2015,In_259,In_613);
nor U2016 (N_2016,In_236,In_337);
or U2017 (N_2017,In_690,In_1331);
nand U2018 (N_2018,In_292,In_984);
xnor U2019 (N_2019,In_1412,In_603);
xnor U2020 (N_2020,In_669,In_1268);
nor U2021 (N_2021,In_179,In_1304);
xnor U2022 (N_2022,In_1312,In_614);
xnor U2023 (N_2023,In_738,In_1321);
nor U2024 (N_2024,In_175,In_435);
nor U2025 (N_2025,In_79,In_64);
xnor U2026 (N_2026,In_1440,In_91);
or U2027 (N_2027,In_959,In_1344);
nor U2028 (N_2028,In_1097,In_1131);
and U2029 (N_2029,In_625,In_741);
and U2030 (N_2030,In_1268,In_141);
nor U2031 (N_2031,In_823,In_955);
nand U2032 (N_2032,In_812,In_1072);
and U2033 (N_2033,In_485,In_1414);
nor U2034 (N_2034,In_531,In_1205);
nand U2035 (N_2035,In_1005,In_1352);
or U2036 (N_2036,In_1354,In_277);
nor U2037 (N_2037,In_659,In_256);
nand U2038 (N_2038,In_950,In_471);
nand U2039 (N_2039,In_1489,In_542);
nand U2040 (N_2040,In_740,In_70);
nor U2041 (N_2041,In_1380,In_1056);
nand U2042 (N_2042,In_1318,In_587);
or U2043 (N_2043,In_189,In_1070);
and U2044 (N_2044,In_866,In_240);
or U2045 (N_2045,In_1298,In_222);
and U2046 (N_2046,In_1028,In_483);
nor U2047 (N_2047,In_600,In_965);
xor U2048 (N_2048,In_115,In_995);
xnor U2049 (N_2049,In_1259,In_1326);
and U2050 (N_2050,In_1250,In_508);
and U2051 (N_2051,In_225,In_542);
xnor U2052 (N_2052,In_284,In_200);
xnor U2053 (N_2053,In_515,In_1116);
nand U2054 (N_2054,In_144,In_1283);
nand U2055 (N_2055,In_253,In_1067);
nor U2056 (N_2056,In_348,In_1130);
xnor U2057 (N_2057,In_1478,In_516);
xor U2058 (N_2058,In_1341,In_712);
xor U2059 (N_2059,In_1431,In_1011);
nor U2060 (N_2060,In_1147,In_833);
nor U2061 (N_2061,In_799,In_786);
xor U2062 (N_2062,In_1371,In_1269);
or U2063 (N_2063,In_804,In_1128);
nand U2064 (N_2064,In_674,In_169);
nand U2065 (N_2065,In_1160,In_319);
and U2066 (N_2066,In_853,In_805);
xnor U2067 (N_2067,In_688,In_690);
and U2068 (N_2068,In_1474,In_1294);
nor U2069 (N_2069,In_925,In_854);
nand U2070 (N_2070,In_712,In_1207);
and U2071 (N_2071,In_1123,In_1033);
nor U2072 (N_2072,In_81,In_1491);
nand U2073 (N_2073,In_1161,In_44);
xor U2074 (N_2074,In_949,In_1278);
nand U2075 (N_2075,In_1492,In_653);
nand U2076 (N_2076,In_617,In_190);
or U2077 (N_2077,In_1206,In_676);
and U2078 (N_2078,In_1318,In_859);
nor U2079 (N_2079,In_1028,In_381);
nand U2080 (N_2080,In_209,In_410);
nand U2081 (N_2081,In_145,In_864);
xor U2082 (N_2082,In_134,In_431);
and U2083 (N_2083,In_938,In_494);
xor U2084 (N_2084,In_589,In_79);
and U2085 (N_2085,In_1100,In_424);
xor U2086 (N_2086,In_1375,In_420);
nand U2087 (N_2087,In_291,In_674);
nor U2088 (N_2088,In_219,In_582);
nand U2089 (N_2089,In_506,In_431);
xor U2090 (N_2090,In_455,In_723);
and U2091 (N_2091,In_693,In_1094);
or U2092 (N_2092,In_177,In_202);
or U2093 (N_2093,In_1482,In_1351);
xnor U2094 (N_2094,In_4,In_1277);
xor U2095 (N_2095,In_72,In_1426);
nor U2096 (N_2096,In_56,In_80);
xnor U2097 (N_2097,In_723,In_1251);
or U2098 (N_2098,In_1272,In_479);
nor U2099 (N_2099,In_1086,In_1408);
xor U2100 (N_2100,In_832,In_198);
xor U2101 (N_2101,In_1261,In_260);
nand U2102 (N_2102,In_1152,In_675);
and U2103 (N_2103,In_285,In_1035);
nor U2104 (N_2104,In_919,In_1456);
nand U2105 (N_2105,In_1468,In_617);
or U2106 (N_2106,In_241,In_1302);
and U2107 (N_2107,In_1417,In_662);
or U2108 (N_2108,In_175,In_1089);
xor U2109 (N_2109,In_613,In_1459);
and U2110 (N_2110,In_668,In_998);
xor U2111 (N_2111,In_1085,In_745);
and U2112 (N_2112,In_939,In_963);
nand U2113 (N_2113,In_518,In_1363);
xnor U2114 (N_2114,In_781,In_637);
or U2115 (N_2115,In_136,In_5);
nor U2116 (N_2116,In_1179,In_1263);
nand U2117 (N_2117,In_376,In_1398);
and U2118 (N_2118,In_1334,In_1084);
nand U2119 (N_2119,In_1494,In_1104);
nor U2120 (N_2120,In_944,In_811);
nand U2121 (N_2121,In_1015,In_1293);
xnor U2122 (N_2122,In_1377,In_786);
and U2123 (N_2123,In_395,In_1389);
nand U2124 (N_2124,In_1245,In_328);
nand U2125 (N_2125,In_1372,In_374);
nand U2126 (N_2126,In_612,In_893);
xnor U2127 (N_2127,In_534,In_763);
nand U2128 (N_2128,In_1070,In_691);
and U2129 (N_2129,In_1165,In_239);
and U2130 (N_2130,In_1229,In_550);
or U2131 (N_2131,In_844,In_379);
or U2132 (N_2132,In_202,In_902);
or U2133 (N_2133,In_668,In_999);
xor U2134 (N_2134,In_1494,In_1499);
nand U2135 (N_2135,In_374,In_873);
and U2136 (N_2136,In_127,In_71);
and U2137 (N_2137,In_111,In_678);
or U2138 (N_2138,In_10,In_376);
nand U2139 (N_2139,In_584,In_588);
or U2140 (N_2140,In_166,In_1168);
nand U2141 (N_2141,In_1188,In_67);
or U2142 (N_2142,In_647,In_1211);
xnor U2143 (N_2143,In_1017,In_878);
nand U2144 (N_2144,In_11,In_225);
nand U2145 (N_2145,In_895,In_428);
xnor U2146 (N_2146,In_513,In_1144);
or U2147 (N_2147,In_1267,In_339);
or U2148 (N_2148,In_478,In_3);
nand U2149 (N_2149,In_1448,In_33);
and U2150 (N_2150,In_714,In_932);
and U2151 (N_2151,In_1053,In_468);
nor U2152 (N_2152,In_381,In_1451);
nor U2153 (N_2153,In_27,In_342);
nand U2154 (N_2154,In_525,In_1281);
nand U2155 (N_2155,In_1356,In_624);
nand U2156 (N_2156,In_123,In_975);
xnor U2157 (N_2157,In_738,In_710);
nor U2158 (N_2158,In_247,In_392);
nor U2159 (N_2159,In_656,In_1084);
nor U2160 (N_2160,In_1248,In_422);
and U2161 (N_2161,In_783,In_1366);
nand U2162 (N_2162,In_941,In_609);
nor U2163 (N_2163,In_711,In_41);
nor U2164 (N_2164,In_843,In_1145);
xnor U2165 (N_2165,In_521,In_794);
nor U2166 (N_2166,In_767,In_1028);
nand U2167 (N_2167,In_1168,In_504);
xor U2168 (N_2168,In_174,In_1065);
xor U2169 (N_2169,In_1342,In_66);
xnor U2170 (N_2170,In_204,In_177);
xor U2171 (N_2171,In_222,In_1192);
and U2172 (N_2172,In_1200,In_1186);
or U2173 (N_2173,In_1080,In_506);
and U2174 (N_2174,In_947,In_91);
xnor U2175 (N_2175,In_1339,In_1268);
xnor U2176 (N_2176,In_973,In_607);
and U2177 (N_2177,In_898,In_749);
and U2178 (N_2178,In_792,In_1218);
xor U2179 (N_2179,In_54,In_135);
or U2180 (N_2180,In_315,In_231);
xor U2181 (N_2181,In_285,In_929);
or U2182 (N_2182,In_122,In_971);
xor U2183 (N_2183,In_1130,In_1425);
and U2184 (N_2184,In_202,In_936);
and U2185 (N_2185,In_570,In_60);
nor U2186 (N_2186,In_761,In_21);
and U2187 (N_2187,In_1072,In_453);
nor U2188 (N_2188,In_828,In_1197);
xor U2189 (N_2189,In_16,In_992);
or U2190 (N_2190,In_816,In_1401);
nor U2191 (N_2191,In_1116,In_1123);
nor U2192 (N_2192,In_1206,In_156);
xnor U2193 (N_2193,In_547,In_729);
nor U2194 (N_2194,In_564,In_430);
nor U2195 (N_2195,In_172,In_695);
nand U2196 (N_2196,In_796,In_373);
nor U2197 (N_2197,In_1002,In_232);
nor U2198 (N_2198,In_292,In_343);
and U2199 (N_2199,In_736,In_1430);
or U2200 (N_2200,In_85,In_657);
nor U2201 (N_2201,In_1382,In_1089);
nor U2202 (N_2202,In_112,In_118);
nor U2203 (N_2203,In_480,In_898);
xor U2204 (N_2204,In_1304,In_159);
nor U2205 (N_2205,In_1295,In_1109);
or U2206 (N_2206,In_395,In_177);
nor U2207 (N_2207,In_499,In_1230);
xnor U2208 (N_2208,In_361,In_812);
or U2209 (N_2209,In_1285,In_1349);
or U2210 (N_2210,In_487,In_1215);
nand U2211 (N_2211,In_1102,In_1035);
xor U2212 (N_2212,In_1174,In_17);
xnor U2213 (N_2213,In_1373,In_452);
and U2214 (N_2214,In_114,In_1146);
xnor U2215 (N_2215,In_91,In_1215);
or U2216 (N_2216,In_259,In_1194);
nor U2217 (N_2217,In_1020,In_1191);
and U2218 (N_2218,In_1299,In_742);
and U2219 (N_2219,In_439,In_60);
and U2220 (N_2220,In_464,In_1104);
nor U2221 (N_2221,In_1398,In_1406);
and U2222 (N_2222,In_1115,In_324);
nor U2223 (N_2223,In_351,In_320);
nor U2224 (N_2224,In_934,In_371);
nor U2225 (N_2225,In_1353,In_1096);
nor U2226 (N_2226,In_249,In_862);
or U2227 (N_2227,In_665,In_567);
or U2228 (N_2228,In_932,In_790);
nand U2229 (N_2229,In_262,In_257);
nor U2230 (N_2230,In_1325,In_910);
and U2231 (N_2231,In_142,In_812);
nand U2232 (N_2232,In_471,In_1015);
or U2233 (N_2233,In_1449,In_1046);
xnor U2234 (N_2234,In_1140,In_209);
nor U2235 (N_2235,In_1189,In_269);
or U2236 (N_2236,In_1305,In_1393);
or U2237 (N_2237,In_1244,In_393);
nor U2238 (N_2238,In_1481,In_1171);
or U2239 (N_2239,In_1321,In_764);
or U2240 (N_2240,In_759,In_729);
and U2241 (N_2241,In_1168,In_652);
and U2242 (N_2242,In_858,In_1137);
and U2243 (N_2243,In_1185,In_718);
xnor U2244 (N_2244,In_1098,In_981);
and U2245 (N_2245,In_765,In_1463);
xnor U2246 (N_2246,In_170,In_599);
or U2247 (N_2247,In_513,In_413);
nor U2248 (N_2248,In_313,In_96);
xor U2249 (N_2249,In_29,In_1150);
or U2250 (N_2250,In_1048,In_1260);
nor U2251 (N_2251,In_820,In_1023);
nor U2252 (N_2252,In_785,In_671);
nor U2253 (N_2253,In_21,In_805);
nor U2254 (N_2254,In_1395,In_628);
and U2255 (N_2255,In_291,In_1374);
nor U2256 (N_2256,In_323,In_754);
xnor U2257 (N_2257,In_8,In_201);
or U2258 (N_2258,In_42,In_325);
nand U2259 (N_2259,In_1186,In_1002);
nand U2260 (N_2260,In_529,In_754);
nand U2261 (N_2261,In_798,In_38);
and U2262 (N_2262,In_1181,In_384);
xor U2263 (N_2263,In_244,In_697);
and U2264 (N_2264,In_26,In_1018);
xor U2265 (N_2265,In_1350,In_1370);
nor U2266 (N_2266,In_548,In_73);
nand U2267 (N_2267,In_1398,In_918);
or U2268 (N_2268,In_964,In_689);
nand U2269 (N_2269,In_784,In_1357);
and U2270 (N_2270,In_1083,In_1272);
nor U2271 (N_2271,In_1332,In_381);
and U2272 (N_2272,In_1129,In_1185);
or U2273 (N_2273,In_1092,In_420);
xor U2274 (N_2274,In_741,In_1253);
and U2275 (N_2275,In_725,In_1125);
nand U2276 (N_2276,In_1235,In_1088);
nor U2277 (N_2277,In_232,In_268);
and U2278 (N_2278,In_49,In_1376);
xnor U2279 (N_2279,In_1357,In_1070);
nor U2280 (N_2280,In_1136,In_942);
nor U2281 (N_2281,In_557,In_1349);
xor U2282 (N_2282,In_289,In_441);
nand U2283 (N_2283,In_1430,In_334);
nand U2284 (N_2284,In_317,In_638);
and U2285 (N_2285,In_51,In_1467);
nand U2286 (N_2286,In_374,In_600);
xor U2287 (N_2287,In_1330,In_209);
nand U2288 (N_2288,In_384,In_447);
or U2289 (N_2289,In_1035,In_1241);
and U2290 (N_2290,In_675,In_57);
and U2291 (N_2291,In_228,In_327);
or U2292 (N_2292,In_834,In_724);
nand U2293 (N_2293,In_378,In_931);
nand U2294 (N_2294,In_694,In_491);
or U2295 (N_2295,In_1107,In_821);
or U2296 (N_2296,In_1319,In_484);
xnor U2297 (N_2297,In_872,In_1495);
and U2298 (N_2298,In_690,In_123);
nand U2299 (N_2299,In_566,In_1367);
and U2300 (N_2300,In_716,In_65);
nand U2301 (N_2301,In_868,In_247);
nand U2302 (N_2302,In_166,In_79);
and U2303 (N_2303,In_1374,In_602);
xnor U2304 (N_2304,In_47,In_1360);
and U2305 (N_2305,In_1497,In_1313);
nor U2306 (N_2306,In_271,In_1176);
nor U2307 (N_2307,In_251,In_476);
or U2308 (N_2308,In_1440,In_74);
and U2309 (N_2309,In_769,In_370);
and U2310 (N_2310,In_597,In_1023);
and U2311 (N_2311,In_429,In_718);
or U2312 (N_2312,In_307,In_697);
nand U2313 (N_2313,In_1296,In_107);
xnor U2314 (N_2314,In_1166,In_855);
nor U2315 (N_2315,In_447,In_196);
nand U2316 (N_2316,In_646,In_1378);
nand U2317 (N_2317,In_1113,In_550);
nand U2318 (N_2318,In_907,In_1182);
or U2319 (N_2319,In_476,In_68);
and U2320 (N_2320,In_13,In_330);
xor U2321 (N_2321,In_664,In_520);
and U2322 (N_2322,In_44,In_1340);
or U2323 (N_2323,In_250,In_684);
or U2324 (N_2324,In_1407,In_46);
or U2325 (N_2325,In_366,In_452);
or U2326 (N_2326,In_1062,In_579);
and U2327 (N_2327,In_908,In_1080);
nor U2328 (N_2328,In_1436,In_419);
xor U2329 (N_2329,In_38,In_371);
nor U2330 (N_2330,In_1229,In_813);
nand U2331 (N_2331,In_560,In_161);
nand U2332 (N_2332,In_123,In_1284);
nand U2333 (N_2333,In_316,In_1410);
xnor U2334 (N_2334,In_195,In_830);
or U2335 (N_2335,In_1361,In_207);
nand U2336 (N_2336,In_951,In_779);
or U2337 (N_2337,In_835,In_260);
nor U2338 (N_2338,In_779,In_1217);
or U2339 (N_2339,In_381,In_517);
nand U2340 (N_2340,In_839,In_936);
nor U2341 (N_2341,In_860,In_969);
nand U2342 (N_2342,In_804,In_807);
xor U2343 (N_2343,In_42,In_969);
and U2344 (N_2344,In_63,In_1243);
xnor U2345 (N_2345,In_708,In_268);
nor U2346 (N_2346,In_780,In_1473);
and U2347 (N_2347,In_739,In_545);
and U2348 (N_2348,In_339,In_1246);
nor U2349 (N_2349,In_185,In_957);
and U2350 (N_2350,In_1382,In_987);
nor U2351 (N_2351,In_647,In_390);
nor U2352 (N_2352,In_940,In_1456);
or U2353 (N_2353,In_274,In_1497);
or U2354 (N_2354,In_114,In_974);
and U2355 (N_2355,In_1155,In_474);
or U2356 (N_2356,In_1314,In_721);
nor U2357 (N_2357,In_1463,In_436);
nand U2358 (N_2358,In_1064,In_804);
xnor U2359 (N_2359,In_867,In_636);
xor U2360 (N_2360,In_529,In_1258);
nand U2361 (N_2361,In_985,In_1215);
nand U2362 (N_2362,In_978,In_1407);
and U2363 (N_2363,In_419,In_1075);
or U2364 (N_2364,In_1241,In_1233);
nor U2365 (N_2365,In_1374,In_225);
xnor U2366 (N_2366,In_413,In_58);
nor U2367 (N_2367,In_670,In_23);
nor U2368 (N_2368,In_1419,In_1029);
nand U2369 (N_2369,In_352,In_1416);
nor U2370 (N_2370,In_485,In_874);
or U2371 (N_2371,In_1022,In_1258);
or U2372 (N_2372,In_643,In_1260);
xnor U2373 (N_2373,In_716,In_781);
nor U2374 (N_2374,In_1128,In_1356);
and U2375 (N_2375,In_983,In_699);
xor U2376 (N_2376,In_164,In_583);
nor U2377 (N_2377,In_1177,In_962);
nand U2378 (N_2378,In_7,In_1079);
or U2379 (N_2379,In_409,In_779);
and U2380 (N_2380,In_1152,In_460);
nor U2381 (N_2381,In_337,In_633);
nor U2382 (N_2382,In_1495,In_1176);
or U2383 (N_2383,In_552,In_941);
and U2384 (N_2384,In_1384,In_1433);
or U2385 (N_2385,In_1204,In_1261);
nor U2386 (N_2386,In_1211,In_506);
nand U2387 (N_2387,In_340,In_1497);
xnor U2388 (N_2388,In_150,In_615);
nor U2389 (N_2389,In_946,In_903);
and U2390 (N_2390,In_1427,In_947);
nor U2391 (N_2391,In_279,In_737);
nor U2392 (N_2392,In_1101,In_83);
xor U2393 (N_2393,In_1036,In_201);
or U2394 (N_2394,In_635,In_461);
nor U2395 (N_2395,In_949,In_186);
nand U2396 (N_2396,In_1411,In_549);
and U2397 (N_2397,In_450,In_1141);
and U2398 (N_2398,In_618,In_1346);
nand U2399 (N_2399,In_634,In_714);
or U2400 (N_2400,In_1334,In_1305);
xnor U2401 (N_2401,In_519,In_952);
or U2402 (N_2402,In_303,In_550);
nor U2403 (N_2403,In_192,In_314);
or U2404 (N_2404,In_936,In_588);
xnor U2405 (N_2405,In_1417,In_873);
or U2406 (N_2406,In_953,In_322);
nor U2407 (N_2407,In_703,In_240);
xnor U2408 (N_2408,In_1053,In_969);
and U2409 (N_2409,In_946,In_395);
or U2410 (N_2410,In_808,In_1028);
or U2411 (N_2411,In_1442,In_594);
nand U2412 (N_2412,In_342,In_1057);
nand U2413 (N_2413,In_462,In_160);
xnor U2414 (N_2414,In_468,In_879);
nor U2415 (N_2415,In_376,In_975);
or U2416 (N_2416,In_665,In_356);
nand U2417 (N_2417,In_223,In_256);
and U2418 (N_2418,In_222,In_1200);
or U2419 (N_2419,In_937,In_982);
xnor U2420 (N_2420,In_1276,In_40);
or U2421 (N_2421,In_303,In_697);
nor U2422 (N_2422,In_33,In_544);
nand U2423 (N_2423,In_344,In_53);
nor U2424 (N_2424,In_219,In_665);
xnor U2425 (N_2425,In_1036,In_191);
xor U2426 (N_2426,In_474,In_726);
and U2427 (N_2427,In_860,In_1043);
and U2428 (N_2428,In_90,In_94);
nand U2429 (N_2429,In_566,In_809);
nand U2430 (N_2430,In_600,In_973);
nor U2431 (N_2431,In_360,In_459);
or U2432 (N_2432,In_937,In_597);
nor U2433 (N_2433,In_1473,In_1393);
or U2434 (N_2434,In_654,In_922);
or U2435 (N_2435,In_247,In_419);
and U2436 (N_2436,In_1309,In_1034);
and U2437 (N_2437,In_521,In_356);
nor U2438 (N_2438,In_117,In_991);
or U2439 (N_2439,In_118,In_630);
xor U2440 (N_2440,In_1337,In_748);
nand U2441 (N_2441,In_1096,In_242);
nor U2442 (N_2442,In_72,In_372);
xnor U2443 (N_2443,In_435,In_1118);
or U2444 (N_2444,In_614,In_741);
and U2445 (N_2445,In_1227,In_1281);
nor U2446 (N_2446,In_1425,In_1095);
xnor U2447 (N_2447,In_1200,In_453);
xnor U2448 (N_2448,In_202,In_791);
and U2449 (N_2449,In_1095,In_1314);
or U2450 (N_2450,In_1228,In_1005);
nor U2451 (N_2451,In_774,In_909);
nor U2452 (N_2452,In_616,In_1431);
or U2453 (N_2453,In_301,In_252);
and U2454 (N_2454,In_1238,In_1462);
nor U2455 (N_2455,In_963,In_1007);
nor U2456 (N_2456,In_88,In_1226);
and U2457 (N_2457,In_535,In_770);
nor U2458 (N_2458,In_930,In_883);
nand U2459 (N_2459,In_699,In_450);
xor U2460 (N_2460,In_72,In_381);
nand U2461 (N_2461,In_1431,In_1206);
nor U2462 (N_2462,In_636,In_144);
or U2463 (N_2463,In_769,In_537);
nand U2464 (N_2464,In_1369,In_259);
nand U2465 (N_2465,In_760,In_0);
xnor U2466 (N_2466,In_302,In_1383);
xnor U2467 (N_2467,In_1253,In_455);
xnor U2468 (N_2468,In_312,In_908);
nor U2469 (N_2469,In_382,In_928);
xnor U2470 (N_2470,In_976,In_876);
nand U2471 (N_2471,In_1254,In_1003);
nor U2472 (N_2472,In_1392,In_102);
nor U2473 (N_2473,In_1384,In_602);
nand U2474 (N_2474,In_984,In_998);
and U2475 (N_2475,In_1315,In_1459);
xor U2476 (N_2476,In_151,In_640);
or U2477 (N_2477,In_407,In_95);
nor U2478 (N_2478,In_1081,In_1117);
and U2479 (N_2479,In_1343,In_559);
xnor U2480 (N_2480,In_326,In_344);
nand U2481 (N_2481,In_187,In_1021);
and U2482 (N_2482,In_951,In_423);
or U2483 (N_2483,In_1072,In_270);
or U2484 (N_2484,In_980,In_1124);
nor U2485 (N_2485,In_1048,In_131);
nand U2486 (N_2486,In_302,In_1443);
and U2487 (N_2487,In_1497,In_939);
and U2488 (N_2488,In_866,In_1469);
and U2489 (N_2489,In_701,In_2);
nor U2490 (N_2490,In_1238,In_1116);
or U2491 (N_2491,In_57,In_220);
and U2492 (N_2492,In_376,In_803);
and U2493 (N_2493,In_1142,In_448);
xor U2494 (N_2494,In_1298,In_207);
xnor U2495 (N_2495,In_669,In_772);
xor U2496 (N_2496,In_322,In_381);
or U2497 (N_2497,In_606,In_286);
and U2498 (N_2498,In_789,In_1372);
or U2499 (N_2499,In_1208,In_157);
xor U2500 (N_2500,In_1401,In_560);
xor U2501 (N_2501,In_687,In_861);
nand U2502 (N_2502,In_1217,In_1214);
nor U2503 (N_2503,In_386,In_1453);
and U2504 (N_2504,In_47,In_635);
nand U2505 (N_2505,In_1175,In_189);
xor U2506 (N_2506,In_735,In_164);
and U2507 (N_2507,In_1144,In_1252);
and U2508 (N_2508,In_708,In_1331);
and U2509 (N_2509,In_487,In_524);
nand U2510 (N_2510,In_1488,In_222);
or U2511 (N_2511,In_1143,In_835);
xor U2512 (N_2512,In_671,In_279);
xor U2513 (N_2513,In_765,In_1083);
or U2514 (N_2514,In_569,In_257);
nand U2515 (N_2515,In_130,In_1488);
nand U2516 (N_2516,In_1320,In_1139);
or U2517 (N_2517,In_1026,In_68);
or U2518 (N_2518,In_1222,In_1259);
and U2519 (N_2519,In_88,In_753);
xor U2520 (N_2520,In_646,In_257);
nand U2521 (N_2521,In_312,In_402);
and U2522 (N_2522,In_1278,In_209);
or U2523 (N_2523,In_145,In_45);
or U2524 (N_2524,In_460,In_38);
nand U2525 (N_2525,In_418,In_501);
nand U2526 (N_2526,In_96,In_1013);
xnor U2527 (N_2527,In_872,In_913);
or U2528 (N_2528,In_192,In_1051);
xor U2529 (N_2529,In_1419,In_690);
nor U2530 (N_2530,In_196,In_798);
and U2531 (N_2531,In_622,In_163);
nor U2532 (N_2532,In_1299,In_1366);
nor U2533 (N_2533,In_1392,In_1400);
and U2534 (N_2534,In_198,In_365);
nor U2535 (N_2535,In_570,In_809);
xnor U2536 (N_2536,In_235,In_160);
nand U2537 (N_2537,In_475,In_1049);
and U2538 (N_2538,In_310,In_1063);
and U2539 (N_2539,In_1294,In_317);
xnor U2540 (N_2540,In_857,In_334);
nand U2541 (N_2541,In_841,In_1486);
and U2542 (N_2542,In_444,In_272);
nand U2543 (N_2543,In_128,In_403);
and U2544 (N_2544,In_773,In_182);
xnor U2545 (N_2545,In_1432,In_123);
xor U2546 (N_2546,In_332,In_1125);
nor U2547 (N_2547,In_337,In_498);
or U2548 (N_2548,In_954,In_427);
xor U2549 (N_2549,In_532,In_690);
xnor U2550 (N_2550,In_797,In_1141);
nand U2551 (N_2551,In_179,In_637);
nand U2552 (N_2552,In_271,In_684);
xnor U2553 (N_2553,In_58,In_401);
nor U2554 (N_2554,In_902,In_951);
nor U2555 (N_2555,In_725,In_1353);
or U2556 (N_2556,In_291,In_794);
or U2557 (N_2557,In_491,In_1171);
and U2558 (N_2558,In_1005,In_206);
or U2559 (N_2559,In_682,In_961);
xnor U2560 (N_2560,In_866,In_1310);
and U2561 (N_2561,In_1091,In_1252);
nor U2562 (N_2562,In_1173,In_1400);
xnor U2563 (N_2563,In_1495,In_187);
nor U2564 (N_2564,In_177,In_912);
or U2565 (N_2565,In_98,In_247);
xor U2566 (N_2566,In_97,In_133);
or U2567 (N_2567,In_946,In_1149);
xor U2568 (N_2568,In_1451,In_946);
nor U2569 (N_2569,In_4,In_792);
xor U2570 (N_2570,In_790,In_163);
xor U2571 (N_2571,In_609,In_370);
and U2572 (N_2572,In_959,In_291);
xnor U2573 (N_2573,In_783,In_1409);
nand U2574 (N_2574,In_191,In_1440);
and U2575 (N_2575,In_99,In_1274);
nor U2576 (N_2576,In_422,In_1309);
and U2577 (N_2577,In_861,In_336);
nor U2578 (N_2578,In_307,In_740);
nand U2579 (N_2579,In_729,In_423);
and U2580 (N_2580,In_744,In_1406);
xnor U2581 (N_2581,In_823,In_47);
or U2582 (N_2582,In_550,In_933);
and U2583 (N_2583,In_471,In_983);
or U2584 (N_2584,In_1009,In_301);
nor U2585 (N_2585,In_475,In_901);
nand U2586 (N_2586,In_437,In_272);
and U2587 (N_2587,In_810,In_466);
or U2588 (N_2588,In_666,In_1494);
or U2589 (N_2589,In_421,In_1316);
and U2590 (N_2590,In_1399,In_891);
nand U2591 (N_2591,In_887,In_1318);
or U2592 (N_2592,In_1187,In_588);
nand U2593 (N_2593,In_737,In_699);
and U2594 (N_2594,In_444,In_101);
and U2595 (N_2595,In_1166,In_1346);
nor U2596 (N_2596,In_877,In_146);
or U2597 (N_2597,In_1379,In_1055);
or U2598 (N_2598,In_1450,In_491);
and U2599 (N_2599,In_750,In_210);
and U2600 (N_2600,In_809,In_1091);
and U2601 (N_2601,In_1124,In_284);
nor U2602 (N_2602,In_502,In_75);
nor U2603 (N_2603,In_1079,In_451);
or U2604 (N_2604,In_1208,In_773);
nor U2605 (N_2605,In_614,In_58);
or U2606 (N_2606,In_1214,In_1254);
nand U2607 (N_2607,In_1262,In_506);
or U2608 (N_2608,In_1374,In_900);
xor U2609 (N_2609,In_11,In_265);
or U2610 (N_2610,In_80,In_182);
nor U2611 (N_2611,In_179,In_22);
nand U2612 (N_2612,In_1050,In_792);
nand U2613 (N_2613,In_523,In_622);
nor U2614 (N_2614,In_232,In_488);
nor U2615 (N_2615,In_1437,In_1318);
and U2616 (N_2616,In_11,In_203);
nand U2617 (N_2617,In_638,In_773);
and U2618 (N_2618,In_879,In_81);
nand U2619 (N_2619,In_1269,In_129);
nor U2620 (N_2620,In_1418,In_24);
and U2621 (N_2621,In_1040,In_796);
or U2622 (N_2622,In_1066,In_984);
nand U2623 (N_2623,In_18,In_1372);
nor U2624 (N_2624,In_393,In_1458);
nor U2625 (N_2625,In_1075,In_807);
nand U2626 (N_2626,In_1009,In_696);
nand U2627 (N_2627,In_1073,In_981);
xnor U2628 (N_2628,In_773,In_1115);
and U2629 (N_2629,In_1314,In_676);
nand U2630 (N_2630,In_133,In_1466);
xor U2631 (N_2631,In_841,In_1014);
nand U2632 (N_2632,In_1079,In_137);
nand U2633 (N_2633,In_627,In_1246);
nor U2634 (N_2634,In_1285,In_290);
xor U2635 (N_2635,In_322,In_1316);
nor U2636 (N_2636,In_147,In_1072);
xor U2637 (N_2637,In_414,In_779);
xnor U2638 (N_2638,In_981,In_417);
nor U2639 (N_2639,In_288,In_483);
nor U2640 (N_2640,In_871,In_451);
xnor U2641 (N_2641,In_243,In_1275);
and U2642 (N_2642,In_1030,In_825);
and U2643 (N_2643,In_1008,In_297);
nor U2644 (N_2644,In_312,In_97);
xnor U2645 (N_2645,In_1341,In_611);
and U2646 (N_2646,In_1368,In_1157);
nand U2647 (N_2647,In_1170,In_154);
nand U2648 (N_2648,In_939,In_19);
or U2649 (N_2649,In_429,In_621);
nor U2650 (N_2650,In_756,In_23);
nand U2651 (N_2651,In_918,In_1463);
and U2652 (N_2652,In_729,In_332);
xnor U2653 (N_2653,In_663,In_114);
or U2654 (N_2654,In_1167,In_363);
nand U2655 (N_2655,In_136,In_1016);
nand U2656 (N_2656,In_649,In_341);
xor U2657 (N_2657,In_1345,In_109);
nand U2658 (N_2658,In_88,In_1258);
or U2659 (N_2659,In_661,In_922);
nor U2660 (N_2660,In_190,In_1235);
and U2661 (N_2661,In_1221,In_1348);
and U2662 (N_2662,In_1383,In_454);
nand U2663 (N_2663,In_1231,In_664);
xor U2664 (N_2664,In_905,In_1293);
or U2665 (N_2665,In_1331,In_1017);
nand U2666 (N_2666,In_1488,In_67);
or U2667 (N_2667,In_238,In_750);
or U2668 (N_2668,In_1349,In_733);
xor U2669 (N_2669,In_899,In_1026);
or U2670 (N_2670,In_1324,In_1301);
nand U2671 (N_2671,In_1193,In_727);
nor U2672 (N_2672,In_355,In_1179);
nor U2673 (N_2673,In_706,In_369);
or U2674 (N_2674,In_999,In_331);
or U2675 (N_2675,In_1412,In_598);
or U2676 (N_2676,In_1070,In_1207);
xnor U2677 (N_2677,In_456,In_149);
and U2678 (N_2678,In_1181,In_833);
or U2679 (N_2679,In_955,In_796);
or U2680 (N_2680,In_573,In_722);
nand U2681 (N_2681,In_1464,In_1156);
nor U2682 (N_2682,In_1088,In_39);
or U2683 (N_2683,In_494,In_342);
or U2684 (N_2684,In_592,In_310);
nor U2685 (N_2685,In_1016,In_520);
nor U2686 (N_2686,In_196,In_205);
and U2687 (N_2687,In_874,In_928);
or U2688 (N_2688,In_310,In_420);
or U2689 (N_2689,In_897,In_807);
nand U2690 (N_2690,In_1062,In_7);
or U2691 (N_2691,In_836,In_1461);
and U2692 (N_2692,In_535,In_1024);
and U2693 (N_2693,In_1147,In_919);
and U2694 (N_2694,In_888,In_1227);
and U2695 (N_2695,In_1313,In_344);
and U2696 (N_2696,In_1297,In_1248);
xnor U2697 (N_2697,In_1079,In_574);
and U2698 (N_2698,In_64,In_1267);
or U2699 (N_2699,In_937,In_216);
or U2700 (N_2700,In_589,In_1057);
or U2701 (N_2701,In_1206,In_265);
nor U2702 (N_2702,In_1213,In_1031);
or U2703 (N_2703,In_53,In_528);
nand U2704 (N_2704,In_536,In_150);
or U2705 (N_2705,In_274,In_235);
nor U2706 (N_2706,In_438,In_1072);
nand U2707 (N_2707,In_874,In_358);
nand U2708 (N_2708,In_1323,In_682);
nor U2709 (N_2709,In_776,In_411);
and U2710 (N_2710,In_879,In_25);
nand U2711 (N_2711,In_55,In_226);
nand U2712 (N_2712,In_978,In_280);
xor U2713 (N_2713,In_80,In_598);
xnor U2714 (N_2714,In_722,In_827);
nand U2715 (N_2715,In_375,In_898);
or U2716 (N_2716,In_1322,In_516);
and U2717 (N_2717,In_836,In_347);
nor U2718 (N_2718,In_1220,In_1081);
nand U2719 (N_2719,In_150,In_1491);
and U2720 (N_2720,In_21,In_530);
and U2721 (N_2721,In_319,In_627);
nand U2722 (N_2722,In_1384,In_640);
and U2723 (N_2723,In_1498,In_1012);
xnor U2724 (N_2724,In_676,In_103);
and U2725 (N_2725,In_606,In_1454);
or U2726 (N_2726,In_1373,In_1197);
xnor U2727 (N_2727,In_889,In_1013);
xnor U2728 (N_2728,In_212,In_567);
or U2729 (N_2729,In_817,In_743);
nand U2730 (N_2730,In_1268,In_366);
or U2731 (N_2731,In_1368,In_423);
nand U2732 (N_2732,In_731,In_1378);
or U2733 (N_2733,In_1286,In_914);
nor U2734 (N_2734,In_68,In_1353);
and U2735 (N_2735,In_1093,In_525);
nor U2736 (N_2736,In_1286,In_1273);
xnor U2737 (N_2737,In_1244,In_577);
and U2738 (N_2738,In_781,In_226);
xnor U2739 (N_2739,In_84,In_874);
nor U2740 (N_2740,In_38,In_241);
or U2741 (N_2741,In_345,In_111);
and U2742 (N_2742,In_755,In_473);
and U2743 (N_2743,In_1373,In_78);
or U2744 (N_2744,In_1437,In_1122);
and U2745 (N_2745,In_797,In_1222);
or U2746 (N_2746,In_209,In_571);
xor U2747 (N_2747,In_1207,In_109);
nor U2748 (N_2748,In_1100,In_353);
nand U2749 (N_2749,In_279,In_432);
nor U2750 (N_2750,In_829,In_1186);
or U2751 (N_2751,In_1378,In_1420);
and U2752 (N_2752,In_505,In_1379);
and U2753 (N_2753,In_969,In_1088);
and U2754 (N_2754,In_1321,In_1228);
and U2755 (N_2755,In_1327,In_589);
xnor U2756 (N_2756,In_149,In_66);
nor U2757 (N_2757,In_520,In_274);
nor U2758 (N_2758,In_1112,In_888);
nor U2759 (N_2759,In_657,In_405);
xor U2760 (N_2760,In_1367,In_818);
and U2761 (N_2761,In_1225,In_240);
nand U2762 (N_2762,In_883,In_105);
and U2763 (N_2763,In_97,In_495);
or U2764 (N_2764,In_652,In_1084);
or U2765 (N_2765,In_387,In_893);
and U2766 (N_2766,In_664,In_1022);
nand U2767 (N_2767,In_239,In_611);
xor U2768 (N_2768,In_326,In_1265);
or U2769 (N_2769,In_744,In_1120);
xnor U2770 (N_2770,In_912,In_819);
nor U2771 (N_2771,In_910,In_235);
or U2772 (N_2772,In_159,In_1208);
and U2773 (N_2773,In_531,In_819);
xnor U2774 (N_2774,In_386,In_749);
xnor U2775 (N_2775,In_1021,In_699);
and U2776 (N_2776,In_1295,In_212);
nor U2777 (N_2777,In_527,In_798);
nand U2778 (N_2778,In_62,In_844);
nor U2779 (N_2779,In_1374,In_1383);
nand U2780 (N_2780,In_1335,In_761);
or U2781 (N_2781,In_590,In_777);
xnor U2782 (N_2782,In_1015,In_1294);
nor U2783 (N_2783,In_1076,In_1038);
xnor U2784 (N_2784,In_13,In_888);
and U2785 (N_2785,In_1396,In_1042);
xnor U2786 (N_2786,In_226,In_1132);
or U2787 (N_2787,In_1306,In_1024);
and U2788 (N_2788,In_1424,In_235);
nor U2789 (N_2789,In_1495,In_748);
and U2790 (N_2790,In_1340,In_493);
or U2791 (N_2791,In_1249,In_1462);
nor U2792 (N_2792,In_269,In_405);
nor U2793 (N_2793,In_110,In_238);
xor U2794 (N_2794,In_251,In_780);
or U2795 (N_2795,In_568,In_1083);
and U2796 (N_2796,In_1033,In_363);
nor U2797 (N_2797,In_466,In_811);
or U2798 (N_2798,In_1375,In_377);
or U2799 (N_2799,In_769,In_972);
and U2800 (N_2800,In_491,In_910);
nand U2801 (N_2801,In_102,In_405);
nor U2802 (N_2802,In_1463,In_410);
xnor U2803 (N_2803,In_1437,In_954);
nor U2804 (N_2804,In_438,In_1468);
xnor U2805 (N_2805,In_1095,In_612);
xnor U2806 (N_2806,In_1463,In_1162);
and U2807 (N_2807,In_1450,In_351);
xnor U2808 (N_2808,In_744,In_1152);
nor U2809 (N_2809,In_524,In_349);
xor U2810 (N_2810,In_1263,In_1303);
or U2811 (N_2811,In_203,In_595);
and U2812 (N_2812,In_549,In_499);
xor U2813 (N_2813,In_483,In_140);
or U2814 (N_2814,In_203,In_1376);
nor U2815 (N_2815,In_615,In_684);
and U2816 (N_2816,In_479,In_292);
nor U2817 (N_2817,In_1335,In_1180);
or U2818 (N_2818,In_339,In_1492);
xnor U2819 (N_2819,In_51,In_1074);
nand U2820 (N_2820,In_1080,In_943);
or U2821 (N_2821,In_1490,In_1322);
xor U2822 (N_2822,In_840,In_1256);
xnor U2823 (N_2823,In_1387,In_1032);
nor U2824 (N_2824,In_166,In_89);
or U2825 (N_2825,In_25,In_717);
and U2826 (N_2826,In_1195,In_738);
nand U2827 (N_2827,In_727,In_849);
nor U2828 (N_2828,In_1244,In_837);
or U2829 (N_2829,In_295,In_868);
nor U2830 (N_2830,In_1476,In_770);
nor U2831 (N_2831,In_1105,In_573);
and U2832 (N_2832,In_951,In_1445);
nor U2833 (N_2833,In_496,In_42);
nor U2834 (N_2834,In_672,In_582);
and U2835 (N_2835,In_1286,In_1472);
xor U2836 (N_2836,In_216,In_1172);
and U2837 (N_2837,In_609,In_831);
nand U2838 (N_2838,In_647,In_1260);
xor U2839 (N_2839,In_1077,In_993);
or U2840 (N_2840,In_15,In_1006);
nor U2841 (N_2841,In_1368,In_294);
or U2842 (N_2842,In_736,In_886);
xnor U2843 (N_2843,In_492,In_1129);
or U2844 (N_2844,In_464,In_901);
nand U2845 (N_2845,In_65,In_1185);
xnor U2846 (N_2846,In_385,In_1150);
or U2847 (N_2847,In_1141,In_1019);
nor U2848 (N_2848,In_909,In_1436);
nand U2849 (N_2849,In_1369,In_1446);
xnor U2850 (N_2850,In_1353,In_1044);
nor U2851 (N_2851,In_641,In_1276);
nor U2852 (N_2852,In_430,In_653);
nand U2853 (N_2853,In_1099,In_810);
or U2854 (N_2854,In_17,In_578);
xor U2855 (N_2855,In_62,In_1183);
and U2856 (N_2856,In_757,In_368);
and U2857 (N_2857,In_1458,In_1250);
xor U2858 (N_2858,In_234,In_921);
nand U2859 (N_2859,In_909,In_732);
nor U2860 (N_2860,In_1494,In_1173);
or U2861 (N_2861,In_194,In_388);
nor U2862 (N_2862,In_762,In_427);
nand U2863 (N_2863,In_1342,In_236);
or U2864 (N_2864,In_695,In_155);
nor U2865 (N_2865,In_354,In_432);
or U2866 (N_2866,In_594,In_345);
xor U2867 (N_2867,In_208,In_869);
xnor U2868 (N_2868,In_415,In_951);
and U2869 (N_2869,In_482,In_317);
and U2870 (N_2870,In_1387,In_1393);
and U2871 (N_2871,In_446,In_136);
xnor U2872 (N_2872,In_338,In_27);
or U2873 (N_2873,In_819,In_1249);
nand U2874 (N_2874,In_272,In_1469);
nand U2875 (N_2875,In_489,In_1478);
nand U2876 (N_2876,In_778,In_701);
nand U2877 (N_2877,In_850,In_1066);
nor U2878 (N_2878,In_870,In_643);
or U2879 (N_2879,In_656,In_18);
nor U2880 (N_2880,In_202,In_1129);
or U2881 (N_2881,In_266,In_426);
nor U2882 (N_2882,In_577,In_1284);
and U2883 (N_2883,In_1237,In_1055);
nor U2884 (N_2884,In_1435,In_1448);
and U2885 (N_2885,In_513,In_1363);
nor U2886 (N_2886,In_38,In_223);
nor U2887 (N_2887,In_1256,In_766);
nand U2888 (N_2888,In_454,In_1209);
or U2889 (N_2889,In_1319,In_383);
and U2890 (N_2890,In_158,In_1099);
xor U2891 (N_2891,In_1464,In_1437);
nor U2892 (N_2892,In_745,In_1301);
and U2893 (N_2893,In_724,In_735);
or U2894 (N_2894,In_772,In_1374);
or U2895 (N_2895,In_241,In_1203);
nor U2896 (N_2896,In_906,In_605);
and U2897 (N_2897,In_871,In_324);
nor U2898 (N_2898,In_1175,In_1001);
or U2899 (N_2899,In_259,In_1018);
and U2900 (N_2900,In_1478,In_821);
or U2901 (N_2901,In_476,In_137);
xor U2902 (N_2902,In_797,In_861);
nor U2903 (N_2903,In_106,In_1069);
nand U2904 (N_2904,In_868,In_667);
nor U2905 (N_2905,In_1397,In_775);
nor U2906 (N_2906,In_930,In_1248);
and U2907 (N_2907,In_1083,In_849);
nor U2908 (N_2908,In_122,In_388);
xor U2909 (N_2909,In_72,In_688);
nand U2910 (N_2910,In_110,In_1462);
nor U2911 (N_2911,In_1357,In_930);
nand U2912 (N_2912,In_452,In_1285);
and U2913 (N_2913,In_31,In_1125);
xnor U2914 (N_2914,In_529,In_790);
nor U2915 (N_2915,In_941,In_1362);
and U2916 (N_2916,In_915,In_363);
xnor U2917 (N_2917,In_49,In_257);
nand U2918 (N_2918,In_341,In_774);
and U2919 (N_2919,In_1113,In_90);
nor U2920 (N_2920,In_325,In_950);
or U2921 (N_2921,In_167,In_793);
and U2922 (N_2922,In_42,In_500);
and U2923 (N_2923,In_131,In_605);
and U2924 (N_2924,In_827,In_88);
nand U2925 (N_2925,In_608,In_361);
or U2926 (N_2926,In_279,In_1474);
nand U2927 (N_2927,In_1133,In_902);
and U2928 (N_2928,In_1379,In_67);
nand U2929 (N_2929,In_1285,In_1269);
nand U2930 (N_2930,In_1278,In_1463);
xor U2931 (N_2931,In_934,In_843);
nor U2932 (N_2932,In_1165,In_466);
and U2933 (N_2933,In_558,In_568);
xnor U2934 (N_2934,In_213,In_404);
and U2935 (N_2935,In_1061,In_401);
or U2936 (N_2936,In_1052,In_262);
nor U2937 (N_2937,In_882,In_1359);
nor U2938 (N_2938,In_260,In_504);
xnor U2939 (N_2939,In_433,In_1144);
and U2940 (N_2940,In_1144,In_765);
xor U2941 (N_2941,In_1024,In_120);
and U2942 (N_2942,In_637,In_1283);
or U2943 (N_2943,In_447,In_969);
xnor U2944 (N_2944,In_1389,In_958);
xnor U2945 (N_2945,In_482,In_683);
nor U2946 (N_2946,In_235,In_1270);
nor U2947 (N_2947,In_696,In_319);
xor U2948 (N_2948,In_1191,In_132);
nor U2949 (N_2949,In_1078,In_1108);
nor U2950 (N_2950,In_1220,In_343);
and U2951 (N_2951,In_1477,In_8);
nand U2952 (N_2952,In_658,In_452);
nor U2953 (N_2953,In_884,In_949);
nor U2954 (N_2954,In_706,In_522);
and U2955 (N_2955,In_347,In_353);
nor U2956 (N_2956,In_222,In_697);
and U2957 (N_2957,In_189,In_584);
or U2958 (N_2958,In_1319,In_26);
xnor U2959 (N_2959,In_942,In_1146);
nor U2960 (N_2960,In_359,In_959);
xnor U2961 (N_2961,In_1424,In_303);
nand U2962 (N_2962,In_1397,In_1017);
or U2963 (N_2963,In_1326,In_857);
xor U2964 (N_2964,In_450,In_1077);
or U2965 (N_2965,In_280,In_561);
nor U2966 (N_2966,In_1487,In_176);
nor U2967 (N_2967,In_239,In_977);
nand U2968 (N_2968,In_555,In_835);
xnor U2969 (N_2969,In_134,In_322);
nor U2970 (N_2970,In_400,In_412);
and U2971 (N_2971,In_243,In_1024);
nor U2972 (N_2972,In_664,In_1330);
nor U2973 (N_2973,In_635,In_1288);
xnor U2974 (N_2974,In_1112,In_694);
and U2975 (N_2975,In_1317,In_1132);
nor U2976 (N_2976,In_260,In_363);
or U2977 (N_2977,In_1099,In_404);
nor U2978 (N_2978,In_671,In_1419);
and U2979 (N_2979,In_1233,In_1257);
nor U2980 (N_2980,In_1238,In_475);
or U2981 (N_2981,In_1328,In_314);
nor U2982 (N_2982,In_894,In_301);
xor U2983 (N_2983,In_31,In_674);
nor U2984 (N_2984,In_100,In_65);
xnor U2985 (N_2985,In_1198,In_239);
xnor U2986 (N_2986,In_1065,In_934);
xnor U2987 (N_2987,In_1483,In_999);
nand U2988 (N_2988,In_1427,In_1246);
nor U2989 (N_2989,In_24,In_491);
xor U2990 (N_2990,In_586,In_392);
and U2991 (N_2991,In_1356,In_728);
nor U2992 (N_2992,In_479,In_879);
xor U2993 (N_2993,In_349,In_785);
and U2994 (N_2994,In_1202,In_202);
or U2995 (N_2995,In_874,In_1210);
nor U2996 (N_2996,In_111,In_161);
nor U2997 (N_2997,In_1112,In_1004);
nand U2998 (N_2998,In_1037,In_1150);
or U2999 (N_2999,In_356,In_1352);
or U3000 (N_3000,N_128,N_1315);
and U3001 (N_3001,N_1333,N_922);
nand U3002 (N_3002,N_1915,N_1189);
xor U3003 (N_3003,N_873,N_1789);
or U3004 (N_3004,N_2417,N_720);
xnor U3005 (N_3005,N_2405,N_1110);
nor U3006 (N_3006,N_1016,N_1716);
nor U3007 (N_3007,N_2532,N_1105);
xnor U3008 (N_3008,N_1696,N_2355);
or U3009 (N_3009,N_2108,N_1039);
and U3010 (N_3010,N_1758,N_973);
nand U3011 (N_3011,N_266,N_1944);
xor U3012 (N_3012,N_2648,N_318);
and U3013 (N_3013,N_71,N_1720);
or U3014 (N_3014,N_910,N_244);
nor U3015 (N_3015,N_26,N_1544);
or U3016 (N_3016,N_2041,N_150);
nor U3017 (N_3017,N_1458,N_1381);
xnor U3018 (N_3018,N_159,N_1678);
and U3019 (N_3019,N_1810,N_1380);
nand U3020 (N_3020,N_1558,N_1672);
nand U3021 (N_3021,N_2794,N_970);
xor U3022 (N_3022,N_1060,N_1265);
nor U3023 (N_3023,N_2718,N_224);
nor U3024 (N_3024,N_2698,N_1067);
or U3025 (N_3025,N_2513,N_2706);
nand U3026 (N_3026,N_2072,N_1274);
and U3027 (N_3027,N_327,N_32);
xnor U3028 (N_3028,N_308,N_929);
nor U3029 (N_3029,N_393,N_2805);
nor U3030 (N_3030,N_1909,N_1298);
nand U3031 (N_3031,N_2151,N_2393);
and U3032 (N_3032,N_1943,N_131);
or U3033 (N_3033,N_424,N_918);
and U3034 (N_3034,N_1163,N_1095);
xnor U3035 (N_3035,N_867,N_1719);
nor U3036 (N_3036,N_1974,N_383);
nand U3037 (N_3037,N_2276,N_2837);
and U3038 (N_3038,N_1331,N_2613);
xor U3039 (N_3039,N_2292,N_1545);
and U3040 (N_3040,N_1913,N_117);
or U3041 (N_3041,N_544,N_950);
nor U3042 (N_3042,N_240,N_2947);
and U3043 (N_3043,N_746,N_1538);
nand U3044 (N_3044,N_722,N_2595);
or U3045 (N_3045,N_989,N_1275);
nor U3046 (N_3046,N_493,N_2332);
xor U3047 (N_3047,N_1247,N_2621);
or U3048 (N_3048,N_2295,N_2287);
nor U3049 (N_3049,N_1557,N_302);
xnor U3050 (N_3050,N_761,N_1121);
nand U3051 (N_3051,N_162,N_2551);
and U3052 (N_3052,N_242,N_1806);
and U3053 (N_3053,N_445,N_1084);
xnor U3054 (N_3054,N_875,N_2094);
nand U3055 (N_3055,N_2208,N_2566);
and U3056 (N_3056,N_721,N_1257);
xnor U3057 (N_3057,N_2797,N_123);
xor U3058 (N_3058,N_2778,N_2337);
or U3059 (N_3059,N_285,N_2165);
xor U3060 (N_3060,N_952,N_1066);
xnor U3061 (N_3061,N_887,N_284);
or U3062 (N_3062,N_289,N_2197);
xnor U3063 (N_3063,N_1900,N_41);
and U3064 (N_3064,N_1308,N_2491);
xnor U3065 (N_3065,N_2083,N_1463);
nor U3066 (N_3066,N_1615,N_349);
nor U3067 (N_3067,N_2304,N_1649);
and U3068 (N_3068,N_1712,N_2875);
nor U3069 (N_3069,N_1881,N_264);
xor U3070 (N_3070,N_1813,N_816);
nand U3071 (N_3071,N_1845,N_1908);
nor U3072 (N_3072,N_1144,N_675);
nor U3073 (N_3073,N_651,N_202);
nor U3074 (N_3074,N_699,N_1426);
xnor U3075 (N_3075,N_1435,N_1527);
and U3076 (N_3076,N_2670,N_2173);
nor U3077 (N_3077,N_2011,N_109);
and U3078 (N_3078,N_1848,N_1807);
or U3079 (N_3079,N_1537,N_93);
nand U3080 (N_3080,N_2413,N_314);
and U3081 (N_3081,N_418,N_1541);
nor U3082 (N_3082,N_847,N_1530);
and U3083 (N_3083,N_824,N_569);
nand U3084 (N_3084,N_252,N_1281);
or U3085 (N_3085,N_1759,N_2506);
nand U3086 (N_3086,N_902,N_1085);
nand U3087 (N_3087,N_668,N_1928);
or U3088 (N_3088,N_411,N_1686);
nand U3089 (N_3089,N_1226,N_2635);
nor U3090 (N_3090,N_294,N_864);
xnor U3091 (N_3091,N_2833,N_2178);
xnor U3092 (N_3092,N_707,N_1674);
nor U3093 (N_3093,N_428,N_628);
nor U3094 (N_3094,N_866,N_394);
and U3095 (N_3095,N_487,N_909);
and U3096 (N_3096,N_2075,N_396);
nand U3097 (N_3097,N_2903,N_1570);
xnor U3098 (N_3098,N_2918,N_2463);
or U3099 (N_3099,N_2006,N_263);
or U3100 (N_3100,N_745,N_2110);
nand U3101 (N_3101,N_2367,N_573);
xnor U3102 (N_3102,N_539,N_1555);
or U3103 (N_3103,N_1722,N_164);
nor U3104 (N_3104,N_1309,N_1255);
or U3105 (N_3105,N_163,N_1620);
and U3106 (N_3106,N_2009,N_964);
nor U3107 (N_3107,N_39,N_534);
or U3108 (N_3108,N_642,N_2731);
xor U3109 (N_3109,N_1336,N_138);
and U3110 (N_3110,N_1631,N_1385);
nor U3111 (N_3111,N_384,N_18);
nor U3112 (N_3112,N_1833,N_1977);
or U3113 (N_3113,N_1128,N_1068);
nor U3114 (N_3114,N_1531,N_136);
nor U3115 (N_3115,N_2458,N_1167);
nand U3116 (N_3116,N_494,N_468);
nand U3117 (N_3117,N_2876,N_649);
and U3118 (N_3118,N_739,N_1522);
or U3119 (N_3119,N_566,N_2692);
nand U3120 (N_3120,N_2590,N_2586);
or U3121 (N_3121,N_1931,N_2474);
and U3122 (N_3122,N_2657,N_1376);
and U3123 (N_3123,N_1590,N_1653);
and U3124 (N_3124,N_1891,N_1840);
nand U3125 (N_3125,N_2572,N_1260);
and U3126 (N_3126,N_2607,N_740);
xnor U3127 (N_3127,N_686,N_225);
nor U3128 (N_3128,N_1566,N_541);
nand U3129 (N_3129,N_1476,N_630);
nor U3130 (N_3130,N_1041,N_2995);
nor U3131 (N_3131,N_283,N_485);
and U3132 (N_3132,N_1878,N_220);
nor U3133 (N_3133,N_2166,N_1428);
nand U3134 (N_3134,N_2709,N_650);
or U3135 (N_3135,N_1787,N_2958);
nor U3136 (N_3136,N_236,N_197);
or U3137 (N_3137,N_1697,N_1633);
nand U3138 (N_3138,N_2581,N_319);
xor U3139 (N_3139,N_2564,N_1601);
or U3140 (N_3140,N_2852,N_1811);
or U3141 (N_3141,N_1088,N_10);
nand U3142 (N_3142,N_951,N_1837);
or U3143 (N_3143,N_2519,N_247);
or U3144 (N_3144,N_2668,N_1434);
nor U3145 (N_3145,N_2806,N_1305);
nor U3146 (N_3146,N_611,N_1933);
xnor U3147 (N_3147,N_1728,N_2308);
xor U3148 (N_3148,N_1969,N_342);
or U3149 (N_3149,N_2611,N_2286);
nand U3150 (N_3150,N_2940,N_1859);
nor U3151 (N_3151,N_457,N_2554);
and U3152 (N_3152,N_2125,N_2031);
nand U3153 (N_3153,N_716,N_1488);
nor U3154 (N_3154,N_2071,N_2759);
or U3155 (N_3155,N_1109,N_2705);
and U3156 (N_3156,N_1169,N_2755);
nand U3157 (N_3157,N_286,N_502);
and U3158 (N_3158,N_57,N_2121);
and U3159 (N_3159,N_2100,N_2508);
and U3160 (N_3160,N_2996,N_849);
nor U3161 (N_3161,N_2691,N_776);
nand U3162 (N_3162,N_2733,N_2764);
and U3163 (N_3163,N_2521,N_1356);
or U3164 (N_3164,N_1542,N_1709);
or U3165 (N_3165,N_2485,N_2717);
or U3166 (N_3166,N_246,N_2159);
xnor U3167 (N_3167,N_704,N_2102);
or U3168 (N_3168,N_840,N_2867);
nor U3169 (N_3169,N_801,N_2236);
or U3170 (N_3170,N_1865,N_2756);
nor U3171 (N_3171,N_2863,N_2267);
and U3172 (N_3172,N_1746,N_1718);
and U3173 (N_3173,N_1702,N_2060);
xnor U3174 (N_3174,N_670,N_844);
xnor U3175 (N_3175,N_2965,N_1890);
and U3176 (N_3176,N_1788,N_907);
nand U3177 (N_3177,N_506,N_1991);
and U3178 (N_3178,N_2567,N_615);
nor U3179 (N_3179,N_2969,N_448);
nor U3180 (N_3180,N_309,N_178);
xor U3181 (N_3181,N_2956,N_1057);
and U3182 (N_3182,N_1482,N_895);
nand U3183 (N_3183,N_439,N_731);
nor U3184 (N_3184,N_2408,N_2330);
xnor U3185 (N_3185,N_2241,N_1403);
xor U3186 (N_3186,N_1821,N_1694);
or U3187 (N_3187,N_2317,N_1456);
or U3188 (N_3188,N_2594,N_2128);
nand U3189 (N_3189,N_1370,N_1976);
or U3190 (N_3190,N_1698,N_86);
nand U3191 (N_3191,N_2856,N_85);
and U3192 (N_3192,N_1142,N_1643);
or U3193 (N_3193,N_2623,N_1803);
or U3194 (N_3194,N_831,N_607);
xor U3195 (N_3195,N_84,N_1776);
and U3196 (N_3196,N_712,N_2779);
or U3197 (N_3197,N_2037,N_293);
nand U3198 (N_3198,N_706,N_2199);
and U3199 (N_3199,N_288,N_1159);
or U3200 (N_3200,N_7,N_2460);
and U3201 (N_3201,N_809,N_122);
and U3202 (N_3202,N_2329,N_1736);
nor U3203 (N_3203,N_1401,N_469);
and U3204 (N_3204,N_1300,N_2053);
or U3205 (N_3205,N_324,N_533);
and U3206 (N_3206,N_1139,N_2898);
nand U3207 (N_3207,N_2600,N_1726);
xnor U3208 (N_3208,N_1414,N_190);
xor U3209 (N_3209,N_783,N_1743);
nor U3210 (N_3210,N_671,N_860);
nand U3211 (N_3211,N_1031,N_1096);
nand U3212 (N_3212,N_998,N_2754);
nand U3213 (N_3213,N_1053,N_984);
or U3214 (N_3214,N_956,N_993);
or U3215 (N_3215,N_2095,N_1610);
and U3216 (N_3216,N_981,N_1839);
nor U3217 (N_3217,N_2365,N_258);
xor U3218 (N_3218,N_173,N_530);
xnor U3219 (N_3219,N_1193,N_2872);
and U3220 (N_3220,N_2013,N_612);
nor U3221 (N_3221,N_334,N_2550);
xor U3222 (N_3222,N_900,N_1723);
or U3223 (N_3223,N_1856,N_2750);
nand U3224 (N_3224,N_639,N_2630);
nor U3225 (N_3225,N_2338,N_2989);
nor U3226 (N_3226,N_780,N_728);
nand U3227 (N_3227,N_1972,N_2983);
nor U3228 (N_3228,N_1213,N_908);
nand U3229 (N_3229,N_1582,N_1893);
nand U3230 (N_3230,N_1734,N_2934);
and U3231 (N_3231,N_1009,N_351);
nor U3232 (N_3232,N_1742,N_373);
xor U3233 (N_3233,N_2785,N_856);
or U3234 (N_3234,N_482,N_1543);
or U3235 (N_3235,N_2813,N_1524);
or U3236 (N_3236,N_114,N_564);
xor U3237 (N_3237,N_358,N_2171);
xnor U3238 (N_3238,N_936,N_183);
xor U3239 (N_3239,N_2608,N_1804);
and U3240 (N_3240,N_1655,N_78);
or U3241 (N_3241,N_375,N_473);
or U3242 (N_3242,N_911,N_708);
xor U3243 (N_3243,N_635,N_2161);
or U3244 (N_3244,N_2484,N_2087);
xor U3245 (N_3245,N_2888,N_1155);
and U3246 (N_3246,N_2187,N_2538);
nand U3247 (N_3247,N_2835,N_520);
or U3248 (N_3248,N_1462,N_2185);
and U3249 (N_3249,N_344,N_2993);
nor U3250 (N_3250,N_2163,N_2420);
nor U3251 (N_3251,N_250,N_522);
nor U3252 (N_3252,N_490,N_2959);
nor U3253 (N_3253,N_272,N_518);
nand U3254 (N_3254,N_2857,N_2243);
nand U3255 (N_3255,N_2507,N_1616);
nand U3256 (N_3256,N_1468,N_1831);
and U3257 (N_3257,N_1382,N_374);
xor U3258 (N_3258,N_406,N_2633);
nor U3259 (N_3259,N_2052,N_484);
and U3260 (N_3260,N_462,N_254);
or U3261 (N_3261,N_2781,N_880);
and U3262 (N_3262,N_934,N_2270);
or U3263 (N_3263,N_1835,N_771);
xor U3264 (N_3264,N_2315,N_2544);
and U3265 (N_3265,N_2221,N_2268);
or U3266 (N_3266,N_698,N_1708);
nor U3267 (N_3267,N_2953,N_280);
nor U3268 (N_3268,N_2002,N_2446);
nand U3269 (N_3269,N_95,N_2703);
nand U3270 (N_3270,N_2105,N_1705);
nor U3271 (N_3271,N_843,N_2699);
nor U3272 (N_3272,N_682,N_2146);
nor U3273 (N_3273,N_1076,N_565);
or U3274 (N_3274,N_1337,N_1208);
nand U3275 (N_3275,N_2951,N_2793);
or U3276 (N_3276,N_1612,N_1780);
xnor U3277 (N_3277,N_2689,N_2305);
or U3278 (N_3278,N_231,N_590);
nor U3279 (N_3279,N_1129,N_1763);
nor U3280 (N_3280,N_2658,N_729);
and U3281 (N_3281,N_2497,N_718);
or U3282 (N_3282,N_773,N_2422);
nor U3283 (N_3283,N_2122,N_545);
and U3284 (N_3284,N_1408,N_2476);
xor U3285 (N_3285,N_837,N_17);
and U3286 (N_3286,N_1252,N_1829);
and U3287 (N_3287,N_2941,N_2260);
nor U3288 (N_3288,N_2064,N_2180);
nand U3289 (N_3289,N_2081,N_2138);
and U3290 (N_3290,N_2273,N_2576);
or U3291 (N_3291,N_2148,N_367);
and U3292 (N_3292,N_305,N_1918);
and U3293 (N_3293,N_1323,N_2530);
and U3294 (N_3294,N_2907,N_1999);
or U3295 (N_3295,N_2636,N_1502);
or U3296 (N_3296,N_972,N_1412);
nand U3297 (N_3297,N_1704,N_1945);
xor U3298 (N_3298,N_1437,N_1348);
or U3299 (N_3299,N_2787,N_174);
nand U3300 (N_3300,N_2617,N_295);
xnor U3301 (N_3301,N_2116,N_654);
and U3302 (N_3302,N_2349,N_1367);
and U3303 (N_3303,N_554,N_660);
and U3304 (N_3304,N_647,N_1699);
and U3305 (N_3305,N_583,N_2776);
nor U3306 (N_3306,N_134,N_717);
nor U3307 (N_3307,N_1556,N_2949);
or U3308 (N_3308,N_2548,N_807);
xnor U3309 (N_3309,N_1445,N_229);
nand U3310 (N_3310,N_2826,N_2275);
xnor U3311 (N_3311,N_526,N_863);
nand U3312 (N_3312,N_442,N_2078);
nand U3313 (N_3313,N_1164,N_1225);
nand U3314 (N_3314,N_204,N_232);
and U3315 (N_3315,N_2447,N_663);
or U3316 (N_3316,N_143,N_1083);
nor U3317 (N_3317,N_101,N_507);
xor U3318 (N_3318,N_1082,N_713);
xor U3319 (N_3319,N_1368,N_772);
and U3320 (N_3320,N_207,N_19);
xnor U3321 (N_3321,N_2156,N_2383);
or U3322 (N_3322,N_1559,N_2906);
nand U3323 (N_3323,N_337,N_1117);
or U3324 (N_3324,N_756,N_2024);
nor U3325 (N_3325,N_595,N_711);
and U3326 (N_3326,N_793,N_1132);
and U3327 (N_3327,N_2932,N_2975);
or U3328 (N_3328,N_2091,N_2387);
xnor U3329 (N_3329,N_2112,N_1026);
nand U3330 (N_3330,N_627,N_2864);
or U3331 (N_3331,N_1923,N_1838);
nand U3332 (N_3332,N_1966,N_301);
nand U3333 (N_3333,N_1662,N_62);
xor U3334 (N_3334,N_2526,N_976);
nand U3335 (N_3335,N_2074,N_443);
and U3336 (N_3336,N_2055,N_1395);
or U3337 (N_3337,N_808,N_1015);
xnor U3338 (N_3338,N_1272,N_2374);
nor U3339 (N_3339,N_700,N_2585);
xnor U3340 (N_3340,N_303,N_787);
nand U3341 (N_3341,N_1574,N_1325);
or U3342 (N_3342,N_2588,N_898);
and U3343 (N_3343,N_2676,N_2882);
or U3344 (N_3344,N_2802,N_2749);
or U3345 (N_3345,N_2023,N_2437);
nand U3346 (N_3346,N_1216,N_897);
and U3347 (N_3347,N_2990,N_2854);
and U3348 (N_3348,N_2780,N_139);
xor U3349 (N_3349,N_770,N_1071);
xor U3350 (N_3350,N_400,N_2923);
nor U3351 (N_3351,N_1870,N_2046);
xor U3352 (N_3352,N_1682,N_2369);
nor U3353 (N_3353,N_622,N_1140);
nand U3354 (N_3354,N_2821,N_2038);
and U3355 (N_3355,N_1518,N_491);
and U3356 (N_3356,N_267,N_2597);
or U3357 (N_3357,N_1635,N_1652);
xnor U3358 (N_3358,N_1248,N_999);
nor U3359 (N_3359,N_2825,N_2381);
or U3360 (N_3360,N_23,N_2603);
nand U3361 (N_3361,N_140,N_2090);
and U3362 (N_3362,N_2540,N_1539);
nor U3363 (N_3363,N_1398,N_1072);
and U3364 (N_3364,N_362,N_54);
or U3365 (N_3365,N_24,N_1112);
or U3366 (N_3366,N_724,N_1691);
and U3367 (N_3367,N_629,N_567);
xnor U3368 (N_3368,N_885,N_1321);
and U3369 (N_3369,N_2188,N_2223);
or U3370 (N_3370,N_1078,N_923);
xnor U3371 (N_3371,N_1625,N_2480);
nand U3372 (N_3372,N_2328,N_1191);
xor U3373 (N_3373,N_1391,N_2944);
nand U3374 (N_3374,N_1127,N_1316);
xor U3375 (N_3375,N_1417,N_1819);
or U3376 (N_3376,N_380,N_883);
nor U3377 (N_3377,N_832,N_1930);
nor U3378 (N_3378,N_2865,N_581);
nand U3379 (N_3379,N_737,N_1299);
xor U3380 (N_3380,N_2571,N_1388);
or U3381 (N_3381,N_2625,N_1680);
or U3382 (N_3382,N_2752,N_2683);
and U3383 (N_3383,N_2181,N_2282);
and U3384 (N_3384,N_1232,N_118);
or U3385 (N_3385,N_2533,N_82);
nand U3386 (N_3386,N_2829,N_2517);
or U3387 (N_3387,N_2080,N_2428);
or U3388 (N_3388,N_2306,N_1920);
nand U3389 (N_3389,N_1795,N_2690);
nand U3390 (N_3390,N_2664,N_68);
xnor U3391 (N_3391,N_2909,N_1489);
and U3392 (N_3392,N_1130,N_602);
nor U3393 (N_3393,N_151,N_2744);
xor U3394 (N_3394,N_1498,N_665);
nand U3395 (N_3395,N_407,N_2257);
nand U3396 (N_3396,N_475,N_2723);
or U3397 (N_3397,N_216,N_1800);
and U3398 (N_3398,N_763,N_901);
and U3399 (N_3399,N_1338,N_2757);
or U3400 (N_3400,N_915,N_2920);
and U3401 (N_3401,N_1901,N_13);
or U3402 (N_3402,N_2502,N_1033);
xnor U3403 (N_3403,N_1304,N_437);
nand U3404 (N_3404,N_1007,N_1150);
or U3405 (N_3405,N_2736,N_1098);
nor U3406 (N_3406,N_1809,N_1005);
nand U3407 (N_3407,N_2015,N_402);
and U3408 (N_3408,N_209,N_1032);
xnor U3409 (N_3409,N_1605,N_409);
xnor U3410 (N_3410,N_2774,N_1608);
and U3411 (N_3411,N_975,N_1251);
and U3412 (N_3412,N_2019,N_2106);
xor U3413 (N_3413,N_834,N_429);
nand U3414 (N_3414,N_794,N_2790);
nor U3415 (N_3415,N_2198,N_2596);
xor U3416 (N_3416,N_1285,N_1895);
xnor U3417 (N_3417,N_764,N_2547);
xnor U3418 (N_3418,N_2228,N_1461);
nor U3419 (N_3419,N_2409,N_2356);
nand U3420 (N_3420,N_2704,N_2927);
xor U3421 (N_3421,N_585,N_2195);
and U3422 (N_3422,N_125,N_1429);
or U3423 (N_3423,N_990,N_894);
nor U3424 (N_3424,N_2546,N_2602);
nor U3425 (N_3425,N_890,N_714);
or U3426 (N_3426,N_1409,N_1812);
or U3427 (N_3427,N_2528,N_1301);
nor U3428 (N_3428,N_2832,N_755);
xor U3429 (N_3429,N_1961,N_408);
nand U3430 (N_3430,N_1533,N_1911);
and U3431 (N_3431,N_316,N_1650);
nor U3432 (N_3432,N_683,N_2149);
nor U3433 (N_3433,N_1953,N_447);
and U3434 (N_3434,N_1739,N_2848);
nor U3435 (N_3435,N_1240,N_2461);
and U3436 (N_3436,N_420,N_1173);
xor U3437 (N_3437,N_2777,N_1897);
xor U3438 (N_3438,N_1288,N_653);
or U3439 (N_3439,N_694,N_855);
or U3440 (N_3440,N_2088,N_2845);
or U3441 (N_3441,N_2926,N_2663);
or U3442 (N_3442,N_738,N_22);
xor U3443 (N_3443,N_1310,N_548);
nand U3444 (N_3444,N_2431,N_853);
nand U3445 (N_3445,N_2604,N_2838);
nor U3446 (N_3446,N_1604,N_529);
and U3447 (N_3447,N_92,N_594);
xor U3448 (N_3448,N_1371,N_2186);
xnor U3449 (N_3449,N_2123,N_1287);
or U3450 (N_3450,N_2811,N_978);
nor U3451 (N_3451,N_1532,N_1168);
and U3452 (N_3452,N_1313,N_1174);
and U3453 (N_3453,N_2453,N_2870);
nor U3454 (N_3454,N_2534,N_165);
xor U3455 (N_3455,N_2010,N_2246);
xor U3456 (N_3456,N_2252,N_1182);
nor U3457 (N_3457,N_803,N_70);
nand U3458 (N_3458,N_2039,N_1444);
nand U3459 (N_3459,N_2721,N_1387);
and U3460 (N_3460,N_1552,N_623);
xor U3461 (N_3461,N_1629,N_2593);
nand U3462 (N_3462,N_646,N_932);
or U3463 (N_3463,N_2029,N_387);
xor U3464 (N_3464,N_1153,N_106);
nand U3465 (N_3465,N_1774,N_2890);
and U3466 (N_3466,N_356,N_1214);
or U3467 (N_3467,N_296,N_861);
nor U3468 (N_3468,N_261,N_1035);
or U3469 (N_3469,N_893,N_65);
nand U3470 (N_3470,N_600,N_1896);
nor U3471 (N_3471,N_599,N_1107);
xor U3472 (N_3472,N_638,N_1061);
or U3473 (N_3473,N_1115,N_2982);
xor U3474 (N_3474,N_2573,N_747);
or U3475 (N_3475,N_2849,N_2366);
and U3476 (N_3476,N_2889,N_2057);
nand U3477 (N_3477,N_777,N_1004);
nand U3478 (N_3478,N_1361,N_1090);
or U3479 (N_3479,N_608,N_156);
and U3480 (N_3480,N_1022,N_1714);
xor U3481 (N_3481,N_0,N_1211);
nor U3482 (N_3482,N_1772,N_73);
and U3483 (N_3483,N_188,N_1512);
nand U3484 (N_3484,N_1745,N_2232);
xnor U3485 (N_3485,N_282,N_386);
or U3486 (N_3486,N_1637,N_593);
xnor U3487 (N_3487,N_1656,N_1416);
and U3488 (N_3488,N_2363,N_2824);
nor U3489 (N_3489,N_403,N_2632);
or U3490 (N_3490,N_640,N_2795);
nor U3491 (N_3491,N_2834,N_2912);
or U3492 (N_3492,N_1575,N_658);
and U3493 (N_3493,N_514,N_2871);
nand U3494 (N_3494,N_757,N_696);
or U3495 (N_3495,N_2284,N_63);
xnor U3496 (N_3496,N_954,N_2618);
xnor U3497 (N_3497,N_2743,N_1268);
nor U3498 (N_3498,N_2210,N_876);
xor U3499 (N_3499,N_2599,N_2333);
and U3500 (N_3500,N_2552,N_2799);
or U3501 (N_3501,N_1295,N_1753);
nor U3502 (N_3502,N_2183,N_2720);
nand U3503 (N_3503,N_1506,N_2729);
xnor U3504 (N_3504,N_1449,N_414);
or U3505 (N_3505,N_2772,N_110);
nand U3506 (N_3506,N_2732,N_2584);
or U3507 (N_3507,N_877,N_2073);
and U3508 (N_3508,N_889,N_2293);
nor U3509 (N_3509,N_381,N_1243);
and U3510 (N_3510,N_1148,N_2059);
nor U3511 (N_3511,N_2807,N_774);
and U3512 (N_3512,N_1622,N_1059);
nand U3513 (N_3513,N_2957,N_2237);
or U3514 (N_3514,N_145,N_688);
or U3515 (N_3515,N_2372,N_1581);
and U3516 (N_3516,N_137,N_87);
nor U3517 (N_3517,N_742,N_1319);
xor U3518 (N_3518,N_2414,N_2288);
nand U3519 (N_3519,N_2192,N_1954);
xnor U3520 (N_3520,N_2535,N_931);
nand U3521 (N_3521,N_1711,N_2049);
or U3522 (N_3522,N_1011,N_2179);
nor U3523 (N_3523,N_2443,N_2212);
nor U3524 (N_3524,N_1621,N_2170);
nor U3525 (N_3525,N_208,N_1671);
or U3526 (N_3526,N_2376,N_2402);
nand U3527 (N_3527,N_2970,N_914);
or U3528 (N_3528,N_1647,N_899);
or U3529 (N_3529,N_2244,N_1289);
xnor U3530 (N_3530,N_1554,N_2483);
nand U3531 (N_3531,N_2150,N_2111);
and U3532 (N_3532,N_2459,N_1291);
or U3533 (N_3533,N_1207,N_433);
nor U3534 (N_3534,N_2646,N_2902);
nand U3535 (N_3535,N_1346,N_2406);
and U3536 (N_3536,N_48,N_364);
nor U3537 (N_3537,N_357,N_2649);
or U3538 (N_3538,N_2404,N_2562);
or U3539 (N_3539,N_2822,N_2285);
nand U3540 (N_3540,N_1567,N_477);
or U3541 (N_3541,N_792,N_378);
nor U3542 (N_3542,N_957,N_987);
nand U3543 (N_3543,N_1877,N_360);
or U3544 (N_3544,N_1998,N_819);
or U3545 (N_3545,N_2218,N_1241);
and U3546 (N_3546,N_1220,N_221);
nor U3547 (N_3547,N_821,N_339);
and U3548 (N_3548,N_1990,N_986);
or U3549 (N_3549,N_1204,N_2119);
or U3550 (N_3550,N_1784,N_451);
nor U3551 (N_3551,N_2935,N_1624);
xor U3552 (N_3552,N_1594,N_753);
nor U3553 (N_3553,N_1402,N_2182);
nor U3554 (N_3554,N_2708,N_1343);
or U3555 (N_3555,N_2606,N_1636);
nand U3556 (N_3556,N_2768,N_1170);
xor U3557 (N_3557,N_965,N_1049);
or U3558 (N_3558,N_515,N_865);
nor U3559 (N_3559,N_421,N_1632);
nor U3560 (N_3560,N_1589,N_59);
xor U3561 (N_3561,N_2887,N_1378);
nand U3562 (N_3562,N_715,N_50);
and U3563 (N_3563,N_1038,N_578);
nor U3564 (N_3564,N_2380,N_2309);
or U3565 (N_3565,N_882,N_405);
and U3566 (N_3566,N_2758,N_598);
and U3567 (N_3567,N_939,N_476);
xnor U3568 (N_3568,N_1453,N_2441);
xor U3569 (N_3569,N_2798,N_505);
or U3570 (N_3570,N_350,N_1703);
xor U3571 (N_3571,N_2464,N_1844);
and U3572 (N_3572,N_1854,N_77);
and U3573 (N_3573,N_1825,N_196);
xnor U3574 (N_3574,N_2575,N_2432);
nand U3575 (N_3575,N_1329,N_205);
nor U3576 (N_3576,N_1771,N_105);
nand U3577 (N_3577,N_822,N_363);
xor U3578 (N_3578,N_1431,N_2050);
and U3579 (N_3579,N_1941,N_2921);
nand U3580 (N_3580,N_1266,N_1485);
and U3581 (N_3581,N_104,N_574);
nor U3582 (N_3582,N_1983,N_1874);
nand U3583 (N_3583,N_1793,N_413);
or U3584 (N_3584,N_1946,N_1569);
xnor U3585 (N_3585,N_532,N_1239);
and U3586 (N_3586,N_2735,N_2235);
xnor U3587 (N_3587,N_1392,N_1801);
nor U3588 (N_3588,N_2628,N_925);
nor U3589 (N_3589,N_778,N_80);
nor U3590 (N_3590,N_1166,N_1905);
and U3591 (N_3591,N_2101,N_1572);
or U3592 (N_3592,N_1614,N_1750);
nand U3593 (N_3593,N_1973,N_2323);
xor U3594 (N_3594,N_2714,N_1786);
and U3595 (N_3595,N_1924,N_1227);
xor U3596 (N_3596,N_478,N_2652);
and U3597 (N_3597,N_126,N_2194);
and U3598 (N_3598,N_340,N_1820);
or U3599 (N_3599,N_953,N_2334);
nand U3600 (N_3600,N_2047,N_2650);
nor U3601 (N_3601,N_678,N_1029);
and U3602 (N_3602,N_736,N_726);
xor U3603 (N_3603,N_369,N_2438);
or U3604 (N_3604,N_2737,N_752);
nand U3605 (N_3605,N_2412,N_2434);
nand U3606 (N_3606,N_577,N_366);
and U3607 (N_3607,N_868,N_2997);
or U3608 (N_3608,N_2481,N_582);
and U3609 (N_3609,N_142,N_1183);
or U3610 (N_3610,N_561,N_1988);
xor U3611 (N_3611,N_684,N_2397);
or U3612 (N_3612,N_2964,N_962);
or U3613 (N_3613,N_2984,N_2283);
nand U3614 (N_3614,N_179,N_1981);
nand U3615 (N_3615,N_2620,N_2786);
nand U3616 (N_3616,N_702,N_1154);
xnor U3617 (N_3617,N_276,N_304);
nor U3618 (N_3618,N_750,N_538);
or U3619 (N_3619,N_547,N_2495);
or U3620 (N_3620,N_2727,N_841);
or U3621 (N_3621,N_542,N_1093);
nor U3622 (N_3622,N_1108,N_2615);
xnor U3623 (N_3623,N_230,N_982);
and U3624 (N_3624,N_169,N_869);
nor U3625 (N_3625,N_2605,N_1735);
xnor U3626 (N_3626,N_2814,N_2471);
nor U3627 (N_3627,N_2272,N_619);
and U3628 (N_3628,N_1427,N_1019);
nor U3629 (N_3629,N_64,N_940);
or U3630 (N_3630,N_1536,N_2379);
xor U3631 (N_3631,N_166,N_2390);
nor U3632 (N_3632,N_2130,N_2184);
and U3633 (N_3633,N_2980,N_2679);
xnor U3634 (N_3634,N_132,N_2880);
nor U3635 (N_3635,N_509,N_1406);
or U3636 (N_3636,N_1286,N_2730);
xnor U3637 (N_3637,N_1658,N_2843);
nor U3638 (N_3638,N_557,N_842);
nand U3639 (N_3639,N_1472,N_2800);
nor U3640 (N_3640,N_930,N_1690);
nand U3641 (N_3641,N_217,N_937);
nor U3642 (N_3642,N_2466,N_609);
nand U3643 (N_3643,N_1469,N_1349);
nor U3644 (N_3644,N_2113,N_449);
or U3645 (N_3645,N_1156,N_2142);
and U3646 (N_3646,N_1824,N_1849);
nor U3647 (N_3647,N_2899,N_12);
xnor U3648 (N_3648,N_633,N_1592);
or U3649 (N_3649,N_2477,N_2771);
or U3650 (N_3650,N_100,N_1345);
and U3651 (N_3651,N_1322,N_1092);
xor U3652 (N_3652,N_379,N_974);
nor U3653 (N_3653,N_1675,N_540);
xor U3654 (N_3654,N_1457,N_1205);
and U3655 (N_3655,N_1133,N_346);
and U3656 (N_3656,N_2160,N_2839);
nor U3657 (N_3657,N_685,N_2924);
nor U3658 (N_3658,N_2342,N_2247);
nand U3659 (N_3659,N_1330,N_2092);
nand U3660 (N_3660,N_2908,N_1450);
or U3661 (N_3661,N_2836,N_1695);
nand U3662 (N_3662,N_1467,N_710);
and U3663 (N_3663,N_913,N_2639);
or U3664 (N_3664,N_2988,N_335);
or U3665 (N_3665,N_1249,N_1192);
or U3666 (N_3666,N_928,N_1583);
and U3667 (N_3667,N_2025,N_2051);
nor U3668 (N_3668,N_1358,N_98);
or U3669 (N_3669,N_2335,N_1685);
or U3670 (N_3670,N_588,N_2570);
nand U3671 (N_3671,N_1001,N_170);
nor U3672 (N_3672,N_233,N_2026);
and U3673 (N_3673,N_2249,N_1600);
nand U3674 (N_3674,N_2747,N_1888);
and U3675 (N_3675,N_1935,N_1242);
xor U3676 (N_3676,N_2844,N_2028);
nor U3677 (N_3677,N_354,N_2936);
nor U3678 (N_3678,N_112,N_1146);
or U3679 (N_3679,N_1847,N_1571);
xnor U3680 (N_3680,N_2040,N_1335);
or U3681 (N_3681,N_1513,N_38);
xnor U3682 (N_3682,N_15,N_659);
nand U3683 (N_3683,N_2860,N_2812);
xnor U3684 (N_3684,N_219,N_2364);
nor U3685 (N_3685,N_644,N_2312);
xor U3686 (N_3686,N_1617,N_1884);
xnor U3687 (N_3687,N_669,N_1270);
and U3688 (N_3688,N_2256,N_172);
xor U3689 (N_3689,N_154,N_2700);
xnor U3690 (N_3690,N_631,N_2942);
nor U3691 (N_3691,N_2616,N_37);
xor U3692 (N_3692,N_1306,N_452);
and U3693 (N_3693,N_963,N_2345);
and U3694 (N_3694,N_1375,N_1256);
or U3695 (N_3695,N_489,N_1971);
and U3696 (N_3696,N_2879,N_1000);
xnor U3697 (N_3697,N_226,N_2027);
nand U3698 (N_3698,N_933,N_1120);
and U3699 (N_3699,N_2457,N_1904);
and U3700 (N_3700,N_781,N_1523);
and U3701 (N_3701,N_959,N_2917);
nand U3702 (N_3702,N_96,N_1700);
xor U3703 (N_3703,N_1765,N_1065);
and U3704 (N_3704,N_2893,N_198);
or U3705 (N_3705,N_2298,N_1834);
xnor U3706 (N_3706,N_606,N_701);
or U3707 (N_3707,N_1790,N_74);
xnor U3708 (N_3708,N_1919,N_1777);
nor U3709 (N_3709,N_2642,N_1792);
or U3710 (N_3710,N_674,N_1137);
nor U3711 (N_3711,N_1917,N_320);
xnor U3712 (N_3712,N_1912,N_1195);
or U3713 (N_3713,N_1480,N_31);
xor U3714 (N_3714,N_2577,N_1880);
or U3715 (N_3715,N_528,N_312);
and U3716 (N_3716,N_1796,N_1030);
nand U3717 (N_3717,N_571,N_1390);
xnor U3718 (N_3718,N_2255,N_483);
nor U3719 (N_3719,N_2549,N_1151);
and U3720 (N_3720,N_2654,N_2326);
nand U3721 (N_3721,N_251,N_1002);
and U3722 (N_3722,N_2207,N_2656);
nand U3723 (N_3723,N_1907,N_235);
or U3724 (N_3724,N_1587,N_2745);
or U3725 (N_3725,N_785,N_1339);
or U3726 (N_3726,N_2601,N_2213);
nor U3727 (N_3727,N_2482,N_102);
nor U3728 (N_3728,N_2157,N_1175);
nor U3729 (N_3729,N_1550,N_2514);
and U3730 (N_3730,N_697,N_1364);
xor U3731 (N_3731,N_1645,N_1710);
and U3732 (N_3732,N_1579,N_796);
nand U3733 (N_3733,N_2624,N_817);
or U3734 (N_3734,N_43,N_94);
or U3735 (N_3735,N_789,N_1379);
nor U3736 (N_3736,N_2922,N_2702);
nor U3737 (N_3737,N_1982,N_1184);
xnor U3738 (N_3738,N_2238,N_30);
or U3739 (N_3739,N_791,N_1103);
nor U3740 (N_3740,N_1043,N_1882);
xnor U3741 (N_3741,N_687,N_1673);
or U3742 (N_3742,N_193,N_53);
nor U3743 (N_3743,N_1706,N_501);
xnor U3744 (N_3744,N_1797,N_2271);
xor U3745 (N_3745,N_1866,N_835);
nand U3746 (N_3746,N_332,N_1669);
nor U3747 (N_3747,N_1215,N_657);
and U3748 (N_3748,N_2070,N_60);
xor U3749 (N_3749,N_1619,N_597);
or U3750 (N_3750,N_2543,N_1464);
nor U3751 (N_3751,N_1603,N_2200);
xor U3752 (N_3752,N_1484,N_2377);
nand U3753 (N_3753,N_1363,N_1613);
or U3754 (N_3754,N_300,N_672);
nor U3755 (N_3755,N_2978,N_2569);
or U3756 (N_3756,N_1236,N_2190);
nor U3757 (N_3757,N_27,N_1104);
or U3758 (N_3758,N_1386,N_2353);
nand U3759 (N_3759,N_2933,N_1496);
or U3760 (N_3760,N_2901,N_1280);
and U3761 (N_3761,N_2761,N_1290);
nor U3762 (N_3762,N_624,N_1503);
nor U3763 (N_3763,N_1707,N_1186);
nor U3764 (N_3764,N_1100,N_292);
nand U3765 (N_3765,N_1964,N_1511);
nand U3766 (N_3766,N_1188,N_2559);
xor U3767 (N_3767,N_1725,N_2313);
nor U3768 (N_3768,N_382,N_511);
xnor U3769 (N_3769,N_1607,N_1951);
nand U3770 (N_3770,N_1217,N_830);
nor U3771 (N_3771,N_1246,N_2682);
nand U3772 (N_3772,N_2327,N_2981);
and U3773 (N_3773,N_464,N_906);
and U3774 (N_3774,N_1521,N_2520);
nor U3775 (N_3775,N_238,N_486);
and U3776 (N_3776,N_1125,N_1731);
xnor U3777 (N_3777,N_1161,N_1659);
nand U3778 (N_3778,N_1421,N_415);
or U3779 (N_3779,N_690,N_1876);
or U3780 (N_3780,N_1433,N_1423);
nand U3781 (N_3781,N_329,N_2415);
and U3782 (N_3782,N_456,N_2307);
nand U3783 (N_3783,N_2439,N_1218);
or U3784 (N_3784,N_2203,N_1441);
xor U3785 (N_3785,N_2488,N_601);
nand U3786 (N_3786,N_1741,N_2357);
nor U3787 (N_3787,N_2233,N_440);
xnor U3788 (N_3788,N_1508,N_1074);
or U3789 (N_3789,N_1580,N_1853);
xnor U3790 (N_3790,N_1297,N_127);
and U3791 (N_3791,N_1171,N_874);
xnor U3792 (N_3792,N_1165,N_1606);
or U3793 (N_3793,N_1394,N_944);
nor U3794 (N_3794,N_1419,N_2352);
and U3795 (N_3795,N_948,N_2339);
xnor U3796 (N_3796,N_271,N_2866);
xnor U3797 (N_3797,N_2846,N_790);
or U3798 (N_3798,N_29,N_472);
xnor U3799 (N_3799,N_1692,N_2580);
nand U3800 (N_3800,N_2344,N_148);
or U3801 (N_3801,N_2999,N_2022);
xor U3802 (N_3802,N_307,N_1106);
xnor U3803 (N_3803,N_637,N_2666);
nand U3804 (N_3804,N_2788,N_352);
and U3805 (N_3805,N_1465,N_616);
nor U3806 (N_3806,N_1262,N_1318);
and U3807 (N_3807,N_2472,N_2211);
or U3808 (N_3808,N_1588,N_1194);
xor U3809 (N_3809,N_1762,N_1563);
nor U3810 (N_3810,N_210,N_1048);
nor U3811 (N_3811,N_1230,N_1187);
nand U3812 (N_3812,N_2855,N_1816);
nor U3813 (N_3813,N_1410,N_2395);
nand U3814 (N_3814,N_2877,N_546);
or U3815 (N_3815,N_1564,N_2598);
xnor U3816 (N_3816,N_827,N_278);
nand U3817 (N_3817,N_1025,N_311);
nor U3818 (N_3818,N_1791,N_2398);
or U3819 (N_3819,N_1080,N_2401);
and U3820 (N_3820,N_1354,N_453);
xnor U3821 (N_3821,N_1769,N_2525);
nor U3822 (N_3822,N_1661,N_1979);
xnor U3823 (N_3823,N_833,N_2486);
or U3824 (N_3824,N_1273,N_1963);
or U3825 (N_3825,N_2043,N_370);
nand U3826 (N_3826,N_2152,N_1341);
or U3827 (N_3827,N_1003,N_550);
xnor U3828 (N_3828,N_1827,N_2176);
xor U3829 (N_3829,N_2878,N_2531);
xnor U3830 (N_3830,N_376,N_2214);
xnor U3831 (N_3831,N_1328,N_1850);
xnor U3832 (N_3832,N_2578,N_2225);
nand U3833 (N_3833,N_2452,N_2943);
or U3834 (N_3834,N_2545,N_2892);
nor U3835 (N_3835,N_1118,N_390);
nand U3836 (N_3836,N_2433,N_2801);
and U3837 (N_3837,N_1123,N_2451);
nand U3838 (N_3838,N_2609,N_1069);
nor U3839 (N_3839,N_2189,N_782);
and U3840 (N_3840,N_2399,N_1925);
and U3841 (N_3841,N_317,N_643);
nor U3842 (N_3842,N_1642,N_826);
xnor U3843 (N_3843,N_2579,N_1006);
and U3844 (N_3844,N_553,N_2910);
xor U3845 (N_3845,N_1224,N_260);
or U3846 (N_3846,N_575,N_1611);
or U3847 (N_3847,N_2206,N_969);
nand U3848 (N_3848,N_2322,N_1717);
or U3849 (N_3849,N_1312,N_2020);
nor U3850 (N_3850,N_2741,N_2318);
and U3851 (N_3851,N_786,N_257);
and U3852 (N_3852,N_1491,N_436);
or U3853 (N_3853,N_1626,N_1425);
and U3854 (N_3854,N_1679,N_748);
or U3855 (N_3855,N_441,N_2828);
nor U3856 (N_3856,N_2425,N_2392);
and U3857 (N_3857,N_2217,N_287);
nand U3858 (N_3858,N_395,N_2694);
nand U3859 (N_3859,N_1598,N_2904);
xor U3860 (N_3860,N_1956,N_2201);
xnor U3861 (N_3861,N_1676,N_1903);
nand U3862 (N_3862,N_1396,N_1932);
nand U3863 (N_3863,N_535,N_1374);
nand U3864 (N_3864,N_2841,N_1501);
and U3865 (N_3865,N_1975,N_980);
nor U3866 (N_3866,N_1284,N_1970);
or U3867 (N_3867,N_2725,N_662);
nor U3868 (N_3868,N_1926,N_1770);
or U3869 (N_3869,N_187,N_107);
or U3870 (N_3870,N_1798,N_1768);
nor U3871 (N_3871,N_811,N_153);
nor U3872 (N_3872,N_2266,N_2487);
nand U3873 (N_3873,N_810,N_72);
or U3874 (N_3874,N_2518,N_2222);
nor U3875 (N_3875,N_1681,N_199);
nand U3876 (N_3876,N_2016,N_610);
and U3877 (N_3877,N_2394,N_614);
and U3878 (N_3878,N_503,N_744);
nor U3879 (N_3879,N_760,N_2097);
and U3880 (N_3880,N_499,N_2386);
and U3881 (N_3881,N_1237,N_129);
xnor U3882 (N_3882,N_1263,N_20);
nor U3883 (N_3883,N_203,N_2036);
or U3884 (N_3884,N_2468,N_800);
xor U3885 (N_3885,N_2137,N_338);
nor U3886 (N_3886,N_498,N_977);
or U3887 (N_3887,N_410,N_241);
or U3888 (N_3888,N_1052,N_2655);
or U3889 (N_3889,N_1628,N_1027);
or U3890 (N_3890,N_1460,N_1916);
and U3891 (N_3891,N_2582,N_90);
nor U3892 (N_3892,N_2930,N_119);
and U3893 (N_3893,N_1906,N_2819);
and U3894 (N_3894,N_1677,N_1715);
nand U3895 (N_3895,N_2144,N_2896);
nand U3896 (N_3896,N_69,N_751);
or U3897 (N_3897,N_2715,N_2042);
and U3898 (N_3898,N_784,N_385);
or U3899 (N_3899,N_1993,N_543);
nor U3900 (N_3900,N_2929,N_1063);
or U3901 (N_3901,N_181,N_2175);
nor U3902 (N_3902,N_2003,N_471);
and U3903 (N_3903,N_2454,N_2641);
nand U3904 (N_3904,N_2316,N_1020);
nand U3905 (N_3905,N_1389,N_2331);
nand U3906 (N_3906,N_1326,N_1949);
or U3907 (N_3907,N_1018,N_1206);
nor U3908 (N_3908,N_1311,N_2680);
nor U3909 (N_3909,N_1965,N_1596);
nand U3910 (N_3910,N_1623,N_2048);
nand U3911 (N_3911,N_1828,N_2808);
or U3912 (N_3912,N_1892,N_1757);
nor U3913 (N_3913,N_185,N_2391);
and U3914 (N_3914,N_2587,N_988);
or U3915 (N_3915,N_2204,N_2136);
and U3916 (N_3916,N_1799,N_767);
nor U3917 (N_3917,N_2269,N_2361);
nor U3918 (N_3918,N_1477,N_149);
nand U3919 (N_3919,N_2411,N_416);
nand U3920 (N_3920,N_391,N_1599);
and U3921 (N_3921,N_1448,N_1940);
or U3922 (N_3922,N_2230,N_1823);
xor U3923 (N_3923,N_1573,N_1898);
nand U3924 (N_3924,N_465,N_2129);
and U3925 (N_3925,N_1864,N_2478);
and U3926 (N_3926,N_1576,N_2972);
nand U3927 (N_3927,N_661,N_495);
and U3928 (N_3928,N_435,N_2529);
xor U3929 (N_3929,N_1271,N_958);
or U3930 (N_3930,N_2510,N_1651);
and U3931 (N_3931,N_1727,N_1250);
or U3932 (N_3932,N_2589,N_2127);
nand U3933 (N_3933,N_2007,N_1922);
xor U3934 (N_3934,N_568,N_1440);
and U3935 (N_3935,N_1245,N_2224);
or U3936 (N_3936,N_2169,N_2231);
and U3937 (N_3937,N_2987,N_992);
xnor U3938 (N_3938,N_2076,N_2032);
xnor U3939 (N_3939,N_592,N_2429);
nor U3940 (N_3940,N_2062,N_870);
xor U3941 (N_3941,N_2340,N_2005);
and U3942 (N_3942,N_632,N_1347);
and U3943 (N_3943,N_878,N_1411);
or U3944 (N_3944,N_1055,N_2568);
or U3945 (N_3945,N_1013,N_677);
or U3946 (N_3946,N_1942,N_2823);
xnor U3947 (N_3947,N_6,N_1927);
nand U3948 (N_3948,N_2378,N_967);
nand U3949 (N_3949,N_2004,N_2742);
nand U3950 (N_3950,N_2804,N_620);
nand U3951 (N_3951,N_2289,N_1683);
nand U3952 (N_3952,N_1314,N_2973);
nor U3953 (N_3953,N_1740,N_858);
and U3954 (N_3954,N_1996,N_1064);
and U3955 (N_3955,N_1047,N_734);
or U3956 (N_3956,N_2681,N_519);
xnor U3957 (N_3957,N_115,N_733);
nand U3958 (N_3958,N_2279,N_2358);
nor U3959 (N_3959,N_1439,N_1373);
or U3960 (N_3960,N_946,N_2619);
nand U3961 (N_3961,N_1075,N_766);
or U3962 (N_3962,N_1179,N_2991);
nand U3963 (N_3963,N_2963,N_2325);
or U3964 (N_3964,N_2537,N_345);
and U3965 (N_3965,N_2665,N_804);
and U3966 (N_3966,N_926,N_2440);
or U3967 (N_3967,N_2191,N_2058);
or U3968 (N_3968,N_2631,N_1761);
xnor U3969 (N_3969,N_1755,N_2314);
or U3970 (N_3970,N_2435,N_1939);
or U3971 (N_3971,N_727,N_11);
xnor U3972 (N_3972,N_2061,N_591);
nor U3973 (N_3973,N_2660,N_2133);
and U3974 (N_3974,N_829,N_1102);
nor U3975 (N_3975,N_1826,N_979);
xnor U3976 (N_3976,N_1767,N_589);
nand U3977 (N_3977,N_1221,N_103);
or U3978 (N_3978,N_1654,N_2859);
nor U3979 (N_3979,N_1808,N_239);
or U3980 (N_3980,N_58,N_1202);
nor U3981 (N_3981,N_613,N_513);
xor U3982 (N_3982,N_2385,N_1122);
xnor U3983 (N_3983,N_1149,N_691);
or U3984 (N_3984,N_2977,N_1754);
xor U3985 (N_3985,N_2697,N_1842);
nand U3986 (N_3986,N_2493,N_2045);
nor U3987 (N_3987,N_892,N_596);
xor U3988 (N_3988,N_579,N_1980);
xnor U3989 (N_3989,N_825,N_2897);
nand U3990 (N_3990,N_2536,N_1077);
or U3991 (N_3991,N_2669,N_584);
nor U3992 (N_3992,N_551,N_2767);
xnor U3993 (N_3993,N_2126,N_228);
nor U3994 (N_3994,N_2916,N_941);
nand U3995 (N_3995,N_1293,N_576);
xor U3996 (N_3996,N_1602,N_1910);
or U3997 (N_3997,N_2542,N_2661);
or U3998 (N_3998,N_2634,N_2968);
xnor U3999 (N_3999,N_2278,N_124);
xor U4000 (N_4000,N_1509,N_1180);
nand U4001 (N_4001,N_253,N_2290);
nor U4002 (N_4002,N_1045,N_431);
xnor U4003 (N_4003,N_2719,N_333);
and U4004 (N_4004,N_160,N_921);
or U4005 (N_4005,N_1178,N_1200);
nand U4006 (N_4006,N_177,N_144);
nand U4007 (N_4007,N_2311,N_2976);
xor U4008 (N_4008,N_2251,N_961);
nor U4009 (N_4009,N_1862,N_1887);
nor U4010 (N_4010,N_896,N_732);
nand U4011 (N_4011,N_1099,N_2216);
xnor U4012 (N_4012,N_371,N_175);
nor U4013 (N_4013,N_1360,N_1324);
nand U4014 (N_4014,N_2766,N_1782);
xor U4015 (N_4015,N_943,N_1591);
nor U4016 (N_4016,N_845,N_2971);
xor U4017 (N_4017,N_912,N_168);
xnor U4018 (N_4018,N_2948,N_79);
nor U4019 (N_4019,N_1054,N_51);
or U4020 (N_4020,N_1553,N_1519);
or U4021 (N_4021,N_1259,N_1147);
and U4022 (N_4022,N_2556,N_2030);
xnor U4023 (N_4023,N_1756,N_1586);
or U4024 (N_4024,N_1737,N_1701);
xnor U4025 (N_4025,N_277,N_1668);
xnor U4026 (N_4026,N_496,N_2202);
nor U4027 (N_4027,N_2728,N_512);
nor U4028 (N_4028,N_1008,N_2120);
xor U4029 (N_4029,N_797,N_8);
or U4030 (N_4030,N_2044,N_81);
nand U4031 (N_4031,N_676,N_1446);
nand U4032 (N_4032,N_2881,N_21);
xor U4033 (N_4033,N_1201,N_1665);
or U4034 (N_4034,N_461,N_2645);
xnor U4035 (N_4035,N_2107,N_111);
nor U4036 (N_4036,N_377,N_920);
or U4037 (N_4037,N_2817,N_735);
nor U4038 (N_4038,N_269,N_1101);
and U4039 (N_4039,N_2082,N_2818);
xor U4040 (N_4040,N_872,N_2427);
or U4041 (N_4041,N_2509,N_2869);
nor U4042 (N_4042,N_1902,N_991);
and U4043 (N_4043,N_1119,N_2205);
nor U4044 (N_4044,N_743,N_1014);
nand U4045 (N_4045,N_1021,N_1794);
xor U4046 (N_4046,N_1062,N_2063);
xnor U4047 (N_4047,N_1131,N_2118);
nand U4048 (N_4048,N_1051,N_2820);
and U4049 (N_4049,N_2099,N_1863);
nor U4050 (N_4050,N_1883,N_75);
and U4051 (N_4051,N_2716,N_1365);
xor U4052 (N_4052,N_1929,N_1034);
nor U4053 (N_4053,N_2511,N_1471);
nand U4054 (N_4054,N_2300,N_927);
or U4055 (N_4055,N_2967,N_1766);
nor U4056 (N_4056,N_955,N_2831);
xnor U4057 (N_4057,N_1418,N_1372);
xor U4058 (N_4058,N_2827,N_2638);
or U4059 (N_4059,N_2056,N_749);
xnor U4060 (N_4060,N_857,N_1493);
nor U4061 (N_4061,N_820,N_1967);
or U4062 (N_4062,N_270,N_1393);
and U4063 (N_4063,N_2840,N_1936);
or U4064 (N_4064,N_2359,N_1459);
nand U4065 (N_4065,N_186,N_1618);
or U4066 (N_4066,N_1253,N_516);
nor U4067 (N_4067,N_2114,N_1781);
and U4068 (N_4068,N_1111,N_586);
nand U4069 (N_4069,N_2505,N_1526);
or U4070 (N_4070,N_2693,N_1185);
and U4071 (N_4071,N_227,N_1841);
nor U4072 (N_4072,N_9,N_2900);
nor U4073 (N_4073,N_1950,N_815);
or U4074 (N_4074,N_2089,N_2640);
xor U4075 (N_4075,N_983,N_310);
or U4076 (N_4076,N_605,N_916);
nand U4077 (N_4077,N_1017,N_2370);
or U4078 (N_4078,N_1483,N_985);
nor U4079 (N_4079,N_1640,N_2462);
and U4080 (N_4080,N_33,N_1666);
nand U4081 (N_4081,N_290,N_812);
xor U4082 (N_4082,N_88,N_1957);
xnor U4083 (N_4083,N_2553,N_846);
nor U4084 (N_4084,N_2153,N_1724);
xor U4085 (N_4085,N_2143,N_450);
or U4086 (N_4086,N_960,N_924);
nand U4087 (N_4087,N_1351,N_2675);
and U4088 (N_4088,N_2688,N_2637);
nand U4089 (N_4089,N_1136,N_1436);
xnor U4090 (N_4090,N_2348,N_2263);
xnor U4091 (N_4091,N_1141,N_432);
nand U4092 (N_4092,N_1528,N_1764);
and U4093 (N_4093,N_570,N_2347);
and U4094 (N_4094,N_2291,N_1023);
and U4095 (N_4095,N_1693,N_2250);
nor U4096 (N_4096,N_2384,N_2469);
xor U4097 (N_4097,N_1404,N_1466);
and U4098 (N_4098,N_1229,N_2008);
nor U4099 (N_4099,N_1775,N_888);
nand U4100 (N_4100,N_1353,N_2498);
or U4101 (N_4101,N_2830,N_1369);
nor U4102 (N_4102,N_2301,N_1152);
nand U4103 (N_4103,N_2789,N_1397);
and U4104 (N_4104,N_398,N_141);
or U4105 (N_4105,N_1560,N_1231);
or U4106 (N_4106,N_2426,N_504);
nor U4107 (N_4107,N_2850,N_2847);
or U4108 (N_4108,N_813,N_942);
xnor U4109 (N_4109,N_66,N_2479);
nand U4110 (N_4110,N_2035,N_2489);
nor U4111 (N_4111,N_836,N_1124);
nand U4112 (N_4112,N_2324,N_1495);
nand U4113 (N_4113,N_1079,N_2803);
nand U4114 (N_4114,N_2018,N_2891);
or U4115 (N_4115,N_617,N_2341);
nand U4116 (N_4116,N_412,N_692);
and U4117 (N_4117,N_1042,N_1036);
and U4118 (N_4118,N_2430,N_2911);
or U4119 (N_4119,N_2450,N_1486);
xnor U4120 (N_4120,N_1585,N_113);
xnor U4121 (N_4121,N_2077,N_1487);
nor U4122 (N_4122,N_1451,N_1639);
xnor U4123 (N_4123,N_2791,N_1751);
xnor U4124 (N_4124,N_2219,N_765);
or U4125 (N_4125,N_336,N_1959);
nor U4126 (N_4126,N_1279,N_1050);
or U4127 (N_4127,N_2928,N_2167);
and U4128 (N_4128,N_99,N_1233);
and U4129 (N_4129,N_655,N_997);
or U4130 (N_4130,N_1713,N_1660);
nand U4131 (N_4131,N_741,N_2816);
xor U4132 (N_4132,N_854,N_479);
nor U4133 (N_4133,N_1836,N_2946);
or U4134 (N_4134,N_1667,N_1914);
nand U4135 (N_4135,N_1424,N_2810);
xor U4136 (N_4136,N_1851,N_1578);
nor U4137 (N_4137,N_2245,N_1873);
and U4138 (N_4138,N_1778,N_823);
nor U4139 (N_4139,N_214,N_1212);
xor U4140 (N_4140,N_1627,N_2522);
and U4141 (N_4141,N_2172,N_1359);
or U4142 (N_4142,N_2017,N_839);
nor U4143 (N_4143,N_949,N_1641);
nand U4144 (N_4144,N_1497,N_1505);
and U4145 (N_4145,N_157,N_2261);
nor U4146 (N_4146,N_2610,N_1885);
xor U4147 (N_4147,N_645,N_97);
or U4148 (N_4148,N_779,N_2931);
and U4149 (N_4149,N_281,N_2229);
nand U4150 (N_4150,N_425,N_218);
xnor U4151 (N_4151,N_2504,N_2320);
xor U4152 (N_4152,N_618,N_1377);
nand U4153 (N_4153,N_2734,N_2424);
and U4154 (N_4154,N_1320,N_2473);
or U4155 (N_4155,N_2068,N_1962);
nand U4156 (N_4156,N_206,N_2524);
nand U4157 (N_4157,N_1867,N_556);
nand U4158 (N_4158,N_1773,N_531);
or U4159 (N_4159,N_2612,N_1499);
nor U4160 (N_4160,N_2455,N_392);
or U4161 (N_4161,N_5,N_703);
nor U4162 (N_4162,N_2154,N_133);
nor U4163 (N_4163,N_176,N_2591);
nor U4164 (N_4164,N_180,N_1995);
nor U4165 (N_4165,N_1219,N_2961);
nor U4166 (N_4166,N_2351,N_695);
nand U4167 (N_4167,N_905,N_1779);
and U4168 (N_4168,N_297,N_1987);
nor U4169 (N_4169,N_2416,N_1551);
and U4170 (N_4170,N_1814,N_802);
xnor U4171 (N_4171,N_194,N_2436);
nor U4172 (N_4172,N_681,N_1858);
or U4173 (N_4173,N_1894,N_1138);
nor U4174 (N_4174,N_2673,N_2966);
and U4175 (N_4175,N_1752,N_2858);
xnor U4176 (N_4176,N_189,N_768);
xor U4177 (N_4177,N_1303,N_328);
or U4178 (N_4178,N_2139,N_549);
or U4179 (N_4179,N_862,N_1244);
or U4180 (N_4180,N_1234,N_2065);
xor U4181 (N_4181,N_798,N_2784);
and U4182 (N_4182,N_116,N_2103);
xor U4183 (N_4183,N_404,N_2227);
and U4184 (N_4184,N_2740,N_1760);
nand U4185 (N_4185,N_321,N_2382);
and U4186 (N_4186,N_1664,N_2753);
and U4187 (N_4187,N_273,N_851);
nor U4188 (N_4188,N_2952,N_1730);
and U4189 (N_4189,N_1442,N_1872);
nor U4190 (N_4190,N_167,N_44);
or U4191 (N_4191,N_1948,N_1978);
nand U4192 (N_4192,N_1097,N_1344);
nor U4193 (N_4193,N_2515,N_1366);
nor U4194 (N_4194,N_353,N_1223);
xor U4195 (N_4195,N_426,N_76);
nand U4196 (N_4196,N_1384,N_2034);
nand U4197 (N_4197,N_626,N_2539);
or U4198 (N_4198,N_2937,N_1540);
xor U4199 (N_4199,N_2234,N_347);
xor U4200 (N_4200,N_315,N_759);
xor U4201 (N_4201,N_1430,N_158);
nand U4202 (N_4202,N_2373,N_2475);
or U4203 (N_4203,N_805,N_1432);
nand U4204 (N_4204,N_2240,N_42);
nor U4205 (N_4205,N_348,N_2132);
xor U4206 (N_4206,N_1670,N_161);
nand U4207 (N_4207,N_1630,N_2659);
nand U4208 (N_4208,N_1514,N_2671);
or U4209 (N_4209,N_994,N_2294);
and U4210 (N_4210,N_47,N_1283);
nand U4211 (N_4211,N_152,N_648);
or U4212 (N_4212,N_1783,N_1520);
xor U4213 (N_4213,N_2842,N_89);
nor U4214 (N_4214,N_2945,N_2177);
nand U4215 (N_4215,N_2851,N_1087);
nor U4216 (N_4216,N_46,N_1561);
and U4217 (N_4217,N_2115,N_1937);
and U4218 (N_4218,N_291,N_1609);
xor U4219 (N_4219,N_2258,N_2096);
nor U4220 (N_4220,N_2985,N_438);
nor U4221 (N_4221,N_1992,N_1352);
xnor U4222 (N_4222,N_2319,N_1481);
xor U4223 (N_4223,N_1648,N_1438);
and U4224 (N_4224,N_2492,N_664);
nand U4225 (N_4225,N_1415,N_331);
or U4226 (N_4226,N_2748,N_500);
or U4227 (N_4227,N_2174,N_2501);
xnor U4228 (N_4228,N_1443,N_2389);
and U4229 (N_4229,N_2686,N_2592);
xor U4230 (N_4230,N_562,N_1176);
or U4231 (N_4231,N_1160,N_460);
nand U4232 (N_4232,N_689,N_2296);
and U4233 (N_4233,N_1818,N_1113);
or U4234 (N_4234,N_2894,N_2884);
xor U4235 (N_4235,N_55,N_434);
and U4236 (N_4236,N_1126,N_1802);
nor U4237 (N_4237,N_656,N_1989);
and U4238 (N_4238,N_2117,N_1516);
and U4239 (N_4239,N_2000,N_587);
or U4240 (N_4240,N_818,N_1012);
xnor U4241 (N_4241,N_1340,N_2622);
nor U4242 (N_4242,N_279,N_693);
and U4243 (N_4243,N_1507,N_2277);
nor U4244 (N_4244,N_2131,N_2321);
or U4245 (N_4245,N_1515,N_2512);
or U4246 (N_4246,N_2950,N_1749);
and U4247 (N_4247,N_365,N_1852);
nor U4248 (N_4248,N_2442,N_1947);
xor U4249 (N_4249,N_2992,N_455);
and U4250 (N_4250,N_497,N_2155);
nand U4251 (N_4251,N_2938,N_2695);
nand U4252 (N_4252,N_995,N_2555);
nand U4253 (N_4253,N_2986,N_1952);
nor U4254 (N_4254,N_2914,N_215);
or U4255 (N_4255,N_330,N_2135);
nand U4256 (N_4256,N_2722,N_2014);
or U4257 (N_4257,N_709,N_1327);
and U4258 (N_4258,N_2765,N_2769);
and U4259 (N_4259,N_1584,N_399);
and U4260 (N_4260,N_1209,N_2134);
and U4261 (N_4261,N_322,N_1535);
or U4262 (N_4262,N_1,N_2375);
nor U4263 (N_4263,N_848,N_1399);
nor U4264 (N_4264,N_1413,N_146);
or U4265 (N_4265,N_480,N_1688);
and U4266 (N_4266,N_2998,N_769);
or U4267 (N_4267,N_2713,N_222);
nor U4268 (N_4268,N_1177,N_1843);
or U4269 (N_4269,N_2701,N_1357);
nand U4270 (N_4270,N_2496,N_2647);
and U4271 (N_4271,N_2974,N_2419);
nor U4272 (N_4272,N_2239,N_1549);
xnor U4273 (N_4273,N_313,N_419);
and U4274 (N_4274,N_341,N_2770);
or U4275 (N_4275,N_730,N_1960);
nand U4276 (N_4276,N_680,N_323);
xnor U4277 (N_4277,N_36,N_1282);
nor U4278 (N_4278,N_1733,N_1644);
xor U4279 (N_4279,N_527,N_91);
nand U4280 (N_4280,N_2662,N_2627);
xor U4281 (N_4281,N_135,N_2350);
and U4282 (N_4282,N_996,N_1994);
and U4283 (N_4283,N_466,N_2560);
nor U4284 (N_4284,N_1732,N_1422);
nor U4285 (N_4285,N_1868,N_430);
nor U4286 (N_4286,N_719,N_2674);
nor U4287 (N_4287,N_237,N_2561);
nor U4288 (N_4288,N_2220,N_1235);
xor U4289 (N_4289,N_120,N_2685);
xor U4290 (N_4290,N_2861,N_45);
nor U4291 (N_4291,N_1307,N_1985);
or U4292 (N_4292,N_1238,N_2557);
nand U4293 (N_4293,N_2109,N_1548);
nand U4294 (N_4294,N_1822,N_1747);
xnor U4295 (N_4295,N_2,N_1684);
nand U4296 (N_4296,N_1056,N_2653);
nand U4297 (N_4297,N_243,N_2193);
xnor U4298 (N_4298,N_458,N_2687);
xnor U4299 (N_4299,N_422,N_762);
or U4300 (N_4300,N_563,N_2054);
xor U4301 (N_4301,N_1383,N_871);
or U4302 (N_4302,N_2140,N_2444);
nor U4303 (N_4303,N_1269,N_1070);
xor U4304 (N_4304,N_2418,N_2410);
nand U4305 (N_4305,N_938,N_1490);
nor U4306 (N_4306,N_359,N_1657);
nand U4307 (N_4307,N_368,N_83);
nor U4308 (N_4308,N_2583,N_775);
and U4309 (N_4309,N_1830,N_1500);
nor U4310 (N_4310,N_268,N_2209);
and U4311 (N_4311,N_2067,N_2124);
nor U4312 (N_4312,N_446,N_1086);
or U4313 (N_4313,N_2895,N_1198);
xor U4314 (N_4314,N_61,N_828);
nor U4315 (N_4315,N_234,N_1294);
or U4316 (N_4316,N_397,N_2033);
or U4317 (N_4317,N_274,N_1134);
xor U4318 (N_4318,N_2873,N_555);
xor U4319 (N_4319,N_1886,N_1157);
or U4320 (N_4320,N_1846,N_2684);
and U4321 (N_4321,N_2574,N_1400);
nor U4322 (N_4322,N_2470,N_2739);
and U4323 (N_4323,N_2883,N_1986);
nand U4324 (N_4324,N_2760,N_968);
xor U4325 (N_4325,N_2724,N_1143);
and U4326 (N_4326,N_2815,N_1261);
and U4327 (N_4327,N_2868,N_2644);
and U4328 (N_4328,N_325,N_262);
xor U4329 (N_4329,N_212,N_265);
nand U4330 (N_4330,N_372,N_2403);
xor U4331 (N_4331,N_2141,N_2467);
xor U4332 (N_4332,N_2955,N_2696);
or U4333 (N_4333,N_2226,N_705);
nor U4334 (N_4334,N_2792,N_850);
nand U4335 (N_4335,N_1577,N_971);
or U4336 (N_4336,N_1479,N_1094);
nor U4337 (N_4337,N_603,N_1921);
and U4338 (N_4338,N_2886,N_2565);
nor U4339 (N_4339,N_14,N_1091);
or U4340 (N_4340,N_2085,N_401);
and U4341 (N_4341,N_604,N_459);
or U4342 (N_4342,N_2862,N_2751);
nor U4343 (N_4343,N_2104,N_2421);
nand U4344 (N_4344,N_641,N_945);
nor U4345 (N_4345,N_1420,N_806);
nor U4346 (N_4346,N_1199,N_2796);
nor U4347 (N_4347,N_2853,N_2448);
or U4348 (N_4348,N_1721,N_1494);
nor U4349 (N_4349,N_2297,N_1744);
xor U4350 (N_4350,N_28,N_2905);
or U4351 (N_4351,N_725,N_625);
or U4352 (N_4352,N_256,N_2354);
xnor U4353 (N_4353,N_1470,N_2162);
xor U4354 (N_4354,N_1934,N_1492);
nor U4355 (N_4355,N_2809,N_1258);
and U4356 (N_4356,N_1172,N_1889);
nor U4357 (N_4357,N_2960,N_2168);
nand U4358 (N_4358,N_467,N_389);
or U4359 (N_4359,N_2215,N_2242);
and U4360 (N_4360,N_2494,N_652);
nor U4361 (N_4361,N_966,N_444);
and U4362 (N_4362,N_1646,N_917);
and U4363 (N_4363,N_1815,N_723);
nand U4364 (N_4364,N_1145,N_2523);
nand U4365 (N_4365,N_1196,N_1037);
nor U4366 (N_4366,N_666,N_508);
xor U4367 (N_4367,N_49,N_814);
or U4368 (N_4368,N_879,N_2196);
and U4369 (N_4369,N_2079,N_1871);
and U4370 (N_4370,N_1899,N_2388);
xnor U4371 (N_4371,N_2629,N_1634);
nor U4372 (N_4372,N_147,N_1010);
xor U4373 (N_4373,N_1158,N_2667);
nor U4374 (N_4374,N_524,N_2677);
nor U4375 (N_4375,N_2001,N_884);
nand U4376 (N_4376,N_2310,N_2264);
xor U4377 (N_4377,N_903,N_2913);
or U4378 (N_4378,N_2248,N_1264);
nand U4379 (N_4379,N_2563,N_1857);
and U4380 (N_4380,N_572,N_2302);
and U4381 (N_4381,N_298,N_838);
nor U4382 (N_4382,N_1362,N_2093);
xnor U4383 (N_4383,N_2371,N_2712);
nor U4384 (N_4384,N_2274,N_1955);
xor U4385 (N_4385,N_1562,N_1861);
xnor U4386 (N_4386,N_673,N_1504);
or U4387 (N_4387,N_2874,N_1116);
or U4388 (N_4388,N_423,N_517);
nor U4389 (N_4389,N_2164,N_891);
or U4390 (N_4390,N_510,N_463);
nor U4391 (N_4391,N_2954,N_184);
or U4392 (N_4392,N_1197,N_1355);
and U4393 (N_4393,N_1689,N_1058);
and U4394 (N_4394,N_1474,N_1044);
and U4395 (N_4395,N_523,N_2672);
and U4396 (N_4396,N_2738,N_223);
nor U4397 (N_4397,N_1228,N_1162);
xnor U4398 (N_4398,N_2086,N_211);
nor U4399 (N_4399,N_1277,N_1081);
nand U4400 (N_4400,N_1276,N_2445);
nor U4401 (N_4401,N_1317,N_1875);
xnor U4402 (N_4402,N_470,N_1203);
or U4403 (N_4403,N_200,N_754);
nand U4404 (N_4404,N_2707,N_1342);
or U4405 (N_4405,N_2782,N_2449);
nor U4406 (N_4406,N_40,N_2262);
or U4407 (N_4407,N_2280,N_559);
nor U4408 (N_4408,N_1024,N_2299);
or U4409 (N_4409,N_4,N_1455);
and U4410 (N_4410,N_2069,N_2407);
nand U4411 (N_4411,N_1785,N_171);
or U4412 (N_4412,N_2066,N_2145);
nor U4413 (N_4413,N_2465,N_2541);
nor U4414 (N_4414,N_758,N_788);
and U4415 (N_4415,N_536,N_1089);
nand U4416 (N_4416,N_667,N_1738);
xnor U4417 (N_4417,N_1663,N_2098);
xnor U4418 (N_4418,N_1748,N_1447);
nand U4419 (N_4419,N_474,N_2499);
xnor U4420 (N_4420,N_108,N_2614);
xnor U4421 (N_4421,N_2763,N_1478);
or U4422 (N_4422,N_213,N_454);
nand U4423 (N_4423,N_1546,N_2626);
nand U4424 (N_4424,N_1568,N_881);
nor U4425 (N_4425,N_1114,N_886);
xor U4426 (N_4426,N_634,N_1547);
nor U4427 (N_4427,N_248,N_2281);
nand U4428 (N_4428,N_1028,N_249);
and U4429 (N_4429,N_1473,N_2254);
xnor U4430 (N_4430,N_2678,N_2259);
xnor U4431 (N_4431,N_3,N_552);
and U4432 (N_4432,N_2456,N_2783);
xnor U4433 (N_4433,N_2368,N_1454);
and U4434 (N_4434,N_2396,N_2919);
xnor U4435 (N_4435,N_1254,N_2651);
or U4436 (N_4436,N_1452,N_1817);
nor U4437 (N_4437,N_326,N_2084);
nand U4438 (N_4438,N_121,N_2726);
xnor U4439 (N_4439,N_1958,N_2343);
nor U4440 (N_4440,N_679,N_1222);
nor U4441 (N_4441,N_1938,N_1190);
nand U4442 (N_4442,N_1073,N_492);
nand U4443 (N_4443,N_361,N_306);
nor U4444 (N_4444,N_1278,N_255);
and U4445 (N_4445,N_2915,N_191);
and U4446 (N_4446,N_2490,N_2360);
or U4447 (N_4447,N_2336,N_537);
nand U4448 (N_4448,N_388,N_67);
and U4449 (N_4449,N_481,N_427);
nand U4450 (N_4450,N_2253,N_2710);
xor U4451 (N_4451,N_2773,N_1296);
nor U4452 (N_4452,N_1565,N_2939);
or U4453 (N_4453,N_1869,N_1510);
or U4454 (N_4454,N_275,N_1517);
nand U4455 (N_4455,N_1595,N_2400);
or U4456 (N_4456,N_1805,N_343);
and U4457 (N_4457,N_2147,N_2711);
nor U4458 (N_4458,N_259,N_1135);
and U4459 (N_4459,N_1534,N_1529);
nor U4460 (N_4460,N_1181,N_488);
xnor U4461 (N_4461,N_799,N_1292);
nor U4462 (N_4462,N_2558,N_2021);
and U4463 (N_4463,N_2962,N_155);
nor U4464 (N_4464,N_2925,N_2762);
nand U4465 (N_4465,N_52,N_521);
or U4466 (N_4466,N_2775,N_2303);
xor U4467 (N_4467,N_16,N_2527);
or U4468 (N_4468,N_1267,N_1350);
nand U4469 (N_4469,N_2885,N_580);
xor U4470 (N_4470,N_904,N_525);
nand U4471 (N_4471,N_2500,N_1729);
and U4472 (N_4472,N_1879,N_25);
nand U4473 (N_4473,N_852,N_192);
xnor U4474 (N_4474,N_1525,N_34);
xnor U4475 (N_4475,N_245,N_1984);
nand U4476 (N_4476,N_1638,N_1302);
nor U4477 (N_4477,N_1860,N_35);
nand U4478 (N_4478,N_636,N_195);
and U4479 (N_4479,N_2012,N_201);
and U4480 (N_4480,N_2746,N_2265);
nand U4481 (N_4481,N_560,N_1997);
nand U4482 (N_4482,N_1832,N_1593);
nor U4483 (N_4483,N_2158,N_1405);
nand U4484 (N_4484,N_2503,N_2423);
nand U4485 (N_4485,N_355,N_1046);
nand U4486 (N_4486,N_935,N_1040);
or U4487 (N_4487,N_1475,N_919);
xnor U4488 (N_4488,N_417,N_2362);
and U4489 (N_4489,N_2346,N_2979);
nand U4490 (N_4490,N_1407,N_795);
xnor U4491 (N_4491,N_1855,N_1210);
nand U4492 (N_4492,N_1968,N_621);
or U4493 (N_4493,N_56,N_299);
nor U4494 (N_4494,N_182,N_947);
and U4495 (N_4495,N_2516,N_130);
and U4496 (N_4496,N_1687,N_2994);
nor U4497 (N_4497,N_1332,N_1597);
xnor U4498 (N_4498,N_558,N_1334);
or U4499 (N_4499,N_2643,N_859);
nor U4500 (N_4500,N_2963,N_2441);
or U4501 (N_4501,N_2845,N_2680);
or U4502 (N_4502,N_192,N_365);
xor U4503 (N_4503,N_1490,N_1806);
nor U4504 (N_4504,N_1479,N_1736);
and U4505 (N_4505,N_2244,N_368);
and U4506 (N_4506,N_742,N_1552);
nand U4507 (N_4507,N_2999,N_1393);
xnor U4508 (N_4508,N_2883,N_1646);
or U4509 (N_4509,N_726,N_2747);
and U4510 (N_4510,N_1869,N_1953);
nor U4511 (N_4511,N_2491,N_2927);
xor U4512 (N_4512,N_1681,N_1345);
xnor U4513 (N_4513,N_2813,N_2671);
xor U4514 (N_4514,N_2131,N_2935);
or U4515 (N_4515,N_860,N_187);
or U4516 (N_4516,N_295,N_2802);
and U4517 (N_4517,N_1021,N_1638);
and U4518 (N_4518,N_1558,N_347);
nor U4519 (N_4519,N_1314,N_1533);
nand U4520 (N_4520,N_1610,N_771);
xnor U4521 (N_4521,N_2951,N_2567);
nand U4522 (N_4522,N_2700,N_508);
and U4523 (N_4523,N_621,N_2997);
or U4524 (N_4524,N_617,N_2360);
xor U4525 (N_4525,N_94,N_1921);
xor U4526 (N_4526,N_937,N_253);
xor U4527 (N_4527,N_2397,N_2439);
or U4528 (N_4528,N_279,N_2014);
and U4529 (N_4529,N_2717,N_2841);
or U4530 (N_4530,N_1790,N_2377);
xnor U4531 (N_4531,N_504,N_1066);
nand U4532 (N_4532,N_1617,N_1553);
or U4533 (N_4533,N_2983,N_687);
or U4534 (N_4534,N_63,N_1381);
nand U4535 (N_4535,N_1821,N_989);
and U4536 (N_4536,N_586,N_1480);
nand U4537 (N_4537,N_444,N_1809);
or U4538 (N_4538,N_2356,N_945);
or U4539 (N_4539,N_1446,N_2341);
and U4540 (N_4540,N_1627,N_2085);
or U4541 (N_4541,N_63,N_1325);
and U4542 (N_4542,N_980,N_2139);
and U4543 (N_4543,N_2065,N_1165);
and U4544 (N_4544,N_1236,N_517);
xnor U4545 (N_4545,N_2070,N_693);
nor U4546 (N_4546,N_2659,N_2811);
nand U4547 (N_4547,N_102,N_665);
and U4548 (N_4548,N_356,N_12);
xor U4549 (N_4549,N_1853,N_1877);
and U4550 (N_4550,N_2086,N_1190);
nand U4551 (N_4551,N_251,N_626);
nor U4552 (N_4552,N_964,N_232);
nand U4553 (N_4553,N_2231,N_2089);
nor U4554 (N_4554,N_2172,N_1807);
xnor U4555 (N_4555,N_1173,N_612);
nand U4556 (N_4556,N_1749,N_2654);
or U4557 (N_4557,N_1877,N_977);
and U4558 (N_4558,N_859,N_2922);
nor U4559 (N_4559,N_1244,N_1649);
nor U4560 (N_4560,N_2891,N_307);
and U4561 (N_4561,N_1636,N_2878);
nor U4562 (N_4562,N_1122,N_2702);
and U4563 (N_4563,N_2990,N_1742);
nor U4564 (N_4564,N_719,N_1433);
or U4565 (N_4565,N_347,N_2713);
and U4566 (N_4566,N_1976,N_10);
and U4567 (N_4567,N_1030,N_676);
nor U4568 (N_4568,N_1388,N_145);
or U4569 (N_4569,N_925,N_1240);
and U4570 (N_4570,N_833,N_1555);
and U4571 (N_4571,N_456,N_2628);
and U4572 (N_4572,N_1610,N_2740);
nand U4573 (N_4573,N_2944,N_351);
xor U4574 (N_4574,N_1831,N_2575);
xor U4575 (N_4575,N_967,N_2889);
xor U4576 (N_4576,N_700,N_2436);
and U4577 (N_4577,N_57,N_332);
xor U4578 (N_4578,N_793,N_699);
nand U4579 (N_4579,N_267,N_2274);
xnor U4580 (N_4580,N_537,N_2249);
nor U4581 (N_4581,N_1537,N_908);
nor U4582 (N_4582,N_2679,N_2248);
nand U4583 (N_4583,N_1902,N_2572);
and U4584 (N_4584,N_1350,N_2927);
nand U4585 (N_4585,N_2950,N_296);
nor U4586 (N_4586,N_1332,N_1225);
and U4587 (N_4587,N_101,N_571);
xnor U4588 (N_4588,N_793,N_1414);
nor U4589 (N_4589,N_390,N_231);
and U4590 (N_4590,N_2684,N_198);
nand U4591 (N_4591,N_1564,N_658);
and U4592 (N_4592,N_2584,N_377);
nand U4593 (N_4593,N_1625,N_2048);
or U4594 (N_4594,N_480,N_70);
or U4595 (N_4595,N_1234,N_1833);
or U4596 (N_4596,N_1820,N_1516);
nor U4597 (N_4597,N_1623,N_1454);
nand U4598 (N_4598,N_755,N_2504);
or U4599 (N_4599,N_1096,N_644);
and U4600 (N_4600,N_102,N_784);
nor U4601 (N_4601,N_164,N_954);
and U4602 (N_4602,N_1478,N_1271);
nand U4603 (N_4603,N_999,N_2966);
and U4604 (N_4604,N_1197,N_1187);
or U4605 (N_4605,N_2921,N_1925);
and U4606 (N_4606,N_2842,N_2357);
or U4607 (N_4607,N_34,N_2939);
or U4608 (N_4608,N_949,N_201);
nand U4609 (N_4609,N_68,N_464);
or U4610 (N_4610,N_1409,N_130);
or U4611 (N_4611,N_1804,N_1270);
or U4612 (N_4612,N_1337,N_2532);
nand U4613 (N_4613,N_2269,N_2342);
or U4614 (N_4614,N_1238,N_1376);
nand U4615 (N_4615,N_1601,N_2911);
nor U4616 (N_4616,N_855,N_332);
and U4617 (N_4617,N_2856,N_2521);
and U4618 (N_4618,N_2515,N_1259);
nand U4619 (N_4619,N_1383,N_1141);
nor U4620 (N_4620,N_2428,N_225);
nor U4621 (N_4621,N_2871,N_1304);
nor U4622 (N_4622,N_1213,N_2820);
and U4623 (N_4623,N_296,N_716);
and U4624 (N_4624,N_2440,N_603);
nand U4625 (N_4625,N_2514,N_1442);
and U4626 (N_4626,N_648,N_2808);
xnor U4627 (N_4627,N_1845,N_853);
and U4628 (N_4628,N_2115,N_2179);
xnor U4629 (N_4629,N_2119,N_947);
or U4630 (N_4630,N_402,N_2205);
or U4631 (N_4631,N_2991,N_283);
nand U4632 (N_4632,N_2943,N_1761);
or U4633 (N_4633,N_2930,N_1447);
xor U4634 (N_4634,N_2762,N_2447);
nor U4635 (N_4635,N_95,N_90);
nor U4636 (N_4636,N_2764,N_2167);
or U4637 (N_4637,N_1415,N_2422);
and U4638 (N_4638,N_2725,N_686);
nor U4639 (N_4639,N_1340,N_984);
and U4640 (N_4640,N_1070,N_602);
nor U4641 (N_4641,N_2443,N_1855);
or U4642 (N_4642,N_72,N_2934);
xor U4643 (N_4643,N_2194,N_2413);
and U4644 (N_4644,N_424,N_1234);
xor U4645 (N_4645,N_807,N_58);
nand U4646 (N_4646,N_54,N_974);
nand U4647 (N_4647,N_2265,N_1767);
nor U4648 (N_4648,N_2616,N_2292);
nor U4649 (N_4649,N_2816,N_2232);
and U4650 (N_4650,N_773,N_956);
and U4651 (N_4651,N_312,N_980);
xor U4652 (N_4652,N_1962,N_2609);
and U4653 (N_4653,N_1459,N_2124);
or U4654 (N_4654,N_672,N_983);
nand U4655 (N_4655,N_2625,N_2369);
and U4656 (N_4656,N_2972,N_2974);
nor U4657 (N_4657,N_2884,N_58);
nor U4658 (N_4658,N_1486,N_2716);
nor U4659 (N_4659,N_1719,N_1347);
nor U4660 (N_4660,N_283,N_380);
nand U4661 (N_4661,N_1804,N_2458);
and U4662 (N_4662,N_373,N_1744);
xor U4663 (N_4663,N_485,N_2785);
nor U4664 (N_4664,N_2460,N_2819);
xor U4665 (N_4665,N_988,N_1507);
xnor U4666 (N_4666,N_1851,N_47);
xor U4667 (N_4667,N_385,N_756);
nor U4668 (N_4668,N_2492,N_1261);
and U4669 (N_4669,N_1643,N_2417);
nor U4670 (N_4670,N_392,N_625);
xor U4671 (N_4671,N_1702,N_1986);
nand U4672 (N_4672,N_2423,N_2895);
xor U4673 (N_4673,N_2261,N_2942);
and U4674 (N_4674,N_2272,N_856);
and U4675 (N_4675,N_2379,N_389);
xnor U4676 (N_4676,N_1265,N_787);
or U4677 (N_4677,N_67,N_707);
nand U4678 (N_4678,N_34,N_1063);
nor U4679 (N_4679,N_826,N_229);
nor U4680 (N_4680,N_1539,N_1171);
and U4681 (N_4681,N_1405,N_453);
and U4682 (N_4682,N_772,N_2233);
xnor U4683 (N_4683,N_687,N_2642);
and U4684 (N_4684,N_2516,N_1094);
xnor U4685 (N_4685,N_1141,N_2488);
and U4686 (N_4686,N_2044,N_96);
or U4687 (N_4687,N_1454,N_1427);
or U4688 (N_4688,N_1012,N_1600);
or U4689 (N_4689,N_853,N_2108);
nand U4690 (N_4690,N_2247,N_1982);
nand U4691 (N_4691,N_1101,N_513);
nand U4692 (N_4692,N_1169,N_1161);
or U4693 (N_4693,N_1839,N_546);
nor U4694 (N_4694,N_2225,N_1210);
xor U4695 (N_4695,N_985,N_1936);
or U4696 (N_4696,N_1522,N_1412);
or U4697 (N_4697,N_1369,N_1102);
nor U4698 (N_4698,N_793,N_1660);
and U4699 (N_4699,N_674,N_2419);
xnor U4700 (N_4700,N_2772,N_229);
nand U4701 (N_4701,N_1775,N_734);
nor U4702 (N_4702,N_2895,N_2533);
nand U4703 (N_4703,N_1307,N_263);
and U4704 (N_4704,N_2942,N_536);
nor U4705 (N_4705,N_306,N_1015);
or U4706 (N_4706,N_2547,N_736);
or U4707 (N_4707,N_1947,N_928);
nor U4708 (N_4708,N_2428,N_446);
xnor U4709 (N_4709,N_2546,N_2333);
nand U4710 (N_4710,N_2655,N_820);
and U4711 (N_4711,N_86,N_1317);
xnor U4712 (N_4712,N_1778,N_1422);
nand U4713 (N_4713,N_1854,N_2689);
nor U4714 (N_4714,N_1567,N_148);
nand U4715 (N_4715,N_871,N_1779);
or U4716 (N_4716,N_2131,N_842);
and U4717 (N_4717,N_2418,N_1544);
nand U4718 (N_4718,N_2310,N_1152);
or U4719 (N_4719,N_2352,N_2050);
xor U4720 (N_4720,N_2487,N_2361);
and U4721 (N_4721,N_591,N_372);
xor U4722 (N_4722,N_2086,N_2634);
nor U4723 (N_4723,N_857,N_593);
or U4724 (N_4724,N_2701,N_2863);
nor U4725 (N_4725,N_25,N_1501);
xnor U4726 (N_4726,N_970,N_2971);
or U4727 (N_4727,N_1981,N_572);
xor U4728 (N_4728,N_265,N_92);
and U4729 (N_4729,N_1774,N_1981);
xnor U4730 (N_4730,N_1354,N_2534);
nor U4731 (N_4731,N_2901,N_830);
nor U4732 (N_4732,N_2374,N_1348);
or U4733 (N_4733,N_2451,N_2204);
and U4734 (N_4734,N_2747,N_1532);
nor U4735 (N_4735,N_2065,N_913);
and U4736 (N_4736,N_1847,N_2490);
or U4737 (N_4737,N_1388,N_185);
nor U4738 (N_4738,N_2628,N_1186);
or U4739 (N_4739,N_2416,N_2872);
xor U4740 (N_4740,N_50,N_1644);
nand U4741 (N_4741,N_826,N_2319);
or U4742 (N_4742,N_2555,N_980);
nand U4743 (N_4743,N_1906,N_1707);
and U4744 (N_4744,N_886,N_838);
nor U4745 (N_4745,N_1964,N_2852);
xnor U4746 (N_4746,N_2710,N_220);
nand U4747 (N_4747,N_2404,N_895);
xor U4748 (N_4748,N_953,N_2251);
nand U4749 (N_4749,N_2174,N_908);
or U4750 (N_4750,N_2025,N_316);
and U4751 (N_4751,N_667,N_58);
nor U4752 (N_4752,N_2900,N_2087);
and U4753 (N_4753,N_1895,N_1575);
nand U4754 (N_4754,N_1213,N_1280);
nand U4755 (N_4755,N_327,N_1083);
or U4756 (N_4756,N_1268,N_2820);
nand U4757 (N_4757,N_439,N_1664);
nand U4758 (N_4758,N_132,N_2658);
nand U4759 (N_4759,N_2149,N_2012);
nand U4760 (N_4760,N_2501,N_2763);
nor U4761 (N_4761,N_2926,N_2848);
or U4762 (N_4762,N_2665,N_1308);
xnor U4763 (N_4763,N_2481,N_19);
nand U4764 (N_4764,N_1781,N_344);
and U4765 (N_4765,N_2350,N_2969);
nand U4766 (N_4766,N_1485,N_2316);
xor U4767 (N_4767,N_843,N_1752);
and U4768 (N_4768,N_1713,N_2447);
xnor U4769 (N_4769,N_310,N_1945);
nor U4770 (N_4770,N_766,N_1235);
xnor U4771 (N_4771,N_1119,N_2496);
nand U4772 (N_4772,N_2539,N_272);
or U4773 (N_4773,N_1819,N_2653);
or U4774 (N_4774,N_1898,N_960);
xnor U4775 (N_4775,N_1832,N_1774);
or U4776 (N_4776,N_800,N_1601);
or U4777 (N_4777,N_1148,N_770);
or U4778 (N_4778,N_122,N_2387);
nand U4779 (N_4779,N_2864,N_2840);
and U4780 (N_4780,N_1152,N_1447);
or U4781 (N_4781,N_916,N_395);
nor U4782 (N_4782,N_372,N_174);
xor U4783 (N_4783,N_110,N_2232);
xor U4784 (N_4784,N_1949,N_831);
nor U4785 (N_4785,N_1970,N_1230);
or U4786 (N_4786,N_516,N_2112);
nor U4787 (N_4787,N_36,N_1389);
nor U4788 (N_4788,N_2922,N_681);
or U4789 (N_4789,N_823,N_1972);
or U4790 (N_4790,N_2678,N_367);
and U4791 (N_4791,N_243,N_1314);
xor U4792 (N_4792,N_2095,N_2895);
nand U4793 (N_4793,N_708,N_1383);
or U4794 (N_4794,N_731,N_2081);
and U4795 (N_4795,N_2039,N_801);
nor U4796 (N_4796,N_365,N_1649);
and U4797 (N_4797,N_1788,N_2113);
nand U4798 (N_4798,N_2045,N_2247);
and U4799 (N_4799,N_640,N_2475);
nand U4800 (N_4800,N_1924,N_1033);
or U4801 (N_4801,N_2941,N_236);
xnor U4802 (N_4802,N_1964,N_685);
xnor U4803 (N_4803,N_1948,N_296);
nor U4804 (N_4804,N_2433,N_1108);
and U4805 (N_4805,N_2017,N_1353);
or U4806 (N_4806,N_1684,N_2793);
or U4807 (N_4807,N_2622,N_751);
xnor U4808 (N_4808,N_1711,N_2671);
and U4809 (N_4809,N_1488,N_2526);
nand U4810 (N_4810,N_1165,N_396);
xor U4811 (N_4811,N_2762,N_1089);
and U4812 (N_4812,N_221,N_2430);
and U4813 (N_4813,N_2940,N_180);
or U4814 (N_4814,N_816,N_1126);
nor U4815 (N_4815,N_1572,N_1555);
xnor U4816 (N_4816,N_489,N_1642);
xnor U4817 (N_4817,N_173,N_1559);
nand U4818 (N_4818,N_778,N_1015);
nand U4819 (N_4819,N_697,N_314);
xnor U4820 (N_4820,N_1114,N_1633);
nand U4821 (N_4821,N_641,N_1399);
nor U4822 (N_4822,N_869,N_53);
and U4823 (N_4823,N_1448,N_2856);
xnor U4824 (N_4824,N_1115,N_86);
and U4825 (N_4825,N_2098,N_671);
and U4826 (N_4826,N_2909,N_82);
or U4827 (N_4827,N_1939,N_422);
xnor U4828 (N_4828,N_2397,N_2613);
or U4829 (N_4829,N_1574,N_728);
and U4830 (N_4830,N_1442,N_1470);
xor U4831 (N_4831,N_2862,N_1172);
and U4832 (N_4832,N_2289,N_1796);
nor U4833 (N_4833,N_2888,N_1507);
nand U4834 (N_4834,N_528,N_1605);
and U4835 (N_4835,N_800,N_2882);
or U4836 (N_4836,N_1855,N_2875);
nor U4837 (N_4837,N_594,N_100);
xor U4838 (N_4838,N_189,N_2592);
nand U4839 (N_4839,N_2534,N_1945);
nand U4840 (N_4840,N_841,N_601);
xor U4841 (N_4841,N_641,N_1391);
nand U4842 (N_4842,N_2149,N_2646);
nand U4843 (N_4843,N_2714,N_1522);
or U4844 (N_4844,N_2919,N_2721);
and U4845 (N_4845,N_2758,N_635);
xnor U4846 (N_4846,N_2239,N_1085);
nand U4847 (N_4847,N_2287,N_1785);
and U4848 (N_4848,N_1497,N_828);
xnor U4849 (N_4849,N_116,N_1558);
nor U4850 (N_4850,N_2196,N_668);
and U4851 (N_4851,N_1608,N_902);
and U4852 (N_4852,N_1135,N_1435);
nor U4853 (N_4853,N_2615,N_2953);
nor U4854 (N_4854,N_2723,N_1904);
or U4855 (N_4855,N_649,N_2400);
and U4856 (N_4856,N_2028,N_792);
and U4857 (N_4857,N_407,N_1630);
or U4858 (N_4858,N_2008,N_662);
and U4859 (N_4859,N_2151,N_2411);
or U4860 (N_4860,N_2434,N_1455);
nand U4861 (N_4861,N_2627,N_2657);
xor U4862 (N_4862,N_2105,N_418);
xnor U4863 (N_4863,N_2588,N_1327);
or U4864 (N_4864,N_1439,N_2318);
or U4865 (N_4865,N_1454,N_398);
or U4866 (N_4866,N_2758,N_140);
nand U4867 (N_4867,N_2000,N_196);
xor U4868 (N_4868,N_958,N_553);
nor U4869 (N_4869,N_2678,N_2969);
nor U4870 (N_4870,N_168,N_1512);
nor U4871 (N_4871,N_1842,N_2028);
or U4872 (N_4872,N_1258,N_197);
nand U4873 (N_4873,N_821,N_27);
xnor U4874 (N_4874,N_2211,N_2246);
or U4875 (N_4875,N_2311,N_2253);
or U4876 (N_4876,N_1504,N_2913);
xnor U4877 (N_4877,N_1298,N_2649);
xnor U4878 (N_4878,N_238,N_2820);
and U4879 (N_4879,N_537,N_848);
or U4880 (N_4880,N_705,N_1908);
xnor U4881 (N_4881,N_1950,N_117);
xnor U4882 (N_4882,N_204,N_689);
and U4883 (N_4883,N_2297,N_1369);
or U4884 (N_4884,N_837,N_1588);
xor U4885 (N_4885,N_2439,N_2122);
and U4886 (N_4886,N_2113,N_1465);
xnor U4887 (N_4887,N_1491,N_758);
and U4888 (N_4888,N_1080,N_2279);
nor U4889 (N_4889,N_242,N_2873);
nand U4890 (N_4890,N_1350,N_609);
or U4891 (N_4891,N_983,N_1787);
nand U4892 (N_4892,N_893,N_1975);
nand U4893 (N_4893,N_2820,N_1023);
nor U4894 (N_4894,N_2348,N_2916);
xnor U4895 (N_4895,N_2826,N_1114);
nand U4896 (N_4896,N_1194,N_1001);
and U4897 (N_4897,N_713,N_997);
xor U4898 (N_4898,N_1604,N_2862);
nand U4899 (N_4899,N_1447,N_2285);
nand U4900 (N_4900,N_2125,N_914);
nand U4901 (N_4901,N_975,N_2928);
and U4902 (N_4902,N_736,N_673);
nand U4903 (N_4903,N_2982,N_1422);
or U4904 (N_4904,N_86,N_243);
xnor U4905 (N_4905,N_2895,N_2059);
or U4906 (N_4906,N_2904,N_728);
nand U4907 (N_4907,N_1145,N_138);
nor U4908 (N_4908,N_491,N_1406);
and U4909 (N_4909,N_1814,N_892);
nand U4910 (N_4910,N_2585,N_466);
xnor U4911 (N_4911,N_2161,N_63);
or U4912 (N_4912,N_2724,N_1757);
nand U4913 (N_4913,N_2413,N_1583);
nor U4914 (N_4914,N_1565,N_1329);
nor U4915 (N_4915,N_2425,N_2748);
nand U4916 (N_4916,N_1603,N_501);
or U4917 (N_4917,N_224,N_2403);
or U4918 (N_4918,N_2700,N_1917);
or U4919 (N_4919,N_699,N_2947);
nor U4920 (N_4920,N_1646,N_1189);
nand U4921 (N_4921,N_1872,N_1959);
nor U4922 (N_4922,N_2566,N_1841);
or U4923 (N_4923,N_1571,N_1717);
and U4924 (N_4924,N_2919,N_971);
or U4925 (N_4925,N_409,N_1607);
and U4926 (N_4926,N_609,N_715);
nor U4927 (N_4927,N_552,N_454);
or U4928 (N_4928,N_524,N_2202);
or U4929 (N_4929,N_807,N_866);
xnor U4930 (N_4930,N_1210,N_2772);
and U4931 (N_4931,N_333,N_794);
nand U4932 (N_4932,N_120,N_206);
nor U4933 (N_4933,N_1352,N_1033);
or U4934 (N_4934,N_2464,N_1114);
and U4935 (N_4935,N_2782,N_165);
nor U4936 (N_4936,N_2641,N_1756);
nor U4937 (N_4937,N_2866,N_1396);
and U4938 (N_4938,N_2358,N_831);
nor U4939 (N_4939,N_1220,N_720);
or U4940 (N_4940,N_2027,N_414);
xnor U4941 (N_4941,N_809,N_1156);
nand U4942 (N_4942,N_109,N_2239);
nor U4943 (N_4943,N_1214,N_988);
nor U4944 (N_4944,N_2985,N_2885);
or U4945 (N_4945,N_193,N_2275);
nand U4946 (N_4946,N_2056,N_2348);
xnor U4947 (N_4947,N_957,N_1686);
nand U4948 (N_4948,N_2755,N_920);
xnor U4949 (N_4949,N_1896,N_281);
and U4950 (N_4950,N_1292,N_2293);
and U4951 (N_4951,N_1696,N_2626);
xor U4952 (N_4952,N_2748,N_135);
xor U4953 (N_4953,N_2283,N_87);
or U4954 (N_4954,N_2515,N_644);
or U4955 (N_4955,N_1640,N_1259);
and U4956 (N_4956,N_2498,N_1576);
nand U4957 (N_4957,N_1397,N_394);
nand U4958 (N_4958,N_352,N_1423);
nor U4959 (N_4959,N_2596,N_2864);
and U4960 (N_4960,N_1354,N_227);
xnor U4961 (N_4961,N_64,N_119);
nand U4962 (N_4962,N_2436,N_1558);
or U4963 (N_4963,N_944,N_992);
nor U4964 (N_4964,N_1884,N_2516);
or U4965 (N_4965,N_1199,N_2032);
nor U4966 (N_4966,N_2572,N_629);
nand U4967 (N_4967,N_2940,N_307);
nand U4968 (N_4968,N_2449,N_1406);
nand U4969 (N_4969,N_1313,N_2262);
or U4970 (N_4970,N_1002,N_699);
nor U4971 (N_4971,N_1428,N_2435);
xnor U4972 (N_4972,N_1852,N_467);
nor U4973 (N_4973,N_822,N_1455);
and U4974 (N_4974,N_1692,N_2450);
xnor U4975 (N_4975,N_2929,N_1243);
xor U4976 (N_4976,N_90,N_1989);
nand U4977 (N_4977,N_1816,N_2190);
xnor U4978 (N_4978,N_2735,N_1751);
or U4979 (N_4979,N_2704,N_1076);
or U4980 (N_4980,N_1435,N_1329);
xnor U4981 (N_4981,N_2124,N_2985);
and U4982 (N_4982,N_1100,N_336);
nand U4983 (N_4983,N_1223,N_1330);
nor U4984 (N_4984,N_1476,N_203);
or U4985 (N_4985,N_2635,N_2714);
nand U4986 (N_4986,N_675,N_2069);
and U4987 (N_4987,N_1561,N_2879);
nand U4988 (N_4988,N_1009,N_803);
or U4989 (N_4989,N_1460,N_863);
nand U4990 (N_4990,N_483,N_2688);
nor U4991 (N_4991,N_2417,N_2335);
nor U4992 (N_4992,N_2863,N_2108);
nor U4993 (N_4993,N_1518,N_77);
nor U4994 (N_4994,N_2598,N_1083);
or U4995 (N_4995,N_1315,N_2679);
and U4996 (N_4996,N_2032,N_2242);
and U4997 (N_4997,N_1794,N_2337);
nand U4998 (N_4998,N_1265,N_863);
nor U4999 (N_4999,N_2636,N_703);
nor U5000 (N_5000,N_1966,N_2946);
or U5001 (N_5001,N_1658,N_1578);
nor U5002 (N_5002,N_376,N_1034);
and U5003 (N_5003,N_1590,N_198);
nor U5004 (N_5004,N_1496,N_1903);
nand U5005 (N_5005,N_1682,N_1844);
or U5006 (N_5006,N_1478,N_1737);
nor U5007 (N_5007,N_49,N_469);
nand U5008 (N_5008,N_1504,N_465);
nor U5009 (N_5009,N_1679,N_2666);
nand U5010 (N_5010,N_1666,N_2670);
nor U5011 (N_5011,N_2611,N_2857);
xor U5012 (N_5012,N_2646,N_1316);
or U5013 (N_5013,N_2731,N_1135);
or U5014 (N_5014,N_282,N_1458);
or U5015 (N_5015,N_2499,N_2735);
xor U5016 (N_5016,N_1347,N_1535);
nand U5017 (N_5017,N_434,N_1819);
or U5018 (N_5018,N_1733,N_2333);
and U5019 (N_5019,N_488,N_1483);
nand U5020 (N_5020,N_2783,N_1294);
xnor U5021 (N_5021,N_2663,N_1607);
nand U5022 (N_5022,N_1700,N_1454);
nand U5023 (N_5023,N_163,N_1581);
xor U5024 (N_5024,N_390,N_1692);
and U5025 (N_5025,N_2072,N_2364);
and U5026 (N_5026,N_2084,N_169);
nand U5027 (N_5027,N_1615,N_2623);
or U5028 (N_5028,N_1271,N_2154);
and U5029 (N_5029,N_2315,N_2219);
or U5030 (N_5030,N_860,N_485);
nand U5031 (N_5031,N_1941,N_757);
nand U5032 (N_5032,N_2118,N_760);
and U5033 (N_5033,N_2570,N_2225);
nor U5034 (N_5034,N_2538,N_1345);
and U5035 (N_5035,N_590,N_2384);
nor U5036 (N_5036,N_2990,N_1233);
or U5037 (N_5037,N_2327,N_1764);
nand U5038 (N_5038,N_2924,N_743);
nor U5039 (N_5039,N_318,N_1385);
xnor U5040 (N_5040,N_177,N_160);
or U5041 (N_5041,N_1692,N_274);
nand U5042 (N_5042,N_819,N_524);
and U5043 (N_5043,N_988,N_371);
xnor U5044 (N_5044,N_1162,N_2153);
and U5045 (N_5045,N_670,N_1131);
nand U5046 (N_5046,N_1043,N_155);
or U5047 (N_5047,N_665,N_2270);
xnor U5048 (N_5048,N_2994,N_1087);
and U5049 (N_5049,N_1898,N_945);
xor U5050 (N_5050,N_1883,N_1536);
nor U5051 (N_5051,N_1856,N_190);
nand U5052 (N_5052,N_37,N_998);
or U5053 (N_5053,N_1487,N_1559);
nor U5054 (N_5054,N_2705,N_1260);
nor U5055 (N_5055,N_270,N_128);
nor U5056 (N_5056,N_1586,N_963);
and U5057 (N_5057,N_197,N_58);
and U5058 (N_5058,N_570,N_2805);
nand U5059 (N_5059,N_2688,N_1252);
or U5060 (N_5060,N_2,N_1866);
or U5061 (N_5061,N_1521,N_1079);
xor U5062 (N_5062,N_2608,N_2512);
xnor U5063 (N_5063,N_59,N_1383);
or U5064 (N_5064,N_2706,N_1632);
nor U5065 (N_5065,N_457,N_224);
xnor U5066 (N_5066,N_919,N_1507);
or U5067 (N_5067,N_2819,N_1369);
xnor U5068 (N_5068,N_2916,N_356);
and U5069 (N_5069,N_1159,N_1478);
nor U5070 (N_5070,N_1383,N_1485);
and U5071 (N_5071,N_1041,N_1514);
nand U5072 (N_5072,N_2067,N_2009);
and U5073 (N_5073,N_920,N_2990);
nand U5074 (N_5074,N_2662,N_2624);
nand U5075 (N_5075,N_2988,N_418);
and U5076 (N_5076,N_38,N_1941);
nand U5077 (N_5077,N_2971,N_2600);
and U5078 (N_5078,N_367,N_1862);
xnor U5079 (N_5079,N_2683,N_2342);
and U5080 (N_5080,N_1298,N_276);
nor U5081 (N_5081,N_1913,N_1946);
or U5082 (N_5082,N_757,N_2293);
nor U5083 (N_5083,N_1036,N_2057);
and U5084 (N_5084,N_1695,N_2372);
nand U5085 (N_5085,N_1757,N_1759);
nand U5086 (N_5086,N_50,N_144);
xnor U5087 (N_5087,N_2292,N_199);
nand U5088 (N_5088,N_1425,N_2787);
or U5089 (N_5089,N_2449,N_1304);
and U5090 (N_5090,N_1415,N_753);
nor U5091 (N_5091,N_2132,N_836);
or U5092 (N_5092,N_1899,N_2249);
and U5093 (N_5093,N_996,N_2878);
xor U5094 (N_5094,N_2006,N_2585);
nor U5095 (N_5095,N_1167,N_1080);
and U5096 (N_5096,N_701,N_2103);
and U5097 (N_5097,N_2546,N_1745);
or U5098 (N_5098,N_1660,N_2921);
or U5099 (N_5099,N_2358,N_1994);
xor U5100 (N_5100,N_2359,N_1674);
nor U5101 (N_5101,N_338,N_455);
xor U5102 (N_5102,N_2993,N_542);
or U5103 (N_5103,N_1345,N_785);
nor U5104 (N_5104,N_2029,N_481);
xnor U5105 (N_5105,N_2514,N_951);
or U5106 (N_5106,N_1612,N_81);
nand U5107 (N_5107,N_1808,N_918);
nor U5108 (N_5108,N_2858,N_2899);
nor U5109 (N_5109,N_910,N_2245);
xnor U5110 (N_5110,N_1029,N_1421);
or U5111 (N_5111,N_458,N_1432);
nor U5112 (N_5112,N_2611,N_507);
and U5113 (N_5113,N_1274,N_2618);
or U5114 (N_5114,N_2400,N_1988);
nor U5115 (N_5115,N_1087,N_14);
and U5116 (N_5116,N_693,N_867);
nand U5117 (N_5117,N_1697,N_546);
nand U5118 (N_5118,N_2405,N_2012);
nand U5119 (N_5119,N_2280,N_1899);
xor U5120 (N_5120,N_1598,N_425);
nor U5121 (N_5121,N_1653,N_2550);
or U5122 (N_5122,N_54,N_944);
xor U5123 (N_5123,N_2723,N_2240);
or U5124 (N_5124,N_1432,N_131);
and U5125 (N_5125,N_1831,N_1142);
or U5126 (N_5126,N_1750,N_1092);
nor U5127 (N_5127,N_2635,N_1329);
nor U5128 (N_5128,N_1173,N_834);
nand U5129 (N_5129,N_2038,N_1958);
nor U5130 (N_5130,N_372,N_1275);
xnor U5131 (N_5131,N_1919,N_2328);
xnor U5132 (N_5132,N_1018,N_1379);
and U5133 (N_5133,N_2764,N_37);
nand U5134 (N_5134,N_1444,N_1588);
and U5135 (N_5135,N_738,N_2318);
xnor U5136 (N_5136,N_930,N_1480);
or U5137 (N_5137,N_2127,N_790);
and U5138 (N_5138,N_2269,N_1960);
nand U5139 (N_5139,N_2426,N_1290);
nor U5140 (N_5140,N_119,N_380);
nand U5141 (N_5141,N_2659,N_375);
or U5142 (N_5142,N_676,N_976);
nand U5143 (N_5143,N_873,N_1914);
and U5144 (N_5144,N_709,N_726);
or U5145 (N_5145,N_615,N_283);
nor U5146 (N_5146,N_840,N_559);
nand U5147 (N_5147,N_1628,N_968);
nor U5148 (N_5148,N_1384,N_1986);
xnor U5149 (N_5149,N_379,N_1978);
or U5150 (N_5150,N_260,N_254);
xor U5151 (N_5151,N_857,N_733);
and U5152 (N_5152,N_1646,N_1031);
or U5153 (N_5153,N_535,N_1563);
nand U5154 (N_5154,N_151,N_371);
xor U5155 (N_5155,N_2648,N_1424);
and U5156 (N_5156,N_1795,N_650);
xnor U5157 (N_5157,N_2898,N_2670);
and U5158 (N_5158,N_262,N_1567);
and U5159 (N_5159,N_1272,N_856);
xnor U5160 (N_5160,N_1784,N_2338);
nor U5161 (N_5161,N_202,N_1374);
nand U5162 (N_5162,N_1798,N_1406);
xor U5163 (N_5163,N_1771,N_2110);
nor U5164 (N_5164,N_597,N_574);
xor U5165 (N_5165,N_327,N_1351);
or U5166 (N_5166,N_865,N_1232);
or U5167 (N_5167,N_2176,N_1744);
nor U5168 (N_5168,N_2152,N_308);
xor U5169 (N_5169,N_1203,N_2414);
and U5170 (N_5170,N_2798,N_516);
nand U5171 (N_5171,N_286,N_10);
xnor U5172 (N_5172,N_958,N_2692);
and U5173 (N_5173,N_459,N_2301);
nor U5174 (N_5174,N_1638,N_842);
nor U5175 (N_5175,N_649,N_80);
or U5176 (N_5176,N_2934,N_2768);
and U5177 (N_5177,N_862,N_1716);
or U5178 (N_5178,N_1718,N_545);
xor U5179 (N_5179,N_1503,N_528);
or U5180 (N_5180,N_914,N_268);
nor U5181 (N_5181,N_894,N_2930);
and U5182 (N_5182,N_1812,N_1487);
nand U5183 (N_5183,N_473,N_1983);
nor U5184 (N_5184,N_130,N_2851);
or U5185 (N_5185,N_38,N_901);
or U5186 (N_5186,N_281,N_2643);
and U5187 (N_5187,N_510,N_2854);
nor U5188 (N_5188,N_1492,N_1512);
nand U5189 (N_5189,N_2356,N_84);
xor U5190 (N_5190,N_1218,N_1799);
xor U5191 (N_5191,N_1022,N_1464);
and U5192 (N_5192,N_205,N_574);
or U5193 (N_5193,N_850,N_2554);
and U5194 (N_5194,N_667,N_1638);
xor U5195 (N_5195,N_2175,N_1570);
nor U5196 (N_5196,N_997,N_1093);
nor U5197 (N_5197,N_2765,N_1421);
xnor U5198 (N_5198,N_855,N_2378);
and U5199 (N_5199,N_2563,N_2761);
xor U5200 (N_5200,N_642,N_1570);
or U5201 (N_5201,N_2634,N_1329);
xnor U5202 (N_5202,N_2036,N_2691);
or U5203 (N_5203,N_1853,N_806);
nand U5204 (N_5204,N_2465,N_2886);
nor U5205 (N_5205,N_2434,N_2558);
nand U5206 (N_5206,N_1884,N_618);
nor U5207 (N_5207,N_1430,N_1177);
and U5208 (N_5208,N_1671,N_1181);
or U5209 (N_5209,N_285,N_2759);
nor U5210 (N_5210,N_2830,N_1618);
nor U5211 (N_5211,N_2401,N_954);
nor U5212 (N_5212,N_1017,N_280);
xor U5213 (N_5213,N_2703,N_760);
or U5214 (N_5214,N_273,N_291);
xor U5215 (N_5215,N_459,N_1302);
nand U5216 (N_5216,N_2205,N_45);
nor U5217 (N_5217,N_517,N_1502);
nand U5218 (N_5218,N_785,N_213);
or U5219 (N_5219,N_2661,N_448);
nand U5220 (N_5220,N_2900,N_1423);
nand U5221 (N_5221,N_2211,N_275);
nor U5222 (N_5222,N_1639,N_577);
xnor U5223 (N_5223,N_1241,N_2899);
nand U5224 (N_5224,N_682,N_1428);
or U5225 (N_5225,N_664,N_408);
nor U5226 (N_5226,N_396,N_21);
nand U5227 (N_5227,N_2085,N_2490);
xnor U5228 (N_5228,N_2829,N_1532);
xor U5229 (N_5229,N_93,N_2796);
xor U5230 (N_5230,N_496,N_238);
nand U5231 (N_5231,N_161,N_1589);
nand U5232 (N_5232,N_2676,N_517);
nand U5233 (N_5233,N_2399,N_2924);
xor U5234 (N_5234,N_1639,N_1302);
xnor U5235 (N_5235,N_1428,N_1780);
or U5236 (N_5236,N_209,N_2138);
nand U5237 (N_5237,N_1015,N_2519);
xor U5238 (N_5238,N_564,N_1824);
or U5239 (N_5239,N_60,N_283);
and U5240 (N_5240,N_2013,N_2785);
or U5241 (N_5241,N_1546,N_1058);
xnor U5242 (N_5242,N_1398,N_1166);
or U5243 (N_5243,N_2631,N_1370);
or U5244 (N_5244,N_336,N_2406);
or U5245 (N_5245,N_790,N_1800);
and U5246 (N_5246,N_1309,N_1938);
nor U5247 (N_5247,N_885,N_1892);
nand U5248 (N_5248,N_2240,N_2023);
nand U5249 (N_5249,N_768,N_2247);
and U5250 (N_5250,N_2124,N_1299);
or U5251 (N_5251,N_1595,N_1933);
nand U5252 (N_5252,N_1984,N_819);
or U5253 (N_5253,N_2684,N_2840);
xnor U5254 (N_5254,N_296,N_2451);
and U5255 (N_5255,N_2339,N_2703);
xor U5256 (N_5256,N_2562,N_2852);
and U5257 (N_5257,N_2986,N_2321);
or U5258 (N_5258,N_1888,N_672);
nor U5259 (N_5259,N_1687,N_202);
and U5260 (N_5260,N_564,N_2229);
nand U5261 (N_5261,N_823,N_714);
or U5262 (N_5262,N_350,N_2463);
nand U5263 (N_5263,N_1489,N_2636);
xnor U5264 (N_5264,N_867,N_275);
or U5265 (N_5265,N_1484,N_1164);
and U5266 (N_5266,N_2256,N_2326);
or U5267 (N_5267,N_39,N_150);
and U5268 (N_5268,N_2015,N_360);
nor U5269 (N_5269,N_701,N_2635);
nor U5270 (N_5270,N_1064,N_582);
nand U5271 (N_5271,N_2259,N_1037);
and U5272 (N_5272,N_2824,N_1105);
and U5273 (N_5273,N_1746,N_1102);
nand U5274 (N_5274,N_93,N_2830);
and U5275 (N_5275,N_354,N_2546);
nor U5276 (N_5276,N_2491,N_2372);
nor U5277 (N_5277,N_2219,N_1092);
nand U5278 (N_5278,N_2402,N_1677);
and U5279 (N_5279,N_977,N_2204);
nand U5280 (N_5280,N_2115,N_1855);
nor U5281 (N_5281,N_1894,N_2547);
nor U5282 (N_5282,N_2367,N_2777);
nor U5283 (N_5283,N_2319,N_252);
and U5284 (N_5284,N_1217,N_158);
nor U5285 (N_5285,N_1681,N_1198);
or U5286 (N_5286,N_1586,N_2454);
and U5287 (N_5287,N_2154,N_837);
nand U5288 (N_5288,N_118,N_2484);
nor U5289 (N_5289,N_589,N_2757);
and U5290 (N_5290,N_1860,N_1258);
xor U5291 (N_5291,N_251,N_2104);
and U5292 (N_5292,N_1646,N_1735);
nor U5293 (N_5293,N_2558,N_1654);
nand U5294 (N_5294,N_326,N_2258);
xnor U5295 (N_5295,N_1334,N_223);
xnor U5296 (N_5296,N_1047,N_2436);
xor U5297 (N_5297,N_2532,N_1687);
xnor U5298 (N_5298,N_829,N_480);
and U5299 (N_5299,N_1498,N_1341);
and U5300 (N_5300,N_1803,N_1816);
or U5301 (N_5301,N_109,N_2516);
nand U5302 (N_5302,N_1268,N_375);
and U5303 (N_5303,N_2482,N_1060);
nand U5304 (N_5304,N_608,N_581);
or U5305 (N_5305,N_426,N_2909);
nor U5306 (N_5306,N_2836,N_591);
or U5307 (N_5307,N_77,N_486);
nand U5308 (N_5308,N_635,N_660);
and U5309 (N_5309,N_814,N_1045);
and U5310 (N_5310,N_2291,N_739);
or U5311 (N_5311,N_995,N_846);
nand U5312 (N_5312,N_1847,N_1035);
or U5313 (N_5313,N_149,N_2724);
and U5314 (N_5314,N_2507,N_421);
and U5315 (N_5315,N_2730,N_1146);
nand U5316 (N_5316,N_570,N_2384);
and U5317 (N_5317,N_1199,N_1925);
nor U5318 (N_5318,N_2873,N_2705);
nand U5319 (N_5319,N_1212,N_2476);
nor U5320 (N_5320,N_2317,N_393);
or U5321 (N_5321,N_2286,N_3);
nand U5322 (N_5322,N_1641,N_922);
and U5323 (N_5323,N_634,N_2697);
nor U5324 (N_5324,N_2368,N_705);
xor U5325 (N_5325,N_2676,N_1050);
or U5326 (N_5326,N_1645,N_450);
and U5327 (N_5327,N_2576,N_1604);
nand U5328 (N_5328,N_1673,N_1481);
nor U5329 (N_5329,N_1771,N_89);
xor U5330 (N_5330,N_1227,N_2619);
or U5331 (N_5331,N_2262,N_2591);
and U5332 (N_5332,N_322,N_2340);
or U5333 (N_5333,N_285,N_2654);
nand U5334 (N_5334,N_2343,N_1709);
and U5335 (N_5335,N_587,N_796);
and U5336 (N_5336,N_586,N_2883);
or U5337 (N_5337,N_786,N_1961);
nand U5338 (N_5338,N_901,N_1633);
and U5339 (N_5339,N_2395,N_611);
nor U5340 (N_5340,N_2339,N_2668);
xor U5341 (N_5341,N_386,N_2773);
nand U5342 (N_5342,N_1705,N_1826);
nor U5343 (N_5343,N_414,N_1906);
nand U5344 (N_5344,N_343,N_965);
or U5345 (N_5345,N_634,N_1236);
nand U5346 (N_5346,N_2365,N_1143);
nor U5347 (N_5347,N_972,N_1169);
nand U5348 (N_5348,N_103,N_1758);
xnor U5349 (N_5349,N_2543,N_1998);
nor U5350 (N_5350,N_1186,N_1635);
nor U5351 (N_5351,N_1905,N_748);
and U5352 (N_5352,N_1324,N_1015);
or U5353 (N_5353,N_1863,N_41);
and U5354 (N_5354,N_690,N_2570);
nand U5355 (N_5355,N_2358,N_469);
nor U5356 (N_5356,N_2311,N_2532);
and U5357 (N_5357,N_2538,N_1293);
nand U5358 (N_5358,N_944,N_22);
nor U5359 (N_5359,N_2788,N_2353);
and U5360 (N_5360,N_2421,N_1675);
nor U5361 (N_5361,N_807,N_2696);
or U5362 (N_5362,N_858,N_2672);
nand U5363 (N_5363,N_1187,N_1420);
xor U5364 (N_5364,N_756,N_1359);
xor U5365 (N_5365,N_1849,N_1459);
or U5366 (N_5366,N_1800,N_1592);
and U5367 (N_5367,N_1961,N_2964);
or U5368 (N_5368,N_895,N_1939);
or U5369 (N_5369,N_2633,N_471);
nand U5370 (N_5370,N_1384,N_1437);
nand U5371 (N_5371,N_2218,N_2904);
nand U5372 (N_5372,N_1879,N_632);
nor U5373 (N_5373,N_2237,N_2314);
xor U5374 (N_5374,N_79,N_2251);
nand U5375 (N_5375,N_2500,N_1938);
xnor U5376 (N_5376,N_2892,N_1240);
nor U5377 (N_5377,N_2408,N_1800);
nand U5378 (N_5378,N_2751,N_576);
or U5379 (N_5379,N_208,N_825);
xor U5380 (N_5380,N_326,N_1956);
xor U5381 (N_5381,N_938,N_2482);
and U5382 (N_5382,N_2060,N_2588);
nand U5383 (N_5383,N_577,N_400);
xnor U5384 (N_5384,N_7,N_1633);
xor U5385 (N_5385,N_2381,N_362);
and U5386 (N_5386,N_2439,N_2485);
and U5387 (N_5387,N_2745,N_1546);
xor U5388 (N_5388,N_2825,N_972);
nand U5389 (N_5389,N_1375,N_838);
nand U5390 (N_5390,N_218,N_847);
nor U5391 (N_5391,N_2342,N_1532);
or U5392 (N_5392,N_338,N_840);
or U5393 (N_5393,N_2818,N_1433);
xnor U5394 (N_5394,N_1350,N_302);
or U5395 (N_5395,N_1018,N_101);
nor U5396 (N_5396,N_2189,N_1997);
nand U5397 (N_5397,N_38,N_2037);
nand U5398 (N_5398,N_2312,N_398);
or U5399 (N_5399,N_2621,N_76);
and U5400 (N_5400,N_321,N_126);
xnor U5401 (N_5401,N_2376,N_552);
xnor U5402 (N_5402,N_2227,N_98);
xor U5403 (N_5403,N_2573,N_2582);
and U5404 (N_5404,N_1537,N_1320);
nand U5405 (N_5405,N_1529,N_23);
nor U5406 (N_5406,N_2324,N_1719);
or U5407 (N_5407,N_1277,N_138);
nand U5408 (N_5408,N_1099,N_1260);
or U5409 (N_5409,N_2803,N_676);
nand U5410 (N_5410,N_1108,N_2603);
xnor U5411 (N_5411,N_2278,N_222);
nand U5412 (N_5412,N_249,N_2803);
xnor U5413 (N_5413,N_103,N_1944);
or U5414 (N_5414,N_1782,N_2384);
and U5415 (N_5415,N_351,N_184);
and U5416 (N_5416,N_1763,N_812);
and U5417 (N_5417,N_1901,N_773);
xnor U5418 (N_5418,N_2414,N_1658);
nor U5419 (N_5419,N_2428,N_1604);
nor U5420 (N_5420,N_1226,N_2511);
nor U5421 (N_5421,N_1630,N_1090);
or U5422 (N_5422,N_1939,N_2690);
nor U5423 (N_5423,N_410,N_2250);
nor U5424 (N_5424,N_2596,N_2194);
nor U5425 (N_5425,N_2498,N_2401);
nor U5426 (N_5426,N_1278,N_1149);
or U5427 (N_5427,N_732,N_892);
xor U5428 (N_5428,N_1754,N_1173);
xnor U5429 (N_5429,N_377,N_2172);
xor U5430 (N_5430,N_1324,N_316);
nand U5431 (N_5431,N_2782,N_768);
or U5432 (N_5432,N_1911,N_2335);
nand U5433 (N_5433,N_2860,N_818);
nor U5434 (N_5434,N_1823,N_2457);
xnor U5435 (N_5435,N_1404,N_2978);
or U5436 (N_5436,N_1224,N_2807);
xnor U5437 (N_5437,N_2097,N_2637);
and U5438 (N_5438,N_2050,N_2579);
xnor U5439 (N_5439,N_1657,N_1596);
nand U5440 (N_5440,N_464,N_2449);
or U5441 (N_5441,N_2371,N_2627);
nor U5442 (N_5442,N_235,N_526);
or U5443 (N_5443,N_2632,N_302);
and U5444 (N_5444,N_1320,N_2836);
nor U5445 (N_5445,N_992,N_1349);
xor U5446 (N_5446,N_1384,N_2689);
xnor U5447 (N_5447,N_1244,N_1005);
or U5448 (N_5448,N_1027,N_2947);
and U5449 (N_5449,N_568,N_2217);
xnor U5450 (N_5450,N_2194,N_1390);
xnor U5451 (N_5451,N_280,N_2964);
or U5452 (N_5452,N_1120,N_999);
or U5453 (N_5453,N_2746,N_380);
and U5454 (N_5454,N_2827,N_2031);
or U5455 (N_5455,N_2738,N_952);
or U5456 (N_5456,N_1477,N_2714);
and U5457 (N_5457,N_2988,N_2299);
or U5458 (N_5458,N_1491,N_1689);
nand U5459 (N_5459,N_2982,N_2561);
or U5460 (N_5460,N_2431,N_1659);
and U5461 (N_5461,N_2497,N_250);
nor U5462 (N_5462,N_2206,N_2828);
or U5463 (N_5463,N_1993,N_1246);
xnor U5464 (N_5464,N_225,N_1334);
and U5465 (N_5465,N_2438,N_2963);
and U5466 (N_5466,N_2112,N_1170);
or U5467 (N_5467,N_152,N_1063);
nor U5468 (N_5468,N_2425,N_2486);
or U5469 (N_5469,N_197,N_420);
or U5470 (N_5470,N_1209,N_2490);
nand U5471 (N_5471,N_1120,N_2608);
xor U5472 (N_5472,N_1288,N_1800);
xor U5473 (N_5473,N_1946,N_2407);
or U5474 (N_5474,N_2039,N_1319);
and U5475 (N_5475,N_761,N_1722);
xnor U5476 (N_5476,N_1230,N_2050);
nor U5477 (N_5477,N_1571,N_2613);
and U5478 (N_5478,N_2020,N_1261);
and U5479 (N_5479,N_239,N_121);
xnor U5480 (N_5480,N_179,N_114);
nor U5481 (N_5481,N_2914,N_343);
xor U5482 (N_5482,N_547,N_1658);
or U5483 (N_5483,N_154,N_2205);
nand U5484 (N_5484,N_2766,N_2972);
xnor U5485 (N_5485,N_2521,N_534);
xor U5486 (N_5486,N_1238,N_872);
or U5487 (N_5487,N_2749,N_997);
nand U5488 (N_5488,N_315,N_2905);
or U5489 (N_5489,N_711,N_2903);
nand U5490 (N_5490,N_335,N_1417);
and U5491 (N_5491,N_394,N_1581);
and U5492 (N_5492,N_1976,N_1882);
xnor U5493 (N_5493,N_68,N_409);
nor U5494 (N_5494,N_1326,N_1801);
and U5495 (N_5495,N_1484,N_2368);
or U5496 (N_5496,N_934,N_2730);
xor U5497 (N_5497,N_1223,N_852);
nand U5498 (N_5498,N_2319,N_2558);
xnor U5499 (N_5499,N_2682,N_1046);
xnor U5500 (N_5500,N_524,N_972);
xnor U5501 (N_5501,N_1481,N_2657);
nand U5502 (N_5502,N_1905,N_2264);
and U5503 (N_5503,N_2795,N_2400);
and U5504 (N_5504,N_2568,N_2367);
nor U5505 (N_5505,N_222,N_1361);
or U5506 (N_5506,N_1406,N_1907);
nor U5507 (N_5507,N_2917,N_1234);
xor U5508 (N_5508,N_911,N_1054);
and U5509 (N_5509,N_323,N_346);
and U5510 (N_5510,N_1516,N_2071);
nand U5511 (N_5511,N_2241,N_414);
nor U5512 (N_5512,N_354,N_701);
and U5513 (N_5513,N_2081,N_2833);
nor U5514 (N_5514,N_626,N_2277);
or U5515 (N_5515,N_2660,N_2441);
nand U5516 (N_5516,N_2230,N_2739);
nor U5517 (N_5517,N_2037,N_1883);
nand U5518 (N_5518,N_2485,N_2149);
nor U5519 (N_5519,N_1024,N_2957);
nand U5520 (N_5520,N_461,N_2862);
nor U5521 (N_5521,N_2793,N_176);
nor U5522 (N_5522,N_2835,N_1588);
and U5523 (N_5523,N_1587,N_1982);
nand U5524 (N_5524,N_2335,N_1668);
or U5525 (N_5525,N_1374,N_1450);
nor U5526 (N_5526,N_1754,N_2632);
and U5527 (N_5527,N_2150,N_220);
or U5528 (N_5528,N_872,N_1575);
and U5529 (N_5529,N_2432,N_2416);
xor U5530 (N_5530,N_1277,N_2997);
nor U5531 (N_5531,N_1883,N_1559);
nand U5532 (N_5532,N_2754,N_1563);
and U5533 (N_5533,N_2444,N_2778);
and U5534 (N_5534,N_1452,N_1140);
xor U5535 (N_5535,N_2222,N_1724);
nor U5536 (N_5536,N_1380,N_1997);
or U5537 (N_5537,N_2718,N_730);
xnor U5538 (N_5538,N_1899,N_519);
nand U5539 (N_5539,N_1426,N_103);
nand U5540 (N_5540,N_2386,N_2707);
nor U5541 (N_5541,N_466,N_541);
and U5542 (N_5542,N_2730,N_128);
and U5543 (N_5543,N_838,N_1231);
xor U5544 (N_5544,N_1212,N_2531);
or U5545 (N_5545,N_2393,N_916);
nand U5546 (N_5546,N_382,N_1141);
and U5547 (N_5547,N_655,N_1477);
nor U5548 (N_5548,N_1358,N_1196);
and U5549 (N_5549,N_2063,N_1438);
or U5550 (N_5550,N_1882,N_134);
nand U5551 (N_5551,N_2627,N_2581);
nor U5552 (N_5552,N_2227,N_2709);
xnor U5553 (N_5553,N_2258,N_598);
nor U5554 (N_5554,N_1361,N_2932);
nand U5555 (N_5555,N_308,N_1756);
nand U5556 (N_5556,N_1337,N_638);
and U5557 (N_5557,N_1477,N_946);
nor U5558 (N_5558,N_996,N_2649);
xor U5559 (N_5559,N_1662,N_2024);
and U5560 (N_5560,N_1156,N_2582);
and U5561 (N_5561,N_2474,N_1609);
nor U5562 (N_5562,N_2242,N_1421);
and U5563 (N_5563,N_2483,N_2407);
xnor U5564 (N_5564,N_828,N_2386);
nand U5565 (N_5565,N_2652,N_78);
nor U5566 (N_5566,N_2827,N_458);
xor U5567 (N_5567,N_2489,N_448);
xor U5568 (N_5568,N_2224,N_2072);
and U5569 (N_5569,N_2105,N_1610);
nand U5570 (N_5570,N_111,N_825);
nand U5571 (N_5571,N_2909,N_2391);
nor U5572 (N_5572,N_441,N_1504);
and U5573 (N_5573,N_2952,N_1294);
nand U5574 (N_5574,N_34,N_1284);
nor U5575 (N_5575,N_2531,N_811);
or U5576 (N_5576,N_502,N_187);
xnor U5577 (N_5577,N_790,N_1405);
and U5578 (N_5578,N_2072,N_875);
nor U5579 (N_5579,N_2518,N_2610);
nor U5580 (N_5580,N_2695,N_701);
or U5581 (N_5581,N_870,N_2226);
nand U5582 (N_5582,N_1998,N_2684);
and U5583 (N_5583,N_2886,N_682);
or U5584 (N_5584,N_333,N_858);
and U5585 (N_5585,N_2424,N_2715);
nor U5586 (N_5586,N_863,N_1043);
and U5587 (N_5587,N_2260,N_578);
nand U5588 (N_5588,N_1652,N_1207);
and U5589 (N_5589,N_2029,N_781);
nand U5590 (N_5590,N_2946,N_1221);
nor U5591 (N_5591,N_2056,N_2605);
nor U5592 (N_5592,N_372,N_1937);
or U5593 (N_5593,N_1361,N_1445);
or U5594 (N_5594,N_2698,N_1479);
nand U5595 (N_5595,N_1101,N_2963);
nand U5596 (N_5596,N_2450,N_1917);
nor U5597 (N_5597,N_328,N_639);
nor U5598 (N_5598,N_1358,N_2475);
nand U5599 (N_5599,N_732,N_2993);
xor U5600 (N_5600,N_1297,N_69);
or U5601 (N_5601,N_1740,N_1229);
and U5602 (N_5602,N_709,N_2797);
and U5603 (N_5603,N_2743,N_2033);
or U5604 (N_5604,N_533,N_1278);
nor U5605 (N_5605,N_1574,N_784);
nand U5606 (N_5606,N_175,N_1979);
nand U5607 (N_5607,N_1191,N_2127);
nor U5608 (N_5608,N_206,N_581);
or U5609 (N_5609,N_59,N_945);
nor U5610 (N_5610,N_353,N_283);
nor U5611 (N_5611,N_2876,N_152);
nand U5612 (N_5612,N_2356,N_1892);
nor U5613 (N_5613,N_1585,N_1207);
xor U5614 (N_5614,N_137,N_1399);
and U5615 (N_5615,N_639,N_1343);
nor U5616 (N_5616,N_2559,N_1384);
and U5617 (N_5617,N_2998,N_1445);
or U5618 (N_5618,N_383,N_1225);
nand U5619 (N_5619,N_1741,N_1170);
xor U5620 (N_5620,N_177,N_679);
and U5621 (N_5621,N_1581,N_2590);
or U5622 (N_5622,N_1250,N_1631);
or U5623 (N_5623,N_2729,N_740);
or U5624 (N_5624,N_1269,N_2827);
nor U5625 (N_5625,N_849,N_1535);
or U5626 (N_5626,N_958,N_84);
nand U5627 (N_5627,N_2,N_2367);
xnor U5628 (N_5628,N_644,N_627);
xor U5629 (N_5629,N_1836,N_279);
or U5630 (N_5630,N_2727,N_805);
nand U5631 (N_5631,N_1942,N_1146);
nand U5632 (N_5632,N_1958,N_2291);
and U5633 (N_5633,N_2617,N_2724);
nor U5634 (N_5634,N_2408,N_2306);
or U5635 (N_5635,N_2976,N_1307);
nand U5636 (N_5636,N_1809,N_18);
or U5637 (N_5637,N_870,N_2198);
nand U5638 (N_5638,N_1697,N_650);
nor U5639 (N_5639,N_2413,N_2080);
nor U5640 (N_5640,N_2256,N_1722);
nor U5641 (N_5641,N_2963,N_395);
or U5642 (N_5642,N_211,N_1826);
and U5643 (N_5643,N_1043,N_267);
and U5644 (N_5644,N_2599,N_2699);
and U5645 (N_5645,N_2611,N_37);
and U5646 (N_5646,N_1738,N_2812);
nand U5647 (N_5647,N_2235,N_1910);
and U5648 (N_5648,N_2083,N_812);
nand U5649 (N_5649,N_2722,N_1153);
nand U5650 (N_5650,N_2765,N_227);
nand U5651 (N_5651,N_2309,N_1335);
or U5652 (N_5652,N_988,N_611);
and U5653 (N_5653,N_482,N_350);
xor U5654 (N_5654,N_191,N_1208);
nor U5655 (N_5655,N_929,N_2355);
or U5656 (N_5656,N_1161,N_2778);
or U5657 (N_5657,N_747,N_1858);
xnor U5658 (N_5658,N_278,N_1290);
nand U5659 (N_5659,N_993,N_370);
nand U5660 (N_5660,N_2458,N_2043);
nor U5661 (N_5661,N_2248,N_2946);
nor U5662 (N_5662,N_420,N_2100);
xnor U5663 (N_5663,N_2706,N_2057);
and U5664 (N_5664,N_1539,N_2074);
and U5665 (N_5665,N_1397,N_857);
nand U5666 (N_5666,N_1549,N_2339);
or U5667 (N_5667,N_2937,N_2489);
nor U5668 (N_5668,N_1362,N_474);
and U5669 (N_5669,N_1421,N_971);
xnor U5670 (N_5670,N_1180,N_1657);
nor U5671 (N_5671,N_1919,N_157);
nand U5672 (N_5672,N_1132,N_919);
or U5673 (N_5673,N_2214,N_2588);
nand U5674 (N_5674,N_428,N_34);
nand U5675 (N_5675,N_115,N_2009);
or U5676 (N_5676,N_114,N_1188);
nand U5677 (N_5677,N_591,N_160);
nor U5678 (N_5678,N_1585,N_2935);
or U5679 (N_5679,N_494,N_1791);
nand U5680 (N_5680,N_1750,N_2552);
and U5681 (N_5681,N_284,N_2733);
nor U5682 (N_5682,N_2886,N_30);
nor U5683 (N_5683,N_883,N_2926);
xnor U5684 (N_5684,N_401,N_2896);
xnor U5685 (N_5685,N_1860,N_815);
or U5686 (N_5686,N_1656,N_733);
or U5687 (N_5687,N_2670,N_2507);
or U5688 (N_5688,N_1748,N_2123);
or U5689 (N_5689,N_1844,N_1920);
nor U5690 (N_5690,N_2496,N_1537);
nand U5691 (N_5691,N_2472,N_1703);
or U5692 (N_5692,N_1533,N_1343);
nor U5693 (N_5693,N_2970,N_2144);
or U5694 (N_5694,N_2065,N_343);
xor U5695 (N_5695,N_1049,N_2463);
or U5696 (N_5696,N_1786,N_2909);
and U5697 (N_5697,N_317,N_1120);
xnor U5698 (N_5698,N_1603,N_793);
and U5699 (N_5699,N_2574,N_2979);
xnor U5700 (N_5700,N_2830,N_1784);
xnor U5701 (N_5701,N_903,N_2052);
or U5702 (N_5702,N_2900,N_671);
or U5703 (N_5703,N_907,N_2151);
xnor U5704 (N_5704,N_539,N_2466);
or U5705 (N_5705,N_2444,N_404);
and U5706 (N_5706,N_2501,N_2034);
or U5707 (N_5707,N_2232,N_2839);
nor U5708 (N_5708,N_205,N_1138);
nand U5709 (N_5709,N_942,N_1809);
or U5710 (N_5710,N_146,N_1575);
nor U5711 (N_5711,N_959,N_2956);
nand U5712 (N_5712,N_1913,N_2211);
nor U5713 (N_5713,N_365,N_406);
xnor U5714 (N_5714,N_1308,N_1771);
xnor U5715 (N_5715,N_355,N_2494);
nand U5716 (N_5716,N_1078,N_1759);
nor U5717 (N_5717,N_1446,N_400);
and U5718 (N_5718,N_1139,N_830);
and U5719 (N_5719,N_1293,N_286);
nor U5720 (N_5720,N_1605,N_2569);
xor U5721 (N_5721,N_1916,N_504);
nand U5722 (N_5722,N_1537,N_2571);
xor U5723 (N_5723,N_1220,N_1968);
or U5724 (N_5724,N_1210,N_2470);
nor U5725 (N_5725,N_2021,N_318);
or U5726 (N_5726,N_803,N_1489);
or U5727 (N_5727,N_1410,N_2993);
nor U5728 (N_5728,N_2075,N_1190);
or U5729 (N_5729,N_1831,N_359);
or U5730 (N_5730,N_2467,N_574);
and U5731 (N_5731,N_160,N_2270);
nand U5732 (N_5732,N_1,N_1448);
nor U5733 (N_5733,N_2541,N_1996);
nand U5734 (N_5734,N_36,N_606);
and U5735 (N_5735,N_489,N_2322);
and U5736 (N_5736,N_2738,N_758);
or U5737 (N_5737,N_2869,N_2481);
or U5738 (N_5738,N_1111,N_1021);
nand U5739 (N_5739,N_2051,N_1682);
and U5740 (N_5740,N_1401,N_553);
nor U5741 (N_5741,N_1070,N_808);
xnor U5742 (N_5742,N_2757,N_2491);
nand U5743 (N_5743,N_2438,N_535);
and U5744 (N_5744,N_2035,N_1080);
or U5745 (N_5745,N_529,N_880);
xnor U5746 (N_5746,N_2612,N_2351);
nor U5747 (N_5747,N_1449,N_39);
or U5748 (N_5748,N_297,N_2354);
nor U5749 (N_5749,N_364,N_2639);
or U5750 (N_5750,N_2773,N_2859);
xnor U5751 (N_5751,N_806,N_1748);
and U5752 (N_5752,N_1945,N_1400);
nor U5753 (N_5753,N_1500,N_2313);
and U5754 (N_5754,N_1755,N_116);
and U5755 (N_5755,N_1518,N_669);
and U5756 (N_5756,N_1518,N_1992);
nand U5757 (N_5757,N_2127,N_126);
or U5758 (N_5758,N_1367,N_245);
xor U5759 (N_5759,N_355,N_1440);
or U5760 (N_5760,N_2112,N_1812);
and U5761 (N_5761,N_1387,N_2209);
nor U5762 (N_5762,N_572,N_1096);
and U5763 (N_5763,N_2607,N_1251);
and U5764 (N_5764,N_629,N_733);
or U5765 (N_5765,N_1961,N_2128);
xnor U5766 (N_5766,N_604,N_2307);
nand U5767 (N_5767,N_864,N_1331);
nand U5768 (N_5768,N_400,N_2300);
and U5769 (N_5769,N_83,N_1062);
nor U5770 (N_5770,N_2007,N_1148);
nor U5771 (N_5771,N_970,N_2896);
xor U5772 (N_5772,N_2594,N_80);
and U5773 (N_5773,N_2224,N_2001);
or U5774 (N_5774,N_2426,N_2938);
xor U5775 (N_5775,N_2440,N_113);
xnor U5776 (N_5776,N_768,N_1079);
and U5777 (N_5777,N_2752,N_315);
or U5778 (N_5778,N_1304,N_2568);
and U5779 (N_5779,N_139,N_2670);
nand U5780 (N_5780,N_1919,N_423);
nand U5781 (N_5781,N_2796,N_737);
or U5782 (N_5782,N_782,N_692);
and U5783 (N_5783,N_2130,N_912);
nand U5784 (N_5784,N_675,N_1026);
nor U5785 (N_5785,N_1334,N_1343);
or U5786 (N_5786,N_1722,N_1863);
nor U5787 (N_5787,N_2917,N_2525);
nand U5788 (N_5788,N_1105,N_1181);
and U5789 (N_5789,N_1999,N_1046);
and U5790 (N_5790,N_1983,N_1945);
nor U5791 (N_5791,N_2679,N_964);
xnor U5792 (N_5792,N_1797,N_311);
or U5793 (N_5793,N_160,N_1660);
xor U5794 (N_5794,N_984,N_749);
nand U5795 (N_5795,N_29,N_98);
xnor U5796 (N_5796,N_259,N_1180);
nor U5797 (N_5797,N_529,N_960);
or U5798 (N_5798,N_367,N_1489);
nand U5799 (N_5799,N_2235,N_136);
xnor U5800 (N_5800,N_722,N_364);
xor U5801 (N_5801,N_1471,N_2901);
or U5802 (N_5802,N_1473,N_2055);
xnor U5803 (N_5803,N_2284,N_698);
nor U5804 (N_5804,N_1891,N_1435);
and U5805 (N_5805,N_326,N_267);
xnor U5806 (N_5806,N_2176,N_0);
nor U5807 (N_5807,N_2411,N_2955);
nor U5808 (N_5808,N_391,N_2725);
and U5809 (N_5809,N_1375,N_81);
and U5810 (N_5810,N_1832,N_1749);
and U5811 (N_5811,N_362,N_466);
nand U5812 (N_5812,N_2623,N_898);
nand U5813 (N_5813,N_197,N_1634);
xor U5814 (N_5814,N_282,N_144);
xor U5815 (N_5815,N_95,N_1779);
xnor U5816 (N_5816,N_2130,N_88);
nand U5817 (N_5817,N_568,N_718);
xnor U5818 (N_5818,N_528,N_493);
xnor U5819 (N_5819,N_1610,N_446);
xnor U5820 (N_5820,N_1391,N_1839);
and U5821 (N_5821,N_1185,N_750);
xnor U5822 (N_5822,N_353,N_2921);
xnor U5823 (N_5823,N_2952,N_2764);
and U5824 (N_5824,N_1175,N_425);
or U5825 (N_5825,N_2818,N_1881);
nand U5826 (N_5826,N_1659,N_153);
xor U5827 (N_5827,N_2285,N_2212);
xor U5828 (N_5828,N_1786,N_704);
and U5829 (N_5829,N_494,N_332);
or U5830 (N_5830,N_1593,N_319);
nand U5831 (N_5831,N_662,N_2222);
or U5832 (N_5832,N_659,N_2563);
or U5833 (N_5833,N_1262,N_74);
or U5834 (N_5834,N_1218,N_1169);
xnor U5835 (N_5835,N_752,N_1867);
nand U5836 (N_5836,N_1209,N_981);
xor U5837 (N_5837,N_1246,N_342);
and U5838 (N_5838,N_562,N_1864);
nor U5839 (N_5839,N_1172,N_859);
nor U5840 (N_5840,N_627,N_438);
or U5841 (N_5841,N_581,N_2559);
nor U5842 (N_5842,N_2368,N_391);
and U5843 (N_5843,N_438,N_2132);
nand U5844 (N_5844,N_619,N_556);
or U5845 (N_5845,N_2176,N_151);
and U5846 (N_5846,N_673,N_1728);
xnor U5847 (N_5847,N_287,N_308);
nand U5848 (N_5848,N_792,N_1049);
xor U5849 (N_5849,N_1350,N_2509);
xnor U5850 (N_5850,N_765,N_2298);
xnor U5851 (N_5851,N_970,N_2044);
or U5852 (N_5852,N_2986,N_2280);
nor U5853 (N_5853,N_1838,N_2114);
nand U5854 (N_5854,N_2708,N_2761);
xnor U5855 (N_5855,N_1495,N_2151);
xnor U5856 (N_5856,N_2570,N_1427);
nor U5857 (N_5857,N_2963,N_963);
nand U5858 (N_5858,N_145,N_364);
or U5859 (N_5859,N_1064,N_1618);
xnor U5860 (N_5860,N_945,N_2853);
nor U5861 (N_5861,N_1216,N_350);
and U5862 (N_5862,N_926,N_1902);
or U5863 (N_5863,N_1987,N_2746);
and U5864 (N_5864,N_1628,N_2974);
and U5865 (N_5865,N_722,N_519);
and U5866 (N_5866,N_1761,N_9);
xnor U5867 (N_5867,N_1973,N_2531);
nor U5868 (N_5868,N_665,N_1810);
nor U5869 (N_5869,N_2287,N_366);
or U5870 (N_5870,N_2622,N_2917);
xnor U5871 (N_5871,N_829,N_264);
xnor U5872 (N_5872,N_69,N_2979);
or U5873 (N_5873,N_752,N_1830);
nand U5874 (N_5874,N_2755,N_1580);
or U5875 (N_5875,N_2816,N_1978);
nand U5876 (N_5876,N_338,N_2350);
nand U5877 (N_5877,N_2182,N_2249);
and U5878 (N_5878,N_1423,N_742);
or U5879 (N_5879,N_1704,N_1127);
and U5880 (N_5880,N_939,N_2281);
xor U5881 (N_5881,N_523,N_2810);
or U5882 (N_5882,N_729,N_188);
and U5883 (N_5883,N_1337,N_938);
or U5884 (N_5884,N_2247,N_1141);
nand U5885 (N_5885,N_350,N_534);
nor U5886 (N_5886,N_2918,N_2201);
nor U5887 (N_5887,N_1649,N_2218);
nor U5888 (N_5888,N_2054,N_2851);
nor U5889 (N_5889,N_1206,N_2205);
xnor U5890 (N_5890,N_125,N_778);
xor U5891 (N_5891,N_658,N_700);
and U5892 (N_5892,N_1064,N_1648);
or U5893 (N_5893,N_2212,N_2006);
xnor U5894 (N_5894,N_1080,N_2506);
xor U5895 (N_5895,N_2592,N_2567);
nor U5896 (N_5896,N_349,N_2429);
or U5897 (N_5897,N_1320,N_1418);
nor U5898 (N_5898,N_85,N_1542);
xor U5899 (N_5899,N_287,N_2639);
or U5900 (N_5900,N_1775,N_564);
nand U5901 (N_5901,N_726,N_624);
and U5902 (N_5902,N_2153,N_1889);
xnor U5903 (N_5903,N_2702,N_1096);
or U5904 (N_5904,N_2671,N_2513);
and U5905 (N_5905,N_1694,N_1718);
or U5906 (N_5906,N_2267,N_1810);
nand U5907 (N_5907,N_2315,N_101);
nor U5908 (N_5908,N_334,N_2524);
nand U5909 (N_5909,N_197,N_1812);
nand U5910 (N_5910,N_2255,N_2416);
xor U5911 (N_5911,N_809,N_2968);
or U5912 (N_5912,N_696,N_2921);
xor U5913 (N_5913,N_339,N_423);
nand U5914 (N_5914,N_155,N_2668);
nor U5915 (N_5915,N_460,N_1329);
xor U5916 (N_5916,N_1459,N_518);
xnor U5917 (N_5917,N_2191,N_381);
and U5918 (N_5918,N_359,N_34);
nor U5919 (N_5919,N_1559,N_259);
or U5920 (N_5920,N_1983,N_2162);
nor U5921 (N_5921,N_2014,N_2704);
xnor U5922 (N_5922,N_1898,N_1200);
xnor U5923 (N_5923,N_1174,N_747);
nand U5924 (N_5924,N_455,N_2983);
nor U5925 (N_5925,N_2368,N_1606);
nor U5926 (N_5926,N_1430,N_2131);
xor U5927 (N_5927,N_2013,N_469);
and U5928 (N_5928,N_1430,N_897);
nand U5929 (N_5929,N_2272,N_2710);
or U5930 (N_5930,N_2503,N_1895);
nor U5931 (N_5931,N_1964,N_1739);
nand U5932 (N_5932,N_2243,N_395);
and U5933 (N_5933,N_377,N_1977);
nor U5934 (N_5934,N_2349,N_1977);
nand U5935 (N_5935,N_2011,N_1507);
or U5936 (N_5936,N_1994,N_227);
and U5937 (N_5937,N_14,N_1054);
and U5938 (N_5938,N_1720,N_1065);
nor U5939 (N_5939,N_196,N_257);
xnor U5940 (N_5940,N_1658,N_827);
nand U5941 (N_5941,N_1608,N_181);
and U5942 (N_5942,N_365,N_2943);
and U5943 (N_5943,N_1348,N_701);
nand U5944 (N_5944,N_1958,N_2702);
or U5945 (N_5945,N_1134,N_2175);
nor U5946 (N_5946,N_1367,N_2128);
nor U5947 (N_5947,N_2523,N_373);
xor U5948 (N_5948,N_1021,N_2829);
or U5949 (N_5949,N_2247,N_211);
nor U5950 (N_5950,N_2802,N_653);
xnor U5951 (N_5951,N_1846,N_2148);
and U5952 (N_5952,N_2779,N_2745);
nand U5953 (N_5953,N_2045,N_1358);
nand U5954 (N_5954,N_1615,N_1314);
nor U5955 (N_5955,N_764,N_1932);
and U5956 (N_5956,N_1855,N_1882);
nand U5957 (N_5957,N_1554,N_1079);
nor U5958 (N_5958,N_2103,N_1098);
nor U5959 (N_5959,N_846,N_1884);
xnor U5960 (N_5960,N_881,N_2265);
xor U5961 (N_5961,N_2457,N_2934);
nand U5962 (N_5962,N_421,N_2383);
xnor U5963 (N_5963,N_2689,N_2176);
and U5964 (N_5964,N_1394,N_2586);
or U5965 (N_5965,N_1306,N_153);
xor U5966 (N_5966,N_2670,N_1707);
and U5967 (N_5967,N_2328,N_1425);
xor U5968 (N_5968,N_626,N_2358);
and U5969 (N_5969,N_659,N_826);
or U5970 (N_5970,N_2081,N_261);
nor U5971 (N_5971,N_2087,N_2667);
xnor U5972 (N_5972,N_1218,N_744);
nor U5973 (N_5973,N_883,N_427);
xnor U5974 (N_5974,N_2624,N_2130);
nor U5975 (N_5975,N_2451,N_795);
nand U5976 (N_5976,N_834,N_121);
or U5977 (N_5977,N_227,N_1085);
or U5978 (N_5978,N_2555,N_2047);
and U5979 (N_5979,N_2299,N_1033);
and U5980 (N_5980,N_1527,N_2784);
and U5981 (N_5981,N_2594,N_2642);
and U5982 (N_5982,N_1992,N_456);
xnor U5983 (N_5983,N_2858,N_1585);
xnor U5984 (N_5984,N_10,N_571);
and U5985 (N_5985,N_1653,N_660);
or U5986 (N_5986,N_177,N_11);
and U5987 (N_5987,N_1078,N_1967);
and U5988 (N_5988,N_70,N_1240);
xnor U5989 (N_5989,N_2866,N_2794);
nor U5990 (N_5990,N_24,N_2985);
or U5991 (N_5991,N_2189,N_2733);
nor U5992 (N_5992,N_699,N_1843);
and U5993 (N_5993,N_1784,N_199);
nand U5994 (N_5994,N_2956,N_1636);
nor U5995 (N_5995,N_2998,N_1917);
nand U5996 (N_5996,N_598,N_1811);
nor U5997 (N_5997,N_894,N_1101);
xor U5998 (N_5998,N_1566,N_2500);
xor U5999 (N_5999,N_2054,N_589);
and U6000 (N_6000,N_3174,N_4347);
nand U6001 (N_6001,N_4993,N_4974);
and U6002 (N_6002,N_4073,N_5914);
nor U6003 (N_6003,N_3220,N_5430);
or U6004 (N_6004,N_4415,N_5217);
or U6005 (N_6005,N_4524,N_5770);
xnor U6006 (N_6006,N_4820,N_4301);
nand U6007 (N_6007,N_3270,N_5036);
and U6008 (N_6008,N_4568,N_5684);
nand U6009 (N_6009,N_3005,N_5298);
or U6010 (N_6010,N_3304,N_5370);
or U6011 (N_6011,N_5310,N_5131);
nand U6012 (N_6012,N_3349,N_3172);
or U6013 (N_6013,N_3689,N_3440);
and U6014 (N_6014,N_3140,N_4865);
or U6015 (N_6015,N_5241,N_3061);
nor U6016 (N_6016,N_4324,N_3554);
or U6017 (N_6017,N_3859,N_5208);
or U6018 (N_6018,N_4293,N_5820);
nand U6019 (N_6019,N_5561,N_5919);
and U6020 (N_6020,N_5396,N_4922);
xnor U6021 (N_6021,N_4026,N_3238);
xor U6022 (N_6022,N_3804,N_5194);
xor U6023 (N_6023,N_3371,N_5883);
nand U6024 (N_6024,N_4245,N_4903);
or U6025 (N_6025,N_3396,N_3613);
nand U6026 (N_6026,N_4286,N_5360);
and U6027 (N_6027,N_3053,N_5921);
or U6028 (N_6028,N_5052,N_4751);
and U6029 (N_6029,N_4621,N_4655);
and U6030 (N_6030,N_4425,N_3322);
nor U6031 (N_6031,N_4667,N_3260);
and U6032 (N_6032,N_4696,N_4926);
and U6033 (N_6033,N_3427,N_3160);
or U6034 (N_6034,N_3205,N_4866);
xor U6035 (N_6035,N_3827,N_3048);
and U6036 (N_6036,N_5617,N_3555);
and U6037 (N_6037,N_3101,N_5595);
and U6038 (N_6038,N_5281,N_3411);
and U6039 (N_6039,N_5659,N_4398);
xor U6040 (N_6040,N_5057,N_5511);
nand U6041 (N_6041,N_3051,N_5748);
or U6042 (N_6042,N_4101,N_3120);
and U6043 (N_6043,N_3444,N_3478);
or U6044 (N_6044,N_4914,N_3650);
and U6045 (N_6045,N_4904,N_4342);
or U6046 (N_6046,N_5510,N_3452);
nor U6047 (N_6047,N_4143,N_3082);
nand U6048 (N_6048,N_4118,N_4290);
nand U6049 (N_6049,N_4658,N_4016);
nand U6050 (N_6050,N_4268,N_3907);
xnor U6051 (N_6051,N_4647,N_4089);
nor U6052 (N_6052,N_5264,N_4367);
xnor U6053 (N_6053,N_5005,N_5892);
xor U6054 (N_6054,N_5946,N_4446);
and U6055 (N_6055,N_4729,N_4876);
nand U6056 (N_6056,N_3321,N_5765);
nand U6057 (N_6057,N_4085,N_4172);
nor U6058 (N_6058,N_3248,N_5314);
nand U6059 (N_6059,N_4808,N_4202);
nand U6060 (N_6060,N_3562,N_4784);
nor U6061 (N_6061,N_4777,N_3295);
xor U6062 (N_6062,N_4705,N_4780);
and U6063 (N_6063,N_5466,N_3951);
nand U6064 (N_6064,N_3932,N_3878);
nor U6065 (N_6065,N_5101,N_5709);
xnor U6066 (N_6066,N_3041,N_4084);
nor U6067 (N_6067,N_4478,N_5687);
and U6068 (N_6068,N_5816,N_4765);
nand U6069 (N_6069,N_5917,N_4279);
or U6070 (N_6070,N_5995,N_5837);
xor U6071 (N_6071,N_5810,N_5184);
xor U6072 (N_6072,N_3818,N_3251);
and U6073 (N_6073,N_5918,N_4919);
nand U6074 (N_6074,N_5358,N_4976);
nor U6075 (N_6075,N_5368,N_5296);
nand U6076 (N_6076,N_3151,N_5961);
or U6077 (N_6077,N_5300,N_4468);
xor U6078 (N_6078,N_4594,N_4657);
nor U6079 (N_6079,N_5244,N_3007);
xor U6080 (N_6080,N_3741,N_5996);
and U6081 (N_6081,N_5708,N_4372);
nand U6082 (N_6082,N_4029,N_5222);
xor U6083 (N_6083,N_4044,N_4300);
or U6084 (N_6084,N_3156,N_3568);
and U6085 (N_6085,N_4994,N_5204);
nand U6086 (N_6086,N_4136,N_4381);
xnor U6087 (N_6087,N_5098,N_4989);
xnor U6088 (N_6088,N_4275,N_5138);
nor U6089 (N_6089,N_3313,N_3374);
nand U6090 (N_6090,N_3791,N_5092);
xnor U6091 (N_6091,N_3638,N_5929);
or U6092 (N_6092,N_5809,N_5291);
nand U6093 (N_6093,N_3730,N_5255);
xnor U6094 (N_6094,N_4664,N_5063);
and U6095 (N_6095,N_4206,N_5814);
and U6096 (N_6096,N_3345,N_4127);
and U6097 (N_6097,N_5160,N_5355);
or U6098 (N_6098,N_5972,N_3953);
or U6099 (N_6099,N_4819,N_3290);
xnor U6100 (N_6100,N_5514,N_5307);
nor U6101 (N_6101,N_4411,N_5849);
or U6102 (N_6102,N_3422,N_4007);
or U6103 (N_6103,N_3144,N_5970);
nand U6104 (N_6104,N_5539,N_3527);
nor U6105 (N_6105,N_4811,N_5905);
and U6106 (N_6106,N_4687,N_5379);
nor U6107 (N_6107,N_5349,N_4023);
and U6108 (N_6108,N_3912,N_4449);
and U6109 (N_6109,N_3428,N_3375);
nor U6110 (N_6110,N_5115,N_4821);
or U6111 (N_6111,N_3446,N_4863);
and U6112 (N_6112,N_5382,N_5186);
or U6113 (N_6113,N_4852,N_5832);
nand U6114 (N_6114,N_3213,N_3426);
nor U6115 (N_6115,N_5532,N_4831);
or U6116 (N_6116,N_3919,N_4075);
nor U6117 (N_6117,N_4875,N_5018);
nand U6118 (N_6118,N_3563,N_4115);
nor U6119 (N_6119,N_5344,N_3343);
nor U6120 (N_6120,N_5326,N_3712);
nor U6121 (N_6121,N_4389,N_4661);
or U6122 (N_6122,N_3024,N_4295);
xor U6123 (N_6123,N_5676,N_4582);
and U6124 (N_6124,N_5259,N_3692);
xor U6125 (N_6125,N_3910,N_4538);
nand U6126 (N_6126,N_4548,N_4169);
nor U6127 (N_6127,N_5537,N_5183);
nor U6128 (N_6128,N_5383,N_3696);
or U6129 (N_6129,N_3887,N_3548);
nand U6130 (N_6130,N_4596,N_3207);
or U6131 (N_6131,N_4608,N_4618);
or U6132 (N_6132,N_4428,N_4317);
nand U6133 (N_6133,N_3350,N_3999);
nor U6134 (N_6134,N_5085,N_4839);
and U6135 (N_6135,N_4900,N_3690);
nor U6136 (N_6136,N_3166,N_5262);
and U6137 (N_6137,N_5414,N_3641);
xnor U6138 (N_6138,N_5710,N_3064);
xor U6139 (N_6139,N_5844,N_3462);
and U6140 (N_6140,N_4972,N_4378);
or U6141 (N_6141,N_4199,N_3871);
and U6142 (N_6142,N_3489,N_3386);
nor U6143 (N_6143,N_5263,N_3844);
or U6144 (N_6144,N_4196,N_4540);
nor U6145 (N_6145,N_5666,N_5951);
nand U6146 (N_6146,N_4114,N_3116);
or U6147 (N_6147,N_4802,N_5873);
and U6148 (N_6148,N_5726,N_5641);
xor U6149 (N_6149,N_4028,N_3333);
nor U6150 (N_6150,N_4727,N_3433);
xor U6151 (N_6151,N_5622,N_4410);
nand U6152 (N_6152,N_4401,N_3264);
nor U6153 (N_6153,N_5534,N_5243);
nor U6154 (N_6154,N_5673,N_5866);
xor U6155 (N_6155,N_5412,N_5863);
and U6156 (N_6156,N_4605,N_5031);
nand U6157 (N_6157,N_3508,N_3453);
and U6158 (N_6158,N_4208,N_3931);
xor U6159 (N_6159,N_4453,N_5000);
and U6160 (N_6160,N_4774,N_3947);
and U6161 (N_6161,N_5491,N_4187);
or U6162 (N_6162,N_3403,N_4690);
nand U6163 (N_6163,N_5274,N_5670);
nor U6164 (N_6164,N_3731,N_5689);
and U6165 (N_6165,N_4219,N_5719);
or U6166 (N_6166,N_3753,N_4640);
nand U6167 (N_6167,N_5768,N_4178);
nand U6168 (N_6168,N_5394,N_3896);
nand U6169 (N_6169,N_5955,N_3188);
xor U6170 (N_6170,N_4339,N_5916);
and U6171 (N_6171,N_4315,N_4986);
or U6172 (N_6172,N_5322,N_5724);
xor U6173 (N_6173,N_5904,N_4527);
nand U6174 (N_6174,N_5247,N_4792);
and U6175 (N_6175,N_3732,N_5419);
nand U6176 (N_6176,N_4750,N_5044);
or U6177 (N_6177,N_4234,N_5427);
nand U6178 (N_6178,N_4135,N_4346);
or U6179 (N_6179,N_5251,N_3477);
and U6180 (N_6180,N_4319,N_4726);
or U6181 (N_6181,N_3836,N_5949);
nand U6182 (N_6182,N_3379,N_5745);
or U6183 (N_6183,N_4982,N_4981);
or U6184 (N_6184,N_3627,N_4395);
nor U6185 (N_6185,N_3894,N_3222);
nand U6186 (N_6186,N_4805,N_4668);
and U6187 (N_6187,N_3869,N_5070);
or U6188 (N_6188,N_3498,N_3214);
nor U6189 (N_6189,N_3451,N_5010);
xor U6190 (N_6190,N_4785,N_5354);
nand U6191 (N_6191,N_5371,N_3749);
or U6192 (N_6192,N_5406,N_5680);
nand U6193 (N_6193,N_5216,N_4559);
nand U6194 (N_6194,N_5749,N_4710);
nand U6195 (N_6195,N_5701,N_5476);
and U6196 (N_6196,N_5341,N_5829);
xor U6197 (N_6197,N_4261,N_4890);
or U6198 (N_6198,N_4649,N_5359);
nand U6199 (N_6199,N_5718,N_4050);
or U6200 (N_6200,N_5176,N_4814);
or U6201 (N_6201,N_5214,N_5668);
xor U6202 (N_6202,N_5535,N_5425);
or U6203 (N_6203,N_4100,N_5267);
and U6204 (N_6204,N_3317,N_5619);
nand U6205 (N_6205,N_4120,N_3868);
xor U6206 (N_6206,N_4355,N_3078);
and U6207 (N_6207,N_4297,N_4375);
nand U6208 (N_6208,N_3042,N_5597);
xnor U6209 (N_6209,N_5975,N_3835);
or U6210 (N_6210,N_5640,N_5774);
nor U6211 (N_6211,N_4112,N_3806);
and U6212 (N_6212,N_4498,N_5757);
nor U6213 (N_6213,N_4393,N_5694);
or U6214 (N_6214,N_3590,N_5367);
and U6215 (N_6215,N_5474,N_5058);
nand U6216 (N_6216,N_5332,N_4654);
nand U6217 (N_6217,N_3037,N_5885);
nor U6218 (N_6218,N_4590,N_3625);
or U6219 (N_6219,N_3980,N_5831);
and U6220 (N_6220,N_4862,N_4723);
nand U6221 (N_6221,N_3305,N_5090);
and U6222 (N_6222,N_5562,N_5703);
xnor U6223 (N_6223,N_5522,N_5422);
xnor U6224 (N_6224,N_5236,N_5315);
nor U6225 (N_6225,N_5911,N_5203);
xnor U6226 (N_6226,N_4359,N_3927);
or U6227 (N_6227,N_4666,N_5894);
nand U6228 (N_6228,N_3470,N_3083);
nand U6229 (N_6229,N_3173,N_3786);
and U6230 (N_6230,N_5893,N_5880);
and U6231 (N_6231,N_3978,N_4604);
or U6232 (N_6232,N_4364,N_3697);
and U6233 (N_6233,N_3162,N_3103);
nand U6234 (N_6234,N_4117,N_5155);
or U6235 (N_6235,N_4479,N_3917);
and U6236 (N_6236,N_4844,N_3329);
and U6237 (N_6237,N_5448,N_4015);
nand U6238 (N_6238,N_5954,N_4846);
nand U6239 (N_6239,N_5449,N_3062);
or U6240 (N_6240,N_4243,N_3545);
xor U6241 (N_6241,N_3181,N_4368);
nand U6242 (N_6242,N_4108,N_4283);
nor U6243 (N_6243,N_3584,N_4333);
and U6244 (N_6244,N_4140,N_4996);
nand U6245 (N_6245,N_4060,N_3959);
xnor U6246 (N_6246,N_3010,N_3955);
xor U6247 (N_6247,N_5128,N_5960);
nor U6248 (N_6248,N_3232,N_3038);
nor U6249 (N_6249,N_4139,N_5346);
and U6250 (N_6250,N_5769,N_4851);
or U6251 (N_6251,N_4492,N_5845);
and U6252 (N_6252,N_4675,N_3977);
and U6253 (N_6253,N_3595,N_5363);
nand U6254 (N_6254,N_4741,N_4350);
xor U6255 (N_6255,N_3898,N_5118);
nor U6256 (N_6256,N_3035,N_3788);
nor U6257 (N_6257,N_4277,N_4848);
or U6258 (N_6258,N_4326,N_4464);
or U6259 (N_6259,N_3157,N_3210);
nor U6260 (N_6260,N_3825,N_3909);
and U6261 (N_6261,N_4435,N_5096);
xor U6262 (N_6262,N_3292,N_3594);
nor U6263 (N_6263,N_4032,N_3273);
nand U6264 (N_6264,N_5876,N_4874);
xor U6265 (N_6265,N_5145,N_5408);
or U6266 (N_6266,N_3876,N_5311);
and U6267 (N_6267,N_5032,N_3920);
or U6268 (N_6268,N_3642,N_4629);
xor U6269 (N_6269,N_3380,N_5189);
nand U6270 (N_6270,N_5702,N_5191);
nor U6271 (N_6271,N_3285,N_4505);
xnor U6272 (N_6272,N_5907,N_3124);
and U6273 (N_6273,N_5665,N_5607);
and U6274 (N_6274,N_3149,N_4081);
or U6275 (N_6275,N_3893,N_3676);
nor U6276 (N_6276,N_5693,N_3347);
nand U6277 (N_6277,N_5125,N_4676);
and U6278 (N_6278,N_5662,N_4466);
nor U6279 (N_6279,N_5426,N_3670);
and U6280 (N_6280,N_4545,N_5223);
xnor U6281 (N_6281,N_5402,N_4915);
nor U6282 (N_6282,N_4531,N_4790);
nor U6283 (N_6283,N_4309,N_4220);
and U6284 (N_6284,N_3579,N_4603);
nand U6285 (N_6285,N_4623,N_5543);
nand U6286 (N_6286,N_4991,N_3407);
nand U6287 (N_6287,N_5669,N_3722);
nand U6288 (N_6288,N_5750,N_4635);
and U6289 (N_6289,N_4701,N_3972);
nor U6290 (N_6290,N_5813,N_4461);
nor U6291 (N_6291,N_4336,N_4971);
nor U6292 (N_6292,N_3376,N_3808);
xnor U6293 (N_6293,N_3123,N_4241);
or U6294 (N_6294,N_3571,N_5477);
and U6295 (N_6295,N_3762,N_4209);
or U6296 (N_6296,N_4533,N_5283);
nand U6297 (N_6297,N_5171,N_5054);
or U6298 (N_6298,N_3537,N_3298);
nand U6299 (N_6299,N_3725,N_5868);
or U6300 (N_6300,N_3984,N_5004);
xor U6301 (N_6301,N_4049,N_5481);
and U6302 (N_6302,N_5802,N_5871);
xnor U6303 (N_6303,N_3943,N_3688);
and U6304 (N_6304,N_5029,N_4168);
xnor U6305 (N_6305,N_4402,N_5112);
nor U6306 (N_6306,N_4685,N_4223);
nor U6307 (N_6307,N_3939,N_4602);
or U6308 (N_6308,N_3644,N_4636);
xnor U6309 (N_6309,N_4950,N_5901);
and U6310 (N_6310,N_4110,N_5050);
or U6311 (N_6311,N_3723,N_4953);
xnor U6312 (N_6312,N_4632,N_3565);
or U6313 (N_6313,N_3837,N_5533);
xor U6314 (N_6314,N_3367,N_4769);
nor U6315 (N_6315,N_5772,N_3889);
nand U6316 (N_6316,N_4263,N_3040);
or U6317 (N_6317,N_3814,N_3208);
xnor U6318 (N_6318,N_3332,N_3283);
and U6319 (N_6319,N_3095,N_5446);
nand U6320 (N_6320,N_4376,N_3683);
xor U6321 (N_6321,N_4537,N_3559);
or U6322 (N_6322,N_5898,N_3022);
nor U6323 (N_6323,N_4789,N_5407);
nor U6324 (N_6324,N_4691,N_3501);
and U6325 (N_6325,N_5526,N_4008);
or U6326 (N_6326,N_3311,N_5019);
nor U6327 (N_6327,N_3771,N_5698);
xnor U6328 (N_6328,N_4191,N_3388);
and U6329 (N_6329,N_4362,N_4961);
xor U6330 (N_6330,N_5172,N_5423);
and U6331 (N_6331,N_3268,N_3202);
or U6332 (N_6332,N_5922,N_4672);
nand U6333 (N_6333,N_3507,N_3539);
or U6334 (N_6334,N_5177,N_5691);
and U6335 (N_6335,N_4124,N_4956);
nand U6336 (N_6336,N_4762,N_3085);
nor U6337 (N_6337,N_3246,N_4121);
nand U6338 (N_6338,N_3057,N_5158);
nor U6339 (N_6339,N_5834,N_3556);
nor U6340 (N_6340,N_4680,N_5139);
nor U6341 (N_6341,N_3335,N_3073);
or U6342 (N_6342,N_3713,N_4233);
or U6343 (N_6343,N_4157,N_5720);
and U6344 (N_6344,N_4891,N_3118);
and U6345 (N_6345,N_4166,N_3602);
nor U6346 (N_6346,N_3715,N_5799);
or U6347 (N_6347,N_5879,N_4975);
or U6348 (N_6348,N_5023,N_5178);
nor U6349 (N_6349,N_3765,N_3533);
xnor U6350 (N_6350,N_5489,N_4700);
nor U6351 (N_6351,N_5478,N_3829);
nor U6352 (N_6352,N_3253,N_3293);
and U6353 (N_6353,N_3986,N_3634);
nand U6354 (N_6354,N_3574,N_4096);
or U6355 (N_6355,N_3025,N_3785);
nand U6356 (N_6356,N_4589,N_3243);
xnor U6357 (N_6357,N_5571,N_5727);
nor U6358 (N_6358,N_5209,N_4467);
xor U6359 (N_6359,N_3740,N_3846);
nor U6360 (N_6360,N_3551,N_3011);
or U6361 (N_6361,N_3099,N_4962);
nor U6362 (N_6362,N_5912,N_5103);
nor U6363 (N_6363,N_4583,N_4005);
and U6364 (N_6364,N_4645,N_4144);
nand U6365 (N_6365,N_5605,N_5121);
nand U6366 (N_6366,N_3708,N_4817);
nor U6367 (N_6367,N_4896,N_5159);
or U6368 (N_6368,N_5626,N_4386);
nor U6369 (N_6369,N_4718,N_4195);
and U6370 (N_6370,N_3774,N_4493);
or U6371 (N_6371,N_4334,N_5685);
nor U6372 (N_6372,N_5974,N_3935);
nand U6373 (N_6373,N_5592,N_4642);
or U6374 (N_6374,N_4593,N_3342);
nor U6375 (N_6375,N_5723,N_3815);
or U6376 (N_6376,N_4773,N_5705);
or U6377 (N_6377,N_5494,N_3589);
nand U6378 (N_6378,N_3975,N_3463);
nand U6379 (N_6379,N_3661,N_3534);
nor U6380 (N_6380,N_4039,N_4057);
or U6381 (N_6381,N_4422,N_4019);
nor U6382 (N_6382,N_4850,N_5903);
xnor U6383 (N_6383,N_4958,N_5574);
and U6384 (N_6384,N_4794,N_4371);
or U6385 (N_6385,N_4237,N_3849);
or U6386 (N_6386,N_3145,N_4899);
xor U6387 (N_6387,N_5324,N_5087);
or U6388 (N_6388,N_4743,N_4541);
and U6389 (N_6389,N_3354,N_3664);
xor U6390 (N_6390,N_3398,N_5590);
nor U6391 (N_6391,N_5039,N_4697);
and U6392 (N_6392,N_4514,N_4704);
and U6393 (N_6393,N_4998,N_5431);
and U6394 (N_6394,N_4104,N_3677);
nand U6395 (N_6395,N_3237,N_3831);
nor U6396 (N_6396,N_3699,N_3484);
and U6397 (N_6397,N_4943,N_3421);
and U6398 (N_6398,N_3126,N_4829);
nor U6399 (N_6399,N_3934,N_5345);
nand U6400 (N_6400,N_5753,N_4949);
nor U6401 (N_6401,N_5199,N_3230);
and U6402 (N_6402,N_3737,N_3900);
or U6403 (N_6403,N_5973,N_3231);
xnor U6404 (N_6404,N_4679,N_5920);
or U6405 (N_6405,N_4179,N_3834);
or U6406 (N_6406,N_5471,N_3466);
xor U6407 (N_6407,N_3619,N_4278);
nand U6408 (N_6408,N_4225,N_5195);
and U6409 (N_6409,N_3526,N_3944);
nand U6410 (N_6410,N_5456,N_3903);
nor U6411 (N_6411,N_4526,N_5940);
and U6412 (N_6412,N_5787,N_3643);
and U6413 (N_6413,N_3266,N_3987);
and U6414 (N_6414,N_3582,N_3503);
nand U6415 (N_6415,N_4487,N_3397);
nor U6416 (N_6416,N_5167,N_5529);
xnor U6417 (N_6417,N_3921,N_5240);
xor U6418 (N_6418,N_3183,N_3826);
and U6419 (N_6419,N_5289,N_3916);
or U6420 (N_6420,N_3993,N_4292);
nor U6421 (N_6421,N_4353,N_3573);
xnor U6422 (N_6422,N_3113,N_3610);
nand U6423 (N_6423,N_3023,N_3154);
nor U6424 (N_6424,N_3132,N_5763);
nand U6425 (N_6425,N_5157,N_4149);
and U6426 (N_6426,N_4391,N_5323);
xor U6427 (N_6427,N_5984,N_5721);
and U6428 (N_6428,N_4581,N_5869);
xnor U6429 (N_6429,N_3707,N_4033);
or U6430 (N_6430,N_3393,N_3585);
xor U6431 (N_6431,N_4451,N_3756);
nor U6432 (N_6432,N_4055,N_4271);
or U6433 (N_6433,N_5601,N_3392);
xor U6434 (N_6434,N_4929,N_4427);
or U6435 (N_6435,N_4959,N_4358);
xor U6436 (N_6436,N_5677,N_4069);
nand U6437 (N_6437,N_3450,N_3262);
and U6438 (N_6438,N_3069,N_4426);
nor U6439 (N_6439,N_5499,N_3164);
nor U6440 (N_6440,N_4474,N_4830);
xnor U6441 (N_6441,N_3307,N_5821);
nand U6442 (N_6442,N_5127,N_5957);
nand U6443 (N_6443,N_5303,N_5452);
or U6444 (N_6444,N_4652,N_4923);
nor U6445 (N_6445,N_3254,N_4551);
xnor U6446 (N_6446,N_5470,N_4739);
and U6447 (N_6447,N_5674,N_5416);
and U6448 (N_6448,N_4898,N_5563);
xnor U6449 (N_6449,N_5890,N_4614);
or U6450 (N_6450,N_5950,N_3226);
xor U6451 (N_6451,N_4062,N_3192);
xor U6452 (N_6452,N_4942,N_3983);
and U6453 (N_6453,N_4713,N_4554);
and U6454 (N_6454,N_3217,N_3245);
or U6455 (N_6455,N_3119,N_3234);
or U6456 (N_6456,N_5305,N_4258);
or U6457 (N_6457,N_3044,N_4622);
nor U6458 (N_6458,N_3077,N_3971);
nor U6459 (N_6459,N_5982,N_3564);
xnor U6460 (N_6460,N_3654,N_4071);
nor U6461 (N_6461,N_3607,N_4163);
and U6462 (N_6462,N_3056,N_5288);
and U6463 (N_6463,N_4014,N_5738);
and U6464 (N_6464,N_4494,N_5862);
xnor U6465 (N_6465,N_4103,N_3855);
or U6466 (N_6466,N_5608,N_5699);
or U6467 (N_6467,N_5553,N_4306);
and U6468 (N_6468,N_4226,N_4842);
and U6469 (N_6469,N_4077,N_4086);
xor U6470 (N_6470,N_3286,N_3402);
xnor U6471 (N_6471,N_5006,N_3122);
nand U6472 (N_6472,N_3914,N_3684);
nor U6473 (N_6473,N_4348,N_3714);
nand U6474 (N_6474,N_3369,N_5190);
and U6475 (N_6475,N_3851,N_3008);
nor U6476 (N_6476,N_3760,N_3500);
xor U6477 (N_6477,N_4951,N_5867);
nand U6478 (N_6478,N_4930,N_4323);
nor U6479 (N_6479,N_4369,N_5811);
xor U6480 (N_6480,N_4617,N_5325);
xnor U6481 (N_6481,N_3055,N_4325);
nand U6482 (N_6482,N_4484,N_5953);
nand U6483 (N_6483,N_4260,N_5554);
nor U6484 (N_6484,N_5261,N_5164);
and U6485 (N_6485,N_3686,N_3097);
nor U6486 (N_6486,N_3705,N_5501);
or U6487 (N_6487,N_4512,N_4677);
xor U6488 (N_6488,N_5304,N_5623);
or U6489 (N_6489,N_5882,N_5061);
or U6490 (N_6490,N_3609,N_5111);
and U6491 (N_6491,N_5077,N_4519);
xnor U6492 (N_6492,N_3631,N_4877);
nand U6493 (N_6493,N_4611,N_5317);
and U6494 (N_6494,N_3612,N_3356);
nor U6495 (N_6495,N_3263,N_4291);
or U6496 (N_6496,N_4417,N_3088);
nor U6497 (N_6497,N_5339,N_3365);
nand U6498 (N_6498,N_5716,N_3219);
nand U6499 (N_6499,N_3561,N_4782);
nand U6500 (N_6500,N_5518,N_4760);
nand U6501 (N_6501,N_3576,N_3995);
and U6502 (N_6502,N_5338,N_3938);
xnor U6503 (N_6503,N_3351,N_3456);
and U6504 (N_6504,N_3769,N_3480);
nand U6505 (N_6505,N_4285,N_5736);
or U6506 (N_6506,N_5507,N_5095);
and U6507 (N_6507,N_5279,N_4074);
or U6508 (N_6508,N_3599,N_3068);
or U6509 (N_6509,N_5462,N_5512);
xnor U6510 (N_6510,N_4404,N_3139);
or U6511 (N_6511,N_5104,N_5743);
and U6512 (N_6512,N_5761,N_5651);
or U6513 (N_6513,N_5784,N_5132);
or U6514 (N_6514,N_4201,N_5170);
xnor U6515 (N_6515,N_4310,N_5088);
xnor U6516 (N_6516,N_4129,N_5333);
and U6517 (N_6517,N_5365,N_3530);
or U6518 (N_6518,N_3792,N_5116);
xor U6519 (N_6519,N_3577,N_3021);
or U6520 (N_6520,N_4341,N_3430);
nand U6521 (N_6521,N_5780,N_4634);
nand U6522 (N_6522,N_3221,N_3710);
xor U6523 (N_6523,N_3373,N_5520);
nor U6524 (N_6524,N_4812,N_4088);
xor U6525 (N_6525,N_3086,N_4637);
xnor U6526 (N_6526,N_3974,N_4833);
nor U6527 (N_6527,N_5642,N_3867);
and U6528 (N_6528,N_3761,N_5963);
nor U6529 (N_6529,N_5292,N_5071);
or U6530 (N_6530,N_5286,N_4270);
or U6531 (N_6531,N_4354,N_3355);
or U6532 (N_6532,N_3464,N_4884);
and U6533 (N_6533,N_4518,N_5927);
or U6534 (N_6534,N_4099,N_4732);
or U6535 (N_6535,N_3515,N_3108);
and U6536 (N_6536,N_4340,N_3875);
nor U6537 (N_6537,N_3143,N_4043);
nor U6538 (N_6538,N_4119,N_5487);
or U6539 (N_6539,N_4630,N_5516);
xor U6540 (N_6540,N_4337,N_4544);
nor U6541 (N_6541,N_4836,N_3146);
xnor U6542 (N_6542,N_5447,N_5541);
or U6543 (N_6543,N_3678,N_4162);
and U6544 (N_6544,N_4365,N_4298);
xnor U6545 (N_6545,N_3617,N_4414);
nor U6546 (N_6546,N_5219,N_5313);
or U6547 (N_6547,N_3493,N_5925);
and U6548 (N_6548,N_5483,N_4528);
and U6549 (N_6549,N_5731,N_4217);
nand U6550 (N_6550,N_5372,N_4565);
xor U6551 (N_6551,N_3338,N_4186);
or U6552 (N_6552,N_4746,N_4387);
and U6553 (N_6553,N_4221,N_4892);
nor U6554 (N_6554,N_5337,N_5188);
xnor U6555 (N_6555,N_4154,N_3637);
and U6556 (N_6556,N_3755,N_4431);
nor U6557 (N_6557,N_3158,N_5334);
and U6558 (N_6558,N_4535,N_5897);
nor U6559 (N_6559,N_3925,N_5454);
and U6560 (N_6560,N_3820,N_4717);
nor U6561 (N_6561,N_4207,N_3523);
nor U6562 (N_6562,N_5275,N_5415);
xnor U6563 (N_6563,N_4601,N_3628);
nand U6564 (N_6564,N_4625,N_4469);
nor U6565 (N_6565,N_5475,N_5403);
nand U6566 (N_6566,N_3331,N_5833);
nor U6567 (N_6567,N_5788,N_3906);
nand U6568 (N_6568,N_5253,N_5968);
or U6569 (N_6569,N_5173,N_4242);
xnor U6570 (N_6570,N_4631,N_3796);
nor U6571 (N_6571,N_5126,N_3323);
and U6572 (N_6572,N_3454,N_4770);
nand U6573 (N_6573,N_4361,N_5065);
nand U6574 (N_6574,N_4273,N_3779);
nor U6575 (N_6575,N_4859,N_3425);
or U6576 (N_6576,N_4236,N_3784);
xnor U6577 (N_6577,N_4065,N_5295);
nand U6578 (N_6578,N_4030,N_4006);
nor U6579 (N_6579,N_3279,N_5435);
or U6580 (N_6580,N_5181,N_4265);
and U6581 (N_6581,N_5515,N_5524);
or U6582 (N_6582,N_3996,N_3315);
nand U6583 (N_6583,N_3667,N_5997);
and U6584 (N_6584,N_5540,N_3775);
nand U6585 (N_6585,N_5956,N_3873);
or U6586 (N_6586,N_5631,N_4947);
xnor U6587 (N_6587,N_5751,N_3541);
or U6588 (N_6588,N_4441,N_5037);
or U6589 (N_6589,N_3165,N_4181);
nor U6590 (N_6590,N_5823,N_3176);
and U6591 (N_6591,N_4460,N_3724);
nor U6592 (N_6592,N_4834,N_4161);
or U6593 (N_6593,N_4098,N_4920);
nor U6594 (N_6594,N_4379,N_4786);
nand U6595 (N_6595,N_3810,N_4203);
nor U6596 (N_6596,N_5606,N_4861);
nand U6597 (N_6597,N_5506,N_4902);
xor U6598 (N_6598,N_3294,N_3957);
nor U6599 (N_6599,N_4627,N_5969);
and U6600 (N_6600,N_3491,N_5992);
xnor U6601 (N_6601,N_3362,N_4613);
xnor U6602 (N_6602,N_4970,N_3695);
xnor U6603 (N_6603,N_4380,N_3389);
nand U6604 (N_6604,N_4893,N_5934);
or U6605 (N_6605,N_5260,N_5798);
nand U6606 (N_6606,N_4706,N_4068);
xnor U6607 (N_6607,N_3239,N_4552);
nand U6608 (N_6608,N_3320,N_5205);
and U6609 (N_6609,N_5301,N_4374);
xor U6610 (N_6610,N_3218,N_3289);
and U6611 (N_6611,N_5858,N_5433);
or U6612 (N_6612,N_3032,N_5977);
nand U6613 (N_6613,N_3240,N_3027);
xor U6614 (N_6614,N_5331,N_5479);
nand U6615 (N_6615,N_4889,N_3029);
nand U6616 (N_6616,N_4281,N_4759);
nor U6617 (N_6617,N_3096,N_5812);
and U6618 (N_6618,N_3344,N_3666);
or U6619 (N_6619,N_5231,N_4228);
nand U6620 (N_6620,N_5612,N_4758);
xor U6621 (N_6621,N_3671,N_4502);
xnor U6622 (N_6622,N_3009,N_5616);
nand U6623 (N_6623,N_3155,N_4447);
xor U6624 (N_6624,N_3704,N_3940);
nor U6625 (N_6625,N_4327,N_5434);
or U6626 (N_6626,N_3105,N_4092);
and U6627 (N_6627,N_4433,N_4213);
nand U6628 (N_6628,N_5566,N_4620);
and U6629 (N_6629,N_3874,N_4311);
nand U6630 (N_6630,N_5583,N_3864);
and U6631 (N_6631,N_4571,N_5660);
nand U6632 (N_6632,N_5110,N_5046);
or U6633 (N_6633,N_4979,N_4267);
or U6634 (N_6634,N_4344,N_5979);
and U6635 (N_6635,N_5076,N_5129);
nand U6636 (N_6636,N_4113,N_4338);
and U6637 (N_6637,N_3383,N_3828);
nand U6638 (N_6638,N_5464,N_4232);
or U6639 (N_6639,N_5681,N_4097);
and U6640 (N_6640,N_4156,N_4072);
nor U6641 (N_6641,N_4815,N_3458);
xnor U6642 (N_6642,N_4147,N_3242);
or U6643 (N_6643,N_5130,N_4964);
nor U6644 (N_6644,N_3719,N_3161);
xor U6645 (N_6645,N_5308,N_5108);
xnor U6646 (N_6646,N_5525,N_5610);
nand U6647 (N_6647,N_5269,N_5836);
xor U6648 (N_6648,N_4418,N_5040);
nand U6649 (N_6649,N_4320,N_3865);
and U6650 (N_6650,N_5149,N_5923);
nand U6651 (N_6651,N_3832,N_4259);
nand U6652 (N_6652,N_4197,N_4488);
or U6653 (N_6653,N_4343,N_3381);
and U6654 (N_6654,N_4035,N_5624);
nand U6655 (N_6655,N_5227,N_4128);
or U6656 (N_6656,N_3870,N_4251);
and U6657 (N_6657,N_4992,N_4105);
or U6658 (N_6658,N_4448,N_3000);
xor U6659 (N_6659,N_3117,N_4516);
nor U6660 (N_6660,N_5544,N_3647);
xor U6661 (N_6661,N_3110,N_3496);
nand U6662 (N_6662,N_4579,N_4173);
and U6663 (N_6663,N_4763,N_5842);
and U6664 (N_6664,N_5793,N_3840);
and U6665 (N_6665,N_5218,N_3182);
or U6666 (N_6666,N_4977,N_5819);
xnor U6667 (N_6667,N_3540,N_3558);
or U6668 (N_6668,N_4235,N_5055);
or U6669 (N_6669,N_5795,N_5667);
and U6670 (N_6670,N_3622,N_5166);
and U6671 (N_6671,N_5079,N_3013);
nand U6672 (N_6672,N_4529,N_5759);
xnor U6673 (N_6673,N_5484,N_5732);
or U6674 (N_6674,N_5206,N_5321);
or U6675 (N_6675,N_4412,N_5193);
and U6676 (N_6676,N_3016,N_5713);
and U6677 (N_6677,N_4560,N_5007);
and U6678 (N_6678,N_4034,N_3131);
and U6679 (N_6679,N_4853,N_3060);
nor U6680 (N_6680,N_3017,N_3227);
nor U6681 (N_6681,N_3824,N_4330);
xnor U6682 (N_6682,N_5654,N_5900);
and U6683 (N_6683,N_5895,N_5146);
nand U6684 (N_6684,N_3979,N_3212);
xor U6685 (N_6685,N_5143,N_4669);
or U6686 (N_6686,N_5201,N_3359);
nor U6687 (N_6687,N_3969,N_5652);
and U6688 (N_6688,N_3448,N_5690);
nand U6689 (N_6689,N_3716,N_4257);
and U6690 (N_6690,N_5441,N_3481);
nor U6691 (N_6691,N_3701,N_4305);
xnor U6692 (N_6692,N_3316,N_3128);
nor U6693 (N_6693,N_5550,N_3424);
or U6694 (N_6694,N_3702,N_5852);
xnor U6695 (N_6695,N_4886,N_3111);
nand U6696 (N_6696,N_3706,N_4037);
or U6697 (N_6697,N_3432,N_3391);
nand U6698 (N_6698,N_5635,N_3768);
nor U6699 (N_6699,N_5947,N_5741);
or U6700 (N_6700,N_4803,N_4490);
xor U6701 (N_6701,N_3882,N_3129);
and U6702 (N_6702,N_5059,N_5265);
nand U6703 (N_6703,N_5397,N_3633);
nand U6704 (N_6704,N_3656,N_4564);
nor U6705 (N_6705,N_5033,N_3908);
xnor U6706 (N_6706,N_4737,N_3981);
or U6707 (N_6707,N_3598,N_4542);
nor U6708 (N_6708,N_4753,N_3312);
xor U6709 (N_6709,N_5517,N_5644);
xnor U6710 (N_6710,N_4747,N_4046);
xor U6711 (N_6711,N_3885,N_3754);
or U6712 (N_6712,N_3521,N_4673);
nand U6713 (N_6713,N_3621,N_3728);
nand U6714 (N_6714,N_3361,N_3127);
or U6715 (N_6715,N_5413,N_5386);
and U6716 (N_6716,N_3052,N_4423);
and U6717 (N_6717,N_4721,N_5498);
and U6718 (N_6718,N_5043,N_4437);
and U6719 (N_6719,N_3891,N_4239);
nor U6720 (N_6720,N_5082,N_3629);
nor U6721 (N_6721,N_5568,N_3079);
nand U6722 (N_6722,N_4159,N_3206);
xnor U6723 (N_6723,N_5928,N_3600);
nand U6724 (N_6724,N_3282,N_5547);
xor U6725 (N_6725,N_3623,N_4445);
and U6726 (N_6726,N_5924,N_4858);
and U6727 (N_6727,N_3203,N_5656);
xor U6728 (N_6728,N_5822,N_5380);
nand U6729 (N_6729,N_5234,N_4405);
nand U6730 (N_6730,N_3962,N_4388);
or U6731 (N_6731,N_4659,N_5230);
and U6732 (N_6732,N_3512,N_3905);
or U6733 (N_6733,N_4816,N_5393);
xnor U6734 (N_6734,N_5560,N_5276);
nor U6735 (N_6735,N_4473,N_4501);
nand U6736 (N_6736,N_3640,N_4586);
and U6737 (N_6737,N_4849,N_3353);
nor U6738 (N_6738,N_4775,N_3982);
or U6739 (N_6739,N_5437,N_4767);
nand U6740 (N_6740,N_3843,N_4331);
and U6741 (N_6741,N_4254,N_4048);
xor U6742 (N_6742,N_5729,N_5049);
or U6743 (N_6743,N_3404,N_5327);
or U6744 (N_6744,N_4184,N_3074);
nand U6745 (N_6745,N_3297,N_4522);
or U6746 (N_6746,N_4553,N_4656);
and U6747 (N_6747,N_4738,N_5357);
and U6748 (N_6748,N_5362,N_3299);
and U6749 (N_6749,N_5991,N_4966);
nand U6750 (N_6750,N_4722,N_5714);
xor U6751 (N_6751,N_4024,N_5490);
xor U6752 (N_6752,N_4177,N_4955);
nand U6753 (N_6753,N_4931,N_4663);
nand U6754 (N_6754,N_4692,N_3605);
or U6755 (N_6755,N_4878,N_4555);
nor U6756 (N_6756,N_4296,N_4521);
nand U6757 (N_6757,N_3646,N_3517);
or U6758 (N_6758,N_5266,N_5843);
or U6759 (N_6759,N_4894,N_5342);
nor U6760 (N_6760,N_5211,N_4133);
xor U6761 (N_6761,N_3937,N_4733);
nand U6762 (N_6762,N_3036,N_5707);
and U6763 (N_6763,N_4079,N_5133);
or U6764 (N_6764,N_5488,N_3592);
nor U6765 (N_6765,N_4495,N_5122);
xnor U6766 (N_6766,N_4598,N_4965);
and U6767 (N_6767,N_4735,N_5715);
and U6768 (N_6768,N_4755,N_3436);
or U6769 (N_6769,N_4682,N_3204);
nor U6770 (N_6770,N_4095,N_3822);
or U6771 (N_6771,N_4252,N_4796);
or U6772 (N_6772,N_3946,N_4204);
or U6773 (N_6773,N_5519,N_3949);
xnor U6774 (N_6774,N_4091,N_5746);
nor U6775 (N_6775,N_3058,N_4255);
nand U6776 (N_6776,N_5229,N_4240);
and U6777 (N_6777,N_4002,N_5021);
and U6778 (N_6778,N_4934,N_5081);
and U6779 (N_6779,N_3416,N_4748);
xor U6780 (N_6780,N_3141,N_3596);
nor U6781 (N_6781,N_3802,N_4709);
nand U6782 (N_6782,N_4216,N_4508);
nand U6783 (N_6783,N_4230,N_5609);
nor U6784 (N_6784,N_3468,N_3926);
nand U6785 (N_6785,N_4719,N_3472);
and U6786 (N_6786,N_5378,N_3072);
nor U6787 (N_6787,N_3325,N_4507);
and U6788 (N_6788,N_3445,N_4653);
or U6789 (N_6789,N_5683,N_4517);
and U6790 (N_6790,N_3043,N_3115);
and U6791 (N_6791,N_4396,N_3618);
xnor U6792 (N_6792,N_5783,N_4616);
and U6793 (N_6793,N_5444,N_5998);
and U6794 (N_6794,N_5528,N_4665);
nand U6795 (N_6795,N_4575,N_5556);
and U6796 (N_6796,N_3505,N_3136);
xnor U6797 (N_6797,N_3764,N_3520);
xor U6798 (N_6798,N_3193,N_3763);
nand U6799 (N_6799,N_5792,N_4563);
nor U6800 (N_6800,N_3012,N_5232);
xnor U6801 (N_6801,N_4573,N_4927);
and U6802 (N_6802,N_4394,N_5356);
nand U6803 (N_6803,N_4182,N_4983);
nand U6804 (N_6804,N_5717,N_5235);
nor U6805 (N_6805,N_4795,N_3685);
or U6806 (N_6806,N_3789,N_5962);
nor U6807 (N_6807,N_5889,N_3734);
nand U6808 (N_6808,N_5679,N_3588);
nor U6809 (N_6809,N_3265,N_4641);
and U6810 (N_6810,N_5739,N_5830);
nand U6811 (N_6811,N_5596,N_4578);
nor U6812 (N_6812,N_5187,N_4695);
xnor U6813 (N_6813,N_5971,N_5069);
xnor U6814 (N_6814,N_3660,N_3319);
and U6815 (N_6815,N_3039,N_5016);
nor U6816 (N_6816,N_3153,N_5817);
nor U6817 (N_6817,N_4744,N_5249);
xnor U6818 (N_6818,N_4307,N_5555);
xnor U6819 (N_6819,N_4756,N_3601);
nor U6820 (N_6820,N_5045,N_5084);
xor U6821 (N_6821,N_4871,N_5604);
nor U6822 (N_6822,N_5585,N_5752);
xnor U6823 (N_6823,N_5864,N_3006);
or U6824 (N_6824,N_3190,N_4606);
xnor U6825 (N_6825,N_4167,N_3090);
nor U6826 (N_6826,N_3566,N_4153);
nor U6827 (N_6827,N_4452,N_3271);
nand U6828 (N_6828,N_4357,N_4662);
xor U6829 (N_6829,N_4826,N_3360);
or U6830 (N_6830,N_3314,N_4185);
or U6831 (N_6831,N_5252,N_5801);
and U6832 (N_6832,N_5099,N_4229);
nor U6833 (N_6833,N_5695,N_3457);
nand U6834 (N_6834,N_4823,N_4266);
xnor U6835 (N_6835,N_4776,N_4087);
xnor U6836 (N_6836,N_5926,N_5646);
nand U6837 (N_6837,N_5404,N_5319);
xnor U6838 (N_6838,N_5302,N_4377);
xnor U6839 (N_6839,N_4716,N_5042);
xor U6840 (N_6840,N_3195,N_5818);
or U6841 (N_6841,N_3358,N_5366);
nand U6842 (N_6842,N_5008,N_3967);
xor U6843 (N_6843,N_4471,N_3990);
nand U6844 (N_6844,N_4810,N_4556);
or U6845 (N_6845,N_4651,N_3506);
and U6846 (N_6846,N_3339,N_3394);
and U6847 (N_6847,N_5593,N_3483);
nand U6848 (N_6848,N_5142,N_4000);
nor U6849 (N_6849,N_5579,N_5391);
and U6850 (N_6850,N_5620,N_4908);
nand U6851 (N_6851,N_4058,N_4688);
xnor U6852 (N_6852,N_4045,N_5053);
or U6853 (N_6853,N_5041,N_4840);
nor U6854 (N_6854,N_5887,N_3729);
and U6855 (N_6855,N_3429,N_4458);
xnor U6856 (N_6856,N_4720,N_5500);
nand U6857 (N_6857,N_3606,N_3630);
and U6858 (N_6858,N_5496,N_3777);
or U6859 (N_6859,N_5469,N_3280);
xor U6860 (N_6860,N_3557,N_3682);
and U6861 (N_6861,N_3845,N_4264);
and U6862 (N_6862,N_3542,N_3420);
and U6863 (N_6863,N_4131,N_5156);
nand U6864 (N_6864,N_3693,N_4698);
and U6865 (N_6865,N_5467,N_3033);
xnor U6866 (N_6866,N_5712,N_4749);
or U6867 (N_6867,N_5361,N_4013);
or U6868 (N_6868,N_3614,N_3067);
nor U6869 (N_6869,N_4945,N_4392);
xor U6870 (N_6870,N_4939,N_3275);
nor U6871 (N_6871,N_5486,N_3310);
xnor U6872 (N_6872,N_3758,N_5848);
or U6873 (N_6873,N_5075,N_4482);
and U6874 (N_6874,N_5803,N_3408);
nor U6875 (N_6875,N_4480,N_5134);
nor U6876 (N_6876,N_5896,N_5048);
xor U6877 (N_6877,N_5591,N_5256);
nand U6878 (N_6878,N_5747,N_5440);
nand U6879 (N_6879,N_5373,N_3378);
or U6880 (N_6880,N_4496,N_3336);
xor U6881 (N_6881,N_5841,N_5003);
or U6882 (N_6882,N_4813,N_3899);
or U6883 (N_6883,N_4703,N_3087);
and U6884 (N_6884,N_5012,N_5144);
nand U6885 (N_6885,N_5881,N_4912);
and U6886 (N_6886,N_5530,N_5865);
and U6887 (N_6887,N_3604,N_3431);
and U6888 (N_6888,N_3401,N_3308);
and U6889 (N_6889,N_5932,N_3163);
or U6890 (N_6890,N_4788,N_4825);
nand U6891 (N_6891,N_5151,N_4940);
and U6892 (N_6892,N_5755,N_5468);
nor U6893 (N_6893,N_3743,N_3570);
nor U6894 (N_6894,N_4901,N_3186);
and U6895 (N_6895,N_3511,N_4070);
xnor U6896 (N_6896,N_3945,N_5329);
or U6897 (N_6897,N_5827,N_5424);
nand U6898 (N_6898,N_4130,N_3886);
nor U6899 (N_6899,N_4160,N_4056);
nand U6900 (N_6900,N_4066,N_5148);
nor U6901 (N_6901,N_4909,N_3364);
or U6902 (N_6902,N_3284,N_3687);
and U6903 (N_6903,N_4999,N_4051);
xor U6904 (N_6904,N_4595,N_4352);
and U6905 (N_6905,N_5450,N_5443);
nand U6906 (N_6906,N_5587,N_5874);
xor U6907 (N_6907,N_3502,N_4456);
nand U6908 (N_6908,N_4436,N_5941);
nor U6909 (N_6909,N_5141,N_5603);
nor U6910 (N_6910,N_5210,N_3236);
and U6911 (N_6911,N_4078,N_4549);
and U6912 (N_6912,N_5870,N_4314);
xnor U6913 (N_6913,N_4938,N_3998);
nor U6914 (N_6914,N_5401,N_4536);
nand U6915 (N_6915,N_4740,N_4443);
xnor U6916 (N_6916,N_5771,N_3257);
nor U6917 (N_6917,N_5137,N_4546);
nand U6918 (N_6918,N_4933,N_5559);
xnor U6919 (N_6919,N_5083,N_5692);
nand U6920 (N_6920,N_5711,N_5576);
xnor U6921 (N_6921,N_4332,N_3581);
nand U6922 (N_6922,N_4222,N_5014);
nor U6923 (N_6923,N_4520,N_5891);
nand U6924 (N_6924,N_4109,N_5066);
nor U6925 (N_6925,N_5776,N_3302);
and U6926 (N_6926,N_3798,N_5777);
or U6927 (N_6927,N_3435,N_4928);
nand U6928 (N_6928,N_3340,N_3892);
or U6929 (N_6929,N_5290,N_5114);
nand U6930 (N_6930,N_3989,N_5760);
and U6931 (N_6931,N_4978,N_5438);
nand U6932 (N_6932,N_5785,N_4607);
nand U6933 (N_6933,N_5429,N_4022);
and U6934 (N_6934,N_5728,N_4211);
or U6935 (N_6935,N_4318,N_3964);
nand U6936 (N_6936,N_4457,N_5808);
or U6937 (N_6937,N_5465,N_4500);
nand U6938 (N_6938,N_4585,N_3471);
nor U6939 (N_6939,N_3721,N_3224);
xnor U6940 (N_6940,N_5197,N_4567);
xnor U6941 (N_6941,N_4885,N_5459);
or U6942 (N_6942,N_4322,N_4116);
xnor U6943 (N_6943,N_5634,N_5800);
nand U6944 (N_6944,N_4561,N_4800);
nor U6945 (N_6945,N_5945,N_3639);
or U6946 (N_6946,N_5985,N_3277);
xor U6947 (N_6947,N_4384,N_4076);
xnor U6948 (N_6948,N_5457,N_5521);
or U6949 (N_6949,N_3341,N_3014);
nand U6950 (N_6950,N_3963,N_5988);
nand U6951 (N_6951,N_3004,N_4486);
nand U6952 (N_6952,N_5615,N_4122);
and U6953 (N_6953,N_4960,N_3560);
and U6954 (N_6954,N_3080,N_5268);
and U6955 (N_6955,N_4403,N_3583);
nor U6956 (N_6956,N_4155,N_4399);
and U6957 (N_6957,N_5725,N_5578);
xnor U6958 (N_6958,N_5038,N_4303);
nor U6959 (N_6959,N_3778,N_4093);
or U6960 (N_6960,N_3019,N_4509);
nor U6961 (N_6961,N_5091,N_5445);
or U6962 (N_6962,N_4137,N_4106);
nor U6963 (N_6963,N_5278,N_5569);
nand U6964 (N_6964,N_3410,N_5418);
or U6965 (N_6965,N_4503,N_5846);
and U6966 (N_6966,N_5855,N_3318);
nor U6967 (N_6967,N_3084,N_5549);
xnor U6968 (N_6968,N_3071,N_5948);
nor U6969 (N_6969,N_4968,N_4227);
nor U6970 (N_6970,N_4249,N_3958);
and U6971 (N_6971,N_3549,N_5854);
nand U6972 (N_6972,N_4280,N_4791);
and U6973 (N_6973,N_4476,N_5002);
nor U6974 (N_6974,N_4455,N_5913);
nand U6975 (N_6975,N_3492,N_5257);
or U6976 (N_6976,N_3180,N_5875);
nor U6977 (N_6977,N_3653,N_4752);
xnor U6978 (N_6978,N_5545,N_5013);
and U6979 (N_6979,N_3648,N_4990);
nor U6980 (N_6980,N_5976,N_4860);
and U6981 (N_6981,N_4082,N_3346);
nand U6982 (N_6982,N_3680,N_3961);
nand U6983 (N_6983,N_4638,N_4312);
and U6984 (N_6984,N_3418,N_5886);
nor U6985 (N_6985,N_3759,N_5850);
xor U6986 (N_6986,N_3766,N_3673);
or U6987 (N_6987,N_3098,N_4052);
nor U6988 (N_6988,N_3720,N_3296);
nand U6989 (N_6989,N_4158,N_3904);
or U6990 (N_6990,N_3495,N_5909);
and U6991 (N_6991,N_3194,N_5056);
and U6992 (N_6992,N_3992,N_5686);
nor U6993 (N_6993,N_5312,N_3665);
or U6994 (N_6994,N_5285,N_3544);
and U6995 (N_6995,N_5064,N_4530);
xor U6996 (N_6996,N_3928,N_3244);
nand U6997 (N_6997,N_3229,N_4001);
or U6998 (N_6998,N_3901,N_4799);
and U6999 (N_6999,N_5789,N_5105);
and U7000 (N_7000,N_5024,N_4424);
xor U7001 (N_7001,N_3399,N_3550);
nand U7002 (N_7002,N_4600,N_3148);
nand U7003 (N_7003,N_5618,N_3881);
or U7004 (N_7004,N_4597,N_3247);
or U7005 (N_7005,N_4856,N_5835);
or U7006 (N_7006,N_3848,N_5233);
or U7007 (N_7007,N_3547,N_3104);
and U7008 (N_7008,N_5967,N_5978);
xor U7009 (N_7009,N_3276,N_3552);
xnor U7010 (N_7010,N_5207,N_5794);
and U7011 (N_7011,N_4793,N_5224);
nand U7012 (N_7012,N_4550,N_5097);
xnor U7013 (N_7013,N_3861,N_5527);
and U7014 (N_7014,N_4778,N_4702);
and U7015 (N_7015,N_5706,N_5025);
nor U7016 (N_7016,N_3094,N_4783);
or U7017 (N_7017,N_5542,N_5102);
nor U7018 (N_7018,N_3615,N_3328);
and U7019 (N_7019,N_5805,N_5781);
xor U7020 (N_7020,N_5558,N_5733);
nand U7021 (N_7021,N_3479,N_3047);
or U7022 (N_7022,N_5485,N_5026);
xnor U7023 (N_7023,N_3872,N_3197);
xor U7024 (N_7024,N_3985,N_4806);
nand U7025 (N_7025,N_3249,N_4250);
xnor U7026 (N_7026,N_4083,N_4730);
nand U7027 (N_7027,N_5815,N_4351);
xor U7028 (N_7028,N_3438,N_3434);
nor U7029 (N_7029,N_3015,N_5136);
xnor U7030 (N_7030,N_5213,N_4807);
or U7031 (N_7031,N_4683,N_4845);
nor U7032 (N_7032,N_3626,N_4818);
or U7033 (N_7033,N_5581,N_3138);
nand U7034 (N_7034,N_3973,N_3059);
or U7035 (N_7035,N_4020,N_3070);
xor U7036 (N_7036,N_4841,N_4644);
or U7037 (N_7037,N_5696,N_4011);
nand U7038 (N_7038,N_3142,N_5473);
and U7039 (N_7039,N_4957,N_5153);
xor U7040 (N_7040,N_5826,N_5455);
xor U7041 (N_7041,N_3258,N_4218);
or U7042 (N_7042,N_3694,N_4400);
or U7043 (N_7043,N_3469,N_4165);
xnor U7044 (N_7044,N_4897,N_4025);
and U7045 (N_7045,N_3941,N_5200);
or U7046 (N_7046,N_5294,N_5451);
or U7047 (N_7047,N_3968,N_5299);
and U7048 (N_7048,N_4316,N_4497);
and U7049 (N_7049,N_4366,N_5492);
nand U7050 (N_7050,N_5154,N_5636);
nor U7051 (N_7051,N_4674,N_3952);
nor U7052 (N_7052,N_4772,N_4276);
and U7053 (N_7053,N_5080,N_3709);
nand U7054 (N_7054,N_3461,N_5860);
or U7055 (N_7055,N_3474,N_3591);
and U7056 (N_7056,N_5389,N_3532);
nand U7057 (N_7057,N_3167,N_3439);
nand U7058 (N_7058,N_3135,N_3587);
nor U7059 (N_7059,N_5258,N_3102);
xor U7060 (N_7060,N_3300,N_5824);
or U7061 (N_7061,N_3281,N_5015);
nand U7062 (N_7062,N_5536,N_4409);
xnor U7063 (N_7063,N_4299,N_3216);
or U7064 (N_7064,N_5987,N_5671);
nand U7065 (N_7065,N_5775,N_4736);
or U7066 (N_7066,N_5306,N_5704);
nand U7067 (N_7067,N_5377,N_5375);
and U7068 (N_7068,N_3772,N_3184);
xnor U7069 (N_7069,N_3482,N_4125);
xnor U7070 (N_7070,N_4385,N_5239);
nand U7071 (N_7071,N_4855,N_4274);
nor U7072 (N_7072,N_4801,N_4712);
xnor U7073 (N_7073,N_4183,N_5119);
nand U7074 (N_7074,N_3267,N_5938);
and U7075 (N_7075,N_3200,N_4798);
nand U7076 (N_7076,N_3924,N_4764);
nand U7077 (N_7077,N_3807,N_3902);
or U7078 (N_7078,N_4193,N_3201);
and U7079 (N_7079,N_5364,N_4432);
and U7080 (N_7080,N_4715,N_3897);
and U7081 (N_7081,N_4728,N_5878);
nand U7082 (N_7082,N_5548,N_3235);
and U7083 (N_7083,N_5573,N_4080);
and U7084 (N_7084,N_4599,N_3179);
nand U7085 (N_7085,N_4731,N_3950);
nand U7086 (N_7086,N_4477,N_3717);
xor U7087 (N_7087,N_4188,N_3177);
nand U7088 (N_7088,N_3109,N_3488);
nor U7089 (N_7089,N_5185,N_4383);
or U7090 (N_7090,N_5387,N_4724);
nand U7091 (N_7091,N_5564,N_3800);
nor U7092 (N_7092,N_4040,N_5621);
nand U7093 (N_7093,N_3050,N_3134);
nand U7094 (N_7094,N_5580,N_4935);
nand U7095 (N_7095,N_4910,N_4932);
and U7096 (N_7096,N_5990,N_3054);
and U7097 (N_7097,N_3757,N_5594);
or U7098 (N_7098,N_3400,N_3781);
or U7099 (N_7099,N_3748,N_5163);
nand U7100 (N_7100,N_5242,N_3799);
nor U7101 (N_7101,N_3228,N_3954);
xor U7102 (N_7102,N_5570,N_3711);
nor U7103 (N_7103,N_4141,N_5730);
xor U7104 (N_7104,N_3911,N_5073);
or U7105 (N_7105,N_4111,N_3269);
or U7106 (N_7106,N_4539,N_4988);
nand U7107 (N_7107,N_4918,N_4138);
and U7108 (N_7108,N_5093,N_5179);
xnor U7109 (N_7109,N_3994,N_3357);
and U7110 (N_7110,N_3168,N_3572);
or U7111 (N_7111,N_4880,N_3272);
nor U7112 (N_7112,N_5027,N_3274);
or U7113 (N_7113,N_4454,N_4835);
nand U7114 (N_7114,N_4192,N_4003);
nand U7115 (N_7115,N_5400,N_4626);
nor U7116 (N_7116,N_4174,N_5320);
nand U7117 (N_7117,N_4576,N_5502);
and U7118 (N_7118,N_5627,N_5202);
nand U7119 (N_7119,N_5884,N_5086);
nor U7120 (N_7120,N_5182,N_3516);
xnor U7121 (N_7121,N_3624,N_4504);
and U7122 (N_7122,N_4246,N_5196);
or U7123 (N_7123,N_4646,N_5328);
nor U7124 (N_7124,N_4725,N_3569);
or U7125 (N_7125,N_3372,N_3409);
xnor U7126 (N_7126,N_5347,N_5986);
and U7127 (N_7127,N_3742,N_4440);
nor U7128 (N_7128,N_5246,N_3189);
nor U7129 (N_7129,N_3884,N_3089);
nand U7130 (N_7130,N_5442,N_3567);
and U7131 (N_7131,N_3801,N_4180);
and U7132 (N_7132,N_5089,N_3918);
xnor U7133 (N_7133,N_5284,N_5238);
nor U7134 (N_7134,N_3337,N_5390);
and U7135 (N_7135,N_3960,N_4294);
and U7136 (N_7136,N_5432,N_5552);
and U7137 (N_7137,N_4963,N_3513);
or U7138 (N_7138,N_4382,N_3663);
and U7139 (N_7139,N_5688,N_4969);
xor U7140 (N_7140,N_4036,N_4150);
xnor U7141 (N_7141,N_3783,N_4205);
or U7142 (N_7142,N_3863,N_5174);
xnor U7143 (N_7143,N_3412,N_5226);
or U7144 (N_7144,N_4462,N_4054);
and U7145 (N_7145,N_4973,N_3538);
and U7146 (N_7146,N_3578,N_4911);
nand U7147 (N_7147,N_3866,N_3460);
nor U7148 (N_7148,N_5348,N_5017);
xnor U7149 (N_7149,N_5565,N_4921);
xnor U7150 (N_7150,N_5124,N_4420);
xnor U7151 (N_7151,N_5152,N_3854);
or U7152 (N_7152,N_5958,N_5655);
nand U7153 (N_7153,N_3833,N_4421);
or U7154 (N_7154,N_3652,N_4574);
and U7155 (N_7155,N_3830,N_4038);
nand U7156 (N_7156,N_4847,N_3467);
nand U7157 (N_7157,N_4824,N_5779);
or U7158 (N_7158,N_4944,N_5113);
nor U7159 (N_7159,N_5806,N_4882);
nand U7160 (N_7160,N_4936,N_3301);
or U7161 (N_7161,N_4714,N_4742);
and U7162 (N_7162,N_5392,N_4407);
nor U7163 (N_7163,N_5629,N_3813);
and U7164 (N_7164,N_3738,N_5650);
and U7165 (N_7165,N_3256,N_5352);
or U7166 (N_7166,N_5856,N_3797);
nand U7167 (N_7167,N_3334,N_3209);
xor U7168 (N_7168,N_3535,N_3669);
or U7169 (N_7169,N_3794,N_5020);
or U7170 (N_7170,N_3745,N_3419);
or U7171 (N_7171,N_4491,N_5678);
and U7172 (N_7172,N_4463,N_3137);
nor U7173 (N_7173,N_5586,N_3853);
nor U7174 (N_7174,N_5277,N_4010);
or U7175 (N_7175,N_4624,N_5734);
xor U7176 (N_7176,N_5840,N_5993);
nor U7177 (N_7177,N_5538,N_5744);
or U7178 (N_7178,N_5754,N_4145);
nor U7179 (N_7179,N_5523,N_4543);
nand U7180 (N_7180,N_5939,N_3787);
or U7181 (N_7181,N_5272,N_5742);
or U7182 (N_7182,N_4588,N_3159);
or U7183 (N_7183,N_5790,N_5271);
nor U7184 (N_7184,N_5933,N_5758);
or U7185 (N_7185,N_5028,N_4304);
xor U7186 (N_7186,N_3817,N_4061);
and U7187 (N_7187,N_4289,N_3028);
and U7188 (N_7188,N_4438,N_5482);
nor U7189 (N_7189,N_3726,N_3841);
nor U7190 (N_7190,N_5582,N_3065);
nand U7191 (N_7191,N_4633,N_4937);
and U7192 (N_7192,N_4390,N_5428);
nor U7193 (N_7193,N_5417,N_4869);
nor U7194 (N_7194,N_3169,N_3658);
nand U7195 (N_7195,N_5847,N_4987);
xor U7196 (N_7196,N_5630,N_5767);
and U7197 (N_7197,N_3133,N_5600);
and U7198 (N_7198,N_4827,N_4360);
or U7199 (N_7199,N_4693,N_3674);
and U7200 (N_7200,N_4572,N_3002);
xnor U7201 (N_7201,N_4017,N_4288);
or U7202 (N_7202,N_3651,N_4459);
nand U7203 (N_7203,N_3437,N_5123);
or U7204 (N_7204,N_3326,N_4284);
xor U7205 (N_7205,N_5248,N_3150);
nor U7206 (N_7206,N_5220,N_4754);
or U7207 (N_7207,N_5756,N_3211);
nand U7208 (N_7208,N_3991,N_4525);
xor U7209 (N_7209,N_3703,N_5381);
nor U7210 (N_7210,N_3838,N_4557);
nor U7211 (N_7211,N_5225,N_3847);
nand U7212 (N_7212,N_5409,N_3575);
nand U7213 (N_7213,N_5343,N_3368);
or U7214 (N_7214,N_3727,N_3611);
or U7215 (N_7215,N_5700,N_5989);
nor U7216 (N_7216,N_3782,N_5658);
xor U7217 (N_7217,N_3241,N_3812);
xor U7218 (N_7218,N_5336,N_4429);
and U7219 (N_7219,N_4699,N_3198);
nand U7220 (N_7220,N_5613,N_3524);
nor U7221 (N_7221,N_4123,N_4857);
nor U7222 (N_7222,N_4335,N_4906);
nor U7223 (N_7223,N_4854,N_5175);
nand U7224 (N_7224,N_3635,N_5797);
and U7225 (N_7225,N_3553,N_5150);
nand U7226 (N_7226,N_4707,N_4689);
and U7227 (N_7227,N_3586,N_4408);
nor U7228 (N_7228,N_5237,N_3839);
and U7229 (N_7229,N_5637,N_5796);
or U7230 (N_7230,N_5994,N_3691);
or U7231 (N_7231,N_3956,N_3816);
or U7232 (N_7232,N_3805,N_4102);
or U7233 (N_7233,N_4247,N_5369);
or U7234 (N_7234,N_4888,N_3225);
nand U7235 (N_7235,N_4570,N_3092);
xnor U7236 (N_7236,N_4628,N_4126);
xor U7237 (N_7237,N_4577,N_3850);
nor U7238 (N_7238,N_5335,N_3405);
or U7239 (N_7239,N_3883,N_5663);
nand U7240 (N_7240,N_3441,N_5791);
xnor U7241 (N_7241,N_5952,N_3395);
or U7242 (N_7242,N_4609,N_4483);
xor U7243 (N_7243,N_5643,N_5577);
xnor U7244 (N_7244,N_5664,N_4694);
nor U7245 (N_7245,N_3442,N_4870);
xnor U7246 (N_7246,N_5458,N_3093);
xnor U7247 (N_7247,N_3175,N_3773);
xor U7248 (N_7248,N_5460,N_4547);
nor U7249 (N_7249,N_3860,N_4797);
xor U7250 (N_7250,N_3529,N_5106);
nor U7251 (N_7251,N_4916,N_4828);
and U7252 (N_7252,N_3423,N_3933);
nor U7253 (N_7253,N_3348,N_3288);
or U7254 (N_7254,N_3966,N_4761);
nor U7255 (N_7255,N_5647,N_5395);
xnor U7256 (N_7256,N_3494,N_5872);
xor U7257 (N_7257,N_5350,N_3031);
and U7258 (N_7258,N_5051,N_5117);
or U7259 (N_7259,N_3473,N_5888);
xor U7260 (N_7260,N_4781,N_3735);
nor U7261 (N_7261,N_5215,N_4321);
xnor U7262 (N_7262,N_4643,N_3948);
and U7263 (N_7263,N_5825,N_3443);
nand U7264 (N_7264,N_5735,N_5161);
nor U7265 (N_7265,N_4941,N_5120);
nor U7266 (N_7266,N_5461,N_4146);
xor U7267 (N_7267,N_4681,N_3655);
nor U7268 (N_7268,N_4948,N_5245);
nand U7269 (N_7269,N_3739,N_4619);
and U7270 (N_7270,N_3049,N_5661);
nor U7271 (N_7271,N_4612,N_3449);
nor U7272 (N_7272,N_4881,N_4349);
and U7273 (N_7273,N_3856,N_4954);
nor U7274 (N_7274,N_4804,N_4107);
xnor U7275 (N_7275,N_4256,N_5983);
nand U7276 (N_7276,N_3034,N_5653);
xnor U7277 (N_7277,N_3215,N_4470);
and U7278 (N_7278,N_4822,N_3385);
or U7279 (N_7279,N_4506,N_4650);
and U7280 (N_7280,N_3915,N_5353);
nand U7281 (N_7281,N_5935,N_4444);
nand U7282 (N_7282,N_4809,N_3632);
and U7283 (N_7283,N_3030,N_3608);
xnor U7284 (N_7284,N_5480,N_5931);
and U7285 (N_7285,N_3718,N_4868);
nand U7286 (N_7286,N_5318,N_4231);
nor U7287 (N_7287,N_5682,N_4925);
xor U7288 (N_7288,N_5838,N_5162);
and U7289 (N_7289,N_4132,N_5633);
and U7290 (N_7290,N_5857,N_4995);
and U7291 (N_7291,N_3510,N_3147);
nand U7292 (N_7292,N_3857,N_4895);
nor U7293 (N_7293,N_5282,N_5140);
and U7294 (N_7294,N_4708,N_3823);
nor U7295 (N_7295,N_4985,N_4734);
or U7296 (N_7296,N_3662,N_3152);
nand U7297 (N_7297,N_4370,N_3895);
and U7298 (N_7298,N_5001,N_3852);
nor U7299 (N_7299,N_3649,N_3776);
nand U7300 (N_7300,N_4329,N_4442);
nand U7301 (N_7301,N_4151,N_3780);
xnor U7302 (N_7302,N_4879,N_5169);
nand U7303 (N_7303,N_4090,N_3106);
and U7304 (N_7304,N_5493,N_3657);
or U7305 (N_7305,N_4450,N_5764);
nor U7306 (N_7306,N_5740,N_4711);
and U7307 (N_7307,N_4566,N_5067);
nand U7308 (N_7308,N_3747,N_4837);
and U7309 (N_7309,N_5060,N_3370);
nor U7310 (N_7310,N_5034,N_4021);
and U7311 (N_7311,N_5463,N_3858);
xnor U7312 (N_7312,N_5495,N_4485);
xnor U7313 (N_7313,N_5877,N_4610);
and U7314 (N_7314,N_4867,N_5807);
nand U7315 (N_7315,N_4094,N_5944);
or U7316 (N_7316,N_4967,N_5965);
and U7317 (N_7317,N_3842,N_5228);
xnor U7318 (N_7318,N_3580,N_4244);
and U7319 (N_7319,N_5930,N_3645);
nand U7320 (N_7320,N_5804,N_3976);
and U7321 (N_7321,N_3879,N_3026);
xor U7322 (N_7322,N_4027,N_5453);
nand U7323 (N_7323,N_5649,N_4434);
and U7324 (N_7324,N_5270,N_5531);
nor U7325 (N_7325,N_3698,N_4887);
and U7326 (N_7326,N_4047,N_4907);
nor U7327 (N_7327,N_3767,N_3191);
or U7328 (N_7328,N_5309,N_5910);
nand U7329 (N_7329,N_5384,N_3485);
or U7330 (N_7330,N_4328,N_3821);
and U7331 (N_7331,N_3672,N_5420);
and U7332 (N_7332,N_4439,N_3751);
nor U7333 (N_7333,N_3306,N_4170);
xor U7334 (N_7334,N_4373,N_5906);
xnor U7335 (N_7335,N_3121,N_4534);
or U7336 (N_7336,N_4175,N_3100);
nor U7337 (N_7337,N_5588,N_5672);
nor U7338 (N_7338,N_3546,N_4041);
and U7339 (N_7339,N_5546,N_3803);
and U7340 (N_7340,N_4481,N_5011);
nor U7341 (N_7341,N_5602,N_5410);
nand U7342 (N_7342,N_5628,N_5981);
or U7343 (N_7343,N_4984,N_4592);
xor U7344 (N_7344,N_3913,N_3363);
or U7345 (N_7345,N_5773,N_3465);
or U7346 (N_7346,N_5374,N_5297);
nor U7347 (N_7347,N_4639,N_4562);
nand U7348 (N_7348,N_4214,N_5330);
or U7349 (N_7349,N_5221,N_5385);
nand U7350 (N_7350,N_4248,N_4745);
nand U7351 (N_7351,N_3965,N_3675);
nand U7352 (N_7352,N_4511,N_4843);
nand U7353 (N_7353,N_5280,N_4768);
nor U7354 (N_7354,N_4042,N_3366);
and U7355 (N_7355,N_3170,N_4671);
or U7356 (N_7356,N_5078,N_4142);
xnor U7357 (N_7357,N_4883,N_5503);
xor U7358 (N_7358,N_3811,N_5722);
and U7359 (N_7359,N_3790,N_5899);
nand U7360 (N_7360,N_5405,N_5632);
and U7361 (N_7361,N_3988,N_4660);
and U7362 (N_7362,N_3597,N_4532);
xnor U7363 (N_7363,N_3303,N_3417);
nor U7364 (N_7364,N_5851,N_5639);
or U7365 (N_7365,N_4018,N_3250);
nand U7366 (N_7366,N_5135,N_5959);
or U7367 (N_7367,N_5697,N_3259);
or U7368 (N_7368,N_3233,N_4569);
and U7369 (N_7369,N_4952,N_3045);
and U7370 (N_7370,N_4872,N_5421);
xor U7371 (N_7371,N_5351,N_5942);
or U7372 (N_7372,N_3620,N_3929);
nor U7373 (N_7373,N_4686,N_5762);
and U7374 (N_7374,N_4670,N_3387);
and U7375 (N_7375,N_3525,N_5035);
or U7376 (N_7376,N_4363,N_5094);
xor U7377 (N_7377,N_4430,N_5611);
xnor U7378 (N_7378,N_5047,N_4917);
nand U7379 (N_7379,N_3795,N_4997);
nand U7380 (N_7380,N_5411,N_4648);
xor U7381 (N_7381,N_4063,N_3770);
xor U7382 (N_7382,N_3514,N_3475);
nand U7383 (N_7383,N_5839,N_5645);
and U7384 (N_7384,N_4472,N_5782);
nor U7385 (N_7385,N_5068,N_3668);
or U7386 (N_7386,N_5504,N_4282);
nor U7387 (N_7387,N_5497,N_3187);
nor U7388 (N_7388,N_3130,N_4215);
nor U7389 (N_7389,N_4171,N_3890);
and U7390 (N_7390,N_5853,N_3476);
xor U7391 (N_7391,N_4465,N_3819);
and U7392 (N_7392,N_3888,N_4031);
xor U7393 (N_7393,N_3261,N_5648);
xor U7394 (N_7394,N_4584,N_3352);
xnor U7395 (N_7395,N_5439,N_3455);
nand U7396 (N_7396,N_5388,N_4397);
or U7397 (N_7397,N_3793,N_4134);
nor U7398 (N_7398,N_3309,N_4345);
or U7399 (N_7399,N_3287,N_3930);
nor U7400 (N_7400,N_3877,N_3291);
nand U7401 (N_7401,N_5074,N_5589);
nand U7402 (N_7402,N_3942,N_4832);
or U7403 (N_7403,N_5287,N_3486);
or U7404 (N_7404,N_5786,N_4272);
xnor U7405 (N_7405,N_5943,N_5572);
nor U7406 (N_7406,N_4873,N_3196);
xnor U7407 (N_7407,N_4510,N_5964);
nand U7408 (N_7408,N_5168,N_5737);
xor U7409 (N_7409,N_4864,N_4515);
or U7410 (N_7410,N_4009,N_4946);
or U7411 (N_7411,N_3384,N_4757);
nor U7412 (N_7412,N_4302,N_4591);
xnor U7413 (N_7413,N_4313,N_3414);
and U7414 (N_7414,N_3528,N_5598);
or U7415 (N_7415,N_4053,N_3063);
or U7416 (N_7416,N_4489,N_5062);
and U7417 (N_7417,N_4200,N_5293);
or U7418 (N_7418,N_3616,N_5859);
and U7419 (N_7419,N_3752,N_3603);
nor U7420 (N_7420,N_3278,N_3076);
and U7421 (N_7421,N_4064,N_4164);
nor U7422 (N_7422,N_3178,N_5508);
xnor U7423 (N_7423,N_3066,N_3330);
xor U7424 (N_7424,N_5436,N_5505);
or U7425 (N_7425,N_4308,N_3415);
and U7426 (N_7426,N_4905,N_5638);
and U7427 (N_7427,N_5192,N_3922);
nor U7428 (N_7428,N_3744,N_4212);
xor U7429 (N_7429,N_3593,N_4615);
nor U7430 (N_7430,N_3809,N_3255);
or U7431 (N_7431,N_4684,N_3199);
nor U7432 (N_7432,N_3923,N_4190);
or U7433 (N_7433,N_4253,N_3543);
xor U7434 (N_7434,N_5551,N_3862);
and U7435 (N_7435,N_4766,N_3382);
nand U7436 (N_7436,N_4587,N_3390);
or U7437 (N_7437,N_3114,N_4419);
and U7438 (N_7438,N_5107,N_3746);
xnor U7439 (N_7439,N_5908,N_5509);
nand U7440 (N_7440,N_5273,N_4012);
nand U7441 (N_7441,N_3406,N_4475);
nor U7442 (N_7442,N_4148,N_5937);
xor U7443 (N_7443,N_5399,N_5902);
and U7444 (N_7444,N_3459,N_5030);
nor U7445 (N_7445,N_3518,N_3750);
nand U7446 (N_7446,N_5398,N_4771);
and U7447 (N_7447,N_4262,N_5022);
and U7448 (N_7448,N_4059,N_4194);
xnor U7449 (N_7449,N_5147,N_3880);
nor U7450 (N_7450,N_4067,N_3125);
and U7451 (N_7451,N_3223,N_3700);
xnor U7452 (N_7452,N_3327,N_5472);
nand U7453 (N_7453,N_5254,N_4176);
or U7454 (N_7454,N_5513,N_5072);
or U7455 (N_7455,N_5165,N_5180);
xnor U7456 (N_7456,N_5657,N_3112);
nor U7457 (N_7457,N_3736,N_4913);
xor U7458 (N_7458,N_3252,N_3447);
and U7459 (N_7459,N_3497,N_4678);
or U7460 (N_7460,N_4189,N_5575);
xor U7461 (N_7461,N_3185,N_4416);
nor U7462 (N_7462,N_4580,N_5557);
or U7463 (N_7463,N_5109,N_3001);
or U7464 (N_7464,N_5009,N_3970);
nor U7465 (N_7465,N_3679,N_5625);
or U7466 (N_7466,N_4787,N_5861);
or U7467 (N_7467,N_4499,N_5100);
or U7468 (N_7468,N_3324,N_5980);
xnor U7469 (N_7469,N_3936,N_5567);
and U7470 (N_7470,N_3487,N_5828);
and U7471 (N_7471,N_3075,N_4838);
nand U7472 (N_7472,N_3504,N_5999);
nand U7473 (N_7473,N_5212,N_3659);
nand U7474 (N_7474,N_4413,N_4238);
or U7475 (N_7475,N_3018,N_5599);
nor U7476 (N_7476,N_4924,N_3636);
nor U7477 (N_7477,N_4356,N_3536);
xnor U7478 (N_7478,N_4779,N_3046);
xnor U7479 (N_7479,N_3997,N_4558);
or U7480 (N_7480,N_4287,N_3091);
nand U7481 (N_7481,N_4980,N_3681);
or U7482 (N_7482,N_3531,N_4152);
and U7483 (N_7483,N_5376,N_3490);
nand U7484 (N_7484,N_3509,N_4523);
nand U7485 (N_7485,N_5198,N_3522);
nand U7486 (N_7486,N_3413,N_3020);
and U7487 (N_7487,N_4004,N_5778);
nand U7488 (N_7488,N_3171,N_3107);
and U7489 (N_7489,N_4224,N_5966);
xor U7490 (N_7490,N_5250,N_5915);
nand U7491 (N_7491,N_5936,N_4406);
xnor U7492 (N_7492,N_3377,N_5614);
nand U7493 (N_7493,N_3499,N_4513);
xnor U7494 (N_7494,N_4210,N_5766);
nor U7495 (N_7495,N_4198,N_5316);
nor U7496 (N_7496,N_5675,N_3733);
nor U7497 (N_7497,N_3081,N_4269);
xor U7498 (N_7498,N_5584,N_5340);
and U7499 (N_7499,N_3003,N_3519);
or U7500 (N_7500,N_5764,N_4083);
nor U7501 (N_7501,N_5980,N_3028);
xnor U7502 (N_7502,N_4213,N_5534);
or U7503 (N_7503,N_3839,N_5050);
or U7504 (N_7504,N_4791,N_5688);
xnor U7505 (N_7505,N_5335,N_5672);
nand U7506 (N_7506,N_3963,N_5277);
and U7507 (N_7507,N_5321,N_4830);
nand U7508 (N_7508,N_4827,N_5696);
nor U7509 (N_7509,N_4339,N_5328);
xnor U7510 (N_7510,N_5620,N_4752);
and U7511 (N_7511,N_4410,N_3360);
nand U7512 (N_7512,N_5363,N_5410);
nor U7513 (N_7513,N_4273,N_3072);
or U7514 (N_7514,N_4024,N_4874);
nand U7515 (N_7515,N_3375,N_5857);
nor U7516 (N_7516,N_4467,N_4481);
and U7517 (N_7517,N_5505,N_3874);
nor U7518 (N_7518,N_4522,N_3185);
xnor U7519 (N_7519,N_5903,N_5103);
nor U7520 (N_7520,N_5288,N_5353);
xnor U7521 (N_7521,N_5540,N_5341);
and U7522 (N_7522,N_5351,N_3112);
and U7523 (N_7523,N_3713,N_4122);
and U7524 (N_7524,N_4950,N_5327);
nand U7525 (N_7525,N_3789,N_3992);
and U7526 (N_7526,N_4969,N_5580);
or U7527 (N_7527,N_3875,N_4783);
nand U7528 (N_7528,N_4034,N_4062);
nand U7529 (N_7529,N_3091,N_5608);
nand U7530 (N_7530,N_5984,N_3305);
nor U7531 (N_7531,N_4592,N_5628);
or U7532 (N_7532,N_4542,N_5424);
nand U7533 (N_7533,N_4200,N_3650);
nor U7534 (N_7534,N_4184,N_3601);
or U7535 (N_7535,N_4421,N_4074);
nor U7536 (N_7536,N_4489,N_5028);
nand U7537 (N_7537,N_3343,N_4666);
nor U7538 (N_7538,N_4667,N_4207);
nand U7539 (N_7539,N_3235,N_4548);
or U7540 (N_7540,N_5525,N_4399);
nand U7541 (N_7541,N_4905,N_4371);
nand U7542 (N_7542,N_4756,N_5746);
nand U7543 (N_7543,N_5087,N_4257);
nand U7544 (N_7544,N_3998,N_4686);
nor U7545 (N_7545,N_3244,N_3293);
nand U7546 (N_7546,N_5975,N_5836);
xnor U7547 (N_7547,N_3409,N_5658);
nand U7548 (N_7548,N_4820,N_5551);
xnor U7549 (N_7549,N_3053,N_3888);
nor U7550 (N_7550,N_3820,N_5781);
xor U7551 (N_7551,N_3211,N_5021);
and U7552 (N_7552,N_5290,N_5317);
or U7553 (N_7553,N_3753,N_4212);
and U7554 (N_7554,N_4621,N_4878);
or U7555 (N_7555,N_4467,N_5060);
nand U7556 (N_7556,N_5359,N_4613);
nor U7557 (N_7557,N_3457,N_5027);
nand U7558 (N_7558,N_3357,N_4506);
xor U7559 (N_7559,N_5487,N_5418);
nand U7560 (N_7560,N_4151,N_4352);
and U7561 (N_7561,N_3547,N_4851);
nand U7562 (N_7562,N_4812,N_4112);
and U7563 (N_7563,N_3398,N_4584);
and U7564 (N_7564,N_3767,N_3531);
nand U7565 (N_7565,N_3667,N_4064);
or U7566 (N_7566,N_4437,N_3975);
xor U7567 (N_7567,N_5848,N_5980);
nor U7568 (N_7568,N_4890,N_5909);
or U7569 (N_7569,N_5727,N_4396);
nand U7570 (N_7570,N_3116,N_5233);
and U7571 (N_7571,N_5225,N_4905);
nor U7572 (N_7572,N_3577,N_3162);
and U7573 (N_7573,N_5972,N_3303);
xor U7574 (N_7574,N_5899,N_3329);
nor U7575 (N_7575,N_3951,N_3964);
and U7576 (N_7576,N_3639,N_4770);
nand U7577 (N_7577,N_5515,N_4904);
or U7578 (N_7578,N_5222,N_5978);
nor U7579 (N_7579,N_3849,N_5739);
xnor U7580 (N_7580,N_5247,N_4697);
xnor U7581 (N_7581,N_5664,N_5686);
xnor U7582 (N_7582,N_4212,N_3773);
nor U7583 (N_7583,N_5941,N_4896);
and U7584 (N_7584,N_4362,N_5822);
nor U7585 (N_7585,N_5615,N_4845);
or U7586 (N_7586,N_4085,N_4522);
and U7587 (N_7587,N_4122,N_3139);
or U7588 (N_7588,N_3285,N_4502);
and U7589 (N_7589,N_5817,N_5703);
or U7590 (N_7590,N_4803,N_4160);
or U7591 (N_7591,N_5854,N_4207);
or U7592 (N_7592,N_3020,N_3127);
nor U7593 (N_7593,N_3283,N_4266);
nor U7594 (N_7594,N_5278,N_5894);
or U7595 (N_7595,N_3385,N_4053);
nor U7596 (N_7596,N_5335,N_5604);
nor U7597 (N_7597,N_4298,N_5888);
xnor U7598 (N_7598,N_5281,N_4743);
nor U7599 (N_7599,N_4187,N_4351);
xor U7600 (N_7600,N_3107,N_4740);
nor U7601 (N_7601,N_5195,N_5582);
or U7602 (N_7602,N_3439,N_3919);
nand U7603 (N_7603,N_4820,N_4137);
nand U7604 (N_7604,N_5635,N_5585);
and U7605 (N_7605,N_4971,N_5942);
nand U7606 (N_7606,N_4067,N_5121);
xor U7607 (N_7607,N_4982,N_5696);
xnor U7608 (N_7608,N_5995,N_3891);
nand U7609 (N_7609,N_5761,N_4528);
and U7610 (N_7610,N_4773,N_4302);
and U7611 (N_7611,N_5862,N_4508);
nand U7612 (N_7612,N_3719,N_5594);
or U7613 (N_7613,N_4794,N_4068);
xnor U7614 (N_7614,N_3035,N_3918);
and U7615 (N_7615,N_3092,N_5252);
xor U7616 (N_7616,N_3632,N_5470);
and U7617 (N_7617,N_5599,N_5291);
xnor U7618 (N_7618,N_4497,N_4254);
nor U7619 (N_7619,N_5429,N_5716);
nor U7620 (N_7620,N_5618,N_4332);
nor U7621 (N_7621,N_4019,N_3275);
and U7622 (N_7622,N_3713,N_5460);
nand U7623 (N_7623,N_3126,N_4685);
xor U7624 (N_7624,N_5871,N_5171);
nor U7625 (N_7625,N_3883,N_3485);
and U7626 (N_7626,N_3655,N_4726);
or U7627 (N_7627,N_3065,N_3428);
nand U7628 (N_7628,N_4565,N_3381);
nand U7629 (N_7629,N_5376,N_3389);
nand U7630 (N_7630,N_4649,N_4560);
or U7631 (N_7631,N_3341,N_5129);
and U7632 (N_7632,N_5967,N_4439);
nor U7633 (N_7633,N_3329,N_4935);
or U7634 (N_7634,N_5502,N_4572);
nor U7635 (N_7635,N_4602,N_4407);
xnor U7636 (N_7636,N_4568,N_4153);
and U7637 (N_7637,N_5166,N_5651);
or U7638 (N_7638,N_4989,N_3045);
nor U7639 (N_7639,N_3261,N_4222);
nor U7640 (N_7640,N_5582,N_3617);
nand U7641 (N_7641,N_3413,N_4210);
or U7642 (N_7642,N_4002,N_5443);
xnor U7643 (N_7643,N_3687,N_3681);
or U7644 (N_7644,N_3803,N_4236);
xor U7645 (N_7645,N_3076,N_5176);
xor U7646 (N_7646,N_3261,N_5549);
xnor U7647 (N_7647,N_5124,N_5077);
nor U7648 (N_7648,N_4957,N_5193);
nand U7649 (N_7649,N_4397,N_4263);
nand U7650 (N_7650,N_4243,N_4244);
nor U7651 (N_7651,N_5397,N_4127);
xnor U7652 (N_7652,N_4827,N_3696);
or U7653 (N_7653,N_3000,N_3976);
or U7654 (N_7654,N_4172,N_4511);
or U7655 (N_7655,N_4357,N_4800);
nand U7656 (N_7656,N_5376,N_3728);
nor U7657 (N_7657,N_5290,N_4650);
or U7658 (N_7658,N_5367,N_4568);
xor U7659 (N_7659,N_4976,N_5088);
and U7660 (N_7660,N_3504,N_3129);
nor U7661 (N_7661,N_3050,N_3209);
nand U7662 (N_7662,N_3388,N_4761);
or U7663 (N_7663,N_3669,N_3941);
and U7664 (N_7664,N_5618,N_3187);
and U7665 (N_7665,N_5909,N_4826);
nor U7666 (N_7666,N_5125,N_5472);
nand U7667 (N_7667,N_5308,N_4038);
and U7668 (N_7668,N_4287,N_4752);
nand U7669 (N_7669,N_5319,N_5147);
or U7670 (N_7670,N_4773,N_4536);
or U7671 (N_7671,N_3462,N_4656);
or U7672 (N_7672,N_4023,N_3386);
nor U7673 (N_7673,N_3917,N_4698);
and U7674 (N_7674,N_3975,N_3172);
nand U7675 (N_7675,N_4623,N_3778);
nand U7676 (N_7676,N_5178,N_5863);
nor U7677 (N_7677,N_3027,N_3196);
nand U7678 (N_7678,N_5290,N_5671);
and U7679 (N_7679,N_3965,N_5001);
and U7680 (N_7680,N_4761,N_3871);
or U7681 (N_7681,N_3307,N_5452);
nor U7682 (N_7682,N_5119,N_3041);
nand U7683 (N_7683,N_4764,N_4728);
and U7684 (N_7684,N_4213,N_4666);
and U7685 (N_7685,N_5825,N_3955);
nand U7686 (N_7686,N_3153,N_5273);
nand U7687 (N_7687,N_5995,N_4490);
nor U7688 (N_7688,N_5944,N_3672);
or U7689 (N_7689,N_3821,N_4508);
nand U7690 (N_7690,N_4050,N_3084);
nor U7691 (N_7691,N_5614,N_3425);
xor U7692 (N_7692,N_4601,N_3966);
or U7693 (N_7693,N_3165,N_3060);
and U7694 (N_7694,N_4296,N_3990);
xor U7695 (N_7695,N_5353,N_5726);
and U7696 (N_7696,N_4736,N_4155);
nand U7697 (N_7697,N_4420,N_4732);
nand U7698 (N_7698,N_5871,N_4709);
or U7699 (N_7699,N_3822,N_4942);
or U7700 (N_7700,N_4292,N_3037);
nor U7701 (N_7701,N_3564,N_5606);
xnor U7702 (N_7702,N_5610,N_4759);
or U7703 (N_7703,N_4739,N_4856);
and U7704 (N_7704,N_3764,N_5678);
nand U7705 (N_7705,N_4897,N_5262);
xnor U7706 (N_7706,N_5587,N_5772);
xnor U7707 (N_7707,N_3761,N_3484);
or U7708 (N_7708,N_3758,N_3409);
nand U7709 (N_7709,N_3230,N_5677);
nor U7710 (N_7710,N_5818,N_4817);
nor U7711 (N_7711,N_4688,N_4550);
and U7712 (N_7712,N_3780,N_5054);
or U7713 (N_7713,N_4477,N_3119);
xor U7714 (N_7714,N_3516,N_5860);
xor U7715 (N_7715,N_5786,N_5740);
and U7716 (N_7716,N_5957,N_5432);
nand U7717 (N_7717,N_5746,N_4539);
nand U7718 (N_7718,N_4575,N_4835);
or U7719 (N_7719,N_5977,N_5806);
and U7720 (N_7720,N_3172,N_3434);
or U7721 (N_7721,N_4841,N_4326);
xnor U7722 (N_7722,N_5582,N_3789);
nand U7723 (N_7723,N_3135,N_4619);
nor U7724 (N_7724,N_5263,N_3494);
nand U7725 (N_7725,N_5499,N_3497);
xor U7726 (N_7726,N_4456,N_5061);
or U7727 (N_7727,N_5394,N_4014);
or U7728 (N_7728,N_3259,N_4481);
nand U7729 (N_7729,N_3888,N_5981);
or U7730 (N_7730,N_5485,N_4617);
nand U7731 (N_7731,N_5989,N_4921);
and U7732 (N_7732,N_3125,N_5820);
xor U7733 (N_7733,N_5675,N_3040);
or U7734 (N_7734,N_5636,N_3673);
or U7735 (N_7735,N_4159,N_5823);
nand U7736 (N_7736,N_4243,N_5524);
xor U7737 (N_7737,N_3713,N_3273);
nand U7738 (N_7738,N_4039,N_4403);
or U7739 (N_7739,N_3399,N_5639);
xor U7740 (N_7740,N_4282,N_4319);
or U7741 (N_7741,N_3744,N_3827);
nor U7742 (N_7742,N_3847,N_4481);
or U7743 (N_7743,N_3992,N_3312);
nor U7744 (N_7744,N_5538,N_4540);
or U7745 (N_7745,N_5120,N_3839);
xnor U7746 (N_7746,N_5898,N_3894);
nand U7747 (N_7747,N_4542,N_5929);
nand U7748 (N_7748,N_5907,N_5249);
and U7749 (N_7749,N_5178,N_3663);
and U7750 (N_7750,N_3094,N_3568);
xnor U7751 (N_7751,N_5979,N_5005);
or U7752 (N_7752,N_3190,N_5608);
nor U7753 (N_7753,N_5341,N_4851);
nor U7754 (N_7754,N_4622,N_4791);
xnor U7755 (N_7755,N_4135,N_3324);
and U7756 (N_7756,N_5087,N_5953);
xor U7757 (N_7757,N_3432,N_3073);
nand U7758 (N_7758,N_4726,N_5547);
xor U7759 (N_7759,N_5279,N_4711);
nor U7760 (N_7760,N_5397,N_3879);
xnor U7761 (N_7761,N_3255,N_3861);
and U7762 (N_7762,N_5930,N_5433);
and U7763 (N_7763,N_4684,N_4586);
or U7764 (N_7764,N_3070,N_5852);
xnor U7765 (N_7765,N_3303,N_5169);
nand U7766 (N_7766,N_3096,N_4212);
xnor U7767 (N_7767,N_3043,N_4386);
nor U7768 (N_7768,N_5858,N_5425);
and U7769 (N_7769,N_5234,N_3074);
nand U7770 (N_7770,N_5230,N_4832);
nand U7771 (N_7771,N_3490,N_3801);
or U7772 (N_7772,N_3988,N_4643);
xnor U7773 (N_7773,N_3562,N_5735);
nand U7774 (N_7774,N_4698,N_5247);
nor U7775 (N_7775,N_3211,N_4639);
nand U7776 (N_7776,N_5772,N_5430);
nor U7777 (N_7777,N_3752,N_3646);
or U7778 (N_7778,N_4199,N_4161);
nor U7779 (N_7779,N_4924,N_4655);
nand U7780 (N_7780,N_4859,N_4203);
and U7781 (N_7781,N_3555,N_3061);
or U7782 (N_7782,N_5230,N_5867);
nor U7783 (N_7783,N_5303,N_3345);
xnor U7784 (N_7784,N_5836,N_5724);
and U7785 (N_7785,N_4081,N_5695);
nor U7786 (N_7786,N_4554,N_3108);
nor U7787 (N_7787,N_5236,N_4944);
nand U7788 (N_7788,N_3231,N_3598);
xnor U7789 (N_7789,N_4870,N_5768);
nand U7790 (N_7790,N_5929,N_3388);
nor U7791 (N_7791,N_5058,N_5002);
or U7792 (N_7792,N_4189,N_3749);
nor U7793 (N_7793,N_4024,N_5342);
or U7794 (N_7794,N_3803,N_3970);
or U7795 (N_7795,N_5721,N_3403);
nor U7796 (N_7796,N_3453,N_3181);
xnor U7797 (N_7797,N_4788,N_3201);
nor U7798 (N_7798,N_4415,N_3415);
nor U7799 (N_7799,N_3463,N_3193);
nand U7800 (N_7800,N_4116,N_3267);
nor U7801 (N_7801,N_5335,N_4909);
and U7802 (N_7802,N_3667,N_3702);
xnor U7803 (N_7803,N_4582,N_5568);
nor U7804 (N_7804,N_3599,N_4136);
xnor U7805 (N_7805,N_5325,N_5092);
xnor U7806 (N_7806,N_5380,N_4415);
or U7807 (N_7807,N_3289,N_4268);
nor U7808 (N_7808,N_3676,N_5292);
xor U7809 (N_7809,N_5229,N_5519);
nand U7810 (N_7810,N_5702,N_5258);
or U7811 (N_7811,N_5116,N_3720);
or U7812 (N_7812,N_3297,N_3361);
xor U7813 (N_7813,N_3544,N_5402);
or U7814 (N_7814,N_5091,N_3846);
and U7815 (N_7815,N_5167,N_3190);
nor U7816 (N_7816,N_3838,N_3483);
or U7817 (N_7817,N_5060,N_3734);
nor U7818 (N_7818,N_5450,N_5275);
or U7819 (N_7819,N_5728,N_5814);
nand U7820 (N_7820,N_4857,N_5771);
xnor U7821 (N_7821,N_3915,N_4512);
or U7822 (N_7822,N_5365,N_5102);
or U7823 (N_7823,N_4068,N_5598);
nor U7824 (N_7824,N_5440,N_4947);
or U7825 (N_7825,N_4651,N_3191);
nor U7826 (N_7826,N_3509,N_3414);
or U7827 (N_7827,N_4681,N_3846);
nand U7828 (N_7828,N_4371,N_4662);
or U7829 (N_7829,N_5115,N_5393);
nand U7830 (N_7830,N_5715,N_3148);
and U7831 (N_7831,N_5292,N_4484);
or U7832 (N_7832,N_3553,N_5412);
xor U7833 (N_7833,N_3530,N_3112);
or U7834 (N_7834,N_4267,N_3519);
xnor U7835 (N_7835,N_3987,N_3265);
and U7836 (N_7836,N_5456,N_4774);
nor U7837 (N_7837,N_4559,N_3834);
nand U7838 (N_7838,N_5845,N_3460);
nand U7839 (N_7839,N_5989,N_4624);
nor U7840 (N_7840,N_4014,N_5015);
xnor U7841 (N_7841,N_4684,N_5227);
nor U7842 (N_7842,N_3346,N_5573);
xnor U7843 (N_7843,N_4777,N_3839);
xnor U7844 (N_7844,N_3886,N_5425);
xnor U7845 (N_7845,N_5018,N_4883);
nand U7846 (N_7846,N_4268,N_5857);
and U7847 (N_7847,N_5178,N_3979);
or U7848 (N_7848,N_4893,N_4488);
or U7849 (N_7849,N_4943,N_5335);
xnor U7850 (N_7850,N_4211,N_4461);
nand U7851 (N_7851,N_3183,N_4774);
and U7852 (N_7852,N_4338,N_4789);
nand U7853 (N_7853,N_4987,N_4049);
nand U7854 (N_7854,N_5213,N_3878);
or U7855 (N_7855,N_5197,N_5135);
or U7856 (N_7856,N_3861,N_4006);
nand U7857 (N_7857,N_3300,N_3499);
and U7858 (N_7858,N_5472,N_4722);
and U7859 (N_7859,N_4756,N_4446);
nand U7860 (N_7860,N_5500,N_4311);
nor U7861 (N_7861,N_4851,N_5695);
and U7862 (N_7862,N_5293,N_3380);
or U7863 (N_7863,N_4473,N_4323);
nor U7864 (N_7864,N_5195,N_5730);
nor U7865 (N_7865,N_4156,N_5852);
and U7866 (N_7866,N_4211,N_5525);
nand U7867 (N_7867,N_3364,N_5161);
or U7868 (N_7868,N_4434,N_3638);
xor U7869 (N_7869,N_4165,N_3529);
nand U7870 (N_7870,N_4160,N_3897);
nand U7871 (N_7871,N_3259,N_3784);
nand U7872 (N_7872,N_4474,N_3079);
or U7873 (N_7873,N_3301,N_4678);
nand U7874 (N_7874,N_5647,N_4524);
and U7875 (N_7875,N_3176,N_4134);
or U7876 (N_7876,N_4534,N_5214);
nand U7877 (N_7877,N_5815,N_4568);
xnor U7878 (N_7878,N_4410,N_5864);
or U7879 (N_7879,N_4544,N_4841);
or U7880 (N_7880,N_3289,N_5264);
nand U7881 (N_7881,N_5827,N_3166);
xnor U7882 (N_7882,N_4932,N_5063);
nand U7883 (N_7883,N_4283,N_5430);
or U7884 (N_7884,N_5868,N_3011);
nor U7885 (N_7885,N_4983,N_3389);
nor U7886 (N_7886,N_5951,N_3502);
nand U7887 (N_7887,N_5963,N_5433);
or U7888 (N_7888,N_5568,N_4699);
xor U7889 (N_7889,N_4005,N_5699);
xor U7890 (N_7890,N_4702,N_5813);
nand U7891 (N_7891,N_5058,N_4889);
or U7892 (N_7892,N_3154,N_3529);
nor U7893 (N_7893,N_5729,N_5195);
nand U7894 (N_7894,N_3705,N_4436);
nor U7895 (N_7895,N_3197,N_4731);
nor U7896 (N_7896,N_5045,N_5185);
xnor U7897 (N_7897,N_4380,N_4599);
nand U7898 (N_7898,N_5670,N_3156);
nand U7899 (N_7899,N_5230,N_4408);
nor U7900 (N_7900,N_3040,N_4324);
nor U7901 (N_7901,N_3979,N_3948);
nor U7902 (N_7902,N_5933,N_3153);
nand U7903 (N_7903,N_5181,N_3361);
and U7904 (N_7904,N_5420,N_5464);
nand U7905 (N_7905,N_5627,N_3704);
xnor U7906 (N_7906,N_3777,N_3597);
nand U7907 (N_7907,N_5898,N_3754);
nand U7908 (N_7908,N_3316,N_4798);
or U7909 (N_7909,N_3706,N_3590);
xor U7910 (N_7910,N_5206,N_3607);
and U7911 (N_7911,N_5135,N_4966);
nand U7912 (N_7912,N_4315,N_3234);
and U7913 (N_7913,N_4345,N_3369);
and U7914 (N_7914,N_5045,N_5162);
nand U7915 (N_7915,N_5982,N_3610);
nor U7916 (N_7916,N_4220,N_5418);
or U7917 (N_7917,N_4185,N_3530);
nand U7918 (N_7918,N_4257,N_5150);
xor U7919 (N_7919,N_3993,N_4293);
xor U7920 (N_7920,N_5817,N_5603);
nor U7921 (N_7921,N_5777,N_3253);
and U7922 (N_7922,N_3172,N_3028);
xnor U7923 (N_7923,N_4309,N_4911);
and U7924 (N_7924,N_3974,N_3293);
and U7925 (N_7925,N_5065,N_5227);
xor U7926 (N_7926,N_3844,N_3327);
or U7927 (N_7927,N_3431,N_4023);
nor U7928 (N_7928,N_5940,N_3402);
or U7929 (N_7929,N_3251,N_5560);
xor U7930 (N_7930,N_5293,N_3124);
and U7931 (N_7931,N_4419,N_3953);
nand U7932 (N_7932,N_5368,N_5454);
nand U7933 (N_7933,N_4631,N_4114);
xor U7934 (N_7934,N_3319,N_5447);
nor U7935 (N_7935,N_4918,N_4738);
nor U7936 (N_7936,N_4395,N_4956);
xnor U7937 (N_7937,N_5441,N_5078);
or U7938 (N_7938,N_5102,N_5469);
or U7939 (N_7939,N_3800,N_5122);
xnor U7940 (N_7940,N_3907,N_4922);
xor U7941 (N_7941,N_3431,N_5518);
and U7942 (N_7942,N_4168,N_5899);
nor U7943 (N_7943,N_5868,N_4744);
nand U7944 (N_7944,N_3418,N_3061);
or U7945 (N_7945,N_5467,N_5028);
or U7946 (N_7946,N_3455,N_4761);
nor U7947 (N_7947,N_5779,N_4013);
xor U7948 (N_7948,N_5968,N_4098);
nor U7949 (N_7949,N_3632,N_5032);
nand U7950 (N_7950,N_4839,N_5213);
xnor U7951 (N_7951,N_3296,N_3678);
and U7952 (N_7952,N_5051,N_3854);
and U7953 (N_7953,N_4411,N_4496);
nor U7954 (N_7954,N_4003,N_4024);
xnor U7955 (N_7955,N_5961,N_5601);
nand U7956 (N_7956,N_4550,N_3201);
nor U7957 (N_7957,N_4234,N_4224);
xor U7958 (N_7958,N_5893,N_5468);
and U7959 (N_7959,N_4846,N_4786);
nor U7960 (N_7960,N_3269,N_5305);
nor U7961 (N_7961,N_3936,N_3615);
nor U7962 (N_7962,N_4146,N_3340);
and U7963 (N_7963,N_4797,N_3575);
nand U7964 (N_7964,N_4521,N_4736);
or U7965 (N_7965,N_5422,N_4860);
nor U7966 (N_7966,N_3694,N_5798);
and U7967 (N_7967,N_5536,N_5848);
nor U7968 (N_7968,N_3173,N_5479);
and U7969 (N_7969,N_3382,N_3362);
nand U7970 (N_7970,N_3056,N_5299);
and U7971 (N_7971,N_3816,N_5909);
nor U7972 (N_7972,N_4310,N_5524);
xor U7973 (N_7973,N_4289,N_4462);
nand U7974 (N_7974,N_3517,N_5857);
and U7975 (N_7975,N_4288,N_5493);
xor U7976 (N_7976,N_4378,N_4489);
and U7977 (N_7977,N_4230,N_5517);
or U7978 (N_7978,N_5522,N_5919);
xor U7979 (N_7979,N_4001,N_5765);
nand U7980 (N_7980,N_4136,N_5678);
xor U7981 (N_7981,N_5188,N_3626);
xor U7982 (N_7982,N_5358,N_3311);
or U7983 (N_7983,N_3627,N_5721);
nand U7984 (N_7984,N_4654,N_4663);
nor U7985 (N_7985,N_3313,N_4126);
nand U7986 (N_7986,N_3084,N_4323);
nand U7987 (N_7987,N_4486,N_3417);
or U7988 (N_7988,N_4854,N_4220);
or U7989 (N_7989,N_5735,N_3422);
xor U7990 (N_7990,N_4034,N_3345);
nand U7991 (N_7991,N_4762,N_5365);
and U7992 (N_7992,N_3941,N_3815);
and U7993 (N_7993,N_5679,N_3913);
nor U7994 (N_7994,N_5195,N_3623);
nor U7995 (N_7995,N_5979,N_4912);
and U7996 (N_7996,N_4554,N_4935);
or U7997 (N_7997,N_4845,N_4123);
nand U7998 (N_7998,N_3264,N_3566);
xnor U7999 (N_7999,N_3986,N_3136);
and U8000 (N_8000,N_5051,N_4584);
or U8001 (N_8001,N_4858,N_4378);
and U8002 (N_8002,N_3147,N_3425);
nor U8003 (N_8003,N_3966,N_5897);
xnor U8004 (N_8004,N_4180,N_5432);
xnor U8005 (N_8005,N_3385,N_5381);
nand U8006 (N_8006,N_3643,N_3525);
nor U8007 (N_8007,N_3978,N_3653);
xor U8008 (N_8008,N_5342,N_3656);
nor U8009 (N_8009,N_4812,N_3891);
nor U8010 (N_8010,N_3792,N_3890);
xnor U8011 (N_8011,N_4888,N_4308);
nand U8012 (N_8012,N_4382,N_4242);
or U8013 (N_8013,N_4292,N_5333);
or U8014 (N_8014,N_3234,N_3728);
xor U8015 (N_8015,N_5078,N_3773);
and U8016 (N_8016,N_5959,N_4461);
or U8017 (N_8017,N_5407,N_3835);
xor U8018 (N_8018,N_4419,N_3223);
nand U8019 (N_8019,N_5870,N_4766);
or U8020 (N_8020,N_4123,N_3826);
nand U8021 (N_8021,N_4474,N_4994);
nor U8022 (N_8022,N_4234,N_4528);
xnor U8023 (N_8023,N_3342,N_5317);
nand U8024 (N_8024,N_5972,N_3472);
or U8025 (N_8025,N_5920,N_3875);
xnor U8026 (N_8026,N_4464,N_4101);
nor U8027 (N_8027,N_3759,N_3092);
or U8028 (N_8028,N_5088,N_4286);
or U8029 (N_8029,N_3980,N_5314);
xnor U8030 (N_8030,N_3132,N_5874);
nor U8031 (N_8031,N_4326,N_4194);
nor U8032 (N_8032,N_5945,N_3611);
xnor U8033 (N_8033,N_3738,N_3381);
and U8034 (N_8034,N_5414,N_5768);
or U8035 (N_8035,N_5005,N_3102);
and U8036 (N_8036,N_5782,N_3102);
and U8037 (N_8037,N_5421,N_5872);
nand U8038 (N_8038,N_4211,N_5296);
nand U8039 (N_8039,N_5574,N_4996);
nor U8040 (N_8040,N_4024,N_4521);
or U8041 (N_8041,N_5198,N_5430);
nand U8042 (N_8042,N_3805,N_5384);
and U8043 (N_8043,N_4777,N_4726);
and U8044 (N_8044,N_4136,N_5835);
nor U8045 (N_8045,N_4525,N_3930);
or U8046 (N_8046,N_5742,N_4485);
nor U8047 (N_8047,N_4623,N_3582);
xnor U8048 (N_8048,N_4282,N_4691);
and U8049 (N_8049,N_4824,N_5237);
and U8050 (N_8050,N_5500,N_4021);
nor U8051 (N_8051,N_4418,N_3393);
nand U8052 (N_8052,N_5247,N_3115);
xor U8053 (N_8053,N_3405,N_4495);
and U8054 (N_8054,N_3067,N_3848);
xor U8055 (N_8055,N_4627,N_4490);
nand U8056 (N_8056,N_4548,N_5529);
nor U8057 (N_8057,N_4976,N_5093);
nor U8058 (N_8058,N_4699,N_3939);
and U8059 (N_8059,N_3895,N_3706);
xor U8060 (N_8060,N_5693,N_5109);
nand U8061 (N_8061,N_3384,N_4116);
nor U8062 (N_8062,N_3260,N_4687);
and U8063 (N_8063,N_3801,N_5976);
and U8064 (N_8064,N_5174,N_5937);
nor U8065 (N_8065,N_3922,N_3384);
xnor U8066 (N_8066,N_4940,N_4998);
nor U8067 (N_8067,N_5392,N_4694);
and U8068 (N_8068,N_4147,N_5506);
and U8069 (N_8069,N_3661,N_4986);
xnor U8070 (N_8070,N_5501,N_4060);
nand U8071 (N_8071,N_3732,N_5242);
nand U8072 (N_8072,N_4418,N_3280);
nand U8073 (N_8073,N_4461,N_5415);
or U8074 (N_8074,N_4440,N_3483);
xor U8075 (N_8075,N_5111,N_5153);
nor U8076 (N_8076,N_4045,N_3461);
and U8077 (N_8077,N_5142,N_3816);
xnor U8078 (N_8078,N_3137,N_4147);
xnor U8079 (N_8079,N_4148,N_5392);
and U8080 (N_8080,N_3167,N_4440);
nor U8081 (N_8081,N_3299,N_4463);
or U8082 (N_8082,N_5387,N_3191);
nor U8083 (N_8083,N_3268,N_4100);
nand U8084 (N_8084,N_4078,N_3640);
or U8085 (N_8085,N_5510,N_4109);
or U8086 (N_8086,N_4311,N_4270);
xnor U8087 (N_8087,N_5224,N_5160);
and U8088 (N_8088,N_3495,N_4449);
or U8089 (N_8089,N_5756,N_5610);
nand U8090 (N_8090,N_3737,N_4996);
nor U8091 (N_8091,N_5130,N_5940);
and U8092 (N_8092,N_5616,N_5048);
nand U8093 (N_8093,N_3334,N_3340);
or U8094 (N_8094,N_5709,N_3873);
nor U8095 (N_8095,N_4900,N_5976);
and U8096 (N_8096,N_3366,N_3443);
and U8097 (N_8097,N_3414,N_3855);
nand U8098 (N_8098,N_5378,N_3598);
and U8099 (N_8099,N_3262,N_5286);
xnor U8100 (N_8100,N_3381,N_5758);
nand U8101 (N_8101,N_5047,N_3724);
nor U8102 (N_8102,N_5441,N_5891);
or U8103 (N_8103,N_3369,N_4024);
and U8104 (N_8104,N_5280,N_4409);
nand U8105 (N_8105,N_3067,N_3698);
xnor U8106 (N_8106,N_5775,N_5553);
xor U8107 (N_8107,N_4048,N_5715);
and U8108 (N_8108,N_5677,N_3567);
or U8109 (N_8109,N_4380,N_3151);
and U8110 (N_8110,N_4434,N_5926);
xor U8111 (N_8111,N_4291,N_3748);
nor U8112 (N_8112,N_4855,N_4127);
nor U8113 (N_8113,N_3378,N_3902);
and U8114 (N_8114,N_5573,N_3438);
xor U8115 (N_8115,N_4168,N_3865);
nand U8116 (N_8116,N_3036,N_4247);
xor U8117 (N_8117,N_3991,N_5501);
and U8118 (N_8118,N_4287,N_4681);
nor U8119 (N_8119,N_5146,N_5763);
nor U8120 (N_8120,N_3077,N_4496);
and U8121 (N_8121,N_5776,N_3921);
or U8122 (N_8122,N_3584,N_5762);
or U8123 (N_8123,N_4874,N_4510);
or U8124 (N_8124,N_4847,N_5860);
nand U8125 (N_8125,N_4664,N_3988);
nor U8126 (N_8126,N_3947,N_5963);
nand U8127 (N_8127,N_4554,N_5806);
xnor U8128 (N_8128,N_5204,N_5600);
and U8129 (N_8129,N_4703,N_3787);
and U8130 (N_8130,N_3047,N_5672);
nor U8131 (N_8131,N_4072,N_3705);
nand U8132 (N_8132,N_3492,N_4404);
and U8133 (N_8133,N_4257,N_3909);
or U8134 (N_8134,N_3554,N_4515);
or U8135 (N_8135,N_5491,N_4995);
nor U8136 (N_8136,N_5951,N_3361);
nor U8137 (N_8137,N_3652,N_5695);
or U8138 (N_8138,N_4097,N_5338);
xor U8139 (N_8139,N_3770,N_3455);
nor U8140 (N_8140,N_4245,N_5253);
xnor U8141 (N_8141,N_3161,N_4435);
nand U8142 (N_8142,N_5819,N_4353);
xnor U8143 (N_8143,N_4486,N_4213);
nand U8144 (N_8144,N_5572,N_5964);
xor U8145 (N_8145,N_3991,N_3347);
or U8146 (N_8146,N_5385,N_4159);
xor U8147 (N_8147,N_4288,N_5351);
nand U8148 (N_8148,N_4721,N_3335);
or U8149 (N_8149,N_5402,N_3590);
nor U8150 (N_8150,N_4312,N_5547);
nand U8151 (N_8151,N_4959,N_4441);
and U8152 (N_8152,N_5579,N_5016);
xnor U8153 (N_8153,N_4366,N_5804);
and U8154 (N_8154,N_5450,N_5872);
nor U8155 (N_8155,N_5920,N_5896);
nand U8156 (N_8156,N_5084,N_4723);
nand U8157 (N_8157,N_5641,N_5794);
and U8158 (N_8158,N_3535,N_5633);
and U8159 (N_8159,N_3814,N_4571);
nor U8160 (N_8160,N_3991,N_3707);
nand U8161 (N_8161,N_3467,N_3182);
nor U8162 (N_8162,N_5759,N_3849);
nand U8163 (N_8163,N_5321,N_5802);
nor U8164 (N_8164,N_4091,N_5630);
and U8165 (N_8165,N_5264,N_3065);
xor U8166 (N_8166,N_3710,N_4098);
nand U8167 (N_8167,N_5708,N_4286);
nor U8168 (N_8168,N_3287,N_4913);
and U8169 (N_8169,N_4692,N_5362);
and U8170 (N_8170,N_4533,N_3289);
nor U8171 (N_8171,N_3545,N_4995);
or U8172 (N_8172,N_5613,N_3847);
or U8173 (N_8173,N_5927,N_3115);
nand U8174 (N_8174,N_3988,N_3310);
or U8175 (N_8175,N_4199,N_3205);
or U8176 (N_8176,N_4779,N_3508);
nand U8177 (N_8177,N_3822,N_4859);
nand U8178 (N_8178,N_5951,N_3105);
nor U8179 (N_8179,N_5805,N_5547);
xnor U8180 (N_8180,N_4573,N_4423);
or U8181 (N_8181,N_3036,N_3356);
xor U8182 (N_8182,N_5911,N_3795);
nand U8183 (N_8183,N_5917,N_3995);
or U8184 (N_8184,N_3980,N_4260);
and U8185 (N_8185,N_4966,N_4024);
nand U8186 (N_8186,N_3099,N_4390);
or U8187 (N_8187,N_3450,N_5388);
and U8188 (N_8188,N_3550,N_4680);
nand U8189 (N_8189,N_5827,N_4748);
nor U8190 (N_8190,N_5678,N_4823);
nor U8191 (N_8191,N_3589,N_5914);
nor U8192 (N_8192,N_3631,N_5316);
or U8193 (N_8193,N_5103,N_5664);
or U8194 (N_8194,N_3231,N_5318);
xor U8195 (N_8195,N_5221,N_5890);
or U8196 (N_8196,N_5858,N_4219);
nand U8197 (N_8197,N_5985,N_4298);
and U8198 (N_8198,N_3169,N_3185);
xor U8199 (N_8199,N_3872,N_5284);
or U8200 (N_8200,N_3605,N_5035);
xor U8201 (N_8201,N_3158,N_3270);
nor U8202 (N_8202,N_5588,N_5309);
and U8203 (N_8203,N_5732,N_4620);
or U8204 (N_8204,N_4817,N_3851);
or U8205 (N_8205,N_3758,N_3878);
nor U8206 (N_8206,N_3109,N_3240);
nor U8207 (N_8207,N_5056,N_4470);
nand U8208 (N_8208,N_3086,N_4429);
nand U8209 (N_8209,N_3295,N_4483);
nor U8210 (N_8210,N_3735,N_5327);
and U8211 (N_8211,N_3590,N_4372);
nor U8212 (N_8212,N_4011,N_3558);
nand U8213 (N_8213,N_5448,N_3801);
or U8214 (N_8214,N_3617,N_3226);
nand U8215 (N_8215,N_4285,N_3439);
nand U8216 (N_8216,N_5320,N_4321);
nor U8217 (N_8217,N_5700,N_5104);
nand U8218 (N_8218,N_5484,N_3033);
or U8219 (N_8219,N_5102,N_3752);
and U8220 (N_8220,N_5244,N_3706);
xnor U8221 (N_8221,N_4115,N_4620);
nand U8222 (N_8222,N_5013,N_5700);
xnor U8223 (N_8223,N_3224,N_4682);
or U8224 (N_8224,N_3891,N_3498);
xor U8225 (N_8225,N_3513,N_3729);
xnor U8226 (N_8226,N_3712,N_5408);
nand U8227 (N_8227,N_4850,N_5626);
nand U8228 (N_8228,N_5475,N_5910);
and U8229 (N_8229,N_4257,N_4966);
and U8230 (N_8230,N_4266,N_4547);
nor U8231 (N_8231,N_3364,N_4892);
nand U8232 (N_8232,N_4907,N_4426);
nand U8233 (N_8233,N_4935,N_3373);
xor U8234 (N_8234,N_4571,N_5127);
xnor U8235 (N_8235,N_4203,N_5077);
and U8236 (N_8236,N_3794,N_3169);
nand U8237 (N_8237,N_3091,N_5278);
or U8238 (N_8238,N_5330,N_4789);
xor U8239 (N_8239,N_5193,N_4156);
or U8240 (N_8240,N_3577,N_3188);
and U8241 (N_8241,N_5897,N_4539);
nand U8242 (N_8242,N_5139,N_5615);
nand U8243 (N_8243,N_4514,N_5035);
or U8244 (N_8244,N_5709,N_3518);
and U8245 (N_8245,N_5483,N_5322);
xnor U8246 (N_8246,N_5878,N_5371);
nor U8247 (N_8247,N_5670,N_4207);
or U8248 (N_8248,N_5368,N_3999);
xnor U8249 (N_8249,N_3884,N_4146);
or U8250 (N_8250,N_3381,N_4029);
and U8251 (N_8251,N_5160,N_3434);
nor U8252 (N_8252,N_5466,N_3747);
and U8253 (N_8253,N_5215,N_4424);
nand U8254 (N_8254,N_4958,N_4238);
or U8255 (N_8255,N_4438,N_5780);
and U8256 (N_8256,N_5736,N_4042);
and U8257 (N_8257,N_4523,N_5966);
nand U8258 (N_8258,N_5835,N_4803);
xnor U8259 (N_8259,N_4249,N_5926);
or U8260 (N_8260,N_4975,N_5100);
and U8261 (N_8261,N_3798,N_3847);
nand U8262 (N_8262,N_5350,N_5189);
xnor U8263 (N_8263,N_5270,N_4150);
nand U8264 (N_8264,N_5241,N_3560);
xnor U8265 (N_8265,N_4232,N_3983);
xnor U8266 (N_8266,N_5117,N_3473);
or U8267 (N_8267,N_4361,N_3067);
nor U8268 (N_8268,N_4290,N_5035);
or U8269 (N_8269,N_4822,N_4029);
and U8270 (N_8270,N_5672,N_5323);
or U8271 (N_8271,N_4858,N_5208);
xor U8272 (N_8272,N_3366,N_3469);
or U8273 (N_8273,N_3262,N_5395);
xnor U8274 (N_8274,N_3522,N_3750);
xnor U8275 (N_8275,N_3743,N_4071);
and U8276 (N_8276,N_5151,N_5955);
and U8277 (N_8277,N_3643,N_5047);
and U8278 (N_8278,N_5330,N_3114);
xnor U8279 (N_8279,N_3580,N_3721);
xnor U8280 (N_8280,N_5905,N_5419);
and U8281 (N_8281,N_5598,N_4556);
or U8282 (N_8282,N_4156,N_5527);
nor U8283 (N_8283,N_4044,N_4563);
xor U8284 (N_8284,N_5269,N_4567);
or U8285 (N_8285,N_3056,N_4077);
or U8286 (N_8286,N_3267,N_4289);
and U8287 (N_8287,N_4824,N_5830);
nand U8288 (N_8288,N_3372,N_5343);
or U8289 (N_8289,N_3835,N_4029);
nand U8290 (N_8290,N_5602,N_4299);
or U8291 (N_8291,N_4432,N_4381);
or U8292 (N_8292,N_5435,N_5911);
xor U8293 (N_8293,N_5645,N_3929);
xor U8294 (N_8294,N_4484,N_4076);
xor U8295 (N_8295,N_3074,N_5365);
xor U8296 (N_8296,N_4472,N_3499);
and U8297 (N_8297,N_4916,N_3187);
nor U8298 (N_8298,N_5922,N_3555);
xnor U8299 (N_8299,N_4574,N_5020);
nor U8300 (N_8300,N_5296,N_5900);
or U8301 (N_8301,N_4494,N_5489);
or U8302 (N_8302,N_3754,N_3730);
nor U8303 (N_8303,N_4745,N_3915);
and U8304 (N_8304,N_3901,N_4104);
nand U8305 (N_8305,N_4458,N_4453);
xor U8306 (N_8306,N_4624,N_5660);
nand U8307 (N_8307,N_4310,N_5921);
nand U8308 (N_8308,N_4167,N_3690);
nor U8309 (N_8309,N_3886,N_4722);
nand U8310 (N_8310,N_4019,N_3345);
nor U8311 (N_8311,N_4944,N_5511);
xor U8312 (N_8312,N_4326,N_3815);
xor U8313 (N_8313,N_5452,N_3339);
xnor U8314 (N_8314,N_3955,N_4279);
or U8315 (N_8315,N_4455,N_4771);
and U8316 (N_8316,N_4503,N_5434);
or U8317 (N_8317,N_3970,N_3584);
nor U8318 (N_8318,N_4425,N_3649);
xnor U8319 (N_8319,N_4133,N_4710);
nand U8320 (N_8320,N_5781,N_5745);
or U8321 (N_8321,N_5081,N_4532);
xnor U8322 (N_8322,N_3084,N_5438);
nor U8323 (N_8323,N_3789,N_3512);
xnor U8324 (N_8324,N_4532,N_4959);
xnor U8325 (N_8325,N_4519,N_4476);
nor U8326 (N_8326,N_5467,N_4588);
or U8327 (N_8327,N_3432,N_3450);
xnor U8328 (N_8328,N_4528,N_5733);
and U8329 (N_8329,N_5542,N_3715);
nand U8330 (N_8330,N_3175,N_5374);
xor U8331 (N_8331,N_3126,N_5158);
xor U8332 (N_8332,N_5099,N_3989);
and U8333 (N_8333,N_3423,N_3937);
nor U8334 (N_8334,N_5755,N_3555);
nand U8335 (N_8335,N_5757,N_5462);
and U8336 (N_8336,N_5726,N_5175);
or U8337 (N_8337,N_3533,N_5464);
and U8338 (N_8338,N_4701,N_3800);
or U8339 (N_8339,N_4070,N_3163);
nand U8340 (N_8340,N_3022,N_3954);
and U8341 (N_8341,N_3408,N_5441);
and U8342 (N_8342,N_3093,N_3390);
nor U8343 (N_8343,N_3672,N_5187);
and U8344 (N_8344,N_4356,N_4710);
and U8345 (N_8345,N_5979,N_5756);
nand U8346 (N_8346,N_3420,N_4241);
nor U8347 (N_8347,N_5125,N_3615);
nand U8348 (N_8348,N_3059,N_3130);
nor U8349 (N_8349,N_4557,N_5964);
and U8350 (N_8350,N_3497,N_5105);
nand U8351 (N_8351,N_4735,N_5373);
nand U8352 (N_8352,N_4714,N_4629);
nor U8353 (N_8353,N_4265,N_5612);
xor U8354 (N_8354,N_4779,N_3367);
xnor U8355 (N_8355,N_4938,N_3329);
and U8356 (N_8356,N_3464,N_4873);
nor U8357 (N_8357,N_3320,N_3865);
nor U8358 (N_8358,N_5037,N_4172);
and U8359 (N_8359,N_3718,N_5624);
nand U8360 (N_8360,N_3872,N_5888);
nor U8361 (N_8361,N_3139,N_5094);
nor U8362 (N_8362,N_3823,N_5216);
xnor U8363 (N_8363,N_4154,N_4014);
nand U8364 (N_8364,N_3287,N_4539);
xor U8365 (N_8365,N_4256,N_3053);
or U8366 (N_8366,N_4316,N_5120);
xnor U8367 (N_8367,N_3066,N_3802);
xor U8368 (N_8368,N_4335,N_3036);
nand U8369 (N_8369,N_5535,N_5021);
and U8370 (N_8370,N_4417,N_3493);
xnor U8371 (N_8371,N_4038,N_5839);
or U8372 (N_8372,N_5694,N_3031);
or U8373 (N_8373,N_5716,N_5419);
nand U8374 (N_8374,N_4800,N_3779);
or U8375 (N_8375,N_5355,N_4139);
nand U8376 (N_8376,N_5824,N_5908);
nand U8377 (N_8377,N_4802,N_3445);
or U8378 (N_8378,N_3818,N_4787);
nand U8379 (N_8379,N_4418,N_3667);
or U8380 (N_8380,N_5140,N_5038);
xor U8381 (N_8381,N_3835,N_4442);
nand U8382 (N_8382,N_4684,N_4461);
nor U8383 (N_8383,N_5624,N_4439);
or U8384 (N_8384,N_5117,N_3157);
xor U8385 (N_8385,N_3153,N_3184);
and U8386 (N_8386,N_3236,N_4740);
xor U8387 (N_8387,N_3457,N_5797);
and U8388 (N_8388,N_3265,N_4744);
xnor U8389 (N_8389,N_3117,N_5106);
and U8390 (N_8390,N_4210,N_4898);
or U8391 (N_8391,N_4287,N_5434);
xor U8392 (N_8392,N_4592,N_3624);
xor U8393 (N_8393,N_5148,N_4991);
xor U8394 (N_8394,N_5461,N_4627);
and U8395 (N_8395,N_5556,N_3458);
xnor U8396 (N_8396,N_4153,N_4218);
nand U8397 (N_8397,N_4369,N_5393);
nand U8398 (N_8398,N_3979,N_4924);
and U8399 (N_8399,N_5681,N_4790);
or U8400 (N_8400,N_3608,N_3117);
and U8401 (N_8401,N_4547,N_4784);
and U8402 (N_8402,N_3204,N_5664);
nand U8403 (N_8403,N_3057,N_3653);
xnor U8404 (N_8404,N_5529,N_5771);
nor U8405 (N_8405,N_3911,N_3537);
and U8406 (N_8406,N_4781,N_5432);
nand U8407 (N_8407,N_5629,N_3696);
or U8408 (N_8408,N_5176,N_3172);
and U8409 (N_8409,N_3669,N_4298);
xor U8410 (N_8410,N_3648,N_3195);
and U8411 (N_8411,N_3381,N_3006);
and U8412 (N_8412,N_3467,N_4157);
and U8413 (N_8413,N_3955,N_3035);
or U8414 (N_8414,N_5665,N_4459);
nand U8415 (N_8415,N_3798,N_4039);
or U8416 (N_8416,N_5424,N_5602);
or U8417 (N_8417,N_3938,N_4793);
nand U8418 (N_8418,N_5833,N_5566);
nor U8419 (N_8419,N_5210,N_4973);
nand U8420 (N_8420,N_4696,N_4650);
and U8421 (N_8421,N_4937,N_4422);
and U8422 (N_8422,N_3093,N_5907);
and U8423 (N_8423,N_4410,N_5228);
xnor U8424 (N_8424,N_5599,N_3691);
and U8425 (N_8425,N_5423,N_4866);
nor U8426 (N_8426,N_5355,N_5929);
or U8427 (N_8427,N_3808,N_5996);
xor U8428 (N_8428,N_5198,N_3528);
nor U8429 (N_8429,N_5892,N_5878);
or U8430 (N_8430,N_3665,N_5559);
nor U8431 (N_8431,N_3565,N_4626);
and U8432 (N_8432,N_3169,N_4371);
xnor U8433 (N_8433,N_3500,N_5284);
nand U8434 (N_8434,N_4478,N_3898);
nand U8435 (N_8435,N_5117,N_5021);
xor U8436 (N_8436,N_4321,N_3409);
and U8437 (N_8437,N_4703,N_3323);
and U8438 (N_8438,N_5678,N_4596);
and U8439 (N_8439,N_4793,N_5874);
xnor U8440 (N_8440,N_4594,N_5552);
or U8441 (N_8441,N_4141,N_4672);
or U8442 (N_8442,N_3371,N_4659);
and U8443 (N_8443,N_5768,N_3184);
xnor U8444 (N_8444,N_5359,N_5834);
xnor U8445 (N_8445,N_3961,N_4285);
or U8446 (N_8446,N_3651,N_3436);
nand U8447 (N_8447,N_4537,N_3643);
or U8448 (N_8448,N_4839,N_3344);
or U8449 (N_8449,N_4552,N_3115);
nor U8450 (N_8450,N_5360,N_4480);
or U8451 (N_8451,N_5602,N_4177);
and U8452 (N_8452,N_5180,N_4198);
nor U8453 (N_8453,N_3641,N_3486);
or U8454 (N_8454,N_5448,N_4585);
nor U8455 (N_8455,N_4634,N_5385);
or U8456 (N_8456,N_4844,N_3847);
xor U8457 (N_8457,N_5222,N_4837);
xnor U8458 (N_8458,N_4201,N_4635);
or U8459 (N_8459,N_3289,N_4881);
nand U8460 (N_8460,N_3189,N_3717);
nor U8461 (N_8461,N_3128,N_4372);
nand U8462 (N_8462,N_5700,N_3787);
or U8463 (N_8463,N_5019,N_5147);
nor U8464 (N_8464,N_5466,N_3482);
xnor U8465 (N_8465,N_4964,N_3600);
nand U8466 (N_8466,N_4623,N_4644);
xor U8467 (N_8467,N_4968,N_4595);
and U8468 (N_8468,N_4914,N_3291);
and U8469 (N_8469,N_5963,N_3088);
or U8470 (N_8470,N_4102,N_5512);
and U8471 (N_8471,N_3688,N_5740);
nor U8472 (N_8472,N_4325,N_3596);
nor U8473 (N_8473,N_4576,N_3876);
or U8474 (N_8474,N_4455,N_5382);
or U8475 (N_8475,N_3096,N_3881);
or U8476 (N_8476,N_3425,N_5284);
nor U8477 (N_8477,N_3353,N_4573);
nor U8478 (N_8478,N_4564,N_4915);
and U8479 (N_8479,N_4846,N_5863);
nand U8480 (N_8480,N_5076,N_3639);
xnor U8481 (N_8481,N_5872,N_3584);
or U8482 (N_8482,N_3588,N_4755);
nand U8483 (N_8483,N_3884,N_5060);
or U8484 (N_8484,N_3157,N_3996);
and U8485 (N_8485,N_5594,N_5700);
nor U8486 (N_8486,N_3282,N_4010);
or U8487 (N_8487,N_4464,N_4144);
nor U8488 (N_8488,N_3424,N_4713);
nor U8489 (N_8489,N_3491,N_5887);
nor U8490 (N_8490,N_4503,N_5046);
and U8491 (N_8491,N_4012,N_5999);
nor U8492 (N_8492,N_5426,N_5259);
and U8493 (N_8493,N_3801,N_4418);
xnor U8494 (N_8494,N_5882,N_4704);
and U8495 (N_8495,N_5812,N_5075);
xor U8496 (N_8496,N_3924,N_4932);
xnor U8497 (N_8497,N_4218,N_3797);
xnor U8498 (N_8498,N_5045,N_5467);
nand U8499 (N_8499,N_5403,N_4909);
and U8500 (N_8500,N_3358,N_3927);
or U8501 (N_8501,N_4162,N_3143);
nor U8502 (N_8502,N_3845,N_3903);
nor U8503 (N_8503,N_3962,N_5780);
nor U8504 (N_8504,N_5118,N_4089);
and U8505 (N_8505,N_4575,N_5249);
xnor U8506 (N_8506,N_5778,N_4220);
or U8507 (N_8507,N_5606,N_4300);
nor U8508 (N_8508,N_3232,N_3882);
nand U8509 (N_8509,N_4734,N_3034);
and U8510 (N_8510,N_5086,N_4310);
nand U8511 (N_8511,N_5627,N_4250);
and U8512 (N_8512,N_4948,N_3659);
and U8513 (N_8513,N_5302,N_5753);
nand U8514 (N_8514,N_4988,N_5987);
and U8515 (N_8515,N_3531,N_3697);
or U8516 (N_8516,N_5247,N_3532);
nor U8517 (N_8517,N_3822,N_4426);
nand U8518 (N_8518,N_5953,N_3984);
nor U8519 (N_8519,N_5488,N_5295);
nor U8520 (N_8520,N_5036,N_4339);
nor U8521 (N_8521,N_3880,N_3765);
nor U8522 (N_8522,N_3849,N_5608);
or U8523 (N_8523,N_5348,N_5649);
nor U8524 (N_8524,N_3628,N_4699);
nand U8525 (N_8525,N_3766,N_3059);
or U8526 (N_8526,N_5022,N_4864);
nor U8527 (N_8527,N_5580,N_3657);
and U8528 (N_8528,N_4480,N_4066);
or U8529 (N_8529,N_5249,N_3848);
xor U8530 (N_8530,N_4003,N_3168);
or U8531 (N_8531,N_4783,N_5868);
nand U8532 (N_8532,N_3201,N_3071);
nor U8533 (N_8533,N_5063,N_3029);
nand U8534 (N_8534,N_3786,N_5123);
and U8535 (N_8535,N_5126,N_5783);
nand U8536 (N_8536,N_4174,N_5441);
xor U8537 (N_8537,N_5873,N_4811);
nand U8538 (N_8538,N_3940,N_3840);
nand U8539 (N_8539,N_5339,N_5359);
or U8540 (N_8540,N_4400,N_5462);
nor U8541 (N_8541,N_5051,N_3950);
or U8542 (N_8542,N_3263,N_4703);
or U8543 (N_8543,N_4655,N_3939);
or U8544 (N_8544,N_4130,N_5305);
nand U8545 (N_8545,N_4732,N_4138);
and U8546 (N_8546,N_5087,N_4881);
nor U8547 (N_8547,N_5377,N_5374);
or U8548 (N_8548,N_3774,N_5862);
nand U8549 (N_8549,N_4091,N_3111);
xnor U8550 (N_8550,N_4260,N_4534);
xor U8551 (N_8551,N_5839,N_4643);
xor U8552 (N_8552,N_4432,N_4227);
and U8553 (N_8553,N_5208,N_3940);
xnor U8554 (N_8554,N_4935,N_5087);
or U8555 (N_8555,N_5513,N_3555);
and U8556 (N_8556,N_5865,N_3952);
nor U8557 (N_8557,N_4789,N_4526);
and U8558 (N_8558,N_3682,N_3105);
xor U8559 (N_8559,N_4651,N_5661);
or U8560 (N_8560,N_5683,N_3584);
or U8561 (N_8561,N_4652,N_4256);
or U8562 (N_8562,N_4453,N_3109);
nand U8563 (N_8563,N_5697,N_4248);
xnor U8564 (N_8564,N_4020,N_3468);
nand U8565 (N_8565,N_3572,N_5177);
nor U8566 (N_8566,N_5377,N_4589);
and U8567 (N_8567,N_4224,N_4539);
xor U8568 (N_8568,N_3666,N_4274);
nor U8569 (N_8569,N_4169,N_3010);
xnor U8570 (N_8570,N_5408,N_4420);
and U8571 (N_8571,N_4358,N_3795);
nand U8572 (N_8572,N_3769,N_4207);
nor U8573 (N_8573,N_3625,N_3056);
nor U8574 (N_8574,N_3507,N_5827);
and U8575 (N_8575,N_3523,N_3833);
nand U8576 (N_8576,N_4105,N_3161);
xnor U8577 (N_8577,N_3920,N_4593);
and U8578 (N_8578,N_5345,N_5703);
nor U8579 (N_8579,N_5743,N_4829);
and U8580 (N_8580,N_4842,N_3812);
xnor U8581 (N_8581,N_5777,N_3939);
nor U8582 (N_8582,N_5438,N_4487);
nor U8583 (N_8583,N_4687,N_4756);
nand U8584 (N_8584,N_4124,N_4250);
or U8585 (N_8585,N_5312,N_4844);
xnor U8586 (N_8586,N_4727,N_5069);
nand U8587 (N_8587,N_4362,N_4151);
nand U8588 (N_8588,N_5379,N_4127);
nor U8589 (N_8589,N_4248,N_5995);
nor U8590 (N_8590,N_3051,N_3810);
or U8591 (N_8591,N_5135,N_5151);
nand U8592 (N_8592,N_3470,N_3950);
or U8593 (N_8593,N_4412,N_5309);
or U8594 (N_8594,N_5892,N_4322);
nand U8595 (N_8595,N_3636,N_3841);
nor U8596 (N_8596,N_3049,N_4203);
or U8597 (N_8597,N_4247,N_3121);
and U8598 (N_8598,N_5740,N_5951);
nor U8599 (N_8599,N_3837,N_3746);
nor U8600 (N_8600,N_4328,N_4382);
xor U8601 (N_8601,N_3883,N_3421);
and U8602 (N_8602,N_3323,N_4236);
nand U8603 (N_8603,N_4164,N_5648);
and U8604 (N_8604,N_3132,N_3911);
or U8605 (N_8605,N_4923,N_4494);
xor U8606 (N_8606,N_5033,N_4310);
nand U8607 (N_8607,N_4614,N_5511);
nor U8608 (N_8608,N_5650,N_3316);
and U8609 (N_8609,N_5253,N_4401);
nor U8610 (N_8610,N_4987,N_5420);
nor U8611 (N_8611,N_5033,N_3777);
or U8612 (N_8612,N_4297,N_5715);
nor U8613 (N_8613,N_3614,N_5290);
nand U8614 (N_8614,N_5008,N_5577);
nand U8615 (N_8615,N_3448,N_3415);
xor U8616 (N_8616,N_5495,N_4664);
nand U8617 (N_8617,N_4412,N_5464);
or U8618 (N_8618,N_4927,N_3647);
nor U8619 (N_8619,N_5301,N_3165);
or U8620 (N_8620,N_5449,N_4450);
and U8621 (N_8621,N_3710,N_5360);
nor U8622 (N_8622,N_3398,N_4468);
nor U8623 (N_8623,N_4797,N_5153);
xnor U8624 (N_8624,N_3172,N_3856);
nor U8625 (N_8625,N_3376,N_4226);
or U8626 (N_8626,N_5218,N_3974);
xor U8627 (N_8627,N_5180,N_4707);
xnor U8628 (N_8628,N_4730,N_5291);
and U8629 (N_8629,N_4921,N_4866);
and U8630 (N_8630,N_4168,N_4665);
xnor U8631 (N_8631,N_3838,N_5839);
or U8632 (N_8632,N_5601,N_5509);
or U8633 (N_8633,N_5838,N_3927);
nand U8634 (N_8634,N_4651,N_5709);
nand U8635 (N_8635,N_3275,N_4324);
nor U8636 (N_8636,N_4376,N_5198);
nor U8637 (N_8637,N_4787,N_3114);
and U8638 (N_8638,N_3032,N_4193);
nor U8639 (N_8639,N_3049,N_4721);
nor U8640 (N_8640,N_3715,N_3039);
or U8641 (N_8641,N_5295,N_5710);
nand U8642 (N_8642,N_4335,N_3900);
or U8643 (N_8643,N_3447,N_4213);
and U8644 (N_8644,N_3653,N_4089);
or U8645 (N_8645,N_3978,N_4680);
nor U8646 (N_8646,N_3483,N_5288);
and U8647 (N_8647,N_4804,N_5827);
xor U8648 (N_8648,N_5342,N_5274);
nand U8649 (N_8649,N_5847,N_5732);
or U8650 (N_8650,N_4082,N_4639);
xnor U8651 (N_8651,N_4259,N_4274);
and U8652 (N_8652,N_3104,N_5118);
nand U8653 (N_8653,N_4458,N_4699);
and U8654 (N_8654,N_3463,N_5509);
nor U8655 (N_8655,N_4705,N_5783);
xnor U8656 (N_8656,N_3231,N_3566);
nand U8657 (N_8657,N_5285,N_4141);
and U8658 (N_8658,N_4931,N_5263);
xor U8659 (N_8659,N_4343,N_3279);
and U8660 (N_8660,N_5477,N_3645);
nand U8661 (N_8661,N_4005,N_3693);
nor U8662 (N_8662,N_4403,N_3904);
nand U8663 (N_8663,N_4183,N_4509);
and U8664 (N_8664,N_5510,N_4116);
and U8665 (N_8665,N_5882,N_4591);
or U8666 (N_8666,N_3392,N_4928);
nand U8667 (N_8667,N_3421,N_3808);
nor U8668 (N_8668,N_4462,N_5718);
nor U8669 (N_8669,N_4405,N_3266);
and U8670 (N_8670,N_3704,N_4035);
or U8671 (N_8671,N_3835,N_4875);
or U8672 (N_8672,N_4816,N_5473);
and U8673 (N_8673,N_5678,N_4664);
nor U8674 (N_8674,N_4217,N_5231);
or U8675 (N_8675,N_3281,N_3110);
nor U8676 (N_8676,N_5743,N_3332);
nor U8677 (N_8677,N_5526,N_4907);
and U8678 (N_8678,N_3651,N_4793);
or U8679 (N_8679,N_3382,N_3676);
and U8680 (N_8680,N_4859,N_5128);
nand U8681 (N_8681,N_3730,N_3183);
or U8682 (N_8682,N_4574,N_5342);
nand U8683 (N_8683,N_3569,N_4324);
and U8684 (N_8684,N_5256,N_5831);
nand U8685 (N_8685,N_5944,N_4115);
xnor U8686 (N_8686,N_3314,N_4453);
and U8687 (N_8687,N_5457,N_4178);
and U8688 (N_8688,N_3681,N_5531);
or U8689 (N_8689,N_5924,N_4756);
and U8690 (N_8690,N_3787,N_4857);
xnor U8691 (N_8691,N_3760,N_5739);
nor U8692 (N_8692,N_3466,N_3653);
nand U8693 (N_8693,N_3204,N_4168);
nor U8694 (N_8694,N_4139,N_3636);
xnor U8695 (N_8695,N_4116,N_4777);
nor U8696 (N_8696,N_4420,N_5356);
nor U8697 (N_8697,N_5708,N_5883);
or U8698 (N_8698,N_5239,N_3178);
and U8699 (N_8699,N_5146,N_3875);
xor U8700 (N_8700,N_4707,N_4143);
and U8701 (N_8701,N_4981,N_5013);
nand U8702 (N_8702,N_3045,N_5658);
nor U8703 (N_8703,N_3648,N_3652);
or U8704 (N_8704,N_4292,N_3226);
nand U8705 (N_8705,N_5074,N_4982);
or U8706 (N_8706,N_5592,N_5048);
or U8707 (N_8707,N_4382,N_3854);
nor U8708 (N_8708,N_4477,N_4205);
or U8709 (N_8709,N_4341,N_3476);
xor U8710 (N_8710,N_4437,N_3136);
or U8711 (N_8711,N_4451,N_3966);
nand U8712 (N_8712,N_4943,N_4948);
xnor U8713 (N_8713,N_3079,N_4299);
nor U8714 (N_8714,N_5132,N_5864);
nor U8715 (N_8715,N_4296,N_5231);
nand U8716 (N_8716,N_4105,N_4863);
xor U8717 (N_8717,N_4709,N_4855);
or U8718 (N_8718,N_4681,N_4390);
xnor U8719 (N_8719,N_4953,N_4307);
and U8720 (N_8720,N_5938,N_5199);
or U8721 (N_8721,N_4831,N_5909);
xor U8722 (N_8722,N_5943,N_4201);
or U8723 (N_8723,N_3719,N_5152);
or U8724 (N_8724,N_5121,N_5160);
nand U8725 (N_8725,N_5009,N_3658);
xnor U8726 (N_8726,N_5967,N_5959);
and U8727 (N_8727,N_5233,N_4564);
or U8728 (N_8728,N_3153,N_5017);
nand U8729 (N_8729,N_4130,N_3559);
xnor U8730 (N_8730,N_3151,N_5217);
nor U8731 (N_8731,N_4662,N_4611);
or U8732 (N_8732,N_5154,N_4413);
nand U8733 (N_8733,N_4851,N_5877);
or U8734 (N_8734,N_5592,N_4191);
xor U8735 (N_8735,N_3995,N_4867);
xnor U8736 (N_8736,N_5594,N_5680);
or U8737 (N_8737,N_4228,N_3974);
nand U8738 (N_8738,N_4097,N_3108);
xnor U8739 (N_8739,N_5576,N_4869);
xor U8740 (N_8740,N_4699,N_4658);
nor U8741 (N_8741,N_4622,N_3457);
and U8742 (N_8742,N_3684,N_4974);
nand U8743 (N_8743,N_4144,N_5692);
or U8744 (N_8744,N_3773,N_3711);
nand U8745 (N_8745,N_4983,N_5198);
nor U8746 (N_8746,N_5521,N_3202);
and U8747 (N_8747,N_5308,N_4862);
xor U8748 (N_8748,N_3352,N_4874);
nor U8749 (N_8749,N_4551,N_5505);
xor U8750 (N_8750,N_5837,N_3419);
xnor U8751 (N_8751,N_4493,N_3016);
or U8752 (N_8752,N_5629,N_4928);
and U8753 (N_8753,N_5796,N_3253);
nor U8754 (N_8754,N_4586,N_5165);
and U8755 (N_8755,N_4752,N_3808);
nor U8756 (N_8756,N_5008,N_4021);
and U8757 (N_8757,N_5331,N_3668);
or U8758 (N_8758,N_3771,N_4955);
nor U8759 (N_8759,N_3401,N_3969);
nand U8760 (N_8760,N_4879,N_5700);
and U8761 (N_8761,N_5644,N_3157);
xor U8762 (N_8762,N_4759,N_4940);
xor U8763 (N_8763,N_3401,N_4784);
nor U8764 (N_8764,N_4209,N_3752);
nor U8765 (N_8765,N_4786,N_5017);
xnor U8766 (N_8766,N_5902,N_3277);
nand U8767 (N_8767,N_5065,N_3849);
xnor U8768 (N_8768,N_3737,N_5164);
nor U8769 (N_8769,N_3225,N_4876);
nor U8770 (N_8770,N_4416,N_5884);
and U8771 (N_8771,N_4506,N_5856);
xnor U8772 (N_8772,N_4192,N_4237);
nand U8773 (N_8773,N_3169,N_5843);
or U8774 (N_8774,N_3548,N_3948);
nand U8775 (N_8775,N_4394,N_5494);
and U8776 (N_8776,N_5960,N_3932);
nand U8777 (N_8777,N_5127,N_5317);
and U8778 (N_8778,N_3181,N_5698);
xnor U8779 (N_8779,N_3701,N_3891);
nor U8780 (N_8780,N_3931,N_4556);
xor U8781 (N_8781,N_4661,N_4104);
nor U8782 (N_8782,N_4678,N_4513);
or U8783 (N_8783,N_4004,N_3842);
and U8784 (N_8784,N_3476,N_5298);
nand U8785 (N_8785,N_4932,N_3121);
and U8786 (N_8786,N_3961,N_3922);
nor U8787 (N_8787,N_4405,N_3861);
xor U8788 (N_8788,N_5653,N_5776);
and U8789 (N_8789,N_3582,N_3614);
xnor U8790 (N_8790,N_3057,N_4970);
or U8791 (N_8791,N_3190,N_4907);
xor U8792 (N_8792,N_5133,N_5046);
xor U8793 (N_8793,N_4132,N_4171);
nor U8794 (N_8794,N_3057,N_5483);
nor U8795 (N_8795,N_4225,N_3036);
or U8796 (N_8796,N_5037,N_5504);
xor U8797 (N_8797,N_3641,N_4289);
and U8798 (N_8798,N_3940,N_3132);
and U8799 (N_8799,N_4488,N_5382);
nor U8800 (N_8800,N_3372,N_5582);
xor U8801 (N_8801,N_4176,N_5394);
or U8802 (N_8802,N_4425,N_4771);
xnor U8803 (N_8803,N_5826,N_3498);
and U8804 (N_8804,N_4645,N_5248);
and U8805 (N_8805,N_5404,N_5495);
nor U8806 (N_8806,N_5375,N_4672);
and U8807 (N_8807,N_4212,N_4204);
and U8808 (N_8808,N_5393,N_4725);
xor U8809 (N_8809,N_5478,N_3667);
xnor U8810 (N_8810,N_4086,N_5694);
and U8811 (N_8811,N_3943,N_5823);
xnor U8812 (N_8812,N_3923,N_4244);
xor U8813 (N_8813,N_5786,N_4533);
nand U8814 (N_8814,N_5300,N_3314);
xnor U8815 (N_8815,N_5781,N_4951);
or U8816 (N_8816,N_4299,N_3180);
xor U8817 (N_8817,N_4590,N_4230);
nand U8818 (N_8818,N_5145,N_3397);
xnor U8819 (N_8819,N_4389,N_5948);
nand U8820 (N_8820,N_3623,N_3252);
xnor U8821 (N_8821,N_3314,N_4444);
and U8822 (N_8822,N_3040,N_4222);
nor U8823 (N_8823,N_3620,N_3792);
or U8824 (N_8824,N_4693,N_4618);
or U8825 (N_8825,N_5185,N_4256);
nand U8826 (N_8826,N_3880,N_5242);
or U8827 (N_8827,N_5580,N_5904);
nand U8828 (N_8828,N_4980,N_3513);
and U8829 (N_8829,N_4394,N_3885);
nand U8830 (N_8830,N_5084,N_5378);
nand U8831 (N_8831,N_4424,N_4041);
xnor U8832 (N_8832,N_5472,N_3008);
or U8833 (N_8833,N_3268,N_3688);
xnor U8834 (N_8834,N_5577,N_3162);
nor U8835 (N_8835,N_4948,N_4429);
nand U8836 (N_8836,N_5803,N_5124);
or U8837 (N_8837,N_4004,N_4645);
nor U8838 (N_8838,N_4249,N_3308);
or U8839 (N_8839,N_3643,N_4749);
xnor U8840 (N_8840,N_4999,N_5531);
nor U8841 (N_8841,N_4053,N_4282);
nor U8842 (N_8842,N_5274,N_3669);
xor U8843 (N_8843,N_4172,N_5156);
and U8844 (N_8844,N_5571,N_4170);
nor U8845 (N_8845,N_5535,N_4461);
xor U8846 (N_8846,N_3204,N_5952);
nand U8847 (N_8847,N_3250,N_3950);
nand U8848 (N_8848,N_3858,N_4006);
nand U8849 (N_8849,N_4921,N_4797);
xnor U8850 (N_8850,N_3132,N_3458);
and U8851 (N_8851,N_4705,N_5992);
nand U8852 (N_8852,N_5390,N_5026);
nor U8853 (N_8853,N_3465,N_3610);
or U8854 (N_8854,N_4478,N_3883);
nand U8855 (N_8855,N_4336,N_4003);
nand U8856 (N_8856,N_3928,N_3059);
nand U8857 (N_8857,N_3978,N_3043);
xor U8858 (N_8858,N_5430,N_5443);
nand U8859 (N_8859,N_4154,N_4056);
or U8860 (N_8860,N_3009,N_5654);
and U8861 (N_8861,N_4484,N_4434);
and U8862 (N_8862,N_3394,N_4701);
nor U8863 (N_8863,N_3661,N_4902);
nand U8864 (N_8864,N_3020,N_3291);
or U8865 (N_8865,N_4556,N_4603);
or U8866 (N_8866,N_5837,N_5097);
and U8867 (N_8867,N_3116,N_3281);
nand U8868 (N_8868,N_5877,N_4575);
xor U8869 (N_8869,N_3338,N_4113);
and U8870 (N_8870,N_5999,N_3620);
nand U8871 (N_8871,N_3946,N_4463);
xor U8872 (N_8872,N_4090,N_5976);
xnor U8873 (N_8873,N_3526,N_4989);
or U8874 (N_8874,N_5428,N_3601);
nand U8875 (N_8875,N_3123,N_3309);
xnor U8876 (N_8876,N_4980,N_3665);
nor U8877 (N_8877,N_5071,N_4942);
and U8878 (N_8878,N_4039,N_5532);
or U8879 (N_8879,N_5783,N_5712);
xor U8880 (N_8880,N_5861,N_4031);
nand U8881 (N_8881,N_3728,N_5914);
xor U8882 (N_8882,N_4170,N_3820);
xor U8883 (N_8883,N_3405,N_5980);
nor U8884 (N_8884,N_3592,N_4064);
xor U8885 (N_8885,N_5620,N_5342);
xnor U8886 (N_8886,N_5553,N_3494);
xnor U8887 (N_8887,N_3234,N_4299);
or U8888 (N_8888,N_5745,N_3217);
xor U8889 (N_8889,N_4887,N_4513);
nand U8890 (N_8890,N_5334,N_4433);
and U8891 (N_8891,N_5935,N_5404);
and U8892 (N_8892,N_3867,N_3147);
nor U8893 (N_8893,N_3438,N_4338);
and U8894 (N_8894,N_4598,N_4981);
nand U8895 (N_8895,N_5686,N_4900);
or U8896 (N_8896,N_3523,N_4444);
or U8897 (N_8897,N_4516,N_4818);
xnor U8898 (N_8898,N_4434,N_3073);
xnor U8899 (N_8899,N_4604,N_4497);
and U8900 (N_8900,N_4773,N_3849);
xor U8901 (N_8901,N_3701,N_5748);
or U8902 (N_8902,N_4663,N_4470);
and U8903 (N_8903,N_5557,N_4545);
or U8904 (N_8904,N_3770,N_4572);
and U8905 (N_8905,N_3671,N_5367);
xor U8906 (N_8906,N_4189,N_4163);
or U8907 (N_8907,N_3351,N_4032);
nor U8908 (N_8908,N_5111,N_5739);
nor U8909 (N_8909,N_3386,N_3389);
xor U8910 (N_8910,N_3502,N_3049);
and U8911 (N_8911,N_4233,N_5952);
nor U8912 (N_8912,N_3212,N_4340);
and U8913 (N_8913,N_5326,N_5216);
or U8914 (N_8914,N_4252,N_5441);
nand U8915 (N_8915,N_3767,N_3861);
nor U8916 (N_8916,N_5105,N_5035);
nand U8917 (N_8917,N_3922,N_4808);
and U8918 (N_8918,N_4447,N_5359);
nor U8919 (N_8919,N_4389,N_5147);
and U8920 (N_8920,N_5888,N_5023);
xnor U8921 (N_8921,N_3396,N_5983);
or U8922 (N_8922,N_3947,N_5400);
and U8923 (N_8923,N_3926,N_5965);
or U8924 (N_8924,N_4906,N_3263);
or U8925 (N_8925,N_3990,N_5150);
nor U8926 (N_8926,N_5409,N_4922);
and U8927 (N_8927,N_3092,N_5316);
and U8928 (N_8928,N_3066,N_5008);
and U8929 (N_8929,N_4991,N_4109);
or U8930 (N_8930,N_5930,N_5008);
xor U8931 (N_8931,N_4025,N_3645);
nand U8932 (N_8932,N_5866,N_3081);
or U8933 (N_8933,N_3382,N_5425);
nor U8934 (N_8934,N_4616,N_4889);
xor U8935 (N_8935,N_3098,N_3976);
and U8936 (N_8936,N_3360,N_5349);
or U8937 (N_8937,N_5885,N_3308);
or U8938 (N_8938,N_4097,N_5027);
nand U8939 (N_8939,N_5939,N_4024);
nand U8940 (N_8940,N_4718,N_5321);
or U8941 (N_8941,N_5328,N_5552);
nor U8942 (N_8942,N_5968,N_4838);
nor U8943 (N_8943,N_3408,N_5116);
nand U8944 (N_8944,N_3597,N_5768);
or U8945 (N_8945,N_5337,N_4713);
xnor U8946 (N_8946,N_5075,N_5691);
nor U8947 (N_8947,N_4961,N_3217);
and U8948 (N_8948,N_5583,N_3768);
xnor U8949 (N_8949,N_5328,N_5085);
or U8950 (N_8950,N_4485,N_3138);
nor U8951 (N_8951,N_4010,N_3153);
xor U8952 (N_8952,N_3168,N_5332);
and U8953 (N_8953,N_3974,N_3107);
or U8954 (N_8954,N_4236,N_3774);
or U8955 (N_8955,N_5606,N_3697);
nor U8956 (N_8956,N_4264,N_5868);
nor U8957 (N_8957,N_4992,N_5951);
xnor U8958 (N_8958,N_5689,N_3279);
nor U8959 (N_8959,N_5879,N_4778);
nor U8960 (N_8960,N_5498,N_4566);
nor U8961 (N_8961,N_3327,N_5249);
xor U8962 (N_8962,N_5340,N_5494);
xnor U8963 (N_8963,N_3277,N_3411);
and U8964 (N_8964,N_5847,N_4962);
nor U8965 (N_8965,N_4113,N_3511);
nand U8966 (N_8966,N_4733,N_5213);
nor U8967 (N_8967,N_4374,N_3372);
or U8968 (N_8968,N_4004,N_5333);
nand U8969 (N_8969,N_3387,N_4965);
or U8970 (N_8970,N_5211,N_4391);
nand U8971 (N_8971,N_5072,N_3598);
xor U8972 (N_8972,N_3960,N_3782);
and U8973 (N_8973,N_4659,N_4609);
and U8974 (N_8974,N_3810,N_5729);
nor U8975 (N_8975,N_4995,N_4639);
and U8976 (N_8976,N_5543,N_4235);
nor U8977 (N_8977,N_5778,N_4564);
xor U8978 (N_8978,N_5031,N_5056);
nor U8979 (N_8979,N_3042,N_3753);
nor U8980 (N_8980,N_3396,N_5328);
nand U8981 (N_8981,N_5466,N_5330);
and U8982 (N_8982,N_5642,N_4059);
xor U8983 (N_8983,N_5384,N_4568);
nor U8984 (N_8984,N_5739,N_3192);
or U8985 (N_8985,N_5173,N_5476);
or U8986 (N_8986,N_5683,N_4694);
nor U8987 (N_8987,N_4529,N_3630);
xor U8988 (N_8988,N_4661,N_5948);
nor U8989 (N_8989,N_5884,N_5504);
or U8990 (N_8990,N_3358,N_5995);
or U8991 (N_8991,N_5134,N_3683);
or U8992 (N_8992,N_3243,N_4093);
or U8993 (N_8993,N_5271,N_5295);
xnor U8994 (N_8994,N_4166,N_5525);
nor U8995 (N_8995,N_5329,N_4223);
nand U8996 (N_8996,N_4555,N_3455);
xor U8997 (N_8997,N_5262,N_4749);
xnor U8998 (N_8998,N_5014,N_4317);
nand U8999 (N_8999,N_5027,N_5784);
and U9000 (N_9000,N_7062,N_8975);
nor U9001 (N_9001,N_7740,N_8278);
nor U9002 (N_9002,N_7965,N_8045);
xor U9003 (N_9003,N_8643,N_6238);
or U9004 (N_9004,N_7106,N_6413);
and U9005 (N_9005,N_7754,N_7750);
and U9006 (N_9006,N_8938,N_6407);
nor U9007 (N_9007,N_7635,N_8583);
nor U9008 (N_9008,N_6914,N_8714);
and U9009 (N_9009,N_6030,N_7813);
nand U9010 (N_9010,N_7476,N_7382);
or U9011 (N_9011,N_8561,N_8759);
xor U9012 (N_9012,N_6174,N_6033);
and U9013 (N_9013,N_6760,N_6027);
and U9014 (N_9014,N_8372,N_7160);
nand U9015 (N_9015,N_8517,N_7996);
or U9016 (N_9016,N_6474,N_7795);
and U9017 (N_9017,N_8052,N_6843);
or U9018 (N_9018,N_8082,N_6781);
or U9019 (N_9019,N_7568,N_7920);
xor U9020 (N_9020,N_6092,N_6081);
xor U9021 (N_9021,N_7640,N_8369);
xor U9022 (N_9022,N_6619,N_7811);
nand U9023 (N_9023,N_7064,N_8460);
xor U9024 (N_9024,N_6734,N_7712);
xor U9025 (N_9025,N_8337,N_7852);
and U9026 (N_9026,N_8622,N_7487);
and U9027 (N_9027,N_6193,N_8926);
nor U9028 (N_9028,N_6920,N_7680);
nor U9029 (N_9029,N_8654,N_7542);
xnor U9030 (N_9030,N_7053,N_6487);
nor U9031 (N_9031,N_7516,N_6875);
nand U9032 (N_9032,N_7224,N_7482);
nand U9033 (N_9033,N_7277,N_7925);
nand U9034 (N_9034,N_6683,N_8784);
nor U9035 (N_9035,N_6803,N_7551);
nor U9036 (N_9036,N_7211,N_8144);
and U9037 (N_9037,N_6661,N_7467);
and U9038 (N_9038,N_8010,N_6333);
or U9039 (N_9039,N_8172,N_7851);
nor U9040 (N_9040,N_8981,N_6695);
nand U9041 (N_9041,N_8685,N_7818);
and U9042 (N_9042,N_6464,N_6204);
nor U9043 (N_9043,N_6365,N_6391);
nor U9044 (N_9044,N_7956,N_8693);
nor U9045 (N_9045,N_7961,N_7981);
nor U9046 (N_9046,N_6186,N_6498);
nand U9047 (N_9047,N_8691,N_6199);
xor U9048 (N_9048,N_7258,N_6806);
xor U9049 (N_9049,N_8856,N_6783);
xor U9050 (N_9050,N_7819,N_6115);
or U9051 (N_9051,N_8909,N_8336);
and U9052 (N_9052,N_8824,N_6007);
xor U9053 (N_9053,N_8785,N_6080);
nor U9054 (N_9054,N_6521,N_8702);
or U9055 (N_9055,N_6577,N_7168);
or U9056 (N_9056,N_8948,N_6928);
or U9057 (N_9057,N_6877,N_7355);
and U9058 (N_9058,N_7520,N_8835);
xor U9059 (N_9059,N_8295,N_8412);
and U9060 (N_9060,N_7278,N_6542);
and U9061 (N_9061,N_7580,N_6026);
nand U9062 (N_9062,N_8068,N_6627);
xor U9063 (N_9063,N_7471,N_6158);
xor U9064 (N_9064,N_8611,N_7773);
or U9065 (N_9065,N_8263,N_8904);
or U9066 (N_9066,N_6794,N_7182);
nand U9067 (N_9067,N_8722,N_7664);
and U9068 (N_9068,N_7723,N_7215);
nand U9069 (N_9069,N_8379,N_7026);
nor U9070 (N_9070,N_8270,N_6880);
nor U9071 (N_9071,N_6378,N_6576);
or U9072 (N_9072,N_6190,N_8145);
nor U9073 (N_9073,N_7112,N_7216);
xor U9074 (N_9074,N_6500,N_7140);
or U9075 (N_9075,N_8020,N_7218);
or U9076 (N_9076,N_8380,N_8871);
and U9077 (N_9077,N_8576,N_7674);
nand U9078 (N_9078,N_8457,N_8456);
nor U9079 (N_9079,N_8589,N_7364);
and U9080 (N_9080,N_6131,N_7016);
and U9081 (N_9081,N_8647,N_6573);
or U9082 (N_9082,N_7759,N_8138);
or U9083 (N_9083,N_8772,N_6923);
xor U9084 (N_9084,N_7625,N_8445);
or U9085 (N_9085,N_8406,N_8775);
or U9086 (N_9086,N_6939,N_8916);
xnor U9087 (N_9087,N_8868,N_6927);
xor U9088 (N_9088,N_7057,N_7189);
and U9089 (N_9089,N_6485,N_8829);
xor U9090 (N_9090,N_6738,N_6802);
nor U9091 (N_9091,N_6956,N_8294);
or U9092 (N_9092,N_8653,N_8448);
nor U9093 (N_9093,N_6670,N_7890);
xnor U9094 (N_9094,N_7812,N_8619);
or U9095 (N_9095,N_7830,N_7008);
and U9096 (N_9096,N_6699,N_6947);
and U9097 (N_9097,N_7343,N_7919);
xor U9098 (N_9098,N_6623,N_6785);
xnor U9099 (N_9099,N_6144,N_7496);
nand U9100 (N_9100,N_6646,N_8204);
nand U9101 (N_9101,N_6171,N_6967);
xor U9102 (N_9102,N_6713,N_8341);
or U9103 (N_9103,N_8723,N_7300);
nand U9104 (N_9104,N_6506,N_8164);
or U9105 (N_9105,N_7308,N_8587);
and U9106 (N_9106,N_8849,N_6096);
nor U9107 (N_9107,N_7582,N_6860);
xnor U9108 (N_9108,N_7173,N_7119);
xor U9109 (N_9109,N_8115,N_6814);
nand U9110 (N_9110,N_7775,N_6099);
and U9111 (N_9111,N_6987,N_7589);
xnor U9112 (N_9112,N_7823,N_8519);
or U9113 (N_9113,N_6183,N_6167);
nor U9114 (N_9114,N_7510,N_6525);
nand U9115 (N_9115,N_8347,N_6331);
nand U9116 (N_9116,N_6435,N_7362);
nor U9117 (N_9117,N_7421,N_6882);
or U9118 (N_9118,N_6979,N_7997);
or U9119 (N_9119,N_7495,N_7720);
or U9120 (N_9120,N_8079,N_7011);
xor U9121 (N_9121,N_7394,N_7672);
or U9122 (N_9122,N_6700,N_8421);
nand U9123 (N_9123,N_8348,N_7989);
xnor U9124 (N_9124,N_7730,N_8839);
nand U9125 (N_9125,N_6971,N_8745);
nand U9126 (N_9126,N_6237,N_7484);
xor U9127 (N_9127,N_7452,N_7135);
and U9128 (N_9128,N_6426,N_7100);
nor U9129 (N_9129,N_6303,N_6547);
nor U9130 (N_9130,N_7833,N_7096);
nand U9131 (N_9131,N_6399,N_7425);
xor U9132 (N_9132,N_6757,N_8301);
and U9133 (N_9133,N_6447,N_6504);
or U9134 (N_9134,N_7456,N_8292);
nand U9135 (N_9135,N_6930,N_8417);
and U9136 (N_9136,N_6278,N_6041);
xnor U9137 (N_9137,N_8955,N_6352);
and U9138 (N_9138,N_6336,N_6643);
or U9139 (N_9139,N_8930,N_8530);
and U9140 (N_9140,N_8770,N_6872);
or U9141 (N_9141,N_6664,N_6489);
xnor U9142 (N_9142,N_6091,N_6126);
nand U9143 (N_9143,N_8252,N_7419);
xnor U9144 (N_9144,N_6600,N_7637);
nor U9145 (N_9145,N_7251,N_6034);
nand U9146 (N_9146,N_6090,N_6173);
xnor U9147 (N_9147,N_6924,N_8766);
xor U9148 (N_9148,N_7760,N_7679);
nand U9149 (N_9149,N_6793,N_6773);
and U9150 (N_9150,N_7587,N_8593);
and U9151 (N_9151,N_7172,N_8166);
or U9152 (N_9152,N_7318,N_7017);
or U9153 (N_9153,N_7791,N_8672);
nand U9154 (N_9154,N_6040,N_6739);
nand U9155 (N_9155,N_8580,N_8738);
nor U9156 (N_9156,N_8044,N_6827);
or U9157 (N_9157,N_6214,N_6082);
xnor U9158 (N_9158,N_8487,N_8936);
xor U9159 (N_9159,N_6554,N_6480);
nor U9160 (N_9160,N_6772,N_7843);
xnor U9161 (N_9161,N_6286,N_7237);
or U9162 (N_9162,N_8754,N_8933);
nor U9163 (N_9163,N_8330,N_6965);
nor U9164 (N_9164,N_7719,N_6259);
xor U9165 (N_9165,N_7121,N_6270);
xor U9166 (N_9166,N_7409,N_6644);
and U9167 (N_9167,N_7081,N_7039);
nand U9168 (N_9168,N_7878,N_7884);
or U9169 (N_9169,N_8016,N_7904);
and U9170 (N_9170,N_7391,N_7264);
nor U9171 (N_9171,N_8721,N_7461);
nand U9172 (N_9172,N_6808,N_7731);
nand U9173 (N_9173,N_7560,N_8744);
and U9174 (N_9174,N_6049,N_6654);
xnor U9175 (N_9175,N_7486,N_8377);
and U9176 (N_9176,N_7979,N_6380);
nand U9177 (N_9177,N_8275,N_6166);
nand U9178 (N_9178,N_7359,N_8817);
or U9179 (N_9179,N_7835,N_8283);
and U9180 (N_9180,N_7814,N_8494);
or U9181 (N_9181,N_7159,N_8351);
nand U9182 (N_9182,N_6220,N_6114);
xor U9183 (N_9183,N_8842,N_8409);
and U9184 (N_9184,N_8137,N_6208);
nor U9185 (N_9185,N_8780,N_6453);
and U9186 (N_9186,N_8710,N_6909);
and U9187 (N_9187,N_6377,N_8514);
and U9188 (N_9188,N_7195,N_6146);
nor U9189 (N_9189,N_6598,N_6659);
xnor U9190 (N_9190,N_6574,N_6261);
and U9191 (N_9191,N_7329,N_7181);
and U9192 (N_9192,N_8540,N_8793);
nor U9193 (N_9193,N_7054,N_6089);
and U9194 (N_9194,N_6995,N_8142);
xor U9195 (N_9195,N_6907,N_8995);
nand U9196 (N_9196,N_8814,N_7333);
and U9197 (N_9197,N_6024,N_8777);
nand U9198 (N_9198,N_6735,N_6200);
nand U9199 (N_9199,N_6750,N_8778);
nand U9200 (N_9200,N_6610,N_7663);
nor U9201 (N_9201,N_7762,N_6305);
or U9202 (N_9202,N_7651,N_8902);
xor U9203 (N_9203,N_8528,N_6604);
xnor U9204 (N_9204,N_7044,N_6281);
nor U9205 (N_9205,N_6854,N_8866);
nand U9206 (N_9206,N_6342,N_8152);
or U9207 (N_9207,N_7523,N_8751);
or U9208 (N_9208,N_7065,N_8130);
nor U9209 (N_9209,N_6858,N_7574);
nor U9210 (N_9210,N_6066,N_6561);
xor U9211 (N_9211,N_6910,N_7654);
nand U9212 (N_9212,N_7536,N_7256);
xor U9213 (N_9213,N_7407,N_7309);
xor U9214 (N_9214,N_7125,N_8350);
nor U9215 (N_9215,N_7217,N_6349);
xnor U9216 (N_9216,N_7666,N_6382);
nor U9217 (N_9217,N_6759,N_7398);
nor U9218 (N_9218,N_7204,N_6257);
and U9219 (N_9219,N_6816,N_7102);
xor U9220 (N_9220,N_8570,N_8420);
and U9221 (N_9221,N_6658,N_8931);
or U9222 (N_9222,N_6328,N_7827);
nand U9223 (N_9223,N_6611,N_6931);
or U9224 (N_9224,N_6112,N_8253);
nand U9225 (N_9225,N_7174,N_8542);
nand U9226 (N_9226,N_7103,N_6672);
and U9227 (N_9227,N_7537,N_7269);
and U9228 (N_9228,N_7577,N_8790);
xnor U9229 (N_9229,N_6334,N_7257);
nor U9230 (N_9230,N_8520,N_6478);
xnor U9231 (N_9231,N_6847,N_7807);
xor U9232 (N_9232,N_6481,N_6782);
nor U9233 (N_9233,N_7950,N_7732);
and U9234 (N_9234,N_6652,N_6731);
nand U9235 (N_9235,N_6752,N_7792);
nand U9236 (N_9236,N_8191,N_8617);
or U9237 (N_9237,N_6648,N_8690);
nor U9238 (N_9238,N_6292,N_6933);
or U9239 (N_9239,N_7590,N_6921);
and U9240 (N_9240,N_7639,N_7477);
nor U9241 (N_9241,N_7566,N_8878);
nand U9242 (N_9242,N_7338,N_7626);
or U9243 (N_9243,N_7066,N_7339);
nor U9244 (N_9244,N_6766,N_8281);
and U9245 (N_9245,N_6400,N_6029);
or U9246 (N_9246,N_8492,N_8820);
xor U9247 (N_9247,N_8575,N_6168);
nor U9248 (N_9248,N_8861,N_6720);
or U9249 (N_9249,N_6235,N_8727);
or U9250 (N_9250,N_7271,N_7080);
or U9251 (N_9251,N_8922,N_8217);
nand U9252 (N_9252,N_7959,N_6151);
nand U9253 (N_9253,N_7110,N_6106);
nor U9254 (N_9254,N_8105,N_6818);
and U9255 (N_9255,N_6975,N_6917);
and U9256 (N_9256,N_7085,N_6240);
xor U9257 (N_9257,N_6674,N_6796);
nand U9258 (N_9258,N_6317,N_7446);
or U9259 (N_9259,N_6390,N_8537);
or U9260 (N_9260,N_6934,N_7108);
nor U9261 (N_9261,N_7087,N_8013);
nand U9262 (N_9262,N_6728,N_6557);
nor U9263 (N_9263,N_7186,N_7274);
nand U9264 (N_9264,N_8375,N_8802);
and U9265 (N_9265,N_7652,N_6776);
xnor U9266 (N_9266,N_6104,N_6470);
xor U9267 (N_9267,N_8921,N_8219);
or U9268 (N_9268,N_8085,N_7236);
nand U9269 (N_9269,N_8183,N_7945);
and U9270 (N_9270,N_7192,N_8632);
and U9271 (N_9271,N_7850,N_7417);
nor U9272 (N_9272,N_8107,N_6984);
and U9273 (N_9273,N_6392,N_7290);
and U9274 (N_9274,N_6466,N_6009);
or U9275 (N_9275,N_6530,N_6855);
or U9276 (N_9276,N_8665,N_8504);
or U9277 (N_9277,N_6052,N_6329);
nor U9278 (N_9278,N_6078,N_7994);
or U9279 (N_9279,N_8272,N_7131);
and U9280 (N_9280,N_7794,N_7569);
or U9281 (N_9281,N_8479,N_7378);
xnor U9282 (N_9282,N_8800,N_6068);
or U9283 (N_9283,N_7453,N_8521);
and U9284 (N_9284,N_8658,N_6000);
nand U9285 (N_9285,N_8469,N_6560);
and U9286 (N_9286,N_7126,N_6424);
or U9287 (N_9287,N_6268,N_6957);
and U9288 (N_9288,N_6461,N_7365);
nor U9289 (N_9289,N_7202,N_8651);
xnor U9290 (N_9290,N_7883,N_8401);
or U9291 (N_9291,N_6831,N_7363);
nor U9292 (N_9292,N_8155,N_6551);
nand U9293 (N_9293,N_7433,N_8763);
or U9294 (N_9294,N_7400,N_7943);
xnor U9295 (N_9295,N_8656,N_6602);
xor U9296 (N_9296,N_8361,N_7114);
and U9297 (N_9297,N_8737,N_8355);
xnor U9298 (N_9298,N_8031,N_6339);
xor U9299 (N_9299,N_8503,N_8276);
or U9300 (N_9300,N_8783,N_8990);
and U9301 (N_9301,N_7815,N_7586);
or U9302 (N_9302,N_7752,N_6432);
or U9303 (N_9303,N_7040,N_7306);
nand U9304 (N_9304,N_6203,N_6546);
nor U9305 (N_9305,N_7912,N_8196);
or U9306 (N_9306,N_7886,N_7288);
nand U9307 (N_9307,N_6053,N_8447);
and U9308 (N_9308,N_6275,N_7964);
or U9309 (N_9309,N_7056,N_6362);
xor U9310 (N_9310,N_7464,N_7503);
nor U9311 (N_9311,N_6097,N_7951);
nor U9312 (N_9312,N_8227,N_8764);
nor U9313 (N_9313,N_6215,N_6976);
nor U9314 (N_9314,N_6536,N_8641);
nor U9315 (N_9315,N_7079,N_8884);
nand U9316 (N_9316,N_6476,N_6640);
and U9317 (N_9317,N_8298,N_6636);
xnor U9318 (N_9318,N_8969,N_6673);
xor U9319 (N_9319,N_6310,N_6911);
or U9320 (N_9320,N_8704,N_7060);
or U9321 (N_9321,N_8202,N_6809);
nor U9322 (N_9322,N_7314,N_7233);
nand U9323 (N_9323,N_7069,N_7928);
and U9324 (N_9324,N_8198,N_6491);
xor U9325 (N_9325,N_8439,N_7693);
nand U9326 (N_9326,N_7061,N_6838);
xor U9327 (N_9327,N_7219,N_8951);
and U9328 (N_9328,N_8245,N_8394);
nand U9329 (N_9329,N_8827,N_8919);
and U9330 (N_9330,N_8387,N_7711);
nor U9331 (N_9331,N_7774,N_8065);
or U9332 (N_9332,N_6209,N_6098);
and U9333 (N_9333,N_8747,N_8496);
and U9334 (N_9334,N_7594,N_6490);
xor U9335 (N_9335,N_8176,N_8940);
nand U9336 (N_9336,N_7029,N_8323);
or U9337 (N_9337,N_8433,N_6669);
or U9338 (N_9338,N_7529,N_6058);
xnor U9339 (N_9339,N_6811,N_6260);
and U9340 (N_9340,N_6889,N_7685);
xor U9341 (N_9341,N_7826,N_8961);
or U9342 (N_9342,N_8103,N_8378);
and U9343 (N_9343,N_7983,N_8333);
and U9344 (N_9344,N_6575,N_7638);
xnor U9345 (N_9345,N_8581,N_8937);
xnor U9346 (N_9346,N_6868,N_8434);
nand U9347 (N_9347,N_8384,N_8928);
or U9348 (N_9348,N_8167,N_7379);
nand U9349 (N_9349,N_6888,N_6744);
nor U9350 (N_9350,N_6299,N_7479);
nor U9351 (N_9351,N_6617,N_8335);
nor U9352 (N_9352,N_8881,N_8157);
xor U9353 (N_9353,N_8889,N_6218);
xnor U9354 (N_9354,N_7090,N_6589);
xor U9355 (N_9355,N_8185,N_8660);
and U9356 (N_9356,N_6320,N_7937);
nand U9357 (N_9357,N_7644,N_7848);
xnor U9358 (N_9358,N_8268,N_8950);
or U9359 (N_9359,N_7170,N_6130);
or U9360 (N_9360,N_6002,N_7227);
or U9361 (N_9361,N_8880,N_8236);
nand U9362 (N_9362,N_7776,N_7860);
nand U9363 (N_9363,N_7921,N_6372);
and U9364 (N_9364,N_7028,N_6729);
or U9365 (N_9365,N_8667,N_7361);
or U9366 (N_9366,N_7208,N_8927);
xor U9367 (N_9367,N_8136,N_6608);
nor U9368 (N_9368,N_6925,N_7588);
xor U9369 (N_9369,N_8805,N_7454);
nor U9370 (N_9370,N_6962,N_6724);
and U9371 (N_9371,N_6876,N_8994);
or U9372 (N_9372,N_7035,N_6539);
and U9373 (N_9373,N_8180,N_6411);
nand U9374 (N_9374,N_8140,N_6649);
nand U9375 (N_9375,N_6981,N_8256);
or U9376 (N_9376,N_8767,N_8993);
nand U9377 (N_9377,N_7643,N_6702);
and U9378 (N_9378,N_7357,N_8452);
xor U9379 (N_9379,N_8495,N_6285);
nor U9380 (N_9380,N_7518,N_6745);
nand U9381 (N_9381,N_6348,N_7463);
xnor U9382 (N_9382,N_7345,N_8371);
and U9383 (N_9383,N_6512,N_7713);
or U9384 (N_9384,N_6974,N_8765);
nand U9385 (N_9385,N_6837,N_7962);
or U9386 (N_9386,N_7955,N_6736);
or U9387 (N_9387,N_8794,N_6730);
or U9388 (N_9388,N_7475,N_6195);
nand U9389 (N_9389,N_7787,N_7647);
xor U9390 (N_9390,N_6443,N_7595);
xnor U9391 (N_9391,N_8474,N_7593);
or U9392 (N_9392,N_8037,N_6505);
nor U9393 (N_9393,N_8958,N_8210);
and U9394 (N_9394,N_8870,N_6185);
and U9395 (N_9395,N_7871,N_8139);
nand U9396 (N_9396,N_6792,N_6198);
or U9397 (N_9397,N_8490,N_7443);
and U9398 (N_9398,N_7315,N_8238);
nand U9399 (N_9399,N_7564,N_6395);
nor U9400 (N_9400,N_7058,N_8905);
or U9401 (N_9401,N_7459,N_6890);
and U9402 (N_9402,N_8985,N_7954);
nor U9403 (N_9403,N_8181,N_7384);
or U9404 (N_9404,N_8557,N_7399);
nor U9405 (N_9405,N_6708,N_7451);
nand U9406 (N_9406,N_6276,N_6179);
nand U9407 (N_9407,N_8368,N_7834);
or U9408 (N_9408,N_6944,N_8402);
and U9409 (N_9409,N_8552,N_7411);
nand U9410 (N_9410,N_8682,N_7785);
and U9411 (N_9411,N_7067,N_7386);
nand U9412 (N_9412,N_6621,N_8600);
nor U9413 (N_9413,N_7953,N_6846);
and U9414 (N_9414,N_6634,N_8719);
and U9415 (N_9415,N_8604,N_6594);
nand U9416 (N_9416,N_6895,N_7968);
nand U9417 (N_9417,N_8273,N_6322);
and U9418 (N_9418,N_7323,N_7506);
xor U9419 (N_9419,N_6005,N_6079);
nor U9420 (N_9420,N_7891,N_6851);
or U9421 (N_9421,N_8666,N_6319);
nand U9422 (N_9422,N_6531,N_8113);
nand U9423 (N_9423,N_8771,N_8629);
nor U9424 (N_9424,N_6839,N_6326);
xor U9425 (N_9425,N_7892,N_6685);
xor U9426 (N_9426,N_8529,N_6912);
or U9427 (N_9427,N_8125,N_6946);
nor U9428 (N_9428,N_6398,N_8133);
or U9429 (N_9429,N_8071,N_6219);
and U9430 (N_9430,N_6616,N_6972);
and U9431 (N_9431,N_7700,N_7563);
nand U9432 (N_9432,N_7592,N_8947);
xnor U9433 (N_9433,N_6206,N_6901);
nor U9434 (N_9434,N_7980,N_8399);
and U9435 (N_9435,N_7947,N_6457);
nor U9436 (N_9436,N_8899,N_7686);
and U9437 (N_9437,N_6367,N_6969);
nand U9438 (N_9438,N_6072,N_6763);
xor U9439 (N_9439,N_6264,N_8091);
or U9440 (N_9440,N_8533,N_8513);
or U9441 (N_9441,N_6439,N_7458);
xnor U9442 (N_9442,N_8523,N_6094);
xnor U9443 (N_9443,N_8562,N_6441);
xor U9444 (N_9444,N_7581,N_6897);
nand U9445 (N_9445,N_6711,N_8197);
nor U9446 (N_9446,N_6503,N_8599);
xor U9447 (N_9447,N_7473,N_6801);
nor U9448 (N_9448,N_7782,N_6821);
xnor U9449 (N_9449,N_8486,N_7444);
xnor U9450 (N_9450,N_6228,N_8300);
xnor U9451 (N_9451,N_8935,N_7019);
or U9452 (N_9452,N_6871,N_6891);
or U9453 (N_9453,N_8462,N_8579);
and U9454 (N_9454,N_6823,N_6095);
nand U9455 (N_9455,N_8649,N_8095);
xor U9456 (N_9456,N_8900,N_8644);
and U9457 (N_9457,N_7214,N_7859);
nand U9458 (N_9458,N_7020,N_7049);
or U9459 (N_9459,N_7213,N_8913);
and U9460 (N_9460,N_6288,N_8525);
nand U9461 (N_9461,N_6727,N_7909);
xor U9462 (N_9462,N_7319,N_7764);
or U9463 (N_9463,N_8168,N_6973);
nor U9464 (N_9464,N_6787,N_7063);
and U9465 (N_9465,N_6829,N_6694);
and U9466 (N_9466,N_8694,N_6862);
nor U9467 (N_9467,N_7248,N_8601);
and U9468 (N_9468,N_8920,N_7734);
nand U9469 (N_9469,N_6119,N_7286);
and U9470 (N_9470,N_7367,N_8121);
or U9471 (N_9471,N_7683,N_7350);
and U9472 (N_9472,N_6430,N_7861);
or U9473 (N_9473,N_8606,N_8388);
or U9474 (N_9474,N_8458,N_8189);
and U9475 (N_9475,N_8429,N_8706);
and U9476 (N_9476,N_7511,N_7504);
and U9477 (N_9477,N_7957,N_6881);
xor U9478 (N_9478,N_6110,N_6715);
xor U9479 (N_9479,N_6612,N_8288);
or U9480 (N_9480,N_7462,N_6857);
nor U9481 (N_9481,N_6371,N_6246);
nand U9482 (N_9482,N_6262,N_8858);
nand U9483 (N_9483,N_8652,N_7611);
nor U9484 (N_9484,N_8840,N_7768);
or U9485 (N_9485,N_6475,N_6631);
nand U9486 (N_9486,N_7371,N_6893);
nor U9487 (N_9487,N_6105,N_7562);
and U9488 (N_9488,N_6747,N_7841);
or U9489 (N_9489,N_6263,N_7423);
nand U9490 (N_9490,N_6982,N_8602);
nand U9491 (N_9491,N_7847,N_6103);
nand U9492 (N_9492,N_8973,N_7245);
xor U9493 (N_9493,N_8354,N_8170);
nor U9494 (N_9494,N_7880,N_7326);
nor U9495 (N_9495,N_6990,N_8732);
or U9496 (N_9496,N_8148,N_7844);
nand U9497 (N_9497,N_8382,N_6603);
nand U9498 (N_9498,N_6705,N_7519);
nor U9499 (N_9499,N_6315,N_8852);
nand U9500 (N_9500,N_6379,N_8679);
nand U9501 (N_9501,N_7703,N_8532);
nor U9502 (N_9502,N_8012,N_6120);
or U9503 (N_9503,N_7353,N_8264);
xor U9504 (N_9504,N_6704,N_6438);
or U9505 (N_9505,N_6225,N_6836);
xor U9506 (N_9506,N_7222,N_8470);
and U9507 (N_9507,N_8073,N_8518);
or U9508 (N_9508,N_8297,N_7466);
xnor U9509 (N_9509,N_7781,N_6335);
nand U9510 (N_9510,N_6540,N_6113);
or U9511 (N_9511,N_8662,N_6255);
nor U9512 (N_9512,N_6451,N_8571);
xor U9513 (N_9513,N_7441,N_8488);
nor U9514 (N_9514,N_6865,N_6369);
xnor U9515 (N_9515,N_8590,N_8112);
xnor U9516 (N_9516,N_6687,N_6393);
nand U9517 (N_9517,N_6287,N_8463);
xnor U9518 (N_9518,N_7027,N_7196);
nor U9519 (N_9519,N_8578,N_6375);
or U9520 (N_9520,N_8430,N_8098);
nor U9521 (N_9521,N_7971,N_6015);
nor U9522 (N_9522,N_8165,N_8021);
or U9523 (N_9523,N_7117,N_6389);
nand U9524 (N_9524,N_8159,N_8425);
xnor U9525 (N_9525,N_8316,N_7769);
xor U9526 (N_9526,N_8267,N_7006);
nor U9527 (N_9527,N_7935,N_8246);
and U9528 (N_9528,N_8692,N_7618);
nor U9529 (N_9529,N_7002,N_6093);
nand U9530 (N_9530,N_7415,N_7779);
nor U9531 (N_9531,N_7603,N_7299);
nand U9532 (N_9532,N_7766,N_7148);
xnor U9533 (N_9533,N_7129,N_8186);
or U9534 (N_9534,N_8964,N_8358);
nor U9535 (N_9535,N_7610,N_6992);
nand U9536 (N_9536,N_6807,N_8846);
or U9537 (N_9537,N_7934,N_7938);
nand U9538 (N_9538,N_7911,N_8392);
nor U9539 (N_9539,N_6037,N_8302);
nor U9540 (N_9540,N_6624,N_8768);
or U9541 (N_9541,N_7190,N_8201);
nand U9542 (N_9542,N_8129,N_8405);
or U9543 (N_9543,N_7356,N_6345);
and U9544 (N_9544,N_7923,N_8211);
nor U9545 (N_9545,N_6211,N_7383);
and U9546 (N_9546,N_6591,N_6452);
nor U9547 (N_9547,N_7716,N_7416);
nand U9548 (N_9548,N_8631,N_8143);
or U9549 (N_9549,N_8408,N_7933);
nor U9550 (N_9550,N_8484,N_8828);
nor U9551 (N_9551,N_8806,N_6416);
or U9552 (N_9552,N_6488,N_7366);
or U9553 (N_9553,N_6983,N_7583);
or U9554 (N_9554,N_7553,N_8441);
nor U9555 (N_9555,N_8715,N_8305);
and U9556 (N_9556,N_7757,N_8696);
xnor U9557 (N_9557,N_8548,N_8752);
and U9558 (N_9558,N_8887,N_8932);
or U9559 (N_9559,N_7502,N_7283);
nand U9560 (N_9560,N_6298,N_7557);
and U9561 (N_9561,N_8230,N_6810);
nand U9562 (N_9562,N_8825,N_6295);
or U9563 (N_9563,N_6563,N_7455);
nor U9564 (N_9564,N_8565,N_8195);
nand U9565 (N_9565,N_7033,N_7642);
xor U9566 (N_9566,N_6945,N_6559);
or U9567 (N_9567,N_7662,N_7570);
nor U9568 (N_9568,N_8092,N_6141);
and U9569 (N_9569,N_6012,N_6663);
xor U9570 (N_9570,N_8188,N_7927);
and U9571 (N_9571,N_7648,N_7600);
or U9572 (N_9572,N_7667,N_7426);
and U9573 (N_9573,N_6396,N_8707);
nor U9574 (N_9574,N_6454,N_8385);
or U9575 (N_9575,N_6138,N_7942);
and U9576 (N_9576,N_7083,N_6408);
nor U9577 (N_9577,N_8367,N_8128);
nand U9578 (N_9578,N_8669,N_7347);
and U9579 (N_9579,N_7528,N_7438);
xor U9580 (N_9580,N_8539,N_8339);
and U9581 (N_9581,N_8340,N_8106);
or U9582 (N_9582,N_6397,N_8511);
xnor U9583 (N_9583,N_6020,N_8193);
nand U9584 (N_9584,N_7034,N_7816);
nand U9585 (N_9585,N_8586,N_7849);
or U9586 (N_9586,N_8449,N_8731);
nor U9587 (N_9587,N_7817,N_7887);
nand U9588 (N_9588,N_6999,N_6832);
nand U9589 (N_9589,N_6014,N_6896);
xnor U9590 (N_9590,N_7545,N_7527);
or U9591 (N_9591,N_7540,N_7837);
nor U9592 (N_9592,N_6994,N_6784);
nand U9593 (N_9593,N_7089,N_8228);
nor U9594 (N_9594,N_8062,N_6980);
nand U9595 (N_9595,N_7554,N_6189);
nand U9596 (N_9596,N_7336,N_8972);
xnor U9597 (N_9597,N_6210,N_8035);
or U9598 (N_9598,N_6247,N_6242);
and U9599 (N_9599,N_8365,N_6544);
nand U9600 (N_9600,N_7704,N_6526);
or U9601 (N_9601,N_6472,N_6277);
and U9602 (N_9602,N_6043,N_8551);
or U9603 (N_9603,N_6327,N_8233);
xnor U9604 (N_9604,N_6156,N_8908);
or U9605 (N_9605,N_7440,N_8436);
or U9606 (N_9606,N_8005,N_8568);
and U9607 (N_9607,N_8832,N_7491);
nor U9608 (N_9608,N_8004,N_6509);
nand U9609 (N_9609,N_8424,N_8026);
xor U9610 (N_9610,N_7727,N_8811);
and U9611 (N_9611,N_6493,N_6133);
nand U9612 (N_9612,N_6764,N_6650);
or U9613 (N_9613,N_8847,N_8328);
nand U9614 (N_9614,N_7410,N_7736);
or U9615 (N_9615,N_7913,N_8797);
nand U9616 (N_9616,N_6172,N_6725);
and U9617 (N_9617,N_8573,N_8247);
nor U9618 (N_9618,N_6800,N_8845);
nand U9619 (N_9619,N_8048,N_8427);
nand U9620 (N_9620,N_7952,N_6637);
nor U9621 (N_9621,N_7022,N_6507);
or U9622 (N_9622,N_6028,N_8244);
nor U9623 (N_9623,N_6044,N_8151);
xor U9624 (N_9624,N_7973,N_7810);
nor U9625 (N_9625,N_7744,N_7836);
and U9626 (N_9626,N_8251,N_8404);
xor U9627 (N_9627,N_7993,N_7535);
nor U9628 (N_9628,N_7013,N_6779);
xnor U9629 (N_9629,N_8645,N_8863);
nand U9630 (N_9630,N_8024,N_6709);
or U9631 (N_9631,N_6300,N_7832);
nor U9632 (N_9632,N_6842,N_6176);
nor U9633 (N_9633,N_8924,N_6555);
nand U9634 (N_9634,N_7070,N_6374);
xor U9635 (N_9635,N_7854,N_7790);
nand U9636 (N_9636,N_7068,N_6515);
nor U9637 (N_9637,N_6742,N_8746);
xor U9638 (N_9638,N_7877,N_8739);
nand U9639 (N_9639,N_7289,N_8116);
and U9640 (N_9640,N_7260,N_8971);
xor U9641 (N_9641,N_6948,N_7977);
xnor U9642 (N_9642,N_8218,N_7821);
or U9643 (N_9643,N_7397,N_6127);
nand U9644 (N_9644,N_8989,N_8349);
xnor U9645 (N_9645,N_8419,N_7885);
nand U9646 (N_9646,N_7949,N_7422);
xor U9647 (N_9647,N_8122,N_6344);
nor U9648 (N_9648,N_6826,N_7998);
xnor U9649 (N_9649,N_8014,N_8953);
nand U9650 (N_9650,N_8467,N_7303);
nand U9651 (N_9651,N_6898,N_6191);
nand U9652 (N_9652,N_6062,N_7193);
and U9653 (N_9653,N_8321,N_7758);
nor U9654 (N_9654,N_7252,N_7780);
nand U9655 (N_9655,N_6580,N_8988);
nand U9656 (N_9656,N_7888,N_7230);
and U9657 (N_9657,N_8057,N_7922);
and U9658 (N_9658,N_8946,N_8008);
and U9659 (N_9659,N_6283,N_7803);
nor U9660 (N_9660,N_6306,N_8728);
and U9661 (N_9661,N_7584,N_6224);
xnor U9662 (N_9662,N_6519,N_7197);
xor U9663 (N_9663,N_8705,N_7207);
xor U9664 (N_9664,N_7489,N_8558);
nand U9665 (N_9665,N_7015,N_8837);
nor U9666 (N_9666,N_6364,N_8046);
xor U9667 (N_9667,N_7031,N_6440);
or U9668 (N_9668,N_8515,N_8206);
nor U9669 (N_9669,N_7304,N_7967);
and U9670 (N_9670,N_6100,N_7856);
and U9671 (N_9671,N_6483,N_7948);
or U9672 (N_9672,N_8187,N_6163);
nand U9673 (N_9673,N_8779,N_8455);
and U9674 (N_9674,N_7525,N_8296);
nand U9675 (N_9675,N_7420,N_8120);
and U9676 (N_9676,N_8998,N_7412);
or U9677 (N_9677,N_8997,N_7558);
nand U9678 (N_9678,N_7183,N_6006);
nor U9679 (N_9679,N_8954,N_7374);
nor U9680 (N_9680,N_8844,N_6524);
nand U9681 (N_9681,N_6414,N_6145);
and U9682 (N_9682,N_8547,N_7675);
xnor U9683 (N_9683,N_6692,N_6533);
xnor U9684 (N_9684,N_8076,N_6463);
xnor U9685 (N_9685,N_8984,N_8625);
xnor U9686 (N_9686,N_6588,N_6102);
nor U9687 (N_9687,N_7485,N_6354);
or U9688 (N_9688,N_6537,N_6357);
xor U9689 (N_9689,N_7995,N_8560);
and U9690 (N_9690,N_8326,N_6458);
and U9691 (N_9691,N_8713,N_8291);
nor U9692 (N_9692,N_6869,N_7272);
nand U9693 (N_9693,N_8615,N_8595);
and U9694 (N_9694,N_8249,N_6338);
nand U9695 (N_9695,N_6075,N_6564);
xnor U9696 (N_9696,N_8854,N_8407);
xor U9697 (N_9697,N_7448,N_6892);
nand U9698 (N_9698,N_8101,N_6528);
xor U9699 (N_9699,N_6385,N_7163);
nand U9700 (N_9700,N_8554,N_7924);
nor U9701 (N_9701,N_6997,N_6656);
and U9702 (N_9702,N_6963,N_8212);
nand U9703 (N_9703,N_8670,N_7021);
nor U9704 (N_9704,N_8917,N_7032);
or U9705 (N_9705,N_7717,N_8266);
nand U9706 (N_9706,N_8630,N_7184);
nor U9707 (N_9707,N_7342,N_7344);
nor U9708 (N_9708,N_7188,N_8331);
nor U9709 (N_9709,N_7684,N_8655);
nor U9710 (N_9710,N_8160,N_7437);
or U9711 (N_9711,N_6527,N_7328);
nand U9712 (N_9712,N_8796,N_6459);
nand U9713 (N_9713,N_6290,N_6918);
or U9714 (N_9714,N_8393,N_6873);
xnor U9715 (N_9715,N_8357,N_7284);
or U9716 (N_9716,N_6586,N_8510);
or U9717 (N_9717,N_6121,N_6790);
or U9718 (N_9718,N_6859,N_8996);
nor U9719 (N_9719,N_7387,N_7944);
xor U9720 (N_9720,N_7770,N_6556);
and U9721 (N_9721,N_8531,N_7059);
and U9722 (N_9722,N_6070,N_6952);
nor U9723 (N_9723,N_8755,N_6083);
nor U9724 (N_9724,N_8443,N_8254);
xnor U9725 (N_9725,N_8061,N_8255);
or U9726 (N_9726,N_8327,N_6254);
and U9727 (N_9727,N_8444,N_8559);
nand U9728 (N_9728,N_6330,N_8248);
nor U9729 (N_9729,N_6403,N_8414);
or U9730 (N_9730,N_6848,N_6795);
or U9731 (N_9731,N_7742,N_7429);
and U9732 (N_9732,N_8535,N_6579);
xnor U9733 (N_9733,N_6422,N_6054);
nand U9734 (N_9734,N_6835,N_6943);
or U9735 (N_9735,N_8813,N_7940);
or U9736 (N_9736,N_6304,N_8314);
xor U9737 (N_9737,N_6815,N_7646);
nand U9738 (N_9738,N_6508,N_7508);
xnor U9739 (N_9739,N_8282,N_6657);
nor U9740 (N_9740,N_7209,N_8034);
nor U9741 (N_9741,N_8753,N_6545);
nor U9742 (N_9742,N_7442,N_7763);
xnor U9743 (N_9743,N_6819,N_6067);
and U9744 (N_9744,N_6552,N_6383);
xnor U9745 (N_9745,N_6820,N_7312);
nor U9746 (N_9746,N_7706,N_7310);
xor U9747 (N_9747,N_8262,N_8585);
nand U9748 (N_9748,N_8491,N_8308);
and U9749 (N_9749,N_7316,N_7198);
or U9750 (N_9750,N_8851,N_8505);
nand U9751 (N_9751,N_8089,N_8986);
or U9752 (N_9752,N_7656,N_6665);
and U9753 (N_9753,N_7082,N_7512);
or U9754 (N_9754,N_7493,N_6178);
or U9755 (N_9755,N_7632,N_7240);
xnor U9756 (N_9756,N_7918,N_8123);
nor U9757 (N_9757,N_8099,N_8074);
or U9758 (N_9758,N_7320,N_6253);
xnor U9759 (N_9759,N_8250,N_6651);
and U9760 (N_9760,N_7203,N_8161);
or U9761 (N_9761,N_6164,N_7402);
nand U9762 (N_9762,N_6718,N_8237);
xor U9763 (N_9763,N_6756,N_6712);
nor U9764 (N_9764,N_8634,N_7789);
xnor U9765 (N_9765,N_7242,N_7294);
nor U9766 (N_9766,N_7974,N_7043);
or U9767 (N_9767,N_8850,N_8043);
xor U9768 (N_9768,N_7691,N_7929);
and U9769 (N_9769,N_6501,N_7368);
nor U9770 (N_9770,N_8030,N_6456);
nor U9771 (N_9771,N_8208,N_8329);
and U9772 (N_9772,N_6647,N_7111);
nand U9773 (N_9773,N_6597,N_8241);
xnor U9774 (N_9774,N_6477,N_6698);
and U9775 (N_9775,N_6929,N_6970);
and U9776 (N_9776,N_7615,N_6343);
or U9777 (N_9777,N_6086,N_6180);
xnor U9778 (N_9778,N_8042,N_8028);
and U9779 (N_9779,N_7143,N_7986);
or U9780 (N_9780,N_8395,N_8598);
and U9781 (N_9781,N_8774,N_6064);
or U9782 (N_9782,N_7753,N_7517);
or U9783 (N_9783,N_7301,N_8700);
nor U9784 (N_9784,N_7141,N_7205);
and U9785 (N_9785,N_7376,N_8735);
or U9786 (N_9786,N_7285,N_8642);
nand U9787 (N_9787,N_8991,N_8147);
nand U9788 (N_9788,N_8226,N_8810);
and U9789 (N_9789,N_6915,N_8610);
nand U9790 (N_9790,N_8640,N_8929);
nand U9791 (N_9791,N_7468,N_7169);
nand U9792 (N_9792,N_8607,N_7530);
nand U9793 (N_9793,N_8284,N_6427);
and U9794 (N_9794,N_7036,N_7225);
and U9795 (N_9795,N_7559,N_7941);
nand U9796 (N_9796,N_7200,N_8594);
nor U9797 (N_9797,N_6867,N_6032);
xor U9798 (N_9798,N_8169,N_6991);
nand U9799 (N_9799,N_7234,N_6353);
xnor U9800 (N_9800,N_8957,N_7809);
xnor U9801 (N_9801,N_8199,N_8582);
xnor U9802 (N_9802,N_7046,N_7393);
and U9803 (N_9803,N_7171,N_7097);
nor U9804 (N_9804,N_8359,N_6177);
nor U9805 (N_9805,N_7352,N_8431);
xor U9806 (N_9806,N_7388,N_8215);
xor U9807 (N_9807,N_8750,N_6446);
nand U9808 (N_9808,N_6272,N_8192);
and U9809 (N_9809,N_6618,N_6558);
xor U9810 (N_9810,N_7311,N_7436);
nand U9811 (N_9811,N_8104,N_6405);
xor U9812 (N_9812,N_7620,N_6950);
nor U9813 (N_9813,N_7805,N_7302);
xnor U9814 (N_9814,N_7501,N_6894);
or U9815 (N_9815,N_8001,N_8239);
nand U9816 (N_9816,N_6679,N_8628);
nor U9817 (N_9817,N_7802,N_6532);
xor U9818 (N_9818,N_7275,N_8162);
and U9819 (N_9819,N_8362,N_8039);
and U9820 (N_9820,N_7492,N_7162);
nand U9821 (N_9821,N_6157,N_6449);
xor U9822 (N_9822,N_7801,N_6722);
xnor U9823 (N_9823,N_7246,N_6388);
nor U9824 (N_9824,N_7671,N_8078);
or U9825 (N_9825,N_6035,N_7158);
or U9826 (N_9826,N_8674,N_6955);
nor U9827 (N_9827,N_7297,N_7905);
or U9828 (N_9828,N_8966,N_8960);
and U9829 (N_9829,N_7098,N_8481);
xor U9830 (N_9830,N_6084,N_8093);
nand U9831 (N_9831,N_8833,N_6849);
nand U9832 (N_9832,N_8352,N_6958);
xnor U9833 (N_9833,N_8769,N_7091);
xnor U9834 (N_9834,N_6550,N_7337);
nor U9835 (N_9835,N_7406,N_7104);
xnor U9836 (N_9836,N_6038,N_7916);
nor U9837 (N_9837,N_8220,N_8478);
nand U9838 (N_9838,N_7889,N_8886);
nand U9839 (N_9839,N_8689,N_6863);
nand U9840 (N_9840,N_7958,N_8910);
nor U9841 (N_9841,N_8970,N_6118);
xor U9842 (N_9842,N_6142,N_8781);
or U9843 (N_9843,N_7052,N_8923);
nor U9844 (N_9844,N_7372,N_8214);
or U9845 (N_9845,N_7296,N_8687);
xnor U9846 (N_9846,N_6639,N_6641);
nand U9847 (N_9847,N_8830,N_7005);
xnor U9848 (N_9848,N_7866,N_7321);
or U9849 (N_9849,N_6900,N_6337);
and U9850 (N_9850,N_6932,N_8841);
nand U9851 (N_9851,N_7369,N_7992);
nand U9852 (N_9852,N_6680,N_7370);
nor U9853 (N_9853,N_6959,N_8299);
and U9854 (N_9854,N_8224,N_7963);
or U9855 (N_9855,N_8324,N_7699);
nand U9856 (N_9856,N_8111,N_6197);
nand U9857 (N_9857,N_8477,N_7910);
xor U9858 (N_9858,N_7480,N_7221);
xnor U9859 (N_9859,N_8725,N_6232);
nand U9860 (N_9860,N_7778,N_6599);
or U9861 (N_9861,N_8499,N_8067);
nor U9862 (N_9862,N_8126,N_7023);
xor U9863 (N_9863,N_7133,N_8965);
and U9864 (N_9864,N_6737,N_8941);
xnor U9865 (N_9865,N_8307,N_6129);
and U9866 (N_9866,N_6902,N_8280);
nor U9867 (N_9867,N_6107,N_8011);
and U9868 (N_9868,N_6845,N_8915);
nand U9869 (N_9869,N_6222,N_7606);
nand U9870 (N_9870,N_7445,N_7729);
nand U9871 (N_9871,N_8334,N_8967);
and U9872 (N_9872,N_7050,N_6047);
nor U9873 (N_9873,N_6417,N_6977);
and U9874 (N_9874,N_8816,N_6124);
nand U9875 (N_9875,N_7268,N_6048);
nand U9876 (N_9876,N_7403,N_8108);
xnor U9877 (N_9877,N_7726,N_8675);
or U9878 (N_9878,N_8592,N_8673);
nand U9879 (N_9879,N_6025,N_7864);
or U9880 (N_9880,N_7228,N_6125);
xnor U9881 (N_9881,N_6696,N_6935);
or U9882 (N_9882,N_6160,N_8440);
and U9883 (N_9883,N_8555,N_7708);
and U9884 (N_9884,N_8683,N_8446);
nand U9885 (N_9885,N_8003,N_8891);
xor U9886 (N_9886,N_6311,N_6517);
and U9887 (N_9887,N_6150,N_7689);
nand U9888 (N_9888,N_6437,N_8633);
nand U9889 (N_9889,N_8124,N_6961);
nand U9890 (N_9890,N_7199,N_8287);
nand U9891 (N_9891,N_7599,N_6479);
nor U9892 (N_9892,N_6717,N_8259);
or U9893 (N_9893,N_8088,N_8489);
or U9894 (N_9894,N_7602,N_6788);
nand U9895 (N_9895,N_6274,N_8231);
nand U9896 (N_9896,N_8831,N_7435);
or U9897 (N_9897,N_6109,N_8945);
and U9898 (N_9898,N_7003,N_7745);
nand U9899 (N_9899,N_7688,N_8019);
nand U9900 (N_9900,N_6045,N_6817);
nor U9901 (N_9901,N_8789,N_8223);
or U9902 (N_9902,N_7605,N_7165);
and U9903 (N_9903,N_6147,N_6291);
xnor U9904 (N_9904,N_7879,N_6905);
xnor U9905 (N_9905,N_7137,N_7796);
or U9906 (N_9906,N_8860,N_6676);
xor U9907 (N_9907,N_7449,N_8877);
xor U9908 (N_9908,N_6769,N_7325);
nand U9909 (N_9909,N_6908,N_7472);
or U9910 (N_9910,N_6148,N_6721);
xnor U9911 (N_9911,N_6302,N_7546);
xor U9912 (N_9912,N_8080,N_6122);
and U9913 (N_9913,N_6308,N_8338);
nand U9914 (N_9914,N_7743,N_7392);
nor U9915 (N_9915,N_6495,N_7718);
and U9916 (N_9916,N_7255,N_7681);
nand U9917 (N_9917,N_7694,N_6117);
nor U9918 (N_9918,N_8163,N_8040);
xnor U9919 (N_9919,N_6852,N_6833);
or U9920 (N_9920,N_8265,N_7526);
and U9921 (N_9921,N_7722,N_8475);
or U9922 (N_9922,N_7636,N_7874);
and U9923 (N_9923,N_6394,N_7327);
or U9924 (N_9924,N_8471,N_8442);
xor U9925 (N_9925,N_6386,N_6986);
nand U9926 (N_9926,N_8386,N_8591);
nand U9927 (N_9927,N_7340,N_6415);
or U9928 (N_9928,N_6356,N_8260);
or U9929 (N_9929,N_7872,N_6840);
nand U9930 (N_9930,N_7567,N_6153);
or U9931 (N_9931,N_8416,N_6376);
and U9932 (N_9932,N_6684,N_6653);
nor U9933 (N_9933,N_7259,N_6165);
xnor U9934 (N_9934,N_8733,N_7086);
and U9935 (N_9935,N_6010,N_6566);
nor U9936 (N_9936,N_7109,N_8029);
or U9937 (N_9937,N_6543,N_6828);
nor U9938 (N_9938,N_7845,N_8271);
and U9939 (N_9939,N_7867,N_8059);
nand U9940 (N_9940,N_7900,N_8473);
nand U9941 (N_9941,N_6774,N_8526);
xor U9942 (N_9942,N_6402,N_7561);
or U9943 (N_9943,N_7741,N_6570);
nand U9944 (N_9944,N_7447,N_8200);
xor U9945 (N_9945,N_8882,N_6571);
nand U9946 (N_9946,N_6312,N_7804);
or U9947 (N_9947,N_7161,N_6484);
and U9948 (N_9948,N_8597,N_6271);
nand U9949 (N_9949,N_8150,N_7071);
nand U9950 (N_9950,N_6360,N_6710);
and U9951 (N_9951,N_8762,N_7982);
nor U9952 (N_9952,N_8621,N_6701);
nand U9953 (N_9953,N_8179,N_6940);
nand U9954 (N_9954,N_7324,N_7166);
nand U9955 (N_9955,N_7609,N_6226);
or U9956 (N_9956,N_6985,N_6592);
nor U9957 (N_9957,N_6733,N_6581);
nor U9958 (N_9958,N_7122,N_7012);
nand U9959 (N_9959,N_8397,N_6553);
xor U9960 (N_9960,N_7721,N_7707);
and U9961 (N_9961,N_7607,N_6691);
xor U9962 (N_9962,N_7351,N_6625);
nor U9963 (N_9963,N_7360,N_6229);
nor U9964 (N_9964,N_7702,N_6429);
and U9965 (N_9965,N_8843,N_6740);
nor U9966 (N_9966,N_7657,N_6645);
nor U9967 (N_9967,N_8381,N_8522);
or U9968 (N_9968,N_7698,N_8509);
xor U9969 (N_9969,N_6523,N_7024);
or U9970 (N_9970,N_7244,N_8410);
nor U9971 (N_9971,N_7739,N_8549);
and U9972 (N_9972,N_8476,N_8864);
or U9973 (N_9973,N_7358,N_6057);
xnor U9974 (N_9974,N_8345,N_8890);
nand U9975 (N_9975,N_8596,N_6775);
or U9976 (N_9976,N_7630,N_7931);
nand U9977 (N_9977,N_8786,N_7870);
or U9978 (N_9978,N_6620,N_6063);
nand U9979 (N_9979,N_8175,N_8712);
or U9980 (N_9980,N_6187,N_6194);
or U9981 (N_9981,N_8258,N_6978);
xor U9982 (N_9982,N_8678,N_8853);
and U9983 (N_9983,N_8466,N_7926);
and U9984 (N_9984,N_8094,N_8978);
or U9985 (N_9985,N_7127,N_7645);
and U9986 (N_9986,N_7783,N_8072);
nand U9987 (N_9987,N_7800,N_7895);
or U9988 (N_9988,N_6001,N_8154);
or U9989 (N_9989,N_6018,N_7136);
nand U9990 (N_9990,N_7930,N_7243);
or U9991 (N_9991,N_8485,N_8943);
or U9992 (N_9992,N_6233,N_6196);
and U9993 (N_9993,N_7305,N_8390);
or U9994 (N_9994,N_7978,N_6697);
nor U9995 (N_9995,N_6549,N_7538);
nand U9996 (N_9996,N_8896,N_7532);
nand U9997 (N_9997,N_7746,N_8025);
nor U9998 (N_9998,N_6448,N_7682);
nand U9999 (N_9999,N_6071,N_7701);
xor U10000 (N_10000,N_6968,N_7735);
xor U10001 (N_10001,N_8261,N_6903);
and U10002 (N_10002,N_7151,N_6423);
or U10003 (N_10003,N_8782,N_7152);
nor U10004 (N_10004,N_7431,N_8015);
and U10005 (N_10005,N_7088,N_6798);
nand U10006 (N_10006,N_8663,N_8819);
and U10007 (N_10007,N_6850,N_8729);
and U10008 (N_10008,N_8758,N_6886);
nand U10009 (N_10009,N_8541,N_6085);
nand U10010 (N_10010,N_8304,N_7414);
nand U10011 (N_10011,N_7806,N_8438);
xnor U10012 (N_10012,N_8453,N_7346);
and U10013 (N_10013,N_6123,N_8564);
or U10014 (N_10014,N_8545,N_6516);
and U10015 (N_10015,N_7150,N_8740);
xnor U10016 (N_10016,N_6355,N_7481);
or U10017 (N_10017,N_7514,N_6245);
xnor U10018 (N_10018,N_7128,N_8216);
xor U10019 (N_10019,N_6562,N_7670);
nor U10020 (N_10020,N_8711,N_7875);
and U10021 (N_10021,N_7261,N_8171);
nand U10022 (N_10022,N_8637,N_7478);
nor U10023 (N_10023,N_7330,N_7725);
and U10024 (N_10024,N_8315,N_7105);
and U10025 (N_10025,N_6069,N_8680);
nand U10026 (N_10026,N_6743,N_7828);
xor U10027 (N_10027,N_8734,N_6022);
nand U10028 (N_10028,N_8874,N_6004);
xnor U10029 (N_10029,N_7755,N_6021);
nand U10030 (N_10030,N_6780,N_7976);
nand U10031 (N_10031,N_6825,N_8225);
and U10032 (N_10032,N_6993,N_7488);
nand U10033 (N_10033,N_7917,N_8050);
nor U10034 (N_10034,N_6677,N_6938);
nor U10035 (N_10035,N_8624,N_8413);
nor U10036 (N_10036,N_8346,N_7249);
or U10037 (N_10037,N_8627,N_7153);
nand U10038 (N_10038,N_6039,N_7908);
nor U10039 (N_10039,N_6791,N_8418);
and U10040 (N_10040,N_6008,N_8454);
or U10041 (N_10041,N_7270,N_8508);
or U10042 (N_10042,N_8482,N_8671);
or U10043 (N_10043,N_7898,N_7873);
nor U10044 (N_10044,N_8983,N_8240);
or U10045 (N_10045,N_7094,N_6297);
or U10046 (N_10046,N_8736,N_6321);
nand U10047 (N_10047,N_6607,N_8836);
nand U10048 (N_10048,N_6280,N_7045);
or U10049 (N_10049,N_6213,N_8051);
nand U10050 (N_10050,N_7132,N_8450);
and U10051 (N_10051,N_7547,N_8742);
nor U10052 (N_10052,N_7749,N_8077);
nor U10053 (N_10053,N_8376,N_7250);
nor U10054 (N_10054,N_8944,N_7178);
xnor U10055 (N_10055,N_8516,N_8799);
nand U10056 (N_10056,N_8153,N_7858);
nor U10057 (N_10057,N_7465,N_8809);
or U10058 (N_10058,N_8686,N_6428);
xnor U10059 (N_10059,N_7868,N_8982);
and U10060 (N_10060,N_6404,N_8353);
or U10061 (N_10061,N_6541,N_6748);
and U10062 (N_10062,N_7556,N_6132);
xor U10063 (N_10063,N_7317,N_8681);
or U10064 (N_10064,N_8608,N_6221);
and U10065 (N_10065,N_8918,N_7180);
or U10066 (N_10066,N_6137,N_8879);
nor U10067 (N_10067,N_8426,N_8855);
nor U10068 (N_10068,N_6749,N_7001);
nand U10069 (N_10069,N_8177,N_6223);
or U10070 (N_10070,N_8684,N_7404);
or U10071 (N_10071,N_6340,N_7116);
and U10072 (N_10072,N_6381,N_7291);
xor U10073 (N_10073,N_8461,N_8605);
nor U10074 (N_10074,N_7232,N_8527);
and U10075 (N_10075,N_8285,N_7239);
and U10076 (N_10076,N_7548,N_7915);
nor U10077 (N_10077,N_7604,N_8664);
xnor U10078 (N_10078,N_8110,N_6671);
xor U10079 (N_10079,N_6765,N_8761);
and U10080 (N_10080,N_8883,N_7432);
xor U10081 (N_10081,N_7897,N_8325);
nor U10082 (N_10082,N_7018,N_7101);
xor U10083 (N_10083,N_7541,N_8826);
nor U10084 (N_10084,N_6596,N_7000);
xnor U10085 (N_10085,N_6409,N_8942);
nor U10086 (N_10086,N_7907,N_7156);
nor U10087 (N_10087,N_6732,N_7348);
nor U10088 (N_10088,N_8812,N_8501);
and U10089 (N_10089,N_8396,N_6529);
or U10090 (N_10090,N_6864,N_8857);
and U10091 (N_10091,N_8872,N_8614);
nor U10092 (N_10092,N_6017,N_7798);
nand U10093 (N_10093,N_7617,N_7175);
and U10094 (N_10094,N_6184,N_7808);
nand U10095 (N_10095,N_7970,N_8047);
and U10096 (N_10096,N_6217,N_8976);
and U10097 (N_10097,N_8638,N_7226);
xnor U10098 (N_10098,N_7894,N_7533);
or U10099 (N_10099,N_6565,N_8716);
nor U10100 (N_10100,N_7210,N_7784);
xnor U10101 (N_10101,N_6632,N_8135);
nor U10102 (N_10102,N_8109,N_6234);
xor U10103 (N_10103,N_8364,N_6590);
and U10104 (N_10104,N_8563,N_8309);
nand U10105 (N_10105,N_6460,N_6706);
xnor U10106 (N_10106,N_7037,N_7408);
nand U10107 (N_10107,N_8962,N_8117);
xor U10108 (N_10108,N_7185,N_8885);
nand U10109 (N_10109,N_6486,N_6384);
nor U10110 (N_10110,N_7014,N_7373);
nand U10111 (N_10111,N_6301,N_6941);
xor U10112 (N_10112,N_8718,N_7500);
xnor U10113 (N_10113,N_8500,N_6615);
xnor U10114 (N_10114,N_7901,N_8055);
nor U10115 (N_10115,N_6988,N_8572);
xor U10116 (N_10116,N_6282,N_8235);
and U10117 (N_10117,N_8318,N_7146);
nand U10118 (N_10118,N_8834,N_8009);
nor U10119 (N_10119,N_7469,N_7842);
nand U10120 (N_10120,N_6324,N_7544);
and U10121 (N_10121,N_7771,N_6755);
nor U10122 (N_10122,N_8709,N_7659);
xor U10123 (N_10123,N_7292,N_8086);
nand U10124 (N_10124,N_7295,N_8493);
xor U10125 (N_10125,N_8017,N_7380);
and U10126 (N_10126,N_6614,N_8312);
nand U10127 (N_10127,N_8332,N_6425);
nand U10128 (N_10128,N_7591,N_7655);
and U10129 (N_10129,N_8070,N_6442);
xnor U10130 (N_10130,N_8553,N_8290);
nor U10131 (N_10131,N_7187,N_6824);
nand U10132 (N_10132,N_8603,N_8274);
or U10133 (N_10133,N_6605,N_7390);
and U10134 (N_10134,N_6241,N_6587);
nand U10135 (N_10135,N_8934,N_8577);
or U10136 (N_10136,N_8415,N_8914);
xnor U10137 (N_10137,N_7975,N_6626);
or U10138 (N_10138,N_7430,N_8992);
nor U10139 (N_10139,N_7623,N_7266);
nor U10140 (N_10140,N_8313,N_8543);
or U10141 (N_10141,N_8090,N_8963);
xor U10142 (N_10142,N_8000,N_7206);
nand U10143 (N_10143,N_8119,N_7509);
xnor U10144 (N_10144,N_7483,N_7130);
and U10145 (N_10145,N_7756,N_8149);
xor U10146 (N_10146,N_6350,N_6754);
xor U10147 (N_10147,N_6046,N_7914);
or U10148 (N_10148,N_8987,N_7677);
nor U10149 (N_10149,N_6347,N_7238);
nand U10150 (N_10150,N_8760,N_7786);
nand U10151 (N_10151,N_8069,N_8894);
nor U10152 (N_10152,N_8873,N_7123);
nor U10153 (N_10153,N_6568,N_7505);
xnor U10154 (N_10154,N_7999,N_6899);
xnor U10155 (N_10155,N_8584,N_8243);
nor U10156 (N_10156,N_8795,N_6767);
nor U10157 (N_10157,N_6513,N_8888);
xnor U10158 (N_10158,N_6059,N_7960);
or U10159 (N_10159,N_7313,N_6510);
or U10160 (N_10160,N_8049,N_7115);
nand U10161 (N_10161,N_6638,N_8100);
xnor U10162 (N_10162,N_6953,N_8459);
and U10163 (N_10163,N_6822,N_6251);
nor U10164 (N_10164,N_7695,N_6668);
nor U10165 (N_10165,N_6660,N_6471);
nand U10166 (N_10166,N_8127,N_8697);
nor U10167 (N_10167,N_7882,N_8374);
nand U10168 (N_10168,N_6436,N_6841);
nand U10169 (N_10169,N_6885,N_6583);
nand U10170 (N_10170,N_6188,N_7280);
or U10171 (N_10171,N_7513,N_8036);
and U10172 (N_10172,N_7751,N_6289);
nor U10173 (N_10173,N_6535,N_8720);
nand U10174 (N_10174,N_6042,N_8007);
or U10175 (N_10175,N_6622,N_6703);
and U10176 (N_10176,N_8343,N_6431);
xor U10177 (N_10177,N_8056,N_7042);
nand U10178 (N_10178,N_7697,N_8588);
or U10179 (N_10179,N_6804,N_8804);
xor U10180 (N_10180,N_7179,N_7825);
xor U10181 (N_10181,N_8158,N_7549);
xor U10182 (N_10182,N_8311,N_7470);
nor U10183 (N_10183,N_6690,N_6192);
xor U10184 (N_10184,N_6421,N_6050);
nor U10185 (N_10185,N_8618,N_6655);
or U10186 (N_10186,N_6686,N_7263);
or U10187 (N_10187,N_6003,N_6789);
xor U10188 (N_10188,N_7055,N_7418);
or U10189 (N_10189,N_7906,N_8773);
xnor U10190 (N_10190,N_6751,N_7521);
nor U10191 (N_10191,N_6088,N_7253);
xnor U10192 (N_10192,N_6155,N_6323);
nor U10193 (N_10193,N_8134,N_7084);
nor U10194 (N_10194,N_7281,N_8776);
and U10195 (N_10195,N_8222,N_7524);
or U10196 (N_10196,N_8319,N_7838);
xor U10197 (N_10197,N_8808,N_8391);
nor U10198 (N_10198,N_7696,N_7862);
nand U10199 (N_10199,N_8451,N_8613);
or U10200 (N_10200,N_8114,N_6351);
or U10201 (N_10201,N_7575,N_6314);
nor U10202 (N_10202,N_6884,N_6239);
and U10203 (N_10203,N_6258,N_7149);
or U10204 (N_10204,N_8356,N_6279);
or U10205 (N_10205,N_6056,N_6830);
xor U10206 (N_10206,N_6922,N_6293);
or U10207 (N_10207,N_7552,N_7896);
nor U10208 (N_10208,N_7831,N_6635);
xor U10209 (N_10209,N_6797,N_8502);
or U10210 (N_10210,N_7939,N_8538);
xnor U10211 (N_10211,N_7522,N_6998);
nand U10212 (N_10212,N_6023,N_6726);
nand U10213 (N_10213,N_6951,N_8084);
nand U10214 (N_10214,N_6578,N_8569);
nor U10215 (N_10215,N_8242,N_7229);
and U10216 (N_10216,N_7235,N_8383);
nor U10217 (N_10217,N_7009,N_8567);
xor U10218 (N_10218,N_7298,N_8703);
nor U10219 (N_10219,N_6111,N_7191);
or U10220 (N_10220,N_6681,N_6919);
nor U10221 (N_10221,N_7668,N_6073);
nor U10222 (N_10222,N_6450,N_7893);
xnor U10223 (N_10223,N_7287,N_7450);
and U10224 (N_10224,N_7167,N_6723);
or U10225 (N_10225,N_7107,N_6406);
and U10226 (N_10226,N_7010,N_8620);
nand U10227 (N_10227,N_6567,N_6230);
or U10228 (N_10228,N_8146,N_7797);
nand U10229 (N_10229,N_8317,N_7331);
nor U10230 (N_10230,N_7863,N_6101);
and U10231 (N_10231,N_8400,N_7714);
or U10232 (N_10232,N_6181,N_8269);
xnor U10233 (N_10233,N_7041,N_8178);
nor U10234 (N_10234,N_7507,N_6445);
and U10235 (N_10235,N_8205,N_8468);
and U10236 (N_10236,N_7658,N_8724);
nor U10237 (N_10237,N_6746,N_6497);
nand U10238 (N_10238,N_8546,N_7571);
nor U10239 (N_10239,N_8363,N_6496);
or U10240 (N_10240,N_6675,N_7048);
nand U10241 (N_10241,N_7124,N_8636);
xnor U10242 (N_10242,N_8743,N_7095);
and U10243 (N_10243,N_6236,N_7220);
xor U10244 (N_10244,N_6373,N_8977);
xnor U10245 (N_10245,N_6595,N_6076);
nor U10246 (N_10246,N_7194,N_7231);
or U10247 (N_10247,N_8898,N_6585);
nand U10248 (N_10248,N_7276,N_6601);
or U10249 (N_10249,N_6309,N_6140);
nor U10250 (N_10250,N_7855,N_7265);
or U10251 (N_10251,N_6169,N_7966);
and U10252 (N_10252,N_8498,N_6482);
nor U10253 (N_10253,N_8506,N_7984);
and U10254 (N_10254,N_6906,N_7988);
and U10255 (N_10255,N_6534,N_7389);
nand U10256 (N_10256,N_8132,N_8903);
xor U10257 (N_10257,N_8821,N_8422);
and U10258 (N_10258,N_7332,N_8952);
and U10259 (N_10259,N_6761,N_7649);
xor U10260 (N_10260,N_6606,N_7857);
xnor U10261 (N_10261,N_7142,N_7650);
xnor U10262 (N_10262,N_6363,N_6051);
nand U10263 (N_10263,N_8959,N_6548);
or U10264 (N_10264,N_7876,N_6256);
nand U10265 (N_10265,N_8370,N_8698);
xnor U10266 (N_10266,N_8194,N_8373);
and U10267 (N_10267,N_8609,N_6856);
or U10268 (N_10268,N_6499,N_6964);
xnor U10269 (N_10269,N_6954,N_8717);
or U10270 (N_10270,N_6294,N_6170);
nor U10271 (N_10271,N_8360,N_6662);
and U10272 (N_10272,N_7025,N_6284);
xnor U10273 (N_10273,N_6966,N_6778);
and U10274 (N_10274,N_7676,N_6401);
and U10275 (N_10275,N_8635,N_8893);
nor U10276 (N_10276,N_7072,N_7120);
xor U10277 (N_10277,N_6332,N_7424);
nand U10278 (N_10278,N_8757,N_6502);
or U10279 (N_10279,N_6741,N_7543);
nor U10280 (N_10280,N_6572,N_8556);
nor U10281 (N_10281,N_7865,N_8064);
or U10282 (N_10282,N_8574,N_6019);
nor U10283 (N_10283,N_8344,N_8435);
and U10284 (N_10284,N_6161,N_8102);
nor U10285 (N_10285,N_7247,N_6613);
nand U10286 (N_10286,N_7322,N_8650);
and U10287 (N_10287,N_8234,N_8293);
xnor U10288 (N_10288,N_8911,N_7820);
and U10289 (N_10289,N_8032,N_6949);
or U10290 (N_10290,N_7665,N_8075);
nor U10291 (N_10291,N_8668,N_6716);
nor U10292 (N_10292,N_7164,N_6244);
xnor U10293 (N_10293,N_8822,N_8616);
or U10294 (N_10294,N_8303,N_8892);
nand U10295 (N_10295,N_8289,N_8999);
and U10296 (N_10296,N_8895,N_7494);
nor U10297 (N_10297,N_7622,N_7673);
nor U10298 (N_10298,N_8699,N_8060);
and U10299 (N_10299,N_7669,N_8848);
or U10300 (N_10300,N_6248,N_7692);
nor U10301 (N_10301,N_7093,N_7201);
xor U10302 (N_10302,N_6883,N_8118);
nor U10303 (N_10303,N_7427,N_6518);
nand U10304 (N_10304,N_7761,N_6473);
and U10305 (N_10305,N_8483,N_6420);
nand U10306 (N_10306,N_6719,N_7531);
nor U10307 (N_10307,N_6936,N_7709);
nand U10308 (N_10308,N_8403,N_6753);
nand U10309 (N_10309,N_8310,N_7793);
nand U10310 (N_10310,N_8906,N_8480);
xor U10311 (N_10311,N_6866,N_8018);
or U10312 (N_10312,N_7678,N_6366);
or U10313 (N_10313,N_8566,N_7428);
nand U10314 (N_10314,N_8097,N_7144);
or U10315 (N_10315,N_8979,N_6061);
xnor U10316 (N_10316,N_6812,N_8464);
or U10317 (N_10317,N_8646,N_7621);
or U10318 (N_10318,N_8803,N_8792);
nand U10319 (N_10319,N_7539,N_8536);
and U10320 (N_10320,N_6216,N_7660);
and U10321 (N_10321,N_7772,N_6996);
and U10322 (N_10322,N_8807,N_6569);
nor U10323 (N_10323,N_6689,N_6762);
nor U10324 (N_10324,N_7903,N_7596);
xor U10325 (N_10325,N_6805,N_8209);
or U10326 (N_10326,N_6688,N_7613);
nand U10327 (N_10327,N_8221,N_7073);
or U10328 (N_10328,N_6777,N_6628);
xnor U10329 (N_10329,N_7047,N_8791);
xor U10330 (N_10330,N_6201,N_7341);
nor U10331 (N_10331,N_6853,N_8398);
nor U10332 (N_10332,N_6707,N_7212);
nor U10333 (N_10333,N_8741,N_6227);
nor U10334 (N_10334,N_7439,N_7777);
and U10335 (N_10335,N_8695,N_7155);
and U10336 (N_10336,N_8956,N_8788);
and U10337 (N_10337,N_7616,N_8006);
xnor U10338 (N_10338,N_7614,N_6584);
or U10339 (N_10339,N_8173,N_8798);
nand U10340 (N_10340,N_7576,N_6444);
xor U10341 (N_10341,N_8968,N_8939);
or U10342 (N_10342,N_7113,N_7030);
or U10343 (N_10343,N_7767,N_8748);
and U10344 (N_10344,N_8058,N_8190);
or U10345 (N_10345,N_8980,N_7254);
or U10346 (N_10346,N_7460,N_6243);
xor U10347 (N_10347,N_6296,N_7572);
nor U10348 (N_10348,N_8730,N_8023);
nor U10349 (N_10349,N_8081,N_6269);
or U10350 (N_10350,N_8862,N_8524);
xor U10351 (N_10351,N_6960,N_7375);
or U10352 (N_10352,N_8229,N_8865);
and U10353 (N_10353,N_7267,N_6682);
or U10354 (N_10354,N_6252,N_6361);
xnor U10355 (N_10355,N_6036,N_6152);
nor U10356 (N_10356,N_7157,N_8184);
or U10357 (N_10357,N_8875,N_8787);
nor U10358 (N_10358,N_8320,N_8912);
nor U10359 (N_10359,N_7633,N_6511);
and U10360 (N_10360,N_7985,N_7273);
and U10361 (N_10361,N_6316,N_7990);
or U10362 (N_10362,N_8342,N_6266);
nand U10363 (N_10363,N_6202,N_6834);
nand U10364 (N_10364,N_7457,N_7498);
nand U10365 (N_10365,N_8676,N_6879);
nand U10366 (N_10366,N_7869,N_6016);
nor U10367 (N_10367,N_7573,N_7765);
xor U10368 (N_10368,N_7334,N_6629);
nor U10369 (N_10369,N_8472,N_7619);
nand U10370 (N_10370,N_8411,N_8639);
nand U10371 (N_10371,N_6265,N_6844);
or U10372 (N_10372,N_8066,N_8876);
and U10373 (N_10373,N_7737,N_6074);
and U10374 (N_10374,N_8612,N_8182);
xnor U10375 (N_10375,N_6514,N_6878);
xor U10376 (N_10376,N_7555,N_6346);
or U10377 (N_10377,N_7748,N_8801);
and U10378 (N_10378,N_7687,N_7690);
or U10379 (N_10379,N_6031,N_7038);
nand U10380 (N_10380,N_7434,N_7822);
and U10381 (N_10381,N_8389,N_6642);
or U10382 (N_10382,N_8701,N_7279);
xor U10383 (N_10383,N_8203,N_6231);
nor U10384 (N_10384,N_7550,N_8207);
nand U10385 (N_10385,N_6520,N_6433);
or U10386 (N_10386,N_7154,N_8437);
and U10387 (N_10387,N_6212,N_7824);
and U10388 (N_10388,N_7612,N_7349);
nand U10389 (N_10389,N_6060,N_6116);
nor U10390 (N_10390,N_7138,N_6318);
nor U10391 (N_10391,N_7601,N_8623);
or U10392 (N_10392,N_8869,N_6307);
and U10393 (N_10393,N_7007,N_7899);
and U10394 (N_10394,N_6077,N_6494);
or U10395 (N_10395,N_6582,N_6538);
nand U10396 (N_10396,N_7092,N_8002);
nor U10397 (N_10397,N_6870,N_8512);
nand U10398 (N_10398,N_6786,N_7715);
xnor U10399 (N_10399,N_6154,N_6410);
xor U10400 (N_10400,N_8544,N_8823);
xor U10401 (N_10401,N_8626,N_8087);
and U10402 (N_10402,N_8815,N_7991);
nand U10403 (N_10403,N_8083,N_7788);
nand U10404 (N_10404,N_7262,N_7932);
nor U10405 (N_10405,N_7223,N_6693);
or U10406 (N_10406,N_6412,N_8131);
nand U10407 (N_10407,N_7139,N_6434);
or U10408 (N_10408,N_6666,N_8054);
nor U10409 (N_10409,N_8141,N_8497);
or U10410 (N_10410,N_6492,N_8465);
or U10411 (N_10411,N_8322,N_6250);
nor U10412 (N_10412,N_8661,N_7585);
nand U10413 (N_10413,N_6462,N_6065);
or U10414 (N_10414,N_6770,N_8659);
nor U10415 (N_10415,N_6273,N_6313);
or U10416 (N_10416,N_6358,N_6249);
and U10417 (N_10417,N_6667,N_6714);
nor U10418 (N_10418,N_7661,N_7413);
nand U10419 (N_10419,N_8756,N_6771);
and U10420 (N_10420,N_6207,N_6904);
nor U10421 (N_10421,N_8174,N_7074);
nor U10422 (N_10422,N_6465,N_8974);
or U10423 (N_10423,N_7381,N_6418);
nor U10424 (N_10424,N_7176,N_6913);
nor U10425 (N_10425,N_6149,N_7946);
nor U10426 (N_10426,N_8534,N_8277);
xor U10427 (N_10427,N_7499,N_7598);
and U10428 (N_10428,N_7631,N_6419);
xnor U10429 (N_10429,N_6135,N_7147);
xnor U10430 (N_10430,N_7134,N_6128);
and U10431 (N_10431,N_7377,N_6522);
and U10432 (N_10432,N_6011,N_7099);
or U10433 (N_10433,N_8366,N_7972);
xnor U10434 (N_10434,N_6887,N_7653);
and U10435 (N_10435,N_8038,N_7078);
xor U10436 (N_10436,N_7396,N_6916);
or U10437 (N_10437,N_6861,N_8859);
xor U10438 (N_10438,N_7799,N_7936);
nor U10439 (N_10439,N_6139,N_8708);
or U10440 (N_10440,N_8867,N_7075);
nand U10441 (N_10441,N_7710,N_7004);
nand U10442 (N_10442,N_6874,N_6013);
nor U10443 (N_10443,N_7118,N_7579);
and U10444 (N_10444,N_7608,N_8063);
or U10445 (N_10445,N_8897,N_6593);
or U10446 (N_10446,N_6359,N_7282);
nand U10447 (N_10447,N_6387,N_7051);
or U10448 (N_10448,N_7724,N_7733);
and U10449 (N_10449,N_7497,N_8096);
nor U10450 (N_10450,N_7881,N_6143);
nand U10451 (N_10451,N_6325,N_6678);
xnor U10452 (N_10452,N_6087,N_8213);
or U10453 (N_10453,N_8818,N_7839);
and U10454 (N_10454,N_7705,N_7401);
xnor U10455 (N_10455,N_8726,N_7578);
or U10456 (N_10456,N_7077,N_7293);
nor U10457 (N_10457,N_8053,N_8432);
or U10458 (N_10458,N_8925,N_7076);
nand U10459 (N_10459,N_8041,N_6937);
or U10460 (N_10460,N_7177,N_6159);
and U10461 (N_10461,N_7597,N_6813);
nor U10462 (N_10462,N_8286,N_7747);
or U10463 (N_10463,N_6205,N_7902);
nor U10464 (N_10464,N_6175,N_7335);
and U10465 (N_10465,N_8022,N_6108);
or U10466 (N_10466,N_6455,N_6267);
or U10467 (N_10467,N_8949,N_7846);
and U10468 (N_10468,N_7641,N_7624);
and U10469 (N_10469,N_8677,N_6609);
nand U10470 (N_10470,N_7728,N_6136);
nor U10471 (N_10471,N_7395,N_7565);
xnor U10472 (N_10472,N_7241,N_6467);
xnor U10473 (N_10473,N_7840,N_7969);
or U10474 (N_10474,N_6942,N_7634);
and U10475 (N_10475,N_6341,N_8507);
xor U10476 (N_10476,N_7385,N_8027);
nand U10477 (N_10477,N_8279,N_8428);
xor U10478 (N_10478,N_6055,N_6469);
and U10479 (N_10479,N_7145,N_6633);
nand U10480 (N_10480,N_6370,N_7987);
xnor U10481 (N_10481,N_8550,N_7307);
nand U10482 (N_10482,N_7627,N_8232);
nand U10483 (N_10483,N_7474,N_6768);
nand U10484 (N_10484,N_7515,N_8648);
and U10485 (N_10485,N_6162,N_8423);
or U10486 (N_10486,N_7405,N_8657);
xnor U10487 (N_10487,N_6926,N_8901);
and U10488 (N_10488,N_8306,N_7534);
nor U10489 (N_10489,N_8156,N_6989);
or U10490 (N_10490,N_8907,N_8688);
or U10491 (N_10491,N_8033,N_8257);
and U10492 (N_10492,N_6630,N_8749);
or U10493 (N_10493,N_6468,N_8838);
and U10494 (N_10494,N_6758,N_7738);
xnor U10495 (N_10495,N_7853,N_6799);
xnor U10496 (N_10496,N_6368,N_6134);
nor U10497 (N_10497,N_7628,N_7490);
nand U10498 (N_10498,N_7629,N_7829);
nand U10499 (N_10499,N_6182,N_7354);
or U10500 (N_10500,N_8889,N_8663);
nand U10501 (N_10501,N_8902,N_7541);
and U10502 (N_10502,N_7141,N_8862);
nor U10503 (N_10503,N_8093,N_6840);
and U10504 (N_10504,N_8169,N_8472);
nor U10505 (N_10505,N_6189,N_8064);
nor U10506 (N_10506,N_7019,N_8486);
nor U10507 (N_10507,N_7930,N_7190);
or U10508 (N_10508,N_7781,N_6237);
nand U10509 (N_10509,N_8789,N_6748);
and U10510 (N_10510,N_7146,N_7747);
xnor U10511 (N_10511,N_6449,N_7412);
or U10512 (N_10512,N_8517,N_8412);
xor U10513 (N_10513,N_7047,N_8098);
nor U10514 (N_10514,N_7411,N_7178);
xor U10515 (N_10515,N_7580,N_7565);
xnor U10516 (N_10516,N_8874,N_7776);
xnor U10517 (N_10517,N_6987,N_7655);
xnor U10518 (N_10518,N_6407,N_6498);
and U10519 (N_10519,N_6028,N_6285);
nor U10520 (N_10520,N_7467,N_7426);
or U10521 (N_10521,N_8930,N_6563);
nor U10522 (N_10522,N_6365,N_6655);
nor U10523 (N_10523,N_6488,N_6326);
xnor U10524 (N_10524,N_8412,N_7725);
nand U10525 (N_10525,N_6192,N_6297);
nand U10526 (N_10526,N_7480,N_7534);
nor U10527 (N_10527,N_6367,N_7201);
xnor U10528 (N_10528,N_7697,N_6615);
or U10529 (N_10529,N_7797,N_6572);
xnor U10530 (N_10530,N_6569,N_6940);
or U10531 (N_10531,N_8510,N_6675);
or U10532 (N_10532,N_6613,N_6064);
xnor U10533 (N_10533,N_7777,N_6066);
nand U10534 (N_10534,N_7713,N_6107);
nand U10535 (N_10535,N_7168,N_7749);
nor U10536 (N_10536,N_7022,N_7048);
xnor U10537 (N_10537,N_6052,N_7573);
xnor U10538 (N_10538,N_6482,N_6013);
nand U10539 (N_10539,N_6486,N_8832);
nor U10540 (N_10540,N_6320,N_6416);
nand U10541 (N_10541,N_8049,N_7002);
nand U10542 (N_10542,N_7261,N_8711);
xnor U10543 (N_10543,N_7552,N_6137);
xor U10544 (N_10544,N_8105,N_8104);
xor U10545 (N_10545,N_6938,N_6897);
and U10546 (N_10546,N_7821,N_8493);
nand U10547 (N_10547,N_7965,N_8602);
nand U10548 (N_10548,N_7888,N_6162);
xnor U10549 (N_10549,N_7761,N_8634);
or U10550 (N_10550,N_7782,N_6099);
nand U10551 (N_10551,N_6599,N_8936);
nand U10552 (N_10552,N_8059,N_6538);
nor U10553 (N_10553,N_6306,N_6007);
or U10554 (N_10554,N_7533,N_8646);
or U10555 (N_10555,N_7632,N_7293);
nand U10556 (N_10556,N_7876,N_7462);
xnor U10557 (N_10557,N_8959,N_8992);
or U10558 (N_10558,N_6894,N_7316);
nor U10559 (N_10559,N_6982,N_6745);
xor U10560 (N_10560,N_7869,N_6583);
and U10561 (N_10561,N_8535,N_8883);
and U10562 (N_10562,N_6819,N_7938);
and U10563 (N_10563,N_6059,N_8252);
nand U10564 (N_10564,N_6311,N_6167);
xor U10565 (N_10565,N_6005,N_6143);
and U10566 (N_10566,N_8479,N_8069);
nor U10567 (N_10567,N_7347,N_6559);
nand U10568 (N_10568,N_6269,N_6520);
xnor U10569 (N_10569,N_8212,N_6362);
nor U10570 (N_10570,N_7369,N_7473);
and U10571 (N_10571,N_7526,N_7772);
xor U10572 (N_10572,N_7328,N_6298);
xor U10573 (N_10573,N_8808,N_6004);
nor U10574 (N_10574,N_7768,N_6248);
nor U10575 (N_10575,N_6306,N_6571);
and U10576 (N_10576,N_6961,N_7797);
or U10577 (N_10577,N_7078,N_8118);
and U10578 (N_10578,N_8191,N_8451);
xnor U10579 (N_10579,N_6447,N_8492);
or U10580 (N_10580,N_6992,N_6834);
nand U10581 (N_10581,N_8626,N_6233);
and U10582 (N_10582,N_8747,N_6854);
nor U10583 (N_10583,N_7290,N_8394);
or U10584 (N_10584,N_7362,N_7691);
xor U10585 (N_10585,N_7391,N_6675);
nand U10586 (N_10586,N_7124,N_7777);
nand U10587 (N_10587,N_6829,N_8744);
nor U10588 (N_10588,N_7840,N_8234);
or U10589 (N_10589,N_6666,N_7322);
and U10590 (N_10590,N_8495,N_7787);
or U10591 (N_10591,N_8750,N_7481);
and U10592 (N_10592,N_8274,N_7371);
and U10593 (N_10593,N_7147,N_7583);
and U10594 (N_10594,N_7305,N_7275);
or U10595 (N_10595,N_6189,N_7714);
and U10596 (N_10596,N_6786,N_6482);
nor U10597 (N_10597,N_7469,N_6437);
nor U10598 (N_10598,N_6509,N_7026);
nor U10599 (N_10599,N_6412,N_8174);
and U10600 (N_10600,N_7240,N_8892);
nand U10601 (N_10601,N_8495,N_6809);
and U10602 (N_10602,N_6551,N_7538);
nor U10603 (N_10603,N_7428,N_7115);
and U10604 (N_10604,N_7132,N_7224);
nand U10605 (N_10605,N_8944,N_6977);
nand U10606 (N_10606,N_7941,N_8469);
nor U10607 (N_10607,N_6200,N_6118);
or U10608 (N_10608,N_6842,N_8760);
nor U10609 (N_10609,N_8940,N_7475);
and U10610 (N_10610,N_8938,N_6149);
and U10611 (N_10611,N_8426,N_8749);
or U10612 (N_10612,N_7516,N_6053);
and U10613 (N_10613,N_6366,N_7362);
or U10614 (N_10614,N_8349,N_6869);
or U10615 (N_10615,N_6315,N_6563);
and U10616 (N_10616,N_8341,N_8475);
xnor U10617 (N_10617,N_6867,N_8701);
xnor U10618 (N_10618,N_6754,N_8660);
or U10619 (N_10619,N_6217,N_6167);
xnor U10620 (N_10620,N_7766,N_8115);
and U10621 (N_10621,N_7014,N_7019);
nand U10622 (N_10622,N_7742,N_6465);
or U10623 (N_10623,N_6823,N_8727);
or U10624 (N_10624,N_7581,N_8357);
nor U10625 (N_10625,N_7485,N_7034);
nor U10626 (N_10626,N_8437,N_6845);
nor U10627 (N_10627,N_6689,N_8789);
and U10628 (N_10628,N_8110,N_6703);
xor U10629 (N_10629,N_6327,N_7955);
and U10630 (N_10630,N_7766,N_8688);
and U10631 (N_10631,N_6582,N_7852);
xnor U10632 (N_10632,N_6575,N_7918);
xor U10633 (N_10633,N_6260,N_7229);
or U10634 (N_10634,N_8425,N_7907);
and U10635 (N_10635,N_6666,N_8697);
nand U10636 (N_10636,N_6673,N_7179);
xor U10637 (N_10637,N_7839,N_7295);
and U10638 (N_10638,N_8289,N_8788);
or U10639 (N_10639,N_8924,N_7360);
nand U10640 (N_10640,N_6435,N_8817);
and U10641 (N_10641,N_7401,N_8061);
xor U10642 (N_10642,N_6404,N_8595);
or U10643 (N_10643,N_7000,N_8639);
nor U10644 (N_10644,N_7725,N_7484);
xor U10645 (N_10645,N_8740,N_7922);
nand U10646 (N_10646,N_8586,N_7323);
nand U10647 (N_10647,N_8386,N_6671);
nor U10648 (N_10648,N_7187,N_8830);
nor U10649 (N_10649,N_8499,N_6662);
nor U10650 (N_10650,N_8169,N_6213);
xor U10651 (N_10651,N_8594,N_7325);
or U10652 (N_10652,N_8743,N_7492);
nor U10653 (N_10653,N_8667,N_8128);
xor U10654 (N_10654,N_7049,N_6866);
nand U10655 (N_10655,N_7923,N_6814);
or U10656 (N_10656,N_7254,N_7660);
or U10657 (N_10657,N_6179,N_7167);
nand U10658 (N_10658,N_7338,N_6041);
xor U10659 (N_10659,N_6937,N_7054);
or U10660 (N_10660,N_8147,N_7885);
nor U10661 (N_10661,N_6203,N_6661);
or U10662 (N_10662,N_7729,N_6647);
nand U10663 (N_10663,N_6303,N_8183);
xnor U10664 (N_10664,N_8429,N_6749);
or U10665 (N_10665,N_7735,N_6121);
xnor U10666 (N_10666,N_7751,N_6597);
xnor U10667 (N_10667,N_7060,N_6074);
and U10668 (N_10668,N_6546,N_6259);
and U10669 (N_10669,N_7829,N_6132);
xor U10670 (N_10670,N_8695,N_7108);
or U10671 (N_10671,N_8169,N_6454);
nand U10672 (N_10672,N_7526,N_6116);
nand U10673 (N_10673,N_7201,N_8142);
nand U10674 (N_10674,N_8095,N_8351);
xnor U10675 (N_10675,N_6099,N_6783);
nand U10676 (N_10676,N_8105,N_8411);
nand U10677 (N_10677,N_7159,N_7712);
xnor U10678 (N_10678,N_8065,N_7465);
xor U10679 (N_10679,N_7467,N_8655);
nor U10680 (N_10680,N_7301,N_6518);
and U10681 (N_10681,N_6694,N_7006);
nor U10682 (N_10682,N_8219,N_8986);
and U10683 (N_10683,N_8091,N_7505);
nand U10684 (N_10684,N_6722,N_8830);
nand U10685 (N_10685,N_6725,N_6263);
nand U10686 (N_10686,N_6771,N_8248);
nand U10687 (N_10687,N_8866,N_7055);
xor U10688 (N_10688,N_6191,N_6115);
nand U10689 (N_10689,N_6181,N_8097);
and U10690 (N_10690,N_6827,N_8346);
and U10691 (N_10691,N_6934,N_7814);
nor U10692 (N_10692,N_8239,N_6616);
and U10693 (N_10693,N_6906,N_6756);
xnor U10694 (N_10694,N_7993,N_7338);
xnor U10695 (N_10695,N_8834,N_6806);
xor U10696 (N_10696,N_7843,N_8021);
nand U10697 (N_10697,N_8681,N_7165);
nand U10698 (N_10698,N_7504,N_6601);
xnor U10699 (N_10699,N_6496,N_8468);
and U10700 (N_10700,N_6415,N_6304);
and U10701 (N_10701,N_8849,N_8777);
or U10702 (N_10702,N_8365,N_8310);
or U10703 (N_10703,N_7428,N_7299);
or U10704 (N_10704,N_7942,N_7474);
nand U10705 (N_10705,N_6026,N_8769);
nor U10706 (N_10706,N_7235,N_7814);
or U10707 (N_10707,N_7973,N_7806);
and U10708 (N_10708,N_7435,N_6406);
or U10709 (N_10709,N_6386,N_8353);
or U10710 (N_10710,N_6173,N_6837);
nand U10711 (N_10711,N_6151,N_8944);
or U10712 (N_10712,N_6869,N_7244);
or U10713 (N_10713,N_8978,N_7041);
nor U10714 (N_10714,N_8099,N_8060);
xor U10715 (N_10715,N_8829,N_8030);
xnor U10716 (N_10716,N_6756,N_7690);
nor U10717 (N_10717,N_6974,N_7467);
and U10718 (N_10718,N_7715,N_6306);
and U10719 (N_10719,N_7413,N_8609);
xor U10720 (N_10720,N_6274,N_6197);
nor U10721 (N_10721,N_7400,N_7133);
and U10722 (N_10722,N_7139,N_7422);
or U10723 (N_10723,N_7711,N_8892);
xnor U10724 (N_10724,N_8665,N_8534);
nand U10725 (N_10725,N_7967,N_8543);
and U10726 (N_10726,N_8535,N_7962);
and U10727 (N_10727,N_8970,N_8051);
nand U10728 (N_10728,N_7997,N_6579);
nand U10729 (N_10729,N_8614,N_8431);
nand U10730 (N_10730,N_6331,N_6782);
and U10731 (N_10731,N_8783,N_6875);
and U10732 (N_10732,N_7973,N_7527);
nand U10733 (N_10733,N_6035,N_8204);
and U10734 (N_10734,N_7558,N_6979);
xnor U10735 (N_10735,N_8065,N_8090);
nand U10736 (N_10736,N_7483,N_8835);
xnor U10737 (N_10737,N_8510,N_8473);
or U10738 (N_10738,N_8725,N_6512);
xor U10739 (N_10739,N_8949,N_7643);
xnor U10740 (N_10740,N_6705,N_8391);
nand U10741 (N_10741,N_7293,N_8180);
nand U10742 (N_10742,N_7952,N_8877);
and U10743 (N_10743,N_7319,N_6445);
or U10744 (N_10744,N_7811,N_7986);
nand U10745 (N_10745,N_8063,N_6964);
xnor U10746 (N_10746,N_6217,N_7042);
xnor U10747 (N_10747,N_8195,N_8274);
and U10748 (N_10748,N_8930,N_7805);
nor U10749 (N_10749,N_7772,N_8912);
or U10750 (N_10750,N_7360,N_6336);
and U10751 (N_10751,N_8313,N_6826);
or U10752 (N_10752,N_6172,N_8016);
or U10753 (N_10753,N_6579,N_6348);
and U10754 (N_10754,N_8057,N_8780);
xnor U10755 (N_10755,N_7333,N_8572);
or U10756 (N_10756,N_6122,N_7627);
nand U10757 (N_10757,N_6845,N_8245);
nor U10758 (N_10758,N_8801,N_8599);
nand U10759 (N_10759,N_8876,N_6058);
nand U10760 (N_10760,N_8671,N_8502);
nor U10761 (N_10761,N_8557,N_8604);
nand U10762 (N_10762,N_6865,N_7246);
and U10763 (N_10763,N_8914,N_8067);
nand U10764 (N_10764,N_7319,N_8842);
xnor U10765 (N_10765,N_7248,N_7897);
nor U10766 (N_10766,N_6810,N_6296);
xnor U10767 (N_10767,N_8780,N_7736);
nor U10768 (N_10768,N_7260,N_8976);
or U10769 (N_10769,N_6021,N_8702);
xor U10770 (N_10770,N_8347,N_7503);
nor U10771 (N_10771,N_6935,N_8413);
or U10772 (N_10772,N_8494,N_8326);
nand U10773 (N_10773,N_6585,N_6732);
nand U10774 (N_10774,N_8286,N_8183);
nor U10775 (N_10775,N_6629,N_7092);
or U10776 (N_10776,N_8421,N_6097);
nor U10777 (N_10777,N_7552,N_8157);
nand U10778 (N_10778,N_6262,N_8396);
nand U10779 (N_10779,N_6563,N_8095);
xnor U10780 (N_10780,N_7925,N_7393);
nand U10781 (N_10781,N_7756,N_7550);
or U10782 (N_10782,N_6021,N_6519);
nor U10783 (N_10783,N_7151,N_6432);
or U10784 (N_10784,N_6801,N_6606);
nand U10785 (N_10785,N_8716,N_7491);
nand U10786 (N_10786,N_6364,N_7386);
xor U10787 (N_10787,N_8946,N_6672);
nand U10788 (N_10788,N_8368,N_7252);
nor U10789 (N_10789,N_7013,N_6967);
nand U10790 (N_10790,N_8500,N_6983);
nand U10791 (N_10791,N_8063,N_8937);
nor U10792 (N_10792,N_8793,N_6027);
nand U10793 (N_10793,N_8680,N_8162);
nand U10794 (N_10794,N_7222,N_6723);
xor U10795 (N_10795,N_7690,N_7824);
and U10796 (N_10796,N_7258,N_7221);
and U10797 (N_10797,N_7307,N_7895);
nor U10798 (N_10798,N_6774,N_7674);
and U10799 (N_10799,N_8172,N_8681);
and U10800 (N_10800,N_8842,N_8662);
nand U10801 (N_10801,N_8720,N_6273);
or U10802 (N_10802,N_6609,N_8021);
nand U10803 (N_10803,N_8769,N_6944);
nor U10804 (N_10804,N_7108,N_7562);
xor U10805 (N_10805,N_7008,N_7702);
nor U10806 (N_10806,N_8136,N_6508);
xnor U10807 (N_10807,N_6051,N_7024);
xnor U10808 (N_10808,N_7455,N_7874);
nor U10809 (N_10809,N_6667,N_6212);
nand U10810 (N_10810,N_6451,N_6490);
xor U10811 (N_10811,N_8698,N_8697);
and U10812 (N_10812,N_8928,N_6604);
or U10813 (N_10813,N_8832,N_7802);
nand U10814 (N_10814,N_6080,N_8609);
xor U10815 (N_10815,N_8801,N_7010);
nor U10816 (N_10816,N_8928,N_7314);
and U10817 (N_10817,N_6164,N_7941);
or U10818 (N_10818,N_8166,N_7851);
nand U10819 (N_10819,N_8582,N_7118);
xor U10820 (N_10820,N_7863,N_6030);
or U10821 (N_10821,N_6815,N_7124);
xnor U10822 (N_10822,N_8113,N_6295);
or U10823 (N_10823,N_8261,N_8776);
nand U10824 (N_10824,N_7297,N_6652);
and U10825 (N_10825,N_8806,N_8821);
and U10826 (N_10826,N_6958,N_7740);
nand U10827 (N_10827,N_6591,N_7673);
and U10828 (N_10828,N_6322,N_6880);
or U10829 (N_10829,N_7256,N_6044);
nor U10830 (N_10830,N_7043,N_8654);
xnor U10831 (N_10831,N_8846,N_8827);
nor U10832 (N_10832,N_8953,N_6964);
and U10833 (N_10833,N_6739,N_6856);
nand U10834 (N_10834,N_7198,N_8889);
nor U10835 (N_10835,N_6706,N_6088);
and U10836 (N_10836,N_7814,N_7993);
xnor U10837 (N_10837,N_7981,N_8380);
nand U10838 (N_10838,N_6580,N_7177);
nand U10839 (N_10839,N_7105,N_6855);
xor U10840 (N_10840,N_6954,N_7860);
nand U10841 (N_10841,N_7795,N_7586);
or U10842 (N_10842,N_7646,N_8143);
or U10843 (N_10843,N_8726,N_7861);
and U10844 (N_10844,N_6153,N_8459);
and U10845 (N_10845,N_8642,N_7892);
nand U10846 (N_10846,N_7160,N_8730);
and U10847 (N_10847,N_7106,N_7180);
or U10848 (N_10848,N_7451,N_6089);
nand U10849 (N_10849,N_8307,N_6541);
nand U10850 (N_10850,N_6263,N_6077);
or U10851 (N_10851,N_7365,N_6074);
xnor U10852 (N_10852,N_7895,N_7450);
nor U10853 (N_10853,N_8337,N_7023);
or U10854 (N_10854,N_8616,N_8509);
nor U10855 (N_10855,N_6858,N_8673);
or U10856 (N_10856,N_8589,N_7276);
xor U10857 (N_10857,N_8323,N_7710);
nor U10858 (N_10858,N_6141,N_8671);
nand U10859 (N_10859,N_6528,N_8911);
and U10860 (N_10860,N_7557,N_6105);
nor U10861 (N_10861,N_8951,N_8433);
or U10862 (N_10862,N_7173,N_6963);
xnor U10863 (N_10863,N_7327,N_7701);
nor U10864 (N_10864,N_6383,N_8416);
and U10865 (N_10865,N_6992,N_7702);
nand U10866 (N_10866,N_8497,N_8511);
xnor U10867 (N_10867,N_6290,N_8095);
or U10868 (N_10868,N_7630,N_7163);
and U10869 (N_10869,N_6369,N_6065);
nand U10870 (N_10870,N_6445,N_7551);
and U10871 (N_10871,N_6296,N_8339);
xnor U10872 (N_10872,N_6797,N_6981);
nand U10873 (N_10873,N_7286,N_6320);
and U10874 (N_10874,N_8418,N_8818);
xor U10875 (N_10875,N_7808,N_8887);
and U10876 (N_10876,N_8584,N_7956);
or U10877 (N_10877,N_7739,N_8747);
and U10878 (N_10878,N_8552,N_6809);
nand U10879 (N_10879,N_7928,N_8974);
and U10880 (N_10880,N_8511,N_6049);
nand U10881 (N_10881,N_8093,N_7363);
and U10882 (N_10882,N_7398,N_6575);
and U10883 (N_10883,N_7598,N_8526);
and U10884 (N_10884,N_8483,N_6535);
nand U10885 (N_10885,N_8800,N_8530);
or U10886 (N_10886,N_7772,N_8228);
or U10887 (N_10887,N_7754,N_6810);
nor U10888 (N_10888,N_8328,N_8683);
nand U10889 (N_10889,N_7669,N_7885);
or U10890 (N_10890,N_6745,N_6394);
nand U10891 (N_10891,N_8336,N_7333);
nand U10892 (N_10892,N_7382,N_7838);
or U10893 (N_10893,N_6410,N_8649);
and U10894 (N_10894,N_8742,N_6096);
nand U10895 (N_10895,N_8744,N_8701);
nand U10896 (N_10896,N_7514,N_8797);
nor U10897 (N_10897,N_8799,N_8855);
or U10898 (N_10898,N_6063,N_7767);
nor U10899 (N_10899,N_7536,N_6107);
nand U10900 (N_10900,N_6303,N_7829);
and U10901 (N_10901,N_7714,N_6046);
or U10902 (N_10902,N_7266,N_8968);
xnor U10903 (N_10903,N_8807,N_7612);
nand U10904 (N_10904,N_6647,N_7416);
xnor U10905 (N_10905,N_8318,N_7217);
nand U10906 (N_10906,N_6096,N_8401);
xor U10907 (N_10907,N_8982,N_8895);
nor U10908 (N_10908,N_6454,N_6648);
nor U10909 (N_10909,N_8184,N_7512);
xnor U10910 (N_10910,N_7157,N_8706);
nor U10911 (N_10911,N_8355,N_7558);
nand U10912 (N_10912,N_7127,N_6931);
or U10913 (N_10913,N_7718,N_7845);
nand U10914 (N_10914,N_6420,N_6085);
and U10915 (N_10915,N_6669,N_6741);
and U10916 (N_10916,N_7970,N_7993);
or U10917 (N_10917,N_7116,N_6472);
and U10918 (N_10918,N_7864,N_7681);
nor U10919 (N_10919,N_6581,N_6216);
or U10920 (N_10920,N_7883,N_7104);
and U10921 (N_10921,N_8889,N_8295);
and U10922 (N_10922,N_6308,N_8541);
or U10923 (N_10923,N_8694,N_6240);
nor U10924 (N_10924,N_7890,N_6632);
nor U10925 (N_10925,N_7002,N_8593);
or U10926 (N_10926,N_7548,N_7595);
nor U10927 (N_10927,N_6525,N_7399);
nand U10928 (N_10928,N_6172,N_6361);
xor U10929 (N_10929,N_7668,N_8965);
nor U10930 (N_10930,N_6201,N_6811);
xnor U10931 (N_10931,N_8645,N_8166);
nor U10932 (N_10932,N_6254,N_6216);
nor U10933 (N_10933,N_6845,N_7087);
nand U10934 (N_10934,N_6872,N_8128);
or U10935 (N_10935,N_7362,N_6606);
and U10936 (N_10936,N_8065,N_6926);
nor U10937 (N_10937,N_7146,N_8785);
or U10938 (N_10938,N_6753,N_7895);
nor U10939 (N_10939,N_7453,N_6124);
nor U10940 (N_10940,N_6150,N_7387);
xor U10941 (N_10941,N_7344,N_7843);
and U10942 (N_10942,N_8886,N_7694);
and U10943 (N_10943,N_6464,N_8199);
or U10944 (N_10944,N_7335,N_7526);
xor U10945 (N_10945,N_8727,N_7580);
xor U10946 (N_10946,N_7520,N_7925);
xor U10947 (N_10947,N_7866,N_6615);
nand U10948 (N_10948,N_6294,N_7839);
nand U10949 (N_10949,N_6506,N_7197);
or U10950 (N_10950,N_6538,N_6721);
xnor U10951 (N_10951,N_6300,N_7418);
nor U10952 (N_10952,N_6875,N_6401);
or U10953 (N_10953,N_7652,N_7387);
nand U10954 (N_10954,N_7873,N_8975);
or U10955 (N_10955,N_7895,N_7491);
and U10956 (N_10956,N_7962,N_6849);
nand U10957 (N_10957,N_8800,N_6943);
xor U10958 (N_10958,N_7856,N_8064);
or U10959 (N_10959,N_6497,N_6294);
xnor U10960 (N_10960,N_6884,N_7519);
xor U10961 (N_10961,N_6169,N_8139);
or U10962 (N_10962,N_6057,N_7944);
xor U10963 (N_10963,N_6425,N_6707);
or U10964 (N_10964,N_8154,N_7302);
and U10965 (N_10965,N_7881,N_8686);
or U10966 (N_10966,N_7189,N_6553);
and U10967 (N_10967,N_8566,N_8409);
nand U10968 (N_10968,N_7007,N_8416);
or U10969 (N_10969,N_7602,N_6985);
nand U10970 (N_10970,N_8892,N_6818);
nor U10971 (N_10971,N_6299,N_6746);
nor U10972 (N_10972,N_8530,N_6007);
nor U10973 (N_10973,N_8854,N_8263);
nor U10974 (N_10974,N_8785,N_7706);
and U10975 (N_10975,N_6292,N_8765);
nand U10976 (N_10976,N_7830,N_6529);
xor U10977 (N_10977,N_6437,N_6830);
and U10978 (N_10978,N_8717,N_8350);
or U10979 (N_10979,N_6962,N_6376);
nor U10980 (N_10980,N_6213,N_8088);
and U10981 (N_10981,N_6164,N_8422);
nand U10982 (N_10982,N_7413,N_6350);
or U10983 (N_10983,N_8630,N_8558);
and U10984 (N_10984,N_8624,N_7661);
nor U10985 (N_10985,N_8075,N_7629);
xor U10986 (N_10986,N_7019,N_8460);
or U10987 (N_10987,N_6862,N_7773);
xnor U10988 (N_10988,N_6120,N_7754);
or U10989 (N_10989,N_8999,N_7669);
and U10990 (N_10990,N_8637,N_8465);
xor U10991 (N_10991,N_6832,N_6206);
nand U10992 (N_10992,N_6051,N_6011);
or U10993 (N_10993,N_6357,N_6777);
or U10994 (N_10994,N_7031,N_8235);
nor U10995 (N_10995,N_6481,N_7002);
nand U10996 (N_10996,N_7159,N_6727);
nor U10997 (N_10997,N_7850,N_7225);
and U10998 (N_10998,N_6517,N_7895);
nor U10999 (N_10999,N_8037,N_8691);
and U11000 (N_11000,N_8299,N_6221);
nor U11001 (N_11001,N_8778,N_8073);
or U11002 (N_11002,N_8564,N_8373);
or U11003 (N_11003,N_6543,N_7501);
xnor U11004 (N_11004,N_8943,N_6785);
or U11005 (N_11005,N_6515,N_6659);
nor U11006 (N_11006,N_6533,N_7186);
nand U11007 (N_11007,N_7536,N_6332);
xnor U11008 (N_11008,N_8052,N_8759);
nand U11009 (N_11009,N_8901,N_6577);
and U11010 (N_11010,N_6442,N_6033);
or U11011 (N_11011,N_7072,N_6924);
or U11012 (N_11012,N_6001,N_6387);
xnor U11013 (N_11013,N_7710,N_6437);
nand U11014 (N_11014,N_6264,N_6401);
xnor U11015 (N_11015,N_6227,N_7972);
nor U11016 (N_11016,N_7966,N_7241);
nand U11017 (N_11017,N_8401,N_6190);
and U11018 (N_11018,N_8008,N_7062);
and U11019 (N_11019,N_7671,N_8172);
nand U11020 (N_11020,N_8122,N_6764);
and U11021 (N_11021,N_6171,N_8982);
xor U11022 (N_11022,N_8552,N_6193);
or U11023 (N_11023,N_7269,N_8607);
xor U11024 (N_11024,N_6520,N_8825);
xnor U11025 (N_11025,N_8406,N_6865);
and U11026 (N_11026,N_7631,N_6339);
nor U11027 (N_11027,N_7048,N_7825);
or U11028 (N_11028,N_8600,N_6780);
nor U11029 (N_11029,N_7927,N_7351);
nor U11030 (N_11030,N_6227,N_7385);
nand U11031 (N_11031,N_7076,N_7081);
or U11032 (N_11032,N_8911,N_8238);
nor U11033 (N_11033,N_7011,N_8711);
nand U11034 (N_11034,N_8168,N_6754);
xnor U11035 (N_11035,N_7093,N_6616);
nand U11036 (N_11036,N_6701,N_6724);
nor U11037 (N_11037,N_6021,N_8124);
xor U11038 (N_11038,N_8576,N_7508);
xnor U11039 (N_11039,N_6951,N_6933);
xnor U11040 (N_11040,N_8730,N_6676);
nor U11041 (N_11041,N_7373,N_8008);
nand U11042 (N_11042,N_8395,N_7347);
nand U11043 (N_11043,N_7510,N_8162);
nor U11044 (N_11044,N_8105,N_6581);
or U11045 (N_11045,N_7590,N_8642);
or U11046 (N_11046,N_7941,N_6407);
xor U11047 (N_11047,N_7223,N_6473);
nor U11048 (N_11048,N_7477,N_8020);
xnor U11049 (N_11049,N_7942,N_7873);
nor U11050 (N_11050,N_8489,N_7523);
or U11051 (N_11051,N_8154,N_8651);
nand U11052 (N_11052,N_8489,N_7536);
or U11053 (N_11053,N_6829,N_6432);
nor U11054 (N_11054,N_7083,N_7491);
or U11055 (N_11055,N_8943,N_6097);
xnor U11056 (N_11056,N_7578,N_8893);
and U11057 (N_11057,N_8596,N_6089);
nand U11058 (N_11058,N_6600,N_6949);
nor U11059 (N_11059,N_8303,N_8291);
nand U11060 (N_11060,N_7493,N_6408);
and U11061 (N_11061,N_7330,N_6787);
nand U11062 (N_11062,N_7499,N_7309);
nand U11063 (N_11063,N_6800,N_6394);
nand U11064 (N_11064,N_8996,N_6586);
nand U11065 (N_11065,N_6043,N_7205);
and U11066 (N_11066,N_7376,N_7266);
xnor U11067 (N_11067,N_6716,N_6401);
or U11068 (N_11068,N_7904,N_6035);
xnor U11069 (N_11069,N_7258,N_7993);
xor U11070 (N_11070,N_8606,N_7029);
or U11071 (N_11071,N_6257,N_7451);
xnor U11072 (N_11072,N_8716,N_8041);
xor U11073 (N_11073,N_6949,N_7447);
or U11074 (N_11074,N_7902,N_6444);
and U11075 (N_11075,N_8160,N_6944);
and U11076 (N_11076,N_6249,N_8766);
or U11077 (N_11077,N_8369,N_8728);
or U11078 (N_11078,N_7700,N_6164);
or U11079 (N_11079,N_6893,N_6334);
and U11080 (N_11080,N_7113,N_8408);
nand U11081 (N_11081,N_8233,N_8222);
and U11082 (N_11082,N_6622,N_6393);
nor U11083 (N_11083,N_6197,N_8312);
nand U11084 (N_11084,N_8981,N_8608);
and U11085 (N_11085,N_8875,N_7247);
nand U11086 (N_11086,N_8172,N_8529);
nor U11087 (N_11087,N_8357,N_8199);
nand U11088 (N_11088,N_8586,N_6433);
nand U11089 (N_11089,N_6456,N_6296);
nor U11090 (N_11090,N_8261,N_7656);
nand U11091 (N_11091,N_8045,N_7685);
and U11092 (N_11092,N_6523,N_7281);
nor U11093 (N_11093,N_8212,N_7920);
nor U11094 (N_11094,N_8974,N_6871);
nor U11095 (N_11095,N_8535,N_7589);
and U11096 (N_11096,N_8288,N_8221);
nor U11097 (N_11097,N_7197,N_7373);
nand U11098 (N_11098,N_7981,N_8815);
nand U11099 (N_11099,N_8714,N_6131);
nor U11100 (N_11100,N_6587,N_6355);
nor U11101 (N_11101,N_7834,N_6505);
or U11102 (N_11102,N_8616,N_7799);
and U11103 (N_11103,N_7374,N_6523);
or U11104 (N_11104,N_7205,N_7438);
xor U11105 (N_11105,N_6625,N_7871);
nand U11106 (N_11106,N_8815,N_6694);
and U11107 (N_11107,N_7522,N_7640);
and U11108 (N_11108,N_8462,N_8756);
or U11109 (N_11109,N_8401,N_8173);
nand U11110 (N_11110,N_7048,N_8670);
and U11111 (N_11111,N_7048,N_8028);
or U11112 (N_11112,N_7426,N_8703);
or U11113 (N_11113,N_6742,N_6573);
nand U11114 (N_11114,N_7486,N_7209);
xor U11115 (N_11115,N_6332,N_8903);
and U11116 (N_11116,N_8841,N_6391);
and U11117 (N_11117,N_6848,N_8807);
nor U11118 (N_11118,N_6997,N_7003);
nand U11119 (N_11119,N_7662,N_7327);
nor U11120 (N_11120,N_7065,N_7078);
xor U11121 (N_11121,N_8423,N_6748);
xor U11122 (N_11122,N_7943,N_7795);
nand U11123 (N_11123,N_8550,N_7736);
nor U11124 (N_11124,N_7252,N_7383);
and U11125 (N_11125,N_8503,N_8777);
nor U11126 (N_11126,N_6785,N_8182);
or U11127 (N_11127,N_8385,N_8295);
or U11128 (N_11128,N_8553,N_7052);
nor U11129 (N_11129,N_7050,N_6619);
nor U11130 (N_11130,N_7065,N_7758);
xnor U11131 (N_11131,N_6329,N_6689);
nand U11132 (N_11132,N_8147,N_6509);
xor U11133 (N_11133,N_7052,N_6628);
and U11134 (N_11134,N_7523,N_6941);
xnor U11135 (N_11135,N_8349,N_7395);
xnor U11136 (N_11136,N_7327,N_8322);
nor U11137 (N_11137,N_6743,N_7134);
or U11138 (N_11138,N_6271,N_8540);
nand U11139 (N_11139,N_7657,N_6966);
or U11140 (N_11140,N_6450,N_7544);
or U11141 (N_11141,N_8465,N_7959);
or U11142 (N_11142,N_6288,N_8985);
nand U11143 (N_11143,N_7219,N_8488);
nor U11144 (N_11144,N_6982,N_7851);
nand U11145 (N_11145,N_7315,N_8165);
or U11146 (N_11146,N_7630,N_8205);
and U11147 (N_11147,N_7893,N_6797);
nor U11148 (N_11148,N_7798,N_8303);
nand U11149 (N_11149,N_6298,N_6236);
or U11150 (N_11150,N_8299,N_6465);
or U11151 (N_11151,N_7410,N_8817);
nor U11152 (N_11152,N_7874,N_6705);
and U11153 (N_11153,N_6602,N_6793);
nand U11154 (N_11154,N_6248,N_8289);
xor U11155 (N_11155,N_6737,N_6453);
and U11156 (N_11156,N_7214,N_7519);
or U11157 (N_11157,N_7459,N_6968);
or U11158 (N_11158,N_8089,N_6719);
nand U11159 (N_11159,N_8094,N_6382);
and U11160 (N_11160,N_7676,N_8229);
or U11161 (N_11161,N_8315,N_7331);
nor U11162 (N_11162,N_6277,N_7827);
nor U11163 (N_11163,N_8906,N_7863);
or U11164 (N_11164,N_7043,N_6589);
and U11165 (N_11165,N_8527,N_7095);
or U11166 (N_11166,N_8181,N_7494);
and U11167 (N_11167,N_7059,N_7282);
nor U11168 (N_11168,N_7503,N_8902);
xnor U11169 (N_11169,N_7768,N_8657);
or U11170 (N_11170,N_8088,N_6006);
xor U11171 (N_11171,N_7958,N_7594);
nand U11172 (N_11172,N_6098,N_6154);
or U11173 (N_11173,N_8233,N_6213);
xor U11174 (N_11174,N_8398,N_6706);
and U11175 (N_11175,N_6443,N_6903);
and U11176 (N_11176,N_6368,N_8054);
or U11177 (N_11177,N_8085,N_7822);
nor U11178 (N_11178,N_7191,N_8260);
xor U11179 (N_11179,N_7323,N_8374);
xor U11180 (N_11180,N_8947,N_8524);
nor U11181 (N_11181,N_7304,N_6159);
or U11182 (N_11182,N_8025,N_7316);
nor U11183 (N_11183,N_7405,N_7303);
xnor U11184 (N_11184,N_7616,N_7454);
and U11185 (N_11185,N_6394,N_6465);
nor U11186 (N_11186,N_7509,N_8678);
nor U11187 (N_11187,N_8849,N_7198);
xor U11188 (N_11188,N_7394,N_6821);
nand U11189 (N_11189,N_8634,N_7568);
or U11190 (N_11190,N_8275,N_6568);
xnor U11191 (N_11191,N_6726,N_8378);
and U11192 (N_11192,N_7653,N_6775);
nand U11193 (N_11193,N_8448,N_6954);
and U11194 (N_11194,N_8424,N_6475);
and U11195 (N_11195,N_8877,N_7083);
xor U11196 (N_11196,N_7236,N_6287);
and U11197 (N_11197,N_7894,N_6059);
nand U11198 (N_11198,N_6307,N_6042);
nand U11199 (N_11199,N_6698,N_6305);
nand U11200 (N_11200,N_7271,N_8900);
or U11201 (N_11201,N_8402,N_8953);
xor U11202 (N_11202,N_8623,N_6444);
nand U11203 (N_11203,N_6353,N_7028);
nand U11204 (N_11204,N_7578,N_7259);
nand U11205 (N_11205,N_6253,N_7773);
nor U11206 (N_11206,N_8444,N_8881);
xnor U11207 (N_11207,N_6365,N_7317);
and U11208 (N_11208,N_6392,N_8707);
nor U11209 (N_11209,N_7337,N_6427);
nand U11210 (N_11210,N_8517,N_8646);
nand U11211 (N_11211,N_7562,N_8989);
or U11212 (N_11212,N_8880,N_7126);
xnor U11213 (N_11213,N_8941,N_6569);
and U11214 (N_11214,N_7921,N_8134);
xor U11215 (N_11215,N_7097,N_7811);
xnor U11216 (N_11216,N_8622,N_6781);
xnor U11217 (N_11217,N_8117,N_8985);
nor U11218 (N_11218,N_8155,N_7494);
and U11219 (N_11219,N_8682,N_8703);
and U11220 (N_11220,N_6795,N_6122);
xor U11221 (N_11221,N_7865,N_6296);
or U11222 (N_11222,N_8071,N_8847);
nor U11223 (N_11223,N_8131,N_7640);
nand U11224 (N_11224,N_8527,N_6999);
xnor U11225 (N_11225,N_8556,N_7667);
or U11226 (N_11226,N_7388,N_7292);
xor U11227 (N_11227,N_6561,N_7168);
nand U11228 (N_11228,N_7521,N_8385);
nand U11229 (N_11229,N_6354,N_6481);
nand U11230 (N_11230,N_6082,N_8497);
nor U11231 (N_11231,N_6429,N_8059);
and U11232 (N_11232,N_8122,N_7499);
or U11233 (N_11233,N_8365,N_6760);
or U11234 (N_11234,N_6754,N_8554);
nor U11235 (N_11235,N_7923,N_6495);
nor U11236 (N_11236,N_7203,N_7189);
nor U11237 (N_11237,N_7819,N_7963);
nand U11238 (N_11238,N_6789,N_7346);
or U11239 (N_11239,N_6284,N_6868);
or U11240 (N_11240,N_7173,N_7386);
xor U11241 (N_11241,N_7751,N_6424);
nand U11242 (N_11242,N_6774,N_7923);
or U11243 (N_11243,N_8430,N_6778);
or U11244 (N_11244,N_7897,N_6078);
nand U11245 (N_11245,N_8933,N_7470);
xor U11246 (N_11246,N_6645,N_6144);
xor U11247 (N_11247,N_6661,N_6890);
or U11248 (N_11248,N_7333,N_8454);
nand U11249 (N_11249,N_8537,N_6016);
or U11250 (N_11250,N_6495,N_7928);
or U11251 (N_11251,N_7657,N_7550);
xnor U11252 (N_11252,N_6587,N_8272);
nor U11253 (N_11253,N_7591,N_6469);
and U11254 (N_11254,N_7971,N_7827);
and U11255 (N_11255,N_8316,N_8991);
or U11256 (N_11256,N_6464,N_6511);
and U11257 (N_11257,N_6461,N_6822);
nand U11258 (N_11258,N_7896,N_7172);
nor U11259 (N_11259,N_7411,N_7833);
nand U11260 (N_11260,N_7951,N_7858);
or U11261 (N_11261,N_7986,N_8530);
nor U11262 (N_11262,N_6735,N_6894);
xnor U11263 (N_11263,N_7908,N_7010);
nand U11264 (N_11264,N_6809,N_7132);
nand U11265 (N_11265,N_7859,N_6305);
nor U11266 (N_11266,N_8186,N_7769);
or U11267 (N_11267,N_8851,N_7505);
and U11268 (N_11268,N_6234,N_7455);
xnor U11269 (N_11269,N_6620,N_8694);
nor U11270 (N_11270,N_8662,N_8912);
or U11271 (N_11271,N_6997,N_6446);
and U11272 (N_11272,N_6894,N_8167);
nand U11273 (N_11273,N_8825,N_7508);
or U11274 (N_11274,N_8985,N_7483);
nor U11275 (N_11275,N_7628,N_7195);
nand U11276 (N_11276,N_7391,N_8702);
or U11277 (N_11277,N_7321,N_7890);
xor U11278 (N_11278,N_7407,N_7041);
or U11279 (N_11279,N_6855,N_7250);
nand U11280 (N_11280,N_7470,N_7226);
nor U11281 (N_11281,N_7377,N_8719);
or U11282 (N_11282,N_7167,N_6449);
and U11283 (N_11283,N_8348,N_7159);
nor U11284 (N_11284,N_8340,N_8569);
and U11285 (N_11285,N_7841,N_7557);
nand U11286 (N_11286,N_7735,N_6386);
xnor U11287 (N_11287,N_8810,N_6759);
and U11288 (N_11288,N_8459,N_8886);
xor U11289 (N_11289,N_6504,N_7977);
xnor U11290 (N_11290,N_8962,N_6860);
nand U11291 (N_11291,N_6717,N_7660);
nand U11292 (N_11292,N_7748,N_6206);
or U11293 (N_11293,N_7292,N_8378);
and U11294 (N_11294,N_7821,N_8102);
or U11295 (N_11295,N_6103,N_6552);
xnor U11296 (N_11296,N_8268,N_6217);
and U11297 (N_11297,N_6577,N_6947);
nand U11298 (N_11298,N_7626,N_8990);
nor U11299 (N_11299,N_8568,N_7714);
nand U11300 (N_11300,N_7223,N_6782);
xor U11301 (N_11301,N_6393,N_6786);
nor U11302 (N_11302,N_7285,N_8385);
nor U11303 (N_11303,N_7404,N_6899);
or U11304 (N_11304,N_6886,N_6679);
xnor U11305 (N_11305,N_7741,N_8718);
and U11306 (N_11306,N_7850,N_6814);
nand U11307 (N_11307,N_8280,N_7458);
or U11308 (N_11308,N_8529,N_8288);
or U11309 (N_11309,N_8098,N_8330);
nand U11310 (N_11310,N_8409,N_7372);
nor U11311 (N_11311,N_8468,N_6355);
and U11312 (N_11312,N_7081,N_6881);
nand U11313 (N_11313,N_6052,N_7048);
and U11314 (N_11314,N_8546,N_7573);
nand U11315 (N_11315,N_8098,N_8604);
xor U11316 (N_11316,N_8529,N_8677);
nand U11317 (N_11317,N_6664,N_8504);
xor U11318 (N_11318,N_8563,N_7193);
or U11319 (N_11319,N_8907,N_6251);
xor U11320 (N_11320,N_6777,N_6646);
nor U11321 (N_11321,N_7807,N_7334);
or U11322 (N_11322,N_7463,N_6370);
nand U11323 (N_11323,N_6647,N_8258);
or U11324 (N_11324,N_6346,N_7229);
xnor U11325 (N_11325,N_7034,N_8563);
xor U11326 (N_11326,N_6524,N_6755);
or U11327 (N_11327,N_7106,N_7136);
nand U11328 (N_11328,N_7588,N_8327);
nor U11329 (N_11329,N_6944,N_8494);
or U11330 (N_11330,N_8893,N_7348);
or U11331 (N_11331,N_7532,N_7665);
or U11332 (N_11332,N_6181,N_8680);
and U11333 (N_11333,N_7662,N_7207);
nor U11334 (N_11334,N_6156,N_7679);
and U11335 (N_11335,N_8538,N_6244);
nor U11336 (N_11336,N_8734,N_8102);
and U11337 (N_11337,N_7421,N_7350);
nor U11338 (N_11338,N_6394,N_6567);
and U11339 (N_11339,N_7129,N_8757);
nand U11340 (N_11340,N_7625,N_6004);
nand U11341 (N_11341,N_6687,N_6074);
xnor U11342 (N_11342,N_8727,N_7557);
xor U11343 (N_11343,N_7338,N_6537);
and U11344 (N_11344,N_8530,N_8369);
nand U11345 (N_11345,N_7746,N_7546);
and U11346 (N_11346,N_8138,N_8144);
and U11347 (N_11347,N_6240,N_8822);
or U11348 (N_11348,N_7216,N_6438);
or U11349 (N_11349,N_7298,N_6332);
xnor U11350 (N_11350,N_8969,N_8328);
nand U11351 (N_11351,N_8414,N_8900);
or U11352 (N_11352,N_7674,N_7256);
or U11353 (N_11353,N_7776,N_8282);
nand U11354 (N_11354,N_8197,N_8641);
nor U11355 (N_11355,N_6638,N_8786);
and U11356 (N_11356,N_6162,N_7818);
xor U11357 (N_11357,N_7720,N_6719);
xnor U11358 (N_11358,N_8744,N_6130);
xor U11359 (N_11359,N_6734,N_6764);
nand U11360 (N_11360,N_6781,N_6726);
and U11361 (N_11361,N_6075,N_7983);
and U11362 (N_11362,N_6075,N_6304);
nor U11363 (N_11363,N_6766,N_8579);
nor U11364 (N_11364,N_6318,N_6113);
or U11365 (N_11365,N_7481,N_6021);
and U11366 (N_11366,N_7314,N_8396);
or U11367 (N_11367,N_7348,N_6693);
or U11368 (N_11368,N_8141,N_7953);
and U11369 (N_11369,N_7355,N_7406);
or U11370 (N_11370,N_6813,N_8747);
nand U11371 (N_11371,N_8366,N_6668);
nand U11372 (N_11372,N_6407,N_6802);
and U11373 (N_11373,N_7497,N_6981);
and U11374 (N_11374,N_7443,N_7270);
or U11375 (N_11375,N_8491,N_8970);
nor U11376 (N_11376,N_6753,N_6764);
xor U11377 (N_11377,N_6451,N_7645);
or U11378 (N_11378,N_8589,N_8734);
and U11379 (N_11379,N_6862,N_7361);
nor U11380 (N_11380,N_8951,N_6255);
nor U11381 (N_11381,N_8297,N_7382);
xor U11382 (N_11382,N_6074,N_7177);
or U11383 (N_11383,N_6811,N_6665);
nand U11384 (N_11384,N_7038,N_8582);
and U11385 (N_11385,N_7736,N_8672);
nand U11386 (N_11386,N_8000,N_7905);
nor U11387 (N_11387,N_7709,N_6510);
and U11388 (N_11388,N_6926,N_7839);
nor U11389 (N_11389,N_8835,N_6277);
nand U11390 (N_11390,N_8473,N_8830);
nand U11391 (N_11391,N_8296,N_8925);
or U11392 (N_11392,N_7025,N_8635);
xnor U11393 (N_11393,N_8788,N_8420);
and U11394 (N_11394,N_6568,N_6923);
nand U11395 (N_11395,N_8623,N_8783);
nor U11396 (N_11396,N_7354,N_7022);
nor U11397 (N_11397,N_8555,N_7560);
nor U11398 (N_11398,N_6312,N_7279);
and U11399 (N_11399,N_8783,N_7489);
and U11400 (N_11400,N_7050,N_7838);
and U11401 (N_11401,N_8709,N_6219);
and U11402 (N_11402,N_8997,N_8240);
xor U11403 (N_11403,N_6153,N_6124);
xor U11404 (N_11404,N_6906,N_8272);
and U11405 (N_11405,N_7736,N_7055);
or U11406 (N_11406,N_8768,N_6788);
or U11407 (N_11407,N_8394,N_7622);
nand U11408 (N_11408,N_6866,N_8869);
or U11409 (N_11409,N_7883,N_7212);
or U11410 (N_11410,N_7036,N_6154);
nor U11411 (N_11411,N_7116,N_8019);
xor U11412 (N_11412,N_6919,N_8411);
nor U11413 (N_11413,N_8056,N_6456);
and U11414 (N_11414,N_8001,N_6294);
nor U11415 (N_11415,N_6244,N_7710);
nor U11416 (N_11416,N_8898,N_6231);
or U11417 (N_11417,N_7716,N_6619);
nand U11418 (N_11418,N_8786,N_7176);
and U11419 (N_11419,N_7723,N_8396);
xor U11420 (N_11420,N_7825,N_8052);
nor U11421 (N_11421,N_6845,N_7982);
nor U11422 (N_11422,N_6684,N_8625);
or U11423 (N_11423,N_8650,N_7690);
xnor U11424 (N_11424,N_8868,N_7467);
xnor U11425 (N_11425,N_6175,N_7586);
or U11426 (N_11426,N_7498,N_6800);
nand U11427 (N_11427,N_6145,N_7187);
and U11428 (N_11428,N_6797,N_6414);
and U11429 (N_11429,N_8059,N_8077);
xor U11430 (N_11430,N_8346,N_6460);
nand U11431 (N_11431,N_8744,N_8160);
nor U11432 (N_11432,N_8736,N_7927);
xnor U11433 (N_11433,N_8429,N_6176);
nor U11434 (N_11434,N_8643,N_6933);
nor U11435 (N_11435,N_8848,N_6277);
xor U11436 (N_11436,N_6694,N_8949);
or U11437 (N_11437,N_6404,N_7281);
and U11438 (N_11438,N_7580,N_6696);
nand U11439 (N_11439,N_6973,N_6428);
and U11440 (N_11440,N_8152,N_7723);
nand U11441 (N_11441,N_6944,N_8179);
and U11442 (N_11442,N_8995,N_8646);
nand U11443 (N_11443,N_7747,N_8511);
or U11444 (N_11444,N_8483,N_8297);
xor U11445 (N_11445,N_8302,N_6939);
nand U11446 (N_11446,N_7879,N_8282);
xnor U11447 (N_11447,N_8144,N_8146);
and U11448 (N_11448,N_8668,N_8217);
or U11449 (N_11449,N_7595,N_8312);
or U11450 (N_11450,N_6750,N_7008);
nand U11451 (N_11451,N_8922,N_6780);
and U11452 (N_11452,N_7661,N_8610);
xnor U11453 (N_11453,N_7798,N_7965);
and U11454 (N_11454,N_6558,N_6764);
nor U11455 (N_11455,N_8004,N_7527);
and U11456 (N_11456,N_6357,N_7228);
nor U11457 (N_11457,N_6836,N_6053);
nand U11458 (N_11458,N_6178,N_6749);
or U11459 (N_11459,N_8503,N_6967);
or U11460 (N_11460,N_7797,N_7027);
or U11461 (N_11461,N_6406,N_8712);
nand U11462 (N_11462,N_6389,N_8757);
nand U11463 (N_11463,N_8682,N_6473);
or U11464 (N_11464,N_6912,N_8057);
nand U11465 (N_11465,N_8424,N_8848);
or U11466 (N_11466,N_6622,N_6512);
nor U11467 (N_11467,N_6778,N_8098);
and U11468 (N_11468,N_6052,N_7810);
or U11469 (N_11469,N_8033,N_7160);
nor U11470 (N_11470,N_6142,N_6315);
or U11471 (N_11471,N_7903,N_8865);
and U11472 (N_11472,N_7125,N_7694);
and U11473 (N_11473,N_8863,N_6993);
and U11474 (N_11474,N_8548,N_6411);
nor U11475 (N_11475,N_7532,N_8083);
nand U11476 (N_11476,N_7407,N_8997);
or U11477 (N_11477,N_6909,N_7925);
nand U11478 (N_11478,N_8108,N_7352);
and U11479 (N_11479,N_8358,N_8236);
nor U11480 (N_11480,N_7668,N_8418);
and U11481 (N_11481,N_8495,N_8076);
xnor U11482 (N_11482,N_8321,N_6454);
xor U11483 (N_11483,N_6386,N_8122);
nand U11484 (N_11484,N_7225,N_6755);
or U11485 (N_11485,N_6467,N_6613);
xnor U11486 (N_11486,N_8304,N_6476);
or U11487 (N_11487,N_6273,N_8667);
or U11488 (N_11488,N_6892,N_6278);
and U11489 (N_11489,N_6341,N_6781);
nand U11490 (N_11490,N_7559,N_8798);
or U11491 (N_11491,N_8003,N_6657);
xnor U11492 (N_11492,N_6721,N_7902);
or U11493 (N_11493,N_8319,N_6296);
xnor U11494 (N_11494,N_6219,N_7289);
and U11495 (N_11495,N_7067,N_8281);
or U11496 (N_11496,N_8853,N_6529);
xnor U11497 (N_11497,N_8348,N_7480);
nand U11498 (N_11498,N_6677,N_8448);
xor U11499 (N_11499,N_8190,N_6613);
nor U11500 (N_11500,N_6382,N_6500);
and U11501 (N_11501,N_8646,N_8247);
xnor U11502 (N_11502,N_7884,N_6110);
nor U11503 (N_11503,N_6724,N_7201);
nand U11504 (N_11504,N_6327,N_6371);
or U11505 (N_11505,N_7368,N_6214);
or U11506 (N_11506,N_6926,N_7841);
and U11507 (N_11507,N_7947,N_6349);
xnor U11508 (N_11508,N_8449,N_7726);
nor U11509 (N_11509,N_6381,N_7406);
nand U11510 (N_11510,N_6902,N_8029);
and U11511 (N_11511,N_7372,N_7291);
nor U11512 (N_11512,N_7903,N_8385);
nand U11513 (N_11513,N_6340,N_8764);
nor U11514 (N_11514,N_8166,N_6980);
nor U11515 (N_11515,N_7611,N_7743);
xor U11516 (N_11516,N_8903,N_7981);
or U11517 (N_11517,N_8913,N_8099);
or U11518 (N_11518,N_7151,N_6546);
or U11519 (N_11519,N_8499,N_7404);
and U11520 (N_11520,N_6642,N_8110);
xor U11521 (N_11521,N_6011,N_6588);
xor U11522 (N_11522,N_6941,N_7840);
nor U11523 (N_11523,N_7952,N_7040);
and U11524 (N_11524,N_8501,N_8750);
nand U11525 (N_11525,N_6598,N_7865);
or U11526 (N_11526,N_8861,N_6133);
xor U11527 (N_11527,N_6336,N_6517);
and U11528 (N_11528,N_7499,N_8735);
and U11529 (N_11529,N_8534,N_7584);
xnor U11530 (N_11530,N_7497,N_7429);
and U11531 (N_11531,N_8334,N_8593);
nor U11532 (N_11532,N_7247,N_8331);
xor U11533 (N_11533,N_6930,N_8440);
nand U11534 (N_11534,N_6090,N_8823);
xor U11535 (N_11535,N_8177,N_6116);
or U11536 (N_11536,N_8495,N_8856);
nor U11537 (N_11537,N_7450,N_7493);
or U11538 (N_11538,N_6903,N_7733);
nand U11539 (N_11539,N_6945,N_7256);
nand U11540 (N_11540,N_8671,N_7136);
nand U11541 (N_11541,N_7431,N_8537);
xor U11542 (N_11542,N_6391,N_7086);
xor U11543 (N_11543,N_8653,N_8577);
nand U11544 (N_11544,N_7115,N_8348);
and U11545 (N_11545,N_6136,N_8351);
and U11546 (N_11546,N_6998,N_7761);
nand U11547 (N_11547,N_6223,N_7562);
or U11548 (N_11548,N_6409,N_8877);
nor U11549 (N_11549,N_8543,N_6791);
nor U11550 (N_11550,N_6447,N_8602);
or U11551 (N_11551,N_7552,N_8726);
nand U11552 (N_11552,N_6148,N_8301);
xnor U11553 (N_11553,N_7644,N_7186);
and U11554 (N_11554,N_8105,N_8972);
nor U11555 (N_11555,N_6054,N_6741);
or U11556 (N_11556,N_6075,N_6662);
xnor U11557 (N_11557,N_8600,N_6807);
xor U11558 (N_11558,N_7078,N_7333);
and U11559 (N_11559,N_8705,N_7688);
and U11560 (N_11560,N_8778,N_8430);
nor U11561 (N_11561,N_7025,N_7467);
or U11562 (N_11562,N_6309,N_7503);
xnor U11563 (N_11563,N_8134,N_7335);
nand U11564 (N_11564,N_8103,N_8751);
and U11565 (N_11565,N_7535,N_7107);
nand U11566 (N_11566,N_6176,N_7602);
xnor U11567 (N_11567,N_8867,N_6401);
nand U11568 (N_11568,N_6633,N_6912);
or U11569 (N_11569,N_8908,N_8634);
xnor U11570 (N_11570,N_8267,N_7026);
nand U11571 (N_11571,N_8295,N_8140);
xor U11572 (N_11572,N_7615,N_6237);
nor U11573 (N_11573,N_7797,N_6423);
and U11574 (N_11574,N_6107,N_7694);
nand U11575 (N_11575,N_8438,N_8996);
nor U11576 (N_11576,N_8342,N_8335);
or U11577 (N_11577,N_7309,N_7469);
nand U11578 (N_11578,N_6796,N_7001);
or U11579 (N_11579,N_7493,N_7854);
or U11580 (N_11580,N_8001,N_8338);
xor U11581 (N_11581,N_8051,N_6844);
and U11582 (N_11582,N_7474,N_6619);
or U11583 (N_11583,N_7953,N_8756);
nand U11584 (N_11584,N_7148,N_7327);
and U11585 (N_11585,N_7932,N_6676);
or U11586 (N_11586,N_7323,N_8678);
nor U11587 (N_11587,N_6258,N_7669);
nand U11588 (N_11588,N_8499,N_8460);
or U11589 (N_11589,N_7979,N_7559);
and U11590 (N_11590,N_8536,N_8722);
nand U11591 (N_11591,N_6140,N_7861);
or U11592 (N_11592,N_7003,N_6060);
and U11593 (N_11593,N_8619,N_6223);
nand U11594 (N_11594,N_7585,N_7496);
or U11595 (N_11595,N_8243,N_6895);
and U11596 (N_11596,N_7306,N_6467);
xnor U11597 (N_11597,N_8673,N_7254);
nand U11598 (N_11598,N_6164,N_8589);
nand U11599 (N_11599,N_6744,N_6577);
or U11600 (N_11600,N_7215,N_8114);
and U11601 (N_11601,N_6565,N_6945);
xor U11602 (N_11602,N_6114,N_7306);
or U11603 (N_11603,N_8847,N_7745);
or U11604 (N_11604,N_8038,N_6343);
xor U11605 (N_11605,N_8974,N_6291);
and U11606 (N_11606,N_6915,N_8344);
nand U11607 (N_11607,N_6905,N_7750);
and U11608 (N_11608,N_7052,N_6051);
and U11609 (N_11609,N_8862,N_6436);
xor U11610 (N_11610,N_6259,N_8534);
xnor U11611 (N_11611,N_8577,N_7832);
or U11612 (N_11612,N_8759,N_6411);
xor U11613 (N_11613,N_8242,N_8996);
or U11614 (N_11614,N_8850,N_7027);
and U11615 (N_11615,N_8925,N_7601);
and U11616 (N_11616,N_7320,N_6991);
and U11617 (N_11617,N_7653,N_7732);
nor U11618 (N_11618,N_6887,N_8126);
nand U11619 (N_11619,N_8917,N_6653);
or U11620 (N_11620,N_7668,N_8428);
and U11621 (N_11621,N_6041,N_6749);
or U11622 (N_11622,N_6170,N_8991);
xor U11623 (N_11623,N_7608,N_6554);
nand U11624 (N_11624,N_6200,N_7540);
nand U11625 (N_11625,N_6271,N_6708);
and U11626 (N_11626,N_7231,N_7064);
or U11627 (N_11627,N_8523,N_7573);
and U11628 (N_11628,N_6791,N_8052);
and U11629 (N_11629,N_6880,N_7255);
or U11630 (N_11630,N_7030,N_8944);
xor U11631 (N_11631,N_8400,N_6618);
nand U11632 (N_11632,N_7713,N_6586);
xor U11633 (N_11633,N_7802,N_8537);
xnor U11634 (N_11634,N_7198,N_7831);
nor U11635 (N_11635,N_6895,N_7353);
xor U11636 (N_11636,N_7310,N_8738);
and U11637 (N_11637,N_6852,N_7606);
nand U11638 (N_11638,N_7608,N_7140);
nand U11639 (N_11639,N_7684,N_8824);
nand U11640 (N_11640,N_8543,N_6672);
xnor U11641 (N_11641,N_6672,N_6908);
xor U11642 (N_11642,N_7086,N_8600);
and U11643 (N_11643,N_8667,N_7197);
xor U11644 (N_11644,N_6908,N_6697);
nand U11645 (N_11645,N_8748,N_7699);
and U11646 (N_11646,N_6097,N_8245);
nor U11647 (N_11647,N_8257,N_6902);
nor U11648 (N_11648,N_7893,N_7120);
nor U11649 (N_11649,N_8611,N_7023);
or U11650 (N_11650,N_8388,N_7145);
nor U11651 (N_11651,N_7166,N_8630);
or U11652 (N_11652,N_6301,N_6280);
or U11653 (N_11653,N_8658,N_6243);
nand U11654 (N_11654,N_7856,N_7535);
nand U11655 (N_11655,N_8703,N_7487);
or U11656 (N_11656,N_8532,N_8240);
and U11657 (N_11657,N_8484,N_7196);
nor U11658 (N_11658,N_6539,N_7855);
nand U11659 (N_11659,N_6922,N_8249);
and U11660 (N_11660,N_6772,N_6593);
nor U11661 (N_11661,N_8404,N_6786);
xnor U11662 (N_11662,N_7626,N_7949);
xor U11663 (N_11663,N_6777,N_8276);
or U11664 (N_11664,N_8026,N_8863);
nand U11665 (N_11665,N_7797,N_8684);
or U11666 (N_11666,N_6859,N_6956);
and U11667 (N_11667,N_6740,N_8734);
xor U11668 (N_11668,N_6788,N_7220);
xnor U11669 (N_11669,N_6793,N_7761);
and U11670 (N_11670,N_8137,N_6814);
and U11671 (N_11671,N_8509,N_6968);
and U11672 (N_11672,N_6052,N_6027);
or U11673 (N_11673,N_7546,N_8672);
and U11674 (N_11674,N_7322,N_8830);
xnor U11675 (N_11675,N_7893,N_8096);
xnor U11676 (N_11676,N_7421,N_7470);
and U11677 (N_11677,N_8623,N_7625);
or U11678 (N_11678,N_6017,N_8169);
nand U11679 (N_11679,N_8195,N_6120);
nor U11680 (N_11680,N_8846,N_8373);
nor U11681 (N_11681,N_8705,N_6211);
xor U11682 (N_11682,N_8601,N_6550);
or U11683 (N_11683,N_6021,N_6583);
nor U11684 (N_11684,N_8455,N_8679);
xor U11685 (N_11685,N_7290,N_6579);
and U11686 (N_11686,N_6564,N_6346);
nor U11687 (N_11687,N_8336,N_7351);
nand U11688 (N_11688,N_7594,N_8325);
and U11689 (N_11689,N_8309,N_6064);
or U11690 (N_11690,N_6580,N_8373);
xnor U11691 (N_11691,N_7684,N_6458);
xnor U11692 (N_11692,N_8321,N_8166);
nand U11693 (N_11693,N_7373,N_7783);
nand U11694 (N_11694,N_7438,N_8456);
xnor U11695 (N_11695,N_7231,N_7537);
nand U11696 (N_11696,N_6027,N_8027);
nor U11697 (N_11697,N_7674,N_6476);
and U11698 (N_11698,N_6079,N_8188);
or U11699 (N_11699,N_7529,N_7333);
nand U11700 (N_11700,N_7593,N_6347);
nand U11701 (N_11701,N_6994,N_7872);
nor U11702 (N_11702,N_7819,N_6470);
and U11703 (N_11703,N_8413,N_8658);
or U11704 (N_11704,N_6503,N_6688);
or U11705 (N_11705,N_7148,N_7392);
xnor U11706 (N_11706,N_6423,N_6614);
nor U11707 (N_11707,N_6107,N_8068);
nor U11708 (N_11708,N_6250,N_7801);
and U11709 (N_11709,N_8228,N_6100);
and U11710 (N_11710,N_8948,N_6206);
xnor U11711 (N_11711,N_7842,N_7289);
xor U11712 (N_11712,N_8496,N_8767);
nor U11713 (N_11713,N_7734,N_8149);
nor U11714 (N_11714,N_6116,N_8407);
nand U11715 (N_11715,N_7036,N_6905);
or U11716 (N_11716,N_7328,N_6463);
or U11717 (N_11717,N_8902,N_6035);
or U11718 (N_11718,N_6312,N_8371);
and U11719 (N_11719,N_6076,N_6292);
or U11720 (N_11720,N_6161,N_7760);
xor U11721 (N_11721,N_8288,N_8537);
xor U11722 (N_11722,N_6293,N_6944);
and U11723 (N_11723,N_8511,N_7116);
nand U11724 (N_11724,N_7899,N_7764);
or U11725 (N_11725,N_7568,N_6080);
or U11726 (N_11726,N_7860,N_7529);
nor U11727 (N_11727,N_7544,N_6576);
nor U11728 (N_11728,N_6846,N_8642);
nor U11729 (N_11729,N_6009,N_6984);
and U11730 (N_11730,N_7060,N_6543);
xor U11731 (N_11731,N_8048,N_7079);
xnor U11732 (N_11732,N_8067,N_8583);
and U11733 (N_11733,N_8182,N_7070);
xnor U11734 (N_11734,N_7372,N_8837);
xor U11735 (N_11735,N_6044,N_7959);
and U11736 (N_11736,N_6666,N_6843);
xor U11737 (N_11737,N_8647,N_6101);
and U11738 (N_11738,N_8015,N_7705);
nand U11739 (N_11739,N_8638,N_8560);
and U11740 (N_11740,N_7599,N_8930);
nand U11741 (N_11741,N_6373,N_7572);
nor U11742 (N_11742,N_6133,N_6268);
or U11743 (N_11743,N_8397,N_6096);
nor U11744 (N_11744,N_6209,N_7138);
nor U11745 (N_11745,N_7285,N_8579);
or U11746 (N_11746,N_7417,N_8966);
and U11747 (N_11747,N_6743,N_6274);
or U11748 (N_11748,N_7089,N_7133);
nand U11749 (N_11749,N_6821,N_7613);
or U11750 (N_11750,N_6520,N_8421);
or U11751 (N_11751,N_6086,N_7626);
nor U11752 (N_11752,N_8122,N_8278);
nor U11753 (N_11753,N_7467,N_7005);
nand U11754 (N_11754,N_6057,N_8907);
xnor U11755 (N_11755,N_6029,N_6126);
xor U11756 (N_11756,N_7253,N_7465);
or U11757 (N_11757,N_6635,N_6315);
and U11758 (N_11758,N_6491,N_7289);
nand U11759 (N_11759,N_7824,N_7518);
or U11760 (N_11760,N_8699,N_6933);
or U11761 (N_11761,N_8315,N_7629);
and U11762 (N_11762,N_7089,N_8251);
and U11763 (N_11763,N_6319,N_6054);
nand U11764 (N_11764,N_8017,N_7488);
xor U11765 (N_11765,N_8764,N_7152);
or U11766 (N_11766,N_8216,N_8502);
nand U11767 (N_11767,N_8406,N_8338);
nor U11768 (N_11768,N_6518,N_7800);
or U11769 (N_11769,N_8623,N_6219);
or U11770 (N_11770,N_6744,N_6362);
xnor U11771 (N_11771,N_7175,N_7996);
xor U11772 (N_11772,N_6915,N_6881);
nor U11773 (N_11773,N_6229,N_8911);
nand U11774 (N_11774,N_8845,N_7987);
and U11775 (N_11775,N_8075,N_7110);
nand U11776 (N_11776,N_7261,N_8528);
and U11777 (N_11777,N_8338,N_6909);
and U11778 (N_11778,N_8224,N_8843);
or U11779 (N_11779,N_6109,N_7228);
or U11780 (N_11780,N_8085,N_8145);
and U11781 (N_11781,N_6724,N_7784);
or U11782 (N_11782,N_6739,N_7046);
or U11783 (N_11783,N_6963,N_6049);
and U11784 (N_11784,N_6346,N_6960);
or U11785 (N_11785,N_8931,N_7602);
nand U11786 (N_11786,N_6961,N_8105);
and U11787 (N_11787,N_8807,N_7114);
and U11788 (N_11788,N_7083,N_7683);
nand U11789 (N_11789,N_6922,N_6792);
and U11790 (N_11790,N_7862,N_6461);
nand U11791 (N_11791,N_6860,N_8847);
and U11792 (N_11792,N_7327,N_7942);
and U11793 (N_11793,N_6686,N_7773);
xnor U11794 (N_11794,N_6861,N_6580);
and U11795 (N_11795,N_6548,N_6364);
xnor U11796 (N_11796,N_8337,N_7693);
or U11797 (N_11797,N_7918,N_8230);
and U11798 (N_11798,N_6286,N_6106);
or U11799 (N_11799,N_7777,N_8649);
and U11800 (N_11800,N_6562,N_8217);
nand U11801 (N_11801,N_7465,N_6152);
nor U11802 (N_11802,N_7580,N_8202);
and U11803 (N_11803,N_6899,N_7861);
nand U11804 (N_11804,N_6087,N_7416);
xnor U11805 (N_11805,N_7789,N_7869);
or U11806 (N_11806,N_7253,N_6617);
nor U11807 (N_11807,N_6387,N_6458);
nand U11808 (N_11808,N_8508,N_6466);
and U11809 (N_11809,N_6502,N_7896);
nand U11810 (N_11810,N_7974,N_7040);
xnor U11811 (N_11811,N_6477,N_8933);
and U11812 (N_11812,N_8888,N_8018);
and U11813 (N_11813,N_7325,N_7882);
nand U11814 (N_11814,N_8544,N_8235);
nand U11815 (N_11815,N_6974,N_8587);
xnor U11816 (N_11816,N_7421,N_6928);
xnor U11817 (N_11817,N_8803,N_6291);
nand U11818 (N_11818,N_6880,N_6857);
or U11819 (N_11819,N_6825,N_8900);
and U11820 (N_11820,N_6775,N_6862);
or U11821 (N_11821,N_8555,N_7043);
nand U11822 (N_11822,N_8373,N_7154);
or U11823 (N_11823,N_8070,N_7614);
nor U11824 (N_11824,N_6324,N_6327);
nand U11825 (N_11825,N_7196,N_7304);
nand U11826 (N_11826,N_6961,N_6121);
xnor U11827 (N_11827,N_8611,N_7471);
nor U11828 (N_11828,N_8507,N_6724);
nand U11829 (N_11829,N_6184,N_7521);
or U11830 (N_11830,N_7074,N_6386);
nor U11831 (N_11831,N_7584,N_7121);
and U11832 (N_11832,N_6456,N_7358);
and U11833 (N_11833,N_7344,N_6796);
or U11834 (N_11834,N_7501,N_8331);
or U11835 (N_11835,N_6623,N_7475);
and U11836 (N_11836,N_6614,N_6161);
xnor U11837 (N_11837,N_6207,N_8874);
and U11838 (N_11838,N_7227,N_7138);
and U11839 (N_11839,N_8507,N_8344);
and U11840 (N_11840,N_6067,N_8368);
xnor U11841 (N_11841,N_8349,N_7273);
and U11842 (N_11842,N_7200,N_6373);
or U11843 (N_11843,N_7645,N_8937);
nand U11844 (N_11844,N_6408,N_6370);
or U11845 (N_11845,N_6843,N_6908);
xor U11846 (N_11846,N_7928,N_8723);
nand U11847 (N_11847,N_7936,N_6100);
nand U11848 (N_11848,N_8723,N_6427);
xnor U11849 (N_11849,N_7522,N_8852);
nor U11850 (N_11850,N_7019,N_8405);
xnor U11851 (N_11851,N_8620,N_6309);
nand U11852 (N_11852,N_7968,N_6921);
and U11853 (N_11853,N_6836,N_7141);
nor U11854 (N_11854,N_6714,N_8995);
nor U11855 (N_11855,N_7907,N_6090);
nand U11856 (N_11856,N_8533,N_6302);
and U11857 (N_11857,N_6010,N_7838);
or U11858 (N_11858,N_6259,N_8478);
xnor U11859 (N_11859,N_7029,N_8386);
nor U11860 (N_11860,N_7592,N_8847);
xor U11861 (N_11861,N_8790,N_8304);
nor U11862 (N_11862,N_6178,N_6485);
or U11863 (N_11863,N_7896,N_8707);
nor U11864 (N_11864,N_6262,N_8218);
xnor U11865 (N_11865,N_8221,N_6634);
and U11866 (N_11866,N_7478,N_8752);
xor U11867 (N_11867,N_7817,N_8299);
nand U11868 (N_11868,N_6959,N_7487);
nand U11869 (N_11869,N_8281,N_8269);
and U11870 (N_11870,N_8347,N_7256);
and U11871 (N_11871,N_7280,N_6079);
nand U11872 (N_11872,N_7791,N_8405);
or U11873 (N_11873,N_6149,N_8298);
xnor U11874 (N_11874,N_7312,N_6757);
nand U11875 (N_11875,N_7803,N_7879);
or U11876 (N_11876,N_8986,N_7428);
nor U11877 (N_11877,N_7111,N_6458);
xnor U11878 (N_11878,N_7609,N_7507);
or U11879 (N_11879,N_7052,N_8217);
xor U11880 (N_11880,N_7832,N_6563);
or U11881 (N_11881,N_6414,N_8228);
xnor U11882 (N_11882,N_8336,N_8174);
nor U11883 (N_11883,N_8464,N_6264);
xor U11884 (N_11884,N_7317,N_6117);
or U11885 (N_11885,N_7835,N_6570);
nor U11886 (N_11886,N_7614,N_7659);
nand U11887 (N_11887,N_7566,N_6848);
nor U11888 (N_11888,N_6836,N_8075);
nor U11889 (N_11889,N_6242,N_7827);
nor U11890 (N_11890,N_7198,N_7590);
nand U11891 (N_11891,N_6676,N_7372);
nor U11892 (N_11892,N_8668,N_6821);
xor U11893 (N_11893,N_7253,N_8519);
xor U11894 (N_11894,N_6672,N_6644);
and U11895 (N_11895,N_7685,N_7266);
and U11896 (N_11896,N_8384,N_6764);
nand U11897 (N_11897,N_6499,N_6464);
or U11898 (N_11898,N_7545,N_8128);
nor U11899 (N_11899,N_8436,N_7358);
nor U11900 (N_11900,N_7953,N_7529);
xnor U11901 (N_11901,N_7321,N_7223);
or U11902 (N_11902,N_6072,N_6352);
and U11903 (N_11903,N_8498,N_7691);
nor U11904 (N_11904,N_7176,N_6184);
nand U11905 (N_11905,N_6461,N_6299);
xor U11906 (N_11906,N_7743,N_7579);
and U11907 (N_11907,N_7940,N_8667);
nor U11908 (N_11908,N_8319,N_7016);
nor U11909 (N_11909,N_6055,N_6247);
nand U11910 (N_11910,N_7274,N_8010);
and U11911 (N_11911,N_7128,N_8435);
xor U11912 (N_11912,N_7639,N_8587);
xor U11913 (N_11913,N_7017,N_6299);
xor U11914 (N_11914,N_7274,N_7978);
xnor U11915 (N_11915,N_6777,N_6141);
nand U11916 (N_11916,N_6202,N_6693);
nor U11917 (N_11917,N_8464,N_8161);
and U11918 (N_11918,N_7728,N_8686);
nand U11919 (N_11919,N_8888,N_7476);
xor U11920 (N_11920,N_7516,N_7312);
xor U11921 (N_11921,N_8258,N_6426);
nor U11922 (N_11922,N_7550,N_7835);
and U11923 (N_11923,N_6968,N_7214);
and U11924 (N_11924,N_7442,N_6331);
or U11925 (N_11925,N_8326,N_7543);
nand U11926 (N_11926,N_6862,N_8321);
xor U11927 (N_11927,N_8685,N_8163);
or U11928 (N_11928,N_6015,N_8118);
nor U11929 (N_11929,N_6512,N_7995);
nor U11930 (N_11930,N_6734,N_7824);
nor U11931 (N_11931,N_8852,N_7453);
or U11932 (N_11932,N_8636,N_8616);
nor U11933 (N_11933,N_8874,N_7421);
nand U11934 (N_11934,N_6071,N_8121);
nand U11935 (N_11935,N_8359,N_8975);
nand U11936 (N_11936,N_8257,N_8433);
xnor U11937 (N_11937,N_7104,N_8781);
or U11938 (N_11938,N_8089,N_7546);
nand U11939 (N_11939,N_7312,N_6264);
nor U11940 (N_11940,N_7868,N_8468);
nor U11941 (N_11941,N_8214,N_6274);
nor U11942 (N_11942,N_6139,N_6841);
or U11943 (N_11943,N_6929,N_8593);
xnor U11944 (N_11944,N_8789,N_7584);
nand U11945 (N_11945,N_6009,N_8196);
or U11946 (N_11946,N_6042,N_8807);
nand U11947 (N_11947,N_6180,N_8100);
xor U11948 (N_11948,N_8468,N_6718);
xor U11949 (N_11949,N_7378,N_6273);
and U11950 (N_11950,N_6247,N_8743);
or U11951 (N_11951,N_8921,N_6807);
or U11952 (N_11952,N_7414,N_7608);
xor U11953 (N_11953,N_6056,N_7288);
nor U11954 (N_11954,N_6375,N_6857);
xnor U11955 (N_11955,N_8462,N_7461);
nor U11956 (N_11956,N_8739,N_8241);
and U11957 (N_11957,N_6464,N_8719);
nand U11958 (N_11958,N_6526,N_7934);
nor U11959 (N_11959,N_6345,N_6971);
nor U11960 (N_11960,N_6476,N_6928);
nor U11961 (N_11961,N_8166,N_6839);
and U11962 (N_11962,N_8342,N_6572);
or U11963 (N_11963,N_7568,N_8888);
or U11964 (N_11964,N_8196,N_8283);
nand U11965 (N_11965,N_8050,N_6260);
and U11966 (N_11966,N_8171,N_8521);
nand U11967 (N_11967,N_8383,N_8478);
xor U11968 (N_11968,N_7255,N_6416);
xnor U11969 (N_11969,N_6863,N_6566);
and U11970 (N_11970,N_7826,N_8339);
or U11971 (N_11971,N_7428,N_7316);
or U11972 (N_11972,N_8702,N_6073);
xor U11973 (N_11973,N_8952,N_8172);
and U11974 (N_11974,N_6433,N_6621);
or U11975 (N_11975,N_8673,N_6667);
xnor U11976 (N_11976,N_7563,N_7464);
xnor U11977 (N_11977,N_8193,N_6888);
and U11978 (N_11978,N_6530,N_8023);
and U11979 (N_11979,N_7236,N_8166);
xnor U11980 (N_11980,N_8920,N_6749);
and U11981 (N_11981,N_6668,N_8671);
and U11982 (N_11982,N_8962,N_6516);
xnor U11983 (N_11983,N_6224,N_8680);
nor U11984 (N_11984,N_6043,N_7513);
nor U11985 (N_11985,N_6100,N_7269);
nor U11986 (N_11986,N_8945,N_8505);
and U11987 (N_11987,N_6988,N_7463);
nor U11988 (N_11988,N_8681,N_6628);
xor U11989 (N_11989,N_8364,N_8158);
and U11990 (N_11990,N_6190,N_8052);
nor U11991 (N_11991,N_7241,N_8014);
and U11992 (N_11992,N_8158,N_8684);
xor U11993 (N_11993,N_7508,N_6980);
nand U11994 (N_11994,N_6666,N_7870);
xor U11995 (N_11995,N_6659,N_8092);
and U11996 (N_11996,N_6277,N_6185);
or U11997 (N_11997,N_7503,N_8264);
xnor U11998 (N_11998,N_8938,N_7381);
nand U11999 (N_11999,N_8391,N_8729);
nor U12000 (N_12000,N_11821,N_10184);
nor U12001 (N_12001,N_9202,N_9070);
nand U12002 (N_12002,N_9660,N_9947);
nor U12003 (N_12003,N_10107,N_9817);
xnor U12004 (N_12004,N_11029,N_9609);
nand U12005 (N_12005,N_10938,N_10222);
nand U12006 (N_12006,N_9510,N_11687);
xor U12007 (N_12007,N_10385,N_11890);
or U12008 (N_12008,N_9822,N_11280);
xnor U12009 (N_12009,N_11377,N_10426);
nor U12010 (N_12010,N_10813,N_11191);
nor U12011 (N_12011,N_10809,N_9071);
nand U12012 (N_12012,N_11321,N_9433);
xor U12013 (N_12013,N_9512,N_11876);
or U12014 (N_12014,N_10988,N_11941);
and U12015 (N_12015,N_9271,N_9062);
nand U12016 (N_12016,N_10878,N_11420);
and U12017 (N_12017,N_10700,N_10658);
nor U12018 (N_12018,N_11038,N_11700);
nor U12019 (N_12019,N_10195,N_9326);
nor U12020 (N_12020,N_11788,N_9905);
and U12021 (N_12021,N_10260,N_11131);
and U12022 (N_12022,N_10987,N_11880);
xnor U12023 (N_12023,N_10905,N_10677);
and U12024 (N_12024,N_11744,N_9385);
xor U12025 (N_12025,N_11680,N_11510);
or U12026 (N_12026,N_11389,N_9221);
and U12027 (N_12027,N_11780,N_10354);
nand U12028 (N_12028,N_10851,N_10580);
xor U12029 (N_12029,N_11889,N_9025);
nand U12030 (N_12030,N_9603,N_11411);
xnor U12031 (N_12031,N_10553,N_11555);
or U12032 (N_12032,N_9834,N_10453);
or U12033 (N_12033,N_9358,N_10512);
nand U12034 (N_12034,N_9377,N_9236);
and U12035 (N_12035,N_11842,N_11532);
xnor U12036 (N_12036,N_11487,N_9327);
nor U12037 (N_12037,N_11175,N_10948);
xor U12038 (N_12038,N_11625,N_9198);
and U12039 (N_12039,N_9415,N_10214);
nor U12040 (N_12040,N_9901,N_9696);
nand U12041 (N_12041,N_10775,N_10893);
or U12042 (N_12042,N_10925,N_9796);
nor U12043 (N_12043,N_11079,N_9953);
or U12044 (N_12044,N_9347,N_9143);
and U12045 (N_12045,N_9223,N_10614);
or U12046 (N_12046,N_10589,N_10029);
nand U12047 (N_12047,N_9148,N_11927);
nand U12048 (N_12048,N_10316,N_9455);
or U12049 (N_12049,N_9361,N_10140);
or U12050 (N_12050,N_10063,N_10175);
nor U12051 (N_12051,N_10120,N_9706);
or U12052 (N_12052,N_9006,N_9515);
xor U12053 (N_12053,N_10365,N_9673);
and U12054 (N_12054,N_10173,N_9081);
xor U12055 (N_12055,N_10145,N_11645);
nand U12056 (N_12056,N_10711,N_11947);
and U12057 (N_12057,N_10479,N_10537);
xnor U12058 (N_12058,N_9781,N_10539);
or U12059 (N_12059,N_9368,N_10875);
nand U12060 (N_12060,N_10480,N_11849);
nor U12061 (N_12061,N_10502,N_10445);
nor U12062 (N_12062,N_11317,N_11310);
or U12063 (N_12063,N_9352,N_10774);
or U12064 (N_12064,N_9357,N_11629);
xor U12065 (N_12065,N_9543,N_11763);
xnor U12066 (N_12066,N_9176,N_11792);
nor U12067 (N_12067,N_9885,N_11058);
and U12068 (N_12068,N_10165,N_11743);
nand U12069 (N_12069,N_9839,N_10628);
nor U12070 (N_12070,N_10257,N_9304);
or U12071 (N_12071,N_10959,N_9344);
xnor U12072 (N_12072,N_11450,N_11202);
and U12073 (N_12073,N_11998,N_9168);
nand U12074 (N_12074,N_11875,N_11279);
xnor U12075 (N_12075,N_9917,N_11395);
nor U12076 (N_12076,N_10467,N_11041);
nor U12077 (N_12077,N_10205,N_10287);
nor U12078 (N_12078,N_10202,N_10003);
xor U12079 (N_12079,N_11285,N_11168);
or U12080 (N_12080,N_10962,N_11047);
nor U12081 (N_12081,N_10956,N_9041);
nor U12082 (N_12082,N_10398,N_11503);
nor U12083 (N_12083,N_9591,N_10719);
nand U12084 (N_12084,N_11009,N_10507);
nor U12085 (N_12085,N_11406,N_11888);
or U12086 (N_12086,N_10309,N_11708);
nand U12087 (N_12087,N_9920,N_9235);
nor U12088 (N_12088,N_11707,N_11380);
nand U12089 (N_12089,N_10736,N_10336);
nor U12090 (N_12090,N_11392,N_10889);
xnor U12091 (N_12091,N_10321,N_11588);
or U12092 (N_12092,N_9274,N_9454);
xnor U12093 (N_12093,N_11526,N_10627);
nor U12094 (N_12094,N_9027,N_10413);
and U12095 (N_12095,N_10028,N_11422);
nand U12096 (N_12096,N_10425,N_11290);
or U12097 (N_12097,N_11263,N_11211);
or U12098 (N_12098,N_11542,N_11097);
nor U12099 (N_12099,N_11940,N_9026);
and U12100 (N_12100,N_10647,N_11346);
nor U12101 (N_12101,N_10492,N_9945);
nor U12102 (N_12102,N_10604,N_11701);
or U12103 (N_12103,N_9316,N_11479);
nor U12104 (N_12104,N_11227,N_10348);
xnor U12105 (N_12105,N_11098,N_9872);
or U12106 (N_12106,N_9576,N_10164);
or U12107 (N_12107,N_11602,N_9575);
or U12108 (N_12108,N_10052,N_9107);
xor U12109 (N_12109,N_10139,N_10543);
nand U12110 (N_12110,N_10887,N_10803);
and U12111 (N_12111,N_10111,N_10181);
xnor U12112 (N_12112,N_10346,N_9932);
nor U12113 (N_12113,N_9560,N_11839);
and U12114 (N_12114,N_11515,N_11275);
and U12115 (N_12115,N_10076,N_9426);
and U12116 (N_12116,N_9808,N_10223);
nor U12117 (N_12117,N_11458,N_11731);
and U12118 (N_12118,N_11613,N_11749);
nand U12119 (N_12119,N_11149,N_10639);
and U12120 (N_12120,N_11809,N_9362);
xor U12121 (N_12121,N_11141,N_11240);
nor U12122 (N_12122,N_9323,N_11699);
nor U12123 (N_12123,N_11081,N_9783);
nand U12124 (N_12124,N_9338,N_10772);
nand U12125 (N_12125,N_10523,N_11461);
or U12126 (N_12126,N_11137,N_10459);
nand U12127 (N_12127,N_11664,N_9131);
xor U12128 (N_12128,N_10421,N_9488);
or U12129 (N_12129,N_9770,N_11987);
nand U12130 (N_12130,N_10780,N_10300);
and U12131 (N_12131,N_11774,N_11896);
nand U12132 (N_12132,N_11087,N_10645);
nand U12133 (N_12133,N_11902,N_9369);
nor U12134 (N_12134,N_10022,N_9302);
nor U12135 (N_12135,N_9757,N_9868);
and U12136 (N_12136,N_11414,N_9043);
nor U12137 (N_12137,N_11383,N_9178);
or U12138 (N_12138,N_9170,N_9634);
xor U12139 (N_12139,N_11019,N_10849);
nor U12140 (N_12140,N_9711,N_10100);
or U12141 (N_12141,N_11897,N_10970);
nand U12142 (N_12142,N_10162,N_9388);
xor U12143 (N_12143,N_9830,N_10037);
nand U12144 (N_12144,N_10693,N_11378);
or U12145 (N_12145,N_11758,N_11078);
and U12146 (N_12146,N_10109,N_9756);
nor U12147 (N_12147,N_9122,N_11017);
nand U12148 (N_12148,N_10822,N_11981);
xnor U12149 (N_12149,N_9249,N_11441);
nor U12150 (N_12150,N_10509,N_9748);
xor U12151 (N_12151,N_10133,N_10108);
nand U12152 (N_12152,N_9187,N_10159);
nand U12153 (N_12153,N_11148,N_9019);
xor U12154 (N_12154,N_9446,N_11466);
xnor U12155 (N_12155,N_10495,N_9538);
or U12156 (N_12156,N_11569,N_9580);
or U12157 (N_12157,N_10606,N_9681);
nand U12158 (N_12158,N_9858,N_10238);
and U12159 (N_12159,N_11570,N_11043);
nand U12160 (N_12160,N_9464,N_11739);
nand U12161 (N_12161,N_10747,N_10437);
and U12162 (N_12162,N_9246,N_10508);
or U12163 (N_12163,N_10123,N_10846);
nand U12164 (N_12164,N_9671,N_9086);
xnor U12165 (N_12165,N_10770,N_11064);
nand U12166 (N_12166,N_10206,N_9517);
nor U12167 (N_12167,N_9355,N_9907);
nor U12168 (N_12168,N_10915,N_11663);
nand U12169 (N_12169,N_10679,N_9418);
nand U12170 (N_12170,N_11410,N_11176);
and U12171 (N_12171,N_11220,N_10446);
or U12172 (N_12172,N_9029,N_9213);
and U12173 (N_12173,N_10654,N_9276);
and U12174 (N_12174,N_10082,N_9685);
and U12175 (N_12175,N_11893,N_11975);
and U12176 (N_12176,N_9118,N_11573);
nand U12177 (N_12177,N_10475,N_9665);
xnor U12178 (N_12178,N_11560,N_11478);
nand U12179 (N_12179,N_11950,N_10835);
and U12180 (N_12180,N_10917,N_10944);
nand U12181 (N_12181,N_9544,N_9547);
xnor U12182 (N_12182,N_11094,N_10496);
and U12183 (N_12183,N_11331,N_9723);
and U12184 (N_12184,N_9733,N_11375);
or U12185 (N_12185,N_10936,N_9986);
or U12186 (N_12186,N_10311,N_9150);
or U12187 (N_12187,N_9373,N_9166);
nand U12188 (N_12188,N_10357,N_11465);
and U12189 (N_12189,N_9930,N_10650);
nand U12190 (N_12190,N_9824,N_10847);
nand U12191 (N_12191,N_9007,N_11761);
and U12192 (N_12192,N_10797,N_10284);
or U12193 (N_12193,N_11257,N_9936);
nand U12194 (N_12194,N_9138,N_11666);
nand U12195 (N_12195,N_11356,N_9261);
or U12196 (N_12196,N_11386,N_9219);
xnor U12197 (N_12197,N_10072,N_9398);
or U12198 (N_12198,N_10296,N_10752);
or U12199 (N_12199,N_11665,N_11160);
nand U12200 (N_12200,N_9184,N_10757);
xor U12201 (N_12201,N_9821,N_11637);
nand U12202 (N_12202,N_10754,N_10833);
nand U12203 (N_12203,N_9744,N_11337);
nand U12204 (N_12204,N_11186,N_10498);
nand U12205 (N_12205,N_9758,N_11514);
nor U12206 (N_12206,N_9195,N_11594);
xnor U12207 (N_12207,N_9906,N_11768);
nand U12208 (N_12208,N_11908,N_11538);
and U12209 (N_12209,N_9766,N_10971);
and U12210 (N_12210,N_11306,N_10248);
xor U12211 (N_12211,N_11471,N_10968);
nor U12212 (N_12212,N_11134,N_11404);
nor U12213 (N_12213,N_10200,N_11883);
or U12214 (N_12214,N_9680,N_11677);
nand U12215 (N_12215,N_10708,N_11568);
xnor U12216 (N_12216,N_11693,N_9899);
or U12217 (N_12217,N_11928,N_9441);
nand U12218 (N_12218,N_11706,N_11624);
nor U12219 (N_12219,N_9975,N_11498);
nor U12220 (N_12220,N_11632,N_10838);
nand U12221 (N_12221,N_11870,N_10471);
nor U12222 (N_12222,N_11233,N_10441);
nor U12223 (N_12223,N_11434,N_9928);
nor U12224 (N_12224,N_10636,N_11686);
nand U12225 (N_12225,N_10622,N_11751);
nand U12226 (N_12226,N_11296,N_9473);
nor U12227 (N_12227,N_9776,N_9628);
nand U12228 (N_12228,N_11436,N_10331);
nand U12229 (N_12229,N_10089,N_9272);
xnor U12230 (N_12230,N_11213,N_9854);
and U12231 (N_12231,N_9755,N_11068);
and U12232 (N_12232,N_10360,N_11630);
or U12233 (N_12233,N_10756,N_9491);
nand U12234 (N_12234,N_10279,N_10949);
xnor U12235 (N_12235,N_10361,N_11991);
nand U12236 (N_12236,N_10420,N_10888);
xnor U12237 (N_12237,N_11104,N_9881);
nor U12238 (N_12238,N_10474,N_10407);
nand U12239 (N_12239,N_9672,N_9039);
nor U12240 (N_12240,N_10583,N_9478);
xor U12241 (N_12241,N_9395,N_9990);
nand U12242 (N_12242,N_9359,N_10596);
and U12243 (N_12243,N_9003,N_9726);
nand U12244 (N_12244,N_9005,N_9466);
or U12245 (N_12245,N_10644,N_9700);
nor U12246 (N_12246,N_10252,N_10669);
or U12247 (N_12247,N_9328,N_9429);
or U12248 (N_12248,N_11453,N_10004);
nand U12249 (N_12249,N_9516,N_10381);
nor U12250 (N_12250,N_10099,N_11584);
or U12251 (N_12251,N_9280,N_10353);
or U12252 (N_12252,N_10375,N_9677);
nor U12253 (N_12253,N_10488,N_9647);
xnor U12254 (N_12254,N_11237,N_10830);
nor U12255 (N_12255,N_9013,N_11370);
nand U12256 (N_12256,N_11865,N_11885);
nand U12257 (N_12257,N_9224,N_9574);
nand U12258 (N_12258,N_10176,N_11848);
xor U12259 (N_12259,N_9957,N_10641);
and U12260 (N_12260,N_9360,N_10380);
nand U12261 (N_12261,N_9052,N_11627);
or U12262 (N_12262,N_9616,N_9773);
xnor U12263 (N_12263,N_9049,N_10114);
or U12264 (N_12264,N_11959,N_9089);
xnor U12265 (N_12265,N_11185,N_9435);
nand U12266 (N_12266,N_9315,N_11869);
and U12267 (N_12267,N_9713,N_11565);
nor U12268 (N_12268,N_11966,N_9165);
nand U12269 (N_12269,N_10799,N_10952);
nor U12270 (N_12270,N_10713,N_9374);
and U12271 (N_12271,N_10691,N_10579);
and U12272 (N_12272,N_10686,N_11485);
nor U12273 (N_12273,N_10870,N_9509);
nor U12274 (N_12274,N_10751,N_11423);
nand U12275 (N_12275,N_9891,N_11641);
nand U12276 (N_12276,N_10303,N_10904);
or U12277 (N_12277,N_11360,N_10388);
or U12278 (N_12278,N_11860,N_10012);
nand U12279 (N_12279,N_11007,N_9633);
nor U12280 (N_12280,N_9286,N_11845);
xnor U12281 (N_12281,N_10092,N_10581);
nand U12282 (N_12282,N_9251,N_10077);
nor U12283 (N_12283,N_9695,N_10951);
and U12284 (N_12284,N_10963,N_11129);
nor U12285 (N_12285,N_10314,N_9849);
or U12286 (N_12286,N_9384,N_11174);
and U12287 (N_12287,N_9785,N_11184);
and U12288 (N_12288,N_10858,N_10027);
nand U12289 (N_12289,N_10439,N_11557);
nor U12290 (N_12290,N_11495,N_10947);
nand U12291 (N_12291,N_10955,N_10500);
xnor U12292 (N_12292,N_10919,N_10794);
and U12293 (N_12293,N_9771,N_9074);
and U12294 (N_12294,N_11506,N_9009);
nand U12295 (N_12295,N_11783,N_10371);
nor U12296 (N_12296,N_11652,N_11742);
xor U12297 (N_12297,N_11543,N_9402);
and U12298 (N_12298,N_10212,N_11578);
nor U12299 (N_12299,N_10170,N_9283);
or U12300 (N_12300,N_11793,N_10069);
xnor U12301 (N_12301,N_9708,N_11784);
nor U12302 (N_12302,N_11766,N_9918);
or U12303 (N_12303,N_9366,N_9867);
or U12304 (N_12304,N_10122,N_11203);
and U12305 (N_12305,N_9730,N_9266);
and U12306 (N_12306,N_9208,N_9277);
nor U12307 (N_12307,N_10544,N_10143);
nand U12308 (N_12308,N_10281,N_11754);
nor U12309 (N_12309,N_11261,N_9507);
and U12310 (N_12310,N_10511,N_11335);
nor U12311 (N_12311,N_11445,N_9400);
xnor U12312 (N_12312,N_10299,N_9793);
xor U12313 (N_12313,N_11446,N_11440);
nor U12314 (N_12314,N_11366,N_10154);
and U12315 (N_12315,N_11427,N_10646);
and U12316 (N_12316,N_10294,N_10487);
nor U12317 (N_12317,N_11956,N_9844);
xnor U12318 (N_12318,N_10050,N_11820);
or U12319 (N_12319,N_9238,N_9980);
and U12320 (N_12320,N_9977,N_10198);
or U12321 (N_12321,N_9556,N_9405);
nor U12322 (N_12322,N_10261,N_9307);
nor U12323 (N_12323,N_11399,N_11651);
or U12324 (N_12324,N_11164,N_11448);
nand U12325 (N_12325,N_10369,N_10249);
or U12326 (N_12326,N_10098,N_9444);
nor U12327 (N_12327,N_10706,N_9060);
or U12328 (N_12328,N_10773,N_9861);
nand U12329 (N_12329,N_10802,N_11143);
xor U12330 (N_12330,N_11026,N_11591);
or U12331 (N_12331,N_10406,N_10734);
nor U12332 (N_12332,N_10358,N_10860);
and U12333 (N_12333,N_11342,N_11486);
nor U12334 (N_12334,N_10672,N_11057);
and U12335 (N_12335,N_11469,N_10091);
xor U12336 (N_12336,N_11330,N_9893);
or U12337 (N_12337,N_10995,N_10486);
or U12338 (N_12338,N_9940,N_9645);
xnor U12339 (N_12339,N_9036,N_9324);
and U12340 (N_12340,N_9349,N_10324);
and U12341 (N_12341,N_9641,N_9869);
nor U12342 (N_12342,N_9088,N_11621);
xnor U12343 (N_12343,N_10183,N_9057);
and U12344 (N_12344,N_11348,N_11313);
and U12345 (N_12345,N_10710,N_10731);
nor U12346 (N_12346,N_9687,N_11190);
and U12347 (N_12347,N_11583,N_9186);
or U12348 (N_12348,N_9779,N_11241);
or U12349 (N_12349,N_10524,N_11121);
nand U12350 (N_12350,N_10259,N_11195);
xor U12351 (N_12351,N_9795,N_11294);
and U12352 (N_12352,N_9200,N_10430);
and U12353 (N_12353,N_9562,N_10810);
nor U12354 (N_12354,N_9226,N_11030);
xor U12355 (N_12355,N_11604,N_11045);
nor U12356 (N_12356,N_10676,N_9911);
nor U12357 (N_12357,N_11850,N_9391);
xnor U12358 (N_12358,N_9784,N_11837);
nand U12359 (N_12359,N_10759,N_9802);
and U12360 (N_12360,N_9637,N_10038);
xnor U12361 (N_12361,N_10827,N_9863);
xnor U12362 (N_12362,N_10116,N_10243);
nand U12363 (N_12363,N_9931,N_10807);
and U12364 (N_12364,N_11250,N_9356);
and U12365 (N_12365,N_11238,N_10855);
nor U12366 (N_12366,N_11738,N_10820);
xor U12367 (N_12367,N_11939,N_11704);
and U12368 (N_12368,N_11268,N_10871);
nand U12369 (N_12369,N_10269,N_11066);
or U12370 (N_12370,N_9119,N_9353);
and U12371 (N_12371,N_10954,N_10315);
or U12372 (N_12372,N_11253,N_10619);
xnor U12373 (N_12373,N_11004,N_10273);
xnor U12374 (N_12374,N_9185,N_10685);
nand U12375 (N_12375,N_10283,N_10872);
nand U12376 (N_12376,N_10244,N_9954);
nor U12377 (N_12377,N_11929,N_11669);
nor U12378 (N_12378,N_11882,N_11281);
nor U12379 (N_12379,N_11553,N_10384);
or U12380 (N_12380,N_10536,N_9476);
nand U12381 (N_12381,N_10044,N_9745);
or U12382 (N_12382,N_9045,N_11925);
nand U12383 (N_12383,N_11985,N_11600);
or U12384 (N_12384,N_11964,N_9629);
xor U12385 (N_12385,N_11125,N_9777);
xor U12386 (N_12386,N_9289,N_10516);
and U12387 (N_12387,N_9558,N_10885);
nand U12388 (N_12388,N_10916,N_9001);
nand U12389 (N_12389,N_11856,N_11033);
or U12390 (N_12390,N_10095,N_9115);
nand U12391 (N_12391,N_9241,N_11868);
and U12392 (N_12392,N_10997,N_10503);
and U12393 (N_12393,N_11472,N_9270);
xor U12394 (N_12394,N_9590,N_11530);
nand U12395 (N_12395,N_10633,N_10841);
nand U12396 (N_12396,N_11177,N_11806);
and U12397 (N_12397,N_9818,N_11921);
xor U12398 (N_12398,N_11886,N_9031);
xnor U12399 (N_12399,N_11249,N_10484);
nor U12400 (N_12400,N_10317,N_10559);
nand U12401 (N_12401,N_11863,N_9508);
and U12402 (N_12402,N_9050,N_10566);
nand U12403 (N_12403,N_9069,N_11451);
and U12404 (N_12404,N_11903,N_11531);
or U12405 (N_12405,N_9703,N_11232);
nand U12406 (N_12406,N_9024,N_11914);
or U12407 (N_12407,N_10340,N_10832);
nor U12408 (N_12408,N_9063,N_11214);
nor U12409 (N_12409,N_10643,N_11101);
nor U12410 (N_12410,N_11502,N_11524);
or U12411 (N_12411,N_11070,N_10921);
nand U12412 (N_12412,N_11271,N_11403);
or U12413 (N_12413,N_11659,N_11229);
nand U12414 (N_12414,N_9305,N_9386);
and U12415 (N_12415,N_11727,N_10093);
or U12416 (N_12416,N_10712,N_11973);
xor U12417 (N_12417,N_9656,N_9260);
nand U12418 (N_12418,N_10873,N_11607);
nand U12419 (N_12419,N_11291,N_10236);
nand U12420 (N_12420,N_11785,N_10527);
or U12421 (N_12421,N_9162,N_9719);
and U12422 (N_12422,N_11599,N_9904);
nor U12423 (N_12423,N_10842,N_9675);
nor U12424 (N_12424,N_11915,N_9743);
xor U12425 (N_12425,N_11936,N_9340);
nor U12426 (N_12426,N_9878,N_9164);
and U12427 (N_12427,N_11954,N_10856);
or U12428 (N_12428,N_9593,N_10704);
nor U12429 (N_12429,N_10137,N_11483);
xor U12430 (N_12430,N_11499,N_9458);
nor U12431 (N_12431,N_10151,N_10352);
nand U12432 (N_12432,N_9919,N_10615);
or U12433 (N_12433,N_10808,N_11831);
nor U12434 (N_12434,N_9104,N_9857);
xor U12435 (N_12435,N_9976,N_11456);
nand U12436 (N_12436,N_9668,N_11264);
nand U12437 (N_12437,N_10033,N_9525);
nand U12438 (N_12438,N_9523,N_9939);
and U12439 (N_12439,N_9984,N_11084);
or U12440 (N_12440,N_10863,N_11857);
nand U12441 (N_12441,N_10094,N_9447);
or U12442 (N_12442,N_10603,N_11273);
nor U12443 (N_12443,N_10339,N_9738);
nand U12444 (N_12444,N_11039,N_9111);
nor U12445 (N_12445,N_11522,N_11254);
or U12446 (N_12446,N_11369,N_9440);
nand U12447 (N_12447,N_10629,N_9659);
and U12448 (N_12448,N_11943,N_11512);
xnor U12449 (N_12449,N_10749,N_10745);
nand U12450 (N_12450,N_11332,N_10974);
or U12451 (N_12451,N_10001,N_9876);
nand U12452 (N_12452,N_10798,N_11178);
and U12453 (N_12453,N_10080,N_10653);
or U12454 (N_12454,N_9434,N_10923);
nor U12455 (N_12455,N_11123,N_10534);
and U12456 (N_12456,N_10229,N_11617);
or U12457 (N_12457,N_9674,N_11697);
nand U12458 (N_12458,N_9715,N_10829);
or U12459 (N_12459,N_11887,N_9459);
nand U12460 (N_12460,N_9564,N_10909);
nand U12461 (N_12461,N_11338,N_11794);
xor U12462 (N_12462,N_10702,N_9573);
nor U12463 (N_12463,N_9942,N_11226);
xor U12464 (N_12464,N_11119,N_11259);
or U12465 (N_12465,N_9650,N_10163);
nor U12466 (N_12466,N_11152,N_10161);
nand U12467 (N_12467,N_11829,N_9790);
or U12468 (N_12468,N_10586,N_9048);
xor U12469 (N_12469,N_9624,N_11089);
xor U12470 (N_12470,N_11192,N_9727);
nand U12471 (N_12471,N_11408,N_10320);
nor U12472 (N_12472,N_11609,N_11668);
or U12473 (N_12473,N_9883,N_11818);
xor U12474 (N_12474,N_10409,N_10592);
and U12475 (N_12475,N_9946,N_11136);
nand U12476 (N_12476,N_9998,N_11135);
nand U12477 (N_12477,N_9910,N_10323);
nor U12478 (N_12478,N_10996,N_9181);
xnor U12479 (N_12479,N_11307,N_11080);
nor U12480 (N_12480,N_11895,N_9462);
xnor U12481 (N_12481,N_10378,N_10518);
xor U12482 (N_12482,N_11655,N_10466);
or U12483 (N_12483,N_9034,N_10631);
nand U12484 (N_12484,N_11405,N_10552);
nand U12485 (N_12485,N_11800,N_11635);
and U12486 (N_12486,N_10760,N_10288);
and U12487 (N_12487,N_11679,N_9787);
nor U12488 (N_12488,N_9064,N_9248);
or U12489 (N_12489,N_10325,N_9643);
and U12490 (N_12490,N_9722,N_9518);
or U12491 (N_12491,N_11963,N_9252);
nand U12492 (N_12492,N_9413,N_11798);
and U12493 (N_12493,N_9520,N_10998);
xnor U12494 (N_12494,N_9401,N_11960);
or U12495 (N_12495,N_10432,N_11830);
nor U12496 (N_12496,N_9684,N_11020);
or U12497 (N_12497,N_11443,N_10876);
nor U12498 (N_12498,N_9683,N_10233);
nand U12499 (N_12499,N_9171,N_10567);
nor U12500 (N_12500,N_9382,N_10698);
xnor U12501 (N_12501,N_11816,N_11646);
nand U12502 (N_12502,N_10550,N_11023);
or U12503 (N_12503,N_9669,N_10359);
and U12504 (N_12504,N_9339,N_10349);
xor U12505 (N_12505,N_10533,N_11899);
nand U12506 (N_12506,N_9416,N_11740);
xor U12507 (N_12507,N_9847,N_11090);
nand U12508 (N_12508,N_10861,N_11319);
xnor U12509 (N_12509,N_10160,N_10035);
nand U12510 (N_12510,N_11803,N_11111);
xor U12511 (N_12511,N_10213,N_10239);
and U12512 (N_12512,N_9090,N_10113);
xnor U12513 (N_12513,N_9310,N_11086);
nand U12514 (N_12514,N_11349,N_10582);
and U12515 (N_12515,N_11207,N_9900);
nor U12516 (N_12516,N_11095,N_10665);
or U12517 (N_12517,N_11329,N_9194);
nand U12518 (N_12518,N_11381,N_11799);
xnor U12519 (N_12519,N_10345,N_11696);
nand U12520 (N_12520,N_11059,N_9354);
or U12521 (N_12521,N_10040,N_11994);
or U12522 (N_12522,N_9113,N_11384);
or U12523 (N_12523,N_10542,N_11563);
nand U12524 (N_12524,N_9761,N_10701);
nor U12525 (N_12525,N_9649,N_10118);
nand U12526 (N_12526,N_9096,N_10156);
nor U12527 (N_12527,N_10984,N_10121);
xnor U12528 (N_12528,N_10966,N_9542);
or U12529 (N_12529,N_9667,N_10455);
nor U12530 (N_12530,N_9321,N_10945);
or U12531 (N_12531,N_9944,N_9581);
and U12532 (N_12532,N_11723,N_10307);
nor U12533 (N_12533,N_10621,N_9425);
and U12534 (N_12534,N_10301,N_11415);
or U12535 (N_12535,N_11496,N_10058);
nand U12536 (N_12536,N_9421,N_11292);
xnor U12537 (N_12537,N_10298,N_9526);
nor U12538 (N_12538,N_10514,N_11374);
nor U12539 (N_12539,N_9160,N_9439);
xnor U12540 (N_12540,N_9091,N_10313);
nand U12541 (N_12541,N_9613,N_9157);
xor U12542 (N_12542,N_10363,N_11367);
xor U12543 (N_12543,N_11912,N_10059);
or U12544 (N_12544,N_10730,N_11935);
or U12545 (N_12545,N_11425,N_10649);
or U12546 (N_12546,N_11222,N_10472);
xnor U12547 (N_12547,N_10986,N_11289);
nand U12548 (N_12548,N_10755,N_9999);
and U12549 (N_12549,N_10482,N_9596);
xor U12550 (N_12550,N_9410,N_9548);
xor U12551 (N_12551,N_9365,N_10196);
nand U12552 (N_12552,N_9094,N_10933);
nor U12553 (N_12553,N_9720,N_9485);
nand U12554 (N_12554,N_10920,N_9499);
and U12555 (N_12555,N_10939,N_10883);
or U12556 (N_12556,N_9460,N_11900);
and U12557 (N_12557,N_10992,N_9066);
nand U12558 (N_12558,N_10836,N_11283);
nor U12559 (N_12559,N_11299,N_11755);
nand U12560 (N_12560,N_9173,N_10043);
xor U12561 (N_12561,N_9909,N_10401);
or U12562 (N_12562,N_9679,N_10785);
xnor U12563 (N_12563,N_11083,N_11246);
nor U12564 (N_12564,N_10535,N_11206);
nor U12565 (N_12565,N_9409,N_10102);
nand U12566 (N_12566,N_11418,N_10418);
xnor U12567 (N_12567,N_11519,N_11357);
nor U12568 (N_12568,N_10167,N_9490);
xor U12569 (N_12569,N_11544,N_10410);
xnor U12570 (N_12570,N_10193,N_9725);
nor U12571 (N_12571,N_9541,N_9303);
xnor U12572 (N_12572,N_10899,N_11351);
or U12573 (N_12573,N_10087,N_11324);
xnor U12574 (N_12574,N_9915,N_11449);
and U12575 (N_12575,N_10744,N_11756);
and U12576 (N_12576,N_10424,N_10814);
nand U12577 (N_12577,N_9970,N_9297);
nor U12578 (N_12578,N_10383,N_9664);
or U12579 (N_12579,N_9080,N_9497);
and U12580 (N_12580,N_10898,N_9461);
nor U12581 (N_12581,N_11682,N_11721);
nor U12582 (N_12582,N_9000,N_11154);
or U12583 (N_12583,N_9100,N_10703);
and U12584 (N_12584,N_9579,N_9626);
and U12585 (N_12585,N_10460,N_9159);
and U12586 (N_12586,N_9230,N_9189);
xor U12587 (N_12587,N_10975,N_11703);
nor U12588 (N_12588,N_10073,N_9619);
or U12589 (N_12589,N_10031,N_11139);
and U12590 (N_12590,N_10746,N_10985);
nand U12591 (N_12591,N_9250,N_10609);
or U12592 (N_12592,N_10548,N_11662);
and U12593 (N_12593,N_11055,N_9422);
or U12594 (N_12594,N_10707,N_10427);
nand U12595 (N_12595,N_10002,N_9570);
nand U12596 (N_12596,N_10519,N_9960);
xor U12597 (N_12597,N_11416,N_10448);
and U12598 (N_12598,N_9196,N_9135);
nor U12599 (N_12599,N_10926,N_10505);
and U12600 (N_12600,N_10819,N_10573);
nand U12601 (N_12601,N_10391,N_11767);
or U12602 (N_12602,N_10209,N_11024);
nand U12603 (N_12603,N_11128,N_10718);
nand U12604 (N_12604,N_9319,N_11093);
and U12605 (N_12605,N_9933,N_11072);
or U12606 (N_12606,N_11158,N_10119);
nor U12607 (N_12607,N_10101,N_9914);
and U12608 (N_12608,N_10738,N_11802);
nor U12609 (N_12609,N_9146,N_9823);
and U12610 (N_12610,N_11690,N_9530);
xnor U12611 (N_12611,N_9463,N_11618);
and U12612 (N_12612,N_11695,N_10918);
xnor U12613 (N_12613,N_10389,N_9482);
nand U12614 (N_12614,N_9934,N_10396);
or U12615 (N_12615,N_11505,N_11776);
nor U12616 (N_12616,N_9145,N_10927);
nor U12617 (N_12617,N_11952,N_9979);
nand U12618 (N_12618,N_9134,N_10452);
nand U12619 (N_12619,N_11710,N_9799);
nor U12620 (N_12620,N_11781,N_10683);
nand U12621 (N_12621,N_9533,N_11488);
nor U12622 (N_12622,N_11537,N_9972);
or U12623 (N_12623,N_10150,N_10379);
or U12624 (N_12624,N_10664,N_11320);
or U12625 (N_12625,N_9183,N_10115);
nor U12626 (N_12626,N_10271,N_11013);
or U12627 (N_12627,N_10066,N_11224);
or U12628 (N_12628,N_11156,N_11293);
nor U12629 (N_12629,N_11122,N_10595);
nand U12630 (N_12630,N_9948,N_10197);
nand U12631 (N_12631,N_9792,N_10494);
nor U12632 (N_12632,N_11096,N_9655);
nand U12633 (N_12633,N_9351,N_11518);
or U12634 (N_12634,N_10210,N_11881);
and U12635 (N_12635,N_11796,N_10659);
nand U12636 (N_12636,N_10364,N_9336);
nand U12637 (N_12637,N_11476,N_9287);
nand U12638 (N_12638,N_9670,N_11521);
nor U12639 (N_12639,N_9594,N_9731);
nand U12640 (N_12640,N_10131,N_9759);
nor U12641 (N_12641,N_11464,N_10616);
nor U12642 (N_12642,N_10791,N_11534);
and U12643 (N_12643,N_9612,N_11942);
nor U12644 (N_12644,N_11658,N_9232);
nand U12645 (N_12645,N_9588,N_10848);
nor U12646 (N_12646,N_10171,N_11576);
and U12647 (N_12647,N_10761,N_10781);
xor U12648 (N_12648,N_11694,N_9896);
or U12649 (N_12649,N_11316,N_11841);
xor U12650 (N_12650,N_10561,N_9584);
and U12651 (N_12651,N_11684,N_11795);
nor U12652 (N_12652,N_9583,N_9965);
nor U12653 (N_12653,N_10967,N_9403);
nor U12654 (N_12654,N_11631,N_9103);
and U12655 (N_12655,N_11194,N_11725);
xnor U12656 (N_12656,N_10220,N_11181);
xor U12657 (N_12657,N_9428,N_11972);
and U12658 (N_12658,N_11874,N_10877);
or U12659 (N_12659,N_10890,N_11718);
and U12660 (N_12660,N_10563,N_9267);
and U12661 (N_12661,N_9231,N_10127);
nand U12662 (N_12662,N_10185,N_10221);
xnor U12663 (N_12663,N_9329,N_9312);
and U12664 (N_12664,N_11620,N_11993);
or U12665 (N_12665,N_10019,N_10800);
nand U12666 (N_12666,N_10668,N_10735);
or U12667 (N_12667,N_11166,N_11219);
nor U12668 (N_12668,N_10577,N_11660);
nand U12669 (N_12669,N_11006,N_9658);
nand U12670 (N_12670,N_11044,N_11817);
or U12671 (N_12671,N_11873,N_9553);
nand U12672 (N_12672,N_10652,N_10117);
nor U12673 (N_12673,N_11601,N_11309);
xor U12674 (N_12674,N_11523,N_10289);
nand U12675 (N_12675,N_11577,N_9245);
and U12676 (N_12676,N_10392,N_10158);
nor U12677 (N_12677,N_9452,N_9767);
nand U12678 (N_12678,N_10640,N_11140);
nand U12679 (N_12679,N_11571,N_9102);
nand U12680 (N_12680,N_11150,N_11813);
nor U12681 (N_12681,N_9663,N_11113);
nor U12682 (N_12682,N_9108,N_9749);
or U12683 (N_12683,N_10681,N_10768);
nand U12684 (N_12684,N_9527,N_11957);
or U12685 (N_12685,N_11183,N_9468);
and U12686 (N_12686,N_10493,N_9436);
and U12687 (N_12687,N_10417,N_10232);
nor U12688 (N_12688,N_9712,N_9314);
nor U12689 (N_12689,N_10034,N_10911);
and U12690 (N_12690,N_11133,N_9742);
or U12691 (N_12691,N_9474,N_9147);
nor U12692 (N_12692,N_9498,N_11714);
xor U12693 (N_12693,N_11990,N_11012);
and U12694 (N_12694,N_10290,N_11872);
xnor U12695 (N_12695,N_9012,N_11851);
or U12696 (N_12696,N_9431,N_9285);
nand U12697 (N_12697,N_9961,N_11737);
or U12698 (N_12698,N_11048,N_11170);
or U12699 (N_12699,N_9804,N_11838);
or U12700 (N_12700,N_11201,N_9851);
nand U12701 (N_12701,N_11566,N_9550);
nand U12702 (N_12702,N_9750,N_11252);
xor U12703 (N_12703,N_11221,N_11974);
nor U12704 (N_12704,N_11234,N_10057);
nor U12705 (N_12705,N_11517,N_11826);
nor U12706 (N_12706,N_11535,N_11529);
nor U12707 (N_12707,N_10018,N_10766);
nor U12708 (N_12708,N_9028,N_11681);
nand U12709 (N_12709,N_11454,N_9775);
nand U12710 (N_12710,N_11269,N_11877);
xor U12711 (N_12711,N_11500,N_9567);
and U12712 (N_12712,N_9692,N_11979);
and U12713 (N_12713,N_9197,N_9618);
xnor U12714 (N_12714,N_10147,N_11462);
xnor U12715 (N_12715,N_9652,N_10610);
nor U12716 (N_12716,N_10786,N_10857);
nand U12717 (N_12717,N_10667,N_9264);
nand U12718 (N_12718,N_10684,N_10136);
nor U12719 (N_12719,N_11243,N_11396);
xor U12720 (N_12720,N_11482,N_10149);
and U12721 (N_12721,N_10520,N_10242);
and U12722 (N_12722,N_10399,N_11824);
nand U12723 (N_12723,N_9813,N_11318);
and U12724 (N_12724,N_9874,N_11236);
xnor U12725 (N_12725,N_9833,N_9158);
xor U12726 (N_12726,N_9780,N_10912);
or U12727 (N_12727,N_10881,N_10742);
and U12728 (N_12728,N_11173,N_9505);
or U12729 (N_12729,N_9617,N_9639);
nand U12730 (N_12730,N_11388,N_9582);
and U12731 (N_12731,N_11142,N_9870);
or U12732 (N_12732,N_10400,N_10587);
or U12733 (N_12733,N_10697,N_10591);
nor U12734 (N_12734,N_9521,N_9177);
or U12735 (N_12735,N_9622,N_9112);
or U12736 (N_12736,N_9335,N_9117);
nor U12737 (N_12737,N_9654,N_11027);
nand U12738 (N_12738,N_9805,N_9500);
nand U12739 (N_12739,N_11759,N_10032);
and U12740 (N_12740,N_11540,N_10138);
or U12741 (N_12741,N_10864,N_10696);
or U12742 (N_12742,N_9534,N_10943);
nand U12743 (N_12743,N_10447,N_11492);
nand U12744 (N_12744,N_9337,N_9532);
and U12745 (N_12745,N_9827,N_10020);
or U12746 (N_12746,N_10465,N_10617);
and U12747 (N_12747,N_10513,N_9008);
nor U12748 (N_12748,N_9554,N_10433);
and U12749 (N_12749,N_9873,N_10230);
and U12750 (N_12750,N_11005,N_11216);
or U12751 (N_12751,N_11716,N_9244);
and U12752 (N_12752,N_10199,N_9424);
or U12753 (N_12753,N_11711,N_11431);
or U12754 (N_12754,N_10913,N_10190);
xor U12755 (N_12755,N_10957,N_10451);
nor U12756 (N_12756,N_11497,N_9222);
or U12757 (N_12757,N_11533,N_11504);
and U12758 (N_12758,N_11944,N_10999);
nand U12759 (N_12759,N_9133,N_11000);
or U12760 (N_12760,N_11352,N_10461);
and U12761 (N_12761,N_9769,N_11373);
or U12762 (N_12762,N_10673,N_11968);
or U12763 (N_12763,N_10546,N_11402);
or U12764 (N_12764,N_11778,N_9974);
nor U12765 (N_12765,N_10727,N_9717);
or U12766 (N_12766,N_9577,N_9815);
and U12767 (N_12767,N_10134,N_10246);
or U12768 (N_12768,N_11467,N_10721);
nand U12769 (N_12769,N_10840,N_11452);
xor U12770 (N_12770,N_9950,N_10788);
nand U12771 (N_12771,N_10688,N_11474);
nand U12772 (N_12772,N_10282,N_11589);
xnor U12773 (N_12773,N_9334,N_10110);
nand U12774 (N_12774,N_10585,N_11003);
nand U12775 (N_12775,N_11597,N_10964);
xor U12776 (N_12776,N_10796,N_11364);
and U12777 (N_12777,N_9894,N_9085);
nor U12778 (N_12778,N_9389,N_9638);
xnor U12779 (N_12779,N_10571,N_10009);
and U12780 (N_12780,N_11484,N_10556);
or U12781 (N_12781,N_10969,N_9798);
and U12782 (N_12782,N_10402,N_9644);
nor U12783 (N_12783,N_9451,N_11145);
and U12784 (N_12784,N_10560,N_10908);
or U12785 (N_12785,N_10010,N_10343);
and U12786 (N_12786,N_9819,N_11391);
nand U12787 (N_12787,N_9606,N_11554);
or U12788 (N_12788,N_11790,N_11671);
or U12789 (N_12789,N_9586,N_10485);
or U12790 (N_12790,N_11109,N_9831);
or U12791 (N_12791,N_10584,N_10090);
nor U12792 (N_12792,N_11720,N_11564);
nand U12793 (N_12793,N_9615,N_11804);
and U12794 (N_12794,N_10694,N_10977);
and U12795 (N_12795,N_10541,N_10739);
nor U12796 (N_12796,N_11223,N_11018);
xnor U12797 (N_12797,N_11341,N_10907);
nor U12798 (N_12798,N_9699,N_9506);
nor U12799 (N_12799,N_11989,N_9994);
nor U12800 (N_12800,N_11955,N_10231);
nand U12801 (N_12801,N_11582,N_11769);
nand U12802 (N_12802,N_11722,N_11475);
nor U12803 (N_12803,N_9363,N_10411);
nand U12804 (N_12804,N_9774,N_9243);
and U12805 (N_12805,N_9912,N_9754);
nor U12806 (N_12806,N_10423,N_10007);
or U12807 (N_12807,N_9437,N_9322);
or U12808 (N_12808,N_11225,N_10790);
and U12809 (N_12809,N_11394,N_9981);
nor U12810 (N_12810,N_11340,N_9772);
xnor U12811 (N_12811,N_10086,N_10714);
nand U12812 (N_12812,N_10347,N_9913);
and U12813 (N_12813,N_10562,N_10978);
or U12814 (N_12814,N_11385,N_11733);
and U12815 (N_12815,N_10950,N_9292);
xnor U12816 (N_12816,N_10333,N_9689);
nand U12817 (N_12817,N_11734,N_11315);
or U12818 (N_12818,N_11525,N_10189);
and U12819 (N_12819,N_10074,N_11053);
or U12820 (N_12820,N_10981,N_9714);
nor U12821 (N_12821,N_10666,N_10264);
and U12822 (N_12822,N_9129,N_11719);
and U12823 (N_12823,N_11477,N_9371);
or U12824 (N_12824,N_10792,N_10601);
xor U12825 (N_12825,N_11147,N_9607);
and U12826 (N_12826,N_11311,N_11644);
and U12827 (N_12827,N_11562,N_11992);
nand U12828 (N_12828,N_10191,N_11067);
nor U12829 (N_12829,N_9149,N_9598);
nor U12830 (N_12830,N_9414,N_10293);
and U12831 (N_12831,N_10517,N_10155);
or U12832 (N_12832,N_10859,N_11235);
nand U12833 (N_12833,N_10085,N_11547);
xnor U12834 (N_12834,N_11163,N_10055);
nand U12835 (N_12835,N_11276,N_9884);
and U12836 (N_12836,N_10036,N_11439);
nor U12837 (N_12837,N_9540,N_9797);
or U12838 (N_12838,N_11035,N_9740);
xnor U12839 (N_12839,N_10663,N_9123);
and U12840 (N_12840,N_11077,N_9288);
and U12841 (N_12841,N_9346,N_10960);
nor U12842 (N_12842,N_10588,N_9380);
or U12843 (N_12843,N_11909,N_10207);
and U12844 (N_12844,N_9067,N_11746);
or U12845 (N_12845,N_10607,N_9204);
or U12846 (N_12846,N_10817,N_11948);
nand U12847 (N_12847,N_10778,N_9988);
nor U12848 (N_12848,N_11390,N_11159);
or U12849 (N_12849,N_9566,N_10724);
nor U12850 (N_12850,N_11429,N_10895);
or U12851 (N_12851,N_9011,N_11932);
xnor U12852 (N_12852,N_11513,N_9101);
or U12853 (N_12853,N_9174,N_9153);
and U12854 (N_12854,N_10549,N_9809);
nor U12855 (N_12855,N_10130,N_10112);
and U12856 (N_12856,N_9483,N_10490);
nand U12857 (N_12857,N_9621,N_9661);
and U12858 (N_12858,N_10733,N_10105);
or U12859 (N_12859,N_10302,N_9640);
and U12860 (N_12860,N_11653,N_9136);
nor U12861 (N_12861,N_11210,N_11917);
xor U12862 (N_12862,N_11215,N_11622);
or U12863 (N_12863,N_10228,N_11779);
or U12864 (N_12864,N_10726,N_10319);
or U12865 (N_12865,N_10373,N_11859);
nor U12866 (N_12866,N_10047,N_9106);
and U12867 (N_12867,N_10103,N_10880);
and U12868 (N_12868,N_9651,N_10891);
nand U12869 (N_12869,N_9099,N_9239);
nand U12870 (N_12870,N_11061,N_10598);
nor U12871 (N_12871,N_11847,N_11258);
and U12872 (N_12872,N_9828,N_11782);
nand U12873 (N_12873,N_10088,N_9037);
nor U12874 (N_12874,N_11353,N_9110);
and U12875 (N_12875,N_11982,N_9215);
or U12876 (N_12876,N_11433,N_11606);
and U12877 (N_12877,N_9800,N_11409);
nor U12878 (N_12878,N_10097,N_11832);
or U12879 (N_12879,N_10262,N_11654);
nor U12880 (N_12880,N_10910,N_9923);
nand U12881 (N_12881,N_10024,N_10692);
nand U12882 (N_12882,N_10211,N_9411);
or U12883 (N_12883,N_10215,N_9922);
xnor U12884 (N_12884,N_9486,N_9093);
or U12885 (N_12885,N_11777,N_9120);
xnor U12886 (N_12886,N_11970,N_9926);
and U12887 (N_12887,N_9376,N_10026);
and U12888 (N_12888,N_10382,N_11301);
nand U12889 (N_12889,N_10204,N_9565);
xor U12890 (N_12890,N_11074,N_11633);
or U12891 (N_12891,N_11082,N_9317);
xor U12892 (N_12892,N_10554,N_9764);
nor U12893 (N_12893,N_11626,N_11421);
nand U12894 (N_12894,N_10266,N_11419);
nand U12895 (N_12895,N_10039,N_9492);
nor U12896 (N_12896,N_11011,N_9741);
or U12897 (N_12897,N_9273,N_11447);
nor U12898 (N_12898,N_10062,N_11730);
nor U12899 (N_12899,N_9599,N_10504);
nand U12900 (N_12900,N_10852,N_10709);
nor U12901 (N_12901,N_9290,N_9806);
nand U12902 (N_12902,N_10661,N_9348);
and U12903 (N_12903,N_9058,N_9890);
nand U12904 (N_12904,N_11032,N_11843);
xor U12905 (N_12905,N_9282,N_9387);
xnor U12906 (N_12906,N_11106,N_9331);
or U12907 (N_12907,N_9545,N_11852);
nand U12908 (N_12908,N_11678,N_10234);
or U12909 (N_12909,N_10732,N_11598);
and U12910 (N_12910,N_10386,N_9379);
and U12911 (N_12911,N_10292,N_10783);
nand U12912 (N_12912,N_11267,N_10270);
or U12913 (N_12913,N_11801,N_9614);
and U12914 (N_12914,N_11541,N_11854);
xnor U12915 (N_12915,N_11247,N_9298);
nand U12916 (N_12916,N_11999,N_11362);
nand U12917 (N_12917,N_9837,N_11536);
and U12918 (N_12918,N_9569,N_10993);
nor U12919 (N_12919,N_9381,N_11894);
or U12920 (N_12920,N_9163,N_9514);
and U12921 (N_12921,N_10805,N_9291);
xor U12922 (N_12922,N_11649,N_10599);
or U12923 (N_12923,N_10953,N_10256);
and U12924 (N_12924,N_10295,N_10777);
nand U12925 (N_12925,N_9350,N_9318);
nand U12926 (N_12926,N_10862,N_11110);
xnor U12927 (N_12927,N_11432,N_9555);
or U12928 (N_12928,N_9557,N_10845);
nand U12929 (N_12929,N_10056,N_11372);
or U12930 (N_12930,N_10458,N_10914);
nand U12931 (N_12931,N_10551,N_9991);
or U12932 (N_12932,N_11918,N_11265);
nand U12933 (N_12933,N_10687,N_10241);
nand U12934 (N_12934,N_9477,N_10416);
and U12935 (N_12935,N_9207,N_9151);
nor U12936 (N_12936,N_9941,N_9571);
nand U12937 (N_12937,N_10310,N_9589);
and U12938 (N_12938,N_11732,N_10982);
nor U12939 (N_12939,N_10811,N_11034);
xnor U12940 (N_12940,N_9887,N_11840);
or U12941 (N_12941,N_9201,N_11274);
xnor U12942 (N_12942,N_11656,N_9778);
and U12943 (N_12943,N_11945,N_11480);
xnor U12944 (N_12944,N_11593,N_11028);
xnor U12945 (N_12945,N_9313,N_11670);
or U12946 (N_12946,N_10868,N_10368);
xnor U12947 (N_12947,N_9816,N_11546);
and U12948 (N_12948,N_11988,N_10332);
and U12949 (N_12949,N_11042,N_9097);
nand U12950 (N_12950,N_11892,N_9646);
xor U12951 (N_12951,N_10897,N_10973);
nand U12952 (N_12952,N_10306,N_10285);
xor U12953 (N_12953,N_10879,N_11595);
or U12954 (N_12954,N_9495,N_9682);
nand U12955 (N_12955,N_9592,N_11673);
xor U12956 (N_12956,N_10729,N_10084);
nor U12957 (N_12957,N_9501,N_9188);
nand U12958 (N_12958,N_11002,N_11073);
and U12959 (N_12959,N_11650,N_11808);
and U12960 (N_12960,N_11172,N_11336);
nor U12961 (N_12961,N_9959,N_11297);
nand U12962 (N_12962,N_10444,N_9531);
nand U12963 (N_12963,N_9632,N_9055);
and U12964 (N_12964,N_11205,N_9973);
or U12965 (N_12965,N_9234,N_11961);
xnor U12966 (N_12966,N_11287,N_9077);
xor U12967 (N_12967,N_9666,N_9789);
or U12968 (N_12968,N_11834,N_11647);
or U12969 (N_12969,N_11151,N_11919);
and U12970 (N_12970,N_11031,N_11085);
xnor U12971 (N_12971,N_9076,N_9330);
xor U12972 (N_12972,N_11619,N_11712);
nor U12973 (N_12973,N_11155,N_10403);
nand U12974 (N_12974,N_9892,N_11551);
xnor U12975 (N_12975,N_10568,N_9059);
xor U12976 (N_12976,N_11260,N_9803);
xnor U12977 (N_12977,N_9636,N_9983);
nor U12978 (N_12978,N_9392,N_10784);
nand U12979 (N_12979,N_9205,N_10000);
nand U12980 (N_12980,N_11334,N_10374);
and U12981 (N_12981,N_9630,N_10637);
xor U12982 (N_12982,N_10575,N_9768);
nor U12983 (N_12983,N_10844,N_10247);
or U12984 (N_12984,N_11702,N_10612);
xnor U12985 (N_12985,N_9484,N_9227);
and U12986 (N_12986,N_10545,N_10976);
and U12987 (N_12987,N_10278,N_9898);
or U12988 (N_12988,N_9927,N_10245);
or U12989 (N_12989,N_10741,N_10787);
nor U12990 (N_12990,N_11494,N_10935);
xor U12991 (N_12991,N_11460,N_9860);
and U12992 (N_12992,N_10837,N_10419);
xnor U12993 (N_12993,N_9127,N_11603);
and U12994 (N_12994,N_11747,N_11969);
and U12995 (N_12995,N_11958,N_10674);
xor U12996 (N_12996,N_11825,N_11197);
xnor U12997 (N_12997,N_9853,N_10179);
nor U12998 (N_12998,N_10395,N_11198);
and U12999 (N_12999,N_11661,N_10608);
nor U13000 (N_13000,N_9061,N_11387);
nand U13001 (N_13001,N_11314,N_11511);
nor U13002 (N_13002,N_9513,N_11811);
and U13003 (N_13003,N_9559,N_9073);
and U13004 (N_13004,N_10670,N_11016);
nor U13005 (N_13005,N_9522,N_11412);
xnor U13006 (N_13006,N_10438,N_9877);
or U13007 (N_13007,N_11949,N_11355);
xor U13008 (N_13008,N_11008,N_9047);
or U13009 (N_13009,N_9210,N_11765);
or U13010 (N_13010,N_11520,N_11208);
or U13011 (N_13011,N_9167,N_11559);
or U13012 (N_13012,N_10824,N_10590);
and U13013 (N_13013,N_10793,N_11088);
nor U13014 (N_13014,N_9889,N_10886);
and U13015 (N_13015,N_9829,N_9442);
xor U13016 (N_13016,N_10224,N_10815);
nand U13017 (N_13017,N_11916,N_11266);
nand U13018 (N_13018,N_9465,N_10605);
nand U13019 (N_13019,N_9015,N_10801);
xor U13020 (N_13020,N_11978,N_11812);
nor U13021 (N_13021,N_11153,N_11014);
and U13022 (N_13022,N_11108,N_10989);
xnor U13023 (N_13023,N_9021,N_10250);
nand U13024 (N_13024,N_10570,N_10940);
or U13025 (N_13025,N_10626,N_11983);
and U13026 (N_13026,N_11438,N_10651);
or U13027 (N_13027,N_9605,N_10569);
nand U13028 (N_13028,N_11228,N_11898);
and U13029 (N_13029,N_9765,N_9469);
xnor U13030 (N_13030,N_9479,N_9218);
and U13031 (N_13031,N_10678,N_10928);
nand U13032 (N_13032,N_9587,N_9952);
xor U13033 (N_13033,N_9840,N_10078);
nand U13034 (N_13034,N_10510,N_9125);
nor U13035 (N_13035,N_10547,N_11371);
and U13036 (N_13036,N_9826,N_10930);
and U13037 (N_13037,N_10146,N_9762);
and U13038 (N_13038,N_9406,N_9438);
nor U13039 (N_13039,N_11288,N_9427);
nor U13040 (N_13040,N_11822,N_11050);
or U13041 (N_13041,N_10538,N_11354);
xor U13042 (N_13042,N_10141,N_9399);
xnor U13043 (N_13043,N_9390,N_10717);
or U13044 (N_13044,N_10483,N_9536);
xnor U13045 (N_13045,N_9496,N_9841);
xor U13046 (N_13046,N_11062,N_9964);
and U13047 (N_13047,N_11907,N_9450);
xor U13048 (N_13048,N_11797,N_11100);
nand U13049 (N_13049,N_9997,N_9126);
nand U13050 (N_13050,N_10440,N_11457);
xor U13051 (N_13051,N_9595,N_10344);
or U13052 (N_13052,N_10894,N_9068);
and U13053 (N_13053,N_9987,N_9002);
or U13054 (N_13054,N_10277,N_10532);
xnor U13055 (N_13055,N_9875,N_10218);
nand U13056 (N_13056,N_10326,N_9152);
and U13057 (N_13057,N_9370,N_11771);
or U13058 (N_13058,N_11325,N_11901);
nor U13059 (N_13059,N_11339,N_10203);
nor U13060 (N_13060,N_10656,N_10528);
xnor U13061 (N_13061,N_11286,N_11561);
nor U13062 (N_13062,N_9702,N_11586);
and U13063 (N_13063,N_9142,N_9432);
xor U13064 (N_13064,N_11272,N_10468);
or U13065 (N_13065,N_10274,N_11397);
and U13066 (N_13066,N_11926,N_9856);
xnor U13067 (N_13067,N_10023,N_10634);
nor U13068 (N_13068,N_11995,N_9836);
or U13069 (N_13069,N_10412,N_10522);
or U13070 (N_13070,N_9375,N_9033);
and U13071 (N_13071,N_9552,N_11063);
nand U13072 (N_13072,N_10017,N_9611);
nor U13073 (N_13073,N_9257,N_10823);
nor U13074 (N_13074,N_11116,N_11775);
xor U13075 (N_13075,N_11118,N_11688);
xnor U13076 (N_13076,N_10462,N_10470);
nand U13077 (N_13077,N_10436,N_11713);
or U13078 (N_13078,N_10624,N_10322);
and U13079 (N_13079,N_10942,N_11507);
nand U13080 (N_13080,N_9378,N_10376);
xnor U13081 (N_13081,N_11853,N_11858);
and U13082 (N_13082,N_10675,N_11819);
nand U13083 (N_13083,N_11413,N_9140);
nor U13084 (N_13084,N_11132,N_10251);
or U13085 (N_13085,N_11327,N_9801);
xnor U13086 (N_13086,N_9179,N_10135);
and U13087 (N_13087,N_11493,N_11962);
xor U13088 (N_13088,N_10901,N_9212);
and U13089 (N_13089,N_10929,N_11862);
and U13090 (N_13090,N_11736,N_10355);
nor U13091 (N_13091,N_10450,N_9888);
and U13092 (N_13092,N_9253,N_9296);
nor U13093 (N_13093,N_9631,N_11835);
xor U13094 (N_13094,N_10834,N_11608);
nor U13095 (N_13095,N_9489,N_9010);
or U13096 (N_13096,N_10902,N_11867);
and U13097 (N_13097,N_11437,N_9503);
nor U13098 (N_13098,N_9480,N_10632);
nor U13099 (N_13099,N_9886,N_9807);
or U13100 (N_13100,N_9698,N_11212);
xnor U13101 (N_13101,N_10068,N_10602);
xor U13102 (N_13102,N_9056,N_11071);
nor U13103 (N_13103,N_11545,N_11001);
nand U13104 (N_13104,N_10327,N_9786);
xnor U13105 (N_13105,N_10414,N_10166);
or U13106 (N_13106,N_10404,N_11065);
xor U13107 (N_13107,N_9082,N_9519);
and U13108 (N_13108,N_10557,N_9838);
or U13109 (N_13109,N_11468,N_10128);
nand U13110 (N_13110,N_10030,N_9443);
or U13111 (N_13111,N_11643,N_11455);
nor U13112 (N_13112,N_9192,N_10083);
nand U13113 (N_13113,N_9214,N_10144);
nand U13114 (N_13114,N_10178,N_11218);
nand U13115 (N_13115,N_9968,N_9051);
or U13116 (N_13116,N_10060,N_9408);
nand U13117 (N_13117,N_11117,N_11861);
xor U13118 (N_13118,N_10106,N_11615);
and U13119 (N_13119,N_9852,N_9278);
nor U13120 (N_13120,N_9897,N_9903);
or U13121 (N_13121,N_11363,N_10572);
and U13122 (N_13122,N_9300,N_9653);
nand U13123 (N_13123,N_11230,N_10818);
xor U13124 (N_13124,N_9453,N_10499);
or U13125 (N_13125,N_9325,N_11144);
nor U13126 (N_13126,N_10258,N_10896);
nor U13127 (N_13127,N_10695,N_9568);
nor U13128 (N_13128,N_9810,N_9585);
xor U13129 (N_13129,N_11786,N_11248);
and U13130 (N_13130,N_11193,N_9814);
and U13131 (N_13131,N_11590,N_10869);
and U13132 (N_13132,N_10152,N_11910);
or U13133 (N_13133,N_11345,N_9343);
and U13134 (N_13134,N_10689,N_10481);
nand U13135 (N_13135,N_11965,N_9467);
nor U13136 (N_13136,N_9812,N_11922);
or U13137 (N_13137,N_9578,N_9263);
nor U13138 (N_13138,N_11091,N_11426);
xnor U13139 (N_13139,N_9943,N_9038);
nor U13140 (N_13140,N_10867,N_10225);
nand U13141 (N_13141,N_9992,N_11764);
and U13142 (N_13142,N_10053,N_11610);
xnor U13143 (N_13143,N_10771,N_11667);
nor U13144 (N_13144,N_9457,N_9608);
nand U13145 (N_13145,N_10994,N_9087);
and U13146 (N_13146,N_10254,N_10892);
nor U13147 (N_13147,N_11574,N_9217);
nor U13148 (N_13148,N_10253,N_11750);
and U13149 (N_13149,N_10265,N_9882);
or U13150 (N_13150,N_10828,N_10489);
and U13151 (N_13151,N_9625,N_9311);
nand U13152 (N_13152,N_10194,N_9763);
and U13153 (N_13153,N_10958,N_10826);
nor U13154 (N_13154,N_9449,N_9751);
and U13155 (N_13155,N_9396,N_11312);
and U13156 (N_13156,N_9342,N_10415);
or U13157 (N_13157,N_10906,N_11326);
or U13158 (N_13158,N_10776,N_11933);
or U13159 (N_13159,N_11398,N_9701);
and U13160 (N_13160,N_9242,N_10387);
xnor U13161 (N_13161,N_9209,N_9258);
or U13162 (N_13162,N_9842,N_9279);
or U13163 (N_13163,N_11146,N_11115);
and U13164 (N_13164,N_11986,N_10337);
nand U13165 (N_13165,N_10866,N_11245);
nand U13166 (N_13166,N_9309,N_11278);
nor U13167 (N_13167,N_11103,N_9448);
xnor U13168 (N_13168,N_10900,N_9023);
nand U13169 (N_13169,N_10046,N_11638);
nor U13170 (N_13170,N_11251,N_10946);
or U13171 (N_13171,N_9121,N_10882);
nand U13172 (N_13172,N_11036,N_11407);
nand U13173 (N_13173,N_10853,N_9206);
nand U13174 (N_13174,N_9825,N_10275);
or U13175 (N_13175,N_10506,N_9284);
nand U13176 (N_13176,N_10821,N_11300);
nor U13177 (N_13177,N_11328,N_10124);
nor U13178 (N_13178,N_10397,N_11698);
and U13179 (N_13179,N_9332,N_9678);
nor U13180 (N_13180,N_11130,N_9030);
nor U13181 (N_13181,N_9233,N_11787);
nand U13182 (N_13182,N_10286,N_11308);
nand U13183 (N_13183,N_9752,N_11728);
and U13184 (N_13184,N_9956,N_9269);
or U13185 (N_13185,N_11376,N_11302);
nand U13186 (N_13186,N_10758,N_9676);
or U13187 (N_13187,N_11905,N_11789);
and U13188 (N_13188,N_9511,N_11509);
nand U13189 (N_13189,N_9394,N_11805);
xor U13190 (N_13190,N_9832,N_11262);
and U13191 (N_13191,N_11640,N_9014);
and U13192 (N_13192,N_11528,N_9095);
nor U13193 (N_13193,N_9604,N_11791);
xor U13194 (N_13194,N_10045,N_11871);
nor U13195 (N_13195,N_11120,N_11692);
nand U13196 (N_13196,N_10825,N_10564);
and U13197 (N_13197,N_10642,N_9423);
nand U13198 (N_13198,N_10874,N_11592);
nor U13199 (N_13199,N_10699,N_11612);
and U13200 (N_13200,N_9493,N_10006);
nor U13201 (N_13201,N_10329,N_11171);
or U13202 (N_13202,N_9254,N_9487);
nor U13203 (N_13203,N_10456,N_9240);
or U13204 (N_13204,N_11891,N_9156);
nor U13205 (N_13205,N_9880,N_10593);
xnor U13206 (N_13206,N_11735,N_9691);
or U13207 (N_13207,N_10597,N_11277);
or U13208 (N_13208,N_10767,N_11165);
nand U13209 (N_13209,N_10350,N_10237);
nand U13210 (N_13210,N_10769,N_10338);
nand U13211 (N_13211,N_9105,N_10016);
nor U13212 (N_13212,N_10526,N_9364);
and U13213 (N_13213,N_9662,N_9098);
or U13214 (N_13214,N_11322,N_9864);
and U13215 (N_13215,N_11911,N_9865);
or U13216 (N_13216,N_11188,N_9978);
or U13217 (N_13217,N_11585,N_11675);
or U13218 (N_13218,N_9697,N_11762);
xor U13219 (N_13219,N_11209,N_9995);
nand U13220 (N_13220,N_11304,N_11967);
xor U13221 (N_13221,N_11284,N_10280);
nand U13222 (N_13222,N_9175,N_9397);
or U13223 (N_13223,N_9921,N_11187);
xor U13224 (N_13224,N_10366,N_11904);
nand U13225 (N_13225,N_10431,N_9845);
or U13226 (N_13226,N_9871,N_11282);
and U13227 (N_13227,N_11056,N_9032);
nor U13228 (N_13228,N_9811,N_9737);
and U13229 (N_13229,N_11864,N_10351);
nand U13230 (N_13230,N_10748,N_11752);
or U13231 (N_13231,N_11138,N_10070);
nor U13232 (N_13232,N_11616,N_11256);
nand U13233 (N_13233,N_9072,N_10555);
nor U13234 (N_13234,N_9220,N_9299);
nor U13235 (N_13235,N_10014,N_10015);
xnor U13236 (N_13236,N_10497,N_9791);
nor U13237 (N_13237,N_10005,N_9128);
xor U13238 (N_13238,N_10722,N_11102);
or U13239 (N_13239,N_9971,N_11879);
xor U13240 (N_13240,N_11015,N_11060);
nand U13241 (N_13241,N_10515,N_11657);
nor U13242 (N_13242,N_10377,N_10096);
nor U13243 (N_13243,N_11717,N_11823);
and U13244 (N_13244,N_10255,N_9137);
or U13245 (N_13245,N_10079,N_11636);
nor U13246 (N_13246,N_9256,N_10263);
or U13247 (N_13247,N_11672,N_9895);
nor U13248 (N_13248,N_11753,N_9237);
nand U13249 (N_13249,N_10680,N_11350);
and U13250 (N_13250,N_11745,N_10157);
xor U13251 (N_13251,N_9109,N_9367);
and U13252 (N_13252,N_9705,N_9846);
nor U13253 (N_13253,N_9383,N_10932);
xor U13254 (N_13254,N_9718,N_9393);
or U13255 (N_13255,N_10367,N_10328);
or U13256 (N_13256,N_11126,N_9627);
xnor U13257 (N_13257,N_10268,N_11473);
or U13258 (N_13258,N_10126,N_9835);
or U13259 (N_13259,N_11976,N_10705);
or U13260 (N_13260,N_9925,N_11980);
nand U13261 (N_13261,N_11358,N_10428);
or U13262 (N_13262,N_9549,N_9989);
or U13263 (N_13263,N_9430,N_10021);
nand U13264 (N_13264,N_11481,N_9929);
xor U13265 (N_13265,N_9372,N_10042);
nor U13266 (N_13266,N_11196,N_11323);
nor U13267 (N_13267,N_11099,N_11729);
nand U13268 (N_13268,N_10142,N_11558);
nand U13269 (N_13269,N_10227,N_10267);
and U13270 (N_13270,N_10075,N_9265);
or U13271 (N_13271,N_10931,N_9404);
and U13272 (N_13272,N_9735,N_10764);
xnor U13273 (N_13273,N_10188,N_10011);
xnor U13274 (N_13274,N_11844,N_10272);
or U13275 (N_13275,N_9229,N_11628);
or U13276 (N_13276,N_11179,N_10903);
xor U13277 (N_13277,N_9294,N_9794);
nand U13278 (N_13278,N_10765,N_10941);
nand U13279 (N_13279,N_9092,N_9020);
xor U13280 (N_13280,N_10529,N_11470);
nor U13281 (N_13281,N_10235,N_10201);
or U13282 (N_13282,N_10750,N_9419);
xnor U13283 (N_13283,N_9139,N_11923);
nand U13284 (N_13284,N_11572,N_9908);
nor U13285 (N_13285,N_11810,N_10186);
nor U13286 (N_13286,N_10865,N_11444);
nor U13287 (N_13287,N_11169,N_10390);
xnor U13288 (N_13288,N_10435,N_11204);
nor U13289 (N_13289,N_11953,N_9199);
nor U13290 (N_13290,N_9046,N_9535);
or U13291 (N_13291,N_11046,N_9193);
nand U13292 (N_13292,N_11435,N_9969);
nor U13293 (N_13293,N_10779,N_9855);
nor U13294 (N_13294,N_10341,N_9301);
and U13295 (N_13295,N_10304,N_11836);
xnor U13296 (N_13296,N_11359,N_10531);
xor U13297 (N_13297,N_9753,N_10334);
nor U13298 (N_13298,N_10723,N_10226);
nand U13299 (N_13299,N_11379,N_10394);
nor U13300 (N_13300,N_9859,N_11833);
nand U13301 (N_13301,N_9600,N_10335);
xor U13302 (N_13302,N_10148,N_9642);
nand U13303 (N_13303,N_9843,N_9537);
nand U13304 (N_13304,N_11760,N_9962);
nand U13305 (N_13305,N_11971,N_9004);
and U13306 (N_13306,N_9016,N_9760);
and U13307 (N_13307,N_10065,N_9345);
and U13308 (N_13308,N_10067,N_10937);
nor U13309 (N_13309,N_11539,N_9191);
and U13310 (N_13310,N_10180,N_10854);
xor U13311 (N_13311,N_11580,N_11605);
xor U13312 (N_13312,N_11946,N_10216);
and U13313 (N_13313,N_9407,N_9295);
nand U13314 (N_13314,N_11689,N_11639);
nor U13315 (N_13315,N_11642,N_11189);
nor U13316 (N_13316,N_9866,N_11773);
nand U13317 (N_13317,N_11180,N_10305);
nor U13318 (N_13318,N_10449,N_9412);
or U13319 (N_13319,N_9848,N_10979);
xor U13320 (N_13320,N_11567,N_11200);
nor U13321 (N_13321,N_10405,N_10922);
or U13322 (N_13322,N_9308,N_9114);
xor U13323 (N_13323,N_9686,N_11579);
nand U13324 (N_13324,N_9546,N_11491);
or U13325 (N_13325,N_9539,N_10443);
and U13326 (N_13326,N_10737,N_9782);
nor U13327 (N_13327,N_10291,N_10187);
xor U13328 (N_13328,N_11124,N_10208);
xnor U13329 (N_13329,N_9475,N_11022);
and U13330 (N_13330,N_11239,N_10276);
or U13331 (N_13331,N_10429,N_9470);
nor U13332 (N_13332,N_10048,N_10715);
xor U13333 (N_13333,N_10972,N_11112);
or U13334 (N_13334,N_10725,N_10623);
and U13335 (N_13335,N_9042,N_9044);
nor U13336 (N_13336,N_9602,N_11596);
and U13337 (N_13337,N_10442,N_11368);
xor U13338 (N_13338,N_10370,N_11244);
nand U13339 (N_13339,N_11075,N_11076);
xor U13340 (N_13340,N_10372,N_9293);
xor U13341 (N_13341,N_10565,N_11365);
or U13342 (N_13342,N_11866,N_11924);
and U13343 (N_13343,N_11676,N_11674);
xnor U13344 (N_13344,N_10576,N_9601);
nor U13345 (N_13345,N_10464,N_10682);
and U13346 (N_13346,N_11162,N_10071);
nand U13347 (N_13347,N_9561,N_10611);
xnor U13348 (N_13348,N_9937,N_9788);
xor U13349 (N_13349,N_9996,N_10648);
xnor U13350 (N_13350,N_9955,N_11107);
and U13351 (N_13351,N_11683,N_10362);
nand U13352 (N_13352,N_11333,N_10172);
or U13353 (N_13353,N_9709,N_11037);
nand U13354 (N_13354,N_9169,N_10312);
xor U13355 (N_13355,N_10831,N_9306);
and U13356 (N_13356,N_9132,N_10219);
nor U13357 (N_13357,N_11295,N_9083);
nand U13358 (N_13358,N_11501,N_10454);
and U13359 (N_13359,N_10469,N_11442);
nor U13360 (N_13360,N_9065,N_10132);
and U13361 (N_13361,N_10934,N_10635);
or U13362 (N_13362,N_11814,N_10806);
or U13363 (N_13363,N_9610,N_10850);
nor U13364 (N_13364,N_11726,N_9182);
or U13365 (N_13365,N_11581,N_10081);
and U13366 (N_13366,N_10816,N_9902);
and U13367 (N_13367,N_10217,N_11424);
xnor U13368 (N_13368,N_9247,N_11741);
xor U13369 (N_13369,N_9078,N_9268);
and U13370 (N_13370,N_11828,N_10980);
or U13371 (N_13371,N_9255,N_10318);
nand U13372 (N_13372,N_10620,N_11347);
nor U13373 (N_13373,N_10720,N_9035);
nand U13374 (N_13374,N_9635,N_11884);
nand U13375 (N_13375,N_10356,N_10013);
or U13376 (N_13376,N_9572,N_10843);
nor U13377 (N_13377,N_9734,N_10177);
nand U13378 (N_13378,N_9967,N_10049);
nand U13379 (N_13379,N_10763,N_11931);
and U13380 (N_13380,N_11401,N_11092);
or U13381 (N_13381,N_9130,N_10740);
xnor U13382 (N_13382,N_10129,N_11114);
nor U13383 (N_13383,N_10839,N_9154);
and U13384 (N_13384,N_10169,N_9172);
nand U13385 (N_13385,N_11748,N_10795);
xor U13386 (N_13386,N_11430,N_11685);
nand U13387 (N_13387,N_11343,N_10308);
nand U13388 (N_13388,N_9916,N_11906);
nor U13389 (N_13389,N_10789,N_10330);
nand U13390 (N_13390,N_9161,N_9124);
xnor U13391 (N_13391,N_11298,N_10990);
xnor U13392 (N_13392,N_10558,N_9850);
or U13393 (N_13393,N_11827,N_9620);
nand U13394 (N_13394,N_9746,N_11508);
or U13395 (N_13395,N_10690,N_9320);
and U13396 (N_13396,N_11556,N_10716);
nor U13397 (N_13397,N_9017,N_9216);
nor U13398 (N_13398,N_10297,N_9958);
xnor U13399 (N_13399,N_9529,N_9079);
nor U13400 (N_13400,N_11937,N_11527);
or U13401 (N_13401,N_11167,N_11715);
nor U13402 (N_13402,N_11913,N_9935);
or U13403 (N_13403,N_10782,N_10728);
nor U13404 (N_13404,N_11951,N_10473);
nand U13405 (N_13405,N_11010,N_9417);
nor U13406 (N_13406,N_9141,N_11382);
nor U13407 (N_13407,N_10525,N_9420);
nand U13408 (N_13408,N_11040,N_11051);
nand U13409 (N_13409,N_11930,N_11575);
nand U13410 (N_13410,N_10463,N_10638);
nor U13411 (N_13411,N_9993,N_11217);
nand U13412 (N_13412,N_9341,N_10477);
xnor U13413 (N_13413,N_10192,N_10041);
nor U13414 (N_13414,N_11400,N_9281);
nor U13415 (N_13415,N_10762,N_9563);
nand U13416 (N_13416,N_10753,N_10812);
or U13417 (N_13417,N_9623,N_9551);
nor U13418 (N_13418,N_11490,N_10884);
xnor U13419 (N_13419,N_10025,N_11587);
and U13420 (N_13420,N_9648,N_9721);
or U13421 (N_13421,N_11691,N_9259);
xor U13422 (N_13422,N_11182,N_11997);
xnor U13423 (N_13423,N_11361,N_9739);
nor U13424 (N_13424,N_10240,N_10540);
xor U13425 (N_13425,N_11516,N_10182);
xor U13426 (N_13426,N_10965,N_10457);
xnor U13427 (N_13427,N_9657,N_10422);
nand U13428 (N_13428,N_11623,N_10804);
nand U13429 (N_13429,N_10125,N_9728);
nor U13430 (N_13430,N_9694,N_11069);
nor U13431 (N_13431,N_9053,N_10961);
nor U13432 (N_13432,N_9456,N_10613);
xor U13433 (N_13433,N_9502,N_10408);
or U13434 (N_13434,N_9985,N_10660);
or U13435 (N_13435,N_11054,N_9716);
or U13436 (N_13436,N_10054,N_10743);
and U13437 (N_13437,N_9228,N_9966);
xor U13438 (N_13438,N_11270,N_9225);
nand U13439 (N_13439,N_9262,N_11105);
or U13440 (N_13440,N_10991,N_11303);
nor U13441 (N_13441,N_10434,N_9690);
nand U13442 (N_13442,N_11709,N_10501);
xor U13443 (N_13443,N_10521,N_11049);
or U13444 (N_13444,N_10594,N_11157);
and U13445 (N_13445,N_11344,N_10008);
or U13446 (N_13446,N_11021,N_9736);
or U13447 (N_13447,N_9862,N_11984);
nand U13448 (N_13448,N_10662,N_11255);
xnor U13449 (N_13449,N_10174,N_11489);
xor U13450 (N_13450,N_9054,N_11878);
or U13451 (N_13451,N_9732,N_9951);
xor U13452 (N_13452,N_11705,N_11938);
nor U13453 (N_13453,N_10491,N_11846);
and U13454 (N_13454,N_10983,N_11977);
and U13455 (N_13455,N_9494,N_11757);
and U13456 (N_13456,N_11549,N_9729);
and U13457 (N_13457,N_11815,N_10671);
nor U13458 (N_13458,N_11634,N_11231);
or U13459 (N_13459,N_9040,N_9022);
or U13460 (N_13460,N_11242,N_9938);
or U13461 (N_13461,N_11459,N_9211);
xnor U13462 (N_13462,N_9018,N_10393);
nand U13463 (N_13463,N_9190,N_9963);
nor U13464 (N_13464,N_11770,N_11772);
xnor U13465 (N_13465,N_11611,N_11724);
or U13466 (N_13466,N_9747,N_9820);
nor U13467 (N_13467,N_10924,N_10478);
or U13468 (N_13468,N_10578,N_9445);
nor U13469 (N_13469,N_9116,N_9879);
nand U13470 (N_13470,N_11052,N_11614);
nor U13471 (N_13471,N_11025,N_9504);
nor U13472 (N_13472,N_9982,N_9471);
nor U13473 (N_13473,N_9924,N_11807);
nand U13474 (N_13474,N_11428,N_10625);
or U13475 (N_13475,N_10104,N_10630);
and U13476 (N_13476,N_9155,N_11161);
or U13477 (N_13477,N_9693,N_10530);
xnor U13478 (N_13478,N_9144,N_10064);
nor U13479 (N_13479,N_10574,N_9688);
nand U13480 (N_13480,N_9084,N_10153);
or U13481 (N_13481,N_11417,N_10051);
or U13482 (N_13482,N_10618,N_9597);
or U13483 (N_13483,N_11934,N_11127);
or U13484 (N_13484,N_9949,N_10600);
and U13485 (N_13485,N_9528,N_11305);
xor U13486 (N_13486,N_11199,N_9481);
xor U13487 (N_13487,N_9724,N_11648);
xor U13488 (N_13488,N_10657,N_11996);
or U13489 (N_13489,N_11548,N_9075);
and U13490 (N_13490,N_9704,N_10476);
or U13491 (N_13491,N_9707,N_9203);
nand U13492 (N_13492,N_11393,N_9333);
or U13493 (N_13493,N_9275,N_9472);
and U13494 (N_13494,N_10342,N_10655);
or U13495 (N_13495,N_11920,N_11855);
and U13496 (N_13496,N_10168,N_9710);
and U13497 (N_13497,N_11550,N_10061);
nor U13498 (N_13498,N_9180,N_11463);
and U13499 (N_13499,N_9524,N_11552);
or U13500 (N_13500,N_9210,N_9722);
and U13501 (N_13501,N_10364,N_11179);
xnor U13502 (N_13502,N_9356,N_9993);
or U13503 (N_13503,N_9801,N_9013);
xnor U13504 (N_13504,N_9134,N_10932);
nand U13505 (N_13505,N_9084,N_10059);
or U13506 (N_13506,N_9749,N_11903);
xor U13507 (N_13507,N_9449,N_9771);
and U13508 (N_13508,N_11721,N_11267);
nor U13509 (N_13509,N_11091,N_9074);
or U13510 (N_13510,N_9189,N_11766);
nor U13511 (N_13511,N_11954,N_11183);
and U13512 (N_13512,N_10360,N_11784);
nand U13513 (N_13513,N_10986,N_9441);
xnor U13514 (N_13514,N_11358,N_9328);
xnor U13515 (N_13515,N_9917,N_9935);
or U13516 (N_13516,N_11245,N_11456);
nand U13517 (N_13517,N_9051,N_11626);
nor U13518 (N_13518,N_10894,N_9516);
and U13519 (N_13519,N_11619,N_11198);
and U13520 (N_13520,N_9775,N_9658);
xnor U13521 (N_13521,N_9942,N_9633);
nand U13522 (N_13522,N_11938,N_9275);
or U13523 (N_13523,N_11261,N_11184);
and U13524 (N_13524,N_11769,N_10961);
xor U13525 (N_13525,N_10486,N_11524);
nand U13526 (N_13526,N_9932,N_9455);
and U13527 (N_13527,N_11293,N_10532);
nand U13528 (N_13528,N_9318,N_10757);
nor U13529 (N_13529,N_9706,N_9027);
nor U13530 (N_13530,N_11122,N_10511);
or U13531 (N_13531,N_9325,N_9177);
nor U13532 (N_13532,N_9431,N_9299);
nor U13533 (N_13533,N_9482,N_9352);
xnor U13534 (N_13534,N_11299,N_10303);
and U13535 (N_13535,N_10988,N_9730);
and U13536 (N_13536,N_9187,N_10441);
or U13537 (N_13537,N_10874,N_11508);
nand U13538 (N_13538,N_10084,N_11360);
nor U13539 (N_13539,N_9142,N_10590);
xnor U13540 (N_13540,N_10918,N_10234);
nand U13541 (N_13541,N_11940,N_10622);
or U13542 (N_13542,N_11480,N_11976);
nand U13543 (N_13543,N_9070,N_9742);
nor U13544 (N_13544,N_11256,N_10706);
and U13545 (N_13545,N_10831,N_10669);
or U13546 (N_13546,N_11069,N_11149);
and U13547 (N_13547,N_9239,N_9242);
or U13548 (N_13548,N_9924,N_10935);
nor U13549 (N_13549,N_10599,N_11246);
and U13550 (N_13550,N_10772,N_11221);
nor U13551 (N_13551,N_10125,N_9001);
and U13552 (N_13552,N_10735,N_9018);
xnor U13553 (N_13553,N_11521,N_11177);
nor U13554 (N_13554,N_9676,N_10861);
and U13555 (N_13555,N_11022,N_11747);
nor U13556 (N_13556,N_11738,N_9086);
nand U13557 (N_13557,N_11116,N_11008);
xnor U13558 (N_13558,N_11689,N_11110);
and U13559 (N_13559,N_10413,N_11197);
or U13560 (N_13560,N_11981,N_11598);
or U13561 (N_13561,N_10245,N_11129);
nor U13562 (N_13562,N_10739,N_10965);
and U13563 (N_13563,N_10759,N_9887);
and U13564 (N_13564,N_11415,N_10497);
xnor U13565 (N_13565,N_10615,N_9390);
nor U13566 (N_13566,N_9126,N_10283);
nor U13567 (N_13567,N_11673,N_10512);
xnor U13568 (N_13568,N_9673,N_11395);
or U13569 (N_13569,N_10905,N_9723);
or U13570 (N_13570,N_11900,N_11043);
xnor U13571 (N_13571,N_10268,N_9367);
nand U13572 (N_13572,N_11313,N_9136);
nand U13573 (N_13573,N_10738,N_11840);
xnor U13574 (N_13574,N_9163,N_9425);
xor U13575 (N_13575,N_9442,N_10773);
xor U13576 (N_13576,N_9052,N_11495);
nor U13577 (N_13577,N_9511,N_10835);
and U13578 (N_13578,N_11921,N_9250);
and U13579 (N_13579,N_9703,N_11806);
nand U13580 (N_13580,N_9033,N_10110);
xnor U13581 (N_13581,N_10794,N_10520);
nand U13582 (N_13582,N_10140,N_11899);
and U13583 (N_13583,N_10062,N_9722);
or U13584 (N_13584,N_11950,N_11753);
xor U13585 (N_13585,N_10992,N_11116);
nor U13586 (N_13586,N_10390,N_11995);
xnor U13587 (N_13587,N_10780,N_11057);
or U13588 (N_13588,N_9623,N_10174);
xnor U13589 (N_13589,N_9097,N_11707);
and U13590 (N_13590,N_9789,N_11831);
nand U13591 (N_13591,N_11084,N_9613);
nor U13592 (N_13592,N_11237,N_10967);
and U13593 (N_13593,N_9448,N_9038);
and U13594 (N_13594,N_9663,N_10168);
or U13595 (N_13595,N_11449,N_11718);
nor U13596 (N_13596,N_10014,N_10904);
and U13597 (N_13597,N_11160,N_10909);
nand U13598 (N_13598,N_11281,N_10789);
nor U13599 (N_13599,N_10401,N_10114);
or U13600 (N_13600,N_10606,N_11277);
nor U13601 (N_13601,N_10277,N_10372);
and U13602 (N_13602,N_9084,N_10615);
or U13603 (N_13603,N_11745,N_11468);
nand U13604 (N_13604,N_11160,N_11337);
nand U13605 (N_13605,N_10111,N_11531);
or U13606 (N_13606,N_10657,N_11699);
and U13607 (N_13607,N_10651,N_9014);
nor U13608 (N_13608,N_9074,N_11110);
and U13609 (N_13609,N_9133,N_10223);
nand U13610 (N_13610,N_11332,N_10198);
nor U13611 (N_13611,N_9700,N_9211);
or U13612 (N_13612,N_10598,N_10340);
and U13613 (N_13613,N_11733,N_10548);
nand U13614 (N_13614,N_10255,N_10373);
nand U13615 (N_13615,N_11797,N_10070);
or U13616 (N_13616,N_11059,N_9761);
or U13617 (N_13617,N_11990,N_10908);
and U13618 (N_13618,N_10485,N_9006);
xnor U13619 (N_13619,N_10539,N_11414);
xnor U13620 (N_13620,N_9110,N_11726);
and U13621 (N_13621,N_11354,N_10670);
or U13622 (N_13622,N_11758,N_11247);
nand U13623 (N_13623,N_10310,N_9787);
nor U13624 (N_13624,N_9768,N_11609);
xnor U13625 (N_13625,N_10013,N_9943);
and U13626 (N_13626,N_9475,N_10030);
or U13627 (N_13627,N_11548,N_11112);
or U13628 (N_13628,N_9354,N_9461);
and U13629 (N_13629,N_9422,N_11589);
and U13630 (N_13630,N_10520,N_9497);
and U13631 (N_13631,N_10299,N_9807);
and U13632 (N_13632,N_10157,N_10933);
nor U13633 (N_13633,N_9979,N_11194);
and U13634 (N_13634,N_9029,N_9106);
and U13635 (N_13635,N_11345,N_11084);
and U13636 (N_13636,N_9137,N_9689);
nor U13637 (N_13637,N_10888,N_11219);
and U13638 (N_13638,N_11986,N_10239);
and U13639 (N_13639,N_10948,N_11629);
or U13640 (N_13640,N_11627,N_10344);
and U13641 (N_13641,N_11765,N_10232);
nand U13642 (N_13642,N_10359,N_9766);
and U13643 (N_13643,N_9790,N_10882);
xor U13644 (N_13644,N_11519,N_10805);
nand U13645 (N_13645,N_11781,N_11619);
or U13646 (N_13646,N_9389,N_11381);
xnor U13647 (N_13647,N_10786,N_10221);
nor U13648 (N_13648,N_10617,N_9939);
or U13649 (N_13649,N_10737,N_9066);
and U13650 (N_13650,N_10558,N_11055);
nand U13651 (N_13651,N_11638,N_9774);
or U13652 (N_13652,N_10488,N_9451);
and U13653 (N_13653,N_9911,N_9371);
nand U13654 (N_13654,N_11701,N_9470);
xor U13655 (N_13655,N_9678,N_11051);
nand U13656 (N_13656,N_10279,N_11911);
nor U13657 (N_13657,N_10778,N_9243);
nand U13658 (N_13658,N_10476,N_11958);
xnor U13659 (N_13659,N_10421,N_11690);
xor U13660 (N_13660,N_11802,N_11820);
or U13661 (N_13661,N_11339,N_10513);
nor U13662 (N_13662,N_11085,N_11114);
or U13663 (N_13663,N_11786,N_9614);
or U13664 (N_13664,N_10510,N_9815);
xor U13665 (N_13665,N_10108,N_9433);
nand U13666 (N_13666,N_10014,N_10527);
and U13667 (N_13667,N_11141,N_10528);
and U13668 (N_13668,N_10913,N_10364);
xor U13669 (N_13669,N_9032,N_10106);
or U13670 (N_13670,N_9613,N_9845);
xor U13671 (N_13671,N_11484,N_10576);
or U13672 (N_13672,N_10397,N_10391);
xor U13673 (N_13673,N_11542,N_9387);
nor U13674 (N_13674,N_11009,N_11476);
nand U13675 (N_13675,N_11771,N_9364);
and U13676 (N_13676,N_9836,N_11846);
nand U13677 (N_13677,N_9038,N_9062);
nand U13678 (N_13678,N_9315,N_9570);
xnor U13679 (N_13679,N_10048,N_11030);
xor U13680 (N_13680,N_11068,N_10592);
nand U13681 (N_13681,N_11754,N_9229);
or U13682 (N_13682,N_9657,N_10479);
nor U13683 (N_13683,N_9427,N_9144);
or U13684 (N_13684,N_10622,N_10232);
or U13685 (N_13685,N_9187,N_9533);
nor U13686 (N_13686,N_9638,N_9332);
or U13687 (N_13687,N_10253,N_11634);
nor U13688 (N_13688,N_9816,N_10903);
or U13689 (N_13689,N_10060,N_11155);
or U13690 (N_13690,N_9231,N_10619);
nand U13691 (N_13691,N_9425,N_10193);
nor U13692 (N_13692,N_10488,N_10632);
and U13693 (N_13693,N_9557,N_11056);
nor U13694 (N_13694,N_11014,N_11972);
xor U13695 (N_13695,N_10191,N_9870);
or U13696 (N_13696,N_9097,N_11449);
nor U13697 (N_13697,N_10122,N_9647);
xor U13698 (N_13698,N_9813,N_10972);
or U13699 (N_13699,N_9007,N_9867);
xnor U13700 (N_13700,N_11336,N_11856);
nand U13701 (N_13701,N_10131,N_11919);
and U13702 (N_13702,N_9939,N_10786);
nand U13703 (N_13703,N_10467,N_9672);
or U13704 (N_13704,N_9498,N_9252);
nand U13705 (N_13705,N_11233,N_9695);
nor U13706 (N_13706,N_9791,N_9687);
xor U13707 (N_13707,N_11856,N_10418);
nand U13708 (N_13708,N_11030,N_11425);
and U13709 (N_13709,N_10029,N_9836);
nand U13710 (N_13710,N_10368,N_10584);
and U13711 (N_13711,N_11670,N_10665);
and U13712 (N_13712,N_11063,N_9611);
xnor U13713 (N_13713,N_9126,N_9705);
or U13714 (N_13714,N_9263,N_9722);
or U13715 (N_13715,N_11548,N_11225);
and U13716 (N_13716,N_10924,N_9387);
nand U13717 (N_13717,N_9888,N_10242);
and U13718 (N_13718,N_11684,N_11902);
xnor U13719 (N_13719,N_9005,N_9724);
xor U13720 (N_13720,N_11823,N_10523);
nand U13721 (N_13721,N_9563,N_11871);
nor U13722 (N_13722,N_9924,N_9181);
nand U13723 (N_13723,N_11742,N_10805);
and U13724 (N_13724,N_10602,N_9302);
or U13725 (N_13725,N_9421,N_11451);
xor U13726 (N_13726,N_10952,N_10777);
or U13727 (N_13727,N_11554,N_10820);
or U13728 (N_13728,N_11862,N_10282);
or U13729 (N_13729,N_10091,N_11761);
nand U13730 (N_13730,N_11217,N_10355);
nor U13731 (N_13731,N_10068,N_11547);
nor U13732 (N_13732,N_10825,N_9276);
and U13733 (N_13733,N_10352,N_11981);
nor U13734 (N_13734,N_10821,N_9333);
and U13735 (N_13735,N_10929,N_10996);
or U13736 (N_13736,N_11652,N_9244);
xor U13737 (N_13737,N_10914,N_11215);
xnor U13738 (N_13738,N_9853,N_10859);
nor U13739 (N_13739,N_10620,N_10757);
or U13740 (N_13740,N_11875,N_9939);
nor U13741 (N_13741,N_11901,N_10635);
xor U13742 (N_13742,N_10915,N_9485);
nor U13743 (N_13743,N_11200,N_10973);
nand U13744 (N_13744,N_9141,N_9437);
nor U13745 (N_13745,N_9753,N_9091);
nand U13746 (N_13746,N_10126,N_9978);
nor U13747 (N_13747,N_11221,N_10401);
nor U13748 (N_13748,N_10272,N_9302);
xnor U13749 (N_13749,N_11280,N_11291);
nand U13750 (N_13750,N_9999,N_11002);
or U13751 (N_13751,N_9299,N_11344);
nand U13752 (N_13752,N_9521,N_9999);
xnor U13753 (N_13753,N_11951,N_11897);
nor U13754 (N_13754,N_11418,N_11572);
or U13755 (N_13755,N_11213,N_9053);
or U13756 (N_13756,N_10769,N_11274);
xor U13757 (N_13757,N_9582,N_10567);
nor U13758 (N_13758,N_9654,N_10376);
nand U13759 (N_13759,N_11219,N_11723);
and U13760 (N_13760,N_10902,N_9542);
nor U13761 (N_13761,N_9401,N_10244);
xnor U13762 (N_13762,N_9041,N_11161);
and U13763 (N_13763,N_11465,N_9245);
xnor U13764 (N_13764,N_11697,N_10504);
nor U13765 (N_13765,N_10243,N_10617);
and U13766 (N_13766,N_11611,N_10117);
or U13767 (N_13767,N_10563,N_10631);
nor U13768 (N_13768,N_9770,N_9147);
xor U13769 (N_13769,N_11327,N_10348);
nor U13770 (N_13770,N_9687,N_11793);
and U13771 (N_13771,N_10072,N_11242);
nand U13772 (N_13772,N_11540,N_11234);
xor U13773 (N_13773,N_11933,N_11007);
nand U13774 (N_13774,N_10463,N_10843);
xnor U13775 (N_13775,N_9294,N_10285);
nor U13776 (N_13776,N_11489,N_10092);
and U13777 (N_13777,N_11684,N_10680);
nand U13778 (N_13778,N_11248,N_10167);
and U13779 (N_13779,N_11946,N_9718);
or U13780 (N_13780,N_10126,N_11112);
or U13781 (N_13781,N_9636,N_9127);
nor U13782 (N_13782,N_10237,N_10605);
and U13783 (N_13783,N_9939,N_11970);
xnor U13784 (N_13784,N_11153,N_9243);
or U13785 (N_13785,N_11208,N_11274);
and U13786 (N_13786,N_11965,N_10329);
nor U13787 (N_13787,N_10467,N_9783);
nor U13788 (N_13788,N_9369,N_10840);
and U13789 (N_13789,N_10966,N_11524);
or U13790 (N_13790,N_11188,N_10181);
nor U13791 (N_13791,N_11339,N_11895);
and U13792 (N_13792,N_11596,N_11606);
nor U13793 (N_13793,N_11610,N_10705);
and U13794 (N_13794,N_9133,N_11445);
nor U13795 (N_13795,N_10112,N_9539);
and U13796 (N_13796,N_11908,N_11395);
and U13797 (N_13797,N_9000,N_10757);
or U13798 (N_13798,N_9190,N_10646);
nor U13799 (N_13799,N_9057,N_10506);
xnor U13800 (N_13800,N_9804,N_9599);
and U13801 (N_13801,N_9945,N_9742);
and U13802 (N_13802,N_11584,N_9505);
xor U13803 (N_13803,N_10595,N_10966);
nor U13804 (N_13804,N_9634,N_9521);
nand U13805 (N_13805,N_10181,N_9377);
nand U13806 (N_13806,N_11972,N_9897);
xor U13807 (N_13807,N_11792,N_10011);
nand U13808 (N_13808,N_11063,N_11316);
xor U13809 (N_13809,N_11108,N_10349);
nand U13810 (N_13810,N_11814,N_9005);
nand U13811 (N_13811,N_9411,N_11301);
and U13812 (N_13812,N_11825,N_10462);
xor U13813 (N_13813,N_10298,N_11559);
xor U13814 (N_13814,N_10612,N_10352);
xor U13815 (N_13815,N_9685,N_9811);
nor U13816 (N_13816,N_9145,N_11437);
xnor U13817 (N_13817,N_10889,N_11248);
or U13818 (N_13818,N_11729,N_9773);
nand U13819 (N_13819,N_10041,N_9515);
nand U13820 (N_13820,N_9770,N_9984);
and U13821 (N_13821,N_9575,N_11516);
nor U13822 (N_13822,N_9343,N_11874);
or U13823 (N_13823,N_11000,N_11469);
nor U13824 (N_13824,N_9754,N_11424);
nand U13825 (N_13825,N_11311,N_9621);
or U13826 (N_13826,N_10100,N_10292);
and U13827 (N_13827,N_9577,N_11318);
or U13828 (N_13828,N_9855,N_11109);
nand U13829 (N_13829,N_9337,N_9016);
and U13830 (N_13830,N_11431,N_11454);
xor U13831 (N_13831,N_9231,N_11963);
xor U13832 (N_13832,N_9351,N_10406);
nor U13833 (N_13833,N_9056,N_9110);
or U13834 (N_13834,N_11003,N_11508);
nor U13835 (N_13835,N_10719,N_11679);
nor U13836 (N_13836,N_10053,N_10393);
nand U13837 (N_13837,N_9137,N_10646);
xor U13838 (N_13838,N_10395,N_11338);
nor U13839 (N_13839,N_10076,N_11647);
and U13840 (N_13840,N_9448,N_9699);
nor U13841 (N_13841,N_9937,N_9418);
or U13842 (N_13842,N_9121,N_10143);
nand U13843 (N_13843,N_11976,N_10013);
or U13844 (N_13844,N_10118,N_10012);
or U13845 (N_13845,N_11492,N_11709);
or U13846 (N_13846,N_10718,N_10824);
nand U13847 (N_13847,N_10310,N_9170);
nor U13848 (N_13848,N_10358,N_9029);
nor U13849 (N_13849,N_11764,N_10275);
or U13850 (N_13850,N_11556,N_9872);
nand U13851 (N_13851,N_10194,N_11995);
nand U13852 (N_13852,N_10081,N_10966);
xor U13853 (N_13853,N_11340,N_10050);
and U13854 (N_13854,N_9092,N_10249);
xnor U13855 (N_13855,N_11632,N_10723);
and U13856 (N_13856,N_10438,N_10443);
or U13857 (N_13857,N_11502,N_9257);
or U13858 (N_13858,N_9461,N_11022);
or U13859 (N_13859,N_11831,N_11659);
nand U13860 (N_13860,N_9999,N_10569);
and U13861 (N_13861,N_11690,N_9432);
xor U13862 (N_13862,N_10980,N_11406);
nor U13863 (N_13863,N_10267,N_10368);
or U13864 (N_13864,N_11099,N_11138);
xor U13865 (N_13865,N_10976,N_11125);
and U13866 (N_13866,N_11830,N_11828);
nor U13867 (N_13867,N_10388,N_10396);
xnor U13868 (N_13868,N_11660,N_9178);
and U13869 (N_13869,N_11013,N_9391);
and U13870 (N_13870,N_9630,N_10461);
xnor U13871 (N_13871,N_10043,N_10353);
or U13872 (N_13872,N_9398,N_11052);
nand U13873 (N_13873,N_11429,N_10344);
nor U13874 (N_13874,N_11143,N_9229);
nor U13875 (N_13875,N_9187,N_9263);
nand U13876 (N_13876,N_9784,N_11659);
or U13877 (N_13877,N_9042,N_11605);
nand U13878 (N_13878,N_11311,N_10704);
xor U13879 (N_13879,N_10072,N_10366);
xor U13880 (N_13880,N_10908,N_9719);
or U13881 (N_13881,N_10782,N_9429);
xor U13882 (N_13882,N_10831,N_11407);
nand U13883 (N_13883,N_10530,N_9842);
nor U13884 (N_13884,N_11479,N_11449);
xnor U13885 (N_13885,N_9481,N_9306);
xor U13886 (N_13886,N_10096,N_10119);
xnor U13887 (N_13887,N_10219,N_11523);
nand U13888 (N_13888,N_9587,N_11682);
and U13889 (N_13889,N_11899,N_9823);
and U13890 (N_13890,N_11062,N_10898);
xor U13891 (N_13891,N_9035,N_9726);
and U13892 (N_13892,N_9005,N_11266);
xnor U13893 (N_13893,N_10745,N_9431);
xor U13894 (N_13894,N_11657,N_11620);
or U13895 (N_13895,N_11785,N_11525);
or U13896 (N_13896,N_10507,N_10483);
xor U13897 (N_13897,N_9563,N_11039);
xor U13898 (N_13898,N_11893,N_11880);
and U13899 (N_13899,N_9657,N_11597);
nand U13900 (N_13900,N_10772,N_10599);
or U13901 (N_13901,N_11394,N_11313);
nand U13902 (N_13902,N_10373,N_9139);
xor U13903 (N_13903,N_10260,N_10987);
nor U13904 (N_13904,N_10995,N_9902);
nand U13905 (N_13905,N_11100,N_11720);
nand U13906 (N_13906,N_11413,N_11907);
or U13907 (N_13907,N_10194,N_9668);
and U13908 (N_13908,N_11588,N_11250);
nand U13909 (N_13909,N_10246,N_11669);
and U13910 (N_13910,N_11642,N_10457);
nor U13911 (N_13911,N_9742,N_11475);
or U13912 (N_13912,N_11106,N_11536);
xor U13913 (N_13913,N_9903,N_9786);
xor U13914 (N_13914,N_9423,N_9137);
xor U13915 (N_13915,N_10603,N_9368);
or U13916 (N_13916,N_11384,N_11751);
xnor U13917 (N_13917,N_10873,N_11308);
and U13918 (N_13918,N_9622,N_11533);
and U13919 (N_13919,N_9708,N_9187);
xnor U13920 (N_13920,N_11627,N_11381);
or U13921 (N_13921,N_9227,N_11428);
and U13922 (N_13922,N_11081,N_9321);
xor U13923 (N_13923,N_10177,N_10827);
nor U13924 (N_13924,N_9721,N_9314);
nand U13925 (N_13925,N_11146,N_10368);
and U13926 (N_13926,N_10083,N_9965);
nor U13927 (N_13927,N_10093,N_10984);
xor U13928 (N_13928,N_10231,N_9229);
or U13929 (N_13929,N_9213,N_11163);
nand U13930 (N_13930,N_11965,N_9497);
nor U13931 (N_13931,N_11754,N_9469);
and U13932 (N_13932,N_9216,N_9341);
and U13933 (N_13933,N_11633,N_9066);
xor U13934 (N_13934,N_10286,N_11000);
xnor U13935 (N_13935,N_11167,N_11834);
nor U13936 (N_13936,N_10173,N_10081);
nand U13937 (N_13937,N_11125,N_10405);
nand U13938 (N_13938,N_9532,N_10921);
xnor U13939 (N_13939,N_11589,N_9984);
xnor U13940 (N_13940,N_9460,N_11757);
xnor U13941 (N_13941,N_9616,N_10731);
xor U13942 (N_13942,N_10558,N_11205);
xnor U13943 (N_13943,N_10211,N_9419);
nor U13944 (N_13944,N_10073,N_9277);
nand U13945 (N_13945,N_11264,N_9534);
nand U13946 (N_13946,N_10033,N_10506);
xor U13947 (N_13947,N_11009,N_9550);
and U13948 (N_13948,N_9528,N_9800);
nor U13949 (N_13949,N_11670,N_9637);
nor U13950 (N_13950,N_10804,N_10056);
and U13951 (N_13951,N_9522,N_9857);
and U13952 (N_13952,N_9160,N_10088);
nand U13953 (N_13953,N_9090,N_9432);
xnor U13954 (N_13954,N_11446,N_9431);
and U13955 (N_13955,N_10571,N_11920);
and U13956 (N_13956,N_10438,N_9025);
and U13957 (N_13957,N_11085,N_9511);
and U13958 (N_13958,N_9015,N_10454);
and U13959 (N_13959,N_9842,N_9859);
or U13960 (N_13960,N_11273,N_10326);
nor U13961 (N_13961,N_9255,N_9374);
xor U13962 (N_13962,N_9517,N_10070);
xor U13963 (N_13963,N_11505,N_10685);
xor U13964 (N_13964,N_11145,N_10071);
nor U13965 (N_13965,N_10354,N_10028);
xor U13966 (N_13966,N_9098,N_11551);
nand U13967 (N_13967,N_10197,N_9923);
and U13968 (N_13968,N_11555,N_11970);
and U13969 (N_13969,N_11011,N_11141);
and U13970 (N_13970,N_10330,N_10400);
xor U13971 (N_13971,N_9823,N_9723);
xor U13972 (N_13972,N_10366,N_9671);
or U13973 (N_13973,N_11143,N_11072);
nand U13974 (N_13974,N_9165,N_10634);
nand U13975 (N_13975,N_11374,N_11884);
nor U13976 (N_13976,N_10487,N_11524);
or U13977 (N_13977,N_11464,N_10741);
nand U13978 (N_13978,N_10286,N_11511);
nor U13979 (N_13979,N_10978,N_11395);
nand U13980 (N_13980,N_10895,N_11653);
nor U13981 (N_13981,N_11362,N_11340);
nor U13982 (N_13982,N_11022,N_10150);
and U13983 (N_13983,N_11184,N_11061);
nand U13984 (N_13984,N_9313,N_10515);
nor U13985 (N_13985,N_9260,N_10677);
nand U13986 (N_13986,N_11428,N_10139);
nand U13987 (N_13987,N_11398,N_11678);
xnor U13988 (N_13988,N_11545,N_11794);
xnor U13989 (N_13989,N_10967,N_9271);
or U13990 (N_13990,N_10401,N_11983);
or U13991 (N_13991,N_11279,N_11210);
or U13992 (N_13992,N_10487,N_9737);
xnor U13993 (N_13993,N_10853,N_10077);
xnor U13994 (N_13994,N_10674,N_11513);
and U13995 (N_13995,N_10424,N_10757);
and U13996 (N_13996,N_10671,N_10315);
and U13997 (N_13997,N_10365,N_9652);
nand U13998 (N_13998,N_10129,N_11020);
nor U13999 (N_13999,N_10802,N_9567);
nand U14000 (N_14000,N_11721,N_11362);
nor U14001 (N_14001,N_11797,N_11038);
nor U14002 (N_14002,N_9928,N_11304);
and U14003 (N_14003,N_10455,N_11808);
nor U14004 (N_14004,N_11818,N_9380);
or U14005 (N_14005,N_11906,N_11745);
and U14006 (N_14006,N_10208,N_9512);
xor U14007 (N_14007,N_9605,N_11712);
nor U14008 (N_14008,N_9171,N_9785);
xor U14009 (N_14009,N_9672,N_11155);
nor U14010 (N_14010,N_10549,N_11937);
xnor U14011 (N_14011,N_10384,N_11974);
xor U14012 (N_14012,N_10782,N_10050);
nand U14013 (N_14013,N_9570,N_9321);
xnor U14014 (N_14014,N_10474,N_9368);
xnor U14015 (N_14015,N_9201,N_9115);
nand U14016 (N_14016,N_9175,N_10373);
xnor U14017 (N_14017,N_9262,N_10351);
or U14018 (N_14018,N_9254,N_10273);
nand U14019 (N_14019,N_11474,N_11743);
nand U14020 (N_14020,N_9230,N_11393);
and U14021 (N_14021,N_9446,N_10513);
and U14022 (N_14022,N_11488,N_11774);
nand U14023 (N_14023,N_11574,N_9096);
nor U14024 (N_14024,N_10256,N_11913);
or U14025 (N_14025,N_9281,N_10947);
nor U14026 (N_14026,N_11708,N_10205);
or U14027 (N_14027,N_10075,N_9263);
or U14028 (N_14028,N_9739,N_10956);
and U14029 (N_14029,N_11059,N_9484);
nor U14030 (N_14030,N_9951,N_9621);
or U14031 (N_14031,N_11973,N_9192);
xnor U14032 (N_14032,N_10983,N_9262);
nor U14033 (N_14033,N_9021,N_11415);
nand U14034 (N_14034,N_9567,N_9068);
or U14035 (N_14035,N_10791,N_9769);
and U14036 (N_14036,N_9982,N_11226);
nand U14037 (N_14037,N_11977,N_9113);
nand U14038 (N_14038,N_10580,N_11275);
or U14039 (N_14039,N_10361,N_10455);
xor U14040 (N_14040,N_9637,N_9755);
or U14041 (N_14041,N_10331,N_9979);
or U14042 (N_14042,N_10254,N_9520);
xor U14043 (N_14043,N_11801,N_9659);
xnor U14044 (N_14044,N_11716,N_11165);
nand U14045 (N_14045,N_9775,N_11079);
nand U14046 (N_14046,N_11206,N_10836);
nor U14047 (N_14047,N_9812,N_10752);
nand U14048 (N_14048,N_9612,N_9236);
xor U14049 (N_14049,N_11658,N_9205);
or U14050 (N_14050,N_9924,N_10159);
or U14051 (N_14051,N_11816,N_9309);
or U14052 (N_14052,N_9506,N_9479);
xnor U14053 (N_14053,N_10402,N_10032);
nor U14054 (N_14054,N_11999,N_11577);
nor U14055 (N_14055,N_11693,N_11333);
nand U14056 (N_14056,N_9341,N_11508);
nor U14057 (N_14057,N_11537,N_9202);
nand U14058 (N_14058,N_9099,N_9646);
and U14059 (N_14059,N_9084,N_9360);
and U14060 (N_14060,N_11925,N_10990);
xor U14061 (N_14061,N_10809,N_9358);
nor U14062 (N_14062,N_11171,N_10937);
nand U14063 (N_14063,N_11779,N_9336);
nand U14064 (N_14064,N_9870,N_10410);
nand U14065 (N_14065,N_11259,N_11498);
or U14066 (N_14066,N_10931,N_11621);
xor U14067 (N_14067,N_9232,N_11102);
nor U14068 (N_14068,N_10664,N_11623);
nor U14069 (N_14069,N_11740,N_11227);
nand U14070 (N_14070,N_10552,N_10462);
nand U14071 (N_14071,N_11552,N_9604);
xnor U14072 (N_14072,N_9131,N_9875);
nor U14073 (N_14073,N_10815,N_9293);
nand U14074 (N_14074,N_11048,N_9813);
nor U14075 (N_14075,N_11542,N_9007);
or U14076 (N_14076,N_11708,N_9170);
and U14077 (N_14077,N_11124,N_9891);
and U14078 (N_14078,N_9569,N_9600);
or U14079 (N_14079,N_10285,N_10933);
xnor U14080 (N_14080,N_10445,N_10387);
nor U14081 (N_14081,N_10143,N_10072);
and U14082 (N_14082,N_11935,N_11700);
nor U14083 (N_14083,N_11602,N_9404);
nand U14084 (N_14084,N_9486,N_9299);
or U14085 (N_14085,N_10989,N_10098);
and U14086 (N_14086,N_9376,N_9550);
xnor U14087 (N_14087,N_10812,N_9834);
xnor U14088 (N_14088,N_10254,N_10087);
xnor U14089 (N_14089,N_10469,N_10232);
xor U14090 (N_14090,N_10405,N_9516);
nand U14091 (N_14091,N_10814,N_11115);
nand U14092 (N_14092,N_11380,N_11403);
nand U14093 (N_14093,N_11754,N_9508);
nand U14094 (N_14094,N_11565,N_11451);
xor U14095 (N_14095,N_11821,N_11953);
nor U14096 (N_14096,N_11339,N_11638);
xor U14097 (N_14097,N_11737,N_10634);
nand U14098 (N_14098,N_11646,N_10080);
and U14099 (N_14099,N_9770,N_10539);
nor U14100 (N_14100,N_9094,N_10474);
nor U14101 (N_14101,N_9154,N_11730);
nand U14102 (N_14102,N_9789,N_11969);
nor U14103 (N_14103,N_10202,N_10396);
nor U14104 (N_14104,N_10502,N_10590);
and U14105 (N_14105,N_10208,N_11078);
nand U14106 (N_14106,N_9076,N_10670);
nor U14107 (N_14107,N_11009,N_9168);
nand U14108 (N_14108,N_9389,N_11022);
and U14109 (N_14109,N_11273,N_11906);
nand U14110 (N_14110,N_10595,N_11720);
xor U14111 (N_14111,N_10882,N_11386);
or U14112 (N_14112,N_11132,N_9884);
or U14113 (N_14113,N_10227,N_10604);
and U14114 (N_14114,N_9492,N_10218);
or U14115 (N_14115,N_10909,N_11617);
and U14116 (N_14116,N_9518,N_11132);
nor U14117 (N_14117,N_11088,N_9990);
and U14118 (N_14118,N_11934,N_11187);
or U14119 (N_14119,N_11431,N_10177);
and U14120 (N_14120,N_10699,N_11287);
nor U14121 (N_14121,N_11332,N_11314);
nand U14122 (N_14122,N_9291,N_9240);
nor U14123 (N_14123,N_11800,N_11303);
and U14124 (N_14124,N_9162,N_11804);
and U14125 (N_14125,N_9017,N_10760);
xor U14126 (N_14126,N_11527,N_9717);
or U14127 (N_14127,N_11922,N_10016);
nor U14128 (N_14128,N_11445,N_11821);
nor U14129 (N_14129,N_9039,N_10569);
nor U14130 (N_14130,N_10175,N_9248);
nor U14131 (N_14131,N_11229,N_11611);
nand U14132 (N_14132,N_10577,N_10679);
or U14133 (N_14133,N_10495,N_10687);
nand U14134 (N_14134,N_9851,N_10908);
nor U14135 (N_14135,N_10183,N_10626);
xor U14136 (N_14136,N_9390,N_10136);
or U14137 (N_14137,N_11140,N_9288);
xnor U14138 (N_14138,N_10038,N_11372);
or U14139 (N_14139,N_9978,N_11235);
or U14140 (N_14140,N_9888,N_9866);
and U14141 (N_14141,N_9537,N_11599);
nand U14142 (N_14142,N_11080,N_11911);
nor U14143 (N_14143,N_10811,N_11045);
nand U14144 (N_14144,N_10431,N_11503);
nand U14145 (N_14145,N_11250,N_11551);
or U14146 (N_14146,N_9887,N_10597);
and U14147 (N_14147,N_10954,N_10180);
or U14148 (N_14148,N_11118,N_11342);
nand U14149 (N_14149,N_11397,N_10586);
or U14150 (N_14150,N_11614,N_9363);
or U14151 (N_14151,N_11038,N_11403);
and U14152 (N_14152,N_11089,N_10900);
and U14153 (N_14153,N_9462,N_11389);
nand U14154 (N_14154,N_11112,N_11587);
nor U14155 (N_14155,N_9263,N_10548);
nand U14156 (N_14156,N_11946,N_10243);
nand U14157 (N_14157,N_9188,N_9366);
nor U14158 (N_14158,N_9334,N_9810);
nand U14159 (N_14159,N_10811,N_10612);
nor U14160 (N_14160,N_11677,N_9398);
or U14161 (N_14161,N_11647,N_11496);
nand U14162 (N_14162,N_10877,N_9906);
and U14163 (N_14163,N_9196,N_10765);
nor U14164 (N_14164,N_10553,N_10443);
and U14165 (N_14165,N_9213,N_10831);
xor U14166 (N_14166,N_9586,N_11789);
nand U14167 (N_14167,N_11593,N_11143);
or U14168 (N_14168,N_11256,N_10294);
nor U14169 (N_14169,N_11801,N_11995);
or U14170 (N_14170,N_11059,N_10002);
xor U14171 (N_14171,N_9990,N_9913);
nand U14172 (N_14172,N_9849,N_10858);
and U14173 (N_14173,N_11029,N_9180);
and U14174 (N_14174,N_10766,N_9000);
or U14175 (N_14175,N_9888,N_10159);
and U14176 (N_14176,N_10683,N_9023);
or U14177 (N_14177,N_10087,N_11650);
or U14178 (N_14178,N_11320,N_11389);
nand U14179 (N_14179,N_9631,N_9060);
and U14180 (N_14180,N_11524,N_10896);
and U14181 (N_14181,N_10138,N_11060);
or U14182 (N_14182,N_11076,N_10526);
nand U14183 (N_14183,N_10602,N_10697);
or U14184 (N_14184,N_11156,N_10668);
nand U14185 (N_14185,N_11631,N_9982);
nand U14186 (N_14186,N_11467,N_10032);
nand U14187 (N_14187,N_9104,N_9049);
nor U14188 (N_14188,N_11401,N_11269);
or U14189 (N_14189,N_9384,N_9807);
and U14190 (N_14190,N_9130,N_11482);
nor U14191 (N_14191,N_11041,N_11068);
nand U14192 (N_14192,N_11179,N_9594);
nor U14193 (N_14193,N_10170,N_10575);
or U14194 (N_14194,N_9809,N_11771);
xnor U14195 (N_14195,N_10949,N_11906);
xor U14196 (N_14196,N_11771,N_11370);
nand U14197 (N_14197,N_10831,N_10737);
and U14198 (N_14198,N_9602,N_10258);
and U14199 (N_14199,N_11954,N_9837);
nand U14200 (N_14200,N_11278,N_10906);
xnor U14201 (N_14201,N_9661,N_9706);
and U14202 (N_14202,N_9394,N_10766);
nand U14203 (N_14203,N_11108,N_9141);
xor U14204 (N_14204,N_9462,N_10188);
and U14205 (N_14205,N_9937,N_9907);
xnor U14206 (N_14206,N_11231,N_10754);
xnor U14207 (N_14207,N_10410,N_11993);
nand U14208 (N_14208,N_11230,N_10386);
nor U14209 (N_14209,N_11592,N_11044);
or U14210 (N_14210,N_9148,N_10637);
xnor U14211 (N_14211,N_10974,N_10929);
and U14212 (N_14212,N_10247,N_10718);
nor U14213 (N_14213,N_10816,N_9755);
nand U14214 (N_14214,N_11794,N_9321);
or U14215 (N_14215,N_11849,N_9958);
and U14216 (N_14216,N_11051,N_10159);
xnor U14217 (N_14217,N_9854,N_9549);
xnor U14218 (N_14218,N_9408,N_9721);
or U14219 (N_14219,N_10671,N_9632);
or U14220 (N_14220,N_11416,N_9127);
and U14221 (N_14221,N_10224,N_10725);
and U14222 (N_14222,N_11523,N_10891);
xor U14223 (N_14223,N_10054,N_10648);
nand U14224 (N_14224,N_9619,N_11631);
nand U14225 (N_14225,N_9158,N_10957);
nand U14226 (N_14226,N_9169,N_11887);
nand U14227 (N_14227,N_10227,N_9136);
xnor U14228 (N_14228,N_10638,N_11088);
or U14229 (N_14229,N_11610,N_10559);
or U14230 (N_14230,N_10003,N_10581);
nand U14231 (N_14231,N_9667,N_11342);
nand U14232 (N_14232,N_11865,N_9368);
and U14233 (N_14233,N_10217,N_9848);
xor U14234 (N_14234,N_9093,N_11775);
or U14235 (N_14235,N_11176,N_10597);
nand U14236 (N_14236,N_10243,N_9440);
xnor U14237 (N_14237,N_11963,N_10803);
or U14238 (N_14238,N_10009,N_11831);
nor U14239 (N_14239,N_9039,N_11030);
nor U14240 (N_14240,N_10198,N_10745);
or U14241 (N_14241,N_10208,N_10023);
nand U14242 (N_14242,N_9280,N_9503);
nor U14243 (N_14243,N_10152,N_10007);
or U14244 (N_14244,N_10555,N_9581);
nor U14245 (N_14245,N_11625,N_9312);
xnor U14246 (N_14246,N_11537,N_11598);
xor U14247 (N_14247,N_11490,N_9383);
nand U14248 (N_14248,N_11678,N_10423);
or U14249 (N_14249,N_10427,N_9315);
nand U14250 (N_14250,N_11525,N_11540);
nor U14251 (N_14251,N_10658,N_9383);
and U14252 (N_14252,N_9643,N_9861);
nor U14253 (N_14253,N_9825,N_9482);
and U14254 (N_14254,N_11943,N_9350);
xnor U14255 (N_14255,N_11339,N_10417);
or U14256 (N_14256,N_11112,N_9238);
and U14257 (N_14257,N_11770,N_9420);
xor U14258 (N_14258,N_11328,N_11467);
xnor U14259 (N_14259,N_10268,N_9838);
nand U14260 (N_14260,N_10707,N_10291);
xnor U14261 (N_14261,N_11643,N_9033);
xor U14262 (N_14262,N_11705,N_11792);
or U14263 (N_14263,N_10795,N_9516);
or U14264 (N_14264,N_10174,N_11057);
or U14265 (N_14265,N_10927,N_11893);
nor U14266 (N_14266,N_9919,N_10184);
and U14267 (N_14267,N_9933,N_10677);
xnor U14268 (N_14268,N_9528,N_11986);
xor U14269 (N_14269,N_9181,N_10396);
nand U14270 (N_14270,N_9096,N_11163);
and U14271 (N_14271,N_9782,N_10643);
nor U14272 (N_14272,N_11410,N_11043);
nor U14273 (N_14273,N_10842,N_9321);
or U14274 (N_14274,N_11568,N_9092);
or U14275 (N_14275,N_9124,N_11361);
xor U14276 (N_14276,N_11553,N_10126);
nor U14277 (N_14277,N_10687,N_10134);
xor U14278 (N_14278,N_9340,N_11941);
nor U14279 (N_14279,N_9273,N_11391);
nand U14280 (N_14280,N_10727,N_9545);
or U14281 (N_14281,N_10529,N_10998);
nor U14282 (N_14282,N_9383,N_10696);
xnor U14283 (N_14283,N_10710,N_9184);
and U14284 (N_14284,N_11145,N_11837);
or U14285 (N_14285,N_11518,N_11179);
xnor U14286 (N_14286,N_9408,N_9981);
or U14287 (N_14287,N_9633,N_11227);
nor U14288 (N_14288,N_11376,N_11825);
or U14289 (N_14289,N_9677,N_11477);
nor U14290 (N_14290,N_11382,N_10264);
nand U14291 (N_14291,N_11263,N_9989);
xnor U14292 (N_14292,N_9763,N_10902);
or U14293 (N_14293,N_9906,N_9102);
xor U14294 (N_14294,N_9711,N_10458);
nor U14295 (N_14295,N_9484,N_9193);
nor U14296 (N_14296,N_10602,N_10095);
nor U14297 (N_14297,N_9843,N_10005);
nand U14298 (N_14298,N_10436,N_10805);
or U14299 (N_14299,N_10895,N_11621);
xnor U14300 (N_14300,N_10810,N_9700);
xor U14301 (N_14301,N_11433,N_10576);
nor U14302 (N_14302,N_9032,N_9077);
nor U14303 (N_14303,N_11386,N_9018);
or U14304 (N_14304,N_11053,N_9263);
and U14305 (N_14305,N_9799,N_11905);
nand U14306 (N_14306,N_11614,N_11455);
xor U14307 (N_14307,N_11974,N_10942);
nand U14308 (N_14308,N_9852,N_9919);
and U14309 (N_14309,N_10508,N_10234);
nor U14310 (N_14310,N_11890,N_10093);
nor U14311 (N_14311,N_10275,N_10676);
or U14312 (N_14312,N_11946,N_10608);
xor U14313 (N_14313,N_10207,N_9696);
nand U14314 (N_14314,N_11388,N_11331);
or U14315 (N_14315,N_10771,N_9225);
nor U14316 (N_14316,N_10304,N_9502);
or U14317 (N_14317,N_10289,N_9614);
nor U14318 (N_14318,N_11340,N_10893);
nand U14319 (N_14319,N_9911,N_9916);
xor U14320 (N_14320,N_11347,N_11466);
or U14321 (N_14321,N_11461,N_11825);
nand U14322 (N_14322,N_9646,N_10823);
nand U14323 (N_14323,N_11893,N_11158);
nor U14324 (N_14324,N_10461,N_9797);
and U14325 (N_14325,N_9471,N_11150);
nor U14326 (N_14326,N_11157,N_9528);
nand U14327 (N_14327,N_10029,N_9121);
nand U14328 (N_14328,N_9700,N_9139);
and U14329 (N_14329,N_9647,N_9808);
xnor U14330 (N_14330,N_11847,N_11951);
nor U14331 (N_14331,N_10719,N_10456);
or U14332 (N_14332,N_9438,N_9783);
xor U14333 (N_14333,N_11282,N_9474);
nand U14334 (N_14334,N_9896,N_10608);
nand U14335 (N_14335,N_10674,N_10797);
xor U14336 (N_14336,N_10043,N_11788);
nand U14337 (N_14337,N_9386,N_10970);
and U14338 (N_14338,N_11941,N_9489);
or U14339 (N_14339,N_10064,N_11305);
and U14340 (N_14340,N_9680,N_10488);
and U14341 (N_14341,N_11721,N_9044);
nand U14342 (N_14342,N_10376,N_10043);
or U14343 (N_14343,N_9632,N_10466);
nand U14344 (N_14344,N_9129,N_11193);
and U14345 (N_14345,N_9152,N_10700);
xor U14346 (N_14346,N_9102,N_9268);
or U14347 (N_14347,N_9079,N_10192);
xnor U14348 (N_14348,N_9813,N_9301);
and U14349 (N_14349,N_11811,N_9605);
nand U14350 (N_14350,N_11497,N_9537);
nor U14351 (N_14351,N_10793,N_9232);
nand U14352 (N_14352,N_9237,N_11936);
and U14353 (N_14353,N_10561,N_9442);
xor U14354 (N_14354,N_11581,N_11571);
xnor U14355 (N_14355,N_10842,N_10248);
xnor U14356 (N_14356,N_9552,N_9563);
nand U14357 (N_14357,N_11597,N_11751);
or U14358 (N_14358,N_9681,N_10166);
nand U14359 (N_14359,N_10593,N_11233);
xnor U14360 (N_14360,N_10141,N_11360);
and U14361 (N_14361,N_10762,N_11802);
and U14362 (N_14362,N_9059,N_9903);
or U14363 (N_14363,N_11713,N_9528);
or U14364 (N_14364,N_10985,N_11964);
xor U14365 (N_14365,N_10223,N_9983);
nand U14366 (N_14366,N_10041,N_9435);
and U14367 (N_14367,N_9696,N_10830);
xor U14368 (N_14368,N_10499,N_11520);
and U14369 (N_14369,N_10899,N_10216);
nor U14370 (N_14370,N_11727,N_9475);
nand U14371 (N_14371,N_10212,N_11404);
or U14372 (N_14372,N_10508,N_9647);
and U14373 (N_14373,N_9712,N_9185);
or U14374 (N_14374,N_9696,N_11398);
or U14375 (N_14375,N_9805,N_9733);
nor U14376 (N_14376,N_11180,N_9189);
nand U14377 (N_14377,N_9466,N_11720);
nor U14378 (N_14378,N_11804,N_11894);
xnor U14379 (N_14379,N_11649,N_10871);
nand U14380 (N_14380,N_11665,N_11591);
or U14381 (N_14381,N_10683,N_10949);
nand U14382 (N_14382,N_10631,N_10609);
and U14383 (N_14383,N_11435,N_10236);
nor U14384 (N_14384,N_10812,N_9723);
nor U14385 (N_14385,N_9506,N_9530);
nand U14386 (N_14386,N_9330,N_10900);
nor U14387 (N_14387,N_10556,N_9994);
nand U14388 (N_14388,N_9159,N_9941);
nor U14389 (N_14389,N_10478,N_11017);
xor U14390 (N_14390,N_9272,N_11255);
or U14391 (N_14391,N_10597,N_10237);
xnor U14392 (N_14392,N_10040,N_11166);
nand U14393 (N_14393,N_11684,N_9431);
or U14394 (N_14394,N_9423,N_10078);
nor U14395 (N_14395,N_9994,N_11527);
xnor U14396 (N_14396,N_11053,N_11103);
nor U14397 (N_14397,N_9472,N_9278);
nand U14398 (N_14398,N_9511,N_9380);
and U14399 (N_14399,N_9258,N_9256);
or U14400 (N_14400,N_10101,N_10082);
xnor U14401 (N_14401,N_9742,N_10296);
and U14402 (N_14402,N_9275,N_9054);
nand U14403 (N_14403,N_9999,N_9560);
and U14404 (N_14404,N_10778,N_9654);
xor U14405 (N_14405,N_9604,N_10698);
nand U14406 (N_14406,N_10911,N_11390);
nand U14407 (N_14407,N_9962,N_11714);
xor U14408 (N_14408,N_10205,N_9370);
and U14409 (N_14409,N_10907,N_9181);
xor U14410 (N_14410,N_11463,N_11364);
xnor U14411 (N_14411,N_11724,N_11181);
and U14412 (N_14412,N_11791,N_11116);
nor U14413 (N_14413,N_9477,N_9046);
nor U14414 (N_14414,N_11439,N_10224);
or U14415 (N_14415,N_11603,N_9590);
or U14416 (N_14416,N_11474,N_10858);
or U14417 (N_14417,N_11944,N_11314);
nor U14418 (N_14418,N_11504,N_9445);
and U14419 (N_14419,N_9737,N_11485);
xor U14420 (N_14420,N_10683,N_10472);
nand U14421 (N_14421,N_10408,N_11913);
and U14422 (N_14422,N_11531,N_9231);
or U14423 (N_14423,N_9413,N_11467);
nand U14424 (N_14424,N_11272,N_9785);
xor U14425 (N_14425,N_11752,N_11616);
and U14426 (N_14426,N_10615,N_9411);
xnor U14427 (N_14427,N_9170,N_11011);
or U14428 (N_14428,N_11069,N_10610);
or U14429 (N_14429,N_10286,N_10453);
or U14430 (N_14430,N_9017,N_10661);
nor U14431 (N_14431,N_9337,N_9455);
xnor U14432 (N_14432,N_11496,N_9016);
nand U14433 (N_14433,N_10536,N_9138);
or U14434 (N_14434,N_11066,N_10954);
nand U14435 (N_14435,N_11290,N_10456);
xor U14436 (N_14436,N_10152,N_9045);
nand U14437 (N_14437,N_11764,N_9221);
and U14438 (N_14438,N_11283,N_10789);
nand U14439 (N_14439,N_10053,N_9916);
nor U14440 (N_14440,N_9892,N_10169);
xnor U14441 (N_14441,N_10004,N_9500);
and U14442 (N_14442,N_11133,N_9990);
nand U14443 (N_14443,N_10188,N_10310);
and U14444 (N_14444,N_10357,N_10747);
or U14445 (N_14445,N_9272,N_10123);
nand U14446 (N_14446,N_10616,N_11209);
nand U14447 (N_14447,N_10148,N_10246);
nor U14448 (N_14448,N_11523,N_9009);
nand U14449 (N_14449,N_11402,N_9820);
xnor U14450 (N_14450,N_10457,N_9391);
and U14451 (N_14451,N_9441,N_11247);
nor U14452 (N_14452,N_9970,N_10944);
nor U14453 (N_14453,N_10719,N_11006);
nor U14454 (N_14454,N_11267,N_9165);
nor U14455 (N_14455,N_11537,N_10194);
xor U14456 (N_14456,N_9322,N_10896);
xor U14457 (N_14457,N_11529,N_10225);
nor U14458 (N_14458,N_9433,N_10003);
nor U14459 (N_14459,N_9704,N_11189);
or U14460 (N_14460,N_10347,N_11394);
or U14461 (N_14461,N_9898,N_10990);
nand U14462 (N_14462,N_11245,N_10480);
or U14463 (N_14463,N_9707,N_11160);
and U14464 (N_14464,N_10832,N_11322);
nand U14465 (N_14465,N_11812,N_9525);
xnor U14466 (N_14466,N_9639,N_9988);
and U14467 (N_14467,N_9639,N_11899);
and U14468 (N_14468,N_11984,N_11080);
xnor U14469 (N_14469,N_11139,N_11766);
or U14470 (N_14470,N_9849,N_10404);
and U14471 (N_14471,N_9036,N_10742);
xor U14472 (N_14472,N_9488,N_10649);
nand U14473 (N_14473,N_9692,N_9642);
and U14474 (N_14474,N_11577,N_11174);
or U14475 (N_14475,N_9632,N_11096);
or U14476 (N_14476,N_11097,N_11793);
nor U14477 (N_14477,N_9953,N_9612);
nor U14478 (N_14478,N_11076,N_10609);
nand U14479 (N_14479,N_10966,N_11665);
nand U14480 (N_14480,N_9473,N_9194);
nor U14481 (N_14481,N_10926,N_11600);
nor U14482 (N_14482,N_10785,N_11974);
xnor U14483 (N_14483,N_10187,N_11254);
or U14484 (N_14484,N_9738,N_11992);
and U14485 (N_14485,N_9645,N_9293);
nand U14486 (N_14486,N_10032,N_11598);
or U14487 (N_14487,N_9075,N_11933);
and U14488 (N_14488,N_10119,N_11302);
and U14489 (N_14489,N_10787,N_11252);
nand U14490 (N_14490,N_10680,N_11724);
and U14491 (N_14491,N_9591,N_10531);
xor U14492 (N_14492,N_9657,N_9970);
xnor U14493 (N_14493,N_10482,N_11728);
nor U14494 (N_14494,N_9566,N_11897);
and U14495 (N_14495,N_10847,N_10795);
xnor U14496 (N_14496,N_9243,N_11973);
or U14497 (N_14497,N_9833,N_9484);
nor U14498 (N_14498,N_11371,N_10890);
and U14499 (N_14499,N_10666,N_9505);
xnor U14500 (N_14500,N_11875,N_11961);
nor U14501 (N_14501,N_10113,N_9805);
or U14502 (N_14502,N_10156,N_9506);
and U14503 (N_14503,N_9579,N_11592);
xnor U14504 (N_14504,N_10234,N_11907);
or U14505 (N_14505,N_9292,N_10710);
nand U14506 (N_14506,N_10899,N_9426);
or U14507 (N_14507,N_9765,N_9143);
or U14508 (N_14508,N_11706,N_10372);
xor U14509 (N_14509,N_9671,N_11926);
or U14510 (N_14510,N_10982,N_10147);
and U14511 (N_14511,N_11079,N_11723);
or U14512 (N_14512,N_9217,N_10732);
and U14513 (N_14513,N_11298,N_9363);
nand U14514 (N_14514,N_10140,N_10446);
nand U14515 (N_14515,N_11664,N_11353);
or U14516 (N_14516,N_11223,N_10785);
nand U14517 (N_14517,N_10043,N_10922);
and U14518 (N_14518,N_10453,N_11425);
or U14519 (N_14519,N_9873,N_11198);
nor U14520 (N_14520,N_10189,N_10998);
nand U14521 (N_14521,N_10952,N_9364);
or U14522 (N_14522,N_10595,N_11251);
or U14523 (N_14523,N_11416,N_10262);
or U14524 (N_14524,N_11712,N_11651);
and U14525 (N_14525,N_10176,N_10325);
nor U14526 (N_14526,N_11972,N_10753);
or U14527 (N_14527,N_11811,N_10288);
nand U14528 (N_14528,N_9880,N_10872);
and U14529 (N_14529,N_11060,N_10356);
xor U14530 (N_14530,N_11293,N_11147);
or U14531 (N_14531,N_11572,N_10359);
xor U14532 (N_14532,N_9500,N_9786);
and U14533 (N_14533,N_11639,N_9037);
and U14534 (N_14534,N_9839,N_10797);
nand U14535 (N_14535,N_10993,N_10335);
xnor U14536 (N_14536,N_10251,N_11542);
or U14537 (N_14537,N_9386,N_11861);
and U14538 (N_14538,N_10662,N_11958);
nand U14539 (N_14539,N_10432,N_11546);
xor U14540 (N_14540,N_11786,N_11951);
nor U14541 (N_14541,N_10373,N_11004);
and U14542 (N_14542,N_9392,N_10755);
nand U14543 (N_14543,N_10877,N_9574);
nand U14544 (N_14544,N_9520,N_11058);
nor U14545 (N_14545,N_9999,N_9781);
or U14546 (N_14546,N_9462,N_10540);
nand U14547 (N_14547,N_11718,N_9113);
and U14548 (N_14548,N_9123,N_11930);
or U14549 (N_14549,N_11800,N_11148);
nor U14550 (N_14550,N_10244,N_11892);
xnor U14551 (N_14551,N_10358,N_10711);
or U14552 (N_14552,N_9770,N_9280);
xor U14553 (N_14553,N_9214,N_11805);
and U14554 (N_14554,N_9752,N_11127);
and U14555 (N_14555,N_9082,N_11167);
and U14556 (N_14556,N_9896,N_11118);
nor U14557 (N_14557,N_10788,N_11438);
nor U14558 (N_14558,N_11624,N_11152);
xor U14559 (N_14559,N_11419,N_9566);
xnor U14560 (N_14560,N_9658,N_9055);
nand U14561 (N_14561,N_9101,N_11036);
or U14562 (N_14562,N_11890,N_11888);
xnor U14563 (N_14563,N_9629,N_11562);
or U14564 (N_14564,N_11330,N_10791);
nand U14565 (N_14565,N_11234,N_10531);
xnor U14566 (N_14566,N_10773,N_9487);
nand U14567 (N_14567,N_10700,N_9147);
xnor U14568 (N_14568,N_9452,N_11260);
xor U14569 (N_14569,N_9761,N_9912);
or U14570 (N_14570,N_10031,N_9341);
or U14571 (N_14571,N_11378,N_10985);
nand U14572 (N_14572,N_10204,N_11860);
and U14573 (N_14573,N_10746,N_11498);
nor U14574 (N_14574,N_9007,N_9333);
or U14575 (N_14575,N_9650,N_10264);
nor U14576 (N_14576,N_10517,N_11463);
and U14577 (N_14577,N_11219,N_11918);
and U14578 (N_14578,N_11173,N_9642);
and U14579 (N_14579,N_10516,N_9229);
and U14580 (N_14580,N_11658,N_10057);
nand U14581 (N_14581,N_11951,N_11231);
and U14582 (N_14582,N_9542,N_9156);
and U14583 (N_14583,N_10189,N_11117);
nand U14584 (N_14584,N_10992,N_10742);
xor U14585 (N_14585,N_9434,N_11955);
nor U14586 (N_14586,N_10491,N_10672);
xor U14587 (N_14587,N_11636,N_11814);
xnor U14588 (N_14588,N_11067,N_10177);
xor U14589 (N_14589,N_11242,N_11394);
and U14590 (N_14590,N_9286,N_10187);
nand U14591 (N_14591,N_9791,N_9684);
nand U14592 (N_14592,N_10140,N_9742);
or U14593 (N_14593,N_11088,N_11605);
xnor U14594 (N_14594,N_9884,N_11329);
or U14595 (N_14595,N_10302,N_10871);
xnor U14596 (N_14596,N_9309,N_11620);
or U14597 (N_14597,N_10261,N_9497);
xor U14598 (N_14598,N_11305,N_10950);
nand U14599 (N_14599,N_10684,N_9162);
and U14600 (N_14600,N_10570,N_10551);
nor U14601 (N_14601,N_11868,N_11140);
and U14602 (N_14602,N_9475,N_9648);
nand U14603 (N_14603,N_11462,N_9278);
xor U14604 (N_14604,N_10151,N_11261);
nand U14605 (N_14605,N_10310,N_10849);
and U14606 (N_14606,N_9223,N_10560);
nor U14607 (N_14607,N_11251,N_11328);
and U14608 (N_14608,N_9797,N_9194);
and U14609 (N_14609,N_11997,N_11120);
nand U14610 (N_14610,N_10270,N_10702);
xnor U14611 (N_14611,N_10075,N_11080);
and U14612 (N_14612,N_9748,N_11489);
and U14613 (N_14613,N_9144,N_9005);
xnor U14614 (N_14614,N_9983,N_9737);
nand U14615 (N_14615,N_10489,N_9585);
or U14616 (N_14616,N_9754,N_10298);
or U14617 (N_14617,N_9887,N_11459);
or U14618 (N_14618,N_10094,N_11401);
and U14619 (N_14619,N_10165,N_10839);
nor U14620 (N_14620,N_9056,N_9683);
nor U14621 (N_14621,N_11092,N_10787);
nand U14622 (N_14622,N_9431,N_10226);
xnor U14623 (N_14623,N_10834,N_9164);
nor U14624 (N_14624,N_9868,N_10910);
and U14625 (N_14625,N_11910,N_11555);
nand U14626 (N_14626,N_9021,N_9740);
or U14627 (N_14627,N_11837,N_11736);
xor U14628 (N_14628,N_11205,N_11020);
or U14629 (N_14629,N_10558,N_10138);
nand U14630 (N_14630,N_9930,N_9898);
and U14631 (N_14631,N_9061,N_10639);
xnor U14632 (N_14632,N_11015,N_11085);
nor U14633 (N_14633,N_9070,N_10481);
nand U14634 (N_14634,N_10345,N_9411);
nor U14635 (N_14635,N_11734,N_11708);
nand U14636 (N_14636,N_10521,N_11664);
xnor U14637 (N_14637,N_10277,N_10151);
and U14638 (N_14638,N_11725,N_10855);
nand U14639 (N_14639,N_11681,N_9381);
and U14640 (N_14640,N_9689,N_10936);
or U14641 (N_14641,N_9734,N_9782);
or U14642 (N_14642,N_9670,N_10987);
and U14643 (N_14643,N_11853,N_10706);
or U14644 (N_14644,N_11095,N_11275);
nor U14645 (N_14645,N_9514,N_11067);
nand U14646 (N_14646,N_11384,N_9818);
xor U14647 (N_14647,N_10999,N_11958);
xnor U14648 (N_14648,N_10382,N_11938);
nand U14649 (N_14649,N_9743,N_11271);
xor U14650 (N_14650,N_11751,N_9694);
xnor U14651 (N_14651,N_9385,N_10241);
and U14652 (N_14652,N_9542,N_11530);
nand U14653 (N_14653,N_9322,N_9400);
and U14654 (N_14654,N_9530,N_10059);
nor U14655 (N_14655,N_11146,N_10697);
nor U14656 (N_14656,N_10081,N_9161);
nor U14657 (N_14657,N_9461,N_9678);
nor U14658 (N_14658,N_9278,N_11944);
or U14659 (N_14659,N_10013,N_9684);
or U14660 (N_14660,N_11500,N_11760);
and U14661 (N_14661,N_9337,N_9188);
xnor U14662 (N_14662,N_10302,N_9521);
or U14663 (N_14663,N_10339,N_9357);
xnor U14664 (N_14664,N_9376,N_10602);
xnor U14665 (N_14665,N_11768,N_11071);
or U14666 (N_14666,N_10763,N_11009);
xnor U14667 (N_14667,N_9434,N_9938);
nor U14668 (N_14668,N_11447,N_10944);
nand U14669 (N_14669,N_9716,N_9525);
or U14670 (N_14670,N_10214,N_9192);
xnor U14671 (N_14671,N_10916,N_10075);
or U14672 (N_14672,N_10102,N_11283);
xnor U14673 (N_14673,N_9631,N_9886);
and U14674 (N_14674,N_10651,N_9824);
xnor U14675 (N_14675,N_11193,N_11007);
and U14676 (N_14676,N_9868,N_11710);
nor U14677 (N_14677,N_11968,N_11762);
xnor U14678 (N_14678,N_11123,N_11808);
xor U14679 (N_14679,N_11830,N_9937);
xor U14680 (N_14680,N_11048,N_10380);
xnor U14681 (N_14681,N_11486,N_11008);
nand U14682 (N_14682,N_11436,N_10378);
and U14683 (N_14683,N_11278,N_9244);
and U14684 (N_14684,N_10254,N_10679);
nand U14685 (N_14685,N_11951,N_9983);
nor U14686 (N_14686,N_11768,N_9826);
or U14687 (N_14687,N_9129,N_9987);
nor U14688 (N_14688,N_11864,N_10732);
nand U14689 (N_14689,N_9724,N_9939);
nand U14690 (N_14690,N_11961,N_10582);
and U14691 (N_14691,N_11844,N_9054);
and U14692 (N_14692,N_10880,N_11854);
nor U14693 (N_14693,N_11448,N_11047);
xnor U14694 (N_14694,N_11267,N_10689);
nor U14695 (N_14695,N_11399,N_10018);
and U14696 (N_14696,N_11058,N_9772);
nor U14697 (N_14697,N_11061,N_10621);
or U14698 (N_14698,N_11077,N_9355);
or U14699 (N_14699,N_10592,N_10390);
nor U14700 (N_14700,N_11333,N_11516);
nand U14701 (N_14701,N_11774,N_9556);
and U14702 (N_14702,N_10484,N_11364);
nand U14703 (N_14703,N_10294,N_10295);
nand U14704 (N_14704,N_11192,N_9924);
nand U14705 (N_14705,N_9827,N_10408);
or U14706 (N_14706,N_11076,N_10134);
nand U14707 (N_14707,N_9554,N_9800);
nand U14708 (N_14708,N_9492,N_11682);
and U14709 (N_14709,N_10921,N_10406);
and U14710 (N_14710,N_10978,N_10050);
nor U14711 (N_14711,N_9596,N_9270);
or U14712 (N_14712,N_11462,N_9322);
nand U14713 (N_14713,N_11058,N_9368);
xnor U14714 (N_14714,N_9727,N_10783);
and U14715 (N_14715,N_10520,N_10714);
xnor U14716 (N_14716,N_9394,N_11570);
xnor U14717 (N_14717,N_11845,N_9393);
nor U14718 (N_14718,N_11739,N_10378);
and U14719 (N_14719,N_11539,N_10759);
xor U14720 (N_14720,N_9096,N_10741);
and U14721 (N_14721,N_11081,N_9602);
xor U14722 (N_14722,N_9385,N_9937);
nand U14723 (N_14723,N_11692,N_11179);
or U14724 (N_14724,N_11280,N_9729);
xnor U14725 (N_14725,N_10165,N_11936);
nor U14726 (N_14726,N_9539,N_10631);
nand U14727 (N_14727,N_10617,N_9314);
nand U14728 (N_14728,N_11909,N_11694);
and U14729 (N_14729,N_9819,N_10827);
and U14730 (N_14730,N_9911,N_9387);
or U14731 (N_14731,N_11601,N_10779);
nand U14732 (N_14732,N_10807,N_10867);
or U14733 (N_14733,N_10923,N_10455);
and U14734 (N_14734,N_10887,N_10815);
and U14735 (N_14735,N_11631,N_10831);
xor U14736 (N_14736,N_9549,N_11972);
and U14737 (N_14737,N_11105,N_11779);
nor U14738 (N_14738,N_9078,N_11553);
and U14739 (N_14739,N_10018,N_10977);
nor U14740 (N_14740,N_9796,N_11756);
xor U14741 (N_14741,N_9100,N_10414);
nand U14742 (N_14742,N_11156,N_10523);
nor U14743 (N_14743,N_10457,N_10960);
and U14744 (N_14744,N_11818,N_10195);
nand U14745 (N_14745,N_10087,N_9563);
nand U14746 (N_14746,N_11503,N_11116);
nor U14747 (N_14747,N_10490,N_11911);
nand U14748 (N_14748,N_10775,N_9107);
xnor U14749 (N_14749,N_11920,N_10467);
nand U14750 (N_14750,N_10084,N_11946);
xnor U14751 (N_14751,N_11188,N_9277);
and U14752 (N_14752,N_10818,N_11376);
or U14753 (N_14753,N_10275,N_9136);
or U14754 (N_14754,N_10916,N_10550);
or U14755 (N_14755,N_10781,N_10078);
nor U14756 (N_14756,N_10459,N_11518);
nand U14757 (N_14757,N_9906,N_10347);
nand U14758 (N_14758,N_11806,N_10202);
or U14759 (N_14759,N_11624,N_9959);
and U14760 (N_14760,N_11822,N_9430);
nor U14761 (N_14761,N_11580,N_9456);
xor U14762 (N_14762,N_11577,N_10617);
or U14763 (N_14763,N_11976,N_9642);
xor U14764 (N_14764,N_10953,N_10981);
or U14765 (N_14765,N_11162,N_11534);
and U14766 (N_14766,N_9081,N_11598);
nor U14767 (N_14767,N_9980,N_9443);
and U14768 (N_14768,N_10664,N_9223);
nor U14769 (N_14769,N_11448,N_10702);
nor U14770 (N_14770,N_9257,N_9513);
xnor U14771 (N_14771,N_11461,N_11475);
or U14772 (N_14772,N_9044,N_9067);
or U14773 (N_14773,N_10558,N_11536);
and U14774 (N_14774,N_9540,N_10297);
and U14775 (N_14775,N_11552,N_10889);
or U14776 (N_14776,N_9478,N_11227);
nor U14777 (N_14777,N_10499,N_11502);
nand U14778 (N_14778,N_11834,N_9652);
xnor U14779 (N_14779,N_9651,N_9001);
xor U14780 (N_14780,N_9722,N_11450);
xor U14781 (N_14781,N_11180,N_11423);
or U14782 (N_14782,N_9476,N_11832);
nor U14783 (N_14783,N_10971,N_11228);
xnor U14784 (N_14784,N_11363,N_9267);
nand U14785 (N_14785,N_9674,N_11623);
nor U14786 (N_14786,N_11699,N_9984);
xor U14787 (N_14787,N_10720,N_10163);
nand U14788 (N_14788,N_11084,N_11115);
and U14789 (N_14789,N_11369,N_9018);
and U14790 (N_14790,N_9212,N_11984);
nor U14791 (N_14791,N_11224,N_10820);
nor U14792 (N_14792,N_10648,N_11283);
or U14793 (N_14793,N_11753,N_11895);
nor U14794 (N_14794,N_10934,N_11708);
nand U14795 (N_14795,N_11439,N_10962);
or U14796 (N_14796,N_10563,N_10192);
nor U14797 (N_14797,N_11209,N_9616);
xor U14798 (N_14798,N_11696,N_9953);
xor U14799 (N_14799,N_11269,N_9558);
and U14800 (N_14800,N_10042,N_11752);
nand U14801 (N_14801,N_11213,N_9144);
nor U14802 (N_14802,N_11199,N_10704);
and U14803 (N_14803,N_9875,N_9566);
or U14804 (N_14804,N_10673,N_10064);
nor U14805 (N_14805,N_10817,N_9405);
or U14806 (N_14806,N_11357,N_11102);
or U14807 (N_14807,N_11920,N_10807);
nand U14808 (N_14808,N_11882,N_10537);
and U14809 (N_14809,N_11929,N_10507);
xnor U14810 (N_14810,N_10223,N_10740);
xor U14811 (N_14811,N_10494,N_9969);
xnor U14812 (N_14812,N_9215,N_10489);
and U14813 (N_14813,N_9743,N_11864);
xnor U14814 (N_14814,N_9161,N_9076);
xnor U14815 (N_14815,N_11166,N_9467);
nor U14816 (N_14816,N_9913,N_11374);
xnor U14817 (N_14817,N_10333,N_9677);
or U14818 (N_14818,N_11908,N_9189);
nor U14819 (N_14819,N_10902,N_11507);
nor U14820 (N_14820,N_10301,N_10099);
nor U14821 (N_14821,N_9981,N_11481);
nor U14822 (N_14822,N_10939,N_10006);
xnor U14823 (N_14823,N_10049,N_10848);
or U14824 (N_14824,N_10072,N_9173);
xor U14825 (N_14825,N_9332,N_10899);
or U14826 (N_14826,N_10365,N_9663);
nor U14827 (N_14827,N_11500,N_10263);
or U14828 (N_14828,N_10355,N_11802);
or U14829 (N_14829,N_10986,N_11577);
nand U14830 (N_14830,N_11090,N_9701);
xnor U14831 (N_14831,N_10980,N_11345);
nand U14832 (N_14832,N_10523,N_10509);
xnor U14833 (N_14833,N_10170,N_11496);
xnor U14834 (N_14834,N_9455,N_9967);
and U14835 (N_14835,N_9364,N_9587);
nand U14836 (N_14836,N_10134,N_9738);
xnor U14837 (N_14837,N_11954,N_9024);
and U14838 (N_14838,N_11198,N_11081);
nand U14839 (N_14839,N_11020,N_10843);
xnor U14840 (N_14840,N_10476,N_10831);
and U14841 (N_14841,N_11603,N_11133);
nor U14842 (N_14842,N_11815,N_10224);
nand U14843 (N_14843,N_9924,N_10431);
nor U14844 (N_14844,N_10663,N_9068);
nand U14845 (N_14845,N_11658,N_10905);
nor U14846 (N_14846,N_10779,N_11135);
xor U14847 (N_14847,N_9030,N_11083);
nor U14848 (N_14848,N_11663,N_11277);
nor U14849 (N_14849,N_9663,N_10452);
and U14850 (N_14850,N_11457,N_10027);
nand U14851 (N_14851,N_9717,N_11571);
or U14852 (N_14852,N_10482,N_11155);
nand U14853 (N_14853,N_11902,N_9739);
nand U14854 (N_14854,N_10922,N_10068);
xor U14855 (N_14855,N_9597,N_11029);
nand U14856 (N_14856,N_9550,N_10175);
or U14857 (N_14857,N_11456,N_9338);
nor U14858 (N_14858,N_10155,N_10129);
nor U14859 (N_14859,N_10959,N_9007);
or U14860 (N_14860,N_11766,N_9540);
nor U14861 (N_14861,N_9879,N_9614);
nand U14862 (N_14862,N_10279,N_10289);
nor U14863 (N_14863,N_11826,N_9548);
or U14864 (N_14864,N_9072,N_10596);
or U14865 (N_14865,N_11780,N_10415);
and U14866 (N_14866,N_10089,N_9309);
nor U14867 (N_14867,N_9937,N_11061);
xor U14868 (N_14868,N_10702,N_9449);
or U14869 (N_14869,N_9229,N_9397);
and U14870 (N_14870,N_9930,N_9113);
nor U14871 (N_14871,N_11698,N_9975);
nand U14872 (N_14872,N_11603,N_9584);
and U14873 (N_14873,N_11322,N_9620);
and U14874 (N_14874,N_11548,N_11421);
xor U14875 (N_14875,N_10407,N_11207);
nand U14876 (N_14876,N_9863,N_9935);
and U14877 (N_14877,N_9535,N_11212);
nor U14878 (N_14878,N_10082,N_11480);
nand U14879 (N_14879,N_9133,N_9111);
and U14880 (N_14880,N_9172,N_9997);
or U14881 (N_14881,N_10152,N_10020);
xnor U14882 (N_14882,N_10935,N_10452);
and U14883 (N_14883,N_10678,N_11641);
or U14884 (N_14884,N_10976,N_9243);
and U14885 (N_14885,N_11973,N_11485);
nor U14886 (N_14886,N_11916,N_10351);
and U14887 (N_14887,N_9687,N_11039);
nand U14888 (N_14888,N_9849,N_9050);
nor U14889 (N_14889,N_11508,N_11985);
or U14890 (N_14890,N_9061,N_11940);
nor U14891 (N_14891,N_11463,N_9928);
nand U14892 (N_14892,N_10334,N_10821);
and U14893 (N_14893,N_11487,N_10126);
and U14894 (N_14894,N_11826,N_9478);
nand U14895 (N_14895,N_9595,N_11258);
nor U14896 (N_14896,N_11238,N_11609);
and U14897 (N_14897,N_9186,N_9889);
nand U14898 (N_14898,N_9540,N_9996);
xnor U14899 (N_14899,N_9741,N_11705);
nand U14900 (N_14900,N_10918,N_10688);
or U14901 (N_14901,N_9597,N_11207);
or U14902 (N_14902,N_9152,N_10588);
or U14903 (N_14903,N_9114,N_11439);
nor U14904 (N_14904,N_11982,N_10200);
or U14905 (N_14905,N_9283,N_10004);
or U14906 (N_14906,N_9618,N_11072);
nor U14907 (N_14907,N_11352,N_11860);
and U14908 (N_14908,N_11678,N_11104);
xnor U14909 (N_14909,N_10635,N_11723);
and U14910 (N_14910,N_9540,N_9942);
or U14911 (N_14911,N_11349,N_11574);
xnor U14912 (N_14912,N_10418,N_11561);
or U14913 (N_14913,N_9407,N_9346);
or U14914 (N_14914,N_10970,N_10549);
nand U14915 (N_14915,N_10958,N_9755);
nand U14916 (N_14916,N_11653,N_9825);
and U14917 (N_14917,N_10744,N_11286);
or U14918 (N_14918,N_10967,N_11094);
xor U14919 (N_14919,N_10202,N_10224);
or U14920 (N_14920,N_9463,N_11622);
nor U14921 (N_14921,N_10220,N_9247);
nand U14922 (N_14922,N_11025,N_11794);
nand U14923 (N_14923,N_10638,N_11931);
or U14924 (N_14924,N_10445,N_11489);
nand U14925 (N_14925,N_9195,N_10753);
nand U14926 (N_14926,N_11988,N_11139);
xor U14927 (N_14927,N_11508,N_9390);
nor U14928 (N_14928,N_9058,N_10448);
or U14929 (N_14929,N_11929,N_10207);
nand U14930 (N_14930,N_10429,N_9622);
or U14931 (N_14931,N_9659,N_9115);
nor U14932 (N_14932,N_11795,N_9162);
nor U14933 (N_14933,N_10723,N_9731);
nor U14934 (N_14934,N_10790,N_9488);
nand U14935 (N_14935,N_11308,N_11101);
nor U14936 (N_14936,N_10478,N_11289);
nand U14937 (N_14937,N_10253,N_9348);
nand U14938 (N_14938,N_11178,N_11110);
xor U14939 (N_14939,N_10366,N_9641);
xor U14940 (N_14940,N_11127,N_10147);
or U14941 (N_14941,N_11384,N_10132);
or U14942 (N_14942,N_10785,N_9406);
and U14943 (N_14943,N_10184,N_11078);
and U14944 (N_14944,N_11749,N_11862);
and U14945 (N_14945,N_11054,N_9999);
xor U14946 (N_14946,N_10823,N_11673);
or U14947 (N_14947,N_10526,N_11572);
nand U14948 (N_14948,N_9528,N_10636);
nor U14949 (N_14949,N_10935,N_10173);
and U14950 (N_14950,N_10937,N_9418);
and U14951 (N_14951,N_9844,N_10457);
and U14952 (N_14952,N_10902,N_9661);
nand U14953 (N_14953,N_10045,N_10392);
nand U14954 (N_14954,N_9505,N_10470);
and U14955 (N_14955,N_9222,N_11359);
xnor U14956 (N_14956,N_9236,N_9708);
nor U14957 (N_14957,N_9227,N_11932);
nor U14958 (N_14958,N_10661,N_11370);
nor U14959 (N_14959,N_11123,N_11610);
nand U14960 (N_14960,N_11445,N_11420);
or U14961 (N_14961,N_10288,N_11711);
nor U14962 (N_14962,N_11500,N_11014);
or U14963 (N_14963,N_9524,N_9683);
or U14964 (N_14964,N_9702,N_11590);
and U14965 (N_14965,N_9967,N_11328);
and U14966 (N_14966,N_9852,N_10449);
or U14967 (N_14967,N_9851,N_11251);
and U14968 (N_14968,N_11863,N_10733);
nand U14969 (N_14969,N_10799,N_10276);
and U14970 (N_14970,N_11864,N_10283);
and U14971 (N_14971,N_10395,N_9099);
nor U14972 (N_14972,N_11012,N_11607);
and U14973 (N_14973,N_9205,N_10859);
or U14974 (N_14974,N_9037,N_10592);
nor U14975 (N_14975,N_9856,N_11493);
nor U14976 (N_14976,N_10896,N_11796);
nand U14977 (N_14977,N_11415,N_9483);
xor U14978 (N_14978,N_9389,N_11052);
xnor U14979 (N_14979,N_10627,N_11929);
nand U14980 (N_14980,N_10893,N_9836);
xor U14981 (N_14981,N_9284,N_11321);
nor U14982 (N_14982,N_11835,N_9695);
and U14983 (N_14983,N_9387,N_9648);
xor U14984 (N_14984,N_9032,N_11382);
xnor U14985 (N_14985,N_9351,N_11403);
or U14986 (N_14986,N_9238,N_10347);
nand U14987 (N_14987,N_11495,N_11615);
and U14988 (N_14988,N_10871,N_11593);
xor U14989 (N_14989,N_11302,N_10180);
or U14990 (N_14990,N_9856,N_11481);
xor U14991 (N_14991,N_11687,N_10188);
xor U14992 (N_14992,N_9909,N_11336);
and U14993 (N_14993,N_10102,N_10908);
and U14994 (N_14994,N_10870,N_9254);
xor U14995 (N_14995,N_10856,N_10484);
or U14996 (N_14996,N_10377,N_10051);
nand U14997 (N_14997,N_10588,N_10878);
or U14998 (N_14998,N_10201,N_10855);
and U14999 (N_14999,N_11656,N_11823);
or UO_0 (O_0,N_13879,N_12076);
or UO_1 (O_1,N_14852,N_14213);
nand UO_2 (O_2,N_14865,N_14098);
nand UO_3 (O_3,N_13784,N_13649);
or UO_4 (O_4,N_13144,N_12267);
nand UO_5 (O_5,N_12516,N_13189);
or UO_6 (O_6,N_13221,N_14818);
and UO_7 (O_7,N_14206,N_13305);
nor UO_8 (O_8,N_13734,N_14186);
or UO_9 (O_9,N_14708,N_12639);
xor UO_10 (O_10,N_13004,N_12419);
nor UO_11 (O_11,N_13196,N_12604);
nand UO_12 (O_12,N_14718,N_13481);
nor UO_13 (O_13,N_14547,N_14975);
and UO_14 (O_14,N_14300,N_14240);
nor UO_15 (O_15,N_14605,N_14507);
or UO_16 (O_16,N_12589,N_14991);
xor UO_17 (O_17,N_13898,N_14824);
and UO_18 (O_18,N_14683,N_14389);
nand UO_19 (O_19,N_14519,N_12576);
xor UO_20 (O_20,N_13187,N_13044);
xor UO_21 (O_21,N_13880,N_12930);
xnor UO_22 (O_22,N_12495,N_12929);
xnor UO_23 (O_23,N_13813,N_13068);
or UO_24 (O_24,N_12425,N_12956);
or UO_25 (O_25,N_14413,N_13341);
xor UO_26 (O_26,N_13599,N_13596);
xor UO_27 (O_27,N_12831,N_12446);
or UO_28 (O_28,N_14575,N_13505);
xnor UO_29 (O_29,N_14280,N_12503);
xnor UO_30 (O_30,N_14781,N_13209);
nand UO_31 (O_31,N_12750,N_13316);
or UO_32 (O_32,N_14782,N_13574);
nand UO_33 (O_33,N_13936,N_14590);
or UO_34 (O_34,N_12209,N_13575);
nor UO_35 (O_35,N_13312,N_13901);
nand UO_36 (O_36,N_14842,N_14680);
and UO_37 (O_37,N_14311,N_12084);
and UO_38 (O_38,N_12479,N_14510);
and UO_39 (O_39,N_12641,N_13143);
and UO_40 (O_40,N_12585,N_14018);
nand UO_41 (O_41,N_14858,N_13247);
and UO_42 (O_42,N_14074,N_12869);
nand UO_43 (O_43,N_12978,N_12122);
or UO_44 (O_44,N_13510,N_12621);
nor UO_45 (O_45,N_14085,N_13122);
nand UO_46 (O_46,N_12325,N_14124);
nor UO_47 (O_47,N_14064,N_13827);
nor UO_48 (O_48,N_14785,N_12655);
or UO_49 (O_49,N_13436,N_13473);
or UO_50 (O_50,N_14863,N_12517);
xor UO_51 (O_51,N_13045,N_14754);
nor UO_52 (O_52,N_13536,N_13294);
and UO_53 (O_53,N_14881,N_12312);
xor UO_54 (O_54,N_13272,N_13113);
nand UO_55 (O_55,N_14360,N_12670);
nand UO_56 (O_56,N_12624,N_14448);
nand UO_57 (O_57,N_13582,N_13521);
or UO_58 (O_58,N_12996,N_12572);
and UO_59 (O_59,N_14674,N_13564);
nand UO_60 (O_60,N_13435,N_14026);
or UO_61 (O_61,N_12509,N_14921);
and UO_62 (O_62,N_12197,N_12347);
or UO_63 (O_63,N_12899,N_12456);
and UO_64 (O_64,N_14182,N_13328);
or UO_65 (O_65,N_14913,N_13591);
or UO_66 (O_66,N_14811,N_14418);
xnor UO_67 (O_67,N_13831,N_14277);
nor UO_68 (O_68,N_13710,N_14832);
xor UO_69 (O_69,N_12870,N_13112);
nor UO_70 (O_70,N_13634,N_12535);
xor UO_71 (O_71,N_13263,N_13335);
or UO_72 (O_72,N_13352,N_13982);
nand UO_73 (O_73,N_14550,N_12969);
nor UO_74 (O_74,N_12098,N_12950);
and UO_75 (O_75,N_13911,N_14211);
xor UO_76 (O_76,N_12276,N_13088);
nor UO_77 (O_77,N_14159,N_12880);
xnor UO_78 (O_78,N_12466,N_14643);
nand UO_79 (O_79,N_14254,N_13141);
xor UO_80 (O_80,N_12571,N_14583);
nand UO_81 (O_81,N_13420,N_13882);
nor UO_82 (O_82,N_13223,N_14039);
nand UO_83 (O_83,N_13943,N_14970);
or UO_84 (O_84,N_12733,N_13958);
and UO_85 (O_85,N_14736,N_13781);
xnor UO_86 (O_86,N_14669,N_12752);
xnor UO_87 (O_87,N_12858,N_14053);
nand UO_88 (O_88,N_12699,N_12687);
and UO_89 (O_89,N_14500,N_14817);
nand UO_90 (O_90,N_12223,N_12949);
xnor UO_91 (O_91,N_14642,N_14685);
nor UO_92 (O_92,N_12926,N_13687);
and UO_93 (O_93,N_13361,N_12669);
nor UO_94 (O_94,N_13327,N_14816);
or UO_95 (O_95,N_12280,N_12512);
xnor UO_96 (O_96,N_12121,N_14305);
nand UO_97 (O_97,N_13688,N_13397);
or UO_98 (O_98,N_13762,N_13383);
and UO_99 (O_99,N_14364,N_13891);
xor UO_100 (O_100,N_13594,N_12593);
or UO_101 (O_101,N_14869,N_12545);
nor UO_102 (O_102,N_12021,N_14025);
nand UO_103 (O_103,N_13254,N_13469);
nand UO_104 (O_104,N_14173,N_13496);
nand UO_105 (O_105,N_13029,N_14788);
or UO_106 (O_106,N_12672,N_12897);
or UO_107 (O_107,N_14363,N_12118);
nor UO_108 (O_108,N_14378,N_12567);
xor UO_109 (O_109,N_12662,N_12795);
and UO_110 (O_110,N_14399,N_14387);
and UO_111 (O_111,N_14215,N_14283);
nor UO_112 (O_112,N_13990,N_12731);
nand UO_113 (O_113,N_12070,N_14814);
xnor UO_114 (O_114,N_14361,N_14796);
xor UO_115 (O_115,N_14222,N_12860);
or UO_116 (O_116,N_12493,N_14797);
nor UO_117 (O_117,N_12413,N_14966);
nand UO_118 (O_118,N_12754,N_14955);
nand UO_119 (O_119,N_13561,N_14640);
nand UO_120 (O_120,N_12316,N_12363);
xnor UO_121 (O_121,N_14326,N_14310);
nor UO_122 (O_122,N_13007,N_13506);
or UO_123 (O_123,N_12382,N_13037);
nand UO_124 (O_124,N_14812,N_13818);
nand UO_125 (O_125,N_14650,N_12263);
or UO_126 (O_126,N_12577,N_14009);
nor UO_127 (O_127,N_12994,N_13315);
nor UO_128 (O_128,N_13150,N_14868);
and UO_129 (O_129,N_14795,N_12849);
or UO_130 (O_130,N_12677,N_14261);
nand UO_131 (O_131,N_13250,N_12380);
xnor UO_132 (O_132,N_13387,N_12295);
nor UO_133 (O_133,N_12887,N_14116);
and UO_134 (O_134,N_13476,N_12195);
nand UO_135 (O_135,N_13136,N_12269);
xor UO_136 (O_136,N_13030,N_13746);
xor UO_137 (O_137,N_12477,N_13282);
xnor UO_138 (O_138,N_13894,N_12022);
nand UO_139 (O_139,N_13376,N_14939);
or UO_140 (O_140,N_12081,N_14257);
xor UO_141 (O_141,N_14647,N_12824);
xnor UO_142 (O_142,N_14931,N_12893);
nor UO_143 (O_143,N_12088,N_13042);
nor UO_144 (O_144,N_12813,N_12551);
xor UO_145 (O_145,N_12163,N_13458);
and UO_146 (O_146,N_13440,N_12037);
nor UO_147 (O_147,N_14096,N_13760);
and UO_148 (O_148,N_13185,N_14901);
nand UO_149 (O_149,N_13468,N_14601);
nand UO_150 (O_150,N_14376,N_12013);
and UO_151 (O_151,N_14433,N_14350);
or UO_152 (O_152,N_14415,N_12698);
and UO_153 (O_153,N_12108,N_13711);
nor UO_154 (O_154,N_12473,N_12270);
and UO_155 (O_155,N_14329,N_12211);
or UO_156 (O_156,N_14295,N_14850);
or UO_157 (O_157,N_12123,N_12898);
and UO_158 (O_158,N_13679,N_13124);
nor UO_159 (O_159,N_14089,N_13805);
xnor UO_160 (O_160,N_14136,N_13200);
nand UO_161 (O_161,N_13585,N_12913);
nor UO_162 (O_162,N_12562,N_13332);
nor UO_163 (O_163,N_12071,N_12638);
nor UO_164 (O_164,N_14620,N_13618);
nand UO_165 (O_165,N_12649,N_14791);
nor UO_166 (O_166,N_13871,N_14828);
or UO_167 (O_167,N_13900,N_12207);
xnor UO_168 (O_168,N_13381,N_14829);
nand UO_169 (O_169,N_14147,N_14823);
nor UO_170 (O_170,N_12632,N_13946);
nand UO_171 (O_171,N_13055,N_14611);
nor UO_172 (O_172,N_13962,N_14593);
nand UO_173 (O_173,N_14174,N_13301);
nor UO_174 (O_174,N_13887,N_14956);
xnor UO_175 (O_175,N_13812,N_12847);
nand UO_176 (O_176,N_13434,N_14489);
or UO_177 (O_177,N_14113,N_14200);
nor UO_178 (O_178,N_14659,N_12251);
xnor UO_179 (O_179,N_14373,N_14558);
nor UO_180 (O_180,N_13096,N_13861);
or UO_181 (O_181,N_12410,N_12900);
nor UO_182 (O_182,N_12254,N_14896);
or UO_183 (O_183,N_14265,N_13388);
nor UO_184 (O_184,N_12620,N_13241);
nand UO_185 (O_185,N_12387,N_12155);
or UO_186 (O_186,N_14471,N_14293);
nor UO_187 (O_187,N_13716,N_14288);
nor UO_188 (O_188,N_12963,N_13296);
nor UO_189 (O_189,N_12566,N_14019);
and UO_190 (O_190,N_14815,N_13104);
nand UO_191 (O_191,N_13409,N_13437);
and UO_192 (O_192,N_13953,N_12379);
or UO_193 (O_193,N_13896,N_14485);
nand UO_194 (O_194,N_13592,N_14016);
and UO_195 (O_195,N_12763,N_12922);
and UO_196 (O_196,N_14641,N_14247);
nand UO_197 (O_197,N_13620,N_13876);
nand UO_198 (O_198,N_13913,N_12218);
nand UO_199 (O_199,N_14224,N_12264);
and UO_200 (O_200,N_13061,N_12600);
nand UO_201 (O_201,N_14972,N_12939);
nor UO_202 (O_202,N_14069,N_13835);
nor UO_203 (O_203,N_12667,N_12819);
nand UO_204 (O_204,N_13291,N_14484);
nand UO_205 (O_205,N_12078,N_14272);
xnor UO_206 (O_206,N_14220,N_13641);
xor UO_207 (O_207,N_14285,N_12005);
xor UO_208 (O_208,N_12330,N_12203);
nor UO_209 (O_209,N_14637,N_14527);
and UO_210 (O_210,N_13833,N_13493);
nand UO_211 (O_211,N_12871,N_13954);
nand UO_212 (O_212,N_14690,N_12353);
or UO_213 (O_213,N_13490,N_14045);
nor UO_214 (O_214,N_13685,N_13370);
or UO_215 (O_215,N_14587,N_12769);
xor UO_216 (O_216,N_14662,N_14099);
nand UO_217 (O_217,N_13147,N_14747);
nor UO_218 (O_218,N_12162,N_13923);
and UO_219 (O_219,N_14193,N_12327);
or UO_220 (O_220,N_14666,N_13067);
and UO_221 (O_221,N_12134,N_12156);
or UO_222 (O_222,N_12644,N_12694);
nor UO_223 (O_223,N_13025,N_14712);
nand UO_224 (O_224,N_13248,N_13557);
or UO_225 (O_225,N_14613,N_14857);
nand UO_226 (O_226,N_13249,N_12782);
nor UO_227 (O_227,N_14320,N_12862);
xnor UO_228 (O_228,N_12696,N_14012);
or UO_229 (O_229,N_13416,N_13190);
and UO_230 (O_230,N_12656,N_12755);
or UO_231 (O_231,N_14615,N_14838);
or UO_232 (O_232,N_13682,N_13443);
or UO_233 (O_233,N_13569,N_13960);
nand UO_234 (O_234,N_14556,N_14450);
and UO_235 (O_235,N_13547,N_13759);
and UO_236 (O_236,N_14059,N_13673);
or UO_237 (O_237,N_12359,N_13427);
and UO_238 (O_238,N_13609,N_13163);
and UO_239 (O_239,N_13662,N_12403);
or UO_240 (O_240,N_13714,N_14733);
nand UO_241 (O_241,N_12390,N_12293);
and UO_242 (O_242,N_13854,N_12085);
and UO_243 (O_243,N_12778,N_14525);
and UO_244 (O_244,N_14580,N_12523);
nand UO_245 (O_245,N_13770,N_13087);
and UO_246 (O_246,N_12398,N_13819);
nand UO_247 (O_247,N_12401,N_13503);
xor UO_248 (O_248,N_13334,N_13377);
nor UO_249 (O_249,N_13981,N_14395);
or UO_250 (O_250,N_13286,N_13179);
or UO_251 (O_251,N_12106,N_14887);
or UO_252 (O_252,N_12925,N_12808);
nor UO_253 (O_253,N_12946,N_14893);
and UO_254 (O_254,N_12643,N_13052);
nor UO_255 (O_255,N_12176,N_14919);
and UO_256 (O_256,N_12362,N_14907);
nor UO_257 (O_257,N_14501,N_13463);
and UO_258 (O_258,N_13053,N_12306);
nand UO_259 (O_259,N_14951,N_12318);
and UO_260 (O_260,N_14630,N_14232);
xnor UO_261 (O_261,N_12232,N_13171);
xnor UO_262 (O_262,N_14977,N_14578);
nor UO_263 (O_263,N_14993,N_14176);
and UO_264 (O_264,N_12091,N_14957);
nor UO_265 (O_265,N_12056,N_14109);
and UO_266 (O_266,N_14051,N_13170);
nand UO_267 (O_267,N_12304,N_14511);
and UO_268 (O_268,N_12611,N_14047);
xnor UO_269 (O_269,N_14199,N_12958);
nor UO_270 (O_270,N_13130,N_12484);
nor UO_271 (O_271,N_12388,N_13489);
nand UO_272 (O_272,N_13173,N_12743);
xnor UO_273 (O_273,N_13169,N_13151);
nor UO_274 (O_274,N_13850,N_12068);
or UO_275 (O_275,N_14462,N_13584);
or UO_276 (O_276,N_14714,N_14923);
nand UO_277 (O_277,N_12335,N_14149);
xnor UO_278 (O_278,N_14629,N_13367);
nand UO_279 (O_279,N_12874,N_14101);
nand UO_280 (O_280,N_14407,N_13390);
xor UO_281 (O_281,N_12031,N_14513);
xor UO_282 (O_282,N_13756,N_14746);
and UO_283 (O_283,N_12099,N_12936);
and UO_284 (O_284,N_14398,N_12185);
and UO_285 (O_285,N_12625,N_13018);
and UO_286 (O_286,N_12674,N_14563);
nor UO_287 (O_287,N_13863,N_12771);
and UO_288 (O_288,N_13043,N_13629);
and UO_289 (O_289,N_14600,N_12038);
nor UO_290 (O_290,N_12829,N_13659);
and UO_291 (O_291,N_13708,N_13253);
or UO_292 (O_292,N_12538,N_14958);
or UO_293 (O_293,N_13127,N_13230);
and UO_294 (O_294,N_13941,N_14655);
nand UO_295 (O_295,N_14313,N_12934);
nand UO_296 (O_296,N_12463,N_14474);
and UO_297 (O_297,N_12710,N_14262);
nand UO_298 (O_298,N_14434,N_13168);
nand UO_299 (O_299,N_13874,N_12530);
and UO_300 (O_300,N_12253,N_12711);
nand UO_301 (O_301,N_14726,N_14700);
or UO_302 (O_302,N_14968,N_12882);
and UO_303 (O_303,N_14458,N_14432);
and UO_304 (O_304,N_12987,N_13276);
or UO_305 (O_305,N_13895,N_14400);
nand UO_306 (O_306,N_13792,N_13661);
nor UO_307 (O_307,N_14306,N_12370);
nand UO_308 (O_308,N_12905,N_13017);
xnor UO_309 (O_309,N_13520,N_12331);
nor UO_310 (O_310,N_12273,N_13353);
xnor UO_311 (O_311,N_13350,N_13695);
xor UO_312 (O_312,N_12149,N_12384);
and UO_313 (O_313,N_14619,N_14379);
or UO_314 (O_314,N_14005,N_12083);
and UO_315 (O_315,N_14806,N_14155);
and UO_316 (O_316,N_12794,N_13146);
and UO_317 (O_317,N_13359,N_14229);
xor UO_318 (O_318,N_12527,N_13743);
nor UO_319 (O_319,N_12651,N_14594);
nand UO_320 (O_320,N_14386,N_13529);
nor UO_321 (O_321,N_12127,N_14710);
xor UO_322 (O_322,N_12957,N_13191);
or UO_323 (O_323,N_12394,N_12903);
and UO_324 (O_324,N_14312,N_14606);
xnor UO_325 (O_325,N_14539,N_14624);
and UO_326 (O_326,N_12909,N_14779);
or UO_327 (O_327,N_13065,N_14266);
and UO_328 (O_328,N_12198,N_14145);
nand UO_329 (O_329,N_13464,N_13100);
and UO_330 (O_330,N_14661,N_13729);
nor UO_331 (O_331,N_13016,N_14031);
or UO_332 (O_332,N_13046,N_12877);
xnor UO_333 (O_333,N_14927,N_12736);
nor UO_334 (O_334,N_14468,N_12361);
nor UO_335 (O_335,N_14275,N_14591);
or UO_336 (O_336,N_14935,N_14340);
xor UO_337 (O_337,N_13578,N_13974);
xor UO_338 (O_338,N_13800,N_13289);
xor UO_339 (O_339,N_13131,N_14439);
nor UO_340 (O_340,N_13844,N_14052);
or UO_341 (O_341,N_14499,N_13862);
or UO_342 (O_342,N_12317,N_13864);
nand UO_343 (O_343,N_13648,N_14227);
nor UO_344 (O_344,N_14372,N_12832);
and UO_345 (O_345,N_14093,N_14212);
and UO_346 (O_346,N_14472,N_12563);
nand UO_347 (O_347,N_13931,N_12690);
nand UO_348 (O_348,N_12402,N_12648);
xnor UO_349 (O_349,N_13393,N_13166);
nor UO_350 (O_350,N_14689,N_13624);
xor UO_351 (O_351,N_13134,N_13456);
and UO_352 (O_352,N_14435,N_13914);
or UO_353 (O_353,N_13319,N_13363);
and UO_354 (O_354,N_12100,N_14820);
or UO_355 (O_355,N_13870,N_14160);
or UO_356 (O_356,N_14307,N_14880);
nand UO_357 (O_357,N_12543,N_14554);
and UO_358 (O_358,N_14354,N_13019);
or UO_359 (O_359,N_14571,N_13300);
and UO_360 (O_360,N_14783,N_12400);
nand UO_361 (O_361,N_14382,N_12916);
nor UO_362 (O_362,N_14548,N_13765);
or UO_363 (O_363,N_12702,N_13174);
nor UO_364 (O_364,N_13322,N_13978);
nor UO_365 (O_365,N_13977,N_14559);
and UO_366 (O_366,N_13331,N_14068);
nand UO_367 (O_367,N_14741,N_12975);
and UO_368 (O_368,N_14759,N_13998);
nor UO_369 (O_369,N_12442,N_12773);
or UO_370 (O_370,N_14339,N_13995);
nor UO_371 (O_371,N_13677,N_13654);
nand UO_372 (O_372,N_13445,N_13604);
or UO_373 (O_373,N_12745,N_13745);
xnor UO_374 (O_374,N_13806,N_14738);
xnor UO_375 (O_375,N_13049,N_13848);
and UO_376 (O_376,N_13769,N_13701);
nor UO_377 (O_377,N_13078,N_12681);
nor UO_378 (O_378,N_13347,N_12820);
or UO_379 (O_379,N_14083,N_13777);
xor UO_380 (O_380,N_14153,N_13533);
nor UO_381 (O_381,N_13114,N_13371);
xnor UO_382 (O_382,N_12812,N_13238);
nor UO_383 (O_383,N_13178,N_13587);
or UO_384 (O_384,N_14327,N_14426);
nand UO_385 (O_385,N_12580,N_14917);
nor UO_386 (O_386,N_14646,N_14065);
or UO_387 (O_387,N_13738,N_12292);
or UO_388 (O_388,N_12894,N_13545);
or UO_389 (O_389,N_14357,N_12979);
and UO_390 (O_390,N_14055,N_13050);
and UO_391 (O_391,N_14050,N_14032);
xor UO_392 (O_392,N_13369,N_12455);
nand UO_393 (O_393,N_13852,N_14317);
and UO_394 (O_394,N_12878,N_14091);
and UO_395 (O_395,N_14625,N_12406);
nand UO_396 (O_396,N_13878,N_12302);
nand UO_397 (O_397,N_12586,N_12855);
or UO_398 (O_398,N_12504,N_12219);
or UO_399 (O_399,N_13015,N_14508);
xnor UO_400 (O_400,N_13040,N_13080);
xnor UO_401 (O_401,N_14902,N_12428);
nor UO_402 (O_402,N_14290,N_12646);
nand UO_403 (O_403,N_14808,N_12998);
xnor UO_404 (O_404,N_13531,N_14839);
xnor UO_405 (O_405,N_13951,N_13284);
nor UO_406 (O_406,N_13077,N_13822);
nor UO_407 (O_407,N_12415,N_13023);
nor UO_408 (O_408,N_13188,N_14813);
nand UO_409 (O_409,N_12461,N_12294);
or UO_410 (O_410,N_12320,N_14589);
and UO_411 (O_411,N_14067,N_13672);
and UO_412 (O_412,N_13089,N_13556);
or UO_413 (O_413,N_12434,N_13773);
nand UO_414 (O_414,N_13345,N_14263);
or UO_415 (O_415,N_12089,N_14592);
nor UO_416 (O_416,N_13081,N_14599);
nor UO_417 (O_417,N_13622,N_12706);
nand UO_418 (O_418,N_12004,N_13889);
or UO_419 (O_419,N_12329,N_13712);
xnor UO_420 (O_420,N_14236,N_13724);
xor UO_421 (O_421,N_14216,N_14139);
xor UO_422 (O_422,N_14429,N_14430);
nor UO_423 (O_423,N_13605,N_12896);
nand UO_424 (O_424,N_14800,N_12212);
nor UO_425 (O_425,N_12953,N_13267);
and UO_426 (O_426,N_12827,N_14664);
nor UO_427 (O_427,N_12407,N_13907);
nor UO_428 (O_428,N_13802,N_12497);
nor UO_429 (O_429,N_13430,N_13326);
xor UO_430 (O_430,N_13501,N_13948);
xnor UO_431 (O_431,N_13926,N_14774);
or UO_432 (O_432,N_12345,N_12045);
xor UO_433 (O_433,N_13843,N_14191);
or UO_434 (O_434,N_12006,N_13433);
nand UO_435 (O_435,N_14447,N_14014);
nand UO_436 (O_436,N_14362,N_14937);
nand UO_437 (O_437,N_12450,N_12568);
or UO_438 (O_438,N_13704,N_12971);
and UO_439 (O_439,N_12346,N_14803);
and UO_440 (O_440,N_13379,N_14870);
or UO_441 (O_441,N_13796,N_14308);
xor UO_442 (O_442,N_14115,N_12046);
xnor UO_443 (O_443,N_14549,N_13094);
or UO_444 (O_444,N_12607,N_12810);
nand UO_445 (O_445,N_13474,N_12749);
and UO_446 (O_446,N_14490,N_12366);
nor UO_447 (O_447,N_14302,N_14208);
nor UO_448 (O_448,N_14322,N_14297);
and UO_449 (O_449,N_13608,N_14449);
or UO_450 (O_450,N_12742,N_14171);
xor UO_451 (O_451,N_12741,N_13680);
and UO_452 (O_452,N_14924,N_14517);
and UO_453 (O_453,N_12385,N_12116);
xor UO_454 (O_454,N_12404,N_14848);
and UO_455 (O_455,N_12853,N_12377);
nor UO_456 (O_456,N_12866,N_13924);
nand UO_457 (O_457,N_12396,N_12510);
nor UO_458 (O_458,N_13942,N_13535);
nor UO_459 (O_459,N_13159,N_13244);
or UO_460 (O_460,N_14244,N_12480);
nand UO_461 (O_461,N_14456,N_12623);
or UO_462 (O_462,N_12471,N_12865);
nor UO_463 (O_463,N_12034,N_13444);
nor UO_464 (O_464,N_14760,N_14201);
nand UO_465 (O_465,N_12222,N_13935);
or UO_466 (O_466,N_13817,N_14932);
xor UO_467 (O_467,N_12933,N_13853);
and UO_468 (O_468,N_14156,N_12774);
nor UO_469 (O_469,N_13071,N_13259);
or UO_470 (O_470,N_12019,N_13588);
nand UO_471 (O_471,N_12823,N_13349);
and UO_472 (O_472,N_12094,N_13856);
and UO_473 (O_473,N_14634,N_13203);
and UO_474 (O_474,N_13062,N_14598);
and UO_475 (O_475,N_14878,N_14041);
and UO_476 (O_476,N_13985,N_12920);
xor UO_477 (O_477,N_12322,N_13145);
xnor UO_478 (O_478,N_12628,N_14343);
nor UO_479 (O_479,N_14509,N_12160);
nand UO_480 (O_480,N_14826,N_12015);
or UO_481 (O_481,N_12053,N_13339);
xor UO_482 (O_482,N_12230,N_12392);
nor UO_483 (O_483,N_14790,N_14677);
nor UO_484 (O_484,N_12546,N_14390);
or UO_485 (O_485,N_12895,N_12744);
nor UO_486 (O_486,N_13499,N_14365);
or UO_487 (O_487,N_13403,N_13251);
xor UO_488 (O_488,N_12337,N_13857);
nand UO_489 (O_489,N_13246,N_12757);
nand UO_490 (O_490,N_14004,N_12086);
or UO_491 (O_491,N_12817,N_12947);
xor UO_492 (O_492,N_14309,N_14369);
and UO_493 (O_493,N_13297,N_13727);
and UO_494 (O_494,N_14202,N_14192);
or UO_495 (O_495,N_14328,N_13512);
nand UO_496 (O_496,N_14737,N_14573);
nand UO_497 (O_497,N_12305,N_14006);
and UO_498 (O_498,N_12368,N_12489);
nand UO_499 (O_499,N_13775,N_14358);
nor UO_500 (O_500,N_12117,N_14488);
nor UO_501 (O_501,N_14008,N_13553);
or UO_502 (O_502,N_14515,N_12940);
or UO_503 (O_503,N_13142,N_14960);
nand UO_504 (O_504,N_12734,N_12863);
nand UO_505 (O_505,N_12216,N_14179);
nor UO_506 (O_506,N_14952,N_12918);
or UO_507 (O_507,N_14844,N_12311);
xor UO_508 (O_508,N_14930,N_14221);
nand UO_509 (O_509,N_12770,N_13082);
and UO_510 (O_510,N_14445,N_13269);
and UO_511 (O_511,N_13664,N_12992);
nor UO_512 (O_512,N_14757,N_12581);
or UO_513 (O_513,N_12919,N_12713);
nand UO_514 (O_514,N_14457,N_12668);
nand UO_515 (O_515,N_12814,N_14794);
and UO_516 (O_516,N_13959,N_13005);
nand UO_517 (O_517,N_13354,N_14516);
xnor UO_518 (O_518,N_13139,N_14775);
xnor UO_519 (O_519,N_14321,N_13616);
and UO_520 (O_520,N_12889,N_14505);
and UO_521 (O_521,N_13274,N_14729);
nor UO_522 (O_522,N_13262,N_12147);
nor UO_523 (O_523,N_12289,N_13175);
or UO_524 (O_524,N_14648,N_13973);
and UO_525 (O_525,N_14483,N_14167);
and UO_526 (O_526,N_14180,N_12186);
xnor UO_527 (O_527,N_13366,N_12412);
or UO_528 (O_528,N_12355,N_14146);
and UO_529 (O_529,N_12879,N_12451);
or UO_530 (O_530,N_14393,N_14999);
nand UO_531 (O_531,N_13351,N_13164);
xnor UO_532 (O_532,N_12448,N_12884);
xor UO_533 (O_533,N_14217,N_12024);
and UO_534 (O_534,N_12389,N_12737);
and UO_535 (O_535,N_13195,N_14873);
xnor UO_536 (O_536,N_13449,N_14036);
nor UO_537 (O_537,N_12608,N_14731);
or UO_538 (O_538,N_14906,N_12338);
xor UO_539 (O_539,N_12221,N_12796);
nand UO_540 (O_540,N_14278,N_12470);
nand UO_541 (O_541,N_13859,N_13807);
and UO_542 (O_542,N_14131,N_12454);
xnor UO_543 (O_543,N_12277,N_12682);
and UO_544 (O_544,N_14503,N_13111);
or UO_545 (O_545,N_12257,N_14140);
xnor UO_546 (O_546,N_14520,N_13517);
and UO_547 (O_547,N_12172,N_12906);
and UO_548 (O_548,N_13543,N_14046);
nor UO_549 (O_549,N_14259,N_14344);
nand UO_550 (O_550,N_14123,N_14479);
and UO_551 (O_551,N_13070,N_12260);
or UO_552 (O_552,N_12891,N_12023);
and UO_553 (O_553,N_14964,N_12844);
or UO_554 (O_554,N_13754,N_14020);
and UO_555 (O_555,N_13971,N_13993);
and UO_556 (O_556,N_14767,N_13903);
and UO_557 (O_557,N_12910,N_14521);
nor UO_558 (O_558,N_14121,N_12067);
xor UO_559 (O_559,N_12788,N_12640);
nand UO_560 (O_560,N_12447,N_13364);
nand UO_561 (O_561,N_14645,N_13218);
nor UO_562 (O_562,N_12615,N_14735);
nor UO_563 (O_563,N_12962,N_13001);
and UO_564 (O_564,N_14532,N_12740);
or UO_565 (O_565,N_12190,N_14094);
and UO_566 (O_566,N_13893,N_13890);
or UO_567 (O_567,N_13683,N_12409);
xnor UO_568 (O_568,N_12433,N_13140);
nand UO_569 (O_569,N_14177,N_12595);
or UO_570 (O_570,N_13283,N_12164);
nand UO_571 (O_571,N_14144,N_12187);
or UO_572 (O_572,N_14506,N_12188);
and UO_573 (O_573,N_14551,N_13108);
nand UO_574 (O_574,N_14453,N_13830);
and UO_575 (O_575,N_13929,N_14953);
or UO_576 (O_576,N_12016,N_14092);
xor UO_577 (O_577,N_12807,N_14577);
xor UO_578 (O_578,N_12914,N_12775);
nor UO_579 (O_579,N_12777,N_14013);
nor UO_580 (O_580,N_14428,N_14205);
or UO_581 (O_581,N_13524,N_14492);
nor UO_582 (O_582,N_12242,N_13758);
nand UO_583 (O_583,N_14112,N_12730);
nand UO_584 (O_584,N_14420,N_13908);
nor UO_585 (O_585,N_14536,N_14560);
xnor UO_586 (O_586,N_13235,N_14477);
and UO_587 (O_587,N_13205,N_13177);
nand UO_588 (O_588,N_14704,N_12797);
and UO_589 (O_589,N_13385,N_13194);
or UO_590 (O_590,N_14294,N_12852);
and UO_591 (O_591,N_13079,N_12281);
nand UO_592 (O_592,N_13619,N_14671);
xor UO_593 (O_593,N_13401,N_13133);
nor UO_594 (O_594,N_12309,N_14565);
nand UO_595 (O_595,N_13744,N_13580);
and UO_596 (O_596,N_12059,N_14895);
nand UO_597 (O_597,N_12705,N_13404);
or UO_598 (O_598,N_13788,N_12453);
and UO_599 (O_599,N_13736,N_12103);
nand UO_600 (O_600,N_13811,N_14256);
and UO_601 (O_601,N_14676,N_13980);
or UO_602 (O_602,N_14657,N_14246);
nor UO_603 (O_603,N_12839,N_12806);
nand UO_604 (O_604,N_14126,N_13638);
and UO_605 (O_605,N_13405,N_13470);
nand UO_606 (O_606,N_14524,N_12042);
nor UO_607 (O_607,N_13928,N_12252);
xor UO_608 (O_608,N_12184,N_14849);
xnor UO_609 (O_609,N_13273,N_13541);
and UO_610 (O_610,N_12986,N_12178);
nor UO_611 (O_611,N_12431,N_12675);
and UO_612 (O_612,N_14002,N_14150);
and UO_613 (O_613,N_14250,N_12590);
or UO_614 (O_614,N_13917,N_13657);
and UO_615 (O_615,N_13920,N_14504);
and UO_616 (O_616,N_14531,N_14172);
nand UO_617 (O_617,N_12718,N_14730);
nand UO_618 (O_618,N_13355,N_12169);
nor UO_619 (O_619,N_14495,N_12429);
nand UO_620 (O_620,N_13697,N_13157);
nor UO_621 (O_621,N_14132,N_12018);
or UO_622 (O_622,N_14860,N_13495);
or UO_623 (O_623,N_12114,N_14441);
and UO_624 (O_624,N_13441,N_13158);
or UO_625 (O_625,N_13829,N_13105);
or UO_626 (O_626,N_12912,N_13181);
nand UO_627 (O_627,N_12000,N_13337);
nor UO_628 (O_628,N_14693,N_14455);
nand UO_629 (O_629,N_13232,N_12700);
or UO_630 (O_630,N_13939,N_13934);
nand UO_631 (O_631,N_12724,N_13497);
nor UO_632 (O_632,N_14552,N_12102);
xor UO_633 (O_633,N_13949,N_12220);
xnor UO_634 (O_634,N_12443,N_14076);
and UO_635 (O_635,N_14612,N_12202);
and UO_636 (O_636,N_13610,N_13500);
and UO_637 (O_637,N_14522,N_14110);
or UO_638 (O_638,N_14128,N_12684);
or UO_639 (O_639,N_13766,N_14185);
or UO_640 (O_640,N_12119,N_12556);
or UO_641 (O_641,N_12805,N_12139);
or UO_642 (O_642,N_13115,N_12514);
nand UO_643 (O_643,N_12151,N_12427);
or UO_644 (O_644,N_12676,N_14804);
or UO_645 (O_645,N_13309,N_13965);
nand UO_646 (O_646,N_14405,N_12165);
or UO_647 (O_647,N_13026,N_14494);
nor UO_648 (O_648,N_12107,N_14946);
or UO_649 (O_649,N_12490,N_12857);
or UO_650 (O_650,N_14748,N_14789);
and UO_651 (O_651,N_13694,N_14000);
or UO_652 (O_652,N_13637,N_13398);
nand UO_653 (O_653,N_12007,N_13975);
xnor UO_654 (O_654,N_14077,N_13008);
xnor UO_655 (O_655,N_13271,N_13325);
or UO_656 (O_656,N_12339,N_13905);
nor UO_657 (O_657,N_13233,N_14151);
xor UO_658 (O_658,N_12228,N_12043);
nor UO_659 (O_659,N_14702,N_12653);
and UO_660 (O_660,N_13129,N_14292);
nor UO_661 (O_661,N_14518,N_13461);
nand UO_662 (O_662,N_14756,N_12395);
nor UO_663 (O_663,N_12137,N_14686);
and UO_664 (O_664,N_14928,N_14978);
nor UO_665 (O_665,N_13285,N_13667);
nor UO_666 (O_666,N_14837,N_12618);
or UO_667 (O_667,N_14740,N_12082);
nand UO_668 (O_668,N_12319,N_12374);
and UO_669 (O_669,N_13860,N_13183);
or UO_670 (O_670,N_14375,N_14443);
xnor UO_671 (O_671,N_13020,N_14567);
nor UO_672 (O_672,N_12739,N_12050);
xor UO_673 (O_673,N_13450,N_14581);
or UO_674 (O_674,N_13035,N_12367);
or UO_675 (O_675,N_13313,N_14371);
and UO_676 (O_676,N_12565,N_13459);
xor UO_677 (O_677,N_13627,N_13795);
and UO_678 (O_678,N_14988,N_13261);
nor UO_679 (O_679,N_12354,N_12719);
nor UO_680 (O_680,N_13036,N_14707);
xor UO_681 (O_681,N_14421,N_13783);
nor UO_682 (O_682,N_14568,N_14476);
nor UO_683 (O_683,N_13421,N_12574);
nor UO_684 (O_684,N_12491,N_14705);
or UO_685 (O_685,N_14761,N_13632);
nand UO_686 (O_686,N_12111,N_14926);
nand UO_687 (O_687,N_13155,N_14905);
nor UO_688 (O_688,N_13323,N_13375);
nand UO_689 (O_689,N_14540,N_12011);
nor UO_690 (O_690,N_13607,N_13032);
nor UO_691 (O_691,N_14900,N_14995);
xor UO_692 (O_692,N_12846,N_14776);
and UO_693 (O_693,N_13663,N_14138);
xor UO_694 (O_694,N_14157,N_13838);
nand UO_695 (O_695,N_14348,N_12032);
xnor UO_696 (O_696,N_13571,N_14985);
xnor UO_697 (O_697,N_12483,N_12033);
or UO_698 (O_698,N_12457,N_14586);
nor UO_699 (O_699,N_12995,N_14243);
nor UO_700 (O_700,N_14537,N_12665);
nand UO_701 (O_701,N_12352,N_12143);
xnor UO_702 (O_702,N_13338,N_14879);
xor UO_703 (O_703,N_13540,N_13215);
xor UO_704 (O_704,N_13333,N_14538);
and UO_705 (O_705,N_13198,N_12553);
nor UO_706 (O_706,N_13565,N_13197);
or UO_707 (O_707,N_12635,N_14561);
nor UO_708 (O_708,N_14385,N_13002);
nor UO_709 (O_709,N_12109,N_13647);
or UO_710 (O_710,N_13799,N_14097);
nor UO_711 (O_711,N_13462,N_12326);
nand UO_712 (O_712,N_14684,N_12161);
nand UO_713 (O_713,N_14024,N_12296);
nand UO_714 (O_714,N_14332,N_13731);
nand UO_715 (O_715,N_14394,N_12980);
xor UO_716 (O_716,N_12183,N_12399);
nor UO_717 (O_717,N_13563,N_14884);
nand UO_718 (O_718,N_14912,N_12942);
and UO_719 (O_719,N_13872,N_14342);
or UO_720 (O_720,N_12179,N_13658);
or UO_721 (O_721,N_13613,N_13307);
and UO_722 (O_722,N_12233,N_14125);
and UO_723 (O_723,N_12213,N_13709);
nand UO_724 (O_724,N_13298,N_12378);
nand UO_725 (O_725,N_12153,N_13324);
or UO_726 (O_726,N_13528,N_14843);
xor UO_727 (O_727,N_14841,N_13368);
and UO_728 (O_728,N_14431,N_12575);
nand UO_729 (O_729,N_14743,N_12226);
or UO_730 (O_730,N_13722,N_14440);
xnor UO_731 (O_731,N_12652,N_12351);
nor UO_732 (O_732,N_14846,N_14831);
nor UO_733 (O_733,N_13693,N_14284);
and UO_734 (O_734,N_13028,N_14341);
nor UO_735 (O_735,N_14467,N_12616);
and UO_736 (O_736,N_12685,N_13389);
or UO_737 (O_737,N_12087,N_12437);
xnor UO_738 (O_738,N_13210,N_12129);
or UO_739 (O_739,N_14523,N_14459);
and UO_740 (O_740,N_12418,N_13847);
or UO_741 (O_741,N_13211,N_13242);
or UO_742 (O_742,N_14106,N_12124);
and UO_743 (O_743,N_13419,N_13834);
and UO_744 (O_744,N_13602,N_12073);
or UO_745 (O_745,N_13356,N_12854);
or UO_746 (O_746,N_13208,N_12915);
nor UO_747 (O_747,N_12265,N_13551);
xor UO_748 (O_748,N_12041,N_12609);
nand UO_749 (O_749,N_14715,N_12521);
xnor UO_750 (O_750,N_12845,N_14230);
nand UO_751 (O_751,N_13522,N_12475);
or UO_752 (O_752,N_12194,N_13066);
nor UO_753 (O_753,N_13794,N_14658);
and UO_754 (O_754,N_12341,N_12416);
and UO_755 (O_755,N_14381,N_12052);
xor UO_756 (O_756,N_12629,N_14722);
xor UO_757 (O_757,N_14904,N_12709);
or UO_758 (O_758,N_12792,N_13428);
and UO_759 (O_759,N_12592,N_14493);
and UO_760 (O_760,N_14725,N_14080);
and UO_761 (O_761,N_13446,N_12815);
nor UO_762 (O_762,N_14396,N_14732);
and UO_763 (O_763,N_14916,N_14920);
and UO_764 (O_764,N_14652,N_12501);
and UO_765 (O_765,N_12044,N_14135);
and UO_766 (O_766,N_13581,N_14940);
nand UO_767 (O_767,N_14534,N_12334);
or UO_768 (O_768,N_13086,N_13986);
nor UO_769 (O_769,N_13635,N_14401);
xnor UO_770 (O_770,N_12240,N_12984);
xnor UO_771 (O_771,N_13888,N_12627);
or UO_772 (O_772,N_14209,N_13280);
and UO_773 (O_773,N_14660,N_14979);
nor UO_774 (O_774,N_14679,N_14347);
or UO_775 (O_775,N_14228,N_12229);
or UO_776 (O_776,N_14784,N_14541);
xnor UO_777 (O_777,N_14351,N_14681);
or UO_778 (O_778,N_12508,N_14810);
xor UO_779 (O_779,N_13382,N_14104);
and UO_780 (O_780,N_14451,N_14442);
or UO_781 (O_781,N_14108,N_12182);
and UO_782 (O_782,N_13733,N_13696);
and UO_783 (O_783,N_12459,N_14406);
xor UO_784 (O_784,N_12868,N_13523);
xnor UO_785 (O_785,N_13400,N_13858);
nand UO_786 (O_786,N_12142,N_13786);
and UO_787 (O_787,N_13636,N_14425);
nand UO_788 (O_788,N_12029,N_13292);
xnor UO_789 (O_789,N_13418,N_14496);
xnor UO_790 (O_790,N_13034,N_14663);
or UO_791 (O_791,N_14316,N_14129);
and UO_792 (O_792,N_12816,N_12313);
xnor UO_793 (O_793,N_12066,N_12283);
xor UO_794 (O_794,N_12558,N_14750);
nand UO_795 (O_795,N_12908,N_13555);
xor UO_796 (O_796,N_13961,N_12074);
xor UO_797 (O_797,N_13655,N_14245);
nand UO_798 (O_798,N_12606,N_13944);
or UO_799 (O_799,N_13562,N_14214);
or UO_800 (O_800,N_13165,N_14632);
xor UO_801 (O_801,N_12077,N_13279);
xnor UO_802 (O_802,N_14130,N_14219);
and UO_803 (O_803,N_12780,N_12636);
and UO_804 (O_804,N_12717,N_14997);
xnor UO_805 (O_805,N_12487,N_13737);
xnor UO_806 (O_806,N_13793,N_12259);
nor UO_807 (O_807,N_14833,N_14235);
nand UO_808 (O_808,N_14535,N_14994);
or UO_809 (O_809,N_14597,N_12666);
or UO_810 (O_810,N_12373,N_14897);
xor UO_811 (O_811,N_13103,N_12247);
xnor UO_812 (O_812,N_14027,N_12488);
or UO_813 (O_813,N_13996,N_12603);
nand UO_814 (O_814,N_12881,N_13386);
and UO_815 (O_815,N_13423,N_13011);
nand UO_816 (O_816,N_14022,N_12208);
and UO_817 (O_817,N_12661,N_13288);
nor UO_818 (O_818,N_13119,N_14996);
nor UO_819 (O_819,N_14945,N_13988);
or UO_820 (O_820,N_12110,N_12993);
xor UO_821 (O_821,N_12943,N_13646);
nor UO_822 (O_822,N_14871,N_13257);
or UO_823 (O_823,N_13947,N_12697);
and UO_824 (O_824,N_12786,N_12729);
nand UO_825 (O_825,N_12917,N_13154);
or UO_826 (O_826,N_13652,N_13161);
or UO_827 (O_827,N_12626,N_12708);
and UO_828 (O_828,N_13399,N_13176);
xor UO_829 (O_829,N_14218,N_14040);
or UO_830 (O_830,N_12650,N_14922);
nand UO_831 (O_831,N_13910,N_13256);
or UO_832 (O_832,N_12132,N_12113);
or UO_833 (O_833,N_12851,N_14918);
xnor UO_834 (O_834,N_13348,N_13358);
nand UO_835 (O_835,N_13832,N_14992);
nor UO_836 (O_836,N_14673,N_14618);
nand UO_837 (O_837,N_13644,N_12452);
or UO_838 (O_838,N_13560,N_13192);
xnor UO_839 (O_839,N_12234,N_12405);
nor UO_840 (O_840,N_12826,N_13748);
xnor UO_841 (O_841,N_12133,N_13810);
and UO_842 (O_842,N_12972,N_14948);
and UO_843 (O_843,N_13207,N_14475);
nand UO_844 (O_844,N_14954,N_13937);
or UO_845 (O_845,N_14621,N_13590);
and UO_846 (O_846,N_13921,N_14909);
nand UO_847 (O_847,N_12010,N_14148);
nand UO_848 (O_848,N_12039,N_13243);
nor UO_849 (O_849,N_12344,N_12536);
xnor UO_850 (O_850,N_12075,N_14260);
or UO_851 (O_851,N_14595,N_14454);
and UO_852 (O_852,N_12602,N_14933);
or UO_853 (O_853,N_14411,N_13791);
nor UO_854 (O_854,N_12300,N_13918);
or UO_855 (O_855,N_12080,N_12735);
or UO_856 (O_856,N_12673,N_14299);
xnor UO_857 (O_857,N_12028,N_13992);
or UO_858 (O_858,N_13845,N_13537);
nor UO_859 (O_859,N_13483,N_12798);
nand UO_860 (O_860,N_14063,N_13699);
nand UO_861 (O_861,N_13031,N_13717);
or UO_862 (O_862,N_12272,N_14042);
and UO_863 (O_863,N_13009,N_14466);
nor UO_864 (O_864,N_12349,N_13270);
nand UO_865 (O_865,N_13706,N_12474);
xor UO_866 (O_866,N_14910,N_14545);
or UO_867 (O_867,N_13255,N_12476);
nand UO_868 (O_868,N_13095,N_14542);
nor UO_869 (O_869,N_13182,N_13180);
or UO_870 (O_870,N_13278,N_12772);
nand UO_871 (O_871,N_13816,N_12840);
nand UO_872 (O_872,N_12255,N_13940);
or UO_873 (O_873,N_13438,N_12040);
nor UO_874 (O_874,N_13933,N_12904);
nor UO_875 (O_875,N_13670,N_13867);
and UO_876 (O_876,N_14969,N_14649);
or UO_877 (O_877,N_12793,N_14114);
and UO_878 (O_878,N_13252,N_12970);
nand UO_879 (O_879,N_12371,N_12564);
nand UO_880 (O_880,N_12482,N_14336);
and UO_881 (O_881,N_12411,N_13308);
and UO_882 (O_882,N_12977,N_14289);
xnor UO_883 (O_883,N_12321,N_12842);
or UO_884 (O_884,N_12008,N_13076);
or UO_885 (O_885,N_12167,N_13484);
or UO_886 (O_886,N_14037,N_14915);
and UO_887 (O_887,N_13329,N_13314);
and UO_888 (O_888,N_13764,N_13373);
nor UO_889 (O_889,N_14203,N_14936);
nand UO_890 (O_890,N_12486,N_12246);
and UO_891 (O_891,N_14773,N_14487);
and UO_892 (O_892,N_13767,N_13703);
nor UO_893 (O_893,N_12460,N_12584);
xor UO_894 (O_894,N_14352,N_12199);
or UO_895 (O_895,N_14675,N_12695);
or UO_896 (O_896,N_13504,N_14274);
nand UO_897 (O_897,N_12054,N_14603);
xor UO_898 (O_898,N_14934,N_13411);
or UO_899 (O_899,N_14298,N_12168);
nor UO_900 (O_900,N_13426,N_12885);
and UO_901 (O_901,N_13260,N_14654);
xor UO_902 (O_902,N_12764,N_12291);
nand UO_903 (O_903,N_13439,N_12515);
xor UO_904 (O_904,N_12631,N_12057);
xnor UO_905 (O_905,N_12502,N_14060);
or UO_906 (O_906,N_13048,N_14082);
or UO_907 (O_907,N_14117,N_14061);
nand UO_908 (O_908,N_13487,N_13803);
nand UO_909 (O_909,N_14058,N_13774);
nand UO_910 (O_910,N_14692,N_13780);
nand UO_911 (O_911,N_13728,N_12314);
nor UO_912 (O_912,N_14579,N_13128);
or UO_913 (O_913,N_14464,N_14667);
or UO_914 (O_914,N_14607,N_12035);
nand UO_915 (O_915,N_14072,N_14264);
and UO_916 (O_916,N_13884,N_12691);
xor UO_917 (O_917,N_13725,N_14727);
xnor UO_918 (O_918,N_13550,N_12464);
nand UO_919 (O_919,N_13808,N_12598);
xor UO_920 (O_920,N_14672,N_12079);
nand UO_921 (O_921,N_13422,N_14947);
and UO_922 (O_922,N_12583,N_14044);
and UO_923 (O_923,N_14742,N_14778);
or UO_924 (O_924,N_13642,N_12250);
and UO_925 (O_925,N_13801,N_14287);
and UO_926 (O_926,N_12126,N_14822);
or UO_927 (O_927,N_13735,N_12727);
and UO_928 (O_928,N_12128,N_12444);
or UO_929 (O_929,N_13669,N_13771);
nand UO_930 (O_930,N_12225,N_13186);
nor UO_931 (O_931,N_12130,N_13213);
nor UO_932 (O_932,N_13881,N_13950);
or UO_933 (O_933,N_13392,N_14980);
and UO_934 (O_934,N_14751,N_12591);
and UO_935 (O_935,N_12105,N_12932);
nand UO_936 (O_936,N_13721,N_12506);
and UO_937 (O_937,N_13626,N_12555);
xnor UO_938 (O_938,N_12065,N_14391);
nor UO_939 (O_939,N_12243,N_13488);
and UO_940 (O_940,N_13372,N_14184);
xnor UO_941 (O_941,N_14196,N_12966);
nor UO_942 (O_942,N_14355,N_13823);
nand UO_943 (O_943,N_13732,N_13006);
nand UO_944 (O_944,N_13047,N_13478);
and UO_945 (O_945,N_13675,N_13425);
or UO_946 (O_946,N_12907,N_13927);
or UO_947 (O_947,N_14353,N_13290);
nand UO_948 (O_948,N_12758,N_14770);
nand UO_949 (O_949,N_14279,N_12890);
and UO_950 (O_950,N_14809,N_14749);
nor UO_951 (O_951,N_14744,N_14001);
nand UO_952 (O_952,N_12048,N_12249);
nand UO_953 (O_953,N_14889,N_12397);
or UO_954 (O_954,N_13098,N_14368);
and UO_955 (O_955,N_12478,N_12955);
or UO_956 (O_956,N_14528,N_12633);
nor UO_957 (O_957,N_13761,N_13494);
or UO_958 (O_958,N_12520,N_13526);
nand UO_959 (O_959,N_12800,N_12554);
nor UO_960 (O_960,N_14769,N_13668);
and UO_961 (O_961,N_14983,N_12492);
or UO_962 (O_962,N_14855,N_13206);
or UO_963 (O_963,N_12340,N_13656);
nor UO_964 (O_964,N_12875,N_13491);
nor UO_965 (O_965,N_13593,N_12214);
and UO_966 (O_966,N_12550,N_14805);
and UO_967 (O_967,N_12818,N_13304);
and UO_968 (O_968,N_12287,N_14491);
nor UO_969 (O_969,N_13212,N_12841);
nor UO_970 (O_970,N_12310,N_13204);
nand UO_971 (O_971,N_12324,N_14141);
or UO_972 (O_972,N_12683,N_13374);
nand UO_973 (O_973,N_13945,N_12290);
or UO_974 (O_974,N_13415,N_12049);
nor UO_975 (O_975,N_12542,N_13193);
or UO_976 (O_976,N_13092,N_13216);
and UO_977 (O_977,N_12825,N_13915);
and UO_978 (O_978,N_13779,N_12002);
nand UO_979 (O_979,N_13265,N_13851);
and UO_980 (O_980,N_14034,N_12712);
nand UO_981 (O_981,N_14929,N_12801);
and UO_982 (O_982,N_12288,N_12544);
nand UO_983 (O_983,N_12157,N_13603);
xnor UO_984 (O_984,N_14419,N_12837);
or UO_985 (O_985,N_13676,N_12645);
xor UO_986 (O_986,N_12500,N_14962);
nor UO_987 (O_987,N_13240,N_12557);
and UO_988 (O_988,N_13597,N_12876);
and UO_989 (O_989,N_12659,N_13601);
or UO_990 (O_990,N_14886,N_13447);
or UO_991 (O_991,N_12193,N_12150);
or UO_992 (O_992,N_12256,N_14728);
xor UO_993 (O_993,N_12507,N_13970);
nand UO_994 (O_994,N_14717,N_13264);
xor UO_995 (O_995,N_14971,N_12017);
nand UO_996 (O_996,N_14622,N_14359);
and UO_997 (O_997,N_12298,N_14502);
xnor UO_998 (O_998,N_14574,N_12738);
nand UO_999 (O_999,N_13293,N_14799);
and UO_1000 (O_1000,N_13739,N_14084);
nand UO_1001 (O_1001,N_12811,N_13755);
nand UO_1002 (O_1002,N_14834,N_14883);
nand UO_1003 (O_1003,N_14720,N_14821);
or UO_1004 (O_1004,N_13919,N_12051);
nand UO_1005 (O_1005,N_12420,N_14584);
xnor UO_1006 (O_1006,N_14291,N_13410);
or UO_1007 (O_1007,N_13828,N_14323);
or UO_1008 (O_1008,N_13472,N_12171);
and UO_1009 (O_1009,N_14859,N_12096);
nor UO_1010 (O_1010,N_14665,N_14553);
or UO_1011 (O_1011,N_14402,N_14062);
or UO_1012 (O_1012,N_12721,N_13226);
nor UO_1013 (O_1013,N_12271,N_12902);
or UO_1014 (O_1014,N_12991,N_12181);
nor UO_1015 (O_1015,N_13966,N_13633);
xnor UO_1016 (O_1016,N_12787,N_13310);
nand UO_1017 (O_1017,N_12622,N_14331);
and UO_1018 (O_1018,N_14758,N_12494);
or UO_1019 (O_1019,N_12505,N_13039);
nand UO_1020 (O_1020,N_13778,N_14807);
xor UO_1021 (O_1021,N_14035,N_14703);
nor UO_1022 (O_1022,N_12967,N_14890);
and UO_1023 (O_1023,N_12999,N_13904);
or UO_1024 (O_1024,N_13306,N_14854);
or UO_1025 (O_1025,N_12548,N_12594);
xnor UO_1026 (O_1026,N_13877,N_14512);
or UO_1027 (O_1027,N_14961,N_14007);
and UO_1028 (O_1028,N_12835,N_13245);
nor UO_1029 (O_1029,N_12261,N_14950);
or UO_1030 (O_1030,N_13640,N_12597);
or UO_1031 (O_1031,N_13227,N_12375);
xor UO_1032 (O_1032,N_12821,N_12693);
xnor UO_1033 (O_1033,N_14417,N_14270);
and UO_1034 (O_1034,N_14569,N_14086);
nor UO_1035 (O_1035,N_14161,N_12496);
xnor UO_1036 (O_1036,N_12688,N_12097);
nand UO_1037 (O_1037,N_13502,N_13757);
xor UO_1038 (O_1038,N_14165,N_12785);
or UO_1039 (O_1039,N_13063,N_13979);
or UO_1040 (O_1040,N_13631,N_12531);
and UO_1041 (O_1041,N_12286,N_13287);
or UO_1042 (O_1042,N_13093,N_13465);
and UO_1043 (O_1043,N_12960,N_12856);
nand UO_1044 (O_1044,N_14461,N_12513);
nand UO_1045 (O_1045,N_12997,N_13074);
nand UO_1046 (O_1046,N_12539,N_14497);
and UO_1047 (O_1047,N_14178,N_14234);
nand UO_1048 (O_1048,N_13651,N_14081);
nand UO_1049 (O_1049,N_14102,N_14898);
or UO_1050 (O_1050,N_12245,N_13653);
nor UO_1051 (O_1051,N_12873,N_12534);
nor UO_1052 (O_1052,N_14301,N_14861);
and UO_1053 (O_1053,N_12159,N_13873);
or UO_1054 (O_1054,N_12215,N_14989);
nor UO_1055 (O_1055,N_14698,N_12141);
or UO_1056 (O_1056,N_12244,N_13660);
xor UO_1057 (O_1057,N_14617,N_13542);
nor UO_1058 (O_1058,N_12760,N_14557);
nor UO_1059 (O_1059,N_12634,N_12174);
and UO_1060 (O_1060,N_12360,N_14987);
and UO_1061 (O_1061,N_14187,N_14631);
or UO_1062 (O_1062,N_13554,N_13424);
nand UO_1063 (O_1063,N_12381,N_13299);
xor UO_1064 (O_1064,N_12266,N_12861);
nand UO_1065 (O_1065,N_14023,N_12988);
and UO_1066 (O_1066,N_12529,N_12948);
xnor UO_1067 (O_1067,N_14636,N_13519);
nor UO_1068 (O_1068,N_12458,N_14043);
or UO_1069 (O_1069,N_14258,N_12937);
xor UO_1070 (O_1070,N_14066,N_13148);
or UO_1071 (O_1071,N_14845,N_12430);
xor UO_1072 (O_1072,N_14410,N_12599);
or UO_1073 (O_1073,N_14482,N_14142);
xor UO_1074 (O_1074,N_12596,N_14276);
nand UO_1075 (O_1075,N_14498,N_14608);
or UO_1076 (O_1076,N_12701,N_12658);
or UO_1077 (O_1077,N_14699,N_12714);
xor UO_1078 (O_1078,N_14653,N_13431);
or UO_1079 (O_1079,N_14835,N_14029);
or UO_1080 (O_1080,N_13362,N_14269);
xnor UO_1081 (O_1081,N_13107,N_14088);
nand UO_1082 (O_1082,N_12759,N_12166);
nor UO_1083 (O_1083,N_12206,N_12679);
and UO_1084 (O_1084,N_13740,N_14588);
nand UO_1085 (O_1085,N_14073,N_13643);
xor UO_1086 (O_1086,N_14183,N_13826);
or UO_1087 (O_1087,N_12072,N_14628);
nor UO_1088 (O_1088,N_13726,N_13222);
or UO_1089 (O_1089,N_13228,N_13022);
xnor UO_1090 (O_1090,N_13573,N_14170);
or UO_1091 (O_1091,N_14555,N_13840);
nand UO_1092 (O_1092,N_12569,N_12686);
nand UO_1093 (O_1093,N_13705,N_13912);
xor UO_1094 (O_1094,N_12438,N_12323);
xnor UO_1095 (O_1095,N_12715,N_12927);
xor UO_1096 (O_1096,N_12647,N_13518);
or UO_1097 (O_1097,N_14514,N_12931);
or UO_1098 (O_1098,N_13224,N_12692);
nor UO_1099 (O_1099,N_12941,N_14324);
nand UO_1100 (O_1100,N_13684,N_12095);
nand UO_1101 (O_1101,N_12533,N_14164);
and UO_1102 (O_1102,N_14753,N_13214);
nand UO_1103 (O_1103,N_12177,N_14974);
xor UO_1104 (O_1104,N_14830,N_12828);
xnor UO_1105 (O_1105,N_12968,N_14210);
or UO_1106 (O_1106,N_12350,N_12125);
nand UO_1107 (O_1107,N_13132,N_13202);
and UO_1108 (O_1108,N_13266,N_13892);
and UO_1109 (O_1109,N_14530,N_14314);
and UO_1110 (O_1110,N_12376,N_14840);
nand UO_1111 (O_1111,N_14610,N_12386);
nor UO_1112 (O_1112,N_12601,N_13027);
nand UO_1113 (O_1113,N_12573,N_12765);
nor UO_1114 (O_1114,N_14452,N_13380);
nand UO_1115 (O_1115,N_13225,N_13815);
xnor UO_1116 (O_1116,N_13678,N_13674);
nand UO_1117 (O_1117,N_14152,N_13234);
and UO_1118 (O_1118,N_14409,N_13258);
or UO_1119 (O_1119,N_13106,N_12060);
and UO_1120 (O_1120,N_13964,N_14465);
xor UO_1121 (O_1121,N_12189,N_12154);
and UO_1122 (O_1122,N_12883,N_13589);
xnor UO_1123 (O_1123,N_13747,N_14762);
and UO_1124 (O_1124,N_13750,N_12945);
nand UO_1125 (O_1125,N_13021,N_13498);
nor UO_1126 (O_1126,N_13681,N_13611);
or UO_1127 (O_1127,N_13956,N_14696);
and UO_1128 (O_1128,N_12131,N_14095);
or UO_1129 (O_1129,N_14925,N_14349);
nor UO_1130 (O_1130,N_13987,N_13220);
xor UO_1131 (O_1131,N_12964,N_12784);
or UO_1132 (O_1132,N_14546,N_14281);
nor UO_1133 (O_1133,N_12369,N_12704);
and UO_1134 (O_1134,N_13110,N_13320);
and UO_1135 (O_1135,N_12990,N_13789);
nor UO_1136 (O_1136,N_14100,N_12924);
nor UO_1137 (O_1137,N_12417,N_13003);
nor UO_1138 (O_1138,N_14544,N_14480);
nor UO_1139 (O_1139,N_12210,N_14333);
or UO_1140 (O_1140,N_12449,N_14423);
and UO_1141 (O_1141,N_12058,N_12258);
or UO_1142 (O_1142,N_12732,N_12408);
or UO_1143 (O_1143,N_14078,N_14422);
or UO_1144 (O_1144,N_12136,N_13558);
nor UO_1145 (O_1145,N_14763,N_14941);
nand UO_1146 (O_1146,N_12722,N_14460);
and UO_1147 (O_1147,N_13559,N_13718);
and UO_1148 (O_1148,N_14876,N_13378);
xnor UO_1149 (O_1149,N_14866,N_12981);
xnor UO_1150 (O_1150,N_13969,N_14446);
and UO_1151 (O_1151,N_12241,N_13125);
xor UO_1152 (O_1152,N_14609,N_14366);
nand UO_1153 (O_1153,N_13010,N_13549);
nand UO_1154 (O_1154,N_13846,N_12112);
or UO_1155 (O_1155,N_14335,N_13689);
nand UO_1156 (O_1156,N_14319,N_13544);
nor UO_1157 (O_1157,N_12173,N_14914);
nor UO_1158 (O_1158,N_14596,N_13809);
xnor UO_1159 (O_1159,N_13702,N_14529);
xnor UO_1160 (O_1160,N_14249,N_14973);
nor UO_1161 (O_1161,N_14638,N_14438);
xnor UO_1162 (O_1162,N_14189,N_14687);
or UO_1163 (O_1163,N_14862,N_14877);
xnor UO_1164 (O_1164,N_12279,N_14682);
nand UO_1165 (O_1165,N_13614,N_13787);
nand UO_1166 (O_1166,N_14242,N_14207);
nand UO_1167 (O_1167,N_14959,N_13365);
xor UO_1168 (O_1168,N_14470,N_13963);
and UO_1169 (O_1169,N_12961,N_13057);
nand UO_1170 (O_1170,N_14345,N_13922);
and UO_1171 (O_1171,N_13790,N_12952);
or UO_1172 (O_1172,N_13013,N_12783);
nand UO_1173 (O_1173,N_12462,N_12432);
and UO_1174 (O_1174,N_14943,N_14436);
and UO_1175 (O_1175,N_13930,N_12192);
or UO_1176 (O_1176,N_12009,N_12802);
or UO_1177 (O_1177,N_14021,N_12923);
and UO_1178 (O_1178,N_12528,N_13033);
or UO_1179 (O_1179,N_14003,N_14414);
nor UO_1180 (O_1180,N_13883,N_14701);
or UO_1181 (O_1181,N_12012,N_12833);
and UO_1182 (O_1182,N_13723,N_14030);
or UO_1183 (O_1183,N_13752,N_12928);
xor UO_1184 (O_1184,N_14416,N_14338);
nand UO_1185 (O_1185,N_12093,N_12976);
or UO_1186 (O_1186,N_12663,N_14190);
xor UO_1187 (O_1187,N_12104,N_12552);
xor UO_1188 (O_1188,N_13839,N_12985);
nor UO_1189 (O_1189,N_13715,N_13268);
or UO_1190 (O_1190,N_12278,N_12836);
or UO_1191 (O_1191,N_13121,N_14644);
xnor UO_1192 (O_1192,N_14071,N_13454);
or UO_1193 (O_1193,N_14856,N_14734);
nand UO_1194 (O_1194,N_12092,N_12422);
and UO_1195 (O_1195,N_13567,N_12055);
and UO_1196 (O_1196,N_12809,N_14162);
xnor UO_1197 (O_1197,N_12191,N_12680);
or UO_1198 (O_1198,N_14982,N_12170);
xor UO_1199 (O_1199,N_14296,N_14798);
nand UO_1200 (O_1200,N_14267,N_13051);
nor UO_1201 (O_1201,N_12781,N_12472);
or UO_1202 (O_1202,N_13413,N_13069);
and UO_1203 (O_1203,N_13628,N_12982);
nor UO_1204 (O_1204,N_12560,N_13156);
or UO_1205 (O_1205,N_13302,N_13041);
xnor UO_1206 (O_1206,N_12282,N_12180);
nand UO_1207 (O_1207,N_13855,N_12158);
nor UO_1208 (O_1208,N_13546,N_14118);
nor UO_1209 (O_1209,N_12791,N_12236);
or UO_1210 (O_1210,N_13797,N_14766);
xnor UO_1211 (O_1211,N_14225,N_13925);
and UO_1212 (O_1212,N_14614,N_13579);
nand UO_1213 (O_1213,N_14231,N_12803);
nand UO_1214 (O_1214,N_13508,N_14105);
xnor UO_1215 (O_1215,N_12549,N_13038);
xor UO_1216 (O_1216,N_12578,N_13231);
and UO_1217 (O_1217,N_14424,N_13467);
or UO_1218 (O_1218,N_13849,N_12657);
nor UO_1219 (O_1219,N_12063,N_13730);
nand UO_1220 (O_1220,N_12973,N_12850);
nand UO_1221 (O_1221,N_13983,N_13152);
or UO_1222 (O_1222,N_14273,N_13477);
or UO_1223 (O_1223,N_13346,N_13471);
or UO_1224 (O_1224,N_12974,N_14721);
nand UO_1225 (O_1225,N_12248,N_14444);
xor UO_1226 (O_1226,N_12027,N_12014);
nand UO_1227 (O_1227,N_14626,N_13515);
nor UO_1228 (O_1228,N_13485,N_12423);
nand UO_1229 (O_1229,N_13906,N_14248);
nand UO_1230 (O_1230,N_14087,N_13568);
xnor UO_1231 (O_1231,N_12747,N_14639);
xnor UO_1232 (O_1232,N_12357,N_12559);
nand UO_1233 (O_1233,N_12468,N_14197);
or UO_1234 (O_1234,N_12834,N_13097);
or UO_1235 (O_1235,N_12238,N_14255);
nor UO_1236 (O_1236,N_13570,N_12499);
xnor UO_1237 (O_1237,N_12001,N_13318);
nand UO_1238 (O_1238,N_12414,N_12061);
and UO_1239 (O_1239,N_12867,N_12872);
nor UO_1240 (O_1240,N_13957,N_14780);
or UO_1241 (O_1241,N_12605,N_13572);
nor UO_1242 (O_1242,N_14853,N_13539);
or UO_1243 (O_1243,N_14286,N_12436);
or UO_1244 (O_1244,N_12756,N_13412);
xnor UO_1245 (O_1245,N_12753,N_13135);
xnor UO_1246 (O_1246,N_12707,N_14564);
nand UO_1247 (O_1247,N_14899,N_13060);
nand UO_1248 (O_1248,N_12231,N_13875);
nand UO_1249 (O_1249,N_14585,N_12547);
or UO_1250 (O_1250,N_14056,N_14572);
or UO_1251 (O_1251,N_13406,N_12391);
or UO_1252 (O_1252,N_13138,N_12003);
nand UO_1253 (O_1253,N_14166,N_12440);
nand UO_1254 (O_1254,N_12954,N_14582);
nand UO_1255 (O_1255,N_12303,N_13479);
nor UO_1256 (O_1256,N_14635,N_13691);
xnor UO_1257 (O_1257,N_14691,N_14801);
nand UO_1258 (O_1258,N_12864,N_13984);
nand UO_1259 (O_1259,N_12789,N_13303);
nor UO_1260 (O_1260,N_14984,N_12285);
xnor UO_1261 (O_1261,N_13277,N_13442);
nor UO_1262 (O_1262,N_14049,N_13630);
and UO_1263 (O_1263,N_12779,N_13576);
nand UO_1264 (O_1264,N_13417,N_14570);
nand UO_1265 (O_1265,N_13606,N_14752);
xnor UO_1266 (O_1266,N_12767,N_13360);
nand UO_1267 (O_1267,N_14127,N_12372);
nand UO_1268 (O_1268,N_13064,N_14891);
or UO_1269 (O_1269,N_13395,N_14226);
or UO_1270 (O_1270,N_13600,N_14694);
or UO_1271 (O_1271,N_13509,N_13749);
or UO_1272 (O_1272,N_13525,N_14033);
nand UO_1273 (O_1273,N_13997,N_14079);
nand UO_1274 (O_1274,N_12299,N_13172);
and UO_1275 (O_1275,N_13219,N_14137);
nand UO_1276 (O_1276,N_14656,N_14168);
or UO_1277 (O_1277,N_12579,N_14633);
nor UO_1278 (O_1278,N_12587,N_13109);
or UO_1279 (O_1279,N_12146,N_13776);
and UO_1280 (O_1280,N_12332,N_14678);
and UO_1281 (O_1281,N_13101,N_14315);
nand UO_1282 (O_1282,N_12275,N_14990);
and UO_1283 (O_1283,N_12911,N_13552);
and UO_1284 (O_1284,N_13090,N_13916);
and UO_1285 (O_1285,N_13394,N_13160);
xnor UO_1286 (O_1286,N_14252,N_12047);
or UO_1287 (O_1287,N_12485,N_12720);
nand UO_1288 (O_1288,N_14836,N_12237);
and UO_1289 (O_1289,N_13012,N_13452);
or UO_1290 (O_1290,N_12138,N_12654);
and UO_1291 (O_1291,N_12642,N_14765);
xnor UO_1292 (O_1292,N_13621,N_12532);
nor UO_1293 (O_1293,N_12703,N_14169);
nor UO_1294 (O_1294,N_13902,N_13024);
nor UO_1295 (O_1295,N_14911,N_12518);
xor UO_1296 (O_1296,N_14268,N_12239);
xnor UO_1297 (O_1297,N_14944,N_14233);
and UO_1298 (O_1298,N_12120,N_12036);
or UO_1299 (O_1299,N_12262,N_14825);
and UO_1300 (O_1300,N_12227,N_14543);
and UO_1301 (O_1301,N_14976,N_13123);
and UO_1302 (O_1302,N_13091,N_13516);
nor UO_1303 (O_1303,N_13407,N_12364);
or UO_1304 (O_1304,N_14602,N_13153);
or UO_1305 (O_1305,N_12441,N_12938);
or UO_1306 (O_1306,N_13825,N_13650);
nand UO_1307 (O_1307,N_14716,N_14237);
or UO_1308 (O_1308,N_13785,N_13866);
or UO_1309 (O_1309,N_13686,N_12689);
nand UO_1310 (O_1310,N_12762,N_12026);
xnor UO_1311 (O_1311,N_14745,N_12610);
xnor UO_1312 (O_1312,N_14318,N_12358);
and UO_1313 (O_1313,N_12561,N_12204);
or UO_1314 (O_1314,N_12196,N_13492);
or UO_1315 (O_1315,N_13707,N_13548);
or UO_1316 (O_1316,N_13598,N_12426);
or UO_1317 (O_1317,N_14892,N_13665);
and UO_1318 (O_1318,N_14238,N_14367);
nor UO_1319 (O_1319,N_13137,N_13475);
and UO_1320 (O_1320,N_12064,N_14473);
xnor UO_1321 (O_1321,N_14325,N_14864);
or UO_1322 (O_1322,N_14851,N_14356);
or UO_1323 (O_1323,N_13084,N_12723);
nor UO_1324 (O_1324,N_13340,N_12421);
and UO_1325 (O_1325,N_13868,N_14154);
and UO_1326 (O_1326,N_12630,N_12424);
nand UO_1327 (O_1327,N_14533,N_13457);
and UO_1328 (O_1328,N_13118,N_13162);
or UO_1329 (O_1329,N_14271,N_14070);
or UO_1330 (O_1330,N_14875,N_13120);
nor UO_1331 (O_1331,N_14872,N_13753);
xnor UO_1332 (O_1332,N_14942,N_13955);
nor UO_1333 (O_1333,N_14015,N_12217);
nand UO_1334 (O_1334,N_12843,N_14623);
and UO_1335 (O_1335,N_14392,N_12541);
and UO_1336 (O_1336,N_14251,N_14894);
xor UO_1337 (O_1337,N_12336,N_13586);
nand UO_1338 (O_1338,N_13989,N_12144);
xnor UO_1339 (O_1339,N_14427,N_13126);
nor UO_1340 (O_1340,N_14133,N_14604);
or UO_1341 (O_1341,N_14981,N_13342);
nor UO_1342 (O_1342,N_14802,N_14711);
nor UO_1343 (O_1343,N_14481,N_12393);
xnor UO_1344 (O_1344,N_12822,N_13886);
and UO_1345 (O_1345,N_12848,N_12268);
or UO_1346 (O_1346,N_14576,N_13577);
xor UO_1347 (O_1347,N_12540,N_14107);
or UO_1348 (O_1348,N_12766,N_14090);
nor UO_1349 (O_1349,N_12888,N_14158);
nand UO_1350 (O_1350,N_14713,N_13448);
nand UO_1351 (O_1351,N_14486,N_14963);
and UO_1352 (O_1352,N_13414,N_13583);
nor UO_1353 (O_1353,N_12859,N_13698);
xor UO_1354 (O_1354,N_13116,N_13692);
nand UO_1355 (O_1355,N_13486,N_12612);
and UO_1356 (O_1356,N_14120,N_12776);
nor UO_1357 (O_1357,N_14223,N_14057);
nor UO_1358 (O_1358,N_13513,N_13899);
xnor UO_1359 (O_1359,N_12965,N_14388);
nand UO_1360 (O_1360,N_14478,N_13058);
nand UO_1361 (O_1361,N_14908,N_12481);
xor UO_1362 (O_1362,N_12307,N_13054);
xor UO_1363 (O_1363,N_13994,N_13281);
nand UO_1364 (O_1364,N_13967,N_12030);
nor UO_1365 (O_1365,N_12498,N_13507);
xnor UO_1366 (O_1366,N_12522,N_12315);
nand UO_1367 (O_1367,N_12297,N_12333);
or UO_1368 (O_1368,N_12435,N_13391);
and UO_1369 (O_1369,N_12200,N_12090);
xor UO_1370 (O_1370,N_12959,N_13014);
or UO_1371 (O_1371,N_13742,N_12152);
or UO_1372 (O_1372,N_14627,N_14241);
and UO_1373 (O_1373,N_14134,N_14403);
xor UO_1374 (O_1374,N_14526,N_12511);
nand UO_1375 (O_1375,N_12140,N_13530);
nand UO_1376 (O_1376,N_12768,N_14437);
and UO_1377 (O_1377,N_13532,N_13645);
or UO_1378 (O_1378,N_14867,N_14755);
nand UO_1379 (O_1379,N_13885,N_12751);
xnor UO_1380 (O_1380,N_13239,N_14463);
or UO_1381 (O_1381,N_13117,N_13869);
nand UO_1382 (O_1382,N_12660,N_12944);
or UO_1383 (O_1383,N_12526,N_13460);
nand UO_1384 (O_1384,N_13321,N_13623);
and UO_1385 (O_1385,N_12062,N_14616);
and UO_1386 (O_1386,N_12135,N_13402);
or UO_1387 (O_1387,N_12637,N_12439);
nor UO_1388 (O_1388,N_14282,N_12524);
nand UO_1389 (O_1389,N_13527,N_13804);
nor UO_1390 (O_1390,N_13837,N_13000);
xor UO_1391 (O_1391,N_12983,N_13999);
and UO_1392 (O_1392,N_13824,N_13932);
nor UO_1393 (O_1393,N_14383,N_13768);
and UO_1394 (O_1394,N_14874,N_13344);
nand UO_1395 (O_1395,N_14986,N_12921);
and UO_1396 (O_1396,N_13538,N_13453);
nor UO_1397 (O_1397,N_13229,N_13897);
or UO_1398 (O_1398,N_12804,N_13842);
or UO_1399 (O_1399,N_13976,N_12342);
and UO_1400 (O_1400,N_12678,N_14380);
and UO_1401 (O_1401,N_14998,N_14739);
xor UO_1402 (O_1402,N_13625,N_14695);
and UO_1403 (O_1403,N_12101,N_13236);
and UO_1404 (O_1404,N_14011,N_12761);
xor UO_1405 (O_1405,N_13798,N_13836);
nand UO_1406 (O_1406,N_14010,N_13511);
or UO_1407 (O_1407,N_14764,N_13615);
xnor UO_1408 (O_1408,N_13275,N_12537);
xor UO_1409 (O_1409,N_12069,N_14404);
nor UO_1410 (O_1410,N_13617,N_13451);
nand UO_1411 (O_1411,N_12148,N_14143);
nand UO_1412 (O_1412,N_14786,N_12469);
and UO_1413 (O_1413,N_14847,N_13566);
xnor UO_1414 (O_1414,N_14777,N_14397);
nand UO_1415 (O_1415,N_14346,N_13085);
xor UO_1416 (O_1416,N_12525,N_14374);
and UO_1417 (O_1417,N_13384,N_14194);
nor UO_1418 (O_1418,N_14017,N_12274);
nand UO_1419 (O_1419,N_14204,N_14949);
or UO_1420 (O_1420,N_14334,N_14706);
nor UO_1421 (O_1421,N_13073,N_13909);
and UO_1422 (O_1422,N_12588,N_13814);
or UO_1423 (O_1423,N_14384,N_12348);
and UO_1424 (O_1424,N_13102,N_13514);
and UO_1425 (O_1425,N_12613,N_12235);
or UO_1426 (O_1426,N_13534,N_13217);
or UO_1427 (O_1427,N_13072,N_12830);
or UO_1428 (O_1428,N_12467,N_13295);
nand UO_1429 (O_1429,N_13056,N_14239);
nor UO_1430 (O_1430,N_13330,N_14377);
or UO_1431 (O_1431,N_13991,N_13201);
or UO_1432 (O_1432,N_12343,N_12951);
nor UO_1433 (O_1433,N_12205,N_13357);
and UO_1434 (O_1434,N_13343,N_14412);
nand UO_1435 (O_1435,N_14175,N_13184);
nor UO_1436 (O_1436,N_12356,N_14195);
nand UO_1437 (O_1437,N_13482,N_12664);
and UO_1438 (O_1438,N_12284,N_14965);
and UO_1439 (O_1439,N_14048,N_13466);
xnor UO_1440 (O_1440,N_12619,N_14054);
nand UO_1441 (O_1441,N_14668,N_13083);
or UO_1442 (O_1442,N_12748,N_12790);
or UO_1443 (O_1443,N_13432,N_13671);
nor UO_1444 (O_1444,N_14188,N_14651);
xor UO_1445 (O_1445,N_14198,N_13317);
or UO_1446 (O_1446,N_12726,N_14709);
and UO_1447 (O_1447,N_14697,N_13199);
nor UO_1448 (O_1448,N_13741,N_13149);
nand UO_1449 (O_1449,N_14827,N_13690);
or UO_1450 (O_1450,N_13167,N_14038);
xnor UO_1451 (O_1451,N_12145,N_12728);
and UO_1452 (O_1452,N_13612,N_13059);
xnor UO_1453 (O_1453,N_14408,N_14337);
nor UO_1454 (O_1454,N_14122,N_13772);
nand UO_1455 (O_1455,N_12328,N_14303);
and UO_1456 (O_1456,N_13408,N_14670);
nand UO_1457 (O_1457,N_14771,N_13099);
nor UO_1458 (O_1458,N_12614,N_13455);
and UO_1459 (O_1459,N_14119,N_12224);
nand UO_1460 (O_1460,N_14885,N_13075);
nand UO_1461 (O_1461,N_13841,N_13719);
nor UO_1462 (O_1462,N_14724,N_12886);
and UO_1463 (O_1463,N_12020,N_12838);
nor UO_1464 (O_1464,N_13480,N_12935);
and UO_1465 (O_1465,N_13952,N_14111);
xor UO_1466 (O_1466,N_13713,N_13821);
and UO_1467 (O_1467,N_12115,N_13700);
xor UO_1468 (O_1468,N_13666,N_13763);
and UO_1469 (O_1469,N_14103,N_14903);
nand UO_1470 (O_1470,N_12025,N_14075);
or UO_1471 (O_1471,N_14469,N_14562);
and UO_1472 (O_1472,N_14330,N_14028);
nand UO_1473 (O_1473,N_14792,N_12892);
and UO_1474 (O_1474,N_13639,N_13938);
xnor UO_1475 (O_1475,N_12725,N_13865);
and UO_1476 (O_1476,N_13595,N_12746);
nor UO_1477 (O_1477,N_12201,N_14819);
and UO_1478 (O_1478,N_14370,N_14793);
or UO_1479 (O_1479,N_12799,N_14882);
or UO_1480 (O_1480,N_13336,N_13782);
nand UO_1481 (O_1481,N_14304,N_12308);
nand UO_1482 (O_1482,N_13237,N_12570);
nand UO_1483 (O_1483,N_12617,N_14181);
nand UO_1484 (O_1484,N_14688,N_14938);
nand UO_1485 (O_1485,N_12365,N_14723);
nand UO_1486 (O_1486,N_14967,N_12671);
xnor UO_1487 (O_1487,N_12175,N_14787);
xnor UO_1488 (O_1488,N_13968,N_14253);
nor UO_1489 (O_1489,N_13311,N_13720);
xor UO_1490 (O_1490,N_12519,N_14566);
and UO_1491 (O_1491,N_12465,N_14768);
or UO_1492 (O_1492,N_12582,N_14888);
xor UO_1493 (O_1493,N_12989,N_14719);
and UO_1494 (O_1494,N_13429,N_13751);
nor UO_1495 (O_1495,N_14772,N_12301);
xor UO_1496 (O_1496,N_14163,N_12901);
nor UO_1497 (O_1497,N_12716,N_12445);
and UO_1498 (O_1498,N_12383,N_13396);
and UO_1499 (O_1499,N_13820,N_13972);
xnor UO_1500 (O_1500,N_12008,N_14593);
nor UO_1501 (O_1501,N_13062,N_13147);
or UO_1502 (O_1502,N_14741,N_13171);
nor UO_1503 (O_1503,N_14356,N_14457);
nor UO_1504 (O_1504,N_13283,N_12821);
and UO_1505 (O_1505,N_12865,N_14343);
or UO_1506 (O_1506,N_12221,N_12179);
nand UO_1507 (O_1507,N_13182,N_13561);
xnor UO_1508 (O_1508,N_12315,N_12691);
xnor UO_1509 (O_1509,N_14100,N_13657);
or UO_1510 (O_1510,N_13355,N_13627);
nor UO_1511 (O_1511,N_14279,N_13216);
nor UO_1512 (O_1512,N_14054,N_12132);
nand UO_1513 (O_1513,N_14578,N_14651);
and UO_1514 (O_1514,N_14865,N_13012);
nor UO_1515 (O_1515,N_12068,N_13561);
or UO_1516 (O_1516,N_14251,N_14642);
nor UO_1517 (O_1517,N_12667,N_12903);
and UO_1518 (O_1518,N_14141,N_12799);
nand UO_1519 (O_1519,N_13740,N_13639);
nor UO_1520 (O_1520,N_13696,N_13643);
xor UO_1521 (O_1521,N_12432,N_13041);
or UO_1522 (O_1522,N_13951,N_12497);
nor UO_1523 (O_1523,N_14310,N_13002);
nor UO_1524 (O_1524,N_14853,N_13737);
nor UO_1525 (O_1525,N_14052,N_13970);
and UO_1526 (O_1526,N_12313,N_13484);
or UO_1527 (O_1527,N_14899,N_14313);
xor UO_1528 (O_1528,N_13855,N_12529);
and UO_1529 (O_1529,N_13068,N_12105);
xnor UO_1530 (O_1530,N_13418,N_12516);
xnor UO_1531 (O_1531,N_12562,N_12813);
xor UO_1532 (O_1532,N_14396,N_13607);
and UO_1533 (O_1533,N_14908,N_14752);
or UO_1534 (O_1534,N_12569,N_13068);
nor UO_1535 (O_1535,N_13811,N_12251);
nand UO_1536 (O_1536,N_14797,N_14563);
or UO_1537 (O_1537,N_12671,N_12678);
or UO_1538 (O_1538,N_13558,N_12575);
and UO_1539 (O_1539,N_12464,N_12841);
nor UO_1540 (O_1540,N_12473,N_13696);
xnor UO_1541 (O_1541,N_13300,N_14214);
xor UO_1542 (O_1542,N_13335,N_14329);
or UO_1543 (O_1543,N_12838,N_13135);
and UO_1544 (O_1544,N_12961,N_14558);
and UO_1545 (O_1545,N_13096,N_12911);
nand UO_1546 (O_1546,N_14670,N_14372);
or UO_1547 (O_1547,N_14009,N_14193);
nand UO_1548 (O_1548,N_12867,N_14848);
and UO_1549 (O_1549,N_14613,N_14206);
nand UO_1550 (O_1550,N_14835,N_12702);
or UO_1551 (O_1551,N_14404,N_12875);
nor UO_1552 (O_1552,N_14810,N_14736);
nand UO_1553 (O_1553,N_14243,N_14490);
nor UO_1554 (O_1554,N_13415,N_14495);
xnor UO_1555 (O_1555,N_14551,N_13340);
and UO_1556 (O_1556,N_14287,N_13067);
nor UO_1557 (O_1557,N_13966,N_13032);
or UO_1558 (O_1558,N_13270,N_13236);
nor UO_1559 (O_1559,N_14283,N_13758);
and UO_1560 (O_1560,N_12055,N_14800);
nand UO_1561 (O_1561,N_13483,N_12469);
and UO_1562 (O_1562,N_13561,N_14992);
xor UO_1563 (O_1563,N_12828,N_14553);
nor UO_1564 (O_1564,N_13972,N_12909);
xnor UO_1565 (O_1565,N_14744,N_14692);
and UO_1566 (O_1566,N_14816,N_13955);
nand UO_1567 (O_1567,N_13167,N_14316);
and UO_1568 (O_1568,N_12689,N_12751);
xor UO_1569 (O_1569,N_14715,N_14133);
and UO_1570 (O_1570,N_14119,N_14955);
nand UO_1571 (O_1571,N_12211,N_12852);
nand UO_1572 (O_1572,N_13964,N_12818);
and UO_1573 (O_1573,N_14092,N_12080);
and UO_1574 (O_1574,N_13147,N_13544);
or UO_1575 (O_1575,N_12311,N_13128);
xnor UO_1576 (O_1576,N_14936,N_12948);
xnor UO_1577 (O_1577,N_13335,N_13529);
and UO_1578 (O_1578,N_13168,N_13238);
nand UO_1579 (O_1579,N_13051,N_13624);
nand UO_1580 (O_1580,N_12935,N_12414);
or UO_1581 (O_1581,N_13899,N_13410);
and UO_1582 (O_1582,N_12691,N_12506);
nor UO_1583 (O_1583,N_14004,N_14587);
nand UO_1584 (O_1584,N_13620,N_14519);
and UO_1585 (O_1585,N_13626,N_14342);
and UO_1586 (O_1586,N_12245,N_12346);
or UO_1587 (O_1587,N_12891,N_14301);
xnor UO_1588 (O_1588,N_13557,N_12490);
or UO_1589 (O_1589,N_13190,N_12210);
or UO_1590 (O_1590,N_13475,N_14908);
or UO_1591 (O_1591,N_14714,N_14014);
or UO_1592 (O_1592,N_12558,N_13414);
and UO_1593 (O_1593,N_13878,N_14142);
nor UO_1594 (O_1594,N_13761,N_14968);
and UO_1595 (O_1595,N_13014,N_12963);
and UO_1596 (O_1596,N_13527,N_14073);
xor UO_1597 (O_1597,N_14257,N_12916);
and UO_1598 (O_1598,N_12165,N_12048);
xnor UO_1599 (O_1599,N_12857,N_12868);
and UO_1600 (O_1600,N_12614,N_14467);
or UO_1601 (O_1601,N_12285,N_12644);
nand UO_1602 (O_1602,N_13488,N_12859);
or UO_1603 (O_1603,N_12420,N_13806);
nor UO_1604 (O_1604,N_14426,N_14847);
xor UO_1605 (O_1605,N_14703,N_12761);
or UO_1606 (O_1606,N_13031,N_12093);
nor UO_1607 (O_1607,N_12765,N_12902);
nor UO_1608 (O_1608,N_14204,N_14054);
nor UO_1609 (O_1609,N_12949,N_14082);
or UO_1610 (O_1610,N_13442,N_13876);
nand UO_1611 (O_1611,N_12761,N_14434);
and UO_1612 (O_1612,N_13711,N_13149);
xor UO_1613 (O_1613,N_14861,N_12027);
nor UO_1614 (O_1614,N_13296,N_14990);
nor UO_1615 (O_1615,N_12138,N_14288);
or UO_1616 (O_1616,N_14729,N_13315);
or UO_1617 (O_1617,N_12951,N_13208);
nand UO_1618 (O_1618,N_13751,N_12283);
nor UO_1619 (O_1619,N_13056,N_12750);
nand UO_1620 (O_1620,N_13439,N_14002);
nor UO_1621 (O_1621,N_12044,N_14310);
xor UO_1622 (O_1622,N_13620,N_12998);
or UO_1623 (O_1623,N_14477,N_13084);
xnor UO_1624 (O_1624,N_13967,N_14086);
and UO_1625 (O_1625,N_13120,N_12994);
or UO_1626 (O_1626,N_13771,N_14818);
or UO_1627 (O_1627,N_14971,N_14052);
and UO_1628 (O_1628,N_14288,N_14554);
xor UO_1629 (O_1629,N_12745,N_12811);
nand UO_1630 (O_1630,N_13181,N_13057);
or UO_1631 (O_1631,N_13244,N_13452);
or UO_1632 (O_1632,N_14538,N_14782);
xnor UO_1633 (O_1633,N_13688,N_12985);
nor UO_1634 (O_1634,N_12541,N_14678);
nand UO_1635 (O_1635,N_14140,N_13796);
nor UO_1636 (O_1636,N_12960,N_14422);
xnor UO_1637 (O_1637,N_13426,N_12909);
nand UO_1638 (O_1638,N_12467,N_13841);
nor UO_1639 (O_1639,N_13717,N_12617);
nor UO_1640 (O_1640,N_12388,N_12769);
nand UO_1641 (O_1641,N_14212,N_13541);
xnor UO_1642 (O_1642,N_14642,N_12355);
nand UO_1643 (O_1643,N_14142,N_14107);
or UO_1644 (O_1644,N_14942,N_12481);
nand UO_1645 (O_1645,N_14422,N_12972);
nand UO_1646 (O_1646,N_12378,N_13344);
nand UO_1647 (O_1647,N_13525,N_12631);
nor UO_1648 (O_1648,N_12259,N_13883);
and UO_1649 (O_1649,N_13079,N_13947);
and UO_1650 (O_1650,N_13681,N_12459);
nor UO_1651 (O_1651,N_13795,N_13807);
or UO_1652 (O_1652,N_14891,N_12544);
xnor UO_1653 (O_1653,N_13493,N_12132);
or UO_1654 (O_1654,N_14011,N_14662);
nor UO_1655 (O_1655,N_13729,N_12121);
xnor UO_1656 (O_1656,N_14408,N_12457);
nand UO_1657 (O_1657,N_14885,N_14219);
and UO_1658 (O_1658,N_13532,N_14619);
nand UO_1659 (O_1659,N_13312,N_14279);
or UO_1660 (O_1660,N_12123,N_13691);
or UO_1661 (O_1661,N_12646,N_12413);
and UO_1662 (O_1662,N_13428,N_14637);
or UO_1663 (O_1663,N_13888,N_14093);
nand UO_1664 (O_1664,N_12406,N_12210);
xor UO_1665 (O_1665,N_14298,N_12928);
and UO_1666 (O_1666,N_12665,N_13801);
or UO_1667 (O_1667,N_13722,N_13555);
nand UO_1668 (O_1668,N_14129,N_12785);
or UO_1669 (O_1669,N_13535,N_13868);
and UO_1670 (O_1670,N_14926,N_12162);
nor UO_1671 (O_1671,N_14676,N_12826);
nor UO_1672 (O_1672,N_12286,N_14247);
and UO_1673 (O_1673,N_13839,N_12244);
xnor UO_1674 (O_1674,N_14936,N_13517);
nor UO_1675 (O_1675,N_12255,N_12580);
xnor UO_1676 (O_1676,N_13081,N_13249);
xor UO_1677 (O_1677,N_14736,N_12131);
nor UO_1678 (O_1678,N_13432,N_12711);
nand UO_1679 (O_1679,N_12071,N_12234);
xnor UO_1680 (O_1680,N_12768,N_12551);
or UO_1681 (O_1681,N_14563,N_12889);
xnor UO_1682 (O_1682,N_13412,N_12904);
and UO_1683 (O_1683,N_14027,N_12173);
or UO_1684 (O_1684,N_13831,N_12751);
and UO_1685 (O_1685,N_14008,N_13584);
and UO_1686 (O_1686,N_14438,N_13812);
xnor UO_1687 (O_1687,N_12317,N_13395);
xnor UO_1688 (O_1688,N_14817,N_13026);
nand UO_1689 (O_1689,N_12541,N_14110);
or UO_1690 (O_1690,N_12764,N_12902);
or UO_1691 (O_1691,N_12659,N_14533);
and UO_1692 (O_1692,N_14237,N_14604);
and UO_1693 (O_1693,N_12838,N_14672);
xor UO_1694 (O_1694,N_12197,N_12327);
nor UO_1695 (O_1695,N_12883,N_12925);
or UO_1696 (O_1696,N_13041,N_12114);
and UO_1697 (O_1697,N_14293,N_12741);
and UO_1698 (O_1698,N_13266,N_12859);
xor UO_1699 (O_1699,N_14614,N_13710);
nor UO_1700 (O_1700,N_14822,N_12648);
nand UO_1701 (O_1701,N_13139,N_12980);
xor UO_1702 (O_1702,N_14447,N_12904);
and UO_1703 (O_1703,N_12708,N_13663);
nand UO_1704 (O_1704,N_12249,N_14890);
nor UO_1705 (O_1705,N_14241,N_12480);
and UO_1706 (O_1706,N_13340,N_12678);
or UO_1707 (O_1707,N_12352,N_13051);
and UO_1708 (O_1708,N_14308,N_12429);
and UO_1709 (O_1709,N_12710,N_14150);
xnor UO_1710 (O_1710,N_14939,N_14919);
xor UO_1711 (O_1711,N_14394,N_13522);
nand UO_1712 (O_1712,N_12614,N_12068);
nand UO_1713 (O_1713,N_14199,N_14700);
xor UO_1714 (O_1714,N_12031,N_14346);
xnor UO_1715 (O_1715,N_12412,N_12040);
and UO_1716 (O_1716,N_13558,N_14430);
xor UO_1717 (O_1717,N_13279,N_12484);
and UO_1718 (O_1718,N_13205,N_12730);
or UO_1719 (O_1719,N_14867,N_13084);
nor UO_1720 (O_1720,N_14136,N_14518);
nor UO_1721 (O_1721,N_13007,N_14601);
or UO_1722 (O_1722,N_14341,N_13156);
nand UO_1723 (O_1723,N_14007,N_12944);
xnor UO_1724 (O_1724,N_12354,N_14258);
and UO_1725 (O_1725,N_14285,N_13906);
and UO_1726 (O_1726,N_12481,N_12879);
or UO_1727 (O_1727,N_14611,N_13373);
nor UO_1728 (O_1728,N_13151,N_13372);
xnor UO_1729 (O_1729,N_12134,N_13670);
or UO_1730 (O_1730,N_14324,N_12571);
nand UO_1731 (O_1731,N_12366,N_13654);
nor UO_1732 (O_1732,N_13599,N_13515);
or UO_1733 (O_1733,N_12389,N_13589);
xor UO_1734 (O_1734,N_13538,N_13145);
nor UO_1735 (O_1735,N_13342,N_12420);
xnor UO_1736 (O_1736,N_12517,N_12794);
xnor UO_1737 (O_1737,N_14286,N_13029);
and UO_1738 (O_1738,N_12389,N_13492);
or UO_1739 (O_1739,N_14651,N_14100);
and UO_1740 (O_1740,N_13394,N_13763);
nor UO_1741 (O_1741,N_14778,N_12256);
or UO_1742 (O_1742,N_14043,N_12939);
and UO_1743 (O_1743,N_12180,N_12869);
nand UO_1744 (O_1744,N_12811,N_13291);
xnor UO_1745 (O_1745,N_14422,N_14881);
nand UO_1746 (O_1746,N_12388,N_13012);
and UO_1747 (O_1747,N_14100,N_14909);
nand UO_1748 (O_1748,N_13915,N_13091);
nor UO_1749 (O_1749,N_12532,N_13642);
xnor UO_1750 (O_1750,N_14966,N_13725);
nor UO_1751 (O_1751,N_14609,N_14454);
nor UO_1752 (O_1752,N_12937,N_12382);
nor UO_1753 (O_1753,N_14627,N_12151);
or UO_1754 (O_1754,N_13193,N_13617);
xnor UO_1755 (O_1755,N_12355,N_14943);
or UO_1756 (O_1756,N_14558,N_12155);
nand UO_1757 (O_1757,N_12917,N_14230);
xnor UO_1758 (O_1758,N_14919,N_12690);
nand UO_1759 (O_1759,N_12197,N_14631);
xor UO_1760 (O_1760,N_14737,N_13045);
nand UO_1761 (O_1761,N_14757,N_12655);
or UO_1762 (O_1762,N_14884,N_12512);
nor UO_1763 (O_1763,N_12953,N_13592);
xnor UO_1764 (O_1764,N_13705,N_14176);
or UO_1765 (O_1765,N_13362,N_13034);
and UO_1766 (O_1766,N_13326,N_14930);
or UO_1767 (O_1767,N_14456,N_12922);
nand UO_1768 (O_1768,N_13090,N_13316);
and UO_1769 (O_1769,N_12055,N_13460);
and UO_1770 (O_1770,N_12921,N_14412);
nor UO_1771 (O_1771,N_12515,N_14183);
nand UO_1772 (O_1772,N_14497,N_14545);
nor UO_1773 (O_1773,N_13680,N_14799);
nor UO_1774 (O_1774,N_12916,N_12770);
xor UO_1775 (O_1775,N_13188,N_13109);
nor UO_1776 (O_1776,N_12199,N_12293);
xor UO_1777 (O_1777,N_13503,N_13447);
nor UO_1778 (O_1778,N_13614,N_12326);
or UO_1779 (O_1779,N_14393,N_12168);
nor UO_1780 (O_1780,N_13424,N_12331);
and UO_1781 (O_1781,N_12868,N_12783);
nor UO_1782 (O_1782,N_13620,N_13789);
nor UO_1783 (O_1783,N_12270,N_14661);
or UO_1784 (O_1784,N_12084,N_14448);
nand UO_1785 (O_1785,N_14539,N_14283);
or UO_1786 (O_1786,N_13971,N_12025);
xnor UO_1787 (O_1787,N_14484,N_12174);
and UO_1788 (O_1788,N_13571,N_13859);
xor UO_1789 (O_1789,N_14736,N_14440);
nor UO_1790 (O_1790,N_12007,N_14920);
or UO_1791 (O_1791,N_12692,N_12645);
and UO_1792 (O_1792,N_13019,N_13768);
nor UO_1793 (O_1793,N_14894,N_14739);
or UO_1794 (O_1794,N_13675,N_13357);
nand UO_1795 (O_1795,N_14405,N_13140);
and UO_1796 (O_1796,N_14678,N_13011);
or UO_1797 (O_1797,N_12849,N_13443);
nand UO_1798 (O_1798,N_14870,N_14568);
nand UO_1799 (O_1799,N_14276,N_13825);
nand UO_1800 (O_1800,N_13388,N_14693);
or UO_1801 (O_1801,N_14786,N_14916);
nand UO_1802 (O_1802,N_13053,N_14004);
xnor UO_1803 (O_1803,N_13188,N_12914);
and UO_1804 (O_1804,N_14032,N_14665);
and UO_1805 (O_1805,N_14619,N_13245);
nor UO_1806 (O_1806,N_12771,N_12301);
xor UO_1807 (O_1807,N_14450,N_13069);
and UO_1808 (O_1808,N_13218,N_13009);
and UO_1809 (O_1809,N_13488,N_13111);
xnor UO_1810 (O_1810,N_14978,N_12690);
and UO_1811 (O_1811,N_12639,N_13559);
and UO_1812 (O_1812,N_13856,N_14333);
nor UO_1813 (O_1813,N_13426,N_12536);
and UO_1814 (O_1814,N_14402,N_14355);
and UO_1815 (O_1815,N_13234,N_14272);
or UO_1816 (O_1816,N_13410,N_13112);
nand UO_1817 (O_1817,N_13358,N_12205);
nand UO_1818 (O_1818,N_14782,N_12014);
or UO_1819 (O_1819,N_12739,N_14895);
and UO_1820 (O_1820,N_12831,N_13947);
or UO_1821 (O_1821,N_13522,N_12088);
nor UO_1822 (O_1822,N_12744,N_13930);
and UO_1823 (O_1823,N_13298,N_13361);
nor UO_1824 (O_1824,N_12003,N_14221);
and UO_1825 (O_1825,N_12525,N_14874);
xor UO_1826 (O_1826,N_13492,N_12706);
nand UO_1827 (O_1827,N_12077,N_13000);
nor UO_1828 (O_1828,N_13610,N_14974);
and UO_1829 (O_1829,N_13908,N_12418);
nor UO_1830 (O_1830,N_14672,N_14137);
xor UO_1831 (O_1831,N_14660,N_13155);
nor UO_1832 (O_1832,N_13520,N_13778);
and UO_1833 (O_1833,N_14709,N_12776);
and UO_1834 (O_1834,N_12261,N_13169);
nand UO_1835 (O_1835,N_14181,N_14443);
nor UO_1836 (O_1836,N_13171,N_14191);
nand UO_1837 (O_1837,N_13624,N_13050);
nor UO_1838 (O_1838,N_14760,N_14724);
nor UO_1839 (O_1839,N_13221,N_14501);
or UO_1840 (O_1840,N_12969,N_12606);
nor UO_1841 (O_1841,N_12432,N_14794);
or UO_1842 (O_1842,N_12045,N_12406);
xnor UO_1843 (O_1843,N_14119,N_12850);
xor UO_1844 (O_1844,N_14386,N_14872);
or UO_1845 (O_1845,N_12744,N_14811);
nand UO_1846 (O_1846,N_14848,N_12919);
nor UO_1847 (O_1847,N_12941,N_12196);
and UO_1848 (O_1848,N_14221,N_13933);
xor UO_1849 (O_1849,N_13125,N_12644);
nand UO_1850 (O_1850,N_12864,N_12647);
xor UO_1851 (O_1851,N_14904,N_12192);
nor UO_1852 (O_1852,N_14489,N_13235);
nor UO_1853 (O_1853,N_12113,N_12833);
xnor UO_1854 (O_1854,N_14927,N_14047);
and UO_1855 (O_1855,N_14192,N_12587);
xor UO_1856 (O_1856,N_13028,N_13670);
nand UO_1857 (O_1857,N_13700,N_12457);
or UO_1858 (O_1858,N_13210,N_14307);
or UO_1859 (O_1859,N_12684,N_14066);
nand UO_1860 (O_1860,N_14059,N_12660);
xor UO_1861 (O_1861,N_12844,N_12609);
or UO_1862 (O_1862,N_13755,N_13728);
and UO_1863 (O_1863,N_12168,N_12930);
or UO_1864 (O_1864,N_13423,N_12704);
xnor UO_1865 (O_1865,N_14516,N_13256);
nand UO_1866 (O_1866,N_12889,N_14066);
or UO_1867 (O_1867,N_14578,N_14046);
nor UO_1868 (O_1868,N_14187,N_14820);
nor UO_1869 (O_1869,N_12543,N_13475);
nand UO_1870 (O_1870,N_12567,N_12031);
or UO_1871 (O_1871,N_12219,N_13496);
xnor UO_1872 (O_1872,N_14362,N_14825);
nand UO_1873 (O_1873,N_13382,N_13198);
nand UO_1874 (O_1874,N_14404,N_12787);
nand UO_1875 (O_1875,N_12168,N_13567);
xnor UO_1876 (O_1876,N_13270,N_13210);
nor UO_1877 (O_1877,N_13871,N_13125);
xnor UO_1878 (O_1878,N_14483,N_14113);
or UO_1879 (O_1879,N_14327,N_13326);
and UO_1880 (O_1880,N_14998,N_12259);
nand UO_1881 (O_1881,N_12177,N_12556);
nor UO_1882 (O_1882,N_14716,N_14850);
nand UO_1883 (O_1883,N_12344,N_12695);
nor UO_1884 (O_1884,N_12547,N_14880);
nand UO_1885 (O_1885,N_13561,N_12657);
or UO_1886 (O_1886,N_12826,N_14543);
xnor UO_1887 (O_1887,N_13757,N_12661);
xor UO_1888 (O_1888,N_12276,N_12824);
xor UO_1889 (O_1889,N_12741,N_14805);
or UO_1890 (O_1890,N_14661,N_13519);
nor UO_1891 (O_1891,N_12671,N_14142);
nor UO_1892 (O_1892,N_13322,N_12362);
nor UO_1893 (O_1893,N_13833,N_12744);
or UO_1894 (O_1894,N_14512,N_12379);
xor UO_1895 (O_1895,N_12785,N_13009);
and UO_1896 (O_1896,N_14279,N_12373);
or UO_1897 (O_1897,N_12396,N_14963);
nand UO_1898 (O_1898,N_12790,N_14706);
xor UO_1899 (O_1899,N_14015,N_12543);
or UO_1900 (O_1900,N_12461,N_13821);
nand UO_1901 (O_1901,N_13648,N_14518);
and UO_1902 (O_1902,N_14604,N_12522);
and UO_1903 (O_1903,N_14896,N_13118);
xnor UO_1904 (O_1904,N_14612,N_13434);
nor UO_1905 (O_1905,N_13489,N_14795);
nor UO_1906 (O_1906,N_14650,N_12749);
xnor UO_1907 (O_1907,N_14795,N_14329);
and UO_1908 (O_1908,N_12234,N_14497);
and UO_1909 (O_1909,N_14399,N_14880);
nand UO_1910 (O_1910,N_13434,N_13283);
nand UO_1911 (O_1911,N_14692,N_13724);
or UO_1912 (O_1912,N_14673,N_13925);
nor UO_1913 (O_1913,N_12549,N_12764);
and UO_1914 (O_1914,N_13215,N_13718);
or UO_1915 (O_1915,N_14234,N_13518);
xnor UO_1916 (O_1916,N_13325,N_14451);
xor UO_1917 (O_1917,N_13306,N_13048);
or UO_1918 (O_1918,N_13049,N_14562);
or UO_1919 (O_1919,N_12671,N_14456);
xor UO_1920 (O_1920,N_13872,N_12718);
and UO_1921 (O_1921,N_13920,N_12535);
or UO_1922 (O_1922,N_13062,N_12477);
nor UO_1923 (O_1923,N_14330,N_14232);
and UO_1924 (O_1924,N_14635,N_12123);
and UO_1925 (O_1925,N_14934,N_13509);
nand UO_1926 (O_1926,N_14024,N_14556);
nor UO_1927 (O_1927,N_14268,N_13767);
nand UO_1928 (O_1928,N_13469,N_13544);
and UO_1929 (O_1929,N_12708,N_12256);
xor UO_1930 (O_1930,N_14594,N_13900);
or UO_1931 (O_1931,N_14800,N_14578);
xnor UO_1932 (O_1932,N_13372,N_12690);
or UO_1933 (O_1933,N_13497,N_13860);
xor UO_1934 (O_1934,N_12312,N_14203);
nand UO_1935 (O_1935,N_13124,N_14958);
or UO_1936 (O_1936,N_14488,N_13529);
nor UO_1937 (O_1937,N_14363,N_12846);
and UO_1938 (O_1938,N_13554,N_13961);
or UO_1939 (O_1939,N_14202,N_13704);
and UO_1940 (O_1940,N_12720,N_14690);
xnor UO_1941 (O_1941,N_12123,N_14581);
nor UO_1942 (O_1942,N_13244,N_13601);
xor UO_1943 (O_1943,N_13556,N_12689);
and UO_1944 (O_1944,N_14219,N_14366);
and UO_1945 (O_1945,N_14607,N_13194);
nor UO_1946 (O_1946,N_13385,N_13121);
or UO_1947 (O_1947,N_14313,N_14269);
or UO_1948 (O_1948,N_14923,N_12578);
nor UO_1949 (O_1949,N_13539,N_12482);
nand UO_1950 (O_1950,N_14758,N_12796);
and UO_1951 (O_1951,N_13363,N_14730);
or UO_1952 (O_1952,N_13993,N_13179);
nor UO_1953 (O_1953,N_12426,N_13733);
nand UO_1954 (O_1954,N_14304,N_12404);
nor UO_1955 (O_1955,N_13066,N_14524);
nand UO_1956 (O_1956,N_13843,N_13459);
nor UO_1957 (O_1957,N_12627,N_14537);
nand UO_1958 (O_1958,N_12969,N_14559);
nand UO_1959 (O_1959,N_12356,N_12649);
xor UO_1960 (O_1960,N_14799,N_14361);
or UO_1961 (O_1961,N_12095,N_12811);
xor UO_1962 (O_1962,N_12994,N_13986);
and UO_1963 (O_1963,N_14449,N_14026);
and UO_1964 (O_1964,N_12198,N_14603);
and UO_1965 (O_1965,N_14143,N_13516);
and UO_1966 (O_1966,N_14965,N_13318);
nand UO_1967 (O_1967,N_12607,N_13856);
or UO_1968 (O_1968,N_13165,N_13819);
nor UO_1969 (O_1969,N_12992,N_14239);
and UO_1970 (O_1970,N_13021,N_12702);
and UO_1971 (O_1971,N_12051,N_12438);
nand UO_1972 (O_1972,N_13197,N_14875);
nor UO_1973 (O_1973,N_12382,N_12925);
xor UO_1974 (O_1974,N_14597,N_13253);
xnor UO_1975 (O_1975,N_13119,N_14363);
or UO_1976 (O_1976,N_14035,N_14482);
or UO_1977 (O_1977,N_14372,N_14694);
or UO_1978 (O_1978,N_14324,N_12959);
or UO_1979 (O_1979,N_13822,N_12892);
and UO_1980 (O_1980,N_13933,N_13017);
and UO_1981 (O_1981,N_13159,N_13070);
or UO_1982 (O_1982,N_13979,N_14432);
xor UO_1983 (O_1983,N_12008,N_13593);
nor UO_1984 (O_1984,N_13213,N_14432);
and UO_1985 (O_1985,N_12334,N_13569);
nand UO_1986 (O_1986,N_12074,N_12877);
nand UO_1987 (O_1987,N_13376,N_14742);
xor UO_1988 (O_1988,N_13609,N_13045);
nor UO_1989 (O_1989,N_12114,N_13145);
and UO_1990 (O_1990,N_13071,N_14595);
nand UO_1991 (O_1991,N_14513,N_12753);
nor UO_1992 (O_1992,N_13203,N_13542);
xnor UO_1993 (O_1993,N_13236,N_13511);
nor UO_1994 (O_1994,N_13118,N_13745);
nor UO_1995 (O_1995,N_12749,N_14948);
and UO_1996 (O_1996,N_13372,N_13786);
and UO_1997 (O_1997,N_12366,N_12185);
or UO_1998 (O_1998,N_13069,N_12560);
xnor UO_1999 (O_1999,N_14422,N_14853);
endmodule