module basic_2000_20000_2500_100_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1630,In_541);
or U1 (N_1,In_1785,In_1397);
nand U2 (N_2,In_1096,In_1171);
xnor U3 (N_3,In_608,In_822);
and U4 (N_4,In_1586,In_335);
nor U5 (N_5,In_95,In_106);
xor U6 (N_6,In_239,In_1257);
or U7 (N_7,In_752,In_1132);
or U8 (N_8,In_101,In_397);
and U9 (N_9,In_209,In_1428);
nor U10 (N_10,In_1468,In_1381);
nand U11 (N_11,In_1239,In_1002);
nor U12 (N_12,In_845,In_1879);
nand U13 (N_13,In_664,In_78);
or U14 (N_14,In_1702,In_1340);
or U15 (N_15,In_346,In_1991);
nor U16 (N_16,In_735,In_185);
nand U17 (N_17,In_1169,In_1367);
and U18 (N_18,In_1634,In_341);
and U19 (N_19,In_1814,In_1260);
xnor U20 (N_20,In_220,In_1598);
nor U21 (N_21,In_787,In_358);
or U22 (N_22,In_1759,In_1844);
or U23 (N_23,In_1607,In_1271);
and U24 (N_24,In_1626,In_797);
nor U25 (N_25,In_1186,In_287);
and U26 (N_26,In_1677,In_833);
nor U27 (N_27,In_514,In_459);
nand U28 (N_28,In_1195,In_715);
and U29 (N_29,In_372,In_1149);
or U30 (N_30,In_1494,In_469);
and U31 (N_31,In_1400,In_666);
nor U32 (N_32,In_1673,In_1245);
nand U33 (N_33,In_1910,In_1901);
nor U34 (N_34,In_173,In_965);
nor U35 (N_35,In_1867,In_629);
nand U36 (N_36,In_1519,In_981);
or U37 (N_37,In_479,In_1776);
or U38 (N_38,In_677,In_223);
nor U39 (N_39,In_1834,In_1732);
nand U40 (N_40,In_1920,In_943);
or U41 (N_41,In_1520,In_138);
nor U42 (N_42,In_1015,In_1316);
or U43 (N_43,In_758,In_1531);
and U44 (N_44,In_1202,In_1424);
or U45 (N_45,In_1456,In_1800);
or U46 (N_46,In_988,In_1762);
or U47 (N_47,In_750,In_927);
and U48 (N_48,In_1538,In_1401);
nand U49 (N_49,In_1114,In_549);
or U50 (N_50,In_236,In_1018);
nand U51 (N_51,In_1486,In_821);
or U52 (N_52,In_278,In_1031);
and U53 (N_53,In_45,In_1729);
or U54 (N_54,In_1223,In_748);
nand U55 (N_55,In_568,In_799);
nor U56 (N_56,In_1258,In_1939);
or U57 (N_57,In_579,In_763);
nor U58 (N_58,In_958,In_7);
and U59 (N_59,In_391,In_892);
xor U60 (N_60,In_131,In_987);
or U61 (N_61,In_1768,In_643);
nand U62 (N_62,In_540,In_290);
and U63 (N_63,In_1268,In_817);
and U64 (N_64,In_1348,In_1074);
or U65 (N_65,In_2,In_61);
nand U66 (N_66,In_1983,In_1530);
and U67 (N_67,In_996,In_681);
or U68 (N_68,In_575,In_414);
or U69 (N_69,In_733,In_779);
and U70 (N_70,In_1948,In_1698);
nand U71 (N_71,In_1502,In_1619);
and U72 (N_72,In_1063,In_1451);
nand U73 (N_73,In_1453,In_1655);
and U74 (N_74,In_382,In_534);
nor U75 (N_75,In_542,In_77);
nor U76 (N_76,In_1387,In_1292);
and U77 (N_77,In_1029,In_910);
nand U78 (N_78,In_1837,In_1462);
or U79 (N_79,In_1856,In_1086);
or U80 (N_80,In_1294,In_675);
nand U81 (N_81,In_297,In_661);
and U82 (N_82,In_1507,In_591);
nand U83 (N_83,In_350,In_1540);
nand U84 (N_84,In_1515,In_8);
or U85 (N_85,In_234,In_1718);
and U86 (N_86,In_513,In_301);
nand U87 (N_87,In_1252,In_360);
or U88 (N_88,In_499,In_1131);
and U89 (N_89,In_1006,In_1500);
nand U90 (N_90,In_1473,In_1106);
and U91 (N_91,In_1383,In_1909);
or U92 (N_92,In_1229,In_464);
or U93 (N_93,In_977,In_1130);
and U94 (N_94,In_316,In_1148);
and U95 (N_95,In_1284,In_744);
nor U96 (N_96,In_896,In_5);
nor U97 (N_97,In_1172,In_873);
nand U98 (N_98,In_1625,In_581);
nand U99 (N_99,In_921,In_94);
and U100 (N_100,In_1911,In_569);
nor U101 (N_101,In_98,In_1405);
nand U102 (N_102,In_764,In_1232);
nand U103 (N_103,In_67,In_1290);
nand U104 (N_104,In_973,In_231);
nand U105 (N_105,In_1103,In_419);
nand U106 (N_106,In_761,In_1893);
nor U107 (N_107,In_1821,In_1080);
or U108 (N_108,In_130,In_1620);
or U109 (N_109,In_1824,In_1512);
nand U110 (N_110,In_1725,In_145);
or U111 (N_111,In_658,In_1108);
and U112 (N_112,In_1224,In_19);
or U113 (N_113,In_1787,In_1988);
xor U114 (N_114,In_1995,In_445);
or U115 (N_115,In_830,In_1140);
xor U116 (N_116,In_984,In_1863);
nor U117 (N_117,In_908,In_1393);
and U118 (N_118,In_1959,In_858);
nand U119 (N_119,In_644,In_1084);
and U120 (N_120,In_1890,In_10);
and U121 (N_121,In_1918,In_1399);
or U122 (N_122,In_1319,In_125);
or U123 (N_123,In_563,In_1222);
and U124 (N_124,In_322,In_877);
nand U125 (N_125,In_1958,In_928);
or U126 (N_126,In_1237,In_1950);
and U127 (N_127,In_1124,In_637);
and U128 (N_128,In_1402,In_51);
nor U129 (N_129,In_1926,In_398);
nand U130 (N_130,In_34,In_823);
and U131 (N_131,In_1985,In_156);
and U132 (N_132,In_783,In_467);
nand U133 (N_133,In_1555,In_1406);
nor U134 (N_134,In_1973,In_948);
nand U135 (N_135,In_665,In_54);
nor U136 (N_136,In_994,In_1280);
nand U137 (N_137,In_843,In_134);
xor U138 (N_138,In_114,In_555);
nand U139 (N_139,In_1164,In_1354);
nor U140 (N_140,In_711,In_47);
or U141 (N_141,In_1806,In_1788);
and U142 (N_142,In_934,In_1672);
or U143 (N_143,In_451,In_168);
and U144 (N_144,In_814,In_1467);
or U145 (N_145,In_1395,In_481);
nor U146 (N_146,In_1639,In_105);
and U147 (N_147,In_876,In_202);
nor U148 (N_148,In_159,In_1009);
nand U149 (N_149,In_250,In_1437);
and U150 (N_150,In_1209,In_1072);
and U151 (N_151,In_771,In_171);
nand U152 (N_152,In_1150,In_1243);
nand U153 (N_153,In_639,In_816);
or U154 (N_154,In_208,In_1325);
nand U155 (N_155,In_359,In_413);
or U156 (N_156,In_1659,In_191);
nor U157 (N_157,In_756,In_1608);
or U158 (N_158,In_43,In_1509);
and U159 (N_159,In_1060,In_431);
nand U160 (N_160,In_309,In_463);
nand U161 (N_161,In_609,In_1668);
nor U162 (N_162,In_147,In_403);
nand U163 (N_163,In_605,In_1658);
nand U164 (N_164,In_1205,In_536);
or U165 (N_165,In_746,In_1366);
and U166 (N_166,In_1102,In_1079);
nor U167 (N_167,In_1070,In_1621);
nand U168 (N_168,In_1611,In_118);
nor U169 (N_169,In_1735,In_1374);
nor U170 (N_170,In_872,In_76);
and U171 (N_171,In_1219,In_636);
or U172 (N_172,In_190,In_857);
or U173 (N_173,In_1891,In_1059);
or U174 (N_174,In_1194,In_1210);
or U175 (N_175,In_74,In_1177);
and U176 (N_176,In_1618,In_1815);
nand U177 (N_177,In_1728,In_699);
or U178 (N_178,In_1185,In_1795);
and U179 (N_179,In_1804,In_380);
and U180 (N_180,In_150,In_228);
nor U181 (N_181,In_1521,In_641);
nor U182 (N_182,In_23,In_275);
or U183 (N_183,In_1827,In_1256);
nor U184 (N_184,In_357,In_659);
or U185 (N_185,In_1946,In_1749);
or U186 (N_186,In_1727,In_697);
or U187 (N_187,In_604,In_660);
nand U188 (N_188,In_577,In_493);
and U189 (N_189,In_1840,In_172);
nor U190 (N_190,In_1645,In_443);
nand U191 (N_191,In_395,In_1774);
and U192 (N_192,In_539,In_1884);
or U193 (N_193,In_1568,In_251);
and U194 (N_194,In_1792,In_1049);
nor U195 (N_195,In_370,In_84);
xnor U196 (N_196,In_1552,In_570);
or U197 (N_197,In_1127,In_1831);
or U198 (N_198,In_1825,In_645);
or U199 (N_199,In_839,In_1599);
nand U200 (N_200,In_1017,In_650);
and U201 (N_201,In_1105,In_1492);
nand U202 (N_202,In_132,In_1949);
nand U203 (N_203,In_1036,In_361);
or U204 (N_204,In_454,In_772);
and U205 (N_205,In_333,In_442);
or U206 (N_206,In_163,In_158);
and U207 (N_207,In_80,In_798);
nand U208 (N_208,In_351,In_435);
nand U209 (N_209,In_635,In_3);
or U210 (N_210,In_808,In_1694);
or U211 (N_211,In_1001,In_1235);
nor U212 (N_212,In_1297,In_1581);
and U213 (N_213,In_527,In_1802);
nand U214 (N_214,In_1320,In_1123);
or U215 (N_215,In_989,In_1772);
or U216 (N_216,In_649,In_1154);
nor U217 (N_217,In_1892,In_1287);
nor U218 (N_218,In_1999,In_551);
and U219 (N_219,In_1925,In_26);
and U220 (N_220,In_433,In_1485);
xor U221 (N_221,In_1887,In_1046);
or U222 (N_222,In_1967,In_606);
or U223 (N_223,In_938,In_647);
or U224 (N_224,In_1035,In_55);
nand U225 (N_225,In_1529,In_1510);
nor U226 (N_226,N_119,In_71);
nor U227 (N_227,N_107,In_982);
nor U228 (N_228,N_101,In_18);
nor U229 (N_229,In_820,In_62);
or U230 (N_230,In_1037,In_809);
and U231 (N_231,In_1679,In_1833);
and U232 (N_232,In_86,In_450);
or U233 (N_233,In_103,In_269);
and U234 (N_234,N_152,In_1048);
nand U235 (N_235,In_1882,In_714);
and U236 (N_236,In_1778,In_1595);
nand U237 (N_237,In_1656,In_1328);
nand U238 (N_238,In_1438,In_1415);
nor U239 (N_239,In_1162,In_438);
and U240 (N_240,In_1556,In_810);
and U241 (N_241,N_89,In_455);
or U242 (N_242,N_120,In_813);
or U243 (N_243,In_1429,In_627);
nand U244 (N_244,In_1902,In_1764);
or U245 (N_245,In_461,In_1935);
nor U246 (N_246,In_367,N_82);
nand U247 (N_247,In_252,N_74);
and U248 (N_248,In_1466,In_837);
and U249 (N_249,In_586,In_501);
nor U250 (N_250,In_1545,In_851);
and U251 (N_251,In_1577,In_1585);
nand U252 (N_252,In_1589,In_1701);
nand U253 (N_253,In_1767,In_1593);
or U254 (N_254,In_1250,In_1300);
nor U255 (N_255,In_1657,N_57);
and U256 (N_256,In_1972,In_1746);
or U257 (N_257,In_262,In_1769);
and U258 (N_258,In_16,In_716);
nand U259 (N_259,In_276,N_41);
nand U260 (N_260,In_705,In_1365);
xor U261 (N_261,In_751,In_471);
and U262 (N_262,N_18,In_1291);
and U263 (N_263,In_175,In_999);
nand U264 (N_264,In_964,In_932);
nand U265 (N_265,In_60,In_707);
nand U266 (N_266,In_386,In_924);
xnor U267 (N_267,In_972,N_162);
nand U268 (N_268,In_352,In_1092);
nand U269 (N_269,N_8,In_1334);
xnor U270 (N_270,In_1176,In_1550);
and U271 (N_271,In_1347,In_1773);
nor U272 (N_272,In_11,In_1894);
and U273 (N_273,In_1110,In_1261);
nand U274 (N_274,In_79,In_127);
or U275 (N_275,In_1078,In_1028);
nand U276 (N_276,In_911,In_1822);
or U277 (N_277,In_1431,N_182);
nor U278 (N_278,In_573,In_1014);
nor U279 (N_279,In_706,In_1790);
and U280 (N_280,In_1075,In_1541);
nor U281 (N_281,In_1551,In_1081);
or U282 (N_282,In_646,In_14);
nor U283 (N_283,In_1118,N_39);
nand U284 (N_284,In_866,In_504);
nor U285 (N_285,In_1004,In_856);
nand U286 (N_286,In_584,In_1179);
xor U287 (N_287,In_441,In_155);
or U288 (N_288,In_1649,In_292);
nor U289 (N_289,In_1687,N_150);
or U290 (N_290,In_1650,In_1571);
and U291 (N_291,N_46,N_67);
nor U292 (N_292,In_1470,In_951);
nand U293 (N_293,In_1643,In_1396);
and U294 (N_294,N_60,In_28);
or U295 (N_295,In_1754,In_247);
nor U296 (N_296,In_1330,In_780);
or U297 (N_297,In_1628,In_766);
nor U298 (N_298,In_684,In_472);
nor U299 (N_299,N_151,In_1566);
and U300 (N_300,In_562,In_238);
or U301 (N_301,In_1495,In_418);
nand U302 (N_302,In_1146,In_1411);
nand U303 (N_303,In_742,In_1906);
nor U304 (N_304,In_253,In_1434);
and U305 (N_305,In_840,In_421);
xnor U306 (N_306,N_145,In_400);
or U307 (N_307,In_151,In_1722);
or U308 (N_308,In_1267,In_363);
nor U309 (N_309,In_1234,In_387);
and U310 (N_310,In_233,In_546);
and U311 (N_311,In_254,In_407);
nand U312 (N_312,In_941,In_1324);
nand U313 (N_313,In_1269,In_1968);
or U314 (N_314,In_126,In_1253);
nor U315 (N_315,In_529,In_850);
and U316 (N_316,N_187,N_176);
or U317 (N_317,In_805,In_1277);
or U318 (N_318,In_204,In_824);
and U319 (N_319,In_1310,In_1713);
nand U320 (N_320,N_100,In_1524);
nor U321 (N_321,In_997,N_139);
nor U322 (N_322,In_1064,In_887);
or U323 (N_323,In_1314,In_588);
and U324 (N_324,In_523,In_920);
or U325 (N_325,In_1090,In_520);
and U326 (N_326,In_483,In_1823);
nor U327 (N_327,In_1012,In_1984);
nor U328 (N_328,In_1885,In_1613);
nor U329 (N_329,In_82,N_117);
or U330 (N_330,In_1323,In_828);
and U331 (N_331,In_1671,N_128);
or U332 (N_332,In_169,In_841);
or U333 (N_333,In_904,In_1872);
or U334 (N_334,In_267,In_1753);
or U335 (N_335,In_974,N_161);
nor U336 (N_336,In_1737,In_1282);
nand U337 (N_337,In_432,In_258);
or U338 (N_338,In_1733,In_1442);
nand U339 (N_339,In_321,In_871);
and U340 (N_340,In_619,In_1848);
or U341 (N_341,In_640,N_54);
nand U342 (N_342,In_1981,In_257);
or U343 (N_343,In_874,In_1311);
or U344 (N_344,In_1359,In_745);
or U345 (N_345,In_564,In_365);
nand U346 (N_346,In_768,In_289);
or U347 (N_347,In_1189,In_1157);
nor U348 (N_348,In_186,N_129);
or U349 (N_349,In_452,In_364);
and U350 (N_350,In_1716,In_1810);
nand U351 (N_351,In_950,In_325);
nand U352 (N_352,In_491,In_1452);
or U353 (N_353,In_1303,In_1919);
or U354 (N_354,In_1780,In_1609);
nor U355 (N_355,In_1944,In_1862);
and U356 (N_356,In_268,In_189);
and U357 (N_357,N_190,In_1850);
nand U358 (N_358,In_1913,In_437);
nor U359 (N_359,In_362,In_1030);
or U360 (N_360,In_389,In_1859);
nand U361 (N_361,In_486,In_1117);
nor U362 (N_362,In_720,N_155);
nand U363 (N_363,In_1970,N_51);
or U364 (N_364,In_1956,In_1854);
or U365 (N_365,In_1249,In_36);
and U366 (N_366,In_1947,In_1994);
and U367 (N_367,In_535,In_980);
and U368 (N_368,N_188,In_1155);
and U369 (N_369,N_158,In_1663);
and U370 (N_370,In_198,In_1475);
nand U371 (N_371,N_196,In_598);
nor U372 (N_372,In_1992,In_853);
or U373 (N_373,In_332,In_500);
nand U374 (N_374,In_1793,In_1040);
nor U375 (N_375,In_59,In_142);
nor U376 (N_376,In_585,In_1481);
and U377 (N_377,In_543,In_1573);
or U378 (N_378,In_905,N_73);
and U379 (N_379,N_146,In_261);
nor U380 (N_380,N_70,In_1213);
or U381 (N_381,In_1665,In_701);
and U382 (N_382,In_1353,In_693);
or U383 (N_383,In_143,In_473);
and U384 (N_384,In_485,In_1914);
nor U385 (N_385,In_424,In_184);
nor U386 (N_386,In_1198,In_765);
nand U387 (N_387,In_1378,In_1895);
nor U388 (N_388,In_305,In_1580);
or U389 (N_389,N_14,In_696);
nor U390 (N_390,In_49,N_44);
or U391 (N_391,In_770,N_148);
or U392 (N_392,In_1109,In_240);
nand U393 (N_393,In_991,In_274);
nand U394 (N_394,In_1041,N_115);
or U395 (N_395,In_256,In_1880);
nand U396 (N_396,In_1480,In_404);
and U397 (N_397,In_1326,In_1047);
nand U398 (N_398,In_1736,In_891);
nor U399 (N_399,N_53,In_458);
nor U400 (N_400,In_1917,In_32);
and U401 (N_401,In_69,In_248);
nor U402 (N_402,In_408,In_669);
nor U403 (N_403,In_1832,In_201);
and U404 (N_404,In_959,In_1864);
nor U405 (N_405,N_291,In_990);
and U406 (N_406,In_271,In_600);
or U407 (N_407,In_152,In_506);
and U408 (N_408,In_323,In_1794);
or U409 (N_409,In_1610,In_1379);
nor U410 (N_410,In_1459,N_43);
or U411 (N_411,In_197,In_283);
nand U412 (N_412,In_246,In_1924);
nand U413 (N_413,In_1542,In_594);
nand U414 (N_414,In_1062,N_265);
nor U415 (N_415,In_961,N_165);
and U416 (N_416,N_375,In_436);
and U417 (N_417,In_157,N_240);
nor U418 (N_418,In_1458,In_1240);
nor U419 (N_419,In_401,N_102);
or U420 (N_420,In_1380,In_1409);
and U421 (N_421,In_578,In_616);
and U422 (N_422,N_368,In_1457);
or U423 (N_423,In_1254,In_122);
nand U424 (N_424,In_1881,In_496);
nand U425 (N_425,In_1433,In_912);
and U426 (N_426,In_1321,In_819);
and U427 (N_427,In_1389,In_1676);
or U428 (N_428,N_278,In_1940);
or U429 (N_429,N_121,In_1122);
and U430 (N_430,In_614,In_480);
nand U431 (N_431,In_657,In_1648);
nand U432 (N_432,In_495,In_144);
and U433 (N_433,In_762,N_305);
nand U434 (N_434,N_124,In_1624);
xnor U435 (N_435,N_232,In_374);
nor U436 (N_436,N_167,In_468);
nor U437 (N_437,N_11,In_1447);
nand U438 (N_438,In_1283,N_153);
nand U439 (N_439,In_1226,In_213);
xor U440 (N_440,In_1805,N_199);
nor U441 (N_441,In_1067,In_1208);
and U442 (N_442,In_794,N_323);
or U443 (N_443,In_1791,In_430);
and U444 (N_444,N_175,N_326);
nor U445 (N_445,In_834,In_1933);
and U446 (N_446,In_119,In_712);
and U447 (N_447,In_1318,In_176);
nand U448 (N_448,N_104,In_427);
nand U449 (N_449,In_1982,In_516);
nor U450 (N_450,In_1307,In_42);
or U451 (N_451,In_1596,In_153);
or U452 (N_452,In_1465,In_1597);
and U453 (N_453,In_470,N_309);
nor U454 (N_454,N_341,In_1076);
nor U455 (N_455,N_72,In_1135);
or U456 (N_456,N_348,In_167);
or U457 (N_457,In_1747,In_1709);
or U458 (N_458,In_849,In_1045);
nand U459 (N_459,N_353,In_1042);
nor U460 (N_460,In_1770,In_273);
nor U461 (N_461,In_1877,In_538);
or U462 (N_462,In_1697,In_1820);
xnor U463 (N_463,In_709,N_223);
and U464 (N_464,In_1474,In_1178);
nand U465 (N_465,In_453,In_703);
and U466 (N_466,In_825,In_610);
nor U467 (N_467,In_314,N_20);
nand U468 (N_468,In_556,In_955);
nor U469 (N_469,In_651,In_1377);
nand U470 (N_470,In_863,In_914);
nor U471 (N_471,In_1721,In_1191);
nor U472 (N_472,In_796,In_25);
and U473 (N_473,N_332,In_893);
nor U474 (N_474,In_331,In_1777);
and U475 (N_475,In_1055,In_1954);
nand U476 (N_476,In_1761,In_818);
or U477 (N_477,In_216,In_970);
nand U478 (N_478,In_882,N_363);
nand U479 (N_479,N_356,N_242);
nand U480 (N_480,In_1175,In_1033);
nor U481 (N_481,In_1121,N_338);
nor U482 (N_482,In_242,N_380);
nand U483 (N_483,In_1870,In_754);
nand U484 (N_484,In_1289,N_324);
and U485 (N_485,N_198,In_1227);
and U486 (N_486,In_907,In_1505);
nor U487 (N_487,In_327,In_1501);
or U488 (N_488,In_1696,In_1591);
or U489 (N_489,N_225,In_1384);
nand U490 (N_490,In_1765,In_1472);
nand U491 (N_491,In_1816,N_284);
nand U492 (N_492,N_173,In_953);
nand U493 (N_493,N_164,In_329);
nand U494 (N_494,N_47,In_1449);
and U495 (N_495,N_127,In_1071);
or U496 (N_496,N_125,N_255);
nand U497 (N_497,In_1225,In_1786);
nor U498 (N_498,In_426,N_29);
or U499 (N_499,N_234,In_531);
nor U500 (N_500,In_1622,In_655);
nor U501 (N_501,In_1276,In_371);
and U502 (N_502,N_275,In_615);
nor U503 (N_503,In_1508,N_210);
or U504 (N_504,In_356,In_245);
nor U505 (N_505,In_1752,N_194);
nand U506 (N_506,In_1050,In_662);
nor U507 (N_507,In_200,N_214);
and U508 (N_508,In_345,In_1666);
and U509 (N_509,In_638,In_883);
nor U510 (N_510,N_163,N_137);
nand U511 (N_511,In_864,N_71);
xor U512 (N_512,In_505,In_402);
or U513 (N_513,In_1535,In_440);
and U514 (N_514,In_1398,In_1313);
or U515 (N_515,N_247,In_1119);
nand U516 (N_516,In_298,N_241);
nand U517 (N_517,In_717,In_1557);
nand U518 (N_518,In_1532,In_689);
nand U519 (N_519,In_1056,In_1927);
nand U520 (N_520,In_1869,In_694);
nand U521 (N_521,In_1362,In_739);
and U522 (N_522,In_303,In_1522);
xnor U523 (N_523,In_668,In_1514);
nor U524 (N_524,N_52,In_336);
nand U525 (N_525,In_1616,In_889);
or U526 (N_526,In_784,In_83);
and U527 (N_527,In_260,In_1897);
or U528 (N_528,In_1385,In_922);
and U529 (N_529,In_1201,In_1315);
and U530 (N_530,In_1717,N_231);
and U531 (N_531,In_1569,In_592);
nand U532 (N_532,In_1000,N_359);
or U533 (N_533,In_1427,In_1945);
or U534 (N_534,N_149,N_393);
nand U535 (N_535,In_207,N_328);
nor U536 (N_536,In_1027,In_511);
or U537 (N_537,N_157,In_785);
nor U538 (N_538,In_396,In_1011);
or U539 (N_539,In_146,N_147);
nand U540 (N_540,In_1503,In_1170);
nor U541 (N_541,N_343,In_1302);
or U542 (N_542,In_1032,In_117);
xor U543 (N_543,In_1811,In_528);
nor U544 (N_544,In_512,In_944);
and U545 (N_545,In_1196,In_963);
and U546 (N_546,In_1113,In_695);
or U547 (N_547,In_1355,In_1711);
and U548 (N_548,In_1461,In_1426);
and U549 (N_549,In_498,In_1068);
nor U550 (N_550,In_317,In_1372);
nor U551 (N_551,In_1295,In_1104);
nor U552 (N_552,In_465,In_1899);
and U553 (N_553,In_1828,In_618);
or U554 (N_554,In_1734,In_1838);
or U555 (N_555,In_710,In_1);
nand U556 (N_556,In_1497,In_462);
nand U557 (N_557,In_700,N_88);
nor U558 (N_558,In_1511,N_350);
nand U559 (N_559,In_931,In_1866);
and U560 (N_560,In_954,In_1638);
nor U561 (N_561,In_439,In_724);
nand U562 (N_562,N_217,In_0);
and U563 (N_563,In_1144,In_381);
nand U564 (N_564,N_33,In_182);
or U565 (N_565,In_740,In_1489);
nand U566 (N_566,In_1136,N_27);
nor U567 (N_567,In_571,In_313);
or U568 (N_568,In_835,In_196);
nand U569 (N_569,In_63,N_349);
or U570 (N_570,In_1338,N_358);
nand U571 (N_571,In_1707,In_1647);
or U572 (N_572,N_379,In_265);
nor U573 (N_573,In_852,In_590);
or U574 (N_574,In_85,N_220);
or U575 (N_575,In_803,In_148);
and U576 (N_576,In_490,In_867);
and U577 (N_577,In_1703,N_342);
or U578 (N_578,In_1414,In_1560);
nor U579 (N_579,In_1259,In_1900);
and U580 (N_580,In_869,In_792);
or U581 (N_581,In_1231,In_1363);
or U582 (N_582,N_269,In_1100);
and U583 (N_583,In_1375,N_233);
and U584 (N_584,In_1187,In_1953);
nor U585 (N_585,In_1923,In_409);
and U586 (N_586,In_222,N_79);
nand U587 (N_587,In_1670,In_1699);
and U588 (N_588,In_1083,In_879);
nand U589 (N_589,In_737,In_295);
nor U590 (N_590,N_108,In_1874);
nor U591 (N_591,In_679,In_149);
or U592 (N_592,N_31,In_1801);
nor U593 (N_593,In_1477,N_7);
and U594 (N_594,In_1023,In_377);
and U595 (N_595,N_78,In_192);
nand U596 (N_596,In_68,In_1843);
nand U597 (N_597,In_1275,In_894);
or U598 (N_598,In_296,N_281);
or U599 (N_599,N_313,In_164);
or U600 (N_600,N_347,In_1561);
nor U601 (N_601,In_1051,N_544);
nand U602 (N_602,In_956,In_895);
nand U603 (N_603,N_403,N_516);
and U604 (N_604,In_671,In_902);
and U605 (N_605,In_1357,In_755);
or U606 (N_606,In_1069,In_993);
and U607 (N_607,N_301,In_1839);
and U608 (N_608,N_490,In_210);
and U609 (N_609,N_2,In_277);
or U610 (N_610,In_1548,In_211);
nand U611 (N_611,In_1653,In_1279);
and U612 (N_612,In_1962,In_1416);
nor U613 (N_613,In_1116,In_1695);
and U614 (N_614,N_365,N_520);
xnor U615 (N_615,In_854,In_1851);
or U616 (N_616,N_451,In_1021);
nor U617 (N_617,In_1662,In_1640);
and U618 (N_618,In_791,In_625);
nor U619 (N_619,In_1444,In_1460);
nand U620 (N_620,In_1570,In_1174);
nand U621 (N_621,N_81,N_45);
nand U622 (N_622,In_1623,In_942);
nand U623 (N_623,In_384,In_4);
and U624 (N_624,In_1601,In_109);
and U625 (N_625,In_1270,N_538);
and U626 (N_626,In_128,In_812);
or U627 (N_627,In_1455,N_470);
or U628 (N_628,In_865,In_141);
nor U629 (N_629,In_1951,In_1675);
nor U630 (N_630,In_890,In_544);
and U631 (N_631,N_96,In_1682);
nand U632 (N_632,In_1487,In_838);
and U633 (N_633,In_1633,N_25);
and U634 (N_634,N_62,In_1281);
and U635 (N_635,N_545,In_1425);
and U636 (N_636,N_110,In_603);
nand U637 (N_637,In_1479,N_514);
or U638 (N_638,In_1533,In_723);
nor U639 (N_639,In_99,N_540);
nand U640 (N_640,In_782,In_1392);
and U641 (N_641,In_565,In_1197);
nand U642 (N_642,N_503,In_800);
or U643 (N_643,In_354,In_1637);
nand U644 (N_644,In_1139,N_221);
xor U645 (N_645,In_793,In_1039);
or U646 (N_646,In_1305,In_1739);
and U647 (N_647,In_1436,N_589);
xnor U648 (N_648,N_271,In_1293);
and U649 (N_649,In_110,In_92);
and U650 (N_650,N_103,N_351);
nor U651 (N_651,In_221,In_861);
or U652 (N_652,N_197,In_1343);
xnor U653 (N_653,N_436,In_1574);
xor U654 (N_654,In_1886,In_179);
or U655 (N_655,N_106,N_412);
and U656 (N_656,N_473,In_1817);
nand U657 (N_657,In_369,In_1274);
and U658 (N_658,In_460,N_504);
nor U659 (N_659,N_140,In_1674);
and U660 (N_660,N_517,In_998);
or U661 (N_661,N_584,N_366);
nor U662 (N_662,In_1719,N_298);
or U663 (N_663,In_1989,In_180);
nand U664 (N_664,N_448,In_1241);
or U665 (N_665,In_1849,In_340);
nand U666 (N_666,In_1807,In_1680);
nor U667 (N_667,N_591,In_1217);
nand U668 (N_668,In_456,In_102);
nand U669 (N_669,N_170,N_245);
nand U670 (N_670,N_431,In_621);
nor U671 (N_671,N_296,In_1077);
nor U672 (N_672,In_1464,N_572);
and U673 (N_673,N_399,In_1403);
or U674 (N_674,In_967,N_524);
or U675 (N_675,N_26,In_1382);
or U676 (N_676,N_280,In_1088);
nor U677 (N_677,N_295,N_258);
and U678 (N_678,In_1246,In_1797);
nand U679 (N_679,In_760,In_1350);
nand U680 (N_680,In_97,N_534);
and U681 (N_681,N_426,N_249);
and U682 (N_682,In_39,In_1912);
nand U683 (N_683,In_1603,In_13);
nand U684 (N_684,In_747,N_464);
and U685 (N_685,In_328,In_1312);
or U686 (N_686,In_1993,In_342);
or U687 (N_687,In_1147,In_1523);
nor U688 (N_688,In_566,N_415);
nor U689 (N_689,In_1053,In_154);
or U690 (N_690,N_476,In_416);
xnor U691 (N_691,In_1527,N_316);
and U692 (N_692,In_1646,In_1288);
or U693 (N_693,N_282,N_30);
and U694 (N_694,In_1654,N_331);
or U695 (N_695,N_310,N_484);
nor U696 (N_696,In_1730,N_568);
nor U697 (N_697,In_1390,In_916);
nor U698 (N_698,In_1490,In_682);
and U699 (N_699,In_378,In_1339);
nor U700 (N_700,N_533,In_1138);
and U701 (N_701,In_741,In_1008);
nand U702 (N_702,N_582,In_757);
nand U703 (N_703,In_1115,In_249);
nand U704 (N_704,In_1562,N_439);
nor U705 (N_705,In_572,N_248);
and U706 (N_706,N_83,In_975);
and U707 (N_707,N_498,In_1043);
or U708 (N_708,N_92,In_1975);
or U709 (N_709,N_475,N_573);
and U710 (N_710,In_38,In_1847);
and U711 (N_711,In_1756,In_1636);
or U712 (N_712,N_510,In_193);
nor U713 (N_713,N_511,In_1974);
nor U714 (N_714,N_37,In_1941);
nand U715 (N_715,In_617,In_1896);
and U716 (N_716,N_450,In_829);
or U717 (N_717,In_1651,In_1484);
and U718 (N_718,In_1929,In_235);
nor U719 (N_719,In_1093,In_1526);
or U720 (N_720,In_596,In_1921);
nand U721 (N_721,N_477,In_1775);
nand U722 (N_722,In_255,N_435);
or U723 (N_723,In_728,In_347);
or U724 (N_724,In_1141,N_537);
nor U725 (N_725,In_1853,N_222);
or U726 (N_726,In_288,In_1212);
nand U727 (N_727,N_559,N_179);
nor U728 (N_728,N_246,N_553);
and U729 (N_729,In_195,N_525);
and U730 (N_730,N_565,In_778);
nor U731 (N_731,In_1743,N_570);
nor U732 (N_732,In_939,N_394);
xnor U733 (N_733,In_489,N_94);
and U734 (N_734,In_875,N_467);
or U735 (N_735,In_1812,N_409);
and U736 (N_736,In_1584,N_432);
and U737 (N_737,In_702,In_65);
and U738 (N_738,In_1265,N_68);
nor U739 (N_739,In_1151,In_597);
nor U740 (N_740,In_1565,In_1748);
nand U741 (N_741,N_65,N_420);
and U742 (N_742,N_543,N_599);
nand U743 (N_743,In_1760,In_507);
nand U744 (N_744,N_404,N_13);
or U745 (N_745,In_399,In_683);
and U746 (N_746,N_169,N_595);
nand U747 (N_747,N_471,In_170);
xnor U748 (N_748,N_91,N_571);
nor U749 (N_749,In_1868,In_96);
nor U750 (N_750,In_1128,In_475);
and U751 (N_751,In_1835,In_214);
or U752 (N_752,N_77,In_1873);
nor U753 (N_753,N_508,N_122);
and U754 (N_754,In_1905,In_123);
and U755 (N_755,N_362,In_1547);
nand U756 (N_756,N_178,In_1327);
nand U757 (N_757,N_262,N_209);
nand U758 (N_758,In_521,N_277);
nand U759 (N_759,N_302,N_21);
nand U760 (N_760,In_530,In_1642);
nor U761 (N_761,N_99,In_1726);
nor U762 (N_762,In_1855,In_429);
nor U763 (N_763,In_1308,N_130);
and U764 (N_764,In_1528,In_722);
nor U765 (N_765,N_93,In_140);
and U766 (N_766,In_1606,N_335);
nor U767 (N_767,In_1052,In_1129);
nand U768 (N_768,In_686,In_919);
nand U769 (N_769,In_1356,In_901);
or U770 (N_770,N_228,In_781);
and U771 (N_771,In_379,In_1809);
and U772 (N_772,In_1738,N_300);
xnor U773 (N_773,N_315,In_48);
nor U774 (N_774,In_1543,N_352);
and U775 (N_775,In_870,In_224);
nand U776 (N_776,In_930,N_42);
or U777 (N_777,In_878,In_1476);
nand U778 (N_778,In_244,In_936);
or U779 (N_779,In_1783,N_274);
nand U780 (N_780,In_81,In_1808);
and U781 (N_781,N_268,In_264);
or U782 (N_782,N_49,N_132);
nor U783 (N_783,In_1038,N_413);
and U784 (N_784,In_1044,N_15);
nand U785 (N_785,In_583,N_141);
and U786 (N_786,In_133,In_1107);
and U787 (N_787,In_420,N_482);
nand U788 (N_788,In_1979,In_915);
nand U789 (N_789,In_1635,In_282);
nor U790 (N_790,In_962,In_1134);
and U791 (N_791,N_17,In_917);
nor U792 (N_792,In_1142,In_1391);
nor U793 (N_793,N_433,N_138);
nand U794 (N_794,In_1394,N_374);
and U795 (N_795,N_590,In_612);
or U796 (N_796,N_286,N_384);
nor U797 (N_797,In_1483,In_1026);
nand U798 (N_798,N_509,In_1563);
or U799 (N_799,In_428,In_1705);
and U800 (N_800,In_1861,N_727);
nand U801 (N_801,In_1161,N_586);
nand U802 (N_802,N_670,In_1333);
or U803 (N_803,N_126,N_105);
nor U804 (N_804,N_397,In_183);
nand U805 (N_805,N_86,N_779);
nand U806 (N_806,N_700,In_1364);
or U807 (N_807,N_613,N_698);
nand U808 (N_808,N_658,N_48);
or U809 (N_809,In_1741,N_769);
and U810 (N_810,N_758,In_553);
nand U811 (N_811,In_926,N_648);
or U812 (N_812,N_741,In_444);
nor U813 (N_813,In_1990,In_135);
and U814 (N_814,In_992,N_34);
nand U815 (N_815,In_492,In_626);
nand U816 (N_816,N_377,N_705);
nor U817 (N_817,N_391,N_547);
or U818 (N_818,In_1661,N_765);
nand U819 (N_819,In_124,N_226);
nand U820 (N_820,In_1536,In_1567);
and U821 (N_821,In_1410,In_56);
nor U822 (N_822,N_123,In_1857);
and U823 (N_823,In_558,N_427);
nor U824 (N_824,In_1054,In_663);
and U825 (N_825,N_364,In_995);
or U826 (N_826,N_483,In_1617);
nand U827 (N_827,N_684,In_1836);
and U828 (N_828,In_1715,N_755);
nand U829 (N_829,In_50,N_405);
or U830 (N_830,In_226,In_482);
and U831 (N_831,N_457,In_383);
nor U832 (N_832,In_339,In_836);
and U833 (N_833,N_402,In_1594);
nor U834 (N_834,N_723,In_53);
nand U835 (N_835,In_749,N_774);
nand U836 (N_836,N_600,In_862);
nor U837 (N_837,In_692,N_395);
and U838 (N_838,In_1221,In_1095);
or U839 (N_839,N_257,In_1331);
nand U840 (N_840,N_729,In_162);
and U841 (N_841,N_263,In_804);
nand U842 (N_842,In_1057,In_1684);
xnor U843 (N_843,In_795,In_826);
nor U844 (N_844,In_1798,In_1430);
nand U845 (N_845,In_687,In_1299);
and U846 (N_846,N_781,In_497);
and U847 (N_847,In_1669,In_1192);
nand U848 (N_848,N_677,In_1034);
or U849 (N_849,N_634,In_1322);
nor U850 (N_850,N_206,N_116);
nor U851 (N_851,N_244,In_30);
or U852 (N_852,In_1263,N_777);
or U853 (N_853,N_761,In_93);
or U854 (N_854,N_685,N_576);
nand U855 (N_855,In_1539,In_1098);
or U856 (N_856,In_1143,In_759);
or U857 (N_857,In_1700,N_501);
nor U858 (N_858,In_1504,N_782);
nand U859 (N_859,N_763,N_493);
nor U860 (N_860,N_75,N_760);
or U861 (N_861,N_676,In_1755);
and U862 (N_862,In_104,N_250);
or U863 (N_863,In_580,In_1407);
or U864 (N_864,N_487,In_1214);
nor U865 (N_865,N_339,In_1332);
nor U866 (N_866,In_9,N_61);
nor U867 (N_867,In_355,In_1386);
and U868 (N_868,N_479,In_1211);
nor U869 (N_869,N_791,N_458);
nand U870 (N_870,N_449,N_160);
or U871 (N_871,In_676,N_715);
and U872 (N_872,N_494,In_393);
or U873 (N_873,N_583,In_1644);
nand U874 (N_874,In_634,In_1010);
or U875 (N_875,In_1066,In_900);
or U876 (N_876,N_767,In_574);
nand U877 (N_877,In_807,In_1204);
nand U878 (N_878,In_726,In_654);
and U879 (N_879,N_647,N_400);
and U880 (N_880,N_645,In_1200);
or U881 (N_881,N_787,In_753);
nand U882 (N_882,In_337,In_227);
and U883 (N_883,In_1830,In_1513);
or U884 (N_884,N_653,N_707);
or U885 (N_885,In_129,In_1306);
or U886 (N_886,In_1976,N_6);
and U887 (N_887,N_492,N_489);
and U888 (N_888,In_1085,In_1614);
and U889 (N_889,N_609,In_215);
nor U890 (N_890,In_1720,In_1163);
nand U891 (N_891,N_603,In_674);
or U892 (N_892,In_503,N_505);
nor U893 (N_893,In_27,N_211);
and U894 (N_894,In_630,N_691);
nand U895 (N_895,N_293,N_76);
xor U896 (N_896,In_1971,In_937);
and U897 (N_897,In_786,In_1525);
nor U898 (N_898,In_422,In_21);
nor U899 (N_899,In_1724,N_632);
and U900 (N_900,In_212,In_623);
nand U901 (N_901,In_1439,In_933);
or U902 (N_902,N_771,N_340);
and U903 (N_903,N_621,N_229);
or U904 (N_904,In_1206,In_57);
and U905 (N_905,N_181,N_444);
nand U906 (N_906,In_731,N_58);
nand U907 (N_907,In_353,N_396);
and U908 (N_908,In_1578,In_1242);
nand U909 (N_909,N_683,N_264);
or U910 (N_910,In_70,In_22);
nor U911 (N_911,In_1714,In_971);
nor U912 (N_912,In_673,In_734);
nand U913 (N_913,N_706,N_243);
or U914 (N_914,N_652,N_614);
nor U915 (N_915,N_114,In_165);
nor U916 (N_916,N_496,In_115);
nor U917 (N_917,In_1168,In_1153);
or U918 (N_918,N_557,In_1368);
nor U919 (N_919,N_183,In_940);
xor U920 (N_920,In_1420,N_193);
or U921 (N_921,N_361,In_308);
nor U922 (N_922,In_690,N_721);
or U923 (N_923,In_1518,In_672);
or U924 (N_924,N_682,In_326);
or U925 (N_925,N_798,N_109);
nor U926 (N_926,In_166,N_797);
or U927 (N_927,In_935,In_366);
or U928 (N_928,N_527,In_1493);
and U929 (N_929,N_354,In_1549);
and U930 (N_930,In_1099,In_1238);
and U931 (N_931,In_1517,In_136);
and U932 (N_932,In_1579,In_1352);
nor U933 (N_933,N_292,In_1228);
nand U934 (N_934,N_689,In_774);
nor U935 (N_935,In_1789,N_306);
nor U936 (N_936,In_802,N_423);
or U937 (N_937,N_97,In_1097);
nor U938 (N_938,In_310,N_334);
nor U939 (N_939,In_1564,N_50);
and U940 (N_940,In_776,In_1193);
or U941 (N_941,In_1781,In_1904);
or U942 (N_942,In_37,In_1966);
nand U943 (N_943,In_302,N_468);
nor U944 (N_944,N_135,In_1329);
nand U945 (N_945,In_537,In_1842);
nand U946 (N_946,In_727,N_549);
and U947 (N_947,In_1019,In_1693);
or U948 (N_948,N_486,N_261);
and U949 (N_949,N_131,N_693);
nor U950 (N_950,N_768,In_846);
or U951 (N_951,In_811,N_333);
or U952 (N_952,In_1344,In_1448);
xor U953 (N_953,In_187,In_1845);
nor U954 (N_954,N_757,N_642);
nor U955 (N_955,In_1987,In_203);
and U956 (N_956,N_12,In_494);
and U957 (N_957,N_500,In_788);
or U958 (N_958,N_239,N_657);
nor U959 (N_959,In_1337,N_154);
and U960 (N_960,In_449,In_622);
and U961 (N_961,In_1898,N_610);
nand U962 (N_962,N_9,In_898);
or U963 (N_963,In_111,N_453);
nor U964 (N_964,In_1089,In_518);
nor U965 (N_965,In_139,In_72);
nor U966 (N_966,In_1692,In_1446);
nand U967 (N_967,In_1137,In_334);
or U968 (N_968,N_546,N_216);
and U969 (N_969,N_536,N_355);
nor U970 (N_970,In_587,In_888);
or U971 (N_971,N_203,N_795);
nand U972 (N_972,In_652,N_98);
nor U973 (N_973,In_1930,N_32);
nor U974 (N_974,N_478,N_376);
and U975 (N_975,N_208,In_285);
and U976 (N_976,In_1218,In_338);
or U977 (N_977,N_722,In_903);
or U978 (N_978,N_608,N_637);
nor U979 (N_979,N_407,N_307);
or U980 (N_980,In_300,In_1683);
and U981 (N_981,In_1370,In_729);
and U982 (N_982,N_668,In_1005);
xor U983 (N_983,N_474,In_1846);
or U984 (N_984,N_620,In_487);
nor U985 (N_985,N_133,In_1445);
or U986 (N_986,In_1203,In_199);
nand U987 (N_987,In_949,In_1373);
nand U988 (N_988,N_789,In_1615);
nand U989 (N_989,In_488,N_273);
nand U990 (N_990,In_160,In_502);
and U991 (N_991,N_236,In_1943);
or U992 (N_992,In_1627,N_535);
nor U993 (N_993,In_17,In_293);
nor U994 (N_994,In_304,N_523);
xnor U995 (N_995,N_564,In_1986);
nor U996 (N_996,In_946,N_134);
and U997 (N_997,N_177,N_437);
or U998 (N_998,In_218,In_548);
nor U999 (N_999,In_1928,N_502);
or U1000 (N_1000,N_731,N_419);
or U1001 (N_1001,N_674,N_136);
and U1002 (N_1002,In_1558,N_687);
nand U1003 (N_1003,N_806,In_1860);
nand U1004 (N_1004,N_252,N_678);
or U1005 (N_1005,N_974,In_1423);
nand U1006 (N_1006,In_161,N_311);
or U1007 (N_1007,N_429,N_702);
nand U1008 (N_1008,N_971,N_174);
nor U1009 (N_1009,In_1082,In_1852);
nor U1010 (N_1010,N_461,In_1706);
nor U1011 (N_1011,In_827,In_789);
nand U1012 (N_1012,N_842,N_605);
nand U1013 (N_1013,In_1158,In_519);
and U1014 (N_1014,N_699,N_909);
or U1015 (N_1015,In_1916,In_561);
and U1016 (N_1016,In_685,In_969);
or U1017 (N_1017,In_509,N_981);
and U1018 (N_1018,In_1199,N_515);
and U1019 (N_1019,N_709,In_842);
nor U1020 (N_1020,In_704,In_522);
and U1021 (N_1021,N_919,N_601);
nor U1022 (N_1022,In_1588,N_770);
nand U1023 (N_1023,In_1272,In_1602);
nand U1024 (N_1024,In_1922,N_863);
nand U1025 (N_1025,N_550,N_751);
nor U1026 (N_1026,In_552,N_562);
or U1027 (N_1027,N_443,N_597);
and U1028 (N_1028,N_911,N_378);
xnor U1029 (N_1029,N_66,N_788);
and U1030 (N_1030,In_595,In_976);
nor U1031 (N_1031,In_1181,N_408);
or U1032 (N_1032,In_1216,In_790);
or U1033 (N_1033,N_784,In_1742);
nand U1034 (N_1034,N_24,In_1803);
or U1035 (N_1035,In_1750,N_688);
nand U1036 (N_1036,In_721,N_993);
or U1037 (N_1037,N_987,N_285);
and U1038 (N_1038,In_478,In_613);
and U1039 (N_1039,N_884,N_626);
or U1040 (N_1040,N_587,N_38);
nand U1041 (N_1041,In_547,N_895);
nor U1042 (N_1042,N_737,In_434);
or U1043 (N_1043,In_599,In_1758);
nand U1044 (N_1044,In_860,In_1419);
nor U1045 (N_1045,N_977,N_695);
nor U1046 (N_1046,In_1779,N_734);
or U1047 (N_1047,In_667,In_1813);
or U1048 (N_1048,N_80,N_186);
nand U1049 (N_1049,In_64,In_557);
nand U1050 (N_1050,N_881,N_907);
or U1051 (N_1051,N_878,N_485);
nor U1052 (N_1052,In_945,N_932);
nor U1053 (N_1053,N_360,In_1546);
and U1054 (N_1054,In_1952,In_263);
nand U1055 (N_1055,In_1369,N_762);
nand U1056 (N_1056,N_838,In_691);
xnor U1057 (N_1057,N_299,N_991);
and U1058 (N_1058,In_1678,N_852);
and U1059 (N_1059,N_808,In_1771);
nand U1060 (N_1060,N_998,In_1304);
nor U1061 (N_1061,In_550,N_816);
or U1062 (N_1062,N_434,N_965);
and U1063 (N_1063,N_36,N_764);
nand U1064 (N_1064,N_866,In_1600);
nor U1065 (N_1065,In_91,N_713);
and U1066 (N_1066,In_1681,N_656);
or U1067 (N_1067,N_792,N_606);
and U1068 (N_1068,N_818,In_1183);
nor U1069 (N_1069,In_1544,N_639);
nor U1070 (N_1070,In_410,N_267);
and U1071 (N_1071,N_171,N_872);
nand U1072 (N_1072,N_959,In_1418);
and U1073 (N_1073,N_594,N_390);
nand U1074 (N_1074,N_55,In_1604);
or U1075 (N_1075,N_980,In_1301);
nor U1076 (N_1076,In_1977,N_819);
or U1077 (N_1077,N_95,In_601);
nor U1078 (N_1078,N_555,N_386);
nand U1079 (N_1079,N_703,In_237);
nor U1080 (N_1080,In_1182,In_855);
nand U1081 (N_1081,N_710,In_412);
nand U1082 (N_1082,N_628,N_815);
nand U1083 (N_1083,N_747,N_994);
nor U1084 (N_1084,N_899,In_1262);
nand U1085 (N_1085,N_22,In_1125);
or U1086 (N_1086,N_480,In_719);
or U1087 (N_1087,N_833,In_266);
nand U1088 (N_1088,N_783,N_195);
or U1089 (N_1089,N_840,N_541);
nand U1090 (N_1090,N_69,N_739);
nor U1091 (N_1091,In_1858,N_716);
or U1092 (N_1092,N_297,In_678);
nor U1093 (N_1093,N_805,N_924);
or U1094 (N_1094,In_848,In_1180);
or U1095 (N_1095,In_229,N_513);
nand U1096 (N_1096,In_526,N_933);
nand U1097 (N_1097,N_166,In_1413);
nand U1098 (N_1098,N_949,In_1016);
and U1099 (N_1099,N_931,N_619);
or U1100 (N_1100,In_1230,N_469);
nand U1101 (N_1101,N_387,N_389);
or U1102 (N_1102,N_327,In_1592);
or U1103 (N_1103,In_1996,N_465);
or U1104 (N_1104,In_801,In_1317);
and U1105 (N_1105,In_633,In_1576);
nand U1106 (N_1106,N_191,In_324);
and U1107 (N_1107,In_307,In_1482);
nand U1108 (N_1108,N_577,N_772);
nor U1109 (N_1109,In_567,In_1932);
or U1110 (N_1110,N_847,In_1435);
or U1111 (N_1111,N_714,In_344);
or U1112 (N_1112,N_927,N_943);
nor U1113 (N_1113,N_854,In_1744);
and U1114 (N_1114,In_1091,In_1961);
or U1115 (N_1115,N_383,In_24);
nand U1116 (N_1116,N_425,N_839);
nand U1117 (N_1117,N_690,In_670);
or U1118 (N_1118,In_315,In_100);
nor U1119 (N_1119,In_405,N_585);
nor U1120 (N_1120,In_385,In_1454);
and U1121 (N_1121,In_767,N_172);
and U1122 (N_1122,In_1233,N_753);
or U1123 (N_1123,In_280,In_390);
nor U1124 (N_1124,N_902,In_736);
nand U1125 (N_1125,N_660,N_865);
or U1126 (N_1126,In_1432,In_628);
or U1127 (N_1127,In_885,N_629);
nor U1128 (N_1128,N_113,In_1112);
or U1129 (N_1129,In_40,N_518);
nand U1130 (N_1130,N_596,In_1931);
and U1131 (N_1131,N_317,N_832);
nor U1132 (N_1132,In_1553,N_883);
and U1133 (N_1133,In_525,In_312);
nor U1134 (N_1134,N_917,N_914);
or U1135 (N_1135,N_424,In_1003);
nand U1136 (N_1136,N_205,N_922);
or U1137 (N_1137,In_219,N_845);
or U1138 (N_1138,In_1516,In_1156);
nand U1139 (N_1139,In_1660,N_851);
or U1140 (N_1140,N_889,In_631);
and U1141 (N_1141,In_582,N_900);
xnor U1142 (N_1142,N_521,N_942);
nand U1143 (N_1143,In_1796,In_1818);
and U1144 (N_1144,In_1799,N_111);
nor U1145 (N_1145,N_958,In_66);
and U1146 (N_1146,In_1740,In_1938);
and U1147 (N_1147,N_843,N_976);
or U1148 (N_1148,N_960,N_717);
and U1149 (N_1149,In_1871,N_891);
nand U1150 (N_1150,N_679,N_823);
nor U1151 (N_1151,In_406,N_921);
nand U1152 (N_1152,N_624,N_827);
nor U1153 (N_1153,In_1488,N_256);
or U1154 (N_1154,N_995,In_205);
nand U1155 (N_1155,N_935,N_488);
or U1156 (N_1156,In_730,N_802);
nand U1157 (N_1157,In_44,N_853);
or U1158 (N_1158,N_370,In_217);
and U1159 (N_1159,N_314,In_899);
nand U1160 (N_1160,In_291,In_1960);
or U1161 (N_1161,N_858,N_112);
and U1162 (N_1162,N_598,In_648);
nand U1163 (N_1163,N_5,N_266);
nand U1164 (N_1164,N_617,N_681);
nor U1165 (N_1165,N_367,In_1471);
and U1166 (N_1166,N_817,In_1371);
or U1167 (N_1167,N_692,N_661);
or U1168 (N_1168,N_822,N_957);
nand U1169 (N_1169,N_979,In_844);
nand U1170 (N_1170,N_901,N_440);
nand U1171 (N_1171,In_968,In_1534);
or U1172 (N_1172,In_286,N_201);
and U1173 (N_1173,In_206,In_1207);
nor U1174 (N_1174,N_336,In_1763);
and U1175 (N_1175,In_602,In_121);
xnor U1176 (N_1176,In_775,N_877);
nor U1177 (N_1177,In_1145,In_1266);
nor U1178 (N_1178,N_807,In_1248);
nor U1179 (N_1179,N_983,In_732);
or U1180 (N_1180,N_322,In_368);
nor U1181 (N_1181,N_497,N_904);
nor U1182 (N_1182,In_376,N_227);
nor U1183 (N_1183,N_812,N_906);
nor U1184 (N_1184,In_1165,N_946);
or U1185 (N_1185,N_887,N_320);
nand U1186 (N_1186,N_430,In_624);
or U1187 (N_1187,N_118,In_446);
nor U1188 (N_1188,In_15,In_985);
nor U1189 (N_1189,N_580,In_457);
or U1190 (N_1190,N_283,N_566);
or U1191 (N_1191,N_144,N_955);
and U1192 (N_1192,N_578,N_903);
or U1193 (N_1193,In_1463,N_40);
nor U1194 (N_1194,In_1590,N_953);
nor U1195 (N_1195,In_725,N_539);
or U1196 (N_1196,N_251,N_659);
and U1197 (N_1197,N_748,In_1689);
nand U1198 (N_1198,N_841,N_913);
and U1199 (N_1199,N_143,N_766);
nand U1200 (N_1200,N_665,N_874);
nor U1201 (N_1201,N_1136,N_1109);
nor U1202 (N_1202,N_720,In_1273);
nor U1203 (N_1203,N_844,N_1196);
nor U1204 (N_1204,N_1043,In_1688);
and U1205 (N_1205,N_219,In_1980);
or U1206 (N_1206,In_1712,N_1019);
nand U1207 (N_1207,N_398,N_588);
and U1208 (N_1208,N_622,N_759);
and U1209 (N_1209,In_847,N_615);
nand U1210 (N_1210,N_918,N_371);
nand U1211 (N_1211,In_73,N_871);
or U1212 (N_1212,N_1000,N_507);
and U1213 (N_1213,N_1194,N_1147);
nand U1214 (N_1214,In_517,N_230);
nand U1215 (N_1215,N_785,In_1309);
nor U1216 (N_1216,In_1013,N_649);
nand U1217 (N_1217,N_466,N_1135);
or U1218 (N_1218,N_1182,N_581);
nand U1219 (N_1219,N_875,N_592);
and U1220 (N_1220,In_1360,N_969);
nand U1221 (N_1221,In_1412,N_1016);
and U1222 (N_1222,N_732,In_35);
nor U1223 (N_1223,N_421,N_575);
nand U1224 (N_1224,N_238,N_928);
nor U1225 (N_1225,In_1358,N_1008);
nor U1226 (N_1226,N_663,In_952);
nand U1227 (N_1227,N_631,In_230);
xor U1228 (N_1228,In_713,N_1118);
and U1229 (N_1229,N_1139,N_1150);
or U1230 (N_1230,N_567,In_279);
nor U1231 (N_1231,N_694,N_529);
or U1232 (N_1232,N_625,N_1005);
or U1233 (N_1233,In_656,N_159);
and U1234 (N_1234,N_930,N_775);
and U1235 (N_1235,N_743,In_1101);
nand U1236 (N_1236,N_1112,N_406);
nor U1237 (N_1237,N_1103,N_460);
and U1238 (N_1238,N_1012,N_825);
or U1239 (N_1239,N_898,In_1915);
or U1240 (N_1240,N_1187,N_63);
and U1241 (N_1241,N_934,N_481);
nand U1242 (N_1242,In_284,N_811);
nand U1243 (N_1243,N_992,In_688);
nand U1244 (N_1244,In_394,In_137);
nor U1245 (N_1245,N_1041,N_1038);
nor U1246 (N_1246,N_290,In_815);
nor U1247 (N_1247,N_654,In_89);
nor U1248 (N_1248,N_1188,N_259);
or U1249 (N_1249,N_1079,N_990);
or U1250 (N_1250,N_373,In_447);
nand U1251 (N_1251,In_957,N_1002);
and U1252 (N_1252,In_1691,N_23);
nor U1253 (N_1253,N_950,N_1031);
and U1254 (N_1254,N_560,In_589);
or U1255 (N_1255,N_1145,N_1124);
nand U1256 (N_1256,N_452,N_321);
or U1257 (N_1257,In_1955,N_963);
and U1258 (N_1258,N_711,N_855);
or U1259 (N_1259,N_1048,In_1341);
and U1260 (N_1260,N_319,N_410);
nor U1261 (N_1261,N_260,N_1160);
and U1262 (N_1262,In_881,In_1704);
or U1263 (N_1263,N_1144,N_204);
and U1264 (N_1264,N_185,In_923);
nand U1265 (N_1265,In_75,In_642);
nor U1266 (N_1266,In_1286,In_1907);
or U1267 (N_1267,N_558,In_1336);
nor U1268 (N_1268,In_593,N_604);
nor U1269 (N_1269,N_1141,N_735);
and U1270 (N_1270,N_530,N_985);
xnor U1271 (N_1271,In_906,N_411);
or U1272 (N_1272,N_422,N_686);
nand U1273 (N_1273,N_1023,In_1408);
nand U1274 (N_1274,N_1007,In_194);
or U1275 (N_1275,N_1026,In_177);
nor U1276 (N_1276,N_1064,In_1641);
nand U1277 (N_1277,N_1137,In_1255);
or U1278 (N_1278,In_1478,In_1506);
nor U1279 (N_1279,N_279,N_641);
and U1280 (N_1280,In_1058,N_801);
nor U1281 (N_1281,N_1100,In_1188);
nor U1282 (N_1282,N_1131,N_728);
or U1283 (N_1283,In_979,In_1664);
or U1284 (N_1284,N_1125,N_870);
and U1285 (N_1285,N_1123,In_1605);
nor U1286 (N_1286,N_392,N_849);
nor U1287 (N_1287,In_1903,N_790);
nor U1288 (N_1288,N_738,N_207);
and U1289 (N_1289,N_941,N_1003);
nand U1290 (N_1290,N_1069,N_1163);
nor U1291 (N_1291,In_1024,In_576);
and U1292 (N_1292,In_88,N_385);
and U1293 (N_1293,In_1889,N_554);
nor U1294 (N_1294,In_806,In_1883);
nor U1295 (N_1295,N_1025,N_929);
and U1296 (N_1296,In_1361,In_868);
nor U1297 (N_1297,N_19,N_1099);
xor U1298 (N_1298,N_876,In_232);
nor U1299 (N_1299,In_320,In_31);
and U1300 (N_1300,In_1346,N_1022);
xnor U1301 (N_1301,N_462,N_719);
nor U1302 (N_1302,In_1167,N_499);
nand U1303 (N_1303,In_1166,N_304);
and U1304 (N_1304,N_1053,In_417);
or U1305 (N_1305,N_1181,In_1978);
and U1306 (N_1306,In_1498,In_1934);
nor U1307 (N_1307,N_1162,N_1128);
nand U1308 (N_1308,In_831,N_701);
or U1309 (N_1309,In_620,N_218);
or U1310 (N_1310,N_84,N_1127);
and U1311 (N_1311,In_1629,In_1685);
or U1312 (N_1312,N_1120,N_671);
nand U1313 (N_1313,In_1583,In_1296);
and U1314 (N_1314,N_526,N_754);
nor U1315 (N_1315,In_1215,In_1007);
nand U1316 (N_1316,N_837,N_947);
or U1317 (N_1317,N_633,In_1686);
nor U1318 (N_1318,N_736,N_879);
nand U1319 (N_1319,In_1667,N_1115);
nor U1320 (N_1320,N_846,N_1178);
or U1321 (N_1321,N_1046,N_1104);
nor U1322 (N_1322,In_1757,In_1417);
and U1323 (N_1323,N_542,In_1491);
nand U1324 (N_1324,N_531,In_1875);
or U1325 (N_1325,N_646,In_1690);
nand U1326 (N_1326,N_1085,N_1094);
nor U1327 (N_1327,N_1082,N_416);
nor U1328 (N_1328,N_16,In_484);
or U1329 (N_1329,N_1070,N_1143);
nand U1330 (N_1330,N_1020,N_1017);
and U1331 (N_1331,N_1186,N_1006);
nor U1332 (N_1332,N_644,In_1936);
nand U1333 (N_1333,N_1074,N_836);
xnor U1334 (N_1334,In_1587,In_978);
or U1335 (N_1335,In_859,In_1878);
and U1336 (N_1336,In_1499,N_744);
or U1337 (N_1337,N_1197,N_90);
nor U1338 (N_1338,In_1349,In_225);
nand U1339 (N_1339,In_1025,In_1582);
and U1340 (N_1340,N_857,N_1170);
or U1341 (N_1341,In_1965,N_794);
and U1342 (N_1342,N_1152,In_343);
nor U1343 (N_1343,In_33,N_569);
nor U1344 (N_1344,N_1174,N_940);
or U1345 (N_1345,N_786,N_289);
or U1346 (N_1346,N_616,N_312);
or U1347 (N_1347,N_456,N_669);
and U1348 (N_1348,N_1151,In_1251);
nand U1349 (N_1349,N_202,In_1120);
and U1350 (N_1350,In_1631,In_777);
and U1351 (N_1351,N_1198,In_1559);
nand U1352 (N_1352,N_778,N_799);
xnor U1353 (N_1353,N_912,N_447);
nand U1354 (N_1354,N_988,In_423);
and U1355 (N_1355,In_108,N_607);
nor U1356 (N_1356,In_348,In_1963);
or U1357 (N_1357,N_1040,In_559);
nor U1358 (N_1358,N_1096,N_551);
xor U1359 (N_1359,N_1062,N_856);
nand U1360 (N_1360,N_897,N_1033);
nand U1361 (N_1361,N_873,In_560);
and U1362 (N_1362,N_612,N_1158);
nor U1363 (N_1363,In_1073,In_1632);
nand U1364 (N_1364,N_664,N_967);
nor U1365 (N_1365,N_10,N_1172);
nor U1366 (N_1366,N_1190,N_829);
nor U1367 (N_1367,N_381,N_886);
nor U1368 (N_1368,N_35,In_1094);
and U1369 (N_1369,N_552,N_1034);
and U1370 (N_1370,N_962,N_3);
nand U1371 (N_1371,N_1078,In_425);
nor U1372 (N_1372,N_997,In_1841);
nand U1373 (N_1373,N_1138,N_1180);
nand U1374 (N_1374,N_809,N_1075);
and U1375 (N_1375,N_978,N_442);
or U1376 (N_1376,N_1156,N_1076);
and U1377 (N_1377,N_372,N_1129);
nand U1378 (N_1378,In_116,N_813);
or U1379 (N_1379,N_253,In_1133);
nand U1380 (N_1380,In_1537,N_1047);
nand U1381 (N_1381,N_696,N_1155);
nand U1382 (N_1382,In_1723,N_495);
or U1383 (N_1383,In_174,N_189);
nor U1384 (N_1384,N_956,In_1554);
nand U1385 (N_1385,N_1189,N_618);
nor U1386 (N_1386,N_1121,In_1422);
or U1387 (N_1387,In_983,N_1061);
and U1388 (N_1388,In_1298,In_1342);
nor U1389 (N_1389,In_1450,In_270);
and U1390 (N_1390,N_330,In_880);
and U1391 (N_1391,In_272,N_1199);
and U1392 (N_1392,N_733,N_1166);
nand U1393 (N_1393,In_607,In_947);
and U1394 (N_1394,In_474,In_188);
and U1395 (N_1395,N_1030,N_506);
and U1396 (N_1396,N_1195,N_672);
nand U1397 (N_1397,In_1335,N_1119);
or U1398 (N_1398,N_563,N_905);
nand U1399 (N_1399,N_445,N_984);
nand U1400 (N_1400,N_1130,N_1014);
nand U1401 (N_1401,N_1175,In_319);
and U1402 (N_1402,N_1091,In_913);
nor U1403 (N_1403,In_178,N_1126);
nor U1404 (N_1404,N_357,N_1263);
or U1405 (N_1405,N_308,N_1208);
or U1406 (N_1406,N_1376,N_1036);
and U1407 (N_1407,N_1290,In_1745);
nor U1408 (N_1408,N_752,N_892);
nor U1409 (N_1409,N_643,N_1185);
nand U1410 (N_1410,N_1060,N_1202);
nor U1411 (N_1411,N_519,N_1146);
and U1412 (N_1412,N_1307,In_510);
nor U1413 (N_1413,N_1207,N_1148);
and U1414 (N_1414,N_1057,N_1374);
or U1415 (N_1415,N_1311,N_1159);
or U1416 (N_1416,N_1359,N_294);
nand U1417 (N_1417,N_925,N_288);
nand U1418 (N_1418,N_1092,N_1279);
or U1419 (N_1419,N_1191,In_1160);
and U1420 (N_1420,N_666,N_1366);
and U1421 (N_1421,N_1122,In_1731);
and U1422 (N_1422,N_746,N_556);
or U1423 (N_1423,In_113,N_848);
nor U1424 (N_1424,N_1063,N_1272);
nand U1425 (N_1425,In_112,N_1059);
and U1426 (N_1426,N_1102,N_999);
nor U1427 (N_1427,N_1111,N_888);
or U1428 (N_1428,N_270,N_749);
and U1429 (N_1429,N_1052,N_868);
or U1430 (N_1430,N_1304,N_814);
nor U1431 (N_1431,N_1,N_894);
nor U1432 (N_1432,In_925,N_1291);
or U1433 (N_1433,In_554,In_1126);
nand U1434 (N_1434,In_769,N_1285);
and U1435 (N_1435,N_1385,N_85);
and U1436 (N_1436,N_1312,N_1330);
nand U1437 (N_1437,N_318,N_1177);
nand U1438 (N_1438,N_1389,N_1325);
or U1439 (N_1439,N_996,N_1357);
nor U1440 (N_1440,N_1090,N_272);
and U1441 (N_1441,In_87,N_1083);
and U1442 (N_1442,N_1204,N_528);
nor U1443 (N_1443,N_1203,N_1273);
nor U1444 (N_1444,N_1349,N_1050);
nor U1445 (N_1445,N_944,In_897);
or U1446 (N_1446,N_915,N_800);
nand U1447 (N_1447,N_1348,N_1303);
nor U1448 (N_1448,N_680,In_986);
nand U1449 (N_1449,In_1022,N_4);
nand U1450 (N_1450,N_1247,N_675);
nor U1451 (N_1451,In_107,N_1230);
nand U1452 (N_1452,N_1319,In_515);
and U1453 (N_1453,N_712,N_1301);
or U1454 (N_1454,N_1254,N_0);
and U1455 (N_1455,N_1027,N_1114);
or U1456 (N_1456,In_411,N_1327);
nor U1457 (N_1457,N_1246,N_635);
nor U1458 (N_1458,N_1337,N_1297);
nor U1459 (N_1459,In_375,N_1149);
xor U1460 (N_1460,N_970,N_1241);
and U1461 (N_1461,N_1183,N_532);
or U1462 (N_1462,N_1066,N_1383);
nand U1463 (N_1463,N_655,N_446);
nand U1464 (N_1464,N_1021,N_951);
and U1465 (N_1465,N_1342,N_1171);
nor U1466 (N_1466,N_1051,N_1264);
or U1467 (N_1467,N_1192,N_945);
nand U1468 (N_1468,In_1264,N_630);
and U1469 (N_1469,N_708,N_742);
and U1470 (N_1470,N_382,N_1044);
nor U1471 (N_1471,N_1110,N_704);
nand U1472 (N_1472,In_1285,N_1328);
and U1473 (N_1473,N_776,In_1496);
or U1474 (N_1474,N_417,N_718);
nand U1475 (N_1475,In_373,N_1169);
nor U1476 (N_1476,In_966,In_1020);
and U1477 (N_1477,N_1333,N_1377);
and U1478 (N_1478,N_1229,N_1350);
and U1479 (N_1479,N_756,In_718);
or U1480 (N_1480,In_90,N_1165);
and U1481 (N_1481,N_1179,N_1098);
nand U1482 (N_1482,N_1373,N_662);
or U1483 (N_1483,N_1347,In_1278);
nor U1484 (N_1484,N_968,In_1190);
nor U1485 (N_1485,N_1355,N_1299);
nand U1486 (N_1486,N_1107,N_673);
nor U1487 (N_1487,N_1266,N_28);
nand U1488 (N_1488,In_708,N_961);
nand U1489 (N_1489,In_1152,In_281);
nor U1490 (N_1490,N_1323,In_12);
or U1491 (N_1491,N_1071,N_1223);
nor U1492 (N_1492,N_730,N_212);
nor U1493 (N_1493,In_1184,N_1390);
nand U1494 (N_1494,N_867,N_428);
xnor U1495 (N_1495,N_1391,N_1340);
nand U1496 (N_1496,N_1240,In_1612);
nor U1497 (N_1497,In_1440,N_623);
or U1498 (N_1498,N_1116,N_973);
and U1499 (N_1499,N_1331,N_1039);
or U1500 (N_1500,N_561,N_1231);
nor U1501 (N_1501,N_454,In_632);
or U1502 (N_1502,In_1404,N_1176);
or U1503 (N_1503,N_1281,N_1300);
nor U1504 (N_1504,N_1269,N_1101);
nand U1505 (N_1505,N_1164,N_1249);
and U1506 (N_1506,In_299,N_1398);
and U1507 (N_1507,N_303,N_1265);
nor U1508 (N_1508,N_455,N_882);
and U1509 (N_1509,N_1388,N_213);
nor U1510 (N_1510,N_810,N_1167);
nor U1511 (N_1511,N_1288,N_1396);
or U1512 (N_1512,N_1346,N_1018);
and U1513 (N_1513,N_1068,In_1173);
nor U1514 (N_1514,In_960,N_1095);
nor U1515 (N_1515,N_803,In_1751);
nand U1516 (N_1516,N_1280,N_1324);
or U1517 (N_1517,N_1219,N_1361);
nor U1518 (N_1518,N_821,N_1093);
and U1519 (N_1519,N_1222,In_311);
or U1520 (N_1520,In_1865,N_796);
or U1521 (N_1521,N_1215,N_1257);
or U1522 (N_1522,N_1042,N_1157);
nor U1523 (N_1523,N_1173,N_329);
and U1524 (N_1524,N_1317,N_1335);
nand U1525 (N_1525,N_579,N_1087);
nand U1526 (N_1526,N_667,N_1213);
or U1527 (N_1527,N_156,N_820);
nor U1528 (N_1528,N_1326,In_1957);
or U1529 (N_1529,In_1244,N_1080);
or U1530 (N_1530,N_1054,In_1829);
or U1531 (N_1531,N_1011,N_56);
and U1532 (N_1532,In_448,N_1239);
or U1533 (N_1533,N_1161,N_200);
nor U1534 (N_1534,N_1108,In_476);
nor U1535 (N_1535,N_1306,N_750);
nand U1536 (N_1536,N_627,N_1345);
and U1537 (N_1537,N_1338,In_1652);
nand U1538 (N_1538,N_1250,N_1226);
nand U1539 (N_1539,N_1261,N_1379);
or U1540 (N_1540,N_1210,N_869);
or U1541 (N_1541,N_235,N_1084);
or U1542 (N_1542,N_937,N_1278);
or U1543 (N_1543,N_650,N_1393);
or U1544 (N_1544,N_1295,N_215);
or U1545 (N_1545,In_243,N_1287);
nor U1546 (N_1546,N_1035,In_1964);
nand U1547 (N_1547,N_864,In_1782);
or U1548 (N_1548,N_638,In_477);
nor U1549 (N_1549,N_337,N_59);
and U1550 (N_1550,N_287,N_1308);
nand U1551 (N_1551,N_1294,N_1097);
and U1552 (N_1552,N_1351,N_1392);
nor U1553 (N_1553,N_1140,N_1216);
nor U1554 (N_1554,In_52,N_1380);
xor U1555 (N_1555,In_1469,N_1233);
xor U1556 (N_1556,N_1344,N_1292);
nor U1557 (N_1557,N_1134,In_330);
or U1558 (N_1558,In_1345,In_1819);
nor U1559 (N_1559,N_1260,In_508);
and U1560 (N_1560,In_1876,N_1321);
and U1561 (N_1561,N_1343,N_740);
or U1562 (N_1562,N_636,In_738);
or U1563 (N_1563,N_1218,N_1224);
nand U1564 (N_1564,N_1086,N_512);
and U1565 (N_1565,In_545,N_1236);
or U1566 (N_1566,N_1358,N_1117);
nor U1567 (N_1567,N_1201,N_1310);
or U1568 (N_1568,N_1386,In_181);
nor U1569 (N_1569,N_908,N_1045);
nand U1570 (N_1570,N_1352,N_345);
nor U1571 (N_1571,N_1243,N_237);
or U1572 (N_1572,N_593,N_834);
nor U1573 (N_1573,N_1235,N_1384);
and U1574 (N_1574,N_850,N_438);
nand U1575 (N_1575,In_1087,In_1766);
nand U1576 (N_1576,N_1154,N_1387);
or U1577 (N_1577,N_1234,In_120);
nand U1578 (N_1578,N_859,N_1399);
and U1579 (N_1579,N_1314,N_964);
nor U1580 (N_1580,In_653,In_1236);
and U1581 (N_1581,N_1360,N_548);
nand U1582 (N_1582,N_1004,In_1247);
and U1583 (N_1583,In_306,N_574);
or U1584 (N_1584,N_224,N_522);
nand U1585 (N_1585,In_1708,N_975);
nor U1586 (N_1586,N_1329,N_1142);
nor U1587 (N_1587,In_773,N_1227);
or U1588 (N_1588,In_524,In_1710);
nand U1589 (N_1589,N_1209,In_294);
nor U1590 (N_1590,N_142,In_1159);
or U1591 (N_1591,N_804,N_1184);
nor U1592 (N_1592,N_916,N_611);
nor U1593 (N_1593,N_1369,N_1309);
nand U1594 (N_1594,In_886,In_241);
and U1595 (N_1595,N_880,In_743);
or U1596 (N_1596,N_1013,N_724);
and U1597 (N_1597,N_936,N_1305);
xor U1598 (N_1598,N_860,N_1320);
and U1599 (N_1599,N_1382,In_58);
and U1600 (N_1600,N_1248,N_1481);
nor U1601 (N_1601,In_1376,N_1514);
nor U1602 (N_1602,N_1284,In_532);
or U1603 (N_1603,N_1408,N_1589);
or U1604 (N_1604,N_1237,N_1401);
and U1605 (N_1605,N_1364,N_1400);
xor U1606 (N_1606,N_1543,N_1277);
or U1607 (N_1607,N_1381,In_1061);
nand U1608 (N_1608,N_184,In_29);
and U1609 (N_1609,N_1522,N_1270);
and U1610 (N_1610,N_1459,N_1286);
nand U1611 (N_1611,N_1423,N_1221);
or U1612 (N_1612,In_1441,In_1421);
nor U1613 (N_1613,N_1554,N_1541);
nand U1614 (N_1614,N_1322,N_1567);
and U1615 (N_1615,N_1550,N_1531);
xnor U1616 (N_1616,N_1353,N_1493);
or U1617 (N_1617,N_1546,N_1556);
nor U1618 (N_1618,N_1512,N_388);
nor U1619 (N_1619,N_1332,N_1534);
nor U1620 (N_1620,In_1065,N_1473);
or U1621 (N_1621,N_726,N_602);
or U1622 (N_1622,N_780,N_1465);
or U1623 (N_1623,N_1507,N_1427);
and U1624 (N_1624,N_1587,In_1572);
and U1625 (N_1625,N_1200,In_1220);
nor U1626 (N_1626,N_1508,N_1477);
nand U1627 (N_1627,N_1523,N_1574);
nor U1628 (N_1628,N_1422,N_254);
nor U1629 (N_1629,N_1572,N_1037);
nand U1630 (N_1630,N_1132,N_1252);
nor U1631 (N_1631,N_1575,N_948);
nand U1632 (N_1632,N_1453,N_192);
nor U1633 (N_1633,N_861,N_1354);
nor U1634 (N_1634,N_1211,N_1205);
or U1635 (N_1635,N_414,N_1450);
nand U1636 (N_1636,N_1479,N_1559);
nand U1637 (N_1637,N_1582,N_1463);
nor U1638 (N_1638,In_1969,N_1245);
or U1639 (N_1639,N_1073,N_1394);
nor U1640 (N_1640,N_1315,N_1560);
or U1641 (N_1641,N_893,In_1997);
nand U1642 (N_1642,N_1429,In_1388);
nor U1643 (N_1643,N_1536,N_1088);
and U1644 (N_1644,N_1526,In_1575);
and U1645 (N_1645,N_1492,N_1500);
nand U1646 (N_1646,N_1505,N_910);
nand U1647 (N_1647,N_1494,N_1501);
nor U1648 (N_1648,N_1417,N_459);
and U1649 (N_1649,In_1111,N_1072);
nor U1650 (N_1650,N_1410,N_418);
nor U1651 (N_1651,N_1545,N_1585);
nor U1652 (N_1652,N_1448,N_1491);
or U1653 (N_1653,N_1225,N_1596);
and U1654 (N_1654,N_1532,N_831);
and U1655 (N_1655,In_884,N_1256);
nand U1656 (N_1656,N_1274,N_1503);
nand U1657 (N_1657,N_697,N_1268);
nand U1658 (N_1658,N_1404,N_828);
nand U1659 (N_1659,In_1443,N_1499);
nand U1660 (N_1660,N_1456,N_1262);
or U1661 (N_1661,N_954,N_1475);
nor U1662 (N_1662,N_1464,N_1533);
or U1663 (N_1663,N_1484,N_1403);
and U1664 (N_1664,N_1573,N_1518);
and U1665 (N_1665,N_1334,N_1524);
or U1666 (N_1666,N_1595,N_1553);
or U1667 (N_1667,N_463,N_1313);
or U1668 (N_1668,N_1395,N_1498);
or U1669 (N_1669,N_1443,N_1597);
and U1670 (N_1670,N_1438,N_1058);
and U1671 (N_1671,N_939,N_1425);
nor U1672 (N_1672,N_1077,N_1462);
or U1673 (N_1673,N_1480,N_1487);
and U1674 (N_1674,N_1571,N_1405);
or U1675 (N_1675,N_1511,N_1547);
nor U1676 (N_1676,N_1133,N_1106);
and U1677 (N_1677,N_640,N_986);
or U1678 (N_1678,N_441,N_1244);
or U1679 (N_1679,N_1586,N_1362);
nor U1680 (N_1680,In_318,In_698);
or U1681 (N_1681,N_1397,N_1506);
nand U1682 (N_1682,N_1544,N_745);
or U1683 (N_1683,N_1253,N_401);
nor U1684 (N_1684,N_1220,N_1413);
nor U1685 (N_1685,N_1460,N_1530);
and U1686 (N_1686,N_1598,N_926);
nand U1687 (N_1687,N_1485,N_1588);
and U1688 (N_1688,N_1549,N_896);
nor U1689 (N_1689,N_1441,N_1497);
and U1690 (N_1690,In_41,N_1591);
and U1691 (N_1691,N_1415,N_64);
or U1692 (N_1692,N_1446,N_491);
and U1693 (N_1693,N_1580,N_344);
and U1694 (N_1694,N_1451,N_1001);
nor U1695 (N_1695,N_1557,N_1555);
nor U1696 (N_1696,N_1442,N_1258);
nor U1697 (N_1697,N_1298,In_392);
and U1698 (N_1698,In_1998,N_966);
and U1699 (N_1699,N_1409,N_1406);
nand U1700 (N_1700,N_1055,N_1206);
nor U1701 (N_1701,N_1593,N_1435);
nand U1702 (N_1702,N_1449,N_1468);
or U1703 (N_1703,N_1193,N_651);
and U1704 (N_1704,N_1529,N_1452);
nand U1705 (N_1705,N_1316,N_1592);
nand U1706 (N_1706,N_1296,N_773);
and U1707 (N_1707,N_1489,N_1370);
or U1708 (N_1708,N_1568,N_1010);
and U1709 (N_1709,N_1081,N_1318);
and U1710 (N_1710,N_1029,N_1421);
or U1711 (N_1711,N_1466,N_1067);
or U1712 (N_1712,N_1414,N_1372);
nand U1713 (N_1713,N_1486,In_533);
and U1714 (N_1714,N_1420,N_1504);
nand U1715 (N_1715,N_1276,N_1434);
or U1716 (N_1716,N_1365,N_1540);
or U1717 (N_1717,N_1283,N_1495);
nor U1718 (N_1718,N_1282,N_1430);
and U1719 (N_1719,N_1551,N_1520);
and U1720 (N_1720,N_1474,In_929);
xnor U1721 (N_1721,N_824,N_1561);
nor U1722 (N_1722,N_1454,N_1168);
nor U1723 (N_1723,N_1552,N_1562);
nor U1724 (N_1724,N_1517,N_1579);
and U1725 (N_1725,N_168,N_1336);
nand U1726 (N_1726,N_1428,N_1476);
and U1727 (N_1727,N_1483,N_1583);
or U1728 (N_1728,N_1289,N_1432);
nand U1729 (N_1729,N_1402,N_1214);
nand U1730 (N_1730,N_1455,N_1032);
or U1731 (N_1731,N_1440,N_1584);
nand U1732 (N_1732,N_1570,In_466);
and U1733 (N_1733,N_1471,N_1407);
and U1734 (N_1734,N_1153,N_1488);
nor U1735 (N_1735,N_1502,N_1436);
nand U1736 (N_1736,In_46,N_1513);
and U1737 (N_1737,In_388,N_1444);
nand U1738 (N_1738,N_1564,N_1519);
nand U1739 (N_1739,N_1293,N_1558);
nand U1740 (N_1740,N_1469,N_1490);
or U1741 (N_1741,In_611,N_972);
nand U1742 (N_1742,In_1942,N_885);
or U1743 (N_1743,N_1510,N_1056);
nand U1744 (N_1744,N_1368,N_1367);
and U1745 (N_1745,N_890,N_1271);
nand U1746 (N_1746,N_1426,N_1302);
nand U1747 (N_1747,In_349,N_1217);
and U1748 (N_1748,N_1535,N_1418);
or U1749 (N_1749,N_1569,N_1251);
and U1750 (N_1750,N_1472,In_832);
nand U1751 (N_1751,N_1212,N_1065);
nand U1752 (N_1752,N_1238,N_1009);
or U1753 (N_1753,N_1539,N_1433);
and U1754 (N_1754,N_1113,N_1563);
nor U1755 (N_1755,N_1024,N_346);
nand U1756 (N_1756,N_1363,N_826);
nor U1757 (N_1757,N_1581,N_1375);
nand U1758 (N_1758,N_1028,N_1482);
nand U1759 (N_1759,N_938,N_1538);
nand U1760 (N_1760,N_1566,N_1089);
and U1761 (N_1761,N_1267,N_1275);
and U1762 (N_1762,N_369,N_830);
nor U1763 (N_1763,N_725,N_1232);
nand U1764 (N_1764,N_1594,In_1908);
nor U1765 (N_1765,In_680,In_20);
nor U1766 (N_1766,N_793,N_923);
nor U1767 (N_1767,N_862,N_1424);
xor U1768 (N_1768,N_1416,N_1470);
nand U1769 (N_1769,N_1255,N_1509);
or U1770 (N_1770,N_1457,N_1439);
nand U1771 (N_1771,N_1458,N_1467);
xor U1772 (N_1772,N_1590,N_1542);
and U1773 (N_1773,N_1521,N_1242);
or U1774 (N_1774,N_1049,N_1525);
or U1775 (N_1775,N_1419,N_1461);
nand U1776 (N_1776,N_1447,N_1478);
nor U1777 (N_1777,N_1528,N_1378);
nor U1778 (N_1778,In_6,N_180);
nor U1779 (N_1779,N_952,N_1412);
nor U1780 (N_1780,N_1431,N_1576);
nand U1781 (N_1781,N_1356,N_1015);
nand U1782 (N_1782,N_1527,In_259);
or U1783 (N_1783,N_1599,N_982);
nand U1784 (N_1784,N_325,N_472);
nor U1785 (N_1785,In_918,In_1937);
or U1786 (N_1786,In_909,N_835);
nand U1787 (N_1787,N_1516,N_1411);
or U1788 (N_1788,N_1537,N_276);
or U1789 (N_1789,N_920,N_1228);
or U1790 (N_1790,N_87,N_989);
nand U1791 (N_1791,N_1496,N_1105);
or U1792 (N_1792,N_1515,In_1888);
and U1793 (N_1793,In_1351,N_1445);
and U1794 (N_1794,N_1339,N_1565);
nand U1795 (N_1795,In_1826,N_1577);
nand U1796 (N_1796,N_1578,N_1437);
and U1797 (N_1797,In_415,In_1784);
nand U1798 (N_1798,N_1341,N_1259);
nand U1799 (N_1799,N_1371,N_1548);
or U1800 (N_1800,N_1635,N_1745);
and U1801 (N_1801,N_1659,N_1734);
and U1802 (N_1802,N_1653,N_1715);
nand U1803 (N_1803,N_1628,N_1743);
nand U1804 (N_1804,N_1638,N_1723);
and U1805 (N_1805,N_1704,N_1768);
and U1806 (N_1806,N_1748,N_1775);
or U1807 (N_1807,N_1660,N_1711);
xnor U1808 (N_1808,N_1735,N_1721);
nand U1809 (N_1809,N_1657,N_1649);
and U1810 (N_1810,N_1761,N_1603);
or U1811 (N_1811,N_1799,N_1644);
nand U1812 (N_1812,N_1687,N_1756);
and U1813 (N_1813,N_1605,N_1690);
and U1814 (N_1814,N_1640,N_1739);
nand U1815 (N_1815,N_1662,N_1624);
and U1816 (N_1816,N_1614,N_1698);
nor U1817 (N_1817,N_1759,N_1630);
xor U1818 (N_1818,N_1620,N_1700);
and U1819 (N_1819,N_1702,N_1648);
and U1820 (N_1820,N_1691,N_1779);
or U1821 (N_1821,N_1697,N_1694);
nor U1822 (N_1822,N_1728,N_1636);
nand U1823 (N_1823,N_1722,N_1616);
and U1824 (N_1824,N_1672,N_1727);
and U1825 (N_1825,N_1777,N_1701);
or U1826 (N_1826,N_1684,N_1661);
or U1827 (N_1827,N_1763,N_1750);
nand U1828 (N_1828,N_1726,N_1766);
nand U1829 (N_1829,N_1714,N_1601);
or U1830 (N_1830,N_1780,N_1781);
and U1831 (N_1831,N_1686,N_1643);
or U1832 (N_1832,N_1683,N_1622);
and U1833 (N_1833,N_1679,N_1736);
and U1834 (N_1834,N_1787,N_1771);
nor U1835 (N_1835,N_1755,N_1619);
nor U1836 (N_1836,N_1774,N_1623);
or U1837 (N_1837,N_1709,N_1767);
nor U1838 (N_1838,N_1789,N_1637);
or U1839 (N_1839,N_1778,N_1741);
and U1840 (N_1840,N_1627,N_1607);
and U1841 (N_1841,N_1754,N_1676);
nor U1842 (N_1842,N_1632,N_1742);
nand U1843 (N_1843,N_1669,N_1772);
or U1844 (N_1844,N_1706,N_1716);
and U1845 (N_1845,N_1703,N_1678);
or U1846 (N_1846,N_1747,N_1606);
or U1847 (N_1847,N_1666,N_1793);
and U1848 (N_1848,N_1729,N_1695);
or U1849 (N_1849,N_1765,N_1696);
xnor U1850 (N_1850,N_1655,N_1617);
nor U1851 (N_1851,N_1674,N_1668);
or U1852 (N_1852,N_1744,N_1783);
and U1853 (N_1853,N_1788,N_1786);
nand U1854 (N_1854,N_1733,N_1677);
or U1855 (N_1855,N_1718,N_1752);
or U1856 (N_1856,N_1708,N_1769);
or U1857 (N_1857,N_1719,N_1737);
or U1858 (N_1858,N_1689,N_1654);
xor U1859 (N_1859,N_1611,N_1773);
and U1860 (N_1860,N_1732,N_1724);
nor U1861 (N_1861,N_1784,N_1699);
nor U1862 (N_1862,N_1758,N_1791);
or U1863 (N_1863,N_1663,N_1629);
nand U1864 (N_1864,N_1664,N_1665);
nor U1865 (N_1865,N_1720,N_1705);
or U1866 (N_1866,N_1681,N_1612);
or U1867 (N_1867,N_1707,N_1785);
and U1868 (N_1868,N_1618,N_1796);
and U1869 (N_1869,N_1667,N_1680);
or U1870 (N_1870,N_1656,N_1639);
or U1871 (N_1871,N_1693,N_1731);
nor U1872 (N_1872,N_1749,N_1646);
nand U1873 (N_1873,N_1682,N_1675);
or U1874 (N_1874,N_1609,N_1751);
or U1875 (N_1875,N_1764,N_1692);
nor U1876 (N_1876,N_1625,N_1713);
nor U1877 (N_1877,N_1797,N_1645);
nand U1878 (N_1878,N_1738,N_1710);
and U1879 (N_1879,N_1730,N_1725);
and U1880 (N_1880,N_1685,N_1740);
nand U1881 (N_1881,N_1652,N_1610);
nor U1882 (N_1882,N_1642,N_1776);
nand U1883 (N_1883,N_1651,N_1600);
and U1884 (N_1884,N_1613,N_1608);
or U1885 (N_1885,N_1798,N_1650);
and U1886 (N_1886,N_1782,N_1658);
nand U1887 (N_1887,N_1621,N_1604);
or U1888 (N_1888,N_1753,N_1688);
xor U1889 (N_1889,N_1757,N_1615);
and U1890 (N_1890,N_1631,N_1647);
or U1891 (N_1891,N_1641,N_1673);
xnor U1892 (N_1892,N_1671,N_1634);
nor U1893 (N_1893,N_1717,N_1770);
nor U1894 (N_1894,N_1746,N_1712);
nor U1895 (N_1895,N_1670,N_1626);
nand U1896 (N_1896,N_1792,N_1602);
nor U1897 (N_1897,N_1790,N_1795);
and U1898 (N_1898,N_1633,N_1762);
nor U1899 (N_1899,N_1794,N_1760);
nor U1900 (N_1900,N_1631,N_1665);
nand U1901 (N_1901,N_1628,N_1786);
nor U1902 (N_1902,N_1644,N_1608);
or U1903 (N_1903,N_1722,N_1749);
nand U1904 (N_1904,N_1761,N_1757);
or U1905 (N_1905,N_1653,N_1639);
nor U1906 (N_1906,N_1658,N_1690);
or U1907 (N_1907,N_1616,N_1743);
and U1908 (N_1908,N_1733,N_1709);
and U1909 (N_1909,N_1623,N_1706);
or U1910 (N_1910,N_1736,N_1640);
nor U1911 (N_1911,N_1787,N_1670);
and U1912 (N_1912,N_1674,N_1758);
and U1913 (N_1913,N_1646,N_1727);
nor U1914 (N_1914,N_1768,N_1790);
and U1915 (N_1915,N_1675,N_1701);
nand U1916 (N_1916,N_1717,N_1701);
nand U1917 (N_1917,N_1764,N_1735);
nor U1918 (N_1918,N_1690,N_1675);
or U1919 (N_1919,N_1692,N_1790);
nor U1920 (N_1920,N_1633,N_1742);
or U1921 (N_1921,N_1785,N_1776);
nand U1922 (N_1922,N_1631,N_1781);
nor U1923 (N_1923,N_1681,N_1615);
or U1924 (N_1924,N_1722,N_1661);
nor U1925 (N_1925,N_1733,N_1690);
or U1926 (N_1926,N_1729,N_1652);
or U1927 (N_1927,N_1665,N_1749);
or U1928 (N_1928,N_1619,N_1624);
or U1929 (N_1929,N_1760,N_1627);
nor U1930 (N_1930,N_1769,N_1618);
xnor U1931 (N_1931,N_1621,N_1630);
xnor U1932 (N_1932,N_1714,N_1609);
nand U1933 (N_1933,N_1654,N_1630);
nor U1934 (N_1934,N_1657,N_1714);
nor U1935 (N_1935,N_1739,N_1784);
nand U1936 (N_1936,N_1740,N_1647);
or U1937 (N_1937,N_1697,N_1719);
xor U1938 (N_1938,N_1635,N_1750);
nor U1939 (N_1939,N_1682,N_1650);
nand U1940 (N_1940,N_1714,N_1665);
nand U1941 (N_1941,N_1670,N_1711);
or U1942 (N_1942,N_1647,N_1656);
or U1943 (N_1943,N_1651,N_1729);
or U1944 (N_1944,N_1769,N_1606);
nand U1945 (N_1945,N_1662,N_1766);
or U1946 (N_1946,N_1780,N_1721);
nand U1947 (N_1947,N_1790,N_1620);
and U1948 (N_1948,N_1718,N_1620);
and U1949 (N_1949,N_1683,N_1669);
nor U1950 (N_1950,N_1724,N_1722);
or U1951 (N_1951,N_1656,N_1644);
nand U1952 (N_1952,N_1731,N_1664);
nand U1953 (N_1953,N_1734,N_1685);
nor U1954 (N_1954,N_1772,N_1724);
nand U1955 (N_1955,N_1768,N_1655);
nor U1956 (N_1956,N_1726,N_1669);
nor U1957 (N_1957,N_1742,N_1603);
nor U1958 (N_1958,N_1624,N_1617);
or U1959 (N_1959,N_1695,N_1748);
nand U1960 (N_1960,N_1647,N_1628);
nor U1961 (N_1961,N_1663,N_1799);
nand U1962 (N_1962,N_1789,N_1771);
and U1963 (N_1963,N_1690,N_1603);
nor U1964 (N_1964,N_1748,N_1686);
nor U1965 (N_1965,N_1689,N_1655);
or U1966 (N_1966,N_1610,N_1792);
nor U1967 (N_1967,N_1742,N_1730);
nor U1968 (N_1968,N_1776,N_1695);
and U1969 (N_1969,N_1624,N_1749);
nand U1970 (N_1970,N_1651,N_1788);
or U1971 (N_1971,N_1714,N_1787);
nand U1972 (N_1972,N_1670,N_1715);
and U1973 (N_1973,N_1750,N_1748);
nand U1974 (N_1974,N_1793,N_1651);
and U1975 (N_1975,N_1735,N_1609);
and U1976 (N_1976,N_1658,N_1713);
or U1977 (N_1977,N_1641,N_1770);
nand U1978 (N_1978,N_1633,N_1606);
nand U1979 (N_1979,N_1729,N_1663);
or U1980 (N_1980,N_1664,N_1715);
nand U1981 (N_1981,N_1671,N_1610);
and U1982 (N_1982,N_1723,N_1790);
and U1983 (N_1983,N_1772,N_1711);
nand U1984 (N_1984,N_1702,N_1736);
nand U1985 (N_1985,N_1660,N_1794);
xnor U1986 (N_1986,N_1614,N_1680);
or U1987 (N_1987,N_1655,N_1681);
and U1988 (N_1988,N_1715,N_1613);
and U1989 (N_1989,N_1681,N_1696);
and U1990 (N_1990,N_1675,N_1637);
nor U1991 (N_1991,N_1621,N_1757);
and U1992 (N_1992,N_1726,N_1756);
or U1993 (N_1993,N_1798,N_1673);
or U1994 (N_1994,N_1735,N_1600);
and U1995 (N_1995,N_1685,N_1619);
nand U1996 (N_1996,N_1713,N_1659);
nand U1997 (N_1997,N_1663,N_1653);
nand U1998 (N_1998,N_1777,N_1688);
nor U1999 (N_1999,N_1728,N_1742);
nand U2000 (N_2000,N_1882,N_1975);
nor U2001 (N_2001,N_1847,N_1979);
nor U2002 (N_2002,N_1926,N_1938);
nor U2003 (N_2003,N_1849,N_1955);
or U2004 (N_2004,N_1890,N_1810);
or U2005 (N_2005,N_1997,N_1807);
or U2006 (N_2006,N_1915,N_1832);
nand U2007 (N_2007,N_1826,N_1827);
and U2008 (N_2008,N_1857,N_1881);
or U2009 (N_2009,N_1806,N_1896);
nor U2010 (N_2010,N_1893,N_1939);
nor U2011 (N_2011,N_1918,N_1987);
or U2012 (N_2012,N_1871,N_1921);
or U2013 (N_2013,N_1998,N_1838);
or U2014 (N_2014,N_1867,N_1984);
xnor U2015 (N_2015,N_1840,N_1949);
nand U2016 (N_2016,N_1801,N_1859);
and U2017 (N_2017,N_1863,N_1972);
nand U2018 (N_2018,N_1854,N_1988);
or U2019 (N_2019,N_1927,N_1917);
nor U2020 (N_2020,N_1866,N_1993);
or U2021 (N_2021,N_1895,N_1865);
and U2022 (N_2022,N_1925,N_1992);
nand U2023 (N_2023,N_1954,N_1873);
and U2024 (N_2024,N_1933,N_1951);
nand U2025 (N_2025,N_1960,N_1967);
nor U2026 (N_2026,N_1870,N_1958);
and U2027 (N_2027,N_1837,N_1875);
nand U2028 (N_2028,N_1853,N_1814);
or U2029 (N_2029,N_1982,N_1942);
nor U2030 (N_2030,N_1858,N_1953);
and U2031 (N_2031,N_1932,N_1985);
or U2032 (N_2032,N_1966,N_1907);
or U2033 (N_2033,N_1891,N_1940);
or U2034 (N_2034,N_1836,N_1821);
nand U2035 (N_2035,N_1959,N_1900);
or U2036 (N_2036,N_1922,N_1941);
nor U2037 (N_2037,N_1983,N_1828);
nand U2038 (N_2038,N_1924,N_1880);
and U2039 (N_2039,N_1971,N_1977);
nor U2040 (N_2040,N_1808,N_1990);
nor U2041 (N_2041,N_1878,N_1934);
nor U2042 (N_2042,N_1835,N_1876);
nor U2043 (N_2043,N_1989,N_1872);
nor U2044 (N_2044,N_1957,N_1906);
nand U2045 (N_2045,N_1823,N_1846);
and U2046 (N_2046,N_1839,N_1825);
or U2047 (N_2047,N_1874,N_1869);
or U2048 (N_2048,N_1976,N_1969);
and U2049 (N_2049,N_1819,N_1913);
or U2050 (N_2050,N_1848,N_1991);
nor U2051 (N_2051,N_1815,N_1868);
and U2052 (N_2052,N_1931,N_1803);
nor U2053 (N_2053,N_1965,N_1944);
and U2054 (N_2054,N_1812,N_1930);
or U2055 (N_2055,N_1898,N_1892);
nor U2056 (N_2056,N_1834,N_1860);
nand U2057 (N_2057,N_1820,N_1946);
nand U2058 (N_2058,N_1816,N_1943);
nand U2059 (N_2059,N_1910,N_1852);
and U2060 (N_2060,N_1888,N_1902);
nor U2061 (N_2061,N_1952,N_1899);
and U2062 (N_2062,N_1811,N_1877);
or U2063 (N_2063,N_1805,N_1978);
nor U2064 (N_2064,N_1862,N_1879);
nor U2065 (N_2065,N_1822,N_1802);
or U2066 (N_2066,N_1861,N_1928);
nor U2067 (N_2067,N_1809,N_1855);
and U2068 (N_2068,N_1980,N_1963);
nand U2069 (N_2069,N_1920,N_1929);
and U2070 (N_2070,N_1883,N_1968);
or U2071 (N_2071,N_1845,N_1914);
nor U2072 (N_2072,N_1850,N_1904);
nor U2073 (N_2073,N_1956,N_1818);
or U2074 (N_2074,N_1843,N_1894);
and U2075 (N_2075,N_1912,N_1889);
nor U2076 (N_2076,N_1973,N_1817);
nand U2077 (N_2077,N_1908,N_1885);
or U2078 (N_2078,N_1830,N_1996);
xnor U2079 (N_2079,N_1804,N_1947);
nand U2080 (N_2080,N_1897,N_1901);
nor U2081 (N_2081,N_1824,N_1903);
nand U2082 (N_2082,N_1962,N_1856);
nand U2083 (N_2083,N_1800,N_1935);
nor U2084 (N_2084,N_1916,N_1936);
and U2085 (N_2085,N_1999,N_1887);
and U2086 (N_2086,N_1864,N_1813);
or U2087 (N_2087,N_1945,N_1884);
nand U2088 (N_2088,N_1986,N_1974);
xor U2089 (N_2089,N_1948,N_1833);
and U2090 (N_2090,N_1842,N_1937);
nand U2091 (N_2091,N_1964,N_1923);
and U2092 (N_2092,N_1829,N_1995);
or U2093 (N_2093,N_1831,N_1919);
nor U2094 (N_2094,N_1950,N_1911);
and U2095 (N_2095,N_1961,N_1994);
and U2096 (N_2096,N_1905,N_1886);
nand U2097 (N_2097,N_1851,N_1981);
nand U2098 (N_2098,N_1844,N_1909);
and U2099 (N_2099,N_1841,N_1970);
nand U2100 (N_2100,N_1810,N_1930);
nand U2101 (N_2101,N_1987,N_1804);
or U2102 (N_2102,N_1845,N_1835);
and U2103 (N_2103,N_1803,N_1935);
or U2104 (N_2104,N_1928,N_1875);
or U2105 (N_2105,N_1945,N_1895);
nor U2106 (N_2106,N_1871,N_1966);
or U2107 (N_2107,N_1901,N_1909);
nor U2108 (N_2108,N_1844,N_1964);
nor U2109 (N_2109,N_1904,N_1974);
or U2110 (N_2110,N_1864,N_1817);
or U2111 (N_2111,N_1968,N_1889);
or U2112 (N_2112,N_1882,N_1823);
or U2113 (N_2113,N_1841,N_1925);
and U2114 (N_2114,N_1807,N_1821);
nor U2115 (N_2115,N_1881,N_1941);
or U2116 (N_2116,N_1911,N_1825);
or U2117 (N_2117,N_1976,N_1900);
and U2118 (N_2118,N_1838,N_1817);
or U2119 (N_2119,N_1844,N_1938);
nor U2120 (N_2120,N_1811,N_1986);
or U2121 (N_2121,N_1822,N_1984);
or U2122 (N_2122,N_1807,N_1857);
and U2123 (N_2123,N_1911,N_1851);
and U2124 (N_2124,N_1960,N_1898);
and U2125 (N_2125,N_1818,N_1929);
nor U2126 (N_2126,N_1820,N_1906);
and U2127 (N_2127,N_1982,N_1921);
or U2128 (N_2128,N_1936,N_1942);
nor U2129 (N_2129,N_1833,N_1956);
nor U2130 (N_2130,N_1848,N_1912);
nor U2131 (N_2131,N_1858,N_1816);
nand U2132 (N_2132,N_1895,N_1906);
and U2133 (N_2133,N_1910,N_1931);
or U2134 (N_2134,N_1943,N_1881);
nand U2135 (N_2135,N_1959,N_1800);
nor U2136 (N_2136,N_1937,N_1942);
nand U2137 (N_2137,N_1883,N_1938);
and U2138 (N_2138,N_1981,N_1838);
or U2139 (N_2139,N_1894,N_1801);
nor U2140 (N_2140,N_1862,N_1898);
nor U2141 (N_2141,N_1952,N_1855);
nand U2142 (N_2142,N_1814,N_1982);
or U2143 (N_2143,N_1885,N_1902);
nand U2144 (N_2144,N_1922,N_1809);
or U2145 (N_2145,N_1867,N_1827);
nor U2146 (N_2146,N_1826,N_1863);
or U2147 (N_2147,N_1890,N_1811);
or U2148 (N_2148,N_1945,N_1855);
or U2149 (N_2149,N_1810,N_1801);
and U2150 (N_2150,N_1825,N_1890);
or U2151 (N_2151,N_1957,N_1933);
and U2152 (N_2152,N_1836,N_1911);
nand U2153 (N_2153,N_1934,N_1808);
or U2154 (N_2154,N_1937,N_1910);
and U2155 (N_2155,N_1852,N_1915);
and U2156 (N_2156,N_1869,N_1988);
nand U2157 (N_2157,N_1899,N_1841);
and U2158 (N_2158,N_1943,N_1990);
and U2159 (N_2159,N_1955,N_1932);
or U2160 (N_2160,N_1939,N_1985);
and U2161 (N_2161,N_1977,N_1963);
nand U2162 (N_2162,N_1805,N_1945);
nand U2163 (N_2163,N_1973,N_1993);
and U2164 (N_2164,N_1930,N_1955);
nor U2165 (N_2165,N_1887,N_1923);
or U2166 (N_2166,N_1812,N_1829);
and U2167 (N_2167,N_1864,N_1808);
nor U2168 (N_2168,N_1962,N_1803);
or U2169 (N_2169,N_1906,N_1951);
nor U2170 (N_2170,N_1861,N_1963);
nor U2171 (N_2171,N_1831,N_1902);
and U2172 (N_2172,N_1991,N_1853);
and U2173 (N_2173,N_1903,N_1899);
nor U2174 (N_2174,N_1886,N_1834);
xor U2175 (N_2175,N_1816,N_1847);
nor U2176 (N_2176,N_1910,N_1851);
nor U2177 (N_2177,N_1802,N_1887);
or U2178 (N_2178,N_1961,N_1806);
xnor U2179 (N_2179,N_1991,N_1886);
xor U2180 (N_2180,N_1993,N_1970);
nor U2181 (N_2181,N_1829,N_1807);
nor U2182 (N_2182,N_1829,N_1928);
nand U2183 (N_2183,N_1957,N_1929);
nor U2184 (N_2184,N_1939,N_1987);
or U2185 (N_2185,N_1948,N_1842);
and U2186 (N_2186,N_1868,N_1819);
nand U2187 (N_2187,N_1962,N_1881);
nand U2188 (N_2188,N_1850,N_1901);
or U2189 (N_2189,N_1941,N_1927);
nor U2190 (N_2190,N_1850,N_1949);
or U2191 (N_2191,N_1881,N_1974);
xor U2192 (N_2192,N_1963,N_1966);
nand U2193 (N_2193,N_1966,N_1912);
nor U2194 (N_2194,N_1824,N_1840);
nand U2195 (N_2195,N_1906,N_1898);
nand U2196 (N_2196,N_1890,N_1973);
nand U2197 (N_2197,N_1869,N_1811);
nand U2198 (N_2198,N_1918,N_1906);
and U2199 (N_2199,N_1815,N_1986);
nor U2200 (N_2200,N_2199,N_2060);
nand U2201 (N_2201,N_2163,N_2072);
nand U2202 (N_2202,N_2136,N_2159);
and U2203 (N_2203,N_2024,N_2005);
xnor U2204 (N_2204,N_2158,N_2022);
nand U2205 (N_2205,N_2080,N_2032);
and U2206 (N_2206,N_2053,N_2054);
nand U2207 (N_2207,N_2188,N_2094);
nand U2208 (N_2208,N_2069,N_2198);
nand U2209 (N_2209,N_2183,N_2011);
nand U2210 (N_2210,N_2192,N_2034);
nand U2211 (N_2211,N_2065,N_2180);
and U2212 (N_2212,N_2195,N_2153);
nor U2213 (N_2213,N_2102,N_2055);
nor U2214 (N_2214,N_2074,N_2157);
and U2215 (N_2215,N_2026,N_2085);
nand U2216 (N_2216,N_2062,N_2048);
or U2217 (N_2217,N_2049,N_2106);
or U2218 (N_2218,N_2045,N_2135);
nand U2219 (N_2219,N_2037,N_2079);
and U2220 (N_2220,N_2082,N_2149);
nand U2221 (N_2221,N_2160,N_2029);
nand U2222 (N_2222,N_2178,N_2111);
or U2223 (N_2223,N_2044,N_2150);
nand U2224 (N_2224,N_2012,N_2186);
nand U2225 (N_2225,N_2015,N_2047);
and U2226 (N_2226,N_2127,N_2025);
nand U2227 (N_2227,N_2021,N_2088);
nand U2228 (N_2228,N_2017,N_2092);
and U2229 (N_2229,N_2139,N_2116);
nor U2230 (N_2230,N_2058,N_2133);
and U2231 (N_2231,N_2078,N_2121);
nand U2232 (N_2232,N_2152,N_2075);
nor U2233 (N_2233,N_2052,N_2042);
nand U2234 (N_2234,N_2130,N_2023);
nand U2235 (N_2235,N_2169,N_2128);
or U2236 (N_2236,N_2089,N_2193);
nor U2237 (N_2237,N_2181,N_2061);
or U2238 (N_2238,N_2165,N_2156);
nand U2239 (N_2239,N_2081,N_2145);
nor U2240 (N_2240,N_2166,N_2105);
nor U2241 (N_2241,N_2134,N_2090);
nor U2242 (N_2242,N_2035,N_2114);
nor U2243 (N_2243,N_2144,N_2103);
nand U2244 (N_2244,N_2190,N_2132);
or U2245 (N_2245,N_2197,N_2126);
nor U2246 (N_2246,N_2138,N_2093);
and U2247 (N_2247,N_2194,N_2039);
nor U2248 (N_2248,N_2027,N_2036);
nor U2249 (N_2249,N_2184,N_2112);
and U2250 (N_2250,N_2108,N_2170);
nor U2251 (N_2251,N_2063,N_2119);
nand U2252 (N_2252,N_2162,N_2175);
nor U2253 (N_2253,N_2123,N_2019);
and U2254 (N_2254,N_2187,N_2142);
nand U2255 (N_2255,N_2057,N_2056);
nor U2256 (N_2256,N_2018,N_2028);
nor U2257 (N_2257,N_2031,N_2115);
and U2258 (N_2258,N_2050,N_2168);
or U2259 (N_2259,N_2174,N_2071);
and U2260 (N_2260,N_2064,N_2004);
and U2261 (N_2261,N_2095,N_2107);
nand U2262 (N_2262,N_2001,N_2124);
and U2263 (N_2263,N_2125,N_2077);
or U2264 (N_2264,N_2148,N_2087);
nand U2265 (N_2265,N_2185,N_2068);
and U2266 (N_2266,N_2118,N_2020);
nand U2267 (N_2267,N_2154,N_2038);
and U2268 (N_2268,N_2141,N_2122);
nor U2269 (N_2269,N_2009,N_2140);
nand U2270 (N_2270,N_2086,N_2117);
nor U2271 (N_2271,N_2059,N_2173);
nor U2272 (N_2272,N_2066,N_2014);
or U2273 (N_2273,N_2167,N_2146);
nor U2274 (N_2274,N_2137,N_2003);
nand U2275 (N_2275,N_2182,N_2164);
nand U2276 (N_2276,N_2171,N_2076);
and U2277 (N_2277,N_2110,N_2101);
nor U2278 (N_2278,N_2070,N_2161);
nor U2279 (N_2279,N_2006,N_2030);
nand U2280 (N_2280,N_2043,N_2051);
nand U2281 (N_2281,N_2013,N_2000);
nor U2282 (N_2282,N_2196,N_2091);
nand U2283 (N_2283,N_2155,N_2084);
nand U2284 (N_2284,N_2151,N_2041);
and U2285 (N_2285,N_2096,N_2104);
nand U2286 (N_2286,N_2007,N_2120);
and U2287 (N_2287,N_2098,N_2172);
nand U2288 (N_2288,N_2002,N_2177);
and U2289 (N_2289,N_2131,N_2100);
and U2290 (N_2290,N_2143,N_2176);
nor U2291 (N_2291,N_2033,N_2010);
or U2292 (N_2292,N_2016,N_2040);
nand U2293 (N_2293,N_2067,N_2008);
nor U2294 (N_2294,N_2189,N_2191);
or U2295 (N_2295,N_2046,N_2073);
nor U2296 (N_2296,N_2179,N_2099);
nor U2297 (N_2297,N_2147,N_2129);
and U2298 (N_2298,N_2083,N_2113);
nor U2299 (N_2299,N_2109,N_2097);
nor U2300 (N_2300,N_2145,N_2065);
and U2301 (N_2301,N_2133,N_2096);
or U2302 (N_2302,N_2167,N_2022);
or U2303 (N_2303,N_2014,N_2104);
xor U2304 (N_2304,N_2045,N_2018);
and U2305 (N_2305,N_2126,N_2196);
xnor U2306 (N_2306,N_2142,N_2034);
nand U2307 (N_2307,N_2085,N_2083);
nor U2308 (N_2308,N_2007,N_2147);
nand U2309 (N_2309,N_2022,N_2007);
nand U2310 (N_2310,N_2069,N_2063);
nor U2311 (N_2311,N_2101,N_2054);
nand U2312 (N_2312,N_2084,N_2198);
or U2313 (N_2313,N_2163,N_2082);
nand U2314 (N_2314,N_2121,N_2054);
nor U2315 (N_2315,N_2053,N_2134);
nor U2316 (N_2316,N_2057,N_2121);
or U2317 (N_2317,N_2195,N_2078);
or U2318 (N_2318,N_2186,N_2110);
and U2319 (N_2319,N_2139,N_2068);
nor U2320 (N_2320,N_2111,N_2142);
nand U2321 (N_2321,N_2184,N_2120);
and U2322 (N_2322,N_2077,N_2176);
or U2323 (N_2323,N_2041,N_2099);
or U2324 (N_2324,N_2172,N_2046);
or U2325 (N_2325,N_2138,N_2084);
or U2326 (N_2326,N_2196,N_2142);
nand U2327 (N_2327,N_2066,N_2016);
xnor U2328 (N_2328,N_2188,N_2023);
nor U2329 (N_2329,N_2184,N_2031);
nand U2330 (N_2330,N_2001,N_2093);
nand U2331 (N_2331,N_2047,N_2040);
nand U2332 (N_2332,N_2142,N_2082);
or U2333 (N_2333,N_2097,N_2044);
nand U2334 (N_2334,N_2041,N_2001);
nand U2335 (N_2335,N_2188,N_2036);
or U2336 (N_2336,N_2153,N_2071);
or U2337 (N_2337,N_2060,N_2165);
or U2338 (N_2338,N_2143,N_2167);
or U2339 (N_2339,N_2174,N_2196);
and U2340 (N_2340,N_2170,N_2191);
or U2341 (N_2341,N_2156,N_2010);
and U2342 (N_2342,N_2123,N_2000);
nand U2343 (N_2343,N_2199,N_2042);
nor U2344 (N_2344,N_2016,N_2108);
nand U2345 (N_2345,N_2065,N_2199);
nor U2346 (N_2346,N_2085,N_2168);
and U2347 (N_2347,N_2037,N_2055);
nand U2348 (N_2348,N_2030,N_2183);
nand U2349 (N_2349,N_2033,N_2022);
and U2350 (N_2350,N_2126,N_2089);
or U2351 (N_2351,N_2043,N_2085);
nor U2352 (N_2352,N_2087,N_2128);
nor U2353 (N_2353,N_2042,N_2102);
or U2354 (N_2354,N_2041,N_2087);
or U2355 (N_2355,N_2012,N_2060);
nor U2356 (N_2356,N_2176,N_2026);
or U2357 (N_2357,N_2151,N_2022);
nor U2358 (N_2358,N_2161,N_2191);
and U2359 (N_2359,N_2181,N_2175);
nand U2360 (N_2360,N_2198,N_2152);
and U2361 (N_2361,N_2140,N_2095);
nor U2362 (N_2362,N_2057,N_2154);
or U2363 (N_2363,N_2008,N_2178);
nor U2364 (N_2364,N_2044,N_2017);
or U2365 (N_2365,N_2116,N_2035);
or U2366 (N_2366,N_2176,N_2066);
and U2367 (N_2367,N_2095,N_2153);
nand U2368 (N_2368,N_2180,N_2071);
nand U2369 (N_2369,N_2160,N_2118);
nand U2370 (N_2370,N_2137,N_2162);
nand U2371 (N_2371,N_2022,N_2078);
nand U2372 (N_2372,N_2026,N_2133);
nor U2373 (N_2373,N_2007,N_2046);
or U2374 (N_2374,N_2036,N_2010);
nor U2375 (N_2375,N_2040,N_2173);
or U2376 (N_2376,N_2189,N_2047);
and U2377 (N_2377,N_2120,N_2121);
and U2378 (N_2378,N_2181,N_2054);
or U2379 (N_2379,N_2026,N_2009);
and U2380 (N_2380,N_2154,N_2104);
or U2381 (N_2381,N_2079,N_2026);
nand U2382 (N_2382,N_2037,N_2028);
nand U2383 (N_2383,N_2001,N_2155);
nor U2384 (N_2384,N_2077,N_2022);
xnor U2385 (N_2385,N_2155,N_2120);
nor U2386 (N_2386,N_2030,N_2197);
or U2387 (N_2387,N_2063,N_2144);
nor U2388 (N_2388,N_2142,N_2011);
nand U2389 (N_2389,N_2075,N_2039);
or U2390 (N_2390,N_2014,N_2174);
or U2391 (N_2391,N_2171,N_2186);
or U2392 (N_2392,N_2011,N_2110);
and U2393 (N_2393,N_2026,N_2104);
nand U2394 (N_2394,N_2102,N_2047);
or U2395 (N_2395,N_2051,N_2003);
nor U2396 (N_2396,N_2182,N_2151);
nand U2397 (N_2397,N_2149,N_2098);
nand U2398 (N_2398,N_2116,N_2046);
or U2399 (N_2399,N_2048,N_2009);
or U2400 (N_2400,N_2305,N_2337);
nor U2401 (N_2401,N_2319,N_2317);
or U2402 (N_2402,N_2277,N_2336);
nor U2403 (N_2403,N_2331,N_2200);
nor U2404 (N_2404,N_2262,N_2368);
nand U2405 (N_2405,N_2315,N_2310);
nand U2406 (N_2406,N_2351,N_2341);
or U2407 (N_2407,N_2306,N_2399);
nor U2408 (N_2408,N_2316,N_2230);
or U2409 (N_2409,N_2298,N_2360);
and U2410 (N_2410,N_2258,N_2376);
xnor U2411 (N_2411,N_2286,N_2361);
nor U2412 (N_2412,N_2215,N_2297);
nor U2413 (N_2413,N_2304,N_2350);
nor U2414 (N_2414,N_2344,N_2364);
nand U2415 (N_2415,N_2342,N_2359);
or U2416 (N_2416,N_2222,N_2375);
or U2417 (N_2417,N_2389,N_2216);
and U2418 (N_2418,N_2202,N_2290);
and U2419 (N_2419,N_2362,N_2203);
or U2420 (N_2420,N_2240,N_2274);
nand U2421 (N_2421,N_2377,N_2296);
nor U2422 (N_2422,N_2205,N_2241);
and U2423 (N_2423,N_2394,N_2221);
or U2424 (N_2424,N_2340,N_2246);
or U2425 (N_2425,N_2392,N_2352);
xnor U2426 (N_2426,N_2268,N_2300);
nor U2427 (N_2427,N_2391,N_2302);
nor U2428 (N_2428,N_2227,N_2294);
nand U2429 (N_2429,N_2272,N_2333);
and U2430 (N_2430,N_2270,N_2214);
nand U2431 (N_2431,N_2243,N_2311);
nand U2432 (N_2432,N_2365,N_2385);
nand U2433 (N_2433,N_2387,N_2212);
and U2434 (N_2434,N_2244,N_2398);
or U2435 (N_2435,N_2312,N_2349);
or U2436 (N_2436,N_2373,N_2252);
nand U2437 (N_2437,N_2223,N_2318);
nor U2438 (N_2438,N_2374,N_2208);
or U2439 (N_2439,N_2369,N_2356);
nand U2440 (N_2440,N_2322,N_2224);
and U2441 (N_2441,N_2313,N_2325);
nor U2442 (N_2442,N_2234,N_2260);
nor U2443 (N_2443,N_2220,N_2379);
nand U2444 (N_2444,N_2232,N_2326);
nand U2445 (N_2445,N_2372,N_2239);
and U2446 (N_2446,N_2238,N_2235);
and U2447 (N_2447,N_2237,N_2284);
and U2448 (N_2448,N_2261,N_2275);
nand U2449 (N_2449,N_2291,N_2345);
or U2450 (N_2450,N_2335,N_2267);
and U2451 (N_2451,N_2281,N_2251);
or U2452 (N_2452,N_2210,N_2242);
nor U2453 (N_2453,N_2219,N_2382);
or U2454 (N_2454,N_2226,N_2236);
nand U2455 (N_2455,N_2330,N_2283);
nand U2456 (N_2456,N_2321,N_2254);
nor U2457 (N_2457,N_2393,N_2282);
nand U2458 (N_2458,N_2299,N_2347);
and U2459 (N_2459,N_2327,N_2295);
and U2460 (N_2460,N_2328,N_2265);
nand U2461 (N_2461,N_2338,N_2201);
and U2462 (N_2462,N_2320,N_2249);
nor U2463 (N_2463,N_2370,N_2264);
and U2464 (N_2464,N_2363,N_2228);
nand U2465 (N_2465,N_2279,N_2371);
and U2466 (N_2466,N_2266,N_2273);
or U2467 (N_2467,N_2358,N_2384);
or U2468 (N_2468,N_2278,N_2396);
nor U2469 (N_2469,N_2378,N_2324);
and U2470 (N_2470,N_2292,N_2388);
and U2471 (N_2471,N_2257,N_2245);
or U2472 (N_2472,N_2381,N_2248);
and U2473 (N_2473,N_2269,N_2263);
nor U2474 (N_2474,N_2307,N_2211);
nand U2475 (N_2475,N_2367,N_2288);
nor U2476 (N_2476,N_2386,N_2383);
or U2477 (N_2477,N_2231,N_2354);
or U2478 (N_2478,N_2247,N_2259);
nand U2479 (N_2479,N_2218,N_2229);
and U2480 (N_2480,N_2253,N_2323);
and U2481 (N_2481,N_2287,N_2213);
nor U2482 (N_2482,N_2353,N_2314);
nand U2483 (N_2483,N_2357,N_2346);
nand U2484 (N_2484,N_2343,N_2303);
nor U2485 (N_2485,N_2329,N_2285);
nor U2486 (N_2486,N_2348,N_2250);
nor U2487 (N_2487,N_2233,N_2390);
nor U2488 (N_2488,N_2217,N_2293);
nand U2489 (N_2489,N_2276,N_2225);
and U2490 (N_2490,N_2256,N_2309);
and U2491 (N_2491,N_2339,N_2301);
nand U2492 (N_2492,N_2206,N_2255);
or U2493 (N_2493,N_2380,N_2355);
or U2494 (N_2494,N_2397,N_2332);
nor U2495 (N_2495,N_2204,N_2207);
nand U2496 (N_2496,N_2289,N_2271);
nor U2497 (N_2497,N_2366,N_2334);
and U2498 (N_2498,N_2209,N_2395);
and U2499 (N_2499,N_2308,N_2280);
nand U2500 (N_2500,N_2392,N_2361);
nand U2501 (N_2501,N_2338,N_2379);
nor U2502 (N_2502,N_2243,N_2252);
nand U2503 (N_2503,N_2355,N_2288);
nor U2504 (N_2504,N_2253,N_2299);
or U2505 (N_2505,N_2285,N_2244);
nand U2506 (N_2506,N_2222,N_2336);
or U2507 (N_2507,N_2354,N_2322);
and U2508 (N_2508,N_2378,N_2289);
or U2509 (N_2509,N_2284,N_2295);
nor U2510 (N_2510,N_2282,N_2274);
and U2511 (N_2511,N_2355,N_2251);
nand U2512 (N_2512,N_2377,N_2317);
nor U2513 (N_2513,N_2250,N_2247);
nor U2514 (N_2514,N_2358,N_2327);
nand U2515 (N_2515,N_2300,N_2390);
or U2516 (N_2516,N_2234,N_2324);
or U2517 (N_2517,N_2269,N_2343);
nand U2518 (N_2518,N_2360,N_2341);
nand U2519 (N_2519,N_2219,N_2247);
xor U2520 (N_2520,N_2270,N_2375);
and U2521 (N_2521,N_2222,N_2329);
nor U2522 (N_2522,N_2328,N_2212);
nor U2523 (N_2523,N_2235,N_2386);
or U2524 (N_2524,N_2305,N_2308);
nand U2525 (N_2525,N_2235,N_2347);
or U2526 (N_2526,N_2304,N_2376);
nand U2527 (N_2527,N_2257,N_2201);
nand U2528 (N_2528,N_2222,N_2256);
and U2529 (N_2529,N_2393,N_2332);
nand U2530 (N_2530,N_2239,N_2396);
nand U2531 (N_2531,N_2363,N_2203);
nor U2532 (N_2532,N_2259,N_2276);
and U2533 (N_2533,N_2261,N_2297);
or U2534 (N_2534,N_2223,N_2283);
nor U2535 (N_2535,N_2240,N_2367);
nor U2536 (N_2536,N_2328,N_2288);
and U2537 (N_2537,N_2390,N_2382);
or U2538 (N_2538,N_2270,N_2396);
nand U2539 (N_2539,N_2363,N_2327);
xnor U2540 (N_2540,N_2315,N_2278);
and U2541 (N_2541,N_2283,N_2275);
nor U2542 (N_2542,N_2391,N_2342);
or U2543 (N_2543,N_2392,N_2326);
nor U2544 (N_2544,N_2296,N_2290);
nor U2545 (N_2545,N_2360,N_2326);
nand U2546 (N_2546,N_2351,N_2309);
and U2547 (N_2547,N_2200,N_2395);
nor U2548 (N_2548,N_2211,N_2246);
and U2549 (N_2549,N_2210,N_2267);
nor U2550 (N_2550,N_2201,N_2296);
nor U2551 (N_2551,N_2372,N_2312);
xor U2552 (N_2552,N_2279,N_2212);
nand U2553 (N_2553,N_2213,N_2298);
and U2554 (N_2554,N_2273,N_2364);
or U2555 (N_2555,N_2238,N_2386);
or U2556 (N_2556,N_2359,N_2387);
nor U2557 (N_2557,N_2397,N_2304);
or U2558 (N_2558,N_2342,N_2393);
nor U2559 (N_2559,N_2331,N_2392);
or U2560 (N_2560,N_2349,N_2286);
nand U2561 (N_2561,N_2243,N_2315);
and U2562 (N_2562,N_2345,N_2325);
nor U2563 (N_2563,N_2364,N_2337);
nor U2564 (N_2564,N_2223,N_2344);
nand U2565 (N_2565,N_2380,N_2370);
nand U2566 (N_2566,N_2279,N_2347);
nand U2567 (N_2567,N_2290,N_2344);
nor U2568 (N_2568,N_2205,N_2357);
xnor U2569 (N_2569,N_2342,N_2246);
nand U2570 (N_2570,N_2361,N_2337);
and U2571 (N_2571,N_2371,N_2359);
nand U2572 (N_2572,N_2394,N_2387);
or U2573 (N_2573,N_2314,N_2347);
nand U2574 (N_2574,N_2242,N_2323);
and U2575 (N_2575,N_2396,N_2279);
nor U2576 (N_2576,N_2250,N_2288);
and U2577 (N_2577,N_2303,N_2220);
or U2578 (N_2578,N_2328,N_2248);
nand U2579 (N_2579,N_2237,N_2359);
or U2580 (N_2580,N_2368,N_2350);
or U2581 (N_2581,N_2384,N_2308);
nor U2582 (N_2582,N_2246,N_2321);
and U2583 (N_2583,N_2383,N_2322);
nor U2584 (N_2584,N_2292,N_2302);
nor U2585 (N_2585,N_2240,N_2326);
nand U2586 (N_2586,N_2398,N_2203);
nor U2587 (N_2587,N_2250,N_2361);
nand U2588 (N_2588,N_2258,N_2235);
nor U2589 (N_2589,N_2308,N_2387);
nor U2590 (N_2590,N_2386,N_2358);
or U2591 (N_2591,N_2377,N_2210);
nor U2592 (N_2592,N_2372,N_2342);
nand U2593 (N_2593,N_2253,N_2392);
nor U2594 (N_2594,N_2208,N_2254);
and U2595 (N_2595,N_2354,N_2289);
nor U2596 (N_2596,N_2279,N_2357);
nand U2597 (N_2597,N_2208,N_2248);
nand U2598 (N_2598,N_2237,N_2233);
xor U2599 (N_2599,N_2295,N_2299);
or U2600 (N_2600,N_2483,N_2430);
and U2601 (N_2601,N_2431,N_2413);
or U2602 (N_2602,N_2502,N_2590);
nor U2603 (N_2603,N_2462,N_2515);
or U2604 (N_2604,N_2579,N_2514);
or U2605 (N_2605,N_2432,N_2442);
nor U2606 (N_2606,N_2500,N_2538);
nor U2607 (N_2607,N_2438,N_2476);
nor U2608 (N_2608,N_2424,N_2480);
or U2609 (N_2609,N_2486,N_2535);
nand U2610 (N_2610,N_2477,N_2578);
nand U2611 (N_2611,N_2420,N_2503);
nand U2612 (N_2612,N_2419,N_2411);
nor U2613 (N_2613,N_2465,N_2415);
and U2614 (N_2614,N_2456,N_2519);
or U2615 (N_2615,N_2494,N_2447);
or U2616 (N_2616,N_2570,N_2541);
nor U2617 (N_2617,N_2402,N_2501);
or U2618 (N_2618,N_2464,N_2416);
and U2619 (N_2619,N_2518,N_2542);
nand U2620 (N_2620,N_2497,N_2532);
and U2621 (N_2621,N_2587,N_2567);
or U2622 (N_2622,N_2548,N_2547);
and U2623 (N_2623,N_2435,N_2482);
and U2624 (N_2624,N_2555,N_2577);
nor U2625 (N_2625,N_2516,N_2466);
xnor U2626 (N_2626,N_2427,N_2487);
nand U2627 (N_2627,N_2546,N_2429);
nand U2628 (N_2628,N_2543,N_2454);
or U2629 (N_2629,N_2531,N_2523);
nor U2630 (N_2630,N_2568,N_2493);
and U2631 (N_2631,N_2457,N_2461);
or U2632 (N_2632,N_2463,N_2560);
and U2633 (N_2633,N_2444,N_2533);
nor U2634 (N_2634,N_2561,N_2537);
and U2635 (N_2635,N_2481,N_2403);
and U2636 (N_2636,N_2484,N_2529);
and U2637 (N_2637,N_2410,N_2414);
and U2638 (N_2638,N_2574,N_2401);
and U2639 (N_2639,N_2556,N_2450);
and U2640 (N_2640,N_2443,N_2545);
nand U2641 (N_2641,N_2460,N_2544);
or U2642 (N_2642,N_2441,N_2525);
nand U2643 (N_2643,N_2508,N_2451);
xor U2644 (N_2644,N_2510,N_2598);
xnor U2645 (N_2645,N_2407,N_2549);
or U2646 (N_2646,N_2520,N_2552);
nand U2647 (N_2647,N_2522,N_2526);
and U2648 (N_2648,N_2473,N_2434);
nor U2649 (N_2649,N_2505,N_2536);
or U2650 (N_2650,N_2474,N_2563);
or U2651 (N_2651,N_2507,N_2490);
and U2652 (N_2652,N_2448,N_2585);
and U2653 (N_2653,N_2580,N_2485);
and U2654 (N_2654,N_2566,N_2557);
nand U2655 (N_2655,N_2495,N_2470);
nand U2656 (N_2656,N_2425,N_2540);
nand U2657 (N_2657,N_2423,N_2586);
or U2658 (N_2658,N_2599,N_2571);
nand U2659 (N_2659,N_2573,N_2565);
or U2660 (N_2660,N_2412,N_2436);
xnor U2661 (N_2661,N_2446,N_2440);
or U2662 (N_2662,N_2452,N_2478);
and U2663 (N_2663,N_2453,N_2489);
or U2664 (N_2664,N_2504,N_2589);
nor U2665 (N_2665,N_2575,N_2592);
nor U2666 (N_2666,N_2553,N_2421);
nor U2667 (N_2667,N_2499,N_2400);
and U2668 (N_2668,N_2539,N_2512);
nand U2669 (N_2669,N_2554,N_2596);
or U2670 (N_2670,N_2594,N_2597);
and U2671 (N_2671,N_2409,N_2591);
or U2672 (N_2672,N_2458,N_2509);
nor U2673 (N_2673,N_2528,N_2517);
nand U2674 (N_2674,N_2471,N_2595);
nand U2675 (N_2675,N_2550,N_2588);
or U2676 (N_2676,N_2521,N_2433);
or U2677 (N_2677,N_2469,N_2459);
and U2678 (N_2678,N_2455,N_2404);
and U2679 (N_2679,N_2475,N_2417);
or U2680 (N_2680,N_2408,N_2422);
nand U2681 (N_2681,N_2488,N_2582);
nand U2682 (N_2682,N_2437,N_2426);
nand U2683 (N_2683,N_2472,N_2564);
and U2684 (N_2684,N_2491,N_2559);
and U2685 (N_2685,N_2449,N_2558);
or U2686 (N_2686,N_2530,N_2551);
nor U2687 (N_2687,N_2584,N_2405);
nand U2688 (N_2688,N_2468,N_2498);
and U2689 (N_2689,N_2439,N_2524);
and U2690 (N_2690,N_2479,N_2496);
and U2691 (N_2691,N_2418,N_2511);
nor U2692 (N_2692,N_2581,N_2428);
nand U2693 (N_2693,N_2467,N_2593);
or U2694 (N_2694,N_2492,N_2576);
or U2695 (N_2695,N_2527,N_2534);
and U2696 (N_2696,N_2406,N_2569);
or U2697 (N_2697,N_2572,N_2583);
or U2698 (N_2698,N_2513,N_2445);
nor U2699 (N_2699,N_2506,N_2562);
and U2700 (N_2700,N_2576,N_2578);
and U2701 (N_2701,N_2544,N_2503);
and U2702 (N_2702,N_2523,N_2591);
or U2703 (N_2703,N_2478,N_2425);
or U2704 (N_2704,N_2561,N_2404);
xnor U2705 (N_2705,N_2400,N_2507);
and U2706 (N_2706,N_2499,N_2574);
nand U2707 (N_2707,N_2486,N_2546);
nand U2708 (N_2708,N_2536,N_2426);
nand U2709 (N_2709,N_2430,N_2570);
nand U2710 (N_2710,N_2518,N_2447);
nor U2711 (N_2711,N_2473,N_2585);
or U2712 (N_2712,N_2562,N_2445);
xor U2713 (N_2713,N_2439,N_2472);
nand U2714 (N_2714,N_2575,N_2492);
nand U2715 (N_2715,N_2532,N_2505);
xnor U2716 (N_2716,N_2476,N_2514);
and U2717 (N_2717,N_2407,N_2498);
nor U2718 (N_2718,N_2538,N_2468);
nand U2719 (N_2719,N_2497,N_2558);
and U2720 (N_2720,N_2575,N_2453);
and U2721 (N_2721,N_2426,N_2419);
nand U2722 (N_2722,N_2549,N_2437);
nand U2723 (N_2723,N_2458,N_2426);
or U2724 (N_2724,N_2455,N_2468);
or U2725 (N_2725,N_2578,N_2552);
and U2726 (N_2726,N_2525,N_2453);
nor U2727 (N_2727,N_2411,N_2455);
and U2728 (N_2728,N_2448,N_2509);
nand U2729 (N_2729,N_2536,N_2496);
and U2730 (N_2730,N_2457,N_2467);
xnor U2731 (N_2731,N_2470,N_2421);
and U2732 (N_2732,N_2511,N_2431);
and U2733 (N_2733,N_2467,N_2506);
or U2734 (N_2734,N_2422,N_2420);
nand U2735 (N_2735,N_2522,N_2542);
xnor U2736 (N_2736,N_2400,N_2535);
or U2737 (N_2737,N_2435,N_2551);
nor U2738 (N_2738,N_2450,N_2564);
or U2739 (N_2739,N_2522,N_2553);
nand U2740 (N_2740,N_2533,N_2506);
and U2741 (N_2741,N_2457,N_2515);
and U2742 (N_2742,N_2415,N_2426);
or U2743 (N_2743,N_2410,N_2571);
or U2744 (N_2744,N_2473,N_2547);
and U2745 (N_2745,N_2564,N_2503);
and U2746 (N_2746,N_2500,N_2572);
or U2747 (N_2747,N_2411,N_2552);
nand U2748 (N_2748,N_2438,N_2496);
or U2749 (N_2749,N_2565,N_2495);
nor U2750 (N_2750,N_2599,N_2526);
nor U2751 (N_2751,N_2430,N_2523);
and U2752 (N_2752,N_2500,N_2532);
nand U2753 (N_2753,N_2433,N_2540);
or U2754 (N_2754,N_2455,N_2554);
and U2755 (N_2755,N_2598,N_2481);
xnor U2756 (N_2756,N_2420,N_2581);
or U2757 (N_2757,N_2520,N_2421);
nand U2758 (N_2758,N_2494,N_2458);
xor U2759 (N_2759,N_2447,N_2562);
xor U2760 (N_2760,N_2439,N_2551);
nor U2761 (N_2761,N_2452,N_2546);
nor U2762 (N_2762,N_2430,N_2432);
or U2763 (N_2763,N_2418,N_2467);
nor U2764 (N_2764,N_2497,N_2523);
nor U2765 (N_2765,N_2455,N_2424);
and U2766 (N_2766,N_2479,N_2573);
or U2767 (N_2767,N_2586,N_2584);
nor U2768 (N_2768,N_2454,N_2508);
or U2769 (N_2769,N_2477,N_2468);
and U2770 (N_2770,N_2547,N_2455);
xor U2771 (N_2771,N_2526,N_2471);
and U2772 (N_2772,N_2582,N_2578);
and U2773 (N_2773,N_2482,N_2416);
xor U2774 (N_2774,N_2457,N_2518);
and U2775 (N_2775,N_2494,N_2461);
nand U2776 (N_2776,N_2401,N_2596);
and U2777 (N_2777,N_2544,N_2574);
or U2778 (N_2778,N_2466,N_2409);
nand U2779 (N_2779,N_2541,N_2446);
and U2780 (N_2780,N_2582,N_2544);
and U2781 (N_2781,N_2405,N_2501);
nor U2782 (N_2782,N_2406,N_2561);
nor U2783 (N_2783,N_2497,N_2440);
and U2784 (N_2784,N_2494,N_2449);
xor U2785 (N_2785,N_2520,N_2483);
xor U2786 (N_2786,N_2599,N_2412);
xnor U2787 (N_2787,N_2455,N_2530);
and U2788 (N_2788,N_2447,N_2487);
nor U2789 (N_2789,N_2461,N_2489);
nand U2790 (N_2790,N_2412,N_2507);
xor U2791 (N_2791,N_2474,N_2443);
nor U2792 (N_2792,N_2497,N_2588);
and U2793 (N_2793,N_2561,N_2478);
or U2794 (N_2794,N_2477,N_2588);
and U2795 (N_2795,N_2597,N_2501);
nor U2796 (N_2796,N_2595,N_2488);
nand U2797 (N_2797,N_2473,N_2536);
nor U2798 (N_2798,N_2590,N_2565);
nand U2799 (N_2799,N_2520,N_2528);
and U2800 (N_2800,N_2665,N_2630);
and U2801 (N_2801,N_2717,N_2649);
and U2802 (N_2802,N_2746,N_2606);
nor U2803 (N_2803,N_2730,N_2753);
nor U2804 (N_2804,N_2791,N_2711);
nor U2805 (N_2805,N_2601,N_2778);
or U2806 (N_2806,N_2703,N_2762);
nand U2807 (N_2807,N_2602,N_2627);
nand U2808 (N_2808,N_2623,N_2666);
and U2809 (N_2809,N_2736,N_2757);
or U2810 (N_2810,N_2744,N_2794);
nand U2811 (N_2811,N_2714,N_2716);
nor U2812 (N_2812,N_2770,N_2715);
nand U2813 (N_2813,N_2752,N_2767);
nor U2814 (N_2814,N_2708,N_2719);
or U2815 (N_2815,N_2650,N_2740);
or U2816 (N_2816,N_2760,N_2782);
nand U2817 (N_2817,N_2648,N_2684);
nor U2818 (N_2818,N_2788,N_2751);
nor U2819 (N_2819,N_2631,N_2655);
or U2820 (N_2820,N_2687,N_2670);
nand U2821 (N_2821,N_2776,N_2734);
nand U2822 (N_2822,N_2609,N_2754);
nand U2823 (N_2823,N_2682,N_2636);
or U2824 (N_2824,N_2619,N_2743);
nor U2825 (N_2825,N_2700,N_2621);
nor U2826 (N_2826,N_2620,N_2722);
nor U2827 (N_2827,N_2728,N_2675);
nor U2828 (N_2828,N_2624,N_2610);
and U2829 (N_2829,N_2646,N_2607);
nand U2830 (N_2830,N_2797,N_2726);
nor U2831 (N_2831,N_2685,N_2629);
and U2832 (N_2832,N_2651,N_2706);
and U2833 (N_2833,N_2733,N_2680);
nand U2834 (N_2834,N_2779,N_2694);
nand U2835 (N_2835,N_2677,N_2738);
and U2836 (N_2836,N_2748,N_2605);
nand U2837 (N_2837,N_2656,N_2669);
or U2838 (N_2838,N_2660,N_2683);
and U2839 (N_2839,N_2635,N_2702);
nor U2840 (N_2840,N_2709,N_2732);
nor U2841 (N_2841,N_2608,N_2707);
nand U2842 (N_2842,N_2790,N_2775);
or U2843 (N_2843,N_2637,N_2737);
or U2844 (N_2844,N_2664,N_2699);
and U2845 (N_2845,N_2673,N_2765);
or U2846 (N_2846,N_2720,N_2676);
or U2847 (N_2847,N_2766,N_2735);
nor U2848 (N_2848,N_2710,N_2771);
nor U2849 (N_2849,N_2786,N_2795);
and U2850 (N_2850,N_2727,N_2686);
nand U2851 (N_2851,N_2789,N_2742);
and U2852 (N_2852,N_2641,N_2640);
or U2853 (N_2853,N_2604,N_2611);
and U2854 (N_2854,N_2663,N_2612);
nor U2855 (N_2855,N_2773,N_2696);
or U2856 (N_2856,N_2704,N_2689);
or U2857 (N_2857,N_2756,N_2643);
nand U2858 (N_2858,N_2741,N_2603);
and U2859 (N_2859,N_2692,N_2614);
or U2860 (N_2860,N_2618,N_2783);
nand U2861 (N_2861,N_2600,N_2718);
nand U2862 (N_2862,N_2647,N_2749);
nand U2863 (N_2863,N_2695,N_2638);
nor U2864 (N_2864,N_2799,N_2780);
nor U2865 (N_2865,N_2693,N_2662);
nand U2866 (N_2866,N_2678,N_2764);
nand U2867 (N_2867,N_2721,N_2793);
nor U2868 (N_2868,N_2747,N_2654);
and U2869 (N_2869,N_2690,N_2633);
nor U2870 (N_2870,N_2645,N_2634);
nand U2871 (N_2871,N_2657,N_2616);
nand U2872 (N_2872,N_2768,N_2626);
and U2873 (N_2873,N_2701,N_2615);
or U2874 (N_2874,N_2617,N_2671);
and U2875 (N_2875,N_2758,N_2652);
and U2876 (N_2876,N_2661,N_2691);
nand U2877 (N_2877,N_2613,N_2798);
nand U2878 (N_2878,N_2784,N_2750);
and U2879 (N_2879,N_2731,N_2755);
nor U2880 (N_2880,N_2628,N_2723);
nand U2881 (N_2881,N_2625,N_2759);
or U2882 (N_2882,N_2658,N_2763);
and U2883 (N_2883,N_2632,N_2792);
nand U2884 (N_2884,N_2769,N_2772);
and U2885 (N_2885,N_2745,N_2653);
or U2886 (N_2886,N_2777,N_2774);
or U2887 (N_2887,N_2697,N_2642);
nor U2888 (N_2888,N_2739,N_2659);
nor U2889 (N_2889,N_2796,N_2688);
or U2890 (N_2890,N_2781,N_2667);
and U2891 (N_2891,N_2713,N_2725);
or U2892 (N_2892,N_2639,N_2679);
or U2893 (N_2893,N_2787,N_2705);
and U2894 (N_2894,N_2761,N_2668);
nor U2895 (N_2895,N_2712,N_2785);
nor U2896 (N_2896,N_2729,N_2644);
or U2897 (N_2897,N_2698,N_2672);
or U2898 (N_2898,N_2724,N_2622);
nor U2899 (N_2899,N_2681,N_2674);
nor U2900 (N_2900,N_2678,N_2676);
nand U2901 (N_2901,N_2706,N_2754);
nand U2902 (N_2902,N_2639,N_2788);
or U2903 (N_2903,N_2648,N_2740);
or U2904 (N_2904,N_2786,N_2756);
or U2905 (N_2905,N_2667,N_2617);
xnor U2906 (N_2906,N_2650,N_2759);
or U2907 (N_2907,N_2778,N_2620);
nor U2908 (N_2908,N_2710,N_2691);
or U2909 (N_2909,N_2670,N_2789);
xnor U2910 (N_2910,N_2705,N_2678);
and U2911 (N_2911,N_2680,N_2626);
or U2912 (N_2912,N_2728,N_2603);
nor U2913 (N_2913,N_2758,N_2736);
or U2914 (N_2914,N_2693,N_2732);
and U2915 (N_2915,N_2671,N_2709);
and U2916 (N_2916,N_2628,N_2762);
nand U2917 (N_2917,N_2753,N_2694);
or U2918 (N_2918,N_2634,N_2741);
nand U2919 (N_2919,N_2645,N_2784);
or U2920 (N_2920,N_2617,N_2777);
nor U2921 (N_2921,N_2673,N_2693);
xnor U2922 (N_2922,N_2647,N_2728);
nor U2923 (N_2923,N_2621,N_2726);
and U2924 (N_2924,N_2742,N_2773);
and U2925 (N_2925,N_2629,N_2696);
nor U2926 (N_2926,N_2706,N_2628);
nand U2927 (N_2927,N_2694,N_2783);
or U2928 (N_2928,N_2784,N_2776);
nand U2929 (N_2929,N_2773,N_2628);
and U2930 (N_2930,N_2765,N_2691);
xor U2931 (N_2931,N_2632,N_2702);
or U2932 (N_2932,N_2736,N_2668);
nand U2933 (N_2933,N_2708,N_2627);
nand U2934 (N_2934,N_2634,N_2612);
or U2935 (N_2935,N_2643,N_2688);
nand U2936 (N_2936,N_2733,N_2604);
nor U2937 (N_2937,N_2659,N_2738);
and U2938 (N_2938,N_2779,N_2742);
nand U2939 (N_2939,N_2634,N_2688);
and U2940 (N_2940,N_2637,N_2654);
and U2941 (N_2941,N_2682,N_2618);
xnor U2942 (N_2942,N_2604,N_2774);
or U2943 (N_2943,N_2640,N_2606);
and U2944 (N_2944,N_2684,N_2747);
and U2945 (N_2945,N_2789,N_2664);
and U2946 (N_2946,N_2695,N_2688);
nand U2947 (N_2947,N_2601,N_2600);
and U2948 (N_2948,N_2774,N_2626);
and U2949 (N_2949,N_2614,N_2661);
nand U2950 (N_2950,N_2651,N_2734);
nand U2951 (N_2951,N_2674,N_2609);
nor U2952 (N_2952,N_2714,N_2664);
nand U2953 (N_2953,N_2649,N_2605);
nand U2954 (N_2954,N_2736,N_2613);
and U2955 (N_2955,N_2798,N_2607);
and U2956 (N_2956,N_2758,N_2770);
or U2957 (N_2957,N_2616,N_2661);
nand U2958 (N_2958,N_2657,N_2612);
nand U2959 (N_2959,N_2674,N_2706);
nand U2960 (N_2960,N_2651,N_2759);
and U2961 (N_2961,N_2603,N_2689);
xor U2962 (N_2962,N_2734,N_2702);
nand U2963 (N_2963,N_2684,N_2709);
nor U2964 (N_2964,N_2771,N_2656);
and U2965 (N_2965,N_2703,N_2715);
and U2966 (N_2966,N_2627,N_2791);
nand U2967 (N_2967,N_2641,N_2763);
nor U2968 (N_2968,N_2627,N_2685);
or U2969 (N_2969,N_2678,N_2795);
nand U2970 (N_2970,N_2708,N_2691);
nand U2971 (N_2971,N_2697,N_2726);
nor U2972 (N_2972,N_2695,N_2748);
nor U2973 (N_2973,N_2735,N_2683);
or U2974 (N_2974,N_2601,N_2637);
and U2975 (N_2975,N_2645,N_2719);
nor U2976 (N_2976,N_2775,N_2678);
nand U2977 (N_2977,N_2728,N_2676);
or U2978 (N_2978,N_2601,N_2748);
and U2979 (N_2979,N_2739,N_2635);
or U2980 (N_2980,N_2659,N_2723);
or U2981 (N_2981,N_2624,N_2657);
nand U2982 (N_2982,N_2691,N_2718);
or U2983 (N_2983,N_2644,N_2607);
nor U2984 (N_2984,N_2703,N_2709);
nand U2985 (N_2985,N_2777,N_2624);
or U2986 (N_2986,N_2718,N_2608);
nand U2987 (N_2987,N_2690,N_2659);
and U2988 (N_2988,N_2696,N_2636);
nor U2989 (N_2989,N_2746,N_2617);
and U2990 (N_2990,N_2694,N_2746);
nor U2991 (N_2991,N_2698,N_2620);
nand U2992 (N_2992,N_2606,N_2757);
and U2993 (N_2993,N_2793,N_2672);
or U2994 (N_2994,N_2610,N_2771);
or U2995 (N_2995,N_2628,N_2600);
or U2996 (N_2996,N_2788,N_2610);
and U2997 (N_2997,N_2777,N_2754);
and U2998 (N_2998,N_2699,N_2660);
and U2999 (N_2999,N_2784,N_2653);
nor U3000 (N_3000,N_2810,N_2859);
and U3001 (N_3001,N_2831,N_2827);
nand U3002 (N_3002,N_2936,N_2807);
nand U3003 (N_3003,N_2874,N_2980);
nand U3004 (N_3004,N_2972,N_2938);
nor U3005 (N_3005,N_2843,N_2814);
or U3006 (N_3006,N_2824,N_2933);
nor U3007 (N_3007,N_2905,N_2985);
nand U3008 (N_3008,N_2925,N_2982);
or U3009 (N_3009,N_2840,N_2947);
nand U3010 (N_3010,N_2823,N_2955);
nand U3011 (N_3011,N_2849,N_2852);
and U3012 (N_3012,N_2954,N_2819);
nor U3013 (N_3013,N_2847,N_2911);
or U3014 (N_3014,N_2987,N_2946);
nor U3015 (N_3015,N_2853,N_2809);
nor U3016 (N_3016,N_2971,N_2945);
or U3017 (N_3017,N_2834,N_2991);
nand U3018 (N_3018,N_2973,N_2901);
or U3019 (N_3019,N_2988,N_2963);
nor U3020 (N_3020,N_2996,N_2943);
nand U3021 (N_3021,N_2895,N_2886);
or U3022 (N_3022,N_2908,N_2956);
nand U3023 (N_3023,N_2885,N_2801);
or U3024 (N_3024,N_2896,N_2941);
and U3025 (N_3025,N_2993,N_2870);
nand U3026 (N_3026,N_2918,N_2957);
or U3027 (N_3027,N_2913,N_2889);
nand U3028 (N_3028,N_2922,N_2898);
nor U3029 (N_3029,N_2872,N_2902);
or U3030 (N_3030,N_2924,N_2999);
nor U3031 (N_3031,N_2854,N_2937);
and U3032 (N_3032,N_2928,N_2959);
and U3033 (N_3033,N_2828,N_2930);
nor U3034 (N_3034,N_2934,N_2805);
and U3035 (N_3035,N_2976,N_2825);
and U3036 (N_3036,N_2960,N_2951);
and U3037 (N_3037,N_2935,N_2906);
and U3038 (N_3038,N_2844,N_2961);
or U3039 (N_3039,N_2888,N_2838);
and U3040 (N_3040,N_2833,N_2931);
and U3041 (N_3041,N_2848,N_2904);
nand U3042 (N_3042,N_2974,N_2952);
nor U3043 (N_3043,N_2989,N_2835);
nor U3044 (N_3044,N_2986,N_2890);
or U3045 (N_3045,N_2837,N_2821);
and U3046 (N_3046,N_2806,N_2968);
and U3047 (N_3047,N_2940,N_2923);
nand U3048 (N_3048,N_2939,N_2871);
nor U3049 (N_3049,N_2846,N_2860);
or U3050 (N_3050,N_2879,N_2892);
xor U3051 (N_3051,N_2893,N_2832);
nor U3052 (N_3052,N_2994,N_2808);
or U3053 (N_3053,N_2851,N_2803);
nor U3054 (N_3054,N_2899,N_2949);
xor U3055 (N_3055,N_2813,N_2950);
nor U3056 (N_3056,N_2897,N_2862);
nand U3057 (N_3057,N_2815,N_2983);
nand U3058 (N_3058,N_2811,N_2962);
and U3059 (N_3059,N_2997,N_2894);
and U3060 (N_3060,N_2900,N_2919);
nand U3061 (N_3061,N_2917,N_2907);
and U3062 (N_3062,N_2975,N_2867);
and U3063 (N_3063,N_2882,N_2912);
nand U3064 (N_3064,N_2878,N_2857);
and U3065 (N_3065,N_2964,N_2884);
nand U3066 (N_3066,N_2802,N_2926);
and U3067 (N_3067,N_2816,N_2812);
nor U3068 (N_3068,N_2869,N_2909);
or U3069 (N_3069,N_2861,N_2842);
or U3070 (N_3070,N_2998,N_2866);
and U3071 (N_3071,N_2864,N_2979);
nand U3072 (N_3072,N_2863,N_2995);
or U3073 (N_3073,N_2829,N_2858);
nor U3074 (N_3074,N_2880,N_2932);
or U3075 (N_3075,N_2883,N_2992);
and U3076 (N_3076,N_2817,N_2826);
nor U3077 (N_3077,N_2914,N_2865);
and U3078 (N_3078,N_2910,N_2984);
nor U3079 (N_3079,N_2948,N_2929);
or U3080 (N_3080,N_2804,N_2881);
or U3081 (N_3081,N_2820,N_2841);
and U3082 (N_3082,N_2942,N_2921);
nor U3083 (N_3083,N_2920,N_2873);
or U3084 (N_3084,N_2927,N_2978);
nor U3085 (N_3085,N_2876,N_2845);
and U3086 (N_3086,N_2877,N_2818);
nand U3087 (N_3087,N_2822,N_2868);
nand U3088 (N_3088,N_2830,N_2990);
and U3089 (N_3089,N_2965,N_2903);
nor U3090 (N_3090,N_2839,N_2887);
nor U3091 (N_3091,N_2856,N_2953);
and U3092 (N_3092,N_2966,N_2967);
nor U3093 (N_3093,N_2915,N_2977);
nand U3094 (N_3094,N_2969,N_2981);
and U3095 (N_3095,N_2850,N_2944);
nand U3096 (N_3096,N_2916,N_2891);
and U3097 (N_3097,N_2970,N_2836);
and U3098 (N_3098,N_2875,N_2855);
and U3099 (N_3099,N_2800,N_2958);
nor U3100 (N_3100,N_2836,N_2831);
nor U3101 (N_3101,N_2991,N_2923);
nor U3102 (N_3102,N_2980,N_2974);
or U3103 (N_3103,N_2895,N_2945);
nor U3104 (N_3104,N_2990,N_2800);
or U3105 (N_3105,N_2807,N_2966);
nand U3106 (N_3106,N_2860,N_2995);
and U3107 (N_3107,N_2837,N_2927);
and U3108 (N_3108,N_2934,N_2926);
and U3109 (N_3109,N_2857,N_2916);
nand U3110 (N_3110,N_2866,N_2925);
nor U3111 (N_3111,N_2961,N_2920);
nor U3112 (N_3112,N_2948,N_2898);
nor U3113 (N_3113,N_2923,N_2802);
nand U3114 (N_3114,N_2877,N_2854);
nand U3115 (N_3115,N_2937,N_2899);
and U3116 (N_3116,N_2814,N_2953);
or U3117 (N_3117,N_2819,N_2957);
and U3118 (N_3118,N_2844,N_2907);
nand U3119 (N_3119,N_2869,N_2965);
nand U3120 (N_3120,N_2855,N_2814);
nand U3121 (N_3121,N_2982,N_2818);
nand U3122 (N_3122,N_2864,N_2925);
nor U3123 (N_3123,N_2999,N_2884);
and U3124 (N_3124,N_2979,N_2950);
or U3125 (N_3125,N_2860,N_2837);
and U3126 (N_3126,N_2879,N_2923);
nand U3127 (N_3127,N_2871,N_2992);
and U3128 (N_3128,N_2982,N_2984);
and U3129 (N_3129,N_2871,N_2808);
or U3130 (N_3130,N_2868,N_2851);
and U3131 (N_3131,N_2995,N_2854);
or U3132 (N_3132,N_2839,N_2809);
nand U3133 (N_3133,N_2874,N_2833);
nand U3134 (N_3134,N_2850,N_2929);
and U3135 (N_3135,N_2990,N_2831);
nand U3136 (N_3136,N_2966,N_2815);
nand U3137 (N_3137,N_2853,N_2981);
and U3138 (N_3138,N_2829,N_2960);
and U3139 (N_3139,N_2861,N_2876);
nand U3140 (N_3140,N_2836,N_2837);
nor U3141 (N_3141,N_2978,N_2815);
and U3142 (N_3142,N_2839,N_2812);
and U3143 (N_3143,N_2993,N_2853);
and U3144 (N_3144,N_2817,N_2998);
or U3145 (N_3145,N_2834,N_2942);
nand U3146 (N_3146,N_2994,N_2918);
nor U3147 (N_3147,N_2965,N_2832);
nand U3148 (N_3148,N_2934,N_2949);
and U3149 (N_3149,N_2868,N_2999);
nand U3150 (N_3150,N_2922,N_2835);
nand U3151 (N_3151,N_2957,N_2856);
and U3152 (N_3152,N_2882,N_2830);
and U3153 (N_3153,N_2953,N_2944);
or U3154 (N_3154,N_2897,N_2919);
or U3155 (N_3155,N_2830,N_2883);
nand U3156 (N_3156,N_2932,N_2885);
nor U3157 (N_3157,N_2979,N_2932);
or U3158 (N_3158,N_2946,N_2876);
nor U3159 (N_3159,N_2820,N_2906);
nor U3160 (N_3160,N_2939,N_2953);
and U3161 (N_3161,N_2970,N_2846);
or U3162 (N_3162,N_2989,N_2943);
or U3163 (N_3163,N_2972,N_2877);
and U3164 (N_3164,N_2837,N_2902);
and U3165 (N_3165,N_2800,N_2904);
nand U3166 (N_3166,N_2892,N_2807);
nand U3167 (N_3167,N_2840,N_2879);
or U3168 (N_3168,N_2823,N_2891);
nor U3169 (N_3169,N_2862,N_2863);
nor U3170 (N_3170,N_2949,N_2895);
and U3171 (N_3171,N_2927,N_2854);
xor U3172 (N_3172,N_2968,N_2979);
and U3173 (N_3173,N_2838,N_2989);
nor U3174 (N_3174,N_2888,N_2948);
nand U3175 (N_3175,N_2955,N_2880);
nand U3176 (N_3176,N_2851,N_2812);
and U3177 (N_3177,N_2891,N_2807);
nor U3178 (N_3178,N_2884,N_2968);
nand U3179 (N_3179,N_2897,N_2983);
nor U3180 (N_3180,N_2961,N_2838);
nand U3181 (N_3181,N_2898,N_2907);
nand U3182 (N_3182,N_2835,N_2867);
and U3183 (N_3183,N_2878,N_2972);
nand U3184 (N_3184,N_2990,N_2928);
nand U3185 (N_3185,N_2835,N_2964);
or U3186 (N_3186,N_2941,N_2813);
nand U3187 (N_3187,N_2949,N_2821);
and U3188 (N_3188,N_2818,N_2843);
and U3189 (N_3189,N_2981,N_2946);
nor U3190 (N_3190,N_2912,N_2894);
and U3191 (N_3191,N_2872,N_2847);
nand U3192 (N_3192,N_2856,N_2813);
nor U3193 (N_3193,N_2949,N_2966);
and U3194 (N_3194,N_2906,N_2842);
or U3195 (N_3195,N_2977,N_2992);
nor U3196 (N_3196,N_2841,N_2888);
nand U3197 (N_3197,N_2984,N_2879);
nor U3198 (N_3198,N_2917,N_2941);
nor U3199 (N_3199,N_2933,N_2891);
or U3200 (N_3200,N_3030,N_3102);
nor U3201 (N_3201,N_3074,N_3063);
nor U3202 (N_3202,N_3125,N_3129);
and U3203 (N_3203,N_3121,N_3033);
and U3204 (N_3204,N_3058,N_3115);
and U3205 (N_3205,N_3167,N_3156);
nor U3206 (N_3206,N_3044,N_3108);
nand U3207 (N_3207,N_3158,N_3169);
nand U3208 (N_3208,N_3154,N_3045);
and U3209 (N_3209,N_3164,N_3008);
nor U3210 (N_3210,N_3029,N_3168);
and U3211 (N_3211,N_3010,N_3061);
and U3212 (N_3212,N_3020,N_3130);
or U3213 (N_3213,N_3054,N_3021);
xor U3214 (N_3214,N_3174,N_3098);
or U3215 (N_3215,N_3134,N_3065);
nor U3216 (N_3216,N_3006,N_3152);
or U3217 (N_3217,N_3079,N_3056);
or U3218 (N_3218,N_3144,N_3180);
nor U3219 (N_3219,N_3175,N_3137);
nand U3220 (N_3220,N_3188,N_3172);
nor U3221 (N_3221,N_3163,N_3135);
nor U3222 (N_3222,N_3072,N_3059);
nand U3223 (N_3223,N_3018,N_3089);
nand U3224 (N_3224,N_3087,N_3017);
or U3225 (N_3225,N_3012,N_3126);
nor U3226 (N_3226,N_3050,N_3091);
or U3227 (N_3227,N_3081,N_3022);
nor U3228 (N_3228,N_3093,N_3109);
nor U3229 (N_3229,N_3042,N_3097);
nand U3230 (N_3230,N_3197,N_3103);
and U3231 (N_3231,N_3067,N_3104);
nand U3232 (N_3232,N_3049,N_3159);
and U3233 (N_3233,N_3016,N_3034);
nand U3234 (N_3234,N_3046,N_3155);
nand U3235 (N_3235,N_3083,N_3119);
or U3236 (N_3236,N_3005,N_3090);
and U3237 (N_3237,N_3062,N_3078);
nand U3238 (N_3238,N_3001,N_3051);
and U3239 (N_3239,N_3000,N_3075);
nand U3240 (N_3240,N_3100,N_3032);
nor U3241 (N_3241,N_3057,N_3092);
nand U3242 (N_3242,N_3182,N_3195);
or U3243 (N_3243,N_3198,N_3181);
nor U3244 (N_3244,N_3039,N_3147);
nand U3245 (N_3245,N_3019,N_3053);
nand U3246 (N_3246,N_3055,N_3040);
or U3247 (N_3247,N_3179,N_3166);
nor U3248 (N_3248,N_3124,N_3086);
nand U3249 (N_3249,N_3114,N_3142);
and U3250 (N_3250,N_3009,N_3190);
nand U3251 (N_3251,N_3069,N_3004);
or U3252 (N_3252,N_3191,N_3048);
nor U3253 (N_3253,N_3196,N_3106);
and U3254 (N_3254,N_3150,N_3025);
nor U3255 (N_3255,N_3096,N_3111);
nor U3256 (N_3256,N_3128,N_3105);
or U3257 (N_3257,N_3002,N_3101);
and U3258 (N_3258,N_3118,N_3047);
nand U3259 (N_3259,N_3070,N_3038);
nor U3260 (N_3260,N_3189,N_3178);
and U3261 (N_3261,N_3066,N_3107);
and U3262 (N_3262,N_3088,N_3173);
or U3263 (N_3263,N_3077,N_3143);
nor U3264 (N_3264,N_3146,N_3171);
nor U3265 (N_3265,N_3199,N_3183);
and U3266 (N_3266,N_3116,N_3043);
nor U3267 (N_3267,N_3145,N_3138);
or U3268 (N_3268,N_3113,N_3064);
or U3269 (N_3269,N_3160,N_3133);
and U3270 (N_3270,N_3148,N_3068);
and U3271 (N_3271,N_3015,N_3071);
nand U3272 (N_3272,N_3136,N_3177);
and U3273 (N_3273,N_3094,N_3193);
nor U3274 (N_3274,N_3139,N_3112);
nand U3275 (N_3275,N_3003,N_3122);
and U3276 (N_3276,N_3085,N_3157);
nor U3277 (N_3277,N_3024,N_3060);
or U3278 (N_3278,N_3011,N_3185);
and U3279 (N_3279,N_3162,N_3170);
nor U3280 (N_3280,N_3110,N_3026);
nor U3281 (N_3281,N_3013,N_3023);
nand U3282 (N_3282,N_3149,N_3014);
and U3283 (N_3283,N_3095,N_3192);
or U3284 (N_3284,N_3076,N_3176);
or U3285 (N_3285,N_3127,N_3099);
and U3286 (N_3286,N_3184,N_3117);
and U3287 (N_3287,N_3194,N_3123);
nand U3288 (N_3288,N_3161,N_3028);
nor U3289 (N_3289,N_3186,N_3165);
nand U3290 (N_3290,N_3084,N_3036);
and U3291 (N_3291,N_3132,N_3140);
and U3292 (N_3292,N_3151,N_3120);
or U3293 (N_3293,N_3035,N_3073);
nand U3294 (N_3294,N_3141,N_3031);
nand U3295 (N_3295,N_3153,N_3082);
xnor U3296 (N_3296,N_3131,N_3080);
nor U3297 (N_3297,N_3052,N_3187);
or U3298 (N_3298,N_3007,N_3041);
nand U3299 (N_3299,N_3027,N_3037);
and U3300 (N_3300,N_3124,N_3136);
or U3301 (N_3301,N_3139,N_3103);
and U3302 (N_3302,N_3134,N_3119);
and U3303 (N_3303,N_3190,N_3104);
nor U3304 (N_3304,N_3063,N_3059);
or U3305 (N_3305,N_3163,N_3186);
nor U3306 (N_3306,N_3071,N_3116);
nor U3307 (N_3307,N_3137,N_3141);
and U3308 (N_3308,N_3126,N_3112);
nand U3309 (N_3309,N_3177,N_3025);
or U3310 (N_3310,N_3008,N_3010);
nor U3311 (N_3311,N_3015,N_3197);
or U3312 (N_3312,N_3184,N_3094);
or U3313 (N_3313,N_3189,N_3017);
and U3314 (N_3314,N_3154,N_3041);
nand U3315 (N_3315,N_3086,N_3173);
or U3316 (N_3316,N_3163,N_3152);
and U3317 (N_3317,N_3036,N_3007);
and U3318 (N_3318,N_3103,N_3142);
and U3319 (N_3319,N_3054,N_3159);
and U3320 (N_3320,N_3095,N_3029);
and U3321 (N_3321,N_3146,N_3172);
or U3322 (N_3322,N_3077,N_3123);
or U3323 (N_3323,N_3153,N_3134);
and U3324 (N_3324,N_3082,N_3106);
xnor U3325 (N_3325,N_3097,N_3148);
nor U3326 (N_3326,N_3061,N_3094);
or U3327 (N_3327,N_3151,N_3018);
nand U3328 (N_3328,N_3083,N_3001);
nand U3329 (N_3329,N_3038,N_3030);
or U3330 (N_3330,N_3144,N_3174);
nand U3331 (N_3331,N_3147,N_3057);
or U3332 (N_3332,N_3081,N_3011);
xor U3333 (N_3333,N_3026,N_3119);
nand U3334 (N_3334,N_3066,N_3127);
and U3335 (N_3335,N_3179,N_3007);
nand U3336 (N_3336,N_3172,N_3176);
nor U3337 (N_3337,N_3127,N_3004);
and U3338 (N_3338,N_3190,N_3148);
xnor U3339 (N_3339,N_3010,N_3119);
nor U3340 (N_3340,N_3195,N_3132);
or U3341 (N_3341,N_3127,N_3176);
nand U3342 (N_3342,N_3175,N_3172);
nor U3343 (N_3343,N_3058,N_3153);
and U3344 (N_3344,N_3182,N_3070);
nor U3345 (N_3345,N_3064,N_3165);
nand U3346 (N_3346,N_3132,N_3133);
and U3347 (N_3347,N_3034,N_3161);
and U3348 (N_3348,N_3132,N_3130);
nor U3349 (N_3349,N_3155,N_3132);
or U3350 (N_3350,N_3197,N_3040);
and U3351 (N_3351,N_3087,N_3151);
or U3352 (N_3352,N_3140,N_3113);
xor U3353 (N_3353,N_3197,N_3088);
nand U3354 (N_3354,N_3123,N_3126);
nand U3355 (N_3355,N_3120,N_3019);
and U3356 (N_3356,N_3064,N_3103);
nor U3357 (N_3357,N_3199,N_3045);
and U3358 (N_3358,N_3063,N_3113);
and U3359 (N_3359,N_3086,N_3037);
and U3360 (N_3360,N_3180,N_3049);
and U3361 (N_3361,N_3091,N_3008);
and U3362 (N_3362,N_3147,N_3080);
nand U3363 (N_3363,N_3190,N_3146);
or U3364 (N_3364,N_3032,N_3157);
or U3365 (N_3365,N_3085,N_3148);
nand U3366 (N_3366,N_3064,N_3169);
and U3367 (N_3367,N_3068,N_3062);
nand U3368 (N_3368,N_3102,N_3134);
nand U3369 (N_3369,N_3051,N_3025);
nand U3370 (N_3370,N_3106,N_3130);
nand U3371 (N_3371,N_3106,N_3098);
nor U3372 (N_3372,N_3018,N_3183);
nand U3373 (N_3373,N_3183,N_3144);
and U3374 (N_3374,N_3195,N_3067);
or U3375 (N_3375,N_3126,N_3097);
nor U3376 (N_3376,N_3167,N_3068);
or U3377 (N_3377,N_3177,N_3045);
or U3378 (N_3378,N_3088,N_3087);
nand U3379 (N_3379,N_3124,N_3029);
xor U3380 (N_3380,N_3006,N_3165);
nor U3381 (N_3381,N_3055,N_3064);
or U3382 (N_3382,N_3090,N_3029);
nand U3383 (N_3383,N_3185,N_3075);
nand U3384 (N_3384,N_3173,N_3103);
nand U3385 (N_3385,N_3108,N_3011);
or U3386 (N_3386,N_3045,N_3117);
and U3387 (N_3387,N_3109,N_3197);
nand U3388 (N_3388,N_3138,N_3004);
and U3389 (N_3389,N_3070,N_3134);
or U3390 (N_3390,N_3126,N_3103);
nand U3391 (N_3391,N_3089,N_3003);
and U3392 (N_3392,N_3073,N_3014);
nand U3393 (N_3393,N_3091,N_3074);
and U3394 (N_3394,N_3120,N_3059);
or U3395 (N_3395,N_3141,N_3100);
or U3396 (N_3396,N_3055,N_3130);
nor U3397 (N_3397,N_3092,N_3107);
nand U3398 (N_3398,N_3168,N_3131);
nand U3399 (N_3399,N_3121,N_3085);
xor U3400 (N_3400,N_3396,N_3234);
and U3401 (N_3401,N_3227,N_3260);
nand U3402 (N_3402,N_3258,N_3253);
nand U3403 (N_3403,N_3340,N_3314);
xor U3404 (N_3404,N_3301,N_3263);
and U3405 (N_3405,N_3341,N_3332);
or U3406 (N_3406,N_3206,N_3369);
and U3407 (N_3407,N_3293,N_3395);
and U3408 (N_3408,N_3245,N_3317);
and U3409 (N_3409,N_3330,N_3384);
and U3410 (N_3410,N_3233,N_3304);
or U3411 (N_3411,N_3343,N_3283);
nor U3412 (N_3412,N_3315,N_3347);
and U3413 (N_3413,N_3281,N_3243);
nor U3414 (N_3414,N_3381,N_3328);
or U3415 (N_3415,N_3289,N_3271);
or U3416 (N_3416,N_3251,N_3345);
and U3417 (N_3417,N_3264,N_3241);
and U3418 (N_3418,N_3364,N_3291);
or U3419 (N_3419,N_3305,N_3244);
nand U3420 (N_3420,N_3398,N_3209);
nor U3421 (N_3421,N_3385,N_3382);
nor U3422 (N_3422,N_3360,N_3259);
and U3423 (N_3423,N_3377,N_3276);
nand U3424 (N_3424,N_3316,N_3339);
nor U3425 (N_3425,N_3371,N_3359);
and U3426 (N_3426,N_3270,N_3326);
and U3427 (N_3427,N_3275,N_3361);
and U3428 (N_3428,N_3204,N_3212);
nor U3429 (N_3429,N_3248,N_3284);
and U3430 (N_3430,N_3287,N_3288);
nor U3431 (N_3431,N_3296,N_3285);
nor U3432 (N_3432,N_3318,N_3363);
nor U3433 (N_3433,N_3297,N_3255);
nand U3434 (N_3434,N_3310,N_3223);
or U3435 (N_3435,N_3246,N_3274);
and U3436 (N_3436,N_3311,N_3213);
or U3437 (N_3437,N_3322,N_3257);
nand U3438 (N_3438,N_3390,N_3354);
or U3439 (N_3439,N_3379,N_3217);
or U3440 (N_3440,N_3324,N_3237);
and U3441 (N_3441,N_3211,N_3373);
nand U3442 (N_3442,N_3374,N_3399);
nor U3443 (N_3443,N_3303,N_3355);
and U3444 (N_3444,N_3273,N_3221);
and U3445 (N_3445,N_3358,N_3334);
and U3446 (N_3446,N_3254,N_3350);
xor U3447 (N_3447,N_3307,N_3392);
or U3448 (N_3448,N_3294,N_3319);
nor U3449 (N_3449,N_3321,N_3376);
nand U3450 (N_3450,N_3279,N_3265);
and U3451 (N_3451,N_3368,N_3214);
and U3452 (N_3452,N_3386,N_3247);
and U3453 (N_3453,N_3277,N_3342);
nor U3454 (N_3454,N_3325,N_3229);
nor U3455 (N_3455,N_3292,N_3240);
or U3456 (N_3456,N_3282,N_3250);
xor U3457 (N_3457,N_3300,N_3308);
nand U3458 (N_3458,N_3261,N_3370);
nor U3459 (N_3459,N_3286,N_3249);
and U3460 (N_3460,N_3346,N_3323);
nor U3461 (N_3461,N_3388,N_3329);
nand U3462 (N_3462,N_3266,N_3335);
and U3463 (N_3463,N_3226,N_3239);
and U3464 (N_3464,N_3256,N_3208);
nor U3465 (N_3465,N_3357,N_3224);
nor U3466 (N_3466,N_3383,N_3356);
nor U3467 (N_3467,N_3366,N_3306);
nor U3468 (N_3468,N_3232,N_3230);
nor U3469 (N_3469,N_3397,N_3268);
and U3470 (N_3470,N_3231,N_3394);
nand U3471 (N_3471,N_3200,N_3298);
or U3472 (N_3472,N_3344,N_3380);
nand U3473 (N_3473,N_3372,N_3216);
nor U3474 (N_3474,N_3336,N_3389);
or U3475 (N_3475,N_3313,N_3210);
nand U3476 (N_3476,N_3367,N_3242);
nor U3477 (N_3477,N_3235,N_3331);
nor U3478 (N_3478,N_3353,N_3201);
or U3479 (N_3479,N_3352,N_3365);
or U3480 (N_3480,N_3262,N_3222);
nand U3481 (N_3481,N_3299,N_3228);
nand U3482 (N_3482,N_3280,N_3236);
nor U3483 (N_3483,N_3391,N_3337);
or U3484 (N_3484,N_3290,N_3338);
nand U3485 (N_3485,N_3202,N_3203);
or U3486 (N_3486,N_3215,N_3320);
nor U3487 (N_3487,N_3218,N_3333);
nand U3488 (N_3488,N_3312,N_3348);
nand U3489 (N_3489,N_3302,N_3278);
and U3490 (N_3490,N_3238,N_3252);
nand U3491 (N_3491,N_3378,N_3309);
and U3492 (N_3492,N_3327,N_3387);
nor U3493 (N_3493,N_3269,N_3272);
xnor U3494 (N_3494,N_3267,N_3220);
nor U3495 (N_3495,N_3393,N_3225);
or U3496 (N_3496,N_3351,N_3349);
nand U3497 (N_3497,N_3362,N_3205);
or U3498 (N_3498,N_3375,N_3295);
nand U3499 (N_3499,N_3219,N_3207);
nand U3500 (N_3500,N_3243,N_3375);
and U3501 (N_3501,N_3232,N_3204);
and U3502 (N_3502,N_3237,N_3263);
nor U3503 (N_3503,N_3378,N_3227);
and U3504 (N_3504,N_3311,N_3203);
or U3505 (N_3505,N_3369,N_3344);
nor U3506 (N_3506,N_3318,N_3202);
nand U3507 (N_3507,N_3383,N_3297);
nor U3508 (N_3508,N_3386,N_3262);
nand U3509 (N_3509,N_3384,N_3227);
and U3510 (N_3510,N_3355,N_3347);
nor U3511 (N_3511,N_3262,N_3246);
and U3512 (N_3512,N_3354,N_3370);
and U3513 (N_3513,N_3313,N_3275);
and U3514 (N_3514,N_3258,N_3264);
nor U3515 (N_3515,N_3344,N_3243);
nand U3516 (N_3516,N_3347,N_3300);
nand U3517 (N_3517,N_3380,N_3224);
or U3518 (N_3518,N_3292,N_3235);
and U3519 (N_3519,N_3258,N_3228);
xor U3520 (N_3520,N_3381,N_3227);
nand U3521 (N_3521,N_3293,N_3239);
nand U3522 (N_3522,N_3204,N_3215);
nor U3523 (N_3523,N_3317,N_3370);
and U3524 (N_3524,N_3334,N_3275);
nand U3525 (N_3525,N_3291,N_3287);
or U3526 (N_3526,N_3238,N_3278);
nor U3527 (N_3527,N_3279,N_3242);
or U3528 (N_3528,N_3350,N_3278);
nor U3529 (N_3529,N_3295,N_3318);
and U3530 (N_3530,N_3317,N_3239);
or U3531 (N_3531,N_3339,N_3277);
nor U3532 (N_3532,N_3208,N_3302);
or U3533 (N_3533,N_3284,N_3234);
or U3534 (N_3534,N_3358,N_3395);
or U3535 (N_3535,N_3257,N_3230);
nor U3536 (N_3536,N_3260,N_3305);
and U3537 (N_3537,N_3305,N_3334);
nor U3538 (N_3538,N_3386,N_3396);
or U3539 (N_3539,N_3310,N_3342);
nand U3540 (N_3540,N_3391,N_3333);
and U3541 (N_3541,N_3379,N_3362);
nand U3542 (N_3542,N_3361,N_3204);
xor U3543 (N_3543,N_3328,N_3264);
nand U3544 (N_3544,N_3257,N_3287);
or U3545 (N_3545,N_3378,N_3323);
nand U3546 (N_3546,N_3294,N_3323);
nand U3547 (N_3547,N_3279,N_3378);
or U3548 (N_3548,N_3262,N_3349);
nor U3549 (N_3549,N_3265,N_3285);
nor U3550 (N_3550,N_3361,N_3358);
and U3551 (N_3551,N_3220,N_3204);
and U3552 (N_3552,N_3331,N_3214);
or U3553 (N_3553,N_3300,N_3343);
nor U3554 (N_3554,N_3273,N_3348);
nor U3555 (N_3555,N_3259,N_3252);
nand U3556 (N_3556,N_3210,N_3259);
xnor U3557 (N_3557,N_3342,N_3213);
or U3558 (N_3558,N_3325,N_3281);
nand U3559 (N_3559,N_3215,N_3285);
nand U3560 (N_3560,N_3271,N_3298);
nand U3561 (N_3561,N_3316,N_3373);
and U3562 (N_3562,N_3349,N_3300);
and U3563 (N_3563,N_3370,N_3294);
nand U3564 (N_3564,N_3205,N_3359);
nand U3565 (N_3565,N_3200,N_3233);
and U3566 (N_3566,N_3252,N_3276);
nand U3567 (N_3567,N_3241,N_3255);
or U3568 (N_3568,N_3303,N_3364);
or U3569 (N_3569,N_3223,N_3242);
and U3570 (N_3570,N_3308,N_3280);
and U3571 (N_3571,N_3352,N_3287);
or U3572 (N_3572,N_3339,N_3385);
nand U3573 (N_3573,N_3216,N_3299);
and U3574 (N_3574,N_3243,N_3349);
nand U3575 (N_3575,N_3366,N_3360);
and U3576 (N_3576,N_3387,N_3334);
and U3577 (N_3577,N_3356,N_3234);
and U3578 (N_3578,N_3295,N_3389);
and U3579 (N_3579,N_3327,N_3352);
nand U3580 (N_3580,N_3380,N_3204);
nand U3581 (N_3581,N_3228,N_3370);
or U3582 (N_3582,N_3255,N_3223);
nor U3583 (N_3583,N_3229,N_3377);
and U3584 (N_3584,N_3352,N_3308);
and U3585 (N_3585,N_3275,N_3206);
and U3586 (N_3586,N_3271,N_3338);
nand U3587 (N_3587,N_3296,N_3367);
nor U3588 (N_3588,N_3235,N_3343);
nand U3589 (N_3589,N_3210,N_3310);
or U3590 (N_3590,N_3359,N_3296);
and U3591 (N_3591,N_3298,N_3392);
xnor U3592 (N_3592,N_3378,N_3254);
nand U3593 (N_3593,N_3340,N_3202);
and U3594 (N_3594,N_3285,N_3314);
nor U3595 (N_3595,N_3233,N_3270);
and U3596 (N_3596,N_3320,N_3309);
or U3597 (N_3597,N_3396,N_3215);
nand U3598 (N_3598,N_3224,N_3385);
nor U3599 (N_3599,N_3319,N_3298);
and U3600 (N_3600,N_3533,N_3560);
nand U3601 (N_3601,N_3597,N_3402);
and U3602 (N_3602,N_3505,N_3486);
and U3603 (N_3603,N_3499,N_3500);
nand U3604 (N_3604,N_3582,N_3407);
and U3605 (N_3605,N_3418,N_3578);
or U3606 (N_3606,N_3550,N_3516);
nor U3607 (N_3607,N_3453,N_3530);
nor U3608 (N_3608,N_3531,N_3542);
nor U3609 (N_3609,N_3408,N_3445);
nor U3610 (N_3610,N_3462,N_3569);
or U3611 (N_3611,N_3434,N_3548);
and U3612 (N_3612,N_3413,N_3591);
or U3613 (N_3613,N_3545,N_3425);
or U3614 (N_3614,N_3441,N_3404);
nor U3615 (N_3615,N_3518,N_3457);
nand U3616 (N_3616,N_3464,N_3543);
and U3617 (N_3617,N_3567,N_3556);
or U3618 (N_3618,N_3594,N_3429);
nand U3619 (N_3619,N_3563,N_3451);
or U3620 (N_3620,N_3561,N_3501);
nand U3621 (N_3621,N_3428,N_3554);
nor U3622 (N_3622,N_3571,N_3463);
or U3623 (N_3623,N_3474,N_3490);
nand U3624 (N_3624,N_3480,N_3482);
nor U3625 (N_3625,N_3519,N_3583);
and U3626 (N_3626,N_3585,N_3485);
nand U3627 (N_3627,N_3452,N_3469);
nand U3628 (N_3628,N_3403,N_3551);
or U3629 (N_3629,N_3491,N_3454);
and U3630 (N_3630,N_3468,N_3443);
and U3631 (N_3631,N_3430,N_3562);
and U3632 (N_3632,N_3587,N_3498);
or U3633 (N_3633,N_3524,N_3546);
or U3634 (N_3634,N_3477,N_3446);
nand U3635 (N_3635,N_3539,N_3461);
and U3636 (N_3636,N_3460,N_3424);
xor U3637 (N_3637,N_3547,N_3431);
nor U3638 (N_3638,N_3590,N_3416);
nor U3639 (N_3639,N_3552,N_3592);
nand U3640 (N_3640,N_3433,N_3510);
and U3641 (N_3641,N_3527,N_3442);
nor U3642 (N_3642,N_3572,N_3577);
nor U3643 (N_3643,N_3419,N_3483);
nand U3644 (N_3644,N_3496,N_3448);
or U3645 (N_3645,N_3450,N_3534);
and U3646 (N_3646,N_3414,N_3525);
xnor U3647 (N_3647,N_3568,N_3432);
nor U3648 (N_3648,N_3536,N_3549);
and U3649 (N_3649,N_3555,N_3508);
and U3650 (N_3650,N_3439,N_3493);
and U3651 (N_3651,N_3580,N_3406);
and U3652 (N_3652,N_3576,N_3514);
or U3653 (N_3653,N_3471,N_3579);
nor U3654 (N_3654,N_3509,N_3478);
and U3655 (N_3655,N_3427,N_3564);
or U3656 (N_3656,N_3589,N_3574);
nor U3657 (N_3657,N_3488,N_3401);
nand U3658 (N_3658,N_3532,N_3517);
nor U3659 (N_3659,N_3558,N_3422);
nor U3660 (N_3660,N_3459,N_3405);
or U3661 (N_3661,N_3476,N_3456);
nor U3662 (N_3662,N_3523,N_3503);
or U3663 (N_3663,N_3540,N_3449);
or U3664 (N_3664,N_3470,N_3455);
nor U3665 (N_3665,N_3467,N_3444);
nor U3666 (N_3666,N_3495,N_3497);
and U3667 (N_3667,N_3410,N_3421);
and U3668 (N_3668,N_3557,N_3420);
nand U3669 (N_3669,N_3595,N_3596);
nand U3670 (N_3670,N_3599,N_3479);
nand U3671 (N_3671,N_3487,N_3400);
and U3672 (N_3672,N_3570,N_3573);
and U3673 (N_3673,N_3438,N_3489);
or U3674 (N_3674,N_3507,N_3411);
or U3675 (N_3675,N_3598,N_3437);
and U3676 (N_3676,N_3521,N_3565);
nand U3677 (N_3677,N_3472,N_3473);
nor U3678 (N_3678,N_3436,N_3440);
nor U3679 (N_3679,N_3586,N_3541);
and U3680 (N_3680,N_3504,N_3584);
nor U3681 (N_3681,N_3494,N_3593);
nand U3682 (N_3682,N_3435,N_3522);
nor U3683 (N_3683,N_3544,N_3484);
nand U3684 (N_3684,N_3538,N_3520);
nand U3685 (N_3685,N_3447,N_3502);
and U3686 (N_3686,N_3458,N_3423);
nand U3687 (N_3687,N_3506,N_3412);
and U3688 (N_3688,N_3475,N_3415);
nor U3689 (N_3689,N_3528,N_3553);
nor U3690 (N_3690,N_3515,N_3535);
and U3691 (N_3691,N_3529,N_3481);
nand U3692 (N_3692,N_3465,N_3426);
and U3693 (N_3693,N_3559,N_3566);
or U3694 (N_3694,N_3417,N_3526);
or U3695 (N_3695,N_3409,N_3512);
or U3696 (N_3696,N_3513,N_3575);
nor U3697 (N_3697,N_3466,N_3537);
and U3698 (N_3698,N_3581,N_3492);
and U3699 (N_3699,N_3588,N_3511);
nor U3700 (N_3700,N_3531,N_3420);
and U3701 (N_3701,N_3442,N_3590);
nor U3702 (N_3702,N_3438,N_3503);
nor U3703 (N_3703,N_3583,N_3510);
or U3704 (N_3704,N_3460,N_3551);
and U3705 (N_3705,N_3478,N_3525);
xnor U3706 (N_3706,N_3472,N_3416);
or U3707 (N_3707,N_3445,N_3412);
nor U3708 (N_3708,N_3440,N_3406);
nand U3709 (N_3709,N_3578,N_3415);
and U3710 (N_3710,N_3418,N_3552);
or U3711 (N_3711,N_3467,N_3513);
or U3712 (N_3712,N_3477,N_3533);
nor U3713 (N_3713,N_3480,N_3573);
nand U3714 (N_3714,N_3426,N_3531);
or U3715 (N_3715,N_3463,N_3562);
nor U3716 (N_3716,N_3475,N_3555);
nand U3717 (N_3717,N_3434,N_3457);
or U3718 (N_3718,N_3548,N_3443);
nor U3719 (N_3719,N_3535,N_3565);
nand U3720 (N_3720,N_3501,N_3558);
or U3721 (N_3721,N_3480,N_3472);
or U3722 (N_3722,N_3524,N_3492);
nor U3723 (N_3723,N_3549,N_3458);
nand U3724 (N_3724,N_3415,N_3543);
nand U3725 (N_3725,N_3457,N_3515);
nand U3726 (N_3726,N_3412,N_3431);
or U3727 (N_3727,N_3595,N_3406);
nand U3728 (N_3728,N_3481,N_3562);
nor U3729 (N_3729,N_3419,N_3410);
nor U3730 (N_3730,N_3577,N_3450);
and U3731 (N_3731,N_3542,N_3454);
or U3732 (N_3732,N_3507,N_3405);
and U3733 (N_3733,N_3437,N_3407);
or U3734 (N_3734,N_3499,N_3510);
nand U3735 (N_3735,N_3496,N_3567);
nand U3736 (N_3736,N_3479,N_3436);
nor U3737 (N_3737,N_3436,N_3583);
nor U3738 (N_3738,N_3423,N_3564);
and U3739 (N_3739,N_3488,N_3449);
or U3740 (N_3740,N_3596,N_3417);
and U3741 (N_3741,N_3465,N_3425);
and U3742 (N_3742,N_3497,N_3514);
or U3743 (N_3743,N_3440,N_3431);
or U3744 (N_3744,N_3591,N_3442);
or U3745 (N_3745,N_3475,N_3454);
and U3746 (N_3746,N_3426,N_3478);
xnor U3747 (N_3747,N_3506,N_3519);
nor U3748 (N_3748,N_3486,N_3409);
nand U3749 (N_3749,N_3548,N_3499);
and U3750 (N_3750,N_3529,N_3557);
and U3751 (N_3751,N_3546,N_3539);
and U3752 (N_3752,N_3473,N_3587);
nand U3753 (N_3753,N_3421,N_3505);
and U3754 (N_3754,N_3484,N_3452);
nor U3755 (N_3755,N_3449,N_3451);
nand U3756 (N_3756,N_3483,N_3410);
nand U3757 (N_3757,N_3516,N_3484);
or U3758 (N_3758,N_3492,N_3494);
and U3759 (N_3759,N_3556,N_3422);
nor U3760 (N_3760,N_3509,N_3440);
nor U3761 (N_3761,N_3582,N_3490);
and U3762 (N_3762,N_3433,N_3453);
nor U3763 (N_3763,N_3577,N_3586);
nor U3764 (N_3764,N_3587,N_3494);
nor U3765 (N_3765,N_3499,N_3448);
and U3766 (N_3766,N_3581,N_3495);
nand U3767 (N_3767,N_3558,N_3424);
or U3768 (N_3768,N_3599,N_3440);
nor U3769 (N_3769,N_3508,N_3473);
nand U3770 (N_3770,N_3591,N_3583);
nor U3771 (N_3771,N_3425,N_3575);
and U3772 (N_3772,N_3533,N_3411);
or U3773 (N_3773,N_3562,N_3407);
or U3774 (N_3774,N_3522,N_3596);
nand U3775 (N_3775,N_3411,N_3477);
nor U3776 (N_3776,N_3467,N_3470);
and U3777 (N_3777,N_3417,N_3510);
and U3778 (N_3778,N_3494,N_3402);
nand U3779 (N_3779,N_3581,N_3519);
and U3780 (N_3780,N_3439,N_3419);
xor U3781 (N_3781,N_3579,N_3488);
and U3782 (N_3782,N_3535,N_3458);
or U3783 (N_3783,N_3588,N_3462);
and U3784 (N_3784,N_3473,N_3586);
and U3785 (N_3785,N_3579,N_3430);
nand U3786 (N_3786,N_3572,N_3545);
or U3787 (N_3787,N_3538,N_3497);
and U3788 (N_3788,N_3459,N_3460);
nor U3789 (N_3789,N_3402,N_3433);
nor U3790 (N_3790,N_3497,N_3533);
xor U3791 (N_3791,N_3568,N_3476);
nor U3792 (N_3792,N_3504,N_3453);
or U3793 (N_3793,N_3462,N_3503);
nor U3794 (N_3794,N_3463,N_3595);
nand U3795 (N_3795,N_3588,N_3597);
and U3796 (N_3796,N_3483,N_3494);
nand U3797 (N_3797,N_3435,N_3402);
and U3798 (N_3798,N_3491,N_3474);
and U3799 (N_3799,N_3419,N_3527);
nand U3800 (N_3800,N_3752,N_3693);
nand U3801 (N_3801,N_3736,N_3765);
nand U3802 (N_3802,N_3708,N_3645);
and U3803 (N_3803,N_3675,N_3643);
nor U3804 (N_3804,N_3767,N_3639);
and U3805 (N_3805,N_3661,N_3760);
nand U3806 (N_3806,N_3705,N_3787);
nand U3807 (N_3807,N_3631,N_3761);
and U3808 (N_3808,N_3759,N_3611);
xor U3809 (N_3809,N_3666,N_3657);
nand U3810 (N_3810,N_3714,N_3637);
or U3811 (N_3811,N_3627,N_3753);
nor U3812 (N_3812,N_3709,N_3758);
nor U3813 (N_3813,N_3775,N_3686);
nand U3814 (N_3814,N_3641,N_3737);
or U3815 (N_3815,N_3707,N_3731);
or U3816 (N_3816,N_3628,N_3704);
nand U3817 (N_3817,N_3679,N_3653);
or U3818 (N_3818,N_3788,N_3642);
nor U3819 (N_3819,N_3744,N_3713);
and U3820 (N_3820,N_3624,N_3687);
nand U3821 (N_3821,N_3689,N_3784);
or U3822 (N_3822,N_3751,N_3727);
nand U3823 (N_3823,N_3778,N_3688);
and U3824 (N_3824,N_3754,N_3663);
nor U3825 (N_3825,N_3667,N_3746);
nor U3826 (N_3826,N_3623,N_3655);
or U3827 (N_3827,N_3699,N_3755);
xor U3828 (N_3828,N_3735,N_3716);
nand U3829 (N_3829,N_3729,N_3664);
or U3830 (N_3830,N_3711,N_3659);
or U3831 (N_3831,N_3660,N_3697);
or U3832 (N_3832,N_3601,N_3681);
nor U3833 (N_3833,N_3656,N_3792);
nand U3834 (N_3834,N_3724,N_3621);
and U3835 (N_3835,N_3715,N_3793);
nor U3836 (N_3836,N_3691,N_3612);
nor U3837 (N_3837,N_3692,N_3644);
nor U3838 (N_3838,N_3682,N_3650);
or U3839 (N_3839,N_3723,N_3622);
and U3840 (N_3840,N_3783,N_3617);
or U3841 (N_3841,N_3694,N_3678);
and U3842 (N_3842,N_3658,N_3618);
xnor U3843 (N_3843,N_3726,N_3683);
and U3844 (N_3844,N_3634,N_3769);
and U3845 (N_3845,N_3721,N_3768);
nand U3846 (N_3846,N_3734,N_3604);
nand U3847 (N_3847,N_3795,N_3670);
xnor U3848 (N_3848,N_3603,N_3668);
nand U3849 (N_3849,N_3698,N_3791);
nor U3850 (N_3850,N_3609,N_3770);
or U3851 (N_3851,N_3733,N_3763);
nor U3852 (N_3852,N_3677,N_3706);
nor U3853 (N_3853,N_3640,N_3756);
and U3854 (N_3854,N_3600,N_3790);
or U3855 (N_3855,N_3798,N_3614);
nor U3856 (N_3856,N_3674,N_3607);
nand U3857 (N_3857,N_3680,N_3685);
nor U3858 (N_3858,N_3749,N_3722);
and U3859 (N_3859,N_3654,N_3613);
nor U3860 (N_3860,N_3796,N_3789);
and U3861 (N_3861,N_3728,N_3771);
xnor U3862 (N_3862,N_3773,N_3700);
nand U3863 (N_3863,N_3635,N_3750);
or U3864 (N_3864,N_3747,N_3636);
nor U3865 (N_3865,N_3647,N_3672);
or U3866 (N_3866,N_3602,N_3738);
and U3867 (N_3867,N_3762,N_3608);
or U3868 (N_3868,N_3730,N_3776);
nand U3869 (N_3869,N_3652,N_3632);
nor U3870 (N_3870,N_3665,N_3777);
and U3871 (N_3871,N_3772,N_3606);
nand U3872 (N_3872,N_3648,N_3732);
and U3873 (N_3873,N_3718,N_3633);
nor U3874 (N_3874,N_3712,N_3702);
nand U3875 (N_3875,N_3799,N_3717);
and U3876 (N_3876,N_3780,N_3649);
and U3877 (N_3877,N_3625,N_3764);
or U3878 (N_3878,N_3748,N_3701);
nor U3879 (N_3879,N_3797,N_3794);
nor U3880 (N_3880,N_3725,N_3651);
and U3881 (N_3881,N_3781,N_3610);
nor U3882 (N_3882,N_3743,N_3719);
and U3883 (N_3883,N_3630,N_3766);
and U3884 (N_3884,N_3615,N_3782);
or U3885 (N_3885,N_3676,N_3745);
or U3886 (N_3886,N_3774,N_3740);
nor U3887 (N_3887,N_3671,N_3662);
xnor U3888 (N_3888,N_3673,N_3605);
nor U3889 (N_3889,N_3669,N_3720);
nand U3890 (N_3890,N_3684,N_3620);
and U3891 (N_3891,N_3741,N_3703);
nand U3892 (N_3892,N_3629,N_3710);
nand U3893 (N_3893,N_3619,N_3690);
nor U3894 (N_3894,N_3695,N_3785);
xor U3895 (N_3895,N_3626,N_3786);
nand U3896 (N_3896,N_3638,N_3616);
nor U3897 (N_3897,N_3739,N_3742);
or U3898 (N_3898,N_3696,N_3779);
nor U3899 (N_3899,N_3646,N_3757);
nor U3900 (N_3900,N_3663,N_3797);
nor U3901 (N_3901,N_3615,N_3605);
or U3902 (N_3902,N_3717,N_3708);
nor U3903 (N_3903,N_3786,N_3708);
nor U3904 (N_3904,N_3603,N_3707);
nor U3905 (N_3905,N_3796,N_3758);
and U3906 (N_3906,N_3773,N_3674);
or U3907 (N_3907,N_3709,N_3708);
or U3908 (N_3908,N_3768,N_3705);
nor U3909 (N_3909,N_3677,N_3734);
and U3910 (N_3910,N_3715,N_3663);
or U3911 (N_3911,N_3786,N_3647);
and U3912 (N_3912,N_3708,N_3775);
xor U3913 (N_3913,N_3788,N_3614);
or U3914 (N_3914,N_3685,N_3616);
and U3915 (N_3915,N_3675,N_3775);
nand U3916 (N_3916,N_3689,N_3688);
and U3917 (N_3917,N_3734,N_3602);
and U3918 (N_3918,N_3602,N_3699);
and U3919 (N_3919,N_3793,N_3683);
nand U3920 (N_3920,N_3698,N_3780);
or U3921 (N_3921,N_3722,N_3710);
nor U3922 (N_3922,N_3729,N_3651);
and U3923 (N_3923,N_3646,N_3782);
nor U3924 (N_3924,N_3781,N_3625);
or U3925 (N_3925,N_3790,N_3691);
nand U3926 (N_3926,N_3662,N_3660);
or U3927 (N_3927,N_3728,N_3672);
nand U3928 (N_3928,N_3721,N_3696);
nand U3929 (N_3929,N_3624,N_3754);
and U3930 (N_3930,N_3764,N_3686);
or U3931 (N_3931,N_3719,N_3658);
and U3932 (N_3932,N_3636,N_3740);
and U3933 (N_3933,N_3644,N_3674);
xnor U3934 (N_3934,N_3642,N_3784);
or U3935 (N_3935,N_3693,N_3621);
nor U3936 (N_3936,N_3765,N_3676);
or U3937 (N_3937,N_3638,N_3693);
nor U3938 (N_3938,N_3786,N_3611);
and U3939 (N_3939,N_3768,N_3671);
nor U3940 (N_3940,N_3711,N_3658);
nor U3941 (N_3941,N_3713,N_3623);
or U3942 (N_3942,N_3675,N_3794);
and U3943 (N_3943,N_3695,N_3784);
xnor U3944 (N_3944,N_3778,N_3788);
and U3945 (N_3945,N_3608,N_3666);
nand U3946 (N_3946,N_3667,N_3749);
or U3947 (N_3947,N_3610,N_3613);
nor U3948 (N_3948,N_3761,N_3619);
and U3949 (N_3949,N_3760,N_3783);
nor U3950 (N_3950,N_3728,N_3701);
nor U3951 (N_3951,N_3707,N_3778);
and U3952 (N_3952,N_3699,N_3702);
nor U3953 (N_3953,N_3798,N_3648);
nor U3954 (N_3954,N_3786,N_3720);
nand U3955 (N_3955,N_3681,N_3650);
nand U3956 (N_3956,N_3786,N_3617);
nor U3957 (N_3957,N_3738,N_3742);
or U3958 (N_3958,N_3628,N_3631);
nor U3959 (N_3959,N_3622,N_3699);
or U3960 (N_3960,N_3684,N_3704);
or U3961 (N_3961,N_3695,N_3715);
and U3962 (N_3962,N_3643,N_3646);
nor U3963 (N_3963,N_3703,N_3635);
or U3964 (N_3964,N_3615,N_3623);
or U3965 (N_3965,N_3789,N_3646);
or U3966 (N_3966,N_3604,N_3658);
and U3967 (N_3967,N_3629,N_3706);
and U3968 (N_3968,N_3691,N_3613);
nor U3969 (N_3969,N_3765,N_3709);
nor U3970 (N_3970,N_3676,N_3619);
and U3971 (N_3971,N_3739,N_3725);
and U3972 (N_3972,N_3684,N_3622);
xnor U3973 (N_3973,N_3645,N_3703);
nand U3974 (N_3974,N_3730,N_3616);
nand U3975 (N_3975,N_3694,N_3628);
and U3976 (N_3976,N_3701,N_3660);
nand U3977 (N_3977,N_3760,N_3767);
nor U3978 (N_3978,N_3648,N_3716);
nand U3979 (N_3979,N_3618,N_3771);
and U3980 (N_3980,N_3763,N_3645);
nor U3981 (N_3981,N_3755,N_3703);
or U3982 (N_3982,N_3737,N_3682);
or U3983 (N_3983,N_3621,N_3751);
nor U3984 (N_3984,N_3714,N_3724);
nor U3985 (N_3985,N_3653,N_3736);
or U3986 (N_3986,N_3710,N_3791);
nor U3987 (N_3987,N_3672,N_3692);
and U3988 (N_3988,N_3600,N_3784);
and U3989 (N_3989,N_3653,N_3624);
xnor U3990 (N_3990,N_3672,N_3673);
and U3991 (N_3991,N_3788,N_3693);
nand U3992 (N_3992,N_3715,N_3686);
nand U3993 (N_3993,N_3740,N_3729);
nand U3994 (N_3994,N_3613,N_3735);
or U3995 (N_3995,N_3704,N_3798);
nand U3996 (N_3996,N_3796,N_3617);
nor U3997 (N_3997,N_3662,N_3708);
or U3998 (N_3998,N_3771,N_3733);
and U3999 (N_3999,N_3603,N_3643);
nor U4000 (N_4000,N_3838,N_3913);
nand U4001 (N_4001,N_3906,N_3802);
or U4002 (N_4002,N_3849,N_3821);
nor U4003 (N_4003,N_3826,N_3901);
nand U4004 (N_4004,N_3841,N_3839);
or U4005 (N_4005,N_3954,N_3816);
nand U4006 (N_4006,N_3822,N_3819);
nor U4007 (N_4007,N_3918,N_3877);
or U4008 (N_4008,N_3870,N_3805);
xnor U4009 (N_4009,N_3938,N_3878);
nand U4010 (N_4010,N_3987,N_3960);
nor U4011 (N_4011,N_3966,N_3976);
nor U4012 (N_4012,N_3833,N_3945);
nor U4013 (N_4013,N_3894,N_3897);
nand U4014 (N_4014,N_3803,N_3977);
or U4015 (N_4015,N_3852,N_3932);
or U4016 (N_4016,N_3971,N_3853);
nand U4017 (N_4017,N_3956,N_3818);
and U4018 (N_4018,N_3921,N_3832);
nor U4019 (N_4019,N_3836,N_3957);
nand U4020 (N_4020,N_3813,N_3898);
nand U4021 (N_4021,N_3824,N_3997);
or U4022 (N_4022,N_3861,N_3990);
and U4023 (N_4023,N_3896,N_3888);
nor U4024 (N_4024,N_3926,N_3893);
or U4025 (N_4025,N_3863,N_3804);
nand U4026 (N_4026,N_3817,N_3912);
nand U4027 (N_4027,N_3992,N_3975);
nor U4028 (N_4028,N_3860,N_3844);
nand U4029 (N_4029,N_3916,N_3949);
or U4030 (N_4030,N_3820,N_3842);
and U4031 (N_4031,N_3808,N_3940);
nand U4032 (N_4032,N_3985,N_3895);
nor U4033 (N_4033,N_3983,N_3953);
nand U4034 (N_4034,N_3995,N_3904);
and U4035 (N_4035,N_3930,N_3947);
nand U4036 (N_4036,N_3955,N_3815);
or U4037 (N_4037,N_3936,N_3811);
nor U4038 (N_4038,N_3825,N_3968);
nand U4039 (N_4039,N_3931,N_3923);
or U4040 (N_4040,N_3874,N_3996);
or U4041 (N_4041,N_3941,N_3812);
and U4042 (N_4042,N_3963,N_3988);
nor U4043 (N_4043,N_3946,N_3908);
and U4044 (N_4044,N_3974,N_3984);
nor U4045 (N_4045,N_3848,N_3880);
nor U4046 (N_4046,N_3886,N_3973);
nor U4047 (N_4047,N_3882,N_3967);
nor U4048 (N_4048,N_3951,N_3847);
nand U4049 (N_4049,N_3905,N_3806);
nand U4050 (N_4050,N_3810,N_3843);
nor U4051 (N_4051,N_3881,N_3837);
nor U4052 (N_4052,N_3937,N_3922);
or U4053 (N_4053,N_3943,N_3828);
nor U4054 (N_4054,N_3899,N_3876);
or U4055 (N_4055,N_3911,N_3920);
and U4056 (N_4056,N_3980,N_3855);
and U4057 (N_4057,N_3934,N_3840);
and U4058 (N_4058,N_3857,N_3950);
nor U4059 (N_4059,N_3903,N_3944);
nand U4060 (N_4060,N_3919,N_3884);
nor U4061 (N_4061,N_3887,N_3994);
or U4062 (N_4062,N_3890,N_3807);
nor U4063 (N_4063,N_3989,N_3969);
and U4064 (N_4064,N_3865,N_3965);
or U4065 (N_4065,N_3979,N_3892);
and U4066 (N_4066,N_3850,N_3928);
and U4067 (N_4067,N_3959,N_3869);
nor U4068 (N_4068,N_3972,N_3889);
nor U4069 (N_4069,N_3962,N_3879);
and U4070 (N_4070,N_3872,N_3866);
nor U4071 (N_4071,N_3999,N_3800);
nand U4072 (N_4072,N_3900,N_3809);
and U4073 (N_4073,N_3891,N_3902);
and U4074 (N_4074,N_3925,N_3873);
nor U4075 (N_4075,N_3875,N_3981);
or U4076 (N_4076,N_3862,N_3935);
nor U4077 (N_4077,N_3914,N_3907);
nor U4078 (N_4078,N_3831,N_3856);
nor U4079 (N_4079,N_3835,N_3834);
nor U4080 (N_4080,N_3964,N_3885);
or U4081 (N_4081,N_3970,N_3929);
nor U4082 (N_4082,N_3958,N_3909);
nand U4083 (N_4083,N_3993,N_3851);
or U4084 (N_4084,N_3915,N_3854);
nand U4085 (N_4085,N_3846,N_3883);
or U4086 (N_4086,N_3991,N_3910);
nor U4087 (N_4087,N_3978,N_3927);
and U4088 (N_4088,N_3952,N_3871);
or U4089 (N_4089,N_3868,N_3942);
or U4090 (N_4090,N_3823,N_3917);
nor U4091 (N_4091,N_3924,N_3933);
or U4092 (N_4092,N_3864,N_3859);
nand U4093 (N_4093,N_3961,N_3829);
and U4094 (N_4094,N_3986,N_3867);
nand U4095 (N_4095,N_3827,N_3830);
nor U4096 (N_4096,N_3982,N_3845);
or U4097 (N_4097,N_3858,N_3814);
nand U4098 (N_4098,N_3948,N_3939);
and U4099 (N_4099,N_3998,N_3801);
and U4100 (N_4100,N_3880,N_3999);
and U4101 (N_4101,N_3815,N_3844);
or U4102 (N_4102,N_3915,N_3926);
nand U4103 (N_4103,N_3892,N_3883);
nor U4104 (N_4104,N_3860,N_3811);
nand U4105 (N_4105,N_3851,N_3957);
or U4106 (N_4106,N_3958,N_3864);
nand U4107 (N_4107,N_3970,N_3979);
and U4108 (N_4108,N_3932,N_3918);
and U4109 (N_4109,N_3854,N_3952);
or U4110 (N_4110,N_3906,N_3949);
nor U4111 (N_4111,N_3866,N_3929);
nor U4112 (N_4112,N_3804,N_3824);
nor U4113 (N_4113,N_3931,N_3866);
and U4114 (N_4114,N_3963,N_3836);
nand U4115 (N_4115,N_3914,N_3801);
and U4116 (N_4116,N_3891,N_3890);
and U4117 (N_4117,N_3829,N_3991);
nor U4118 (N_4118,N_3880,N_3801);
nor U4119 (N_4119,N_3958,N_3903);
and U4120 (N_4120,N_3868,N_3932);
or U4121 (N_4121,N_3974,N_3844);
nand U4122 (N_4122,N_3835,N_3978);
and U4123 (N_4123,N_3817,N_3987);
nand U4124 (N_4124,N_3873,N_3874);
nand U4125 (N_4125,N_3831,N_3987);
or U4126 (N_4126,N_3881,N_3989);
and U4127 (N_4127,N_3913,N_3835);
nor U4128 (N_4128,N_3896,N_3913);
nand U4129 (N_4129,N_3998,N_3991);
or U4130 (N_4130,N_3826,N_3870);
and U4131 (N_4131,N_3973,N_3863);
nand U4132 (N_4132,N_3870,N_3836);
or U4133 (N_4133,N_3816,N_3998);
nand U4134 (N_4134,N_3884,N_3943);
xor U4135 (N_4135,N_3890,N_3941);
or U4136 (N_4136,N_3907,N_3850);
or U4137 (N_4137,N_3877,N_3883);
nand U4138 (N_4138,N_3959,N_3802);
or U4139 (N_4139,N_3843,N_3958);
and U4140 (N_4140,N_3827,N_3900);
and U4141 (N_4141,N_3991,N_3952);
or U4142 (N_4142,N_3998,N_3805);
or U4143 (N_4143,N_3891,N_3811);
or U4144 (N_4144,N_3800,N_3876);
or U4145 (N_4145,N_3867,N_3895);
or U4146 (N_4146,N_3942,N_3864);
and U4147 (N_4147,N_3946,N_3812);
or U4148 (N_4148,N_3865,N_3860);
nand U4149 (N_4149,N_3947,N_3985);
nor U4150 (N_4150,N_3885,N_3921);
nor U4151 (N_4151,N_3903,N_3860);
and U4152 (N_4152,N_3885,N_3961);
nand U4153 (N_4153,N_3987,N_3833);
or U4154 (N_4154,N_3949,N_3909);
xor U4155 (N_4155,N_3907,N_3978);
or U4156 (N_4156,N_3865,N_3985);
and U4157 (N_4157,N_3939,N_3936);
xor U4158 (N_4158,N_3998,N_3919);
or U4159 (N_4159,N_3944,N_3909);
nor U4160 (N_4160,N_3926,N_3993);
or U4161 (N_4161,N_3858,N_3849);
nor U4162 (N_4162,N_3915,N_3920);
or U4163 (N_4163,N_3967,N_3893);
nand U4164 (N_4164,N_3942,N_3865);
and U4165 (N_4165,N_3916,N_3886);
nand U4166 (N_4166,N_3929,N_3864);
and U4167 (N_4167,N_3938,N_3910);
and U4168 (N_4168,N_3925,N_3829);
nor U4169 (N_4169,N_3826,N_3897);
nor U4170 (N_4170,N_3883,N_3920);
and U4171 (N_4171,N_3878,N_3854);
xor U4172 (N_4172,N_3958,N_3815);
nor U4173 (N_4173,N_3971,N_3932);
nor U4174 (N_4174,N_3932,N_3892);
nand U4175 (N_4175,N_3925,N_3825);
or U4176 (N_4176,N_3843,N_3919);
or U4177 (N_4177,N_3910,N_3886);
nand U4178 (N_4178,N_3967,N_3829);
nand U4179 (N_4179,N_3979,N_3932);
or U4180 (N_4180,N_3888,N_3950);
nand U4181 (N_4181,N_3886,N_3941);
and U4182 (N_4182,N_3933,N_3961);
nor U4183 (N_4183,N_3999,N_3973);
and U4184 (N_4184,N_3833,N_3888);
and U4185 (N_4185,N_3833,N_3981);
nor U4186 (N_4186,N_3820,N_3962);
nor U4187 (N_4187,N_3883,N_3918);
nor U4188 (N_4188,N_3951,N_3817);
xnor U4189 (N_4189,N_3976,N_3936);
and U4190 (N_4190,N_3920,N_3912);
or U4191 (N_4191,N_3916,N_3858);
or U4192 (N_4192,N_3991,N_3932);
or U4193 (N_4193,N_3850,N_3920);
and U4194 (N_4194,N_3823,N_3919);
nand U4195 (N_4195,N_3963,N_3815);
or U4196 (N_4196,N_3955,N_3902);
xnor U4197 (N_4197,N_3853,N_3802);
or U4198 (N_4198,N_3906,N_3944);
and U4199 (N_4199,N_3940,N_3886);
nor U4200 (N_4200,N_4057,N_4055);
nand U4201 (N_4201,N_4090,N_4169);
and U4202 (N_4202,N_4024,N_4063);
nor U4203 (N_4203,N_4074,N_4139);
and U4204 (N_4204,N_4165,N_4029);
and U4205 (N_4205,N_4031,N_4132);
nor U4206 (N_4206,N_4120,N_4018);
nor U4207 (N_4207,N_4160,N_4097);
nand U4208 (N_4208,N_4008,N_4065);
nand U4209 (N_4209,N_4193,N_4014);
and U4210 (N_4210,N_4012,N_4115);
or U4211 (N_4211,N_4149,N_4025);
xor U4212 (N_4212,N_4136,N_4013);
or U4213 (N_4213,N_4107,N_4032);
and U4214 (N_4214,N_4003,N_4137);
and U4215 (N_4215,N_4061,N_4166);
and U4216 (N_4216,N_4021,N_4094);
and U4217 (N_4217,N_4062,N_4056);
and U4218 (N_4218,N_4000,N_4142);
nor U4219 (N_4219,N_4030,N_4157);
nand U4220 (N_4220,N_4146,N_4156);
nor U4221 (N_4221,N_4124,N_4079);
nor U4222 (N_4222,N_4150,N_4050);
and U4223 (N_4223,N_4005,N_4070);
and U4224 (N_4224,N_4179,N_4052);
nor U4225 (N_4225,N_4147,N_4022);
nand U4226 (N_4226,N_4197,N_4167);
and U4227 (N_4227,N_4064,N_4006);
nand U4228 (N_4228,N_4010,N_4119);
xor U4229 (N_4229,N_4118,N_4084);
or U4230 (N_4230,N_4026,N_4134);
nor U4231 (N_4231,N_4016,N_4145);
and U4232 (N_4232,N_4130,N_4140);
and U4233 (N_4233,N_4187,N_4182);
and U4234 (N_4234,N_4034,N_4069);
or U4235 (N_4235,N_4045,N_4004);
nand U4236 (N_4236,N_4100,N_4059);
nor U4237 (N_4237,N_4183,N_4190);
or U4238 (N_4238,N_4162,N_4102);
nor U4239 (N_4239,N_4049,N_4173);
nand U4240 (N_4240,N_4088,N_4087);
and U4241 (N_4241,N_4178,N_4048);
nand U4242 (N_4242,N_4066,N_4168);
or U4243 (N_4243,N_4114,N_4108);
nor U4244 (N_4244,N_4199,N_4128);
nor U4245 (N_4245,N_4105,N_4125);
or U4246 (N_4246,N_4185,N_4138);
nor U4247 (N_4247,N_4051,N_4086);
or U4248 (N_4248,N_4080,N_4117);
nor U4249 (N_4249,N_4163,N_4184);
nand U4250 (N_4250,N_4076,N_4151);
or U4251 (N_4251,N_4158,N_4180);
and U4252 (N_4252,N_4152,N_4009);
nor U4253 (N_4253,N_4047,N_4072);
nand U4254 (N_4254,N_4054,N_4155);
and U4255 (N_4255,N_4122,N_4077);
or U4256 (N_4256,N_4020,N_4001);
nand U4257 (N_4257,N_4035,N_4126);
or U4258 (N_4258,N_4133,N_4083);
or U4259 (N_4259,N_4042,N_4177);
nand U4260 (N_4260,N_4104,N_4186);
and U4261 (N_4261,N_4046,N_4044);
nand U4262 (N_4262,N_4110,N_4191);
nand U4263 (N_4263,N_4198,N_4192);
and U4264 (N_4264,N_4175,N_4141);
and U4265 (N_4265,N_4172,N_4002);
nand U4266 (N_4266,N_4127,N_4116);
and U4267 (N_4267,N_4109,N_4040);
nand U4268 (N_4268,N_4196,N_4073);
or U4269 (N_4269,N_4131,N_4148);
xor U4270 (N_4270,N_4041,N_4161);
and U4271 (N_4271,N_4098,N_4113);
nand U4272 (N_4272,N_4007,N_4171);
nand U4273 (N_4273,N_4015,N_4036);
nand U4274 (N_4274,N_4053,N_4060);
nand U4275 (N_4275,N_4101,N_4092);
and U4276 (N_4276,N_4170,N_4176);
nor U4277 (N_4277,N_4058,N_4017);
nor U4278 (N_4278,N_4071,N_4089);
and U4279 (N_4279,N_4091,N_4123);
nor U4280 (N_4280,N_4037,N_4081);
nor U4281 (N_4281,N_4135,N_4144);
or U4282 (N_4282,N_4189,N_4011);
nand U4283 (N_4283,N_4096,N_4111);
nor U4284 (N_4284,N_4174,N_4078);
and U4285 (N_4285,N_4027,N_4085);
or U4286 (N_4286,N_4159,N_4075);
nor U4287 (N_4287,N_4067,N_4068);
or U4288 (N_4288,N_4112,N_4164);
nand U4289 (N_4289,N_4195,N_4103);
nor U4290 (N_4290,N_4033,N_4039);
or U4291 (N_4291,N_4181,N_4095);
nor U4292 (N_4292,N_4099,N_4023);
and U4293 (N_4293,N_4082,N_4106);
or U4294 (N_4294,N_4019,N_4043);
and U4295 (N_4295,N_4153,N_4188);
nand U4296 (N_4296,N_4028,N_4038);
nor U4297 (N_4297,N_4093,N_4121);
or U4298 (N_4298,N_4143,N_4154);
and U4299 (N_4299,N_4129,N_4194);
and U4300 (N_4300,N_4055,N_4026);
nor U4301 (N_4301,N_4133,N_4164);
nand U4302 (N_4302,N_4084,N_4069);
nor U4303 (N_4303,N_4074,N_4014);
or U4304 (N_4304,N_4152,N_4138);
nor U4305 (N_4305,N_4056,N_4072);
nand U4306 (N_4306,N_4052,N_4026);
xnor U4307 (N_4307,N_4093,N_4111);
and U4308 (N_4308,N_4061,N_4143);
nor U4309 (N_4309,N_4014,N_4026);
and U4310 (N_4310,N_4199,N_4150);
xnor U4311 (N_4311,N_4108,N_4002);
nor U4312 (N_4312,N_4190,N_4099);
and U4313 (N_4313,N_4194,N_4157);
and U4314 (N_4314,N_4149,N_4163);
or U4315 (N_4315,N_4063,N_4140);
nor U4316 (N_4316,N_4059,N_4013);
and U4317 (N_4317,N_4149,N_4076);
and U4318 (N_4318,N_4147,N_4144);
nand U4319 (N_4319,N_4147,N_4066);
and U4320 (N_4320,N_4083,N_4137);
and U4321 (N_4321,N_4168,N_4074);
or U4322 (N_4322,N_4120,N_4164);
xnor U4323 (N_4323,N_4111,N_4143);
nand U4324 (N_4324,N_4007,N_4189);
nand U4325 (N_4325,N_4090,N_4089);
and U4326 (N_4326,N_4151,N_4101);
nand U4327 (N_4327,N_4199,N_4012);
nor U4328 (N_4328,N_4171,N_4087);
and U4329 (N_4329,N_4099,N_4154);
or U4330 (N_4330,N_4114,N_4087);
and U4331 (N_4331,N_4176,N_4070);
and U4332 (N_4332,N_4078,N_4086);
nor U4333 (N_4333,N_4058,N_4168);
or U4334 (N_4334,N_4196,N_4083);
and U4335 (N_4335,N_4167,N_4176);
nor U4336 (N_4336,N_4109,N_4019);
nand U4337 (N_4337,N_4141,N_4005);
nand U4338 (N_4338,N_4003,N_4060);
nand U4339 (N_4339,N_4031,N_4090);
and U4340 (N_4340,N_4166,N_4080);
nand U4341 (N_4341,N_4039,N_4021);
nor U4342 (N_4342,N_4184,N_4069);
and U4343 (N_4343,N_4039,N_4149);
and U4344 (N_4344,N_4077,N_4013);
nor U4345 (N_4345,N_4179,N_4092);
nor U4346 (N_4346,N_4129,N_4063);
nor U4347 (N_4347,N_4009,N_4093);
or U4348 (N_4348,N_4118,N_4054);
and U4349 (N_4349,N_4068,N_4159);
or U4350 (N_4350,N_4075,N_4097);
nand U4351 (N_4351,N_4013,N_4049);
or U4352 (N_4352,N_4102,N_4095);
nor U4353 (N_4353,N_4125,N_4109);
nor U4354 (N_4354,N_4116,N_4106);
and U4355 (N_4355,N_4054,N_4154);
nand U4356 (N_4356,N_4168,N_4072);
nor U4357 (N_4357,N_4025,N_4167);
nor U4358 (N_4358,N_4176,N_4002);
or U4359 (N_4359,N_4053,N_4187);
or U4360 (N_4360,N_4026,N_4151);
nand U4361 (N_4361,N_4169,N_4074);
and U4362 (N_4362,N_4117,N_4169);
nor U4363 (N_4363,N_4061,N_4033);
xor U4364 (N_4364,N_4052,N_4084);
nand U4365 (N_4365,N_4018,N_4055);
nor U4366 (N_4366,N_4045,N_4195);
or U4367 (N_4367,N_4120,N_4065);
xnor U4368 (N_4368,N_4065,N_4045);
nand U4369 (N_4369,N_4177,N_4128);
or U4370 (N_4370,N_4186,N_4012);
nor U4371 (N_4371,N_4095,N_4176);
or U4372 (N_4372,N_4153,N_4117);
nor U4373 (N_4373,N_4053,N_4109);
nor U4374 (N_4374,N_4059,N_4118);
nor U4375 (N_4375,N_4062,N_4198);
and U4376 (N_4376,N_4157,N_4145);
and U4377 (N_4377,N_4004,N_4110);
and U4378 (N_4378,N_4101,N_4163);
nand U4379 (N_4379,N_4176,N_4094);
and U4380 (N_4380,N_4010,N_4080);
nand U4381 (N_4381,N_4166,N_4046);
or U4382 (N_4382,N_4105,N_4082);
nor U4383 (N_4383,N_4018,N_4136);
xor U4384 (N_4384,N_4102,N_4049);
nand U4385 (N_4385,N_4099,N_4053);
nor U4386 (N_4386,N_4147,N_4050);
nand U4387 (N_4387,N_4040,N_4138);
nor U4388 (N_4388,N_4041,N_4010);
and U4389 (N_4389,N_4136,N_4176);
and U4390 (N_4390,N_4140,N_4036);
and U4391 (N_4391,N_4037,N_4095);
or U4392 (N_4392,N_4135,N_4165);
and U4393 (N_4393,N_4118,N_4016);
and U4394 (N_4394,N_4098,N_4144);
nor U4395 (N_4395,N_4093,N_4038);
or U4396 (N_4396,N_4106,N_4099);
xnor U4397 (N_4397,N_4095,N_4060);
nand U4398 (N_4398,N_4050,N_4175);
or U4399 (N_4399,N_4016,N_4155);
nand U4400 (N_4400,N_4368,N_4287);
or U4401 (N_4401,N_4240,N_4291);
nand U4402 (N_4402,N_4367,N_4289);
or U4403 (N_4403,N_4327,N_4261);
nor U4404 (N_4404,N_4230,N_4345);
nor U4405 (N_4405,N_4271,N_4294);
nor U4406 (N_4406,N_4236,N_4337);
and U4407 (N_4407,N_4341,N_4312);
or U4408 (N_4408,N_4251,N_4342);
xor U4409 (N_4409,N_4349,N_4295);
nand U4410 (N_4410,N_4210,N_4383);
nand U4411 (N_4411,N_4226,N_4296);
nand U4412 (N_4412,N_4386,N_4375);
nor U4413 (N_4413,N_4288,N_4263);
or U4414 (N_4414,N_4292,N_4250);
nor U4415 (N_4415,N_4352,N_4222);
and U4416 (N_4416,N_4326,N_4385);
and U4417 (N_4417,N_4313,N_4238);
nor U4418 (N_4418,N_4237,N_4213);
and U4419 (N_4419,N_4235,N_4234);
nand U4420 (N_4420,N_4365,N_4243);
and U4421 (N_4421,N_4246,N_4320);
nor U4422 (N_4422,N_4297,N_4394);
or U4423 (N_4423,N_4266,N_4353);
or U4424 (N_4424,N_4225,N_4204);
nand U4425 (N_4425,N_4208,N_4391);
xnor U4426 (N_4426,N_4274,N_4216);
nand U4427 (N_4427,N_4220,N_4227);
or U4428 (N_4428,N_4293,N_4347);
nor U4429 (N_4429,N_4203,N_4336);
nor U4430 (N_4430,N_4300,N_4343);
nand U4431 (N_4431,N_4374,N_4275);
and U4432 (N_4432,N_4315,N_4371);
or U4433 (N_4433,N_4209,N_4378);
or U4434 (N_4434,N_4355,N_4282);
and U4435 (N_4435,N_4369,N_4285);
nor U4436 (N_4436,N_4307,N_4387);
or U4437 (N_4437,N_4223,N_4322);
or U4438 (N_4438,N_4211,N_4305);
or U4439 (N_4439,N_4325,N_4397);
nand U4440 (N_4440,N_4260,N_4389);
or U4441 (N_4441,N_4268,N_4248);
nand U4442 (N_4442,N_4231,N_4351);
nand U4443 (N_4443,N_4366,N_4219);
and U4444 (N_4444,N_4280,N_4247);
nor U4445 (N_4445,N_4255,N_4284);
nand U4446 (N_4446,N_4205,N_4270);
nand U4447 (N_4447,N_4232,N_4324);
and U4448 (N_4448,N_4399,N_4370);
or U4449 (N_4449,N_4241,N_4304);
nor U4450 (N_4450,N_4393,N_4354);
and U4451 (N_4451,N_4317,N_4311);
or U4452 (N_4452,N_4332,N_4356);
or U4453 (N_4453,N_4276,N_4376);
and U4454 (N_4454,N_4279,N_4265);
nor U4455 (N_4455,N_4388,N_4373);
and U4456 (N_4456,N_4212,N_4381);
nor U4457 (N_4457,N_4302,N_4318);
nand U4458 (N_4458,N_4273,N_4364);
nor U4459 (N_4459,N_4286,N_4264);
nor U4460 (N_4460,N_4283,N_4392);
or U4461 (N_4461,N_4301,N_4314);
and U4462 (N_4462,N_4206,N_4290);
and U4463 (N_4463,N_4339,N_4363);
and U4464 (N_4464,N_4396,N_4239);
nand U4465 (N_4465,N_4306,N_4310);
nor U4466 (N_4466,N_4308,N_4244);
nand U4467 (N_4467,N_4303,N_4278);
or U4468 (N_4468,N_4233,N_4331);
and U4469 (N_4469,N_4333,N_4281);
and U4470 (N_4470,N_4358,N_4330);
nand U4471 (N_4471,N_4357,N_4316);
or U4472 (N_4472,N_4379,N_4207);
and U4473 (N_4473,N_4362,N_4253);
or U4474 (N_4474,N_4321,N_4344);
xnor U4475 (N_4475,N_4249,N_4361);
or U4476 (N_4476,N_4346,N_4340);
nand U4477 (N_4477,N_4384,N_4348);
nor U4478 (N_4478,N_4360,N_4262);
nand U4479 (N_4479,N_4272,N_4328);
nor U4480 (N_4480,N_4221,N_4269);
or U4481 (N_4481,N_4259,N_4377);
nor U4482 (N_4482,N_4229,N_4202);
and U4483 (N_4483,N_4299,N_4201);
or U4484 (N_4484,N_4277,N_4382);
and U4485 (N_4485,N_4214,N_4256);
nor U4486 (N_4486,N_4217,N_4224);
nor U4487 (N_4487,N_4372,N_4242);
or U4488 (N_4488,N_4390,N_4200);
and U4489 (N_4489,N_4338,N_4380);
nand U4490 (N_4490,N_4395,N_4335);
and U4491 (N_4491,N_4252,N_4309);
nor U4492 (N_4492,N_4254,N_4329);
and U4493 (N_4493,N_4298,N_4228);
and U4494 (N_4494,N_4359,N_4257);
or U4495 (N_4495,N_4350,N_4245);
nand U4496 (N_4496,N_4267,N_4398);
nor U4497 (N_4497,N_4258,N_4323);
nand U4498 (N_4498,N_4319,N_4334);
and U4499 (N_4499,N_4218,N_4215);
nand U4500 (N_4500,N_4350,N_4311);
nor U4501 (N_4501,N_4236,N_4212);
nand U4502 (N_4502,N_4209,N_4362);
xor U4503 (N_4503,N_4213,N_4377);
nor U4504 (N_4504,N_4266,N_4290);
nand U4505 (N_4505,N_4364,N_4288);
and U4506 (N_4506,N_4255,N_4238);
or U4507 (N_4507,N_4320,N_4373);
and U4508 (N_4508,N_4327,N_4394);
and U4509 (N_4509,N_4290,N_4239);
and U4510 (N_4510,N_4342,N_4218);
and U4511 (N_4511,N_4228,N_4376);
or U4512 (N_4512,N_4223,N_4235);
nor U4513 (N_4513,N_4339,N_4206);
nor U4514 (N_4514,N_4370,N_4317);
nand U4515 (N_4515,N_4258,N_4324);
or U4516 (N_4516,N_4308,N_4366);
xor U4517 (N_4517,N_4280,N_4294);
and U4518 (N_4518,N_4329,N_4349);
nor U4519 (N_4519,N_4294,N_4230);
nor U4520 (N_4520,N_4213,N_4229);
nor U4521 (N_4521,N_4356,N_4328);
nand U4522 (N_4522,N_4271,N_4239);
nand U4523 (N_4523,N_4246,N_4233);
nand U4524 (N_4524,N_4399,N_4284);
nand U4525 (N_4525,N_4247,N_4308);
and U4526 (N_4526,N_4345,N_4255);
nand U4527 (N_4527,N_4341,N_4234);
nand U4528 (N_4528,N_4256,N_4384);
or U4529 (N_4529,N_4269,N_4320);
xnor U4530 (N_4530,N_4320,N_4236);
and U4531 (N_4531,N_4307,N_4330);
or U4532 (N_4532,N_4283,N_4310);
or U4533 (N_4533,N_4351,N_4289);
and U4534 (N_4534,N_4207,N_4319);
and U4535 (N_4535,N_4365,N_4319);
and U4536 (N_4536,N_4303,N_4378);
or U4537 (N_4537,N_4263,N_4220);
xnor U4538 (N_4538,N_4205,N_4268);
nor U4539 (N_4539,N_4247,N_4354);
and U4540 (N_4540,N_4230,N_4335);
nand U4541 (N_4541,N_4210,N_4351);
or U4542 (N_4542,N_4316,N_4364);
or U4543 (N_4543,N_4266,N_4359);
nor U4544 (N_4544,N_4288,N_4277);
or U4545 (N_4545,N_4206,N_4314);
nand U4546 (N_4546,N_4336,N_4326);
or U4547 (N_4547,N_4273,N_4256);
nand U4548 (N_4548,N_4343,N_4341);
nand U4549 (N_4549,N_4372,N_4385);
and U4550 (N_4550,N_4269,N_4266);
nor U4551 (N_4551,N_4342,N_4376);
nand U4552 (N_4552,N_4390,N_4370);
or U4553 (N_4553,N_4390,N_4217);
nor U4554 (N_4554,N_4285,N_4378);
and U4555 (N_4555,N_4295,N_4291);
nand U4556 (N_4556,N_4383,N_4236);
nor U4557 (N_4557,N_4247,N_4303);
nand U4558 (N_4558,N_4356,N_4209);
nand U4559 (N_4559,N_4250,N_4312);
nand U4560 (N_4560,N_4354,N_4234);
or U4561 (N_4561,N_4314,N_4339);
nand U4562 (N_4562,N_4220,N_4334);
or U4563 (N_4563,N_4281,N_4325);
and U4564 (N_4564,N_4306,N_4241);
or U4565 (N_4565,N_4343,N_4269);
nand U4566 (N_4566,N_4259,N_4224);
nand U4567 (N_4567,N_4315,N_4391);
or U4568 (N_4568,N_4221,N_4233);
and U4569 (N_4569,N_4265,N_4229);
or U4570 (N_4570,N_4218,N_4312);
xnor U4571 (N_4571,N_4304,N_4269);
nand U4572 (N_4572,N_4366,N_4212);
nor U4573 (N_4573,N_4236,N_4395);
and U4574 (N_4574,N_4293,N_4336);
or U4575 (N_4575,N_4242,N_4204);
and U4576 (N_4576,N_4232,N_4209);
and U4577 (N_4577,N_4206,N_4331);
nor U4578 (N_4578,N_4307,N_4239);
or U4579 (N_4579,N_4298,N_4290);
nand U4580 (N_4580,N_4373,N_4286);
and U4581 (N_4581,N_4381,N_4303);
nand U4582 (N_4582,N_4349,N_4385);
or U4583 (N_4583,N_4336,N_4383);
nor U4584 (N_4584,N_4265,N_4338);
nor U4585 (N_4585,N_4293,N_4348);
nand U4586 (N_4586,N_4249,N_4359);
and U4587 (N_4587,N_4243,N_4291);
xnor U4588 (N_4588,N_4331,N_4320);
and U4589 (N_4589,N_4387,N_4224);
and U4590 (N_4590,N_4344,N_4295);
nand U4591 (N_4591,N_4273,N_4308);
or U4592 (N_4592,N_4258,N_4364);
nor U4593 (N_4593,N_4236,N_4211);
nor U4594 (N_4594,N_4349,N_4341);
nand U4595 (N_4595,N_4215,N_4361);
nor U4596 (N_4596,N_4360,N_4392);
nor U4597 (N_4597,N_4318,N_4317);
nand U4598 (N_4598,N_4385,N_4222);
nor U4599 (N_4599,N_4381,N_4279);
and U4600 (N_4600,N_4465,N_4459);
nand U4601 (N_4601,N_4422,N_4510);
nand U4602 (N_4602,N_4434,N_4575);
nand U4603 (N_4603,N_4527,N_4586);
nor U4604 (N_4604,N_4568,N_4463);
or U4605 (N_4605,N_4512,N_4594);
nor U4606 (N_4606,N_4438,N_4497);
nand U4607 (N_4607,N_4478,N_4521);
nand U4608 (N_4608,N_4415,N_4508);
nor U4609 (N_4609,N_4519,N_4440);
and U4610 (N_4610,N_4414,N_4444);
nor U4611 (N_4611,N_4416,N_4591);
or U4612 (N_4612,N_4419,N_4539);
nor U4613 (N_4613,N_4493,N_4513);
or U4614 (N_4614,N_4489,N_4569);
or U4615 (N_4615,N_4554,N_4450);
nor U4616 (N_4616,N_4476,N_4542);
nor U4617 (N_4617,N_4411,N_4580);
nor U4618 (N_4618,N_4517,N_4445);
and U4619 (N_4619,N_4564,N_4533);
nor U4620 (N_4620,N_4552,N_4409);
nor U4621 (N_4621,N_4545,N_4437);
nand U4622 (N_4622,N_4590,N_4559);
nand U4623 (N_4623,N_4461,N_4469);
and U4624 (N_4624,N_4441,N_4403);
and U4625 (N_4625,N_4543,N_4511);
xor U4626 (N_4626,N_4496,N_4515);
xor U4627 (N_4627,N_4417,N_4425);
and U4628 (N_4628,N_4506,N_4435);
xor U4629 (N_4629,N_4494,N_4582);
or U4630 (N_4630,N_4531,N_4420);
nor U4631 (N_4631,N_4534,N_4439);
or U4632 (N_4632,N_4442,N_4426);
nor U4633 (N_4633,N_4555,N_4436);
nand U4634 (N_4634,N_4412,N_4585);
nor U4635 (N_4635,N_4593,N_4401);
or U4636 (N_4636,N_4509,N_4479);
nand U4637 (N_4637,N_4576,N_4577);
or U4638 (N_4638,N_4405,N_4486);
nor U4639 (N_4639,N_4562,N_4400);
and U4640 (N_4640,N_4561,N_4464);
and U4641 (N_4641,N_4455,N_4536);
or U4642 (N_4642,N_4483,N_4413);
nand U4643 (N_4643,N_4528,N_4589);
xor U4644 (N_4644,N_4452,N_4443);
nand U4645 (N_4645,N_4516,N_4520);
nor U4646 (N_4646,N_4578,N_4421);
nand U4647 (N_4647,N_4556,N_4427);
nand U4648 (N_4648,N_4495,N_4466);
or U4649 (N_4649,N_4524,N_4433);
xor U4650 (N_4650,N_4423,N_4451);
or U4651 (N_4651,N_4473,N_4565);
and U4652 (N_4652,N_4581,N_4540);
or U4653 (N_4653,N_4404,N_4484);
nor U4654 (N_4654,N_4501,N_4503);
nor U4655 (N_4655,N_4407,N_4453);
and U4656 (N_4656,N_4448,N_4522);
or U4657 (N_4657,N_4566,N_4523);
nand U4658 (N_4658,N_4418,N_4446);
xnor U4659 (N_4659,N_4474,N_4579);
or U4660 (N_4660,N_4507,N_4447);
and U4661 (N_4661,N_4549,N_4526);
nand U4662 (N_4662,N_4588,N_4487);
and U4663 (N_4663,N_4541,N_4550);
and U4664 (N_4664,N_4424,N_4505);
nand U4665 (N_4665,N_4557,N_4514);
and U4666 (N_4666,N_4567,N_4525);
nor U4667 (N_4667,N_4597,N_4502);
or U4668 (N_4668,N_4460,N_4563);
nand U4669 (N_4669,N_4574,N_4530);
nand U4670 (N_4670,N_4406,N_4462);
or U4671 (N_4671,N_4572,N_4471);
or U4672 (N_4672,N_4583,N_4504);
nor U4673 (N_4673,N_4432,N_4429);
nand U4674 (N_4674,N_4475,N_4481);
or U4675 (N_4675,N_4458,N_4498);
nand U4676 (N_4676,N_4537,N_4402);
nand U4677 (N_4677,N_4430,N_4467);
or U4678 (N_4678,N_4454,N_4573);
nor U4679 (N_4679,N_4499,N_4480);
nand U4680 (N_4680,N_4592,N_4410);
nand U4681 (N_4681,N_4532,N_4408);
nand U4682 (N_4682,N_4596,N_4570);
nand U4683 (N_4683,N_4599,N_4571);
nor U4684 (N_4684,N_4477,N_4470);
nand U4685 (N_4685,N_4560,N_4490);
and U4686 (N_4686,N_4529,N_4551);
nand U4687 (N_4687,N_4428,N_4538);
and U4688 (N_4688,N_4535,N_4548);
or U4689 (N_4689,N_4488,N_4544);
nor U4690 (N_4690,N_4485,N_4449);
nor U4691 (N_4691,N_4553,N_4456);
or U4692 (N_4692,N_4482,N_4518);
nand U4693 (N_4693,N_4595,N_4558);
and U4694 (N_4694,N_4472,N_4457);
or U4695 (N_4695,N_4431,N_4598);
nand U4696 (N_4696,N_4500,N_4468);
xnor U4697 (N_4697,N_4546,N_4547);
nor U4698 (N_4698,N_4587,N_4584);
nor U4699 (N_4699,N_4491,N_4492);
and U4700 (N_4700,N_4446,N_4536);
and U4701 (N_4701,N_4543,N_4565);
and U4702 (N_4702,N_4490,N_4549);
and U4703 (N_4703,N_4483,N_4403);
nand U4704 (N_4704,N_4510,N_4460);
or U4705 (N_4705,N_4446,N_4552);
nor U4706 (N_4706,N_4530,N_4501);
or U4707 (N_4707,N_4576,N_4573);
or U4708 (N_4708,N_4407,N_4454);
xor U4709 (N_4709,N_4545,N_4525);
nor U4710 (N_4710,N_4475,N_4427);
nand U4711 (N_4711,N_4596,N_4595);
and U4712 (N_4712,N_4511,N_4496);
nand U4713 (N_4713,N_4495,N_4595);
xor U4714 (N_4714,N_4454,N_4430);
nor U4715 (N_4715,N_4431,N_4549);
and U4716 (N_4716,N_4467,N_4578);
nand U4717 (N_4717,N_4570,N_4488);
and U4718 (N_4718,N_4522,N_4534);
and U4719 (N_4719,N_4514,N_4404);
nand U4720 (N_4720,N_4519,N_4480);
nor U4721 (N_4721,N_4465,N_4485);
or U4722 (N_4722,N_4468,N_4407);
nand U4723 (N_4723,N_4497,N_4529);
nor U4724 (N_4724,N_4563,N_4494);
or U4725 (N_4725,N_4431,N_4508);
and U4726 (N_4726,N_4499,N_4563);
or U4727 (N_4727,N_4516,N_4581);
or U4728 (N_4728,N_4449,N_4551);
nand U4729 (N_4729,N_4539,N_4507);
nor U4730 (N_4730,N_4405,N_4530);
nand U4731 (N_4731,N_4537,N_4541);
or U4732 (N_4732,N_4550,N_4457);
nand U4733 (N_4733,N_4454,N_4495);
xor U4734 (N_4734,N_4409,N_4458);
nand U4735 (N_4735,N_4431,N_4583);
nand U4736 (N_4736,N_4597,N_4584);
nor U4737 (N_4737,N_4455,N_4403);
nor U4738 (N_4738,N_4465,N_4549);
nor U4739 (N_4739,N_4587,N_4434);
and U4740 (N_4740,N_4423,N_4400);
or U4741 (N_4741,N_4460,N_4514);
or U4742 (N_4742,N_4479,N_4527);
and U4743 (N_4743,N_4545,N_4590);
and U4744 (N_4744,N_4442,N_4464);
or U4745 (N_4745,N_4596,N_4487);
xnor U4746 (N_4746,N_4503,N_4444);
nand U4747 (N_4747,N_4409,N_4576);
nand U4748 (N_4748,N_4463,N_4464);
or U4749 (N_4749,N_4492,N_4525);
nand U4750 (N_4750,N_4422,N_4556);
and U4751 (N_4751,N_4568,N_4504);
or U4752 (N_4752,N_4453,N_4430);
nand U4753 (N_4753,N_4455,N_4546);
or U4754 (N_4754,N_4478,N_4487);
nand U4755 (N_4755,N_4467,N_4471);
nand U4756 (N_4756,N_4467,N_4478);
nand U4757 (N_4757,N_4563,N_4542);
nor U4758 (N_4758,N_4480,N_4587);
nand U4759 (N_4759,N_4523,N_4470);
or U4760 (N_4760,N_4447,N_4589);
nor U4761 (N_4761,N_4452,N_4410);
and U4762 (N_4762,N_4434,N_4544);
or U4763 (N_4763,N_4559,N_4463);
nand U4764 (N_4764,N_4570,N_4544);
nor U4765 (N_4765,N_4427,N_4555);
nor U4766 (N_4766,N_4423,N_4467);
or U4767 (N_4767,N_4409,N_4496);
or U4768 (N_4768,N_4450,N_4401);
nand U4769 (N_4769,N_4494,N_4486);
nor U4770 (N_4770,N_4558,N_4518);
nand U4771 (N_4771,N_4584,N_4505);
and U4772 (N_4772,N_4567,N_4521);
and U4773 (N_4773,N_4416,N_4526);
nor U4774 (N_4774,N_4589,N_4569);
nor U4775 (N_4775,N_4527,N_4523);
and U4776 (N_4776,N_4411,N_4562);
nor U4777 (N_4777,N_4441,N_4521);
nor U4778 (N_4778,N_4431,N_4580);
nor U4779 (N_4779,N_4588,N_4480);
nand U4780 (N_4780,N_4536,N_4442);
and U4781 (N_4781,N_4460,N_4583);
nor U4782 (N_4782,N_4546,N_4432);
xor U4783 (N_4783,N_4466,N_4494);
nand U4784 (N_4784,N_4414,N_4494);
and U4785 (N_4785,N_4576,N_4518);
nor U4786 (N_4786,N_4427,N_4474);
and U4787 (N_4787,N_4423,N_4529);
and U4788 (N_4788,N_4438,N_4401);
nand U4789 (N_4789,N_4439,N_4484);
nand U4790 (N_4790,N_4434,N_4597);
and U4791 (N_4791,N_4554,N_4540);
and U4792 (N_4792,N_4496,N_4526);
nand U4793 (N_4793,N_4556,N_4457);
nand U4794 (N_4794,N_4431,N_4566);
nand U4795 (N_4795,N_4574,N_4426);
nor U4796 (N_4796,N_4535,N_4457);
and U4797 (N_4797,N_4529,N_4436);
nand U4798 (N_4798,N_4472,N_4552);
nor U4799 (N_4799,N_4524,N_4488);
nand U4800 (N_4800,N_4730,N_4659);
or U4801 (N_4801,N_4653,N_4783);
nand U4802 (N_4802,N_4614,N_4792);
and U4803 (N_4803,N_4649,N_4746);
xnor U4804 (N_4804,N_4799,N_4698);
nor U4805 (N_4805,N_4761,N_4661);
nand U4806 (N_4806,N_4677,N_4683);
nor U4807 (N_4807,N_4779,N_4611);
or U4808 (N_4808,N_4780,N_4702);
and U4809 (N_4809,N_4737,N_4726);
or U4810 (N_4810,N_4633,N_4766);
or U4811 (N_4811,N_4699,N_4727);
or U4812 (N_4812,N_4763,N_4605);
or U4813 (N_4813,N_4689,N_4708);
or U4814 (N_4814,N_4603,N_4786);
and U4815 (N_4815,N_4640,N_4788);
or U4816 (N_4816,N_4607,N_4753);
nor U4817 (N_4817,N_4688,N_4756);
nor U4818 (N_4818,N_4624,N_4602);
and U4819 (N_4819,N_4666,N_4631);
nand U4820 (N_4820,N_4728,N_4636);
and U4821 (N_4821,N_4774,N_4718);
nand U4822 (N_4822,N_4711,N_4644);
xnor U4823 (N_4823,N_4684,N_4751);
and U4824 (N_4824,N_4608,N_4634);
nand U4825 (N_4825,N_4772,N_4630);
and U4826 (N_4826,N_4771,N_4738);
or U4827 (N_4827,N_4765,N_4669);
or U4828 (N_4828,N_4660,N_4748);
and U4829 (N_4829,N_4662,N_4721);
nand U4830 (N_4830,N_4693,N_4676);
nor U4831 (N_4831,N_4648,N_4674);
and U4832 (N_4832,N_4794,N_4637);
or U4833 (N_4833,N_4638,N_4769);
nor U4834 (N_4834,N_4663,N_4785);
nor U4835 (N_4835,N_4629,N_4675);
nand U4836 (N_4836,N_4620,N_4736);
xor U4837 (N_4837,N_4600,N_4796);
nand U4838 (N_4838,N_4686,N_4628);
nand U4839 (N_4839,N_4705,N_4768);
nand U4840 (N_4840,N_4687,N_4784);
nor U4841 (N_4841,N_4619,N_4673);
or U4842 (N_4842,N_4627,N_4703);
or U4843 (N_4843,N_4715,N_4734);
nor U4844 (N_4844,N_4680,N_4787);
and U4845 (N_4845,N_4606,N_4665);
nor U4846 (N_4846,N_4710,N_4615);
nor U4847 (N_4847,N_4782,N_4621);
nand U4848 (N_4848,N_4760,N_4739);
and U4849 (N_4849,N_4747,N_4613);
and U4850 (N_4850,N_4793,N_4672);
nand U4851 (N_4851,N_4789,N_4729);
nor U4852 (N_4852,N_4623,N_4712);
nand U4853 (N_4853,N_4609,N_4740);
and U4854 (N_4854,N_4668,N_4612);
nor U4855 (N_4855,N_4707,N_4685);
or U4856 (N_4856,N_4670,N_4691);
or U4857 (N_4857,N_4656,N_4758);
nand U4858 (N_4858,N_4724,N_4719);
nand U4859 (N_4859,N_4657,N_4790);
nor U4860 (N_4860,N_4641,N_4639);
nor U4861 (N_4861,N_4642,N_4647);
nor U4862 (N_4862,N_4678,N_4695);
nand U4863 (N_4863,N_4781,N_4692);
xor U4864 (N_4864,N_4749,N_4601);
nand U4865 (N_4865,N_4795,N_4625);
nand U4866 (N_4866,N_4752,N_4731);
nor U4867 (N_4867,N_4770,N_4798);
xor U4868 (N_4868,N_4775,N_4651);
or U4869 (N_4869,N_4755,N_4701);
nand U4870 (N_4870,N_4632,N_4776);
nand U4871 (N_4871,N_4650,N_4744);
and U4872 (N_4872,N_4654,N_4645);
nor U4873 (N_4873,N_4714,N_4618);
nor U4874 (N_4874,N_4754,N_4713);
and U4875 (N_4875,N_4697,N_4646);
and U4876 (N_4876,N_4694,N_4706);
or U4877 (N_4877,N_4635,N_4762);
nand U4878 (N_4878,N_4622,N_4791);
or U4879 (N_4879,N_4696,N_4709);
nand U4880 (N_4880,N_4759,N_4652);
or U4881 (N_4881,N_4723,N_4777);
or U4882 (N_4882,N_4704,N_4750);
or U4883 (N_4883,N_4626,N_4664);
nand U4884 (N_4884,N_4658,N_4733);
or U4885 (N_4885,N_4616,N_4610);
and U4886 (N_4886,N_4655,N_4778);
or U4887 (N_4887,N_4757,N_4681);
nor U4888 (N_4888,N_4720,N_4742);
nand U4889 (N_4889,N_4643,N_4725);
nor U4890 (N_4890,N_4679,N_4741);
nand U4891 (N_4891,N_4700,N_4732);
and U4892 (N_4892,N_4671,N_4604);
or U4893 (N_4893,N_4745,N_4667);
and U4894 (N_4894,N_4797,N_4743);
nand U4895 (N_4895,N_4767,N_4682);
nor U4896 (N_4896,N_4716,N_4717);
nor U4897 (N_4897,N_4722,N_4617);
and U4898 (N_4898,N_4735,N_4690);
nor U4899 (N_4899,N_4764,N_4773);
or U4900 (N_4900,N_4782,N_4788);
nand U4901 (N_4901,N_4743,N_4634);
or U4902 (N_4902,N_4627,N_4621);
nand U4903 (N_4903,N_4748,N_4762);
or U4904 (N_4904,N_4775,N_4706);
and U4905 (N_4905,N_4680,N_4769);
and U4906 (N_4906,N_4742,N_4771);
or U4907 (N_4907,N_4755,N_4605);
nor U4908 (N_4908,N_4755,N_4670);
or U4909 (N_4909,N_4770,N_4721);
and U4910 (N_4910,N_4790,N_4799);
nor U4911 (N_4911,N_4722,N_4624);
nor U4912 (N_4912,N_4735,N_4756);
and U4913 (N_4913,N_4775,N_4787);
or U4914 (N_4914,N_4704,N_4651);
nor U4915 (N_4915,N_4775,N_4631);
or U4916 (N_4916,N_4735,N_4770);
xor U4917 (N_4917,N_4777,N_4765);
or U4918 (N_4918,N_4675,N_4703);
nor U4919 (N_4919,N_4693,N_4738);
and U4920 (N_4920,N_4795,N_4786);
nand U4921 (N_4921,N_4731,N_4712);
and U4922 (N_4922,N_4648,N_4604);
xor U4923 (N_4923,N_4788,N_4787);
or U4924 (N_4924,N_4743,N_4733);
nand U4925 (N_4925,N_4772,N_4662);
nand U4926 (N_4926,N_4712,N_4640);
nor U4927 (N_4927,N_4672,N_4622);
and U4928 (N_4928,N_4635,N_4707);
or U4929 (N_4929,N_4604,N_4698);
nor U4930 (N_4930,N_4785,N_4793);
or U4931 (N_4931,N_4673,N_4685);
and U4932 (N_4932,N_4601,N_4682);
and U4933 (N_4933,N_4795,N_4663);
nor U4934 (N_4934,N_4711,N_4638);
xor U4935 (N_4935,N_4730,N_4797);
nor U4936 (N_4936,N_4641,N_4705);
nand U4937 (N_4937,N_4643,N_4647);
nand U4938 (N_4938,N_4660,N_4616);
nand U4939 (N_4939,N_4667,N_4672);
nor U4940 (N_4940,N_4688,N_4745);
nor U4941 (N_4941,N_4619,N_4778);
and U4942 (N_4942,N_4769,N_4796);
or U4943 (N_4943,N_4780,N_4677);
nand U4944 (N_4944,N_4619,N_4607);
nor U4945 (N_4945,N_4688,N_4625);
xnor U4946 (N_4946,N_4745,N_4795);
nand U4947 (N_4947,N_4691,N_4771);
nor U4948 (N_4948,N_4737,N_4763);
nand U4949 (N_4949,N_4723,N_4715);
and U4950 (N_4950,N_4736,N_4729);
nand U4951 (N_4951,N_4720,N_4601);
nand U4952 (N_4952,N_4768,N_4790);
nand U4953 (N_4953,N_4656,N_4761);
and U4954 (N_4954,N_4687,N_4602);
nor U4955 (N_4955,N_4784,N_4620);
and U4956 (N_4956,N_4729,N_4738);
nand U4957 (N_4957,N_4697,N_4767);
nand U4958 (N_4958,N_4779,N_4663);
or U4959 (N_4959,N_4672,N_4619);
nor U4960 (N_4960,N_4684,N_4756);
nor U4961 (N_4961,N_4798,N_4773);
or U4962 (N_4962,N_4697,N_4737);
or U4963 (N_4963,N_4719,N_4765);
nor U4964 (N_4964,N_4652,N_4771);
nand U4965 (N_4965,N_4738,N_4757);
nand U4966 (N_4966,N_4768,N_4703);
nand U4967 (N_4967,N_4627,N_4622);
nor U4968 (N_4968,N_4710,N_4670);
and U4969 (N_4969,N_4742,N_4725);
nor U4970 (N_4970,N_4713,N_4782);
or U4971 (N_4971,N_4615,N_4604);
or U4972 (N_4972,N_4650,N_4747);
nor U4973 (N_4973,N_4652,N_4614);
nor U4974 (N_4974,N_4664,N_4781);
or U4975 (N_4975,N_4752,N_4725);
and U4976 (N_4976,N_4734,N_4605);
or U4977 (N_4977,N_4711,N_4766);
and U4978 (N_4978,N_4747,N_4632);
and U4979 (N_4979,N_4724,N_4679);
nor U4980 (N_4980,N_4662,N_4727);
nor U4981 (N_4981,N_4685,N_4728);
nand U4982 (N_4982,N_4629,N_4615);
or U4983 (N_4983,N_4617,N_4600);
or U4984 (N_4984,N_4725,N_4661);
or U4985 (N_4985,N_4782,N_4756);
nor U4986 (N_4986,N_4625,N_4791);
nand U4987 (N_4987,N_4728,N_4630);
nand U4988 (N_4988,N_4752,N_4779);
xnor U4989 (N_4989,N_4733,N_4768);
nor U4990 (N_4990,N_4788,N_4666);
nor U4991 (N_4991,N_4657,N_4653);
nand U4992 (N_4992,N_4757,N_4695);
nand U4993 (N_4993,N_4735,N_4744);
and U4994 (N_4994,N_4639,N_4654);
nand U4995 (N_4995,N_4743,N_4681);
or U4996 (N_4996,N_4637,N_4618);
nor U4997 (N_4997,N_4692,N_4646);
nand U4998 (N_4998,N_4641,N_4731);
nand U4999 (N_4999,N_4641,N_4611);
or U5000 (N_5000,N_4930,N_4886);
nand U5001 (N_5001,N_4946,N_4940);
and U5002 (N_5002,N_4983,N_4980);
nor U5003 (N_5003,N_4819,N_4907);
nand U5004 (N_5004,N_4929,N_4884);
nand U5005 (N_5005,N_4936,N_4827);
nor U5006 (N_5006,N_4947,N_4978);
nor U5007 (N_5007,N_4913,N_4993);
and U5008 (N_5008,N_4953,N_4988);
nand U5009 (N_5009,N_4964,N_4891);
nand U5010 (N_5010,N_4896,N_4915);
nor U5011 (N_5011,N_4997,N_4872);
nor U5012 (N_5012,N_4948,N_4898);
and U5013 (N_5013,N_4981,N_4870);
and U5014 (N_5014,N_4899,N_4958);
nand U5015 (N_5015,N_4949,N_4882);
and U5016 (N_5016,N_4877,N_4905);
nor U5017 (N_5017,N_4873,N_4811);
nand U5018 (N_5018,N_4821,N_4863);
or U5019 (N_5019,N_4967,N_4864);
nor U5020 (N_5020,N_4815,N_4977);
or U5021 (N_5021,N_4973,N_4830);
and U5022 (N_5022,N_4808,N_4956);
and U5023 (N_5023,N_4901,N_4817);
nor U5024 (N_5024,N_4893,N_4825);
nand U5025 (N_5025,N_4971,N_4826);
nor U5026 (N_5026,N_4895,N_4854);
and U5027 (N_5027,N_4881,N_4985);
xnor U5028 (N_5028,N_4912,N_4918);
and U5029 (N_5029,N_4810,N_4813);
xnor U5030 (N_5030,N_4911,N_4875);
nand U5031 (N_5031,N_4996,N_4851);
and U5032 (N_5032,N_4920,N_4954);
and U5033 (N_5033,N_4848,N_4922);
or U5034 (N_5034,N_4982,N_4932);
and U5035 (N_5035,N_4968,N_4974);
and U5036 (N_5036,N_4951,N_4857);
and U5037 (N_5037,N_4904,N_4818);
or U5038 (N_5038,N_4855,N_4806);
and U5039 (N_5039,N_4829,N_4916);
nor U5040 (N_5040,N_4871,N_4824);
nor U5041 (N_5041,N_4987,N_4924);
xnor U5042 (N_5042,N_4846,N_4903);
nor U5043 (N_5043,N_4861,N_4931);
and U5044 (N_5044,N_4820,N_4975);
or U5045 (N_5045,N_4942,N_4856);
or U5046 (N_5046,N_4986,N_4945);
nor U5047 (N_5047,N_4853,N_4937);
and U5048 (N_5048,N_4906,N_4850);
nand U5049 (N_5049,N_4805,N_4888);
nor U5050 (N_5050,N_4939,N_4828);
and U5051 (N_5051,N_4897,N_4844);
or U5052 (N_5052,N_4835,N_4803);
or U5053 (N_5053,N_4972,N_4952);
or U5054 (N_5054,N_4832,N_4992);
and U5055 (N_5055,N_4822,N_4837);
nor U5056 (N_5056,N_4860,N_4957);
or U5057 (N_5057,N_4925,N_4921);
nor U5058 (N_5058,N_4943,N_4923);
and U5059 (N_5059,N_4950,N_4814);
nor U5060 (N_5060,N_4935,N_4926);
nand U5061 (N_5061,N_4970,N_4991);
or U5062 (N_5062,N_4847,N_4892);
nor U5063 (N_5063,N_4800,N_4914);
nand U5064 (N_5064,N_4885,N_4878);
nor U5065 (N_5065,N_4879,N_4959);
nand U5066 (N_5066,N_4866,N_4989);
nor U5067 (N_5067,N_4842,N_4840);
or U5068 (N_5068,N_4955,N_4867);
nand U5069 (N_5069,N_4999,N_4816);
and U5070 (N_5070,N_4963,N_4961);
and U5071 (N_5071,N_4910,N_4998);
nand U5072 (N_5072,N_4836,N_4938);
nand U5073 (N_5073,N_4858,N_4839);
xor U5074 (N_5074,N_4928,N_4902);
nor U5075 (N_5075,N_4995,N_4979);
or U5076 (N_5076,N_4976,N_4944);
and U5077 (N_5077,N_4843,N_4809);
nor U5078 (N_5078,N_4941,N_4934);
nand U5079 (N_5079,N_4804,N_4838);
nor U5080 (N_5080,N_4894,N_4984);
and U5081 (N_5081,N_4868,N_4917);
nor U5082 (N_5082,N_4801,N_4969);
nand U5083 (N_5083,N_4859,N_4862);
nor U5084 (N_5084,N_4994,N_4845);
nor U5085 (N_5085,N_4887,N_4889);
nor U5086 (N_5086,N_4841,N_4874);
nor U5087 (N_5087,N_4965,N_4966);
nand U5088 (N_5088,N_4962,N_4933);
or U5089 (N_5089,N_4812,N_4876);
nor U5090 (N_5090,N_4833,N_4927);
and U5091 (N_5091,N_4834,N_4890);
nand U5092 (N_5092,N_4919,N_4880);
nor U5093 (N_5093,N_4869,N_4960);
and U5094 (N_5094,N_4831,N_4865);
and U5095 (N_5095,N_4908,N_4900);
nand U5096 (N_5096,N_4849,N_4990);
nand U5097 (N_5097,N_4807,N_4802);
and U5098 (N_5098,N_4823,N_4909);
nor U5099 (N_5099,N_4852,N_4883);
nor U5100 (N_5100,N_4913,N_4800);
nor U5101 (N_5101,N_4951,N_4990);
or U5102 (N_5102,N_4852,N_4846);
nor U5103 (N_5103,N_4840,N_4904);
nor U5104 (N_5104,N_4920,N_4820);
or U5105 (N_5105,N_4876,N_4959);
nor U5106 (N_5106,N_4833,N_4864);
or U5107 (N_5107,N_4983,N_4925);
or U5108 (N_5108,N_4844,N_4911);
nor U5109 (N_5109,N_4957,N_4972);
and U5110 (N_5110,N_4902,N_4823);
nor U5111 (N_5111,N_4839,N_4863);
nor U5112 (N_5112,N_4988,N_4856);
nand U5113 (N_5113,N_4898,N_4851);
and U5114 (N_5114,N_4862,N_4810);
nor U5115 (N_5115,N_4972,N_4977);
nand U5116 (N_5116,N_4837,N_4937);
nand U5117 (N_5117,N_4890,N_4979);
or U5118 (N_5118,N_4881,N_4868);
and U5119 (N_5119,N_4989,N_4886);
and U5120 (N_5120,N_4979,N_4927);
or U5121 (N_5121,N_4930,N_4942);
or U5122 (N_5122,N_4896,N_4835);
or U5123 (N_5123,N_4962,N_4826);
and U5124 (N_5124,N_4953,N_4903);
nand U5125 (N_5125,N_4921,N_4959);
nor U5126 (N_5126,N_4816,N_4860);
nand U5127 (N_5127,N_4935,N_4827);
nor U5128 (N_5128,N_4862,N_4958);
and U5129 (N_5129,N_4990,N_4915);
nand U5130 (N_5130,N_4905,N_4813);
nand U5131 (N_5131,N_4990,N_4893);
nand U5132 (N_5132,N_4933,N_4821);
or U5133 (N_5133,N_4943,N_4942);
and U5134 (N_5134,N_4988,N_4854);
nand U5135 (N_5135,N_4966,N_4830);
and U5136 (N_5136,N_4899,N_4968);
and U5137 (N_5137,N_4980,N_4848);
and U5138 (N_5138,N_4893,N_4839);
or U5139 (N_5139,N_4987,N_4950);
and U5140 (N_5140,N_4890,N_4932);
or U5141 (N_5141,N_4925,N_4978);
or U5142 (N_5142,N_4921,N_4806);
nor U5143 (N_5143,N_4923,N_4891);
and U5144 (N_5144,N_4903,N_4938);
nor U5145 (N_5145,N_4961,N_4833);
nor U5146 (N_5146,N_4904,N_4905);
nor U5147 (N_5147,N_4853,N_4807);
or U5148 (N_5148,N_4856,N_4996);
nand U5149 (N_5149,N_4902,N_4856);
or U5150 (N_5150,N_4962,N_4966);
nor U5151 (N_5151,N_4836,N_4851);
and U5152 (N_5152,N_4966,N_4943);
and U5153 (N_5153,N_4917,N_4936);
nand U5154 (N_5154,N_4862,N_4979);
nor U5155 (N_5155,N_4942,N_4906);
or U5156 (N_5156,N_4955,N_4970);
nand U5157 (N_5157,N_4831,N_4907);
nand U5158 (N_5158,N_4919,N_4878);
and U5159 (N_5159,N_4958,N_4887);
or U5160 (N_5160,N_4968,N_4869);
nor U5161 (N_5161,N_4976,N_4967);
or U5162 (N_5162,N_4903,N_4880);
nor U5163 (N_5163,N_4897,N_4822);
or U5164 (N_5164,N_4902,N_4895);
and U5165 (N_5165,N_4861,N_4860);
nor U5166 (N_5166,N_4834,N_4953);
and U5167 (N_5167,N_4927,N_4887);
xor U5168 (N_5168,N_4830,N_4922);
nor U5169 (N_5169,N_4956,N_4860);
and U5170 (N_5170,N_4884,N_4869);
or U5171 (N_5171,N_4875,N_4841);
nor U5172 (N_5172,N_4876,N_4992);
nand U5173 (N_5173,N_4909,N_4859);
nor U5174 (N_5174,N_4901,N_4881);
or U5175 (N_5175,N_4963,N_4879);
or U5176 (N_5176,N_4995,N_4828);
or U5177 (N_5177,N_4928,N_4916);
nor U5178 (N_5178,N_4843,N_4968);
nor U5179 (N_5179,N_4905,N_4917);
nand U5180 (N_5180,N_4881,N_4807);
and U5181 (N_5181,N_4810,N_4912);
and U5182 (N_5182,N_4889,N_4858);
nor U5183 (N_5183,N_4915,N_4803);
or U5184 (N_5184,N_4826,N_4934);
and U5185 (N_5185,N_4854,N_4911);
nand U5186 (N_5186,N_4925,N_4971);
or U5187 (N_5187,N_4931,N_4961);
nor U5188 (N_5188,N_4866,N_4947);
and U5189 (N_5189,N_4974,N_4807);
or U5190 (N_5190,N_4806,N_4985);
nor U5191 (N_5191,N_4992,N_4997);
nand U5192 (N_5192,N_4838,N_4835);
nor U5193 (N_5193,N_4975,N_4911);
nand U5194 (N_5194,N_4950,N_4886);
nand U5195 (N_5195,N_4974,N_4813);
or U5196 (N_5196,N_4812,N_4954);
nor U5197 (N_5197,N_4969,N_4894);
xnor U5198 (N_5198,N_4888,N_4939);
and U5199 (N_5199,N_4903,N_4851);
or U5200 (N_5200,N_5053,N_5032);
nor U5201 (N_5201,N_5172,N_5045);
or U5202 (N_5202,N_5096,N_5169);
nand U5203 (N_5203,N_5118,N_5183);
nand U5204 (N_5204,N_5047,N_5198);
or U5205 (N_5205,N_5018,N_5048);
nor U5206 (N_5206,N_5109,N_5072);
xnor U5207 (N_5207,N_5086,N_5008);
nor U5208 (N_5208,N_5091,N_5116);
nand U5209 (N_5209,N_5023,N_5120);
and U5210 (N_5210,N_5154,N_5166);
and U5211 (N_5211,N_5052,N_5014);
or U5212 (N_5212,N_5140,N_5179);
and U5213 (N_5213,N_5020,N_5002);
nand U5214 (N_5214,N_5015,N_5197);
and U5215 (N_5215,N_5163,N_5159);
or U5216 (N_5216,N_5124,N_5035);
nand U5217 (N_5217,N_5027,N_5057);
and U5218 (N_5218,N_5176,N_5126);
or U5219 (N_5219,N_5122,N_5100);
and U5220 (N_5220,N_5142,N_5075);
and U5221 (N_5221,N_5068,N_5152);
or U5222 (N_5222,N_5074,N_5164);
xor U5223 (N_5223,N_5193,N_5061);
and U5224 (N_5224,N_5151,N_5041);
nand U5225 (N_5225,N_5021,N_5175);
nand U5226 (N_5226,N_5055,N_5173);
or U5227 (N_5227,N_5155,N_5016);
and U5228 (N_5228,N_5150,N_5059);
nand U5229 (N_5229,N_5167,N_5121);
and U5230 (N_5230,N_5178,N_5030);
nor U5231 (N_5231,N_5199,N_5099);
and U5232 (N_5232,N_5063,N_5054);
nand U5233 (N_5233,N_5181,N_5135);
or U5234 (N_5234,N_5034,N_5125);
nor U5235 (N_5235,N_5005,N_5180);
nand U5236 (N_5236,N_5132,N_5006);
nand U5237 (N_5237,N_5046,N_5079);
or U5238 (N_5238,N_5190,N_5082);
and U5239 (N_5239,N_5042,N_5105);
nand U5240 (N_5240,N_5094,N_5127);
nor U5241 (N_5241,N_5157,N_5108);
or U5242 (N_5242,N_5113,N_5028);
nand U5243 (N_5243,N_5146,N_5187);
nor U5244 (N_5244,N_5168,N_5103);
and U5245 (N_5245,N_5141,N_5170);
and U5246 (N_5246,N_5087,N_5081);
nand U5247 (N_5247,N_5065,N_5011);
and U5248 (N_5248,N_5145,N_5085);
nand U5249 (N_5249,N_5004,N_5149);
or U5250 (N_5250,N_5038,N_5076);
nand U5251 (N_5251,N_5130,N_5066);
nand U5252 (N_5252,N_5185,N_5069);
nand U5253 (N_5253,N_5097,N_5119);
nand U5254 (N_5254,N_5196,N_5022);
or U5255 (N_5255,N_5123,N_5143);
nor U5256 (N_5256,N_5128,N_5182);
and U5257 (N_5257,N_5037,N_5110);
nor U5258 (N_5258,N_5184,N_5129);
or U5259 (N_5259,N_5115,N_5177);
and U5260 (N_5260,N_5160,N_5165);
nor U5261 (N_5261,N_5114,N_5001);
or U5262 (N_5262,N_5111,N_5117);
and U5263 (N_5263,N_5089,N_5036);
or U5264 (N_5264,N_5013,N_5092);
nand U5265 (N_5265,N_5138,N_5078);
nor U5266 (N_5266,N_5106,N_5049);
nand U5267 (N_5267,N_5186,N_5148);
nor U5268 (N_5268,N_5070,N_5007);
nand U5269 (N_5269,N_5077,N_5024);
nor U5270 (N_5270,N_5031,N_5033);
and U5271 (N_5271,N_5067,N_5073);
or U5272 (N_5272,N_5194,N_5131);
and U5273 (N_5273,N_5161,N_5000);
and U5274 (N_5274,N_5153,N_5058);
nand U5275 (N_5275,N_5010,N_5029);
and U5276 (N_5276,N_5095,N_5084);
nand U5277 (N_5277,N_5195,N_5189);
or U5278 (N_5278,N_5158,N_5192);
xor U5279 (N_5279,N_5019,N_5040);
or U5280 (N_5280,N_5104,N_5050);
and U5281 (N_5281,N_5025,N_5003);
nand U5282 (N_5282,N_5136,N_5134);
nor U5283 (N_5283,N_5051,N_5156);
nand U5284 (N_5284,N_5093,N_5174);
or U5285 (N_5285,N_5071,N_5112);
nand U5286 (N_5286,N_5090,N_5043);
nand U5287 (N_5287,N_5144,N_5060);
nor U5288 (N_5288,N_5171,N_5102);
nand U5289 (N_5289,N_5026,N_5062);
or U5290 (N_5290,N_5137,N_5107);
and U5291 (N_5291,N_5191,N_5101);
and U5292 (N_5292,N_5147,N_5012);
and U5293 (N_5293,N_5009,N_5044);
xnor U5294 (N_5294,N_5162,N_5188);
and U5295 (N_5295,N_5133,N_5056);
nand U5296 (N_5296,N_5139,N_5039);
and U5297 (N_5297,N_5080,N_5098);
or U5298 (N_5298,N_5017,N_5083);
nor U5299 (N_5299,N_5064,N_5088);
and U5300 (N_5300,N_5128,N_5047);
nor U5301 (N_5301,N_5036,N_5098);
nand U5302 (N_5302,N_5122,N_5068);
or U5303 (N_5303,N_5150,N_5009);
nor U5304 (N_5304,N_5073,N_5184);
or U5305 (N_5305,N_5196,N_5164);
and U5306 (N_5306,N_5066,N_5080);
nor U5307 (N_5307,N_5151,N_5003);
or U5308 (N_5308,N_5030,N_5164);
nor U5309 (N_5309,N_5140,N_5076);
and U5310 (N_5310,N_5007,N_5165);
and U5311 (N_5311,N_5177,N_5118);
nor U5312 (N_5312,N_5042,N_5021);
nand U5313 (N_5313,N_5078,N_5050);
and U5314 (N_5314,N_5147,N_5192);
nand U5315 (N_5315,N_5139,N_5057);
nand U5316 (N_5316,N_5103,N_5051);
nor U5317 (N_5317,N_5111,N_5008);
and U5318 (N_5318,N_5051,N_5189);
or U5319 (N_5319,N_5181,N_5017);
or U5320 (N_5320,N_5056,N_5154);
and U5321 (N_5321,N_5158,N_5119);
nand U5322 (N_5322,N_5028,N_5156);
or U5323 (N_5323,N_5066,N_5044);
nand U5324 (N_5324,N_5165,N_5090);
and U5325 (N_5325,N_5005,N_5124);
and U5326 (N_5326,N_5193,N_5165);
and U5327 (N_5327,N_5101,N_5035);
nand U5328 (N_5328,N_5135,N_5090);
or U5329 (N_5329,N_5162,N_5130);
nand U5330 (N_5330,N_5022,N_5091);
and U5331 (N_5331,N_5157,N_5166);
and U5332 (N_5332,N_5074,N_5124);
nand U5333 (N_5333,N_5135,N_5187);
and U5334 (N_5334,N_5034,N_5112);
nand U5335 (N_5335,N_5018,N_5037);
and U5336 (N_5336,N_5097,N_5159);
nor U5337 (N_5337,N_5004,N_5053);
nand U5338 (N_5338,N_5084,N_5129);
nor U5339 (N_5339,N_5189,N_5094);
xnor U5340 (N_5340,N_5196,N_5009);
or U5341 (N_5341,N_5159,N_5071);
or U5342 (N_5342,N_5064,N_5168);
and U5343 (N_5343,N_5174,N_5145);
or U5344 (N_5344,N_5187,N_5175);
nand U5345 (N_5345,N_5013,N_5075);
or U5346 (N_5346,N_5117,N_5094);
or U5347 (N_5347,N_5099,N_5147);
nor U5348 (N_5348,N_5162,N_5104);
nand U5349 (N_5349,N_5144,N_5028);
nor U5350 (N_5350,N_5094,N_5039);
nand U5351 (N_5351,N_5125,N_5168);
nand U5352 (N_5352,N_5098,N_5017);
or U5353 (N_5353,N_5081,N_5032);
or U5354 (N_5354,N_5185,N_5028);
and U5355 (N_5355,N_5161,N_5022);
and U5356 (N_5356,N_5191,N_5063);
and U5357 (N_5357,N_5129,N_5098);
and U5358 (N_5358,N_5007,N_5032);
nand U5359 (N_5359,N_5026,N_5175);
nand U5360 (N_5360,N_5067,N_5121);
nor U5361 (N_5361,N_5011,N_5036);
nor U5362 (N_5362,N_5175,N_5174);
and U5363 (N_5363,N_5097,N_5125);
nand U5364 (N_5364,N_5192,N_5106);
nand U5365 (N_5365,N_5019,N_5074);
nand U5366 (N_5366,N_5115,N_5190);
nor U5367 (N_5367,N_5076,N_5175);
or U5368 (N_5368,N_5105,N_5171);
nand U5369 (N_5369,N_5145,N_5172);
nor U5370 (N_5370,N_5097,N_5140);
and U5371 (N_5371,N_5113,N_5141);
nor U5372 (N_5372,N_5144,N_5078);
and U5373 (N_5373,N_5022,N_5034);
and U5374 (N_5374,N_5076,N_5083);
nand U5375 (N_5375,N_5002,N_5089);
or U5376 (N_5376,N_5098,N_5157);
nor U5377 (N_5377,N_5101,N_5045);
xnor U5378 (N_5378,N_5133,N_5032);
nor U5379 (N_5379,N_5061,N_5137);
or U5380 (N_5380,N_5132,N_5127);
or U5381 (N_5381,N_5128,N_5178);
nand U5382 (N_5382,N_5123,N_5061);
nor U5383 (N_5383,N_5043,N_5143);
and U5384 (N_5384,N_5038,N_5022);
nand U5385 (N_5385,N_5026,N_5084);
and U5386 (N_5386,N_5112,N_5197);
xor U5387 (N_5387,N_5060,N_5120);
or U5388 (N_5388,N_5165,N_5178);
nor U5389 (N_5389,N_5115,N_5113);
or U5390 (N_5390,N_5135,N_5052);
nor U5391 (N_5391,N_5190,N_5139);
nor U5392 (N_5392,N_5034,N_5082);
or U5393 (N_5393,N_5024,N_5167);
and U5394 (N_5394,N_5100,N_5077);
and U5395 (N_5395,N_5187,N_5085);
nor U5396 (N_5396,N_5039,N_5185);
nand U5397 (N_5397,N_5174,N_5053);
nor U5398 (N_5398,N_5153,N_5103);
nand U5399 (N_5399,N_5128,N_5185);
or U5400 (N_5400,N_5352,N_5257);
xor U5401 (N_5401,N_5317,N_5262);
nand U5402 (N_5402,N_5320,N_5380);
nor U5403 (N_5403,N_5231,N_5319);
nor U5404 (N_5404,N_5373,N_5312);
nand U5405 (N_5405,N_5246,N_5349);
nor U5406 (N_5406,N_5266,N_5381);
or U5407 (N_5407,N_5211,N_5329);
or U5408 (N_5408,N_5267,N_5279);
nor U5409 (N_5409,N_5281,N_5280);
or U5410 (N_5410,N_5271,N_5238);
or U5411 (N_5411,N_5214,N_5367);
and U5412 (N_5412,N_5235,N_5393);
nor U5413 (N_5413,N_5276,N_5202);
or U5414 (N_5414,N_5234,N_5375);
and U5415 (N_5415,N_5368,N_5389);
nand U5416 (N_5416,N_5331,N_5362);
and U5417 (N_5417,N_5365,N_5283);
nor U5418 (N_5418,N_5201,N_5251);
nor U5419 (N_5419,N_5307,N_5204);
or U5420 (N_5420,N_5232,N_5203);
or U5421 (N_5421,N_5261,N_5296);
nand U5422 (N_5422,N_5314,N_5219);
nand U5423 (N_5423,N_5341,N_5302);
nor U5424 (N_5424,N_5218,N_5384);
and U5425 (N_5425,N_5294,N_5253);
or U5426 (N_5426,N_5372,N_5209);
and U5427 (N_5427,N_5395,N_5383);
nor U5428 (N_5428,N_5286,N_5321);
and U5429 (N_5429,N_5205,N_5217);
nand U5430 (N_5430,N_5340,N_5228);
or U5431 (N_5431,N_5369,N_5243);
nand U5432 (N_5432,N_5387,N_5354);
xor U5433 (N_5433,N_5297,N_5311);
and U5434 (N_5434,N_5325,N_5363);
nor U5435 (N_5435,N_5248,N_5336);
or U5436 (N_5436,N_5388,N_5298);
nor U5437 (N_5437,N_5345,N_5324);
nand U5438 (N_5438,N_5371,N_5390);
nor U5439 (N_5439,N_5301,N_5364);
and U5440 (N_5440,N_5350,N_5379);
xor U5441 (N_5441,N_5282,N_5288);
nand U5442 (N_5442,N_5338,N_5355);
nand U5443 (N_5443,N_5308,N_5237);
or U5444 (N_5444,N_5377,N_5357);
and U5445 (N_5445,N_5252,N_5318);
nor U5446 (N_5446,N_5240,N_5366);
nor U5447 (N_5447,N_5207,N_5226);
or U5448 (N_5448,N_5332,N_5254);
nor U5449 (N_5449,N_5351,N_5272);
nor U5450 (N_5450,N_5230,N_5374);
or U5451 (N_5451,N_5300,N_5391);
nand U5452 (N_5452,N_5268,N_5326);
nand U5453 (N_5453,N_5322,N_5208);
or U5454 (N_5454,N_5278,N_5200);
nand U5455 (N_5455,N_5275,N_5353);
and U5456 (N_5456,N_5227,N_5273);
xnor U5457 (N_5457,N_5323,N_5291);
xor U5458 (N_5458,N_5210,N_5358);
nand U5459 (N_5459,N_5347,N_5224);
nor U5460 (N_5460,N_5392,N_5225);
xor U5461 (N_5461,N_5335,N_5309);
nand U5462 (N_5462,N_5263,N_5216);
and U5463 (N_5463,N_5292,N_5299);
and U5464 (N_5464,N_5270,N_5333);
and U5465 (N_5465,N_5285,N_5303);
nor U5466 (N_5466,N_5342,N_5360);
nand U5467 (N_5467,N_5290,N_5239);
or U5468 (N_5468,N_5359,N_5394);
or U5469 (N_5469,N_5328,N_5382);
or U5470 (N_5470,N_5274,N_5313);
nand U5471 (N_5471,N_5236,N_5315);
nand U5472 (N_5472,N_5306,N_5293);
nand U5473 (N_5473,N_5304,N_5348);
nand U5474 (N_5474,N_5356,N_5378);
nor U5475 (N_5475,N_5386,N_5310);
nand U5476 (N_5476,N_5220,N_5346);
xor U5477 (N_5477,N_5245,N_5327);
or U5478 (N_5478,N_5206,N_5260);
nor U5479 (N_5479,N_5258,N_5344);
and U5480 (N_5480,N_5249,N_5399);
nor U5481 (N_5481,N_5250,N_5277);
or U5482 (N_5482,N_5337,N_5339);
or U5483 (N_5483,N_5221,N_5397);
and U5484 (N_5484,N_5212,N_5376);
or U5485 (N_5485,N_5330,N_5265);
or U5486 (N_5486,N_5229,N_5223);
and U5487 (N_5487,N_5305,N_5213);
nor U5488 (N_5488,N_5264,N_5295);
and U5489 (N_5489,N_5361,N_5241);
nor U5490 (N_5490,N_5255,N_5222);
and U5491 (N_5491,N_5398,N_5289);
nand U5492 (N_5492,N_5287,N_5256);
nand U5493 (N_5493,N_5284,N_5343);
nand U5494 (N_5494,N_5269,N_5370);
nand U5495 (N_5495,N_5385,N_5242);
or U5496 (N_5496,N_5259,N_5334);
nand U5497 (N_5497,N_5316,N_5215);
or U5498 (N_5498,N_5396,N_5233);
or U5499 (N_5499,N_5247,N_5244);
and U5500 (N_5500,N_5345,N_5259);
and U5501 (N_5501,N_5253,N_5267);
and U5502 (N_5502,N_5392,N_5228);
nor U5503 (N_5503,N_5374,N_5223);
and U5504 (N_5504,N_5385,N_5227);
or U5505 (N_5505,N_5235,N_5247);
and U5506 (N_5506,N_5312,N_5254);
or U5507 (N_5507,N_5222,N_5355);
and U5508 (N_5508,N_5250,N_5203);
and U5509 (N_5509,N_5295,N_5294);
xor U5510 (N_5510,N_5292,N_5214);
nand U5511 (N_5511,N_5312,N_5390);
nor U5512 (N_5512,N_5385,N_5372);
and U5513 (N_5513,N_5364,N_5218);
or U5514 (N_5514,N_5285,N_5355);
and U5515 (N_5515,N_5223,N_5264);
nand U5516 (N_5516,N_5251,N_5370);
nor U5517 (N_5517,N_5334,N_5381);
nand U5518 (N_5518,N_5238,N_5381);
nand U5519 (N_5519,N_5331,N_5215);
and U5520 (N_5520,N_5329,N_5331);
and U5521 (N_5521,N_5267,N_5304);
and U5522 (N_5522,N_5352,N_5210);
or U5523 (N_5523,N_5351,N_5315);
nand U5524 (N_5524,N_5248,N_5379);
or U5525 (N_5525,N_5374,N_5360);
and U5526 (N_5526,N_5297,N_5248);
and U5527 (N_5527,N_5371,N_5234);
nand U5528 (N_5528,N_5201,N_5237);
nand U5529 (N_5529,N_5360,N_5332);
and U5530 (N_5530,N_5348,N_5288);
or U5531 (N_5531,N_5370,N_5276);
or U5532 (N_5532,N_5363,N_5290);
nor U5533 (N_5533,N_5237,N_5303);
or U5534 (N_5534,N_5350,N_5316);
nand U5535 (N_5535,N_5310,N_5201);
or U5536 (N_5536,N_5355,N_5229);
or U5537 (N_5537,N_5362,N_5307);
and U5538 (N_5538,N_5232,N_5364);
nand U5539 (N_5539,N_5235,N_5386);
nand U5540 (N_5540,N_5345,N_5208);
nor U5541 (N_5541,N_5265,N_5314);
xor U5542 (N_5542,N_5267,N_5246);
and U5543 (N_5543,N_5334,N_5337);
nor U5544 (N_5544,N_5290,N_5397);
and U5545 (N_5545,N_5396,N_5341);
nand U5546 (N_5546,N_5319,N_5356);
nand U5547 (N_5547,N_5244,N_5281);
or U5548 (N_5548,N_5373,N_5392);
and U5549 (N_5549,N_5303,N_5202);
or U5550 (N_5550,N_5289,N_5287);
or U5551 (N_5551,N_5336,N_5218);
and U5552 (N_5552,N_5297,N_5251);
nand U5553 (N_5553,N_5252,N_5262);
xor U5554 (N_5554,N_5309,N_5327);
or U5555 (N_5555,N_5276,N_5356);
xor U5556 (N_5556,N_5352,N_5206);
and U5557 (N_5557,N_5289,N_5266);
nor U5558 (N_5558,N_5222,N_5333);
and U5559 (N_5559,N_5292,N_5288);
and U5560 (N_5560,N_5290,N_5208);
nand U5561 (N_5561,N_5305,N_5246);
and U5562 (N_5562,N_5212,N_5345);
nand U5563 (N_5563,N_5238,N_5399);
nand U5564 (N_5564,N_5356,N_5367);
and U5565 (N_5565,N_5254,N_5305);
nor U5566 (N_5566,N_5251,N_5360);
nand U5567 (N_5567,N_5345,N_5206);
nand U5568 (N_5568,N_5303,N_5354);
nand U5569 (N_5569,N_5250,N_5252);
nor U5570 (N_5570,N_5218,N_5208);
nand U5571 (N_5571,N_5281,N_5327);
nor U5572 (N_5572,N_5349,N_5208);
and U5573 (N_5573,N_5275,N_5240);
and U5574 (N_5574,N_5307,N_5303);
and U5575 (N_5575,N_5392,N_5316);
and U5576 (N_5576,N_5296,N_5288);
nand U5577 (N_5577,N_5279,N_5394);
and U5578 (N_5578,N_5271,N_5215);
nand U5579 (N_5579,N_5326,N_5228);
nor U5580 (N_5580,N_5311,N_5218);
and U5581 (N_5581,N_5313,N_5309);
nand U5582 (N_5582,N_5248,N_5281);
xor U5583 (N_5583,N_5274,N_5238);
xnor U5584 (N_5584,N_5261,N_5377);
nand U5585 (N_5585,N_5238,N_5265);
or U5586 (N_5586,N_5275,N_5312);
nand U5587 (N_5587,N_5292,N_5343);
or U5588 (N_5588,N_5247,N_5266);
nand U5589 (N_5589,N_5285,N_5312);
or U5590 (N_5590,N_5381,N_5328);
nand U5591 (N_5591,N_5352,N_5307);
and U5592 (N_5592,N_5334,N_5276);
nor U5593 (N_5593,N_5321,N_5381);
or U5594 (N_5594,N_5207,N_5264);
or U5595 (N_5595,N_5353,N_5280);
and U5596 (N_5596,N_5377,N_5273);
nand U5597 (N_5597,N_5289,N_5236);
nand U5598 (N_5598,N_5217,N_5201);
and U5599 (N_5599,N_5290,N_5389);
nor U5600 (N_5600,N_5566,N_5485);
nand U5601 (N_5601,N_5556,N_5438);
and U5602 (N_5602,N_5504,N_5445);
xor U5603 (N_5603,N_5559,N_5575);
or U5604 (N_5604,N_5529,N_5411);
or U5605 (N_5605,N_5552,N_5507);
or U5606 (N_5606,N_5410,N_5592);
and U5607 (N_5607,N_5549,N_5515);
and U5608 (N_5608,N_5571,N_5520);
nand U5609 (N_5609,N_5464,N_5400);
xnor U5610 (N_5610,N_5589,N_5542);
nand U5611 (N_5611,N_5468,N_5482);
or U5612 (N_5612,N_5490,N_5402);
nand U5613 (N_5613,N_5420,N_5456);
nor U5614 (N_5614,N_5569,N_5429);
nor U5615 (N_5615,N_5534,N_5572);
or U5616 (N_5616,N_5596,N_5498);
nor U5617 (N_5617,N_5412,N_5436);
nor U5618 (N_5618,N_5451,N_5594);
nand U5619 (N_5619,N_5413,N_5554);
or U5620 (N_5620,N_5461,N_5401);
or U5621 (N_5621,N_5519,N_5508);
and U5622 (N_5622,N_5532,N_5422);
nand U5623 (N_5623,N_5593,N_5491);
nand U5624 (N_5624,N_5553,N_5563);
or U5625 (N_5625,N_5417,N_5526);
nor U5626 (N_5626,N_5433,N_5435);
nand U5627 (N_5627,N_5540,N_5557);
or U5628 (N_5628,N_5474,N_5530);
nor U5629 (N_5629,N_5539,N_5460);
and U5630 (N_5630,N_5567,N_5469);
and U5631 (N_5631,N_5478,N_5423);
nand U5632 (N_5632,N_5505,N_5521);
nand U5633 (N_5633,N_5425,N_5579);
nand U5634 (N_5634,N_5470,N_5558);
nand U5635 (N_5635,N_5514,N_5424);
and U5636 (N_5636,N_5555,N_5409);
nand U5637 (N_5637,N_5500,N_5564);
nor U5638 (N_5638,N_5467,N_5568);
nand U5639 (N_5639,N_5450,N_5421);
or U5640 (N_5640,N_5414,N_5443);
nor U5641 (N_5641,N_5546,N_5455);
and U5642 (N_5642,N_5439,N_5502);
and U5643 (N_5643,N_5509,N_5501);
nor U5644 (N_5644,N_5440,N_5403);
nand U5645 (N_5645,N_5516,N_5416);
or U5646 (N_5646,N_5585,N_5475);
nand U5647 (N_5647,N_5426,N_5537);
nor U5648 (N_5648,N_5465,N_5432);
nand U5649 (N_5649,N_5427,N_5495);
nand U5650 (N_5650,N_5544,N_5578);
and U5651 (N_5651,N_5541,N_5570);
xor U5652 (N_5652,N_5430,N_5503);
and U5653 (N_5653,N_5488,N_5506);
and U5654 (N_5654,N_5573,N_5525);
and U5655 (N_5655,N_5582,N_5437);
and U5656 (N_5656,N_5512,N_5448);
and U5657 (N_5657,N_5459,N_5538);
nor U5658 (N_5658,N_5431,N_5595);
and U5659 (N_5659,N_5574,N_5551);
and U5660 (N_5660,N_5598,N_5577);
nor U5661 (N_5661,N_5444,N_5407);
nand U5662 (N_5662,N_5550,N_5536);
nor U5663 (N_5663,N_5547,N_5493);
nand U5664 (N_5664,N_5419,N_5406);
nor U5665 (N_5665,N_5408,N_5418);
nand U5666 (N_5666,N_5489,N_5528);
nor U5667 (N_5667,N_5524,N_5580);
or U5668 (N_5668,N_5587,N_5442);
nand U5669 (N_5669,N_5597,N_5499);
nand U5670 (N_5670,N_5458,N_5484);
nor U5671 (N_5671,N_5449,N_5492);
nor U5672 (N_5672,N_5487,N_5466);
and U5673 (N_5673,N_5513,N_5472);
nor U5674 (N_5674,N_5565,N_5548);
nand U5675 (N_5675,N_5428,N_5457);
nor U5676 (N_5676,N_5446,N_5527);
nand U5677 (N_5677,N_5496,N_5545);
nor U5678 (N_5678,N_5599,N_5497);
and U5679 (N_5679,N_5562,N_5447);
or U5680 (N_5680,N_5480,N_5583);
or U5681 (N_5681,N_5494,N_5576);
and U5682 (N_5682,N_5560,N_5543);
nand U5683 (N_5683,N_5523,N_5481);
nand U5684 (N_5684,N_5477,N_5531);
or U5685 (N_5685,N_5510,N_5588);
nand U5686 (N_5686,N_5441,N_5586);
nand U5687 (N_5687,N_5479,N_5518);
or U5688 (N_5688,N_5462,N_5434);
nor U5689 (N_5689,N_5486,N_5584);
nor U5690 (N_5690,N_5404,N_5591);
xor U5691 (N_5691,N_5452,N_5511);
and U5692 (N_5692,N_5533,N_5405);
nor U5693 (N_5693,N_5471,N_5454);
nand U5694 (N_5694,N_5517,N_5561);
nand U5695 (N_5695,N_5535,N_5463);
nand U5696 (N_5696,N_5415,N_5590);
nand U5697 (N_5697,N_5476,N_5522);
nand U5698 (N_5698,N_5453,N_5483);
and U5699 (N_5699,N_5473,N_5581);
or U5700 (N_5700,N_5599,N_5404);
and U5701 (N_5701,N_5548,N_5462);
nor U5702 (N_5702,N_5516,N_5565);
and U5703 (N_5703,N_5490,N_5574);
xnor U5704 (N_5704,N_5504,N_5494);
nand U5705 (N_5705,N_5462,N_5508);
nand U5706 (N_5706,N_5534,N_5574);
nor U5707 (N_5707,N_5597,N_5451);
nor U5708 (N_5708,N_5493,N_5575);
nand U5709 (N_5709,N_5551,N_5486);
nand U5710 (N_5710,N_5458,N_5448);
or U5711 (N_5711,N_5450,N_5545);
nand U5712 (N_5712,N_5431,N_5458);
and U5713 (N_5713,N_5433,N_5474);
and U5714 (N_5714,N_5430,N_5464);
or U5715 (N_5715,N_5553,N_5539);
and U5716 (N_5716,N_5509,N_5556);
nand U5717 (N_5717,N_5598,N_5465);
or U5718 (N_5718,N_5452,N_5550);
nand U5719 (N_5719,N_5420,N_5592);
and U5720 (N_5720,N_5490,N_5502);
and U5721 (N_5721,N_5438,N_5474);
or U5722 (N_5722,N_5544,N_5447);
nand U5723 (N_5723,N_5534,N_5437);
nand U5724 (N_5724,N_5419,N_5554);
and U5725 (N_5725,N_5559,N_5499);
and U5726 (N_5726,N_5552,N_5491);
nor U5727 (N_5727,N_5506,N_5570);
nand U5728 (N_5728,N_5447,N_5480);
or U5729 (N_5729,N_5594,N_5446);
and U5730 (N_5730,N_5425,N_5457);
nand U5731 (N_5731,N_5436,N_5428);
nor U5732 (N_5732,N_5471,N_5486);
and U5733 (N_5733,N_5590,N_5416);
nor U5734 (N_5734,N_5554,N_5540);
or U5735 (N_5735,N_5597,N_5446);
or U5736 (N_5736,N_5509,N_5409);
nor U5737 (N_5737,N_5534,N_5440);
and U5738 (N_5738,N_5429,N_5431);
nor U5739 (N_5739,N_5451,N_5486);
nand U5740 (N_5740,N_5425,N_5582);
or U5741 (N_5741,N_5468,N_5530);
or U5742 (N_5742,N_5467,N_5440);
nor U5743 (N_5743,N_5533,N_5560);
or U5744 (N_5744,N_5541,N_5562);
or U5745 (N_5745,N_5503,N_5595);
and U5746 (N_5746,N_5493,N_5450);
nand U5747 (N_5747,N_5502,N_5536);
and U5748 (N_5748,N_5460,N_5572);
and U5749 (N_5749,N_5581,N_5481);
or U5750 (N_5750,N_5441,N_5439);
nand U5751 (N_5751,N_5529,N_5599);
and U5752 (N_5752,N_5580,N_5496);
or U5753 (N_5753,N_5512,N_5508);
nor U5754 (N_5754,N_5411,N_5410);
and U5755 (N_5755,N_5579,N_5560);
and U5756 (N_5756,N_5576,N_5480);
nor U5757 (N_5757,N_5530,N_5508);
and U5758 (N_5758,N_5548,N_5497);
nor U5759 (N_5759,N_5579,N_5409);
nand U5760 (N_5760,N_5523,N_5527);
nand U5761 (N_5761,N_5581,N_5548);
or U5762 (N_5762,N_5447,N_5417);
nor U5763 (N_5763,N_5559,N_5598);
or U5764 (N_5764,N_5590,N_5588);
or U5765 (N_5765,N_5596,N_5521);
nor U5766 (N_5766,N_5480,N_5564);
nor U5767 (N_5767,N_5572,N_5541);
or U5768 (N_5768,N_5534,N_5500);
or U5769 (N_5769,N_5585,N_5592);
and U5770 (N_5770,N_5475,N_5453);
nor U5771 (N_5771,N_5599,N_5510);
nand U5772 (N_5772,N_5427,N_5480);
nand U5773 (N_5773,N_5537,N_5479);
and U5774 (N_5774,N_5547,N_5492);
and U5775 (N_5775,N_5519,N_5479);
or U5776 (N_5776,N_5480,N_5470);
nand U5777 (N_5777,N_5577,N_5538);
xor U5778 (N_5778,N_5445,N_5427);
nand U5779 (N_5779,N_5435,N_5591);
nand U5780 (N_5780,N_5468,N_5544);
nor U5781 (N_5781,N_5480,N_5547);
nand U5782 (N_5782,N_5540,N_5414);
nor U5783 (N_5783,N_5487,N_5594);
or U5784 (N_5784,N_5405,N_5593);
nand U5785 (N_5785,N_5553,N_5410);
nor U5786 (N_5786,N_5458,N_5571);
nor U5787 (N_5787,N_5541,N_5555);
nor U5788 (N_5788,N_5586,N_5455);
and U5789 (N_5789,N_5526,N_5537);
and U5790 (N_5790,N_5588,N_5595);
and U5791 (N_5791,N_5520,N_5524);
nor U5792 (N_5792,N_5431,N_5513);
and U5793 (N_5793,N_5586,N_5421);
nand U5794 (N_5794,N_5560,N_5538);
nand U5795 (N_5795,N_5436,N_5590);
or U5796 (N_5796,N_5436,N_5422);
nor U5797 (N_5797,N_5569,N_5490);
nor U5798 (N_5798,N_5421,N_5437);
nor U5799 (N_5799,N_5578,N_5540);
or U5800 (N_5800,N_5622,N_5782);
xnor U5801 (N_5801,N_5688,N_5733);
nand U5802 (N_5802,N_5713,N_5683);
nor U5803 (N_5803,N_5632,N_5728);
nand U5804 (N_5804,N_5630,N_5675);
nand U5805 (N_5805,N_5697,N_5642);
and U5806 (N_5806,N_5605,N_5665);
and U5807 (N_5807,N_5792,N_5742);
or U5808 (N_5808,N_5727,N_5763);
nor U5809 (N_5809,N_5799,N_5724);
nand U5810 (N_5810,N_5721,N_5648);
nor U5811 (N_5811,N_5612,N_5714);
xnor U5812 (N_5812,N_5786,N_5718);
nand U5813 (N_5813,N_5678,N_5762);
nor U5814 (N_5814,N_5626,N_5754);
nor U5815 (N_5815,N_5680,N_5664);
nand U5816 (N_5816,N_5766,N_5757);
and U5817 (N_5817,N_5602,N_5738);
or U5818 (N_5818,N_5791,N_5734);
and U5819 (N_5819,N_5620,N_5679);
nor U5820 (N_5820,N_5759,N_5789);
nand U5821 (N_5821,N_5649,N_5768);
nor U5822 (N_5822,N_5629,N_5627);
nor U5823 (N_5823,N_5659,N_5623);
nor U5824 (N_5824,N_5691,N_5703);
xor U5825 (N_5825,N_5638,N_5744);
nand U5826 (N_5826,N_5600,N_5695);
and U5827 (N_5827,N_5779,N_5621);
nor U5828 (N_5828,N_5652,N_5616);
or U5829 (N_5829,N_5707,N_5774);
nor U5830 (N_5830,N_5756,N_5755);
or U5831 (N_5831,N_5693,N_5641);
xnor U5832 (N_5832,N_5773,N_5715);
and U5833 (N_5833,N_5797,N_5671);
or U5834 (N_5834,N_5706,N_5781);
nand U5835 (N_5835,N_5711,N_5637);
and U5836 (N_5836,N_5702,N_5661);
or U5837 (N_5837,N_5751,N_5731);
nor U5838 (N_5838,N_5723,N_5761);
and U5839 (N_5839,N_5758,N_5760);
nor U5840 (N_5840,N_5701,N_5793);
and U5841 (N_5841,N_5689,N_5677);
nand U5842 (N_5842,N_5694,N_5698);
nand U5843 (N_5843,N_5670,N_5708);
nand U5844 (N_5844,N_5798,N_5609);
or U5845 (N_5845,N_5608,N_5726);
nand U5846 (N_5846,N_5739,N_5692);
nand U5847 (N_5847,N_5636,N_5699);
and U5848 (N_5848,N_5681,N_5788);
nand U5849 (N_5849,N_5777,N_5633);
and U5850 (N_5850,N_5717,N_5783);
or U5851 (N_5851,N_5647,N_5666);
nand U5852 (N_5852,N_5617,N_5684);
nor U5853 (N_5853,N_5639,N_5750);
and U5854 (N_5854,N_5732,N_5624);
and U5855 (N_5855,N_5690,N_5651);
and U5856 (N_5856,N_5614,N_5601);
nor U5857 (N_5857,N_5610,N_5685);
or U5858 (N_5858,N_5730,N_5737);
or U5859 (N_5859,N_5700,N_5769);
nand U5860 (N_5860,N_5729,N_5663);
nand U5861 (N_5861,N_5645,N_5676);
nand U5862 (N_5862,N_5775,N_5667);
nor U5863 (N_5863,N_5720,N_5710);
xor U5864 (N_5864,N_5765,N_5650);
and U5865 (N_5865,N_5719,N_5696);
nor U5866 (N_5866,N_5795,N_5785);
and U5867 (N_5867,N_5716,N_5686);
and U5868 (N_5868,N_5625,N_5736);
or U5869 (N_5869,N_5776,N_5687);
nand U5870 (N_5870,N_5749,N_5669);
or U5871 (N_5871,N_5655,N_5606);
nand U5872 (N_5872,N_5604,N_5635);
xor U5873 (N_5873,N_5787,N_5628);
or U5874 (N_5874,N_5796,N_5725);
and U5875 (N_5875,N_5780,N_5662);
nor U5876 (N_5876,N_5657,N_5673);
and U5877 (N_5877,N_5741,N_5654);
xor U5878 (N_5878,N_5653,N_5640);
and U5879 (N_5879,N_5752,N_5722);
nand U5880 (N_5880,N_5634,N_5770);
nand U5881 (N_5881,N_5613,N_5656);
nand U5882 (N_5882,N_5631,N_5607);
nor U5883 (N_5883,N_5746,N_5764);
or U5884 (N_5884,N_5740,N_5619);
nor U5885 (N_5885,N_5643,N_5747);
or U5886 (N_5886,N_5618,N_5658);
nand U5887 (N_5887,N_5794,N_5735);
or U5888 (N_5888,N_5767,N_5778);
nand U5889 (N_5889,N_5611,N_5745);
nor U5890 (N_5890,N_5712,N_5705);
and U5891 (N_5891,N_5771,N_5668);
and U5892 (N_5892,N_5603,N_5646);
nor U5893 (N_5893,N_5709,N_5672);
or U5894 (N_5894,N_5772,N_5743);
nor U5895 (N_5895,N_5748,N_5704);
or U5896 (N_5896,N_5644,N_5615);
nand U5897 (N_5897,N_5674,N_5682);
nor U5898 (N_5898,N_5790,N_5784);
nand U5899 (N_5899,N_5660,N_5753);
nor U5900 (N_5900,N_5665,N_5709);
nand U5901 (N_5901,N_5686,N_5667);
nand U5902 (N_5902,N_5674,N_5798);
nand U5903 (N_5903,N_5757,N_5718);
or U5904 (N_5904,N_5600,N_5786);
and U5905 (N_5905,N_5722,N_5647);
or U5906 (N_5906,N_5614,N_5773);
and U5907 (N_5907,N_5623,N_5739);
or U5908 (N_5908,N_5681,N_5728);
or U5909 (N_5909,N_5623,N_5612);
or U5910 (N_5910,N_5775,N_5717);
or U5911 (N_5911,N_5794,N_5655);
nor U5912 (N_5912,N_5631,N_5625);
nor U5913 (N_5913,N_5720,N_5769);
nand U5914 (N_5914,N_5788,N_5652);
nand U5915 (N_5915,N_5602,N_5734);
or U5916 (N_5916,N_5758,N_5741);
and U5917 (N_5917,N_5634,N_5749);
and U5918 (N_5918,N_5783,N_5684);
and U5919 (N_5919,N_5734,N_5698);
and U5920 (N_5920,N_5697,N_5795);
nor U5921 (N_5921,N_5786,N_5792);
and U5922 (N_5922,N_5647,N_5640);
nor U5923 (N_5923,N_5761,N_5634);
nand U5924 (N_5924,N_5665,N_5608);
nor U5925 (N_5925,N_5638,N_5737);
nor U5926 (N_5926,N_5628,N_5691);
nand U5927 (N_5927,N_5741,N_5607);
nor U5928 (N_5928,N_5731,N_5636);
and U5929 (N_5929,N_5785,N_5697);
and U5930 (N_5930,N_5790,N_5694);
nand U5931 (N_5931,N_5697,N_5699);
nand U5932 (N_5932,N_5665,N_5657);
xor U5933 (N_5933,N_5762,N_5732);
nor U5934 (N_5934,N_5799,N_5641);
xnor U5935 (N_5935,N_5622,N_5672);
nor U5936 (N_5936,N_5714,N_5716);
and U5937 (N_5937,N_5621,N_5626);
or U5938 (N_5938,N_5640,N_5787);
or U5939 (N_5939,N_5638,N_5732);
nand U5940 (N_5940,N_5627,N_5602);
or U5941 (N_5941,N_5688,N_5600);
and U5942 (N_5942,N_5726,N_5660);
nand U5943 (N_5943,N_5778,N_5757);
nand U5944 (N_5944,N_5635,N_5625);
nor U5945 (N_5945,N_5705,N_5716);
and U5946 (N_5946,N_5743,N_5699);
or U5947 (N_5947,N_5681,N_5640);
nand U5948 (N_5948,N_5684,N_5755);
and U5949 (N_5949,N_5618,N_5746);
nand U5950 (N_5950,N_5785,N_5600);
or U5951 (N_5951,N_5765,N_5602);
nor U5952 (N_5952,N_5750,N_5619);
nand U5953 (N_5953,N_5619,N_5617);
nor U5954 (N_5954,N_5614,N_5629);
or U5955 (N_5955,N_5777,N_5617);
nor U5956 (N_5956,N_5665,N_5766);
nor U5957 (N_5957,N_5618,N_5694);
and U5958 (N_5958,N_5647,N_5682);
or U5959 (N_5959,N_5793,N_5639);
and U5960 (N_5960,N_5605,N_5668);
or U5961 (N_5961,N_5603,N_5709);
nand U5962 (N_5962,N_5698,N_5711);
nand U5963 (N_5963,N_5767,N_5692);
nor U5964 (N_5964,N_5623,N_5692);
and U5965 (N_5965,N_5691,N_5756);
nand U5966 (N_5966,N_5651,N_5755);
nand U5967 (N_5967,N_5753,N_5665);
and U5968 (N_5968,N_5731,N_5770);
nand U5969 (N_5969,N_5758,N_5789);
or U5970 (N_5970,N_5672,N_5678);
or U5971 (N_5971,N_5763,N_5795);
nand U5972 (N_5972,N_5652,N_5711);
and U5973 (N_5973,N_5622,N_5699);
or U5974 (N_5974,N_5672,N_5671);
or U5975 (N_5975,N_5775,N_5701);
and U5976 (N_5976,N_5798,N_5770);
nand U5977 (N_5977,N_5659,N_5772);
nand U5978 (N_5978,N_5610,N_5715);
nand U5979 (N_5979,N_5731,N_5792);
nor U5980 (N_5980,N_5689,N_5675);
or U5981 (N_5981,N_5656,N_5649);
or U5982 (N_5982,N_5678,N_5625);
and U5983 (N_5983,N_5750,N_5613);
and U5984 (N_5984,N_5740,N_5654);
and U5985 (N_5985,N_5659,N_5675);
nand U5986 (N_5986,N_5738,N_5679);
and U5987 (N_5987,N_5655,N_5704);
and U5988 (N_5988,N_5733,N_5631);
and U5989 (N_5989,N_5765,N_5622);
nor U5990 (N_5990,N_5685,N_5677);
or U5991 (N_5991,N_5725,N_5761);
or U5992 (N_5992,N_5717,N_5781);
or U5993 (N_5993,N_5698,N_5684);
nor U5994 (N_5994,N_5709,N_5777);
or U5995 (N_5995,N_5667,N_5798);
or U5996 (N_5996,N_5678,N_5657);
nor U5997 (N_5997,N_5739,N_5604);
nand U5998 (N_5998,N_5798,N_5735);
nand U5999 (N_5999,N_5778,N_5746);
nor U6000 (N_6000,N_5997,N_5946);
nand U6001 (N_6001,N_5921,N_5964);
or U6002 (N_6002,N_5934,N_5912);
nor U6003 (N_6003,N_5988,N_5808);
and U6004 (N_6004,N_5917,N_5911);
nand U6005 (N_6005,N_5959,N_5857);
nand U6006 (N_6006,N_5851,N_5909);
and U6007 (N_6007,N_5989,N_5858);
and U6008 (N_6008,N_5927,N_5925);
or U6009 (N_6009,N_5854,N_5915);
nand U6010 (N_6010,N_5806,N_5816);
nand U6011 (N_6011,N_5969,N_5938);
and U6012 (N_6012,N_5833,N_5812);
nor U6013 (N_6013,N_5862,N_5880);
nand U6014 (N_6014,N_5865,N_5918);
or U6015 (N_6015,N_5931,N_5847);
nor U6016 (N_6016,N_5957,N_5962);
and U6017 (N_6017,N_5945,N_5978);
nor U6018 (N_6018,N_5944,N_5943);
nand U6019 (N_6019,N_5876,N_5924);
and U6020 (N_6020,N_5904,N_5848);
or U6021 (N_6021,N_5830,N_5856);
and U6022 (N_6022,N_5899,N_5984);
or U6023 (N_6023,N_5834,N_5886);
nand U6024 (N_6024,N_5933,N_5855);
nor U6025 (N_6025,N_5824,N_5804);
or U6026 (N_6026,N_5879,N_5845);
nor U6027 (N_6027,N_5956,N_5983);
or U6028 (N_6028,N_5942,N_5908);
nand U6029 (N_6029,N_5872,N_5822);
nand U6030 (N_6030,N_5894,N_5941);
nand U6031 (N_6031,N_5892,N_5844);
nand U6032 (N_6032,N_5860,N_5999);
nor U6033 (N_6033,N_5825,N_5937);
nand U6034 (N_6034,N_5966,N_5866);
nand U6035 (N_6035,N_5967,N_5981);
or U6036 (N_6036,N_5930,N_5965);
nor U6037 (N_6037,N_5987,N_5963);
nand U6038 (N_6038,N_5839,N_5869);
nor U6039 (N_6039,N_5852,N_5803);
nand U6040 (N_6040,N_5827,N_5843);
nand U6041 (N_6041,N_5875,N_5979);
nor U6042 (N_6042,N_5920,N_5951);
nand U6043 (N_6043,N_5829,N_5800);
and U6044 (N_6044,N_5961,N_5823);
and U6045 (N_6045,N_5995,N_5874);
and U6046 (N_6046,N_5914,N_5998);
xor U6047 (N_6047,N_5952,N_5840);
nand U6048 (N_6048,N_5835,N_5992);
nand U6049 (N_6049,N_5898,N_5900);
and U6050 (N_6050,N_5841,N_5850);
nor U6051 (N_6051,N_5871,N_5985);
and U6052 (N_6052,N_5974,N_5810);
and U6053 (N_6053,N_5991,N_5838);
or U6054 (N_6054,N_5814,N_5884);
nor U6055 (N_6055,N_5919,N_5815);
and U6056 (N_6056,N_5958,N_5955);
nor U6057 (N_6057,N_5973,N_5867);
and U6058 (N_6058,N_5878,N_5832);
or U6059 (N_6059,N_5972,N_5936);
nand U6060 (N_6060,N_5913,N_5820);
or U6061 (N_6061,N_5889,N_5895);
nor U6062 (N_6062,N_5885,N_5968);
and U6063 (N_6063,N_5916,N_5928);
nand U6064 (N_6064,N_5935,N_5923);
and U6065 (N_6065,N_5994,N_5986);
or U6066 (N_6066,N_5993,N_5891);
and U6067 (N_6067,N_5883,N_5818);
nor U6068 (N_6068,N_5950,N_5905);
nor U6069 (N_6069,N_5887,N_5870);
nor U6070 (N_6070,N_5976,N_5888);
nand U6071 (N_6071,N_5811,N_5805);
and U6072 (N_6072,N_5849,N_5902);
or U6073 (N_6073,N_5975,N_5901);
nand U6074 (N_6074,N_5907,N_5807);
and U6075 (N_6075,N_5890,N_5922);
nand U6076 (N_6076,N_5877,N_5868);
and U6077 (N_6077,N_5864,N_5881);
nand U6078 (N_6078,N_5947,N_5990);
or U6079 (N_6079,N_5906,N_5903);
nand U6080 (N_6080,N_5982,N_5837);
xnor U6081 (N_6081,N_5897,N_5926);
nand U6082 (N_6082,N_5939,N_5859);
nor U6083 (N_6083,N_5846,N_5802);
nor U6084 (N_6084,N_5960,N_5861);
nand U6085 (N_6085,N_5970,N_5817);
nand U6086 (N_6086,N_5896,N_5971);
nand U6087 (N_6087,N_5953,N_5948);
nand U6088 (N_6088,N_5863,N_5929);
or U6089 (N_6089,N_5821,N_5932);
nand U6090 (N_6090,N_5910,N_5954);
nor U6091 (N_6091,N_5949,N_5826);
nand U6092 (N_6092,N_5873,N_5801);
or U6093 (N_6093,N_5842,N_5980);
nand U6094 (N_6094,N_5809,N_5819);
or U6095 (N_6095,N_5813,N_5940);
and U6096 (N_6096,N_5977,N_5853);
xnor U6097 (N_6097,N_5882,N_5836);
and U6098 (N_6098,N_5831,N_5828);
or U6099 (N_6099,N_5893,N_5996);
or U6100 (N_6100,N_5866,N_5997);
nor U6101 (N_6101,N_5892,N_5929);
or U6102 (N_6102,N_5993,N_5925);
or U6103 (N_6103,N_5889,N_5960);
or U6104 (N_6104,N_5946,N_5977);
and U6105 (N_6105,N_5813,N_5963);
nand U6106 (N_6106,N_5983,N_5980);
nor U6107 (N_6107,N_5901,N_5978);
or U6108 (N_6108,N_5811,N_5953);
or U6109 (N_6109,N_5815,N_5863);
or U6110 (N_6110,N_5916,N_5805);
nor U6111 (N_6111,N_5846,N_5867);
nand U6112 (N_6112,N_5945,N_5987);
nand U6113 (N_6113,N_5873,N_5971);
nand U6114 (N_6114,N_5918,N_5829);
nor U6115 (N_6115,N_5903,N_5966);
nand U6116 (N_6116,N_5812,N_5830);
and U6117 (N_6117,N_5850,N_5977);
and U6118 (N_6118,N_5867,N_5812);
nor U6119 (N_6119,N_5865,N_5916);
or U6120 (N_6120,N_5898,N_5963);
nor U6121 (N_6121,N_5836,N_5806);
nand U6122 (N_6122,N_5970,N_5814);
and U6123 (N_6123,N_5979,N_5824);
and U6124 (N_6124,N_5890,N_5894);
or U6125 (N_6125,N_5995,N_5870);
nor U6126 (N_6126,N_5883,N_5800);
or U6127 (N_6127,N_5800,N_5890);
or U6128 (N_6128,N_5956,N_5835);
nor U6129 (N_6129,N_5867,N_5830);
nand U6130 (N_6130,N_5866,N_5806);
nand U6131 (N_6131,N_5972,N_5833);
nand U6132 (N_6132,N_5821,N_5843);
nor U6133 (N_6133,N_5940,N_5951);
and U6134 (N_6134,N_5863,N_5831);
nor U6135 (N_6135,N_5980,N_5984);
and U6136 (N_6136,N_5908,N_5897);
or U6137 (N_6137,N_5916,N_5919);
nor U6138 (N_6138,N_5909,N_5817);
and U6139 (N_6139,N_5882,N_5883);
and U6140 (N_6140,N_5818,N_5966);
nor U6141 (N_6141,N_5809,N_5900);
nor U6142 (N_6142,N_5997,N_5896);
and U6143 (N_6143,N_5849,N_5938);
or U6144 (N_6144,N_5913,N_5918);
and U6145 (N_6145,N_5881,N_5873);
nand U6146 (N_6146,N_5903,N_5953);
or U6147 (N_6147,N_5804,N_5882);
and U6148 (N_6148,N_5844,N_5866);
nand U6149 (N_6149,N_5812,N_5906);
or U6150 (N_6150,N_5871,N_5975);
or U6151 (N_6151,N_5832,N_5921);
and U6152 (N_6152,N_5956,N_5942);
nand U6153 (N_6153,N_5995,N_5999);
nor U6154 (N_6154,N_5979,N_5841);
or U6155 (N_6155,N_5877,N_5963);
or U6156 (N_6156,N_5887,N_5865);
nand U6157 (N_6157,N_5833,N_5805);
and U6158 (N_6158,N_5888,N_5929);
or U6159 (N_6159,N_5999,N_5866);
nand U6160 (N_6160,N_5883,N_5935);
xnor U6161 (N_6161,N_5967,N_5914);
and U6162 (N_6162,N_5900,N_5974);
or U6163 (N_6163,N_5959,N_5926);
nand U6164 (N_6164,N_5936,N_5818);
or U6165 (N_6165,N_5960,N_5948);
and U6166 (N_6166,N_5889,N_5806);
xnor U6167 (N_6167,N_5872,N_5846);
or U6168 (N_6168,N_5944,N_5903);
nand U6169 (N_6169,N_5892,N_5807);
nand U6170 (N_6170,N_5907,N_5806);
nand U6171 (N_6171,N_5884,N_5992);
and U6172 (N_6172,N_5841,N_5821);
or U6173 (N_6173,N_5949,N_5905);
and U6174 (N_6174,N_5864,N_5854);
nand U6175 (N_6175,N_5915,N_5880);
nand U6176 (N_6176,N_5947,N_5955);
or U6177 (N_6177,N_5839,N_5924);
nand U6178 (N_6178,N_5818,N_5902);
nand U6179 (N_6179,N_5901,N_5878);
nor U6180 (N_6180,N_5821,N_5969);
and U6181 (N_6181,N_5998,N_5836);
nor U6182 (N_6182,N_5847,N_5869);
nor U6183 (N_6183,N_5870,N_5980);
or U6184 (N_6184,N_5916,N_5939);
and U6185 (N_6185,N_5920,N_5861);
or U6186 (N_6186,N_5858,N_5846);
nor U6187 (N_6187,N_5907,N_5853);
or U6188 (N_6188,N_5893,N_5828);
and U6189 (N_6189,N_5973,N_5935);
nand U6190 (N_6190,N_5959,N_5953);
nand U6191 (N_6191,N_5960,N_5857);
nand U6192 (N_6192,N_5908,N_5825);
nor U6193 (N_6193,N_5836,N_5813);
or U6194 (N_6194,N_5915,N_5851);
nor U6195 (N_6195,N_5954,N_5878);
or U6196 (N_6196,N_5973,N_5891);
nand U6197 (N_6197,N_5921,N_5817);
and U6198 (N_6198,N_5942,N_5945);
xor U6199 (N_6199,N_5918,N_5808);
or U6200 (N_6200,N_6084,N_6028);
nand U6201 (N_6201,N_6102,N_6038);
and U6202 (N_6202,N_6106,N_6189);
and U6203 (N_6203,N_6041,N_6197);
and U6204 (N_6204,N_6082,N_6026);
and U6205 (N_6205,N_6121,N_6117);
or U6206 (N_6206,N_6134,N_6186);
or U6207 (N_6207,N_6176,N_6099);
and U6208 (N_6208,N_6172,N_6014);
nand U6209 (N_6209,N_6073,N_6114);
and U6210 (N_6210,N_6013,N_6067);
xnor U6211 (N_6211,N_6177,N_6005);
nor U6212 (N_6212,N_6079,N_6065);
nand U6213 (N_6213,N_6062,N_6123);
or U6214 (N_6214,N_6180,N_6188);
nor U6215 (N_6215,N_6154,N_6072);
and U6216 (N_6216,N_6133,N_6167);
nor U6217 (N_6217,N_6051,N_6126);
or U6218 (N_6218,N_6173,N_6150);
nor U6219 (N_6219,N_6064,N_6088);
nand U6220 (N_6220,N_6178,N_6031);
or U6221 (N_6221,N_6128,N_6116);
nand U6222 (N_6222,N_6037,N_6164);
or U6223 (N_6223,N_6085,N_6015);
or U6224 (N_6224,N_6021,N_6017);
and U6225 (N_6225,N_6045,N_6080);
nor U6226 (N_6226,N_6066,N_6138);
and U6227 (N_6227,N_6100,N_6061);
nand U6228 (N_6228,N_6153,N_6070);
and U6229 (N_6229,N_6196,N_6192);
or U6230 (N_6230,N_6105,N_6027);
nand U6231 (N_6231,N_6130,N_6009);
and U6232 (N_6232,N_6019,N_6174);
nor U6233 (N_6233,N_6094,N_6023);
nand U6234 (N_6234,N_6093,N_6199);
nand U6235 (N_6235,N_6122,N_6056);
nor U6236 (N_6236,N_6004,N_6043);
and U6237 (N_6237,N_6125,N_6077);
nand U6238 (N_6238,N_6163,N_6159);
and U6239 (N_6239,N_6185,N_6120);
or U6240 (N_6240,N_6146,N_6068);
nor U6241 (N_6241,N_6181,N_6198);
and U6242 (N_6242,N_6143,N_6193);
nand U6243 (N_6243,N_6040,N_6145);
nor U6244 (N_6244,N_6109,N_6044);
or U6245 (N_6245,N_6124,N_6054);
nand U6246 (N_6246,N_6097,N_6098);
nand U6247 (N_6247,N_6058,N_6155);
or U6248 (N_6248,N_6086,N_6162);
and U6249 (N_6249,N_6057,N_6137);
nor U6250 (N_6250,N_6144,N_6152);
nor U6251 (N_6251,N_6111,N_6053);
nor U6252 (N_6252,N_6024,N_6087);
and U6253 (N_6253,N_6049,N_6119);
nor U6254 (N_6254,N_6129,N_6112);
or U6255 (N_6255,N_6032,N_6052);
nand U6256 (N_6256,N_6139,N_6131);
nor U6257 (N_6257,N_6010,N_6000);
or U6258 (N_6258,N_6107,N_6029);
or U6259 (N_6259,N_6089,N_6101);
and U6260 (N_6260,N_6169,N_6011);
or U6261 (N_6261,N_6184,N_6060);
nand U6262 (N_6262,N_6103,N_6132);
nand U6263 (N_6263,N_6118,N_6115);
or U6264 (N_6264,N_6050,N_6074);
nand U6265 (N_6265,N_6147,N_6047);
nand U6266 (N_6266,N_6016,N_6075);
nor U6267 (N_6267,N_6170,N_6025);
nand U6268 (N_6268,N_6001,N_6059);
and U6269 (N_6269,N_6175,N_6194);
or U6270 (N_6270,N_6160,N_6113);
nand U6271 (N_6271,N_6149,N_6063);
or U6272 (N_6272,N_6012,N_6158);
and U6273 (N_6273,N_6151,N_6156);
and U6274 (N_6274,N_6161,N_6090);
xor U6275 (N_6275,N_6092,N_6195);
and U6276 (N_6276,N_6165,N_6078);
nor U6277 (N_6277,N_6018,N_6104);
nor U6278 (N_6278,N_6187,N_6039);
nand U6279 (N_6279,N_6071,N_6081);
and U6280 (N_6280,N_6135,N_6191);
and U6281 (N_6281,N_6036,N_6055);
or U6282 (N_6282,N_6141,N_6003);
nand U6283 (N_6283,N_6006,N_6127);
or U6284 (N_6284,N_6048,N_6034);
and U6285 (N_6285,N_6030,N_6110);
nor U6286 (N_6286,N_6033,N_6171);
and U6287 (N_6287,N_6076,N_6002);
or U6288 (N_6288,N_6108,N_6069);
and U6289 (N_6289,N_6142,N_6020);
nand U6290 (N_6290,N_6140,N_6148);
and U6291 (N_6291,N_6035,N_6091);
nand U6292 (N_6292,N_6083,N_6007);
and U6293 (N_6293,N_6182,N_6042);
nand U6294 (N_6294,N_6190,N_6183);
and U6295 (N_6295,N_6166,N_6046);
nand U6296 (N_6296,N_6179,N_6008);
and U6297 (N_6297,N_6095,N_6022);
nor U6298 (N_6298,N_6168,N_6136);
or U6299 (N_6299,N_6157,N_6096);
nor U6300 (N_6300,N_6086,N_6032);
nor U6301 (N_6301,N_6095,N_6159);
and U6302 (N_6302,N_6175,N_6163);
nand U6303 (N_6303,N_6058,N_6037);
nand U6304 (N_6304,N_6010,N_6055);
nor U6305 (N_6305,N_6087,N_6173);
nor U6306 (N_6306,N_6157,N_6005);
nor U6307 (N_6307,N_6116,N_6068);
and U6308 (N_6308,N_6074,N_6075);
and U6309 (N_6309,N_6178,N_6135);
or U6310 (N_6310,N_6063,N_6032);
or U6311 (N_6311,N_6152,N_6169);
nand U6312 (N_6312,N_6076,N_6159);
and U6313 (N_6313,N_6051,N_6076);
nor U6314 (N_6314,N_6135,N_6157);
nand U6315 (N_6315,N_6129,N_6051);
or U6316 (N_6316,N_6021,N_6117);
and U6317 (N_6317,N_6073,N_6184);
nor U6318 (N_6318,N_6138,N_6171);
or U6319 (N_6319,N_6069,N_6083);
nand U6320 (N_6320,N_6064,N_6098);
nor U6321 (N_6321,N_6071,N_6099);
nand U6322 (N_6322,N_6069,N_6028);
or U6323 (N_6323,N_6075,N_6026);
and U6324 (N_6324,N_6139,N_6047);
or U6325 (N_6325,N_6118,N_6056);
or U6326 (N_6326,N_6183,N_6004);
and U6327 (N_6327,N_6189,N_6005);
or U6328 (N_6328,N_6076,N_6047);
nor U6329 (N_6329,N_6152,N_6093);
and U6330 (N_6330,N_6152,N_6080);
nand U6331 (N_6331,N_6196,N_6193);
nand U6332 (N_6332,N_6067,N_6022);
nor U6333 (N_6333,N_6012,N_6011);
and U6334 (N_6334,N_6113,N_6039);
nor U6335 (N_6335,N_6131,N_6123);
nand U6336 (N_6336,N_6140,N_6003);
and U6337 (N_6337,N_6026,N_6146);
and U6338 (N_6338,N_6022,N_6125);
and U6339 (N_6339,N_6144,N_6077);
or U6340 (N_6340,N_6170,N_6112);
nand U6341 (N_6341,N_6087,N_6153);
and U6342 (N_6342,N_6083,N_6065);
nand U6343 (N_6343,N_6012,N_6024);
or U6344 (N_6344,N_6131,N_6067);
and U6345 (N_6345,N_6098,N_6090);
nor U6346 (N_6346,N_6039,N_6117);
nor U6347 (N_6347,N_6081,N_6135);
and U6348 (N_6348,N_6023,N_6117);
and U6349 (N_6349,N_6079,N_6036);
nand U6350 (N_6350,N_6159,N_6148);
nor U6351 (N_6351,N_6041,N_6175);
nor U6352 (N_6352,N_6053,N_6017);
or U6353 (N_6353,N_6050,N_6192);
nand U6354 (N_6354,N_6150,N_6080);
nor U6355 (N_6355,N_6053,N_6130);
nor U6356 (N_6356,N_6124,N_6103);
and U6357 (N_6357,N_6166,N_6040);
nor U6358 (N_6358,N_6186,N_6093);
and U6359 (N_6359,N_6180,N_6051);
and U6360 (N_6360,N_6085,N_6168);
or U6361 (N_6361,N_6069,N_6045);
nand U6362 (N_6362,N_6098,N_6062);
nand U6363 (N_6363,N_6101,N_6126);
nand U6364 (N_6364,N_6047,N_6079);
nor U6365 (N_6365,N_6055,N_6133);
and U6366 (N_6366,N_6039,N_6150);
nand U6367 (N_6367,N_6017,N_6046);
nand U6368 (N_6368,N_6192,N_6060);
nor U6369 (N_6369,N_6055,N_6074);
and U6370 (N_6370,N_6194,N_6055);
nand U6371 (N_6371,N_6170,N_6031);
or U6372 (N_6372,N_6169,N_6123);
nand U6373 (N_6373,N_6147,N_6040);
nor U6374 (N_6374,N_6131,N_6081);
or U6375 (N_6375,N_6046,N_6073);
or U6376 (N_6376,N_6125,N_6089);
nand U6377 (N_6377,N_6176,N_6001);
nor U6378 (N_6378,N_6151,N_6084);
or U6379 (N_6379,N_6192,N_6166);
and U6380 (N_6380,N_6124,N_6119);
nand U6381 (N_6381,N_6163,N_6089);
nor U6382 (N_6382,N_6094,N_6099);
and U6383 (N_6383,N_6155,N_6068);
or U6384 (N_6384,N_6157,N_6117);
and U6385 (N_6385,N_6039,N_6180);
nand U6386 (N_6386,N_6194,N_6087);
nor U6387 (N_6387,N_6011,N_6181);
nor U6388 (N_6388,N_6103,N_6059);
nand U6389 (N_6389,N_6129,N_6038);
or U6390 (N_6390,N_6086,N_6193);
or U6391 (N_6391,N_6140,N_6071);
and U6392 (N_6392,N_6039,N_6006);
nand U6393 (N_6393,N_6014,N_6127);
and U6394 (N_6394,N_6006,N_6076);
and U6395 (N_6395,N_6064,N_6061);
nand U6396 (N_6396,N_6146,N_6105);
or U6397 (N_6397,N_6047,N_6098);
and U6398 (N_6398,N_6101,N_6158);
nand U6399 (N_6399,N_6128,N_6080);
and U6400 (N_6400,N_6235,N_6391);
and U6401 (N_6401,N_6254,N_6212);
nor U6402 (N_6402,N_6279,N_6325);
nor U6403 (N_6403,N_6288,N_6220);
or U6404 (N_6404,N_6280,N_6389);
and U6405 (N_6405,N_6277,N_6306);
or U6406 (N_6406,N_6294,N_6244);
or U6407 (N_6407,N_6207,N_6290);
or U6408 (N_6408,N_6315,N_6388);
nor U6409 (N_6409,N_6338,N_6371);
and U6410 (N_6410,N_6268,N_6312);
or U6411 (N_6411,N_6365,N_6247);
or U6412 (N_6412,N_6282,N_6368);
or U6413 (N_6413,N_6314,N_6305);
nor U6414 (N_6414,N_6348,N_6260);
nor U6415 (N_6415,N_6248,N_6399);
nand U6416 (N_6416,N_6356,N_6215);
or U6417 (N_6417,N_6236,N_6275);
or U6418 (N_6418,N_6224,N_6217);
and U6419 (N_6419,N_6310,N_6237);
and U6420 (N_6420,N_6266,N_6343);
nor U6421 (N_6421,N_6295,N_6345);
and U6422 (N_6422,N_6287,N_6360);
nand U6423 (N_6423,N_6228,N_6239);
and U6424 (N_6424,N_6253,N_6396);
nand U6425 (N_6425,N_6202,N_6203);
or U6426 (N_6426,N_6208,N_6200);
and U6427 (N_6427,N_6308,N_6296);
nor U6428 (N_6428,N_6354,N_6326);
nor U6429 (N_6429,N_6241,N_6289);
nand U6430 (N_6430,N_6256,N_6350);
nand U6431 (N_6431,N_6246,N_6209);
nand U6432 (N_6432,N_6329,N_6250);
and U6433 (N_6433,N_6362,N_6379);
or U6434 (N_6434,N_6249,N_6378);
or U6435 (N_6435,N_6347,N_6227);
nor U6436 (N_6436,N_6251,N_6299);
or U6437 (N_6437,N_6377,N_6327);
and U6438 (N_6438,N_6298,N_6303);
and U6439 (N_6439,N_6206,N_6328);
or U6440 (N_6440,N_6267,N_6272);
and U6441 (N_6441,N_6330,N_6386);
and U6442 (N_6442,N_6398,N_6223);
and U6443 (N_6443,N_6342,N_6361);
nand U6444 (N_6444,N_6286,N_6336);
nor U6445 (N_6445,N_6376,N_6240);
or U6446 (N_6446,N_6264,N_6263);
and U6447 (N_6447,N_6331,N_6384);
nor U6448 (N_6448,N_6380,N_6346);
nand U6449 (N_6449,N_6341,N_6243);
nor U6450 (N_6450,N_6344,N_6383);
nand U6451 (N_6451,N_6234,N_6313);
and U6452 (N_6452,N_6218,N_6238);
nor U6453 (N_6453,N_6231,N_6265);
nor U6454 (N_6454,N_6307,N_6381);
nor U6455 (N_6455,N_6309,N_6349);
and U6456 (N_6456,N_6395,N_6353);
nand U6457 (N_6457,N_6359,N_6393);
nor U6458 (N_6458,N_6304,N_6210);
and U6459 (N_6459,N_6257,N_6339);
and U6460 (N_6460,N_6285,N_6358);
nor U6461 (N_6461,N_6318,N_6211);
and U6462 (N_6462,N_6316,N_6333);
nor U6463 (N_6463,N_6352,N_6382);
and U6464 (N_6464,N_6216,N_6252);
or U6465 (N_6465,N_6233,N_6204);
and U6466 (N_6466,N_6320,N_6261);
nand U6467 (N_6467,N_6387,N_6369);
or U6468 (N_6468,N_6372,N_6324);
nor U6469 (N_6469,N_6269,N_6283);
and U6470 (N_6470,N_6334,N_6300);
nor U6471 (N_6471,N_6242,N_6293);
nor U6472 (N_6472,N_6258,N_6375);
or U6473 (N_6473,N_6255,N_6367);
or U6474 (N_6474,N_6276,N_6245);
nand U6475 (N_6475,N_6230,N_6292);
or U6476 (N_6476,N_6273,N_6225);
nor U6477 (N_6477,N_6373,N_6274);
and U6478 (N_6478,N_6229,N_6278);
or U6479 (N_6479,N_6205,N_6394);
or U6480 (N_6480,N_6232,N_6226);
or U6481 (N_6481,N_6337,N_6302);
nor U6482 (N_6482,N_6222,N_6351);
or U6483 (N_6483,N_6291,N_6284);
nand U6484 (N_6484,N_6385,N_6297);
and U6485 (N_6485,N_6213,N_6355);
and U6486 (N_6486,N_6319,N_6332);
and U6487 (N_6487,N_6281,N_6214);
or U6488 (N_6488,N_6357,N_6262);
or U6489 (N_6489,N_6340,N_6363);
nor U6490 (N_6490,N_6370,N_6323);
and U6491 (N_6491,N_6321,N_6201);
nor U6492 (N_6492,N_6271,N_6301);
or U6493 (N_6493,N_6392,N_6366);
xor U6494 (N_6494,N_6219,N_6364);
nand U6495 (N_6495,N_6270,N_6322);
or U6496 (N_6496,N_6390,N_6311);
nor U6497 (N_6497,N_6397,N_6259);
or U6498 (N_6498,N_6317,N_6335);
and U6499 (N_6499,N_6374,N_6221);
or U6500 (N_6500,N_6395,N_6302);
and U6501 (N_6501,N_6288,N_6310);
and U6502 (N_6502,N_6255,N_6228);
and U6503 (N_6503,N_6234,N_6224);
and U6504 (N_6504,N_6275,N_6221);
or U6505 (N_6505,N_6365,N_6315);
or U6506 (N_6506,N_6389,N_6338);
nand U6507 (N_6507,N_6338,N_6300);
nand U6508 (N_6508,N_6307,N_6233);
or U6509 (N_6509,N_6337,N_6328);
nand U6510 (N_6510,N_6262,N_6299);
nor U6511 (N_6511,N_6228,N_6259);
nor U6512 (N_6512,N_6293,N_6379);
nand U6513 (N_6513,N_6351,N_6384);
and U6514 (N_6514,N_6394,N_6387);
nor U6515 (N_6515,N_6259,N_6357);
nand U6516 (N_6516,N_6226,N_6340);
nor U6517 (N_6517,N_6201,N_6310);
or U6518 (N_6518,N_6320,N_6314);
and U6519 (N_6519,N_6255,N_6204);
nor U6520 (N_6520,N_6297,N_6238);
or U6521 (N_6521,N_6260,N_6282);
nand U6522 (N_6522,N_6246,N_6259);
or U6523 (N_6523,N_6376,N_6362);
and U6524 (N_6524,N_6350,N_6261);
nand U6525 (N_6525,N_6367,N_6237);
and U6526 (N_6526,N_6207,N_6353);
or U6527 (N_6527,N_6269,N_6289);
and U6528 (N_6528,N_6286,N_6330);
and U6529 (N_6529,N_6397,N_6378);
and U6530 (N_6530,N_6273,N_6258);
nand U6531 (N_6531,N_6360,N_6357);
nor U6532 (N_6532,N_6247,N_6304);
xnor U6533 (N_6533,N_6314,N_6368);
nand U6534 (N_6534,N_6345,N_6260);
or U6535 (N_6535,N_6286,N_6314);
nor U6536 (N_6536,N_6264,N_6271);
nand U6537 (N_6537,N_6323,N_6385);
and U6538 (N_6538,N_6268,N_6264);
and U6539 (N_6539,N_6313,N_6233);
and U6540 (N_6540,N_6263,N_6277);
nor U6541 (N_6541,N_6361,N_6202);
nand U6542 (N_6542,N_6348,N_6300);
nand U6543 (N_6543,N_6247,N_6370);
or U6544 (N_6544,N_6340,N_6216);
or U6545 (N_6545,N_6204,N_6268);
nor U6546 (N_6546,N_6306,N_6254);
nor U6547 (N_6547,N_6382,N_6347);
nand U6548 (N_6548,N_6325,N_6354);
nand U6549 (N_6549,N_6388,N_6277);
nor U6550 (N_6550,N_6384,N_6275);
or U6551 (N_6551,N_6312,N_6237);
nor U6552 (N_6552,N_6373,N_6310);
xor U6553 (N_6553,N_6280,N_6222);
or U6554 (N_6554,N_6252,N_6203);
or U6555 (N_6555,N_6279,N_6364);
or U6556 (N_6556,N_6375,N_6386);
nand U6557 (N_6557,N_6396,N_6291);
or U6558 (N_6558,N_6349,N_6252);
nand U6559 (N_6559,N_6361,N_6243);
and U6560 (N_6560,N_6278,N_6382);
xnor U6561 (N_6561,N_6203,N_6241);
and U6562 (N_6562,N_6357,N_6385);
or U6563 (N_6563,N_6337,N_6227);
nand U6564 (N_6564,N_6317,N_6203);
nand U6565 (N_6565,N_6210,N_6399);
nor U6566 (N_6566,N_6358,N_6261);
nand U6567 (N_6567,N_6289,N_6319);
or U6568 (N_6568,N_6342,N_6238);
nor U6569 (N_6569,N_6311,N_6244);
and U6570 (N_6570,N_6301,N_6217);
and U6571 (N_6571,N_6275,N_6341);
and U6572 (N_6572,N_6278,N_6257);
nor U6573 (N_6573,N_6281,N_6209);
nand U6574 (N_6574,N_6283,N_6386);
nor U6575 (N_6575,N_6277,N_6207);
and U6576 (N_6576,N_6342,N_6326);
or U6577 (N_6577,N_6352,N_6276);
or U6578 (N_6578,N_6339,N_6335);
nor U6579 (N_6579,N_6210,N_6379);
nand U6580 (N_6580,N_6309,N_6394);
or U6581 (N_6581,N_6346,N_6273);
nand U6582 (N_6582,N_6217,N_6248);
nand U6583 (N_6583,N_6315,N_6326);
nand U6584 (N_6584,N_6296,N_6317);
or U6585 (N_6585,N_6395,N_6360);
and U6586 (N_6586,N_6299,N_6362);
nor U6587 (N_6587,N_6303,N_6365);
nand U6588 (N_6588,N_6309,N_6323);
nor U6589 (N_6589,N_6229,N_6358);
or U6590 (N_6590,N_6378,N_6309);
and U6591 (N_6591,N_6221,N_6300);
nor U6592 (N_6592,N_6367,N_6291);
nor U6593 (N_6593,N_6373,N_6383);
and U6594 (N_6594,N_6350,N_6375);
and U6595 (N_6595,N_6399,N_6326);
nor U6596 (N_6596,N_6254,N_6358);
nand U6597 (N_6597,N_6378,N_6336);
nor U6598 (N_6598,N_6373,N_6351);
nand U6599 (N_6599,N_6202,N_6240);
or U6600 (N_6600,N_6533,N_6495);
nand U6601 (N_6601,N_6576,N_6483);
nor U6602 (N_6602,N_6553,N_6449);
nand U6603 (N_6603,N_6550,N_6418);
and U6604 (N_6604,N_6549,N_6578);
or U6605 (N_6605,N_6513,N_6420);
nor U6606 (N_6606,N_6589,N_6532);
and U6607 (N_6607,N_6481,N_6564);
and U6608 (N_6608,N_6504,N_6594);
nor U6609 (N_6609,N_6508,N_6456);
or U6610 (N_6610,N_6590,N_6591);
or U6611 (N_6611,N_6493,N_6555);
and U6612 (N_6612,N_6429,N_6443);
or U6613 (N_6613,N_6461,N_6574);
and U6614 (N_6614,N_6520,N_6462);
xor U6615 (N_6615,N_6471,N_6492);
and U6616 (N_6616,N_6527,N_6525);
nor U6617 (N_6617,N_6465,N_6595);
or U6618 (N_6618,N_6415,N_6592);
or U6619 (N_6619,N_6522,N_6544);
nand U6620 (N_6620,N_6587,N_6416);
or U6621 (N_6621,N_6430,N_6423);
nor U6622 (N_6622,N_6466,N_6435);
nand U6623 (N_6623,N_6517,N_6477);
and U6624 (N_6624,N_6455,N_6507);
and U6625 (N_6625,N_6486,N_6516);
xor U6626 (N_6626,N_6511,N_6496);
nand U6627 (N_6627,N_6485,N_6400);
and U6628 (N_6628,N_6568,N_6534);
and U6629 (N_6629,N_6518,N_6472);
or U6630 (N_6630,N_6419,N_6433);
nand U6631 (N_6631,N_6512,N_6505);
nand U6632 (N_6632,N_6523,N_6484);
nor U6633 (N_6633,N_6597,N_6598);
or U6634 (N_6634,N_6599,N_6593);
nand U6635 (N_6635,N_6545,N_6404);
and U6636 (N_6636,N_6441,N_6557);
or U6637 (N_6637,N_6442,N_6478);
nand U6638 (N_6638,N_6579,N_6526);
or U6639 (N_6639,N_6431,N_6451);
nand U6640 (N_6640,N_6436,N_6521);
or U6641 (N_6641,N_6541,N_6539);
nand U6642 (N_6642,N_6446,N_6554);
or U6643 (N_6643,N_6454,N_6586);
nor U6644 (N_6644,N_6596,N_6409);
nor U6645 (N_6645,N_6547,N_6585);
xor U6646 (N_6646,N_6438,N_6542);
nand U6647 (N_6647,N_6566,N_6475);
and U6648 (N_6648,N_6506,N_6488);
and U6649 (N_6649,N_6529,N_6405);
nand U6650 (N_6650,N_6588,N_6536);
or U6651 (N_6651,N_6414,N_6417);
nand U6652 (N_6652,N_6551,N_6490);
or U6653 (N_6653,N_6581,N_6489);
and U6654 (N_6654,N_6439,N_6531);
and U6655 (N_6655,N_6561,N_6571);
or U6656 (N_6656,N_6469,N_6464);
and U6657 (N_6657,N_6425,N_6467);
and U6658 (N_6658,N_6444,N_6580);
nand U6659 (N_6659,N_6575,N_6538);
and U6660 (N_6660,N_6565,N_6445);
or U6661 (N_6661,N_6582,N_6501);
xor U6662 (N_6662,N_6573,N_6452);
and U6663 (N_6663,N_6535,N_6577);
nand U6664 (N_6664,N_6470,N_6432);
xor U6665 (N_6665,N_6509,N_6491);
nor U6666 (N_6666,N_6410,N_6412);
nand U6667 (N_6667,N_6437,N_6559);
xor U6668 (N_6668,N_6552,N_6482);
or U6669 (N_6669,N_6560,N_6546);
nor U6670 (N_6670,N_6479,N_6584);
or U6671 (N_6671,N_6558,N_6572);
and U6672 (N_6672,N_6403,N_6460);
or U6673 (N_6673,N_6515,N_6413);
and U6674 (N_6674,N_6426,N_6424);
or U6675 (N_6675,N_6510,N_6458);
nor U6676 (N_6676,N_6450,N_6459);
or U6677 (N_6677,N_6407,N_6463);
nor U6678 (N_6678,N_6570,N_6480);
nand U6679 (N_6679,N_6448,N_6499);
and U6680 (N_6680,N_6447,N_6548);
nor U6681 (N_6681,N_6476,N_6457);
and U6682 (N_6682,N_6567,N_6524);
nand U6683 (N_6683,N_6408,N_6543);
nand U6684 (N_6684,N_6473,N_6434);
and U6685 (N_6685,N_6422,N_6440);
or U6686 (N_6686,N_6402,N_6497);
nand U6687 (N_6687,N_6421,N_6540);
nor U6688 (N_6688,N_6537,N_6474);
nand U6689 (N_6689,N_6528,N_6427);
nand U6690 (N_6690,N_6563,N_6487);
or U6691 (N_6691,N_6494,N_6583);
and U6692 (N_6692,N_6453,N_6514);
or U6693 (N_6693,N_6503,N_6519);
nor U6694 (N_6694,N_6556,N_6530);
xnor U6695 (N_6695,N_6406,N_6401);
or U6696 (N_6696,N_6562,N_6500);
nor U6697 (N_6697,N_6411,N_6569);
and U6698 (N_6698,N_6428,N_6498);
nor U6699 (N_6699,N_6502,N_6468);
or U6700 (N_6700,N_6489,N_6473);
nand U6701 (N_6701,N_6599,N_6462);
or U6702 (N_6702,N_6415,N_6511);
and U6703 (N_6703,N_6451,N_6457);
or U6704 (N_6704,N_6553,N_6405);
nor U6705 (N_6705,N_6552,N_6466);
nor U6706 (N_6706,N_6577,N_6495);
or U6707 (N_6707,N_6454,N_6521);
or U6708 (N_6708,N_6451,N_6561);
nor U6709 (N_6709,N_6447,N_6420);
xnor U6710 (N_6710,N_6587,N_6476);
nor U6711 (N_6711,N_6497,N_6587);
nand U6712 (N_6712,N_6585,N_6557);
and U6713 (N_6713,N_6550,N_6504);
and U6714 (N_6714,N_6540,N_6450);
or U6715 (N_6715,N_6408,N_6456);
and U6716 (N_6716,N_6569,N_6591);
or U6717 (N_6717,N_6597,N_6507);
nor U6718 (N_6718,N_6557,N_6432);
nor U6719 (N_6719,N_6523,N_6421);
nor U6720 (N_6720,N_6469,N_6565);
and U6721 (N_6721,N_6545,N_6524);
nor U6722 (N_6722,N_6467,N_6519);
or U6723 (N_6723,N_6528,N_6508);
nor U6724 (N_6724,N_6520,N_6422);
xor U6725 (N_6725,N_6527,N_6415);
and U6726 (N_6726,N_6574,N_6426);
and U6727 (N_6727,N_6507,N_6427);
nor U6728 (N_6728,N_6523,N_6577);
nor U6729 (N_6729,N_6575,N_6442);
nor U6730 (N_6730,N_6443,N_6550);
or U6731 (N_6731,N_6459,N_6437);
and U6732 (N_6732,N_6542,N_6575);
or U6733 (N_6733,N_6467,N_6584);
nand U6734 (N_6734,N_6530,N_6455);
nand U6735 (N_6735,N_6482,N_6575);
or U6736 (N_6736,N_6496,N_6573);
nand U6737 (N_6737,N_6547,N_6526);
nor U6738 (N_6738,N_6425,N_6570);
or U6739 (N_6739,N_6450,N_6401);
nand U6740 (N_6740,N_6453,N_6545);
and U6741 (N_6741,N_6580,N_6589);
xor U6742 (N_6742,N_6531,N_6579);
nand U6743 (N_6743,N_6539,N_6469);
nand U6744 (N_6744,N_6441,N_6587);
and U6745 (N_6745,N_6440,N_6469);
and U6746 (N_6746,N_6497,N_6405);
and U6747 (N_6747,N_6422,N_6410);
nor U6748 (N_6748,N_6468,N_6437);
nand U6749 (N_6749,N_6410,N_6518);
or U6750 (N_6750,N_6592,N_6526);
or U6751 (N_6751,N_6598,N_6588);
nand U6752 (N_6752,N_6442,N_6472);
nand U6753 (N_6753,N_6403,N_6512);
and U6754 (N_6754,N_6471,N_6486);
nand U6755 (N_6755,N_6496,N_6434);
or U6756 (N_6756,N_6577,N_6554);
xor U6757 (N_6757,N_6533,N_6536);
nand U6758 (N_6758,N_6587,N_6575);
nand U6759 (N_6759,N_6532,N_6525);
and U6760 (N_6760,N_6425,N_6506);
and U6761 (N_6761,N_6594,N_6593);
nor U6762 (N_6762,N_6492,N_6586);
or U6763 (N_6763,N_6414,N_6486);
or U6764 (N_6764,N_6488,N_6483);
nor U6765 (N_6765,N_6596,N_6444);
or U6766 (N_6766,N_6423,N_6583);
and U6767 (N_6767,N_6595,N_6531);
nor U6768 (N_6768,N_6575,N_6479);
nand U6769 (N_6769,N_6487,N_6497);
and U6770 (N_6770,N_6500,N_6485);
or U6771 (N_6771,N_6521,N_6590);
or U6772 (N_6772,N_6463,N_6594);
nor U6773 (N_6773,N_6508,N_6513);
nor U6774 (N_6774,N_6589,N_6517);
or U6775 (N_6775,N_6576,N_6493);
nor U6776 (N_6776,N_6432,N_6563);
nor U6777 (N_6777,N_6577,N_6403);
or U6778 (N_6778,N_6436,N_6466);
and U6779 (N_6779,N_6434,N_6491);
or U6780 (N_6780,N_6470,N_6462);
nor U6781 (N_6781,N_6462,N_6502);
nor U6782 (N_6782,N_6477,N_6556);
or U6783 (N_6783,N_6546,N_6445);
or U6784 (N_6784,N_6417,N_6410);
or U6785 (N_6785,N_6437,N_6594);
or U6786 (N_6786,N_6473,N_6534);
or U6787 (N_6787,N_6592,N_6434);
or U6788 (N_6788,N_6520,N_6527);
nand U6789 (N_6789,N_6528,N_6572);
nor U6790 (N_6790,N_6493,N_6596);
and U6791 (N_6791,N_6562,N_6535);
and U6792 (N_6792,N_6574,N_6439);
and U6793 (N_6793,N_6545,N_6406);
xnor U6794 (N_6794,N_6543,N_6544);
or U6795 (N_6795,N_6590,N_6426);
nand U6796 (N_6796,N_6481,N_6422);
nor U6797 (N_6797,N_6559,N_6469);
or U6798 (N_6798,N_6572,N_6464);
nand U6799 (N_6799,N_6404,N_6419);
nand U6800 (N_6800,N_6674,N_6604);
nand U6801 (N_6801,N_6779,N_6678);
or U6802 (N_6802,N_6616,N_6795);
and U6803 (N_6803,N_6773,N_6609);
nor U6804 (N_6804,N_6691,N_6719);
nand U6805 (N_6805,N_6607,N_6640);
or U6806 (N_6806,N_6781,N_6642);
and U6807 (N_6807,N_6738,N_6655);
and U6808 (N_6808,N_6650,N_6657);
nand U6809 (N_6809,N_6735,N_6628);
or U6810 (N_6810,N_6767,N_6747);
nor U6811 (N_6811,N_6608,N_6643);
or U6812 (N_6812,N_6702,N_6754);
or U6813 (N_6813,N_6682,N_6714);
and U6814 (N_6814,N_6671,N_6644);
nand U6815 (N_6815,N_6633,N_6725);
or U6816 (N_6816,N_6727,N_6761);
nand U6817 (N_6817,N_6606,N_6664);
or U6818 (N_6818,N_6629,N_6651);
or U6819 (N_6819,N_6740,N_6717);
nor U6820 (N_6820,N_6698,N_6718);
or U6821 (N_6821,N_6611,N_6681);
nor U6822 (N_6822,N_6756,N_6675);
and U6823 (N_6823,N_6677,N_6723);
nand U6824 (N_6824,N_6603,N_6771);
and U6825 (N_6825,N_6656,N_6705);
nor U6826 (N_6826,N_6632,N_6613);
nand U6827 (N_6827,N_6748,N_6783);
nand U6828 (N_6828,N_6744,N_6768);
nor U6829 (N_6829,N_6652,N_6786);
or U6830 (N_6830,N_6764,N_6619);
nor U6831 (N_6831,N_6688,N_6792);
nand U6832 (N_6832,N_6679,N_6623);
and U6833 (N_6833,N_6668,N_6708);
and U6834 (N_6834,N_6791,N_6605);
or U6835 (N_6835,N_6710,N_6711);
nor U6836 (N_6836,N_6745,N_6743);
nor U6837 (N_6837,N_6666,N_6704);
and U6838 (N_6838,N_6615,N_6746);
nor U6839 (N_6839,N_6794,N_6799);
and U6840 (N_6840,N_6760,N_6733);
nand U6841 (N_6841,N_6622,N_6726);
xnor U6842 (N_6842,N_6684,N_6777);
and U6843 (N_6843,N_6729,N_6600);
xor U6844 (N_6844,N_6641,N_6776);
nor U6845 (N_6845,N_6690,N_6638);
nand U6846 (N_6846,N_6687,N_6697);
or U6847 (N_6847,N_6713,N_6766);
nor U6848 (N_6848,N_6672,N_6665);
xnor U6849 (N_6849,N_6654,N_6785);
or U6850 (N_6850,N_6648,N_6653);
nand U6851 (N_6851,N_6649,N_6731);
and U6852 (N_6852,N_6676,N_6692);
and U6853 (N_6853,N_6721,N_6750);
or U6854 (N_6854,N_6601,N_6715);
or U6855 (N_6855,N_6757,N_6749);
and U6856 (N_6856,N_6759,N_6752);
nand U6857 (N_6857,N_6620,N_6670);
nand U6858 (N_6858,N_6765,N_6772);
or U6859 (N_6859,N_6784,N_6669);
xor U6860 (N_6860,N_6780,N_6716);
nor U6861 (N_6861,N_6797,N_6667);
nor U6862 (N_6862,N_6755,N_6775);
and U6863 (N_6863,N_6787,N_6617);
and U6864 (N_6864,N_6722,N_6736);
nand U6865 (N_6865,N_6798,N_6614);
or U6866 (N_6866,N_6753,N_6741);
or U6867 (N_6867,N_6730,N_6630);
nand U6868 (N_6868,N_6790,N_6639);
or U6869 (N_6869,N_6636,N_6732);
nor U6870 (N_6870,N_6796,N_6621);
or U6871 (N_6871,N_6680,N_6637);
nor U6872 (N_6872,N_6770,N_6661);
and U6873 (N_6873,N_6686,N_6782);
nand U6874 (N_6874,N_6724,N_6602);
and U6875 (N_6875,N_6699,N_6631);
and U6876 (N_6876,N_6758,N_6788);
nor U6877 (N_6877,N_6703,N_6763);
and U6878 (N_6878,N_6720,N_6694);
and U6879 (N_6879,N_6751,N_6789);
or U6880 (N_6880,N_6627,N_6663);
and U6881 (N_6881,N_6701,N_6625);
nand U6882 (N_6882,N_6769,N_6673);
or U6883 (N_6883,N_6700,N_6618);
nand U6884 (N_6884,N_6707,N_6660);
nor U6885 (N_6885,N_6734,N_6683);
xor U6886 (N_6886,N_6695,N_6709);
nand U6887 (N_6887,N_6728,N_6706);
xnor U6888 (N_6888,N_6737,N_6662);
nor U6889 (N_6889,N_6659,N_6647);
and U6890 (N_6890,N_6774,N_6793);
or U6891 (N_6891,N_6762,N_6646);
and U6892 (N_6892,N_6693,N_6712);
or U6893 (N_6893,N_6685,N_6610);
nand U6894 (N_6894,N_6624,N_6739);
nor U6895 (N_6895,N_6645,N_6612);
nand U6896 (N_6896,N_6626,N_6658);
nand U6897 (N_6897,N_6778,N_6689);
nand U6898 (N_6898,N_6696,N_6634);
nand U6899 (N_6899,N_6742,N_6635);
nand U6900 (N_6900,N_6794,N_6739);
xor U6901 (N_6901,N_6768,N_6799);
and U6902 (N_6902,N_6768,N_6658);
nor U6903 (N_6903,N_6761,N_6700);
and U6904 (N_6904,N_6753,N_6793);
nand U6905 (N_6905,N_6799,N_6636);
or U6906 (N_6906,N_6604,N_6720);
nor U6907 (N_6907,N_6622,N_6793);
nand U6908 (N_6908,N_6759,N_6615);
and U6909 (N_6909,N_6757,N_6619);
nand U6910 (N_6910,N_6668,N_6788);
and U6911 (N_6911,N_6610,N_6602);
nand U6912 (N_6912,N_6626,N_6799);
or U6913 (N_6913,N_6786,N_6720);
nand U6914 (N_6914,N_6777,N_6662);
and U6915 (N_6915,N_6738,N_6695);
and U6916 (N_6916,N_6682,N_6678);
and U6917 (N_6917,N_6738,N_6626);
nor U6918 (N_6918,N_6667,N_6757);
nand U6919 (N_6919,N_6655,N_6675);
nor U6920 (N_6920,N_6624,N_6740);
or U6921 (N_6921,N_6785,N_6673);
nand U6922 (N_6922,N_6736,N_6621);
nor U6923 (N_6923,N_6765,N_6641);
and U6924 (N_6924,N_6790,N_6741);
and U6925 (N_6925,N_6687,N_6758);
nor U6926 (N_6926,N_6711,N_6686);
nand U6927 (N_6927,N_6690,N_6681);
and U6928 (N_6928,N_6626,N_6753);
and U6929 (N_6929,N_6613,N_6617);
or U6930 (N_6930,N_6688,N_6702);
nand U6931 (N_6931,N_6627,N_6631);
nor U6932 (N_6932,N_6668,N_6772);
nor U6933 (N_6933,N_6745,N_6651);
and U6934 (N_6934,N_6648,N_6690);
or U6935 (N_6935,N_6677,N_6646);
or U6936 (N_6936,N_6692,N_6794);
nand U6937 (N_6937,N_6716,N_6790);
nand U6938 (N_6938,N_6764,N_6617);
or U6939 (N_6939,N_6773,N_6702);
or U6940 (N_6940,N_6668,N_6622);
and U6941 (N_6941,N_6776,N_6706);
and U6942 (N_6942,N_6756,N_6613);
nand U6943 (N_6943,N_6600,N_6644);
nor U6944 (N_6944,N_6696,N_6679);
or U6945 (N_6945,N_6765,N_6627);
and U6946 (N_6946,N_6617,N_6662);
or U6947 (N_6947,N_6712,N_6756);
and U6948 (N_6948,N_6731,N_6781);
and U6949 (N_6949,N_6629,N_6602);
and U6950 (N_6950,N_6687,N_6719);
nor U6951 (N_6951,N_6693,N_6760);
nand U6952 (N_6952,N_6642,N_6794);
nor U6953 (N_6953,N_6731,N_6655);
nand U6954 (N_6954,N_6757,N_6700);
and U6955 (N_6955,N_6749,N_6661);
nor U6956 (N_6956,N_6655,N_6684);
and U6957 (N_6957,N_6718,N_6621);
or U6958 (N_6958,N_6668,N_6662);
nand U6959 (N_6959,N_6604,N_6766);
nand U6960 (N_6960,N_6634,N_6764);
nand U6961 (N_6961,N_6625,N_6699);
or U6962 (N_6962,N_6727,N_6775);
nor U6963 (N_6963,N_6633,N_6704);
nand U6964 (N_6964,N_6647,N_6676);
or U6965 (N_6965,N_6767,N_6792);
or U6966 (N_6966,N_6630,N_6768);
nor U6967 (N_6967,N_6745,N_6635);
or U6968 (N_6968,N_6734,N_6616);
and U6969 (N_6969,N_6686,N_6607);
and U6970 (N_6970,N_6714,N_6710);
nor U6971 (N_6971,N_6653,N_6692);
and U6972 (N_6972,N_6707,N_6756);
nor U6973 (N_6973,N_6613,N_6798);
or U6974 (N_6974,N_6750,N_6618);
or U6975 (N_6975,N_6699,N_6761);
or U6976 (N_6976,N_6652,N_6663);
or U6977 (N_6977,N_6632,N_6602);
nand U6978 (N_6978,N_6603,N_6625);
nor U6979 (N_6979,N_6616,N_6606);
and U6980 (N_6980,N_6619,N_6717);
and U6981 (N_6981,N_6712,N_6644);
nor U6982 (N_6982,N_6611,N_6796);
nor U6983 (N_6983,N_6668,N_6635);
and U6984 (N_6984,N_6739,N_6742);
nor U6985 (N_6985,N_6769,N_6764);
and U6986 (N_6986,N_6660,N_6776);
nand U6987 (N_6987,N_6776,N_6713);
or U6988 (N_6988,N_6657,N_6786);
nand U6989 (N_6989,N_6739,N_6751);
or U6990 (N_6990,N_6713,N_6681);
nand U6991 (N_6991,N_6780,N_6632);
nand U6992 (N_6992,N_6689,N_6631);
or U6993 (N_6993,N_6709,N_6639);
and U6994 (N_6994,N_6676,N_6784);
nor U6995 (N_6995,N_6786,N_6637);
and U6996 (N_6996,N_6797,N_6686);
and U6997 (N_6997,N_6717,N_6742);
nand U6998 (N_6998,N_6754,N_6653);
nor U6999 (N_6999,N_6749,N_6627);
or U7000 (N_7000,N_6972,N_6956);
and U7001 (N_7001,N_6855,N_6865);
and U7002 (N_7002,N_6905,N_6935);
and U7003 (N_7003,N_6928,N_6950);
and U7004 (N_7004,N_6835,N_6947);
or U7005 (N_7005,N_6879,N_6929);
and U7006 (N_7006,N_6953,N_6886);
or U7007 (N_7007,N_6927,N_6993);
nand U7008 (N_7008,N_6961,N_6844);
nand U7009 (N_7009,N_6804,N_6819);
nor U7010 (N_7010,N_6824,N_6943);
or U7011 (N_7011,N_6944,N_6998);
and U7012 (N_7012,N_6901,N_6995);
or U7013 (N_7013,N_6951,N_6881);
nor U7014 (N_7014,N_6888,N_6921);
or U7015 (N_7015,N_6802,N_6955);
nor U7016 (N_7016,N_6911,N_6945);
nand U7017 (N_7017,N_6884,N_6968);
nand U7018 (N_7018,N_6885,N_6827);
or U7019 (N_7019,N_6992,N_6974);
or U7020 (N_7020,N_6948,N_6898);
or U7021 (N_7021,N_6967,N_6848);
nand U7022 (N_7022,N_6839,N_6832);
or U7023 (N_7023,N_6861,N_6949);
nor U7024 (N_7024,N_6803,N_6829);
or U7025 (N_7025,N_6854,N_6979);
nand U7026 (N_7026,N_6999,N_6836);
nand U7027 (N_7027,N_6860,N_6876);
and U7028 (N_7028,N_6871,N_6982);
nand U7029 (N_7029,N_6915,N_6990);
nor U7030 (N_7030,N_6984,N_6913);
nand U7031 (N_7031,N_6908,N_6969);
nand U7032 (N_7032,N_6826,N_6838);
and U7033 (N_7033,N_6882,N_6966);
nand U7034 (N_7034,N_6933,N_6801);
or U7035 (N_7035,N_6852,N_6906);
nand U7036 (N_7036,N_6963,N_6834);
and U7037 (N_7037,N_6907,N_6866);
nand U7038 (N_7038,N_6870,N_6980);
nor U7039 (N_7039,N_6811,N_6914);
nand U7040 (N_7040,N_6846,N_6892);
or U7041 (N_7041,N_6809,N_6930);
and U7042 (N_7042,N_6814,N_6973);
nand U7043 (N_7043,N_6845,N_6987);
and U7044 (N_7044,N_6925,N_6924);
and U7045 (N_7045,N_6878,N_6877);
nand U7046 (N_7046,N_6857,N_6837);
and U7047 (N_7047,N_6828,N_6812);
and U7048 (N_7048,N_6936,N_6981);
nor U7049 (N_7049,N_6899,N_6849);
nand U7050 (N_7050,N_6867,N_6931);
and U7051 (N_7051,N_6988,N_6853);
or U7052 (N_7052,N_6922,N_6895);
nor U7053 (N_7053,N_6850,N_6806);
and U7054 (N_7054,N_6964,N_6900);
nand U7055 (N_7055,N_6940,N_6941);
xor U7056 (N_7056,N_6820,N_6821);
or U7057 (N_7057,N_6986,N_6926);
nand U7058 (N_7058,N_6869,N_6810);
or U7059 (N_7059,N_6958,N_6939);
nor U7060 (N_7060,N_6934,N_6959);
or U7061 (N_7061,N_6863,N_6868);
xor U7062 (N_7062,N_6874,N_6938);
and U7063 (N_7063,N_6887,N_6997);
nor U7064 (N_7064,N_6816,N_6996);
nor U7065 (N_7065,N_6889,N_6912);
nand U7066 (N_7066,N_6965,N_6991);
and U7067 (N_7067,N_6962,N_6893);
or U7068 (N_7068,N_6942,N_6808);
nor U7069 (N_7069,N_6970,N_6872);
or U7070 (N_7070,N_6843,N_6890);
nor U7071 (N_7071,N_6971,N_6957);
nor U7072 (N_7072,N_6946,N_6891);
nor U7073 (N_7073,N_6818,N_6864);
or U7074 (N_7074,N_6875,N_6985);
nor U7075 (N_7075,N_6920,N_6873);
and U7076 (N_7076,N_6918,N_6896);
nor U7077 (N_7077,N_6817,N_6989);
nor U7078 (N_7078,N_6894,N_6960);
or U7079 (N_7079,N_6976,N_6916);
nor U7080 (N_7080,N_6954,N_6851);
or U7081 (N_7081,N_6859,N_6823);
or U7082 (N_7082,N_6932,N_6880);
or U7083 (N_7083,N_6883,N_6897);
nand U7084 (N_7084,N_6847,N_6903);
or U7085 (N_7085,N_6978,N_6858);
nor U7086 (N_7086,N_6841,N_6983);
nand U7087 (N_7087,N_6937,N_6977);
nand U7088 (N_7088,N_6975,N_6952);
xor U7089 (N_7089,N_6862,N_6904);
nor U7090 (N_7090,N_6994,N_6917);
nor U7091 (N_7091,N_6807,N_6825);
or U7092 (N_7092,N_6923,N_6822);
and U7093 (N_7093,N_6842,N_6840);
or U7094 (N_7094,N_6909,N_6910);
nand U7095 (N_7095,N_6805,N_6902);
or U7096 (N_7096,N_6919,N_6813);
or U7097 (N_7097,N_6833,N_6830);
nor U7098 (N_7098,N_6856,N_6800);
and U7099 (N_7099,N_6815,N_6831);
nand U7100 (N_7100,N_6854,N_6925);
or U7101 (N_7101,N_6962,N_6909);
and U7102 (N_7102,N_6870,N_6810);
nor U7103 (N_7103,N_6862,N_6829);
nor U7104 (N_7104,N_6896,N_6967);
or U7105 (N_7105,N_6959,N_6897);
or U7106 (N_7106,N_6980,N_6929);
and U7107 (N_7107,N_6809,N_6861);
or U7108 (N_7108,N_6904,N_6819);
nor U7109 (N_7109,N_6958,N_6880);
nand U7110 (N_7110,N_6803,N_6837);
nand U7111 (N_7111,N_6911,N_6933);
nand U7112 (N_7112,N_6939,N_6922);
nor U7113 (N_7113,N_6941,N_6949);
and U7114 (N_7114,N_6968,N_6897);
or U7115 (N_7115,N_6955,N_6801);
or U7116 (N_7116,N_6993,N_6845);
or U7117 (N_7117,N_6903,N_6937);
nand U7118 (N_7118,N_6917,N_6892);
nor U7119 (N_7119,N_6886,N_6940);
nor U7120 (N_7120,N_6823,N_6868);
nand U7121 (N_7121,N_6836,N_6807);
or U7122 (N_7122,N_6836,N_6816);
nand U7123 (N_7123,N_6814,N_6932);
nand U7124 (N_7124,N_6819,N_6846);
xnor U7125 (N_7125,N_6862,N_6924);
nand U7126 (N_7126,N_6943,N_6901);
and U7127 (N_7127,N_6888,N_6893);
or U7128 (N_7128,N_6810,N_6923);
and U7129 (N_7129,N_6835,N_6920);
nor U7130 (N_7130,N_6998,N_6862);
and U7131 (N_7131,N_6996,N_6824);
or U7132 (N_7132,N_6944,N_6840);
nor U7133 (N_7133,N_6813,N_6802);
and U7134 (N_7134,N_6995,N_6805);
or U7135 (N_7135,N_6913,N_6893);
or U7136 (N_7136,N_6902,N_6855);
nor U7137 (N_7137,N_6827,N_6868);
or U7138 (N_7138,N_6955,N_6882);
and U7139 (N_7139,N_6807,N_6974);
or U7140 (N_7140,N_6849,N_6982);
or U7141 (N_7141,N_6852,N_6934);
or U7142 (N_7142,N_6949,N_6915);
nor U7143 (N_7143,N_6901,N_6986);
nand U7144 (N_7144,N_6873,N_6838);
or U7145 (N_7145,N_6901,N_6860);
nor U7146 (N_7146,N_6893,N_6970);
nor U7147 (N_7147,N_6885,N_6955);
nand U7148 (N_7148,N_6927,N_6978);
nand U7149 (N_7149,N_6964,N_6827);
or U7150 (N_7150,N_6894,N_6858);
and U7151 (N_7151,N_6845,N_6805);
nor U7152 (N_7152,N_6885,N_6943);
and U7153 (N_7153,N_6816,N_6957);
or U7154 (N_7154,N_6887,N_6959);
nand U7155 (N_7155,N_6941,N_6840);
or U7156 (N_7156,N_6930,N_6931);
nor U7157 (N_7157,N_6821,N_6936);
nand U7158 (N_7158,N_6896,N_6899);
or U7159 (N_7159,N_6863,N_6882);
nand U7160 (N_7160,N_6945,N_6845);
and U7161 (N_7161,N_6904,N_6960);
nand U7162 (N_7162,N_6811,N_6984);
nand U7163 (N_7163,N_6882,N_6951);
nor U7164 (N_7164,N_6850,N_6894);
or U7165 (N_7165,N_6951,N_6939);
nand U7166 (N_7166,N_6989,N_6883);
xnor U7167 (N_7167,N_6837,N_6878);
or U7168 (N_7168,N_6925,N_6920);
nor U7169 (N_7169,N_6867,N_6913);
nand U7170 (N_7170,N_6850,N_6945);
or U7171 (N_7171,N_6929,N_6835);
nand U7172 (N_7172,N_6909,N_6852);
and U7173 (N_7173,N_6815,N_6976);
or U7174 (N_7174,N_6948,N_6840);
and U7175 (N_7175,N_6922,N_6860);
or U7176 (N_7176,N_6956,N_6955);
nor U7177 (N_7177,N_6926,N_6812);
nor U7178 (N_7178,N_6988,N_6898);
or U7179 (N_7179,N_6806,N_6813);
or U7180 (N_7180,N_6833,N_6836);
and U7181 (N_7181,N_6956,N_6882);
or U7182 (N_7182,N_6831,N_6808);
nor U7183 (N_7183,N_6813,N_6994);
or U7184 (N_7184,N_6827,N_6976);
or U7185 (N_7185,N_6962,N_6998);
or U7186 (N_7186,N_6845,N_6867);
nor U7187 (N_7187,N_6996,N_6944);
and U7188 (N_7188,N_6805,N_6975);
nand U7189 (N_7189,N_6983,N_6806);
nand U7190 (N_7190,N_6896,N_6988);
nor U7191 (N_7191,N_6894,N_6851);
nand U7192 (N_7192,N_6975,N_6871);
nand U7193 (N_7193,N_6946,N_6980);
or U7194 (N_7194,N_6930,N_6828);
and U7195 (N_7195,N_6901,N_6830);
nand U7196 (N_7196,N_6931,N_6983);
nor U7197 (N_7197,N_6935,N_6860);
or U7198 (N_7198,N_6835,N_6903);
nor U7199 (N_7199,N_6870,N_6860);
or U7200 (N_7200,N_7190,N_7046);
xnor U7201 (N_7201,N_7069,N_7050);
or U7202 (N_7202,N_7136,N_7149);
nor U7203 (N_7203,N_7191,N_7144);
and U7204 (N_7204,N_7185,N_7193);
nand U7205 (N_7205,N_7024,N_7034);
and U7206 (N_7206,N_7169,N_7143);
nand U7207 (N_7207,N_7103,N_7117);
and U7208 (N_7208,N_7062,N_7019);
nor U7209 (N_7209,N_7058,N_7037);
nand U7210 (N_7210,N_7110,N_7151);
nand U7211 (N_7211,N_7048,N_7195);
nor U7212 (N_7212,N_7150,N_7043);
nand U7213 (N_7213,N_7112,N_7056);
nand U7214 (N_7214,N_7168,N_7099);
or U7215 (N_7215,N_7017,N_7086);
nor U7216 (N_7216,N_7145,N_7035);
and U7217 (N_7217,N_7176,N_7119);
nand U7218 (N_7218,N_7005,N_7045);
nor U7219 (N_7219,N_7076,N_7135);
nand U7220 (N_7220,N_7159,N_7125);
nand U7221 (N_7221,N_7036,N_7071);
nand U7222 (N_7222,N_7057,N_7038);
and U7223 (N_7223,N_7118,N_7018);
or U7224 (N_7224,N_7180,N_7002);
or U7225 (N_7225,N_7000,N_7140);
and U7226 (N_7226,N_7192,N_7187);
and U7227 (N_7227,N_7166,N_7148);
nand U7228 (N_7228,N_7108,N_7027);
or U7229 (N_7229,N_7109,N_7165);
and U7230 (N_7230,N_7101,N_7152);
nand U7231 (N_7231,N_7177,N_7132);
nor U7232 (N_7232,N_7011,N_7020);
and U7233 (N_7233,N_7074,N_7006);
and U7234 (N_7234,N_7078,N_7080);
nand U7235 (N_7235,N_7053,N_7022);
nor U7236 (N_7236,N_7033,N_7008);
nand U7237 (N_7237,N_7001,N_7063);
xor U7238 (N_7238,N_7194,N_7023);
or U7239 (N_7239,N_7147,N_7129);
or U7240 (N_7240,N_7072,N_7173);
and U7241 (N_7241,N_7097,N_7095);
or U7242 (N_7242,N_7188,N_7164);
nand U7243 (N_7243,N_7060,N_7041);
nor U7244 (N_7244,N_7088,N_7131);
and U7245 (N_7245,N_7175,N_7123);
or U7246 (N_7246,N_7089,N_7133);
or U7247 (N_7247,N_7160,N_7146);
nor U7248 (N_7248,N_7107,N_7127);
and U7249 (N_7249,N_7092,N_7199);
and U7250 (N_7250,N_7098,N_7137);
or U7251 (N_7251,N_7021,N_7039);
or U7252 (N_7252,N_7007,N_7163);
and U7253 (N_7253,N_7031,N_7126);
or U7254 (N_7254,N_7172,N_7154);
and U7255 (N_7255,N_7104,N_7084);
or U7256 (N_7256,N_7082,N_7087);
or U7257 (N_7257,N_7004,N_7196);
nor U7258 (N_7258,N_7028,N_7061);
nor U7259 (N_7259,N_7156,N_7009);
xor U7260 (N_7260,N_7085,N_7124);
nor U7261 (N_7261,N_7174,N_7029);
nand U7262 (N_7262,N_7070,N_7134);
nand U7263 (N_7263,N_7003,N_7167);
nor U7264 (N_7264,N_7186,N_7114);
and U7265 (N_7265,N_7179,N_7197);
and U7266 (N_7266,N_7161,N_7025);
and U7267 (N_7267,N_7016,N_7051);
and U7268 (N_7268,N_7157,N_7065);
nand U7269 (N_7269,N_7010,N_7183);
and U7270 (N_7270,N_7121,N_7105);
and U7271 (N_7271,N_7064,N_7142);
nand U7272 (N_7272,N_7158,N_7052);
nor U7273 (N_7273,N_7171,N_7130);
nor U7274 (N_7274,N_7115,N_7155);
or U7275 (N_7275,N_7015,N_7083);
nand U7276 (N_7276,N_7032,N_7040);
or U7277 (N_7277,N_7106,N_7102);
or U7278 (N_7278,N_7111,N_7075);
nand U7279 (N_7279,N_7030,N_7077);
xnor U7280 (N_7280,N_7081,N_7055);
and U7281 (N_7281,N_7153,N_7073);
and U7282 (N_7282,N_7054,N_7026);
nor U7283 (N_7283,N_7091,N_7181);
nand U7284 (N_7284,N_7059,N_7096);
nand U7285 (N_7285,N_7162,N_7066);
or U7286 (N_7286,N_7128,N_7116);
nand U7287 (N_7287,N_7014,N_7068);
nor U7288 (N_7288,N_7042,N_7047);
or U7289 (N_7289,N_7044,N_7113);
nand U7290 (N_7290,N_7184,N_7120);
and U7291 (N_7291,N_7013,N_7178);
and U7292 (N_7292,N_7141,N_7012);
and U7293 (N_7293,N_7122,N_7138);
or U7294 (N_7294,N_7182,N_7198);
xnor U7295 (N_7295,N_7079,N_7094);
nor U7296 (N_7296,N_7189,N_7093);
or U7297 (N_7297,N_7100,N_7049);
or U7298 (N_7298,N_7139,N_7170);
xnor U7299 (N_7299,N_7067,N_7090);
or U7300 (N_7300,N_7013,N_7138);
nor U7301 (N_7301,N_7119,N_7181);
nor U7302 (N_7302,N_7069,N_7062);
nor U7303 (N_7303,N_7025,N_7183);
nand U7304 (N_7304,N_7168,N_7143);
nand U7305 (N_7305,N_7020,N_7159);
nor U7306 (N_7306,N_7097,N_7062);
xnor U7307 (N_7307,N_7110,N_7036);
nor U7308 (N_7308,N_7110,N_7182);
nor U7309 (N_7309,N_7114,N_7060);
nand U7310 (N_7310,N_7107,N_7112);
and U7311 (N_7311,N_7042,N_7006);
or U7312 (N_7312,N_7109,N_7044);
nand U7313 (N_7313,N_7158,N_7145);
nor U7314 (N_7314,N_7001,N_7117);
and U7315 (N_7315,N_7099,N_7106);
nor U7316 (N_7316,N_7106,N_7153);
or U7317 (N_7317,N_7110,N_7192);
and U7318 (N_7318,N_7199,N_7005);
or U7319 (N_7319,N_7161,N_7181);
nor U7320 (N_7320,N_7099,N_7122);
or U7321 (N_7321,N_7092,N_7138);
nand U7322 (N_7322,N_7083,N_7142);
nor U7323 (N_7323,N_7105,N_7166);
and U7324 (N_7324,N_7052,N_7182);
nor U7325 (N_7325,N_7058,N_7150);
and U7326 (N_7326,N_7183,N_7181);
xor U7327 (N_7327,N_7198,N_7073);
and U7328 (N_7328,N_7175,N_7143);
xor U7329 (N_7329,N_7156,N_7143);
nor U7330 (N_7330,N_7023,N_7054);
nand U7331 (N_7331,N_7002,N_7178);
nand U7332 (N_7332,N_7147,N_7139);
nor U7333 (N_7333,N_7197,N_7193);
nor U7334 (N_7334,N_7063,N_7100);
nor U7335 (N_7335,N_7100,N_7170);
or U7336 (N_7336,N_7028,N_7148);
nand U7337 (N_7337,N_7089,N_7189);
nor U7338 (N_7338,N_7041,N_7094);
and U7339 (N_7339,N_7049,N_7062);
nor U7340 (N_7340,N_7049,N_7057);
nand U7341 (N_7341,N_7107,N_7000);
nor U7342 (N_7342,N_7150,N_7092);
nand U7343 (N_7343,N_7189,N_7078);
nand U7344 (N_7344,N_7148,N_7165);
and U7345 (N_7345,N_7126,N_7102);
and U7346 (N_7346,N_7025,N_7017);
nor U7347 (N_7347,N_7191,N_7171);
nand U7348 (N_7348,N_7148,N_7135);
nand U7349 (N_7349,N_7175,N_7058);
or U7350 (N_7350,N_7173,N_7098);
nand U7351 (N_7351,N_7189,N_7187);
nand U7352 (N_7352,N_7185,N_7046);
or U7353 (N_7353,N_7184,N_7175);
or U7354 (N_7354,N_7109,N_7054);
nand U7355 (N_7355,N_7188,N_7161);
nand U7356 (N_7356,N_7181,N_7014);
nand U7357 (N_7357,N_7189,N_7117);
or U7358 (N_7358,N_7000,N_7179);
and U7359 (N_7359,N_7016,N_7060);
nor U7360 (N_7360,N_7004,N_7182);
or U7361 (N_7361,N_7160,N_7086);
and U7362 (N_7362,N_7122,N_7182);
or U7363 (N_7363,N_7159,N_7046);
xnor U7364 (N_7364,N_7057,N_7117);
or U7365 (N_7365,N_7076,N_7196);
and U7366 (N_7366,N_7187,N_7156);
or U7367 (N_7367,N_7076,N_7123);
and U7368 (N_7368,N_7183,N_7018);
nor U7369 (N_7369,N_7118,N_7035);
nand U7370 (N_7370,N_7021,N_7019);
and U7371 (N_7371,N_7171,N_7097);
nor U7372 (N_7372,N_7121,N_7046);
or U7373 (N_7373,N_7178,N_7032);
and U7374 (N_7374,N_7009,N_7174);
nor U7375 (N_7375,N_7167,N_7061);
nand U7376 (N_7376,N_7105,N_7110);
nand U7377 (N_7377,N_7018,N_7029);
and U7378 (N_7378,N_7081,N_7025);
or U7379 (N_7379,N_7158,N_7062);
or U7380 (N_7380,N_7137,N_7186);
nand U7381 (N_7381,N_7052,N_7162);
nand U7382 (N_7382,N_7193,N_7021);
and U7383 (N_7383,N_7006,N_7125);
or U7384 (N_7384,N_7185,N_7145);
or U7385 (N_7385,N_7142,N_7191);
nand U7386 (N_7386,N_7193,N_7010);
nand U7387 (N_7387,N_7193,N_7191);
and U7388 (N_7388,N_7164,N_7040);
nand U7389 (N_7389,N_7007,N_7035);
nand U7390 (N_7390,N_7008,N_7000);
and U7391 (N_7391,N_7156,N_7149);
nand U7392 (N_7392,N_7042,N_7026);
and U7393 (N_7393,N_7092,N_7015);
and U7394 (N_7394,N_7081,N_7049);
or U7395 (N_7395,N_7055,N_7036);
nor U7396 (N_7396,N_7165,N_7189);
nand U7397 (N_7397,N_7122,N_7080);
nand U7398 (N_7398,N_7152,N_7163);
and U7399 (N_7399,N_7121,N_7195);
or U7400 (N_7400,N_7384,N_7280);
nor U7401 (N_7401,N_7247,N_7326);
nor U7402 (N_7402,N_7216,N_7312);
nor U7403 (N_7403,N_7235,N_7253);
nand U7404 (N_7404,N_7386,N_7376);
and U7405 (N_7405,N_7282,N_7393);
or U7406 (N_7406,N_7211,N_7274);
nand U7407 (N_7407,N_7308,N_7331);
or U7408 (N_7408,N_7323,N_7379);
and U7409 (N_7409,N_7392,N_7248);
and U7410 (N_7410,N_7267,N_7303);
xnor U7411 (N_7411,N_7349,N_7373);
and U7412 (N_7412,N_7300,N_7311);
nand U7413 (N_7413,N_7277,N_7377);
nor U7414 (N_7414,N_7363,N_7254);
nand U7415 (N_7415,N_7299,N_7321);
nand U7416 (N_7416,N_7297,N_7245);
nor U7417 (N_7417,N_7304,N_7344);
nand U7418 (N_7418,N_7234,N_7309);
nor U7419 (N_7419,N_7342,N_7389);
or U7420 (N_7420,N_7289,N_7357);
and U7421 (N_7421,N_7343,N_7364);
or U7422 (N_7422,N_7292,N_7313);
or U7423 (N_7423,N_7307,N_7334);
or U7424 (N_7424,N_7291,N_7367);
nor U7425 (N_7425,N_7257,N_7325);
and U7426 (N_7426,N_7310,N_7224);
nand U7427 (N_7427,N_7399,N_7258);
or U7428 (N_7428,N_7210,N_7232);
xor U7429 (N_7429,N_7271,N_7330);
and U7430 (N_7430,N_7220,N_7371);
nor U7431 (N_7431,N_7221,N_7388);
and U7432 (N_7432,N_7246,N_7242);
or U7433 (N_7433,N_7238,N_7360);
or U7434 (N_7434,N_7230,N_7239);
or U7435 (N_7435,N_7290,N_7281);
nor U7436 (N_7436,N_7329,N_7298);
nand U7437 (N_7437,N_7215,N_7362);
or U7438 (N_7438,N_7397,N_7279);
nor U7439 (N_7439,N_7315,N_7390);
nor U7440 (N_7440,N_7278,N_7204);
or U7441 (N_7441,N_7340,N_7252);
and U7442 (N_7442,N_7333,N_7328);
nand U7443 (N_7443,N_7263,N_7265);
and U7444 (N_7444,N_7214,N_7207);
nand U7445 (N_7445,N_7370,N_7346);
nand U7446 (N_7446,N_7345,N_7341);
and U7447 (N_7447,N_7203,N_7395);
nor U7448 (N_7448,N_7361,N_7213);
or U7449 (N_7449,N_7259,N_7233);
nor U7450 (N_7450,N_7359,N_7229);
nand U7451 (N_7451,N_7250,N_7375);
nor U7452 (N_7452,N_7305,N_7217);
and U7453 (N_7453,N_7318,N_7355);
nand U7454 (N_7454,N_7222,N_7249);
and U7455 (N_7455,N_7358,N_7372);
and U7456 (N_7456,N_7243,N_7244);
and U7457 (N_7457,N_7284,N_7205);
and U7458 (N_7458,N_7206,N_7332);
and U7459 (N_7459,N_7294,N_7268);
nand U7460 (N_7460,N_7296,N_7208);
and U7461 (N_7461,N_7369,N_7365);
and U7462 (N_7462,N_7200,N_7269);
nand U7463 (N_7463,N_7273,N_7285);
nand U7464 (N_7464,N_7255,N_7236);
nor U7465 (N_7465,N_7382,N_7225);
and U7466 (N_7466,N_7283,N_7251);
and U7467 (N_7467,N_7383,N_7352);
nand U7468 (N_7468,N_7264,N_7356);
nor U7469 (N_7469,N_7385,N_7348);
or U7470 (N_7470,N_7338,N_7260);
or U7471 (N_7471,N_7316,N_7394);
nor U7472 (N_7472,N_7398,N_7314);
nor U7473 (N_7473,N_7347,N_7387);
or U7474 (N_7474,N_7212,N_7261);
and U7475 (N_7475,N_7324,N_7262);
and U7476 (N_7476,N_7380,N_7219);
or U7477 (N_7477,N_7337,N_7288);
or U7478 (N_7478,N_7378,N_7276);
or U7479 (N_7479,N_7354,N_7223);
or U7480 (N_7480,N_7240,N_7339);
or U7481 (N_7481,N_7241,N_7396);
or U7482 (N_7482,N_7295,N_7202);
or U7483 (N_7483,N_7287,N_7231);
nand U7484 (N_7484,N_7327,N_7286);
nor U7485 (N_7485,N_7228,N_7319);
nand U7486 (N_7486,N_7322,N_7256);
or U7487 (N_7487,N_7301,N_7270);
nand U7488 (N_7488,N_7226,N_7391);
and U7489 (N_7489,N_7366,N_7350);
or U7490 (N_7490,N_7320,N_7201);
and U7491 (N_7491,N_7351,N_7293);
nor U7492 (N_7492,N_7237,N_7335);
nand U7493 (N_7493,N_7306,N_7317);
and U7494 (N_7494,N_7266,N_7275);
and U7495 (N_7495,N_7353,N_7381);
and U7496 (N_7496,N_7368,N_7272);
or U7497 (N_7497,N_7336,N_7227);
and U7498 (N_7498,N_7218,N_7209);
or U7499 (N_7499,N_7302,N_7374);
nand U7500 (N_7500,N_7361,N_7200);
and U7501 (N_7501,N_7247,N_7287);
or U7502 (N_7502,N_7261,N_7392);
nand U7503 (N_7503,N_7312,N_7272);
or U7504 (N_7504,N_7269,N_7266);
and U7505 (N_7505,N_7302,N_7375);
or U7506 (N_7506,N_7259,N_7313);
nand U7507 (N_7507,N_7235,N_7392);
nor U7508 (N_7508,N_7288,N_7212);
nand U7509 (N_7509,N_7211,N_7250);
nand U7510 (N_7510,N_7371,N_7222);
nor U7511 (N_7511,N_7244,N_7376);
nand U7512 (N_7512,N_7263,N_7345);
or U7513 (N_7513,N_7319,N_7201);
nor U7514 (N_7514,N_7263,N_7261);
and U7515 (N_7515,N_7398,N_7280);
and U7516 (N_7516,N_7360,N_7247);
nand U7517 (N_7517,N_7205,N_7233);
nand U7518 (N_7518,N_7382,N_7209);
or U7519 (N_7519,N_7201,N_7378);
or U7520 (N_7520,N_7399,N_7274);
nand U7521 (N_7521,N_7235,N_7273);
nor U7522 (N_7522,N_7386,N_7351);
nand U7523 (N_7523,N_7294,N_7395);
nor U7524 (N_7524,N_7288,N_7374);
nor U7525 (N_7525,N_7282,N_7216);
and U7526 (N_7526,N_7280,N_7348);
and U7527 (N_7527,N_7395,N_7219);
nand U7528 (N_7528,N_7286,N_7396);
or U7529 (N_7529,N_7297,N_7330);
nor U7530 (N_7530,N_7319,N_7217);
nand U7531 (N_7531,N_7369,N_7240);
and U7532 (N_7532,N_7310,N_7221);
xor U7533 (N_7533,N_7323,N_7328);
or U7534 (N_7534,N_7223,N_7234);
and U7535 (N_7535,N_7359,N_7356);
and U7536 (N_7536,N_7336,N_7361);
and U7537 (N_7537,N_7296,N_7341);
or U7538 (N_7538,N_7308,N_7208);
or U7539 (N_7539,N_7236,N_7261);
nand U7540 (N_7540,N_7265,N_7239);
nand U7541 (N_7541,N_7298,N_7277);
and U7542 (N_7542,N_7200,N_7242);
nand U7543 (N_7543,N_7233,N_7360);
nor U7544 (N_7544,N_7203,N_7230);
and U7545 (N_7545,N_7256,N_7374);
and U7546 (N_7546,N_7359,N_7255);
and U7547 (N_7547,N_7303,N_7237);
and U7548 (N_7548,N_7249,N_7307);
nor U7549 (N_7549,N_7390,N_7295);
nor U7550 (N_7550,N_7251,N_7278);
nor U7551 (N_7551,N_7301,N_7223);
or U7552 (N_7552,N_7241,N_7237);
or U7553 (N_7553,N_7288,N_7232);
and U7554 (N_7554,N_7305,N_7359);
nand U7555 (N_7555,N_7252,N_7389);
nand U7556 (N_7556,N_7374,N_7356);
nand U7557 (N_7557,N_7350,N_7317);
nand U7558 (N_7558,N_7208,N_7263);
nand U7559 (N_7559,N_7356,N_7312);
or U7560 (N_7560,N_7343,N_7351);
or U7561 (N_7561,N_7397,N_7208);
nand U7562 (N_7562,N_7381,N_7209);
nand U7563 (N_7563,N_7333,N_7226);
or U7564 (N_7564,N_7311,N_7352);
or U7565 (N_7565,N_7331,N_7265);
and U7566 (N_7566,N_7377,N_7381);
and U7567 (N_7567,N_7366,N_7305);
and U7568 (N_7568,N_7335,N_7341);
and U7569 (N_7569,N_7214,N_7345);
nor U7570 (N_7570,N_7309,N_7212);
or U7571 (N_7571,N_7360,N_7267);
nor U7572 (N_7572,N_7226,N_7205);
and U7573 (N_7573,N_7219,N_7257);
and U7574 (N_7574,N_7201,N_7215);
nand U7575 (N_7575,N_7314,N_7300);
nor U7576 (N_7576,N_7289,N_7373);
nand U7577 (N_7577,N_7347,N_7206);
nor U7578 (N_7578,N_7320,N_7379);
nand U7579 (N_7579,N_7355,N_7256);
and U7580 (N_7580,N_7292,N_7323);
or U7581 (N_7581,N_7232,N_7373);
and U7582 (N_7582,N_7359,N_7399);
or U7583 (N_7583,N_7377,N_7296);
or U7584 (N_7584,N_7290,N_7288);
or U7585 (N_7585,N_7336,N_7360);
or U7586 (N_7586,N_7383,N_7359);
nand U7587 (N_7587,N_7259,N_7252);
nand U7588 (N_7588,N_7257,N_7234);
or U7589 (N_7589,N_7367,N_7260);
and U7590 (N_7590,N_7291,N_7289);
nor U7591 (N_7591,N_7206,N_7341);
nand U7592 (N_7592,N_7398,N_7385);
nor U7593 (N_7593,N_7234,N_7379);
nor U7594 (N_7594,N_7360,N_7330);
nor U7595 (N_7595,N_7318,N_7245);
nand U7596 (N_7596,N_7221,N_7236);
nand U7597 (N_7597,N_7300,N_7253);
nor U7598 (N_7598,N_7341,N_7208);
nand U7599 (N_7599,N_7310,N_7248);
nand U7600 (N_7600,N_7447,N_7459);
or U7601 (N_7601,N_7417,N_7463);
nand U7602 (N_7602,N_7584,N_7458);
or U7603 (N_7603,N_7405,N_7531);
nor U7604 (N_7604,N_7595,N_7593);
nor U7605 (N_7605,N_7551,N_7425);
nor U7606 (N_7606,N_7481,N_7577);
nand U7607 (N_7607,N_7498,N_7587);
and U7608 (N_7608,N_7528,N_7484);
nand U7609 (N_7609,N_7557,N_7583);
nor U7610 (N_7610,N_7424,N_7590);
nor U7611 (N_7611,N_7407,N_7454);
nor U7612 (N_7612,N_7455,N_7576);
and U7613 (N_7613,N_7443,N_7538);
nor U7614 (N_7614,N_7439,N_7569);
or U7615 (N_7615,N_7422,N_7536);
or U7616 (N_7616,N_7548,N_7586);
nand U7617 (N_7617,N_7598,N_7568);
nand U7618 (N_7618,N_7433,N_7563);
nor U7619 (N_7619,N_7520,N_7483);
nand U7620 (N_7620,N_7549,N_7490);
and U7621 (N_7621,N_7545,N_7402);
nand U7622 (N_7622,N_7410,N_7527);
nor U7623 (N_7623,N_7512,N_7477);
nand U7624 (N_7624,N_7404,N_7550);
nor U7625 (N_7625,N_7432,N_7599);
or U7626 (N_7626,N_7436,N_7450);
or U7627 (N_7627,N_7581,N_7441);
and U7628 (N_7628,N_7486,N_7501);
nor U7629 (N_7629,N_7438,N_7535);
or U7630 (N_7630,N_7468,N_7591);
nand U7631 (N_7631,N_7554,N_7465);
nand U7632 (N_7632,N_7427,N_7406);
nand U7633 (N_7633,N_7524,N_7502);
or U7634 (N_7634,N_7580,N_7411);
nand U7635 (N_7635,N_7469,N_7567);
and U7636 (N_7636,N_7592,N_7519);
nor U7637 (N_7637,N_7482,N_7420);
nand U7638 (N_7638,N_7491,N_7513);
and U7639 (N_7639,N_7423,N_7456);
nor U7640 (N_7640,N_7471,N_7431);
or U7641 (N_7641,N_7434,N_7594);
or U7642 (N_7642,N_7476,N_7445);
or U7643 (N_7643,N_7552,N_7561);
nor U7644 (N_7644,N_7475,N_7492);
nor U7645 (N_7645,N_7571,N_7559);
nor U7646 (N_7646,N_7564,N_7523);
and U7647 (N_7647,N_7579,N_7509);
nand U7648 (N_7648,N_7573,N_7496);
nor U7649 (N_7649,N_7414,N_7578);
nand U7650 (N_7650,N_7534,N_7572);
nand U7651 (N_7651,N_7495,N_7460);
nor U7652 (N_7652,N_7542,N_7472);
nand U7653 (N_7653,N_7413,N_7547);
nor U7654 (N_7654,N_7400,N_7487);
nand U7655 (N_7655,N_7499,N_7466);
and U7656 (N_7656,N_7588,N_7493);
nor U7657 (N_7657,N_7541,N_7409);
nand U7658 (N_7658,N_7488,N_7589);
or U7659 (N_7659,N_7452,N_7516);
nand U7660 (N_7660,N_7401,N_7480);
nand U7661 (N_7661,N_7530,N_7521);
and U7662 (N_7662,N_7506,N_7470);
nand U7663 (N_7663,N_7555,N_7457);
nand U7664 (N_7664,N_7556,N_7449);
and U7665 (N_7665,N_7515,N_7446);
nor U7666 (N_7666,N_7540,N_7444);
and U7667 (N_7667,N_7442,N_7558);
or U7668 (N_7668,N_7435,N_7461);
and U7669 (N_7669,N_7418,N_7464);
xnor U7670 (N_7670,N_7467,N_7421);
or U7671 (N_7671,N_7504,N_7560);
nor U7672 (N_7672,N_7565,N_7533);
nand U7673 (N_7673,N_7517,N_7494);
and U7674 (N_7674,N_7596,N_7597);
nor U7675 (N_7675,N_7415,N_7507);
nand U7676 (N_7676,N_7462,N_7426);
nor U7677 (N_7677,N_7575,N_7539);
and U7678 (N_7678,N_7505,N_7403);
nor U7679 (N_7679,N_7566,N_7537);
and U7680 (N_7680,N_7544,N_7497);
and U7681 (N_7681,N_7428,N_7430);
nand U7682 (N_7682,N_7546,N_7440);
nor U7683 (N_7683,N_7448,N_7416);
or U7684 (N_7684,N_7451,N_7473);
nand U7685 (N_7685,N_7582,N_7485);
and U7686 (N_7686,N_7500,N_7474);
nand U7687 (N_7687,N_7412,N_7510);
nand U7688 (N_7688,N_7514,N_7511);
or U7689 (N_7689,N_7478,N_7525);
and U7690 (N_7690,N_7526,N_7585);
or U7691 (N_7691,N_7574,N_7518);
or U7692 (N_7692,N_7522,N_7408);
nor U7693 (N_7693,N_7419,N_7532);
and U7694 (N_7694,N_7489,N_7553);
or U7695 (N_7695,N_7570,N_7429);
and U7696 (N_7696,N_7562,N_7479);
nand U7697 (N_7697,N_7508,N_7453);
and U7698 (N_7698,N_7437,N_7529);
or U7699 (N_7699,N_7543,N_7503);
or U7700 (N_7700,N_7548,N_7443);
and U7701 (N_7701,N_7516,N_7459);
nor U7702 (N_7702,N_7555,N_7530);
nor U7703 (N_7703,N_7460,N_7573);
and U7704 (N_7704,N_7457,N_7493);
or U7705 (N_7705,N_7593,N_7416);
or U7706 (N_7706,N_7565,N_7590);
and U7707 (N_7707,N_7577,N_7549);
and U7708 (N_7708,N_7441,N_7502);
or U7709 (N_7709,N_7584,N_7437);
or U7710 (N_7710,N_7491,N_7416);
nand U7711 (N_7711,N_7455,N_7485);
nand U7712 (N_7712,N_7444,N_7564);
nand U7713 (N_7713,N_7531,N_7564);
nor U7714 (N_7714,N_7573,N_7563);
nand U7715 (N_7715,N_7588,N_7483);
or U7716 (N_7716,N_7454,N_7569);
nand U7717 (N_7717,N_7457,N_7414);
nand U7718 (N_7718,N_7455,N_7446);
nand U7719 (N_7719,N_7426,N_7535);
nand U7720 (N_7720,N_7445,N_7559);
or U7721 (N_7721,N_7415,N_7474);
nand U7722 (N_7722,N_7561,N_7455);
nor U7723 (N_7723,N_7472,N_7444);
nor U7724 (N_7724,N_7430,N_7461);
nand U7725 (N_7725,N_7411,N_7461);
nand U7726 (N_7726,N_7408,N_7594);
nor U7727 (N_7727,N_7531,N_7435);
and U7728 (N_7728,N_7477,N_7498);
and U7729 (N_7729,N_7565,N_7486);
nand U7730 (N_7730,N_7582,N_7523);
nand U7731 (N_7731,N_7405,N_7463);
and U7732 (N_7732,N_7448,N_7406);
or U7733 (N_7733,N_7558,N_7445);
and U7734 (N_7734,N_7400,N_7498);
and U7735 (N_7735,N_7435,N_7595);
and U7736 (N_7736,N_7450,N_7425);
nor U7737 (N_7737,N_7528,N_7594);
nor U7738 (N_7738,N_7580,N_7474);
and U7739 (N_7739,N_7565,N_7422);
or U7740 (N_7740,N_7516,N_7453);
nand U7741 (N_7741,N_7589,N_7547);
nor U7742 (N_7742,N_7429,N_7405);
and U7743 (N_7743,N_7498,N_7453);
or U7744 (N_7744,N_7424,N_7594);
nor U7745 (N_7745,N_7480,N_7554);
or U7746 (N_7746,N_7586,N_7401);
and U7747 (N_7747,N_7466,N_7412);
and U7748 (N_7748,N_7461,N_7482);
or U7749 (N_7749,N_7562,N_7547);
nor U7750 (N_7750,N_7597,N_7428);
and U7751 (N_7751,N_7520,N_7433);
or U7752 (N_7752,N_7550,N_7406);
or U7753 (N_7753,N_7528,N_7400);
nor U7754 (N_7754,N_7550,N_7403);
and U7755 (N_7755,N_7571,N_7438);
or U7756 (N_7756,N_7544,N_7589);
nand U7757 (N_7757,N_7479,N_7410);
nand U7758 (N_7758,N_7470,N_7587);
or U7759 (N_7759,N_7449,N_7585);
xor U7760 (N_7760,N_7563,N_7405);
and U7761 (N_7761,N_7407,N_7509);
and U7762 (N_7762,N_7465,N_7469);
nor U7763 (N_7763,N_7443,N_7582);
or U7764 (N_7764,N_7508,N_7516);
or U7765 (N_7765,N_7586,N_7460);
and U7766 (N_7766,N_7531,N_7488);
nor U7767 (N_7767,N_7511,N_7401);
or U7768 (N_7768,N_7555,N_7474);
or U7769 (N_7769,N_7457,N_7496);
or U7770 (N_7770,N_7519,N_7572);
and U7771 (N_7771,N_7551,N_7557);
nor U7772 (N_7772,N_7415,N_7524);
and U7773 (N_7773,N_7448,N_7570);
and U7774 (N_7774,N_7427,N_7413);
nor U7775 (N_7775,N_7580,N_7539);
nand U7776 (N_7776,N_7568,N_7496);
and U7777 (N_7777,N_7407,N_7455);
nor U7778 (N_7778,N_7557,N_7412);
nor U7779 (N_7779,N_7408,N_7525);
nand U7780 (N_7780,N_7521,N_7409);
nor U7781 (N_7781,N_7585,N_7470);
nor U7782 (N_7782,N_7519,N_7443);
or U7783 (N_7783,N_7561,N_7519);
xnor U7784 (N_7784,N_7468,N_7512);
and U7785 (N_7785,N_7418,N_7557);
nand U7786 (N_7786,N_7475,N_7479);
nand U7787 (N_7787,N_7527,N_7417);
and U7788 (N_7788,N_7430,N_7516);
or U7789 (N_7789,N_7422,N_7489);
nor U7790 (N_7790,N_7560,N_7576);
and U7791 (N_7791,N_7481,N_7578);
or U7792 (N_7792,N_7414,N_7477);
nand U7793 (N_7793,N_7576,N_7441);
and U7794 (N_7794,N_7416,N_7479);
nor U7795 (N_7795,N_7468,N_7501);
xor U7796 (N_7796,N_7587,N_7536);
and U7797 (N_7797,N_7556,N_7406);
nor U7798 (N_7798,N_7543,N_7505);
nand U7799 (N_7799,N_7558,N_7425);
or U7800 (N_7800,N_7715,N_7682);
nand U7801 (N_7801,N_7636,N_7612);
nor U7802 (N_7802,N_7649,N_7655);
nor U7803 (N_7803,N_7773,N_7621);
and U7804 (N_7804,N_7762,N_7728);
and U7805 (N_7805,N_7693,N_7615);
and U7806 (N_7806,N_7774,N_7677);
and U7807 (N_7807,N_7635,N_7729);
nand U7808 (N_7808,N_7724,N_7647);
nor U7809 (N_7809,N_7617,N_7618);
or U7810 (N_7810,N_7777,N_7748);
nand U7811 (N_7811,N_7699,N_7720);
and U7812 (N_7812,N_7620,N_7661);
or U7813 (N_7813,N_7611,N_7739);
nor U7814 (N_7814,N_7731,N_7639);
or U7815 (N_7815,N_7722,N_7723);
nand U7816 (N_7816,N_7709,N_7660);
or U7817 (N_7817,N_7604,N_7633);
or U7818 (N_7818,N_7792,N_7798);
or U7819 (N_7819,N_7634,N_7643);
and U7820 (N_7820,N_7678,N_7745);
nand U7821 (N_7821,N_7741,N_7706);
nand U7822 (N_7822,N_7669,N_7656);
or U7823 (N_7823,N_7607,N_7640);
nand U7824 (N_7824,N_7679,N_7630);
and U7825 (N_7825,N_7718,N_7740);
nor U7826 (N_7826,N_7689,N_7673);
nor U7827 (N_7827,N_7624,N_7702);
and U7828 (N_7828,N_7717,N_7714);
or U7829 (N_7829,N_7788,N_7700);
nor U7830 (N_7830,N_7737,N_7756);
or U7831 (N_7831,N_7734,N_7659);
nor U7832 (N_7832,N_7685,N_7730);
xnor U7833 (N_7833,N_7632,N_7654);
nor U7834 (N_7834,N_7776,N_7795);
nor U7835 (N_7835,N_7683,N_7675);
nor U7836 (N_7836,N_7692,N_7786);
and U7837 (N_7837,N_7772,N_7628);
and U7838 (N_7838,N_7753,N_7658);
and U7839 (N_7839,N_7780,N_7645);
nor U7840 (N_7840,N_7775,N_7727);
and U7841 (N_7841,N_7705,N_7627);
nor U7842 (N_7842,N_7642,N_7725);
or U7843 (N_7843,N_7783,N_7694);
or U7844 (N_7844,N_7600,N_7614);
and U7845 (N_7845,N_7619,N_7603);
and U7846 (N_7846,N_7657,N_7651);
nor U7847 (N_7847,N_7668,N_7767);
nand U7848 (N_7848,N_7785,N_7662);
nor U7849 (N_7849,N_7613,N_7744);
and U7850 (N_7850,N_7755,N_7703);
or U7851 (N_7851,N_7644,N_7758);
or U7852 (N_7852,N_7759,N_7770);
and U7853 (N_7853,N_7710,N_7707);
nand U7854 (N_7854,N_7697,N_7719);
xnor U7855 (N_7855,N_7738,N_7631);
or U7856 (N_7856,N_7698,N_7757);
and U7857 (N_7857,N_7778,N_7754);
nand U7858 (N_7858,N_7799,N_7680);
nand U7859 (N_7859,N_7793,N_7676);
nor U7860 (N_7860,N_7794,N_7747);
nor U7861 (N_7861,N_7608,N_7666);
nor U7862 (N_7862,N_7711,N_7781);
nand U7863 (N_7863,N_7746,N_7771);
and U7864 (N_7864,N_7695,N_7687);
nand U7865 (N_7865,N_7686,N_7672);
nand U7866 (N_7866,N_7779,N_7641);
or U7867 (N_7867,N_7696,N_7787);
and U7868 (N_7868,N_7601,N_7796);
and U7869 (N_7869,N_7688,N_7742);
and U7870 (N_7870,N_7623,N_7726);
nor U7871 (N_7871,N_7629,N_7768);
xnor U7872 (N_7872,N_7721,N_7605);
or U7873 (N_7873,N_7766,N_7610);
or U7874 (N_7874,N_7681,N_7789);
nor U7875 (N_7875,N_7797,N_7791);
or U7876 (N_7876,N_7761,N_7637);
and U7877 (N_7877,N_7749,N_7712);
and U7878 (N_7878,N_7790,N_7670);
and U7879 (N_7879,N_7716,N_7732);
and U7880 (N_7880,N_7704,N_7650);
nand U7881 (N_7881,N_7602,N_7648);
or U7882 (N_7882,N_7606,N_7691);
and U7883 (N_7883,N_7733,N_7701);
nor U7884 (N_7884,N_7663,N_7713);
nor U7885 (N_7885,N_7616,N_7674);
or U7886 (N_7886,N_7743,N_7646);
and U7887 (N_7887,N_7622,N_7763);
nand U7888 (N_7888,N_7765,N_7667);
or U7889 (N_7889,N_7769,N_7626);
and U7890 (N_7890,N_7764,N_7784);
nand U7891 (N_7891,N_7735,N_7665);
xnor U7892 (N_7892,N_7736,N_7625);
nor U7893 (N_7893,N_7708,N_7664);
nand U7894 (N_7894,N_7638,N_7609);
or U7895 (N_7895,N_7684,N_7750);
nor U7896 (N_7896,N_7690,N_7782);
nand U7897 (N_7897,N_7652,N_7752);
or U7898 (N_7898,N_7760,N_7751);
and U7899 (N_7899,N_7653,N_7671);
or U7900 (N_7900,N_7744,N_7620);
and U7901 (N_7901,N_7758,N_7787);
nor U7902 (N_7902,N_7753,N_7608);
or U7903 (N_7903,N_7685,N_7775);
and U7904 (N_7904,N_7790,N_7693);
or U7905 (N_7905,N_7609,N_7793);
and U7906 (N_7906,N_7701,N_7661);
or U7907 (N_7907,N_7752,N_7700);
nor U7908 (N_7908,N_7758,N_7770);
nand U7909 (N_7909,N_7702,N_7674);
nor U7910 (N_7910,N_7789,N_7642);
nand U7911 (N_7911,N_7642,N_7684);
and U7912 (N_7912,N_7710,N_7668);
or U7913 (N_7913,N_7618,N_7683);
nor U7914 (N_7914,N_7660,N_7714);
and U7915 (N_7915,N_7755,N_7740);
nand U7916 (N_7916,N_7605,N_7734);
xnor U7917 (N_7917,N_7604,N_7614);
nand U7918 (N_7918,N_7768,N_7665);
nor U7919 (N_7919,N_7762,N_7709);
nor U7920 (N_7920,N_7614,N_7779);
or U7921 (N_7921,N_7697,N_7742);
or U7922 (N_7922,N_7627,N_7735);
nand U7923 (N_7923,N_7768,N_7654);
nand U7924 (N_7924,N_7773,N_7634);
and U7925 (N_7925,N_7699,N_7721);
nor U7926 (N_7926,N_7650,N_7786);
or U7927 (N_7927,N_7658,N_7644);
and U7928 (N_7928,N_7613,N_7683);
and U7929 (N_7929,N_7701,N_7790);
nor U7930 (N_7930,N_7787,N_7610);
xor U7931 (N_7931,N_7612,N_7799);
nand U7932 (N_7932,N_7657,N_7742);
nor U7933 (N_7933,N_7616,N_7712);
nand U7934 (N_7934,N_7754,N_7744);
nand U7935 (N_7935,N_7763,N_7683);
and U7936 (N_7936,N_7698,N_7735);
nand U7937 (N_7937,N_7652,N_7778);
nor U7938 (N_7938,N_7739,N_7620);
or U7939 (N_7939,N_7718,N_7792);
nand U7940 (N_7940,N_7640,N_7778);
and U7941 (N_7941,N_7619,N_7673);
or U7942 (N_7942,N_7714,N_7625);
nand U7943 (N_7943,N_7612,N_7760);
nand U7944 (N_7944,N_7619,N_7746);
and U7945 (N_7945,N_7675,N_7631);
nor U7946 (N_7946,N_7618,N_7766);
or U7947 (N_7947,N_7733,N_7728);
and U7948 (N_7948,N_7618,N_7781);
xnor U7949 (N_7949,N_7651,N_7690);
nand U7950 (N_7950,N_7635,N_7711);
nor U7951 (N_7951,N_7775,N_7669);
or U7952 (N_7952,N_7627,N_7604);
and U7953 (N_7953,N_7753,N_7638);
and U7954 (N_7954,N_7612,N_7679);
nor U7955 (N_7955,N_7734,N_7607);
or U7956 (N_7956,N_7738,N_7655);
nand U7957 (N_7957,N_7655,N_7634);
nand U7958 (N_7958,N_7633,N_7601);
nor U7959 (N_7959,N_7792,N_7781);
and U7960 (N_7960,N_7784,N_7642);
nor U7961 (N_7961,N_7735,N_7697);
or U7962 (N_7962,N_7710,N_7754);
nor U7963 (N_7963,N_7653,N_7650);
nand U7964 (N_7964,N_7786,N_7709);
nor U7965 (N_7965,N_7735,N_7769);
nand U7966 (N_7966,N_7733,N_7756);
and U7967 (N_7967,N_7701,N_7714);
or U7968 (N_7968,N_7659,N_7626);
nand U7969 (N_7969,N_7718,N_7691);
nor U7970 (N_7970,N_7661,N_7668);
nand U7971 (N_7971,N_7759,N_7786);
nor U7972 (N_7972,N_7702,N_7708);
and U7973 (N_7973,N_7737,N_7785);
and U7974 (N_7974,N_7745,N_7712);
nand U7975 (N_7975,N_7734,N_7783);
and U7976 (N_7976,N_7690,N_7605);
and U7977 (N_7977,N_7788,N_7793);
or U7978 (N_7978,N_7623,N_7727);
nand U7979 (N_7979,N_7709,N_7722);
or U7980 (N_7980,N_7696,N_7797);
nor U7981 (N_7981,N_7797,N_7604);
nand U7982 (N_7982,N_7711,N_7777);
nand U7983 (N_7983,N_7610,N_7757);
nor U7984 (N_7984,N_7778,N_7647);
or U7985 (N_7985,N_7798,N_7764);
and U7986 (N_7986,N_7695,N_7705);
xor U7987 (N_7987,N_7603,N_7715);
nand U7988 (N_7988,N_7716,N_7630);
or U7989 (N_7989,N_7793,N_7705);
and U7990 (N_7990,N_7685,N_7751);
nand U7991 (N_7991,N_7653,N_7621);
nor U7992 (N_7992,N_7780,N_7726);
nor U7993 (N_7993,N_7668,N_7728);
or U7994 (N_7994,N_7603,N_7712);
nand U7995 (N_7995,N_7735,N_7604);
or U7996 (N_7996,N_7791,N_7654);
nand U7997 (N_7997,N_7724,N_7753);
nand U7998 (N_7998,N_7700,N_7699);
nand U7999 (N_7999,N_7795,N_7723);
or U8000 (N_8000,N_7936,N_7873);
nand U8001 (N_8001,N_7905,N_7878);
and U8002 (N_8002,N_7982,N_7824);
and U8003 (N_8003,N_7972,N_7814);
and U8004 (N_8004,N_7973,N_7937);
nand U8005 (N_8005,N_7801,N_7996);
or U8006 (N_8006,N_7963,N_7828);
nand U8007 (N_8007,N_7855,N_7871);
nand U8008 (N_8008,N_7991,N_7822);
nor U8009 (N_8009,N_7933,N_7889);
nor U8010 (N_8010,N_7934,N_7805);
nor U8011 (N_8011,N_7912,N_7882);
nor U8012 (N_8012,N_7880,N_7993);
and U8013 (N_8013,N_7924,N_7998);
nand U8014 (N_8014,N_7988,N_7914);
and U8015 (N_8015,N_7955,N_7960);
nand U8016 (N_8016,N_7913,N_7927);
nor U8017 (N_8017,N_7815,N_7986);
and U8018 (N_8018,N_7968,N_7894);
and U8019 (N_8019,N_7921,N_7954);
nor U8020 (N_8020,N_7979,N_7848);
nand U8021 (N_8021,N_7854,N_7881);
nand U8022 (N_8022,N_7803,N_7809);
or U8023 (N_8023,N_7964,N_7910);
nand U8024 (N_8024,N_7835,N_7990);
nor U8025 (N_8025,N_7813,N_7941);
or U8026 (N_8026,N_7950,N_7891);
and U8027 (N_8027,N_7892,N_7944);
and U8028 (N_8028,N_7920,N_7845);
and U8029 (N_8029,N_7800,N_7853);
nand U8030 (N_8030,N_7841,N_7981);
or U8031 (N_8031,N_7816,N_7829);
or U8032 (N_8032,N_7872,N_7930);
and U8033 (N_8033,N_7948,N_7919);
nor U8034 (N_8034,N_7931,N_7818);
and U8035 (N_8035,N_7947,N_7918);
or U8036 (N_8036,N_7866,N_7938);
nor U8037 (N_8037,N_7808,N_7825);
nand U8038 (N_8038,N_7893,N_7847);
or U8039 (N_8039,N_7952,N_7939);
nand U8040 (N_8040,N_7958,N_7884);
nor U8041 (N_8041,N_7940,N_7932);
nor U8042 (N_8042,N_7838,N_7874);
or U8043 (N_8043,N_7886,N_7899);
or U8044 (N_8044,N_7807,N_7970);
and U8045 (N_8045,N_7978,N_7851);
or U8046 (N_8046,N_7975,N_7820);
nor U8047 (N_8047,N_7804,N_7868);
nand U8048 (N_8048,N_7915,N_7840);
and U8049 (N_8049,N_7846,N_7984);
nand U8050 (N_8050,N_7879,N_7834);
or U8051 (N_8051,N_7830,N_7976);
nor U8052 (N_8052,N_7904,N_7859);
nand U8053 (N_8053,N_7965,N_7849);
or U8054 (N_8054,N_7860,N_7877);
nand U8055 (N_8055,N_7898,N_7900);
and U8056 (N_8056,N_7819,N_7967);
and U8057 (N_8057,N_7856,N_7917);
and U8058 (N_8058,N_7928,N_7911);
nor U8059 (N_8059,N_7895,N_7844);
or U8060 (N_8060,N_7858,N_7926);
and U8061 (N_8061,N_7863,N_7922);
and U8062 (N_8062,N_7909,N_7962);
nand U8063 (N_8063,N_7802,N_7806);
and U8064 (N_8064,N_7957,N_7974);
and U8065 (N_8065,N_7817,N_7929);
nand U8066 (N_8066,N_7987,N_7945);
nor U8067 (N_8067,N_7997,N_7999);
and U8068 (N_8068,N_7923,N_7843);
xnor U8069 (N_8069,N_7943,N_7935);
or U8070 (N_8070,N_7980,N_7861);
nand U8071 (N_8071,N_7875,N_7907);
and U8072 (N_8072,N_7869,N_7865);
nor U8073 (N_8073,N_7896,N_7983);
nand U8074 (N_8074,N_7857,N_7885);
and U8075 (N_8075,N_7811,N_7836);
and U8076 (N_8076,N_7832,N_7810);
xnor U8077 (N_8077,N_7827,N_7951);
and U8078 (N_8078,N_7949,N_7902);
and U8079 (N_8079,N_7903,N_7812);
or U8080 (N_8080,N_7916,N_7969);
and U8081 (N_8081,N_7883,N_7897);
or U8082 (N_8082,N_7833,N_7995);
nand U8083 (N_8083,N_7946,N_7867);
xor U8084 (N_8084,N_7831,N_7966);
nand U8085 (N_8085,N_7842,N_7959);
nand U8086 (N_8086,N_7956,N_7864);
or U8087 (N_8087,N_7901,N_7906);
nor U8088 (N_8088,N_7887,N_7826);
nand U8089 (N_8089,N_7852,N_7961);
and U8090 (N_8090,N_7989,N_7890);
nor U8091 (N_8091,N_7837,N_7994);
or U8092 (N_8092,N_7985,N_7977);
or U8093 (N_8093,N_7953,N_7992);
nand U8094 (N_8094,N_7876,N_7823);
or U8095 (N_8095,N_7870,N_7850);
nor U8096 (N_8096,N_7839,N_7862);
nor U8097 (N_8097,N_7888,N_7908);
xnor U8098 (N_8098,N_7821,N_7925);
or U8099 (N_8099,N_7942,N_7971);
and U8100 (N_8100,N_7920,N_7823);
nor U8101 (N_8101,N_7912,N_7842);
or U8102 (N_8102,N_7974,N_7804);
nand U8103 (N_8103,N_7873,N_7802);
and U8104 (N_8104,N_7912,N_7946);
or U8105 (N_8105,N_7890,N_7865);
nor U8106 (N_8106,N_7954,N_7891);
nor U8107 (N_8107,N_7827,N_7891);
nand U8108 (N_8108,N_7877,N_7834);
nor U8109 (N_8109,N_7934,N_7826);
and U8110 (N_8110,N_7816,N_7911);
nand U8111 (N_8111,N_7956,N_7878);
nand U8112 (N_8112,N_7947,N_7952);
nand U8113 (N_8113,N_7955,N_7949);
or U8114 (N_8114,N_7832,N_7835);
or U8115 (N_8115,N_7833,N_7908);
nor U8116 (N_8116,N_7834,N_7880);
nor U8117 (N_8117,N_7922,N_7881);
nand U8118 (N_8118,N_7976,N_7902);
or U8119 (N_8119,N_7878,N_7888);
or U8120 (N_8120,N_7844,N_7811);
or U8121 (N_8121,N_7998,N_7811);
nand U8122 (N_8122,N_7806,N_7903);
nor U8123 (N_8123,N_7832,N_7842);
nor U8124 (N_8124,N_7977,N_7810);
nor U8125 (N_8125,N_7828,N_7827);
nand U8126 (N_8126,N_7998,N_7832);
and U8127 (N_8127,N_7906,N_7892);
or U8128 (N_8128,N_7939,N_7860);
nand U8129 (N_8129,N_7898,N_7822);
and U8130 (N_8130,N_7825,N_7853);
and U8131 (N_8131,N_7993,N_7924);
nand U8132 (N_8132,N_7839,N_7905);
nand U8133 (N_8133,N_7934,N_7979);
or U8134 (N_8134,N_7942,N_7928);
xnor U8135 (N_8135,N_7964,N_7968);
and U8136 (N_8136,N_7960,N_7896);
nor U8137 (N_8137,N_7805,N_7970);
or U8138 (N_8138,N_7940,N_7935);
nand U8139 (N_8139,N_7951,N_7886);
and U8140 (N_8140,N_7908,N_7877);
nand U8141 (N_8141,N_7857,N_7851);
and U8142 (N_8142,N_7970,N_7800);
and U8143 (N_8143,N_7863,N_7804);
or U8144 (N_8144,N_7814,N_7986);
or U8145 (N_8145,N_7854,N_7857);
nand U8146 (N_8146,N_7953,N_7869);
nor U8147 (N_8147,N_7882,N_7891);
nand U8148 (N_8148,N_7840,N_7997);
and U8149 (N_8149,N_7913,N_7809);
nand U8150 (N_8150,N_7982,N_7894);
or U8151 (N_8151,N_7830,N_7961);
nor U8152 (N_8152,N_7981,N_7902);
nor U8153 (N_8153,N_7875,N_7848);
and U8154 (N_8154,N_7843,N_7848);
and U8155 (N_8155,N_7861,N_7819);
and U8156 (N_8156,N_7891,N_7824);
nand U8157 (N_8157,N_7974,N_7809);
or U8158 (N_8158,N_7890,N_7807);
or U8159 (N_8159,N_7964,N_7838);
or U8160 (N_8160,N_7913,N_7933);
nor U8161 (N_8161,N_7976,N_7908);
nand U8162 (N_8162,N_7829,N_7971);
nand U8163 (N_8163,N_7998,N_7803);
and U8164 (N_8164,N_7987,N_7927);
or U8165 (N_8165,N_7929,N_7912);
nand U8166 (N_8166,N_7832,N_7930);
and U8167 (N_8167,N_7935,N_7988);
and U8168 (N_8168,N_7987,N_7856);
or U8169 (N_8169,N_7915,N_7819);
nor U8170 (N_8170,N_7889,N_7879);
nand U8171 (N_8171,N_7966,N_7860);
nor U8172 (N_8172,N_7992,N_7894);
and U8173 (N_8173,N_7942,N_7886);
nor U8174 (N_8174,N_7812,N_7943);
nor U8175 (N_8175,N_7977,N_7815);
nor U8176 (N_8176,N_7938,N_7923);
xor U8177 (N_8177,N_7853,N_7996);
nand U8178 (N_8178,N_7893,N_7997);
or U8179 (N_8179,N_7855,N_7971);
and U8180 (N_8180,N_7847,N_7924);
nand U8181 (N_8181,N_7893,N_7983);
or U8182 (N_8182,N_7975,N_7863);
xnor U8183 (N_8183,N_7831,N_7947);
nor U8184 (N_8184,N_7997,N_7989);
nand U8185 (N_8185,N_7814,N_7849);
or U8186 (N_8186,N_7976,N_7805);
and U8187 (N_8187,N_7823,N_7841);
and U8188 (N_8188,N_7997,N_7907);
nor U8189 (N_8189,N_7866,N_7913);
nand U8190 (N_8190,N_7971,N_7949);
and U8191 (N_8191,N_7982,N_7890);
or U8192 (N_8192,N_7804,N_7858);
nor U8193 (N_8193,N_7864,N_7910);
or U8194 (N_8194,N_7829,N_7951);
and U8195 (N_8195,N_7902,N_7991);
nand U8196 (N_8196,N_7821,N_7979);
nand U8197 (N_8197,N_7865,N_7994);
nor U8198 (N_8198,N_7948,N_7812);
nor U8199 (N_8199,N_7911,N_7848);
nand U8200 (N_8200,N_8036,N_8168);
nand U8201 (N_8201,N_8189,N_8136);
nor U8202 (N_8202,N_8092,N_8040);
nand U8203 (N_8203,N_8021,N_8039);
nor U8204 (N_8204,N_8105,N_8093);
nor U8205 (N_8205,N_8184,N_8109);
and U8206 (N_8206,N_8160,N_8002);
nand U8207 (N_8207,N_8150,N_8033);
nor U8208 (N_8208,N_8190,N_8030);
and U8209 (N_8209,N_8023,N_8082);
nor U8210 (N_8210,N_8078,N_8034);
and U8211 (N_8211,N_8100,N_8108);
nand U8212 (N_8212,N_8120,N_8015);
nand U8213 (N_8213,N_8157,N_8140);
nand U8214 (N_8214,N_8111,N_8080);
or U8215 (N_8215,N_8001,N_8075);
and U8216 (N_8216,N_8122,N_8037);
xor U8217 (N_8217,N_8161,N_8081);
and U8218 (N_8218,N_8155,N_8031);
nand U8219 (N_8219,N_8144,N_8139);
nor U8220 (N_8220,N_8102,N_8091);
nor U8221 (N_8221,N_8097,N_8053);
xor U8222 (N_8222,N_8019,N_8165);
nand U8223 (N_8223,N_8123,N_8198);
nand U8224 (N_8224,N_8171,N_8055);
nand U8225 (N_8225,N_8049,N_8059);
nor U8226 (N_8226,N_8012,N_8096);
nand U8227 (N_8227,N_8045,N_8043);
and U8228 (N_8228,N_8058,N_8011);
nand U8229 (N_8229,N_8000,N_8152);
nor U8230 (N_8230,N_8115,N_8106);
and U8231 (N_8231,N_8065,N_8048);
nand U8232 (N_8232,N_8170,N_8186);
and U8233 (N_8233,N_8143,N_8197);
xor U8234 (N_8234,N_8141,N_8131);
nor U8235 (N_8235,N_8026,N_8164);
nand U8236 (N_8236,N_8013,N_8029);
nor U8237 (N_8237,N_8192,N_8147);
or U8238 (N_8238,N_8191,N_8158);
nand U8239 (N_8239,N_8074,N_8020);
or U8240 (N_8240,N_8159,N_8130);
or U8241 (N_8241,N_8077,N_8128);
nand U8242 (N_8242,N_8148,N_8187);
nand U8243 (N_8243,N_8032,N_8028);
nor U8244 (N_8244,N_8016,N_8008);
and U8245 (N_8245,N_8063,N_8174);
nand U8246 (N_8246,N_8090,N_8062);
or U8247 (N_8247,N_8182,N_8044);
and U8248 (N_8248,N_8151,N_8088);
nor U8249 (N_8249,N_8064,N_8104);
or U8250 (N_8250,N_8134,N_8129);
nand U8251 (N_8251,N_8126,N_8079);
nor U8252 (N_8252,N_8193,N_8073);
nor U8253 (N_8253,N_8010,N_8017);
and U8254 (N_8254,N_8135,N_8112);
nand U8255 (N_8255,N_8173,N_8180);
or U8256 (N_8256,N_8132,N_8099);
nand U8257 (N_8257,N_8114,N_8145);
and U8258 (N_8258,N_8041,N_8098);
nor U8259 (N_8259,N_8133,N_8195);
nand U8260 (N_8260,N_8118,N_8163);
nor U8261 (N_8261,N_8154,N_8061);
nand U8262 (N_8262,N_8054,N_8072);
nand U8263 (N_8263,N_8137,N_8175);
or U8264 (N_8264,N_8003,N_8085);
or U8265 (N_8265,N_8027,N_8076);
and U8266 (N_8266,N_8107,N_8038);
or U8267 (N_8267,N_8156,N_8167);
or U8268 (N_8268,N_8014,N_8095);
or U8269 (N_8269,N_8060,N_8117);
nor U8270 (N_8270,N_8005,N_8166);
nor U8271 (N_8271,N_8046,N_8089);
or U8272 (N_8272,N_8070,N_8185);
nand U8273 (N_8273,N_8125,N_8194);
and U8274 (N_8274,N_8181,N_8047);
and U8275 (N_8275,N_8086,N_8068);
and U8276 (N_8276,N_8103,N_8101);
or U8277 (N_8277,N_8178,N_8177);
or U8278 (N_8278,N_8024,N_8127);
nor U8279 (N_8279,N_8050,N_8196);
or U8280 (N_8280,N_8067,N_8149);
nand U8281 (N_8281,N_8018,N_8022);
nand U8282 (N_8282,N_8042,N_8124);
nor U8283 (N_8283,N_8084,N_8113);
and U8284 (N_8284,N_8138,N_8110);
nor U8285 (N_8285,N_8057,N_8052);
nand U8286 (N_8286,N_8116,N_8119);
or U8287 (N_8287,N_8051,N_8176);
and U8288 (N_8288,N_8007,N_8162);
nand U8289 (N_8289,N_8035,N_8153);
nand U8290 (N_8290,N_8083,N_8172);
and U8291 (N_8291,N_8087,N_8183);
and U8292 (N_8292,N_8069,N_8056);
nor U8293 (N_8293,N_8066,N_8009);
or U8294 (N_8294,N_8199,N_8004);
nand U8295 (N_8295,N_8121,N_8071);
or U8296 (N_8296,N_8006,N_8142);
nand U8297 (N_8297,N_8169,N_8146);
or U8298 (N_8298,N_8094,N_8179);
or U8299 (N_8299,N_8188,N_8025);
nand U8300 (N_8300,N_8042,N_8083);
or U8301 (N_8301,N_8070,N_8142);
and U8302 (N_8302,N_8050,N_8054);
and U8303 (N_8303,N_8148,N_8118);
nor U8304 (N_8304,N_8016,N_8120);
nor U8305 (N_8305,N_8162,N_8108);
or U8306 (N_8306,N_8009,N_8167);
and U8307 (N_8307,N_8110,N_8046);
and U8308 (N_8308,N_8147,N_8072);
nand U8309 (N_8309,N_8117,N_8180);
nor U8310 (N_8310,N_8182,N_8143);
or U8311 (N_8311,N_8139,N_8041);
and U8312 (N_8312,N_8189,N_8135);
nor U8313 (N_8313,N_8172,N_8189);
or U8314 (N_8314,N_8149,N_8085);
or U8315 (N_8315,N_8171,N_8120);
or U8316 (N_8316,N_8189,N_8004);
nor U8317 (N_8317,N_8123,N_8069);
nor U8318 (N_8318,N_8065,N_8164);
nor U8319 (N_8319,N_8053,N_8119);
and U8320 (N_8320,N_8039,N_8189);
nand U8321 (N_8321,N_8116,N_8139);
or U8322 (N_8322,N_8004,N_8184);
and U8323 (N_8323,N_8148,N_8015);
or U8324 (N_8324,N_8070,N_8096);
and U8325 (N_8325,N_8111,N_8175);
and U8326 (N_8326,N_8065,N_8019);
nand U8327 (N_8327,N_8019,N_8155);
or U8328 (N_8328,N_8113,N_8003);
or U8329 (N_8329,N_8008,N_8000);
nand U8330 (N_8330,N_8108,N_8110);
or U8331 (N_8331,N_8073,N_8144);
nor U8332 (N_8332,N_8160,N_8011);
nor U8333 (N_8333,N_8044,N_8108);
nor U8334 (N_8334,N_8193,N_8150);
nor U8335 (N_8335,N_8125,N_8076);
nand U8336 (N_8336,N_8096,N_8158);
nand U8337 (N_8337,N_8011,N_8051);
nor U8338 (N_8338,N_8070,N_8182);
nor U8339 (N_8339,N_8097,N_8108);
nand U8340 (N_8340,N_8004,N_8033);
nand U8341 (N_8341,N_8112,N_8111);
or U8342 (N_8342,N_8098,N_8027);
and U8343 (N_8343,N_8143,N_8089);
nor U8344 (N_8344,N_8155,N_8193);
or U8345 (N_8345,N_8165,N_8046);
nand U8346 (N_8346,N_8077,N_8111);
and U8347 (N_8347,N_8153,N_8189);
and U8348 (N_8348,N_8067,N_8123);
nand U8349 (N_8349,N_8198,N_8046);
nor U8350 (N_8350,N_8067,N_8091);
and U8351 (N_8351,N_8187,N_8073);
nor U8352 (N_8352,N_8176,N_8082);
and U8353 (N_8353,N_8097,N_8010);
nand U8354 (N_8354,N_8069,N_8091);
or U8355 (N_8355,N_8068,N_8107);
nor U8356 (N_8356,N_8194,N_8064);
nor U8357 (N_8357,N_8128,N_8155);
and U8358 (N_8358,N_8104,N_8121);
and U8359 (N_8359,N_8000,N_8039);
and U8360 (N_8360,N_8132,N_8155);
nand U8361 (N_8361,N_8148,N_8120);
or U8362 (N_8362,N_8025,N_8191);
and U8363 (N_8363,N_8143,N_8172);
or U8364 (N_8364,N_8093,N_8127);
and U8365 (N_8365,N_8050,N_8074);
nor U8366 (N_8366,N_8159,N_8116);
and U8367 (N_8367,N_8076,N_8130);
nor U8368 (N_8368,N_8079,N_8004);
and U8369 (N_8369,N_8025,N_8060);
or U8370 (N_8370,N_8078,N_8018);
nor U8371 (N_8371,N_8005,N_8090);
or U8372 (N_8372,N_8186,N_8149);
nor U8373 (N_8373,N_8177,N_8135);
nor U8374 (N_8374,N_8076,N_8011);
or U8375 (N_8375,N_8040,N_8120);
or U8376 (N_8376,N_8028,N_8071);
or U8377 (N_8377,N_8027,N_8179);
and U8378 (N_8378,N_8027,N_8100);
or U8379 (N_8379,N_8070,N_8043);
or U8380 (N_8380,N_8072,N_8099);
nor U8381 (N_8381,N_8091,N_8198);
or U8382 (N_8382,N_8062,N_8183);
nor U8383 (N_8383,N_8091,N_8006);
or U8384 (N_8384,N_8035,N_8050);
nor U8385 (N_8385,N_8199,N_8019);
or U8386 (N_8386,N_8137,N_8150);
nand U8387 (N_8387,N_8034,N_8147);
or U8388 (N_8388,N_8083,N_8147);
and U8389 (N_8389,N_8128,N_8030);
and U8390 (N_8390,N_8194,N_8101);
xnor U8391 (N_8391,N_8147,N_8111);
or U8392 (N_8392,N_8193,N_8035);
or U8393 (N_8393,N_8186,N_8028);
or U8394 (N_8394,N_8124,N_8035);
nand U8395 (N_8395,N_8193,N_8129);
nor U8396 (N_8396,N_8000,N_8070);
nand U8397 (N_8397,N_8184,N_8091);
nor U8398 (N_8398,N_8195,N_8156);
or U8399 (N_8399,N_8170,N_8011);
nand U8400 (N_8400,N_8345,N_8331);
and U8401 (N_8401,N_8275,N_8232);
nand U8402 (N_8402,N_8298,N_8336);
and U8403 (N_8403,N_8216,N_8254);
nor U8404 (N_8404,N_8268,N_8226);
and U8405 (N_8405,N_8330,N_8387);
or U8406 (N_8406,N_8368,N_8349);
or U8407 (N_8407,N_8220,N_8346);
nor U8408 (N_8408,N_8397,N_8255);
or U8409 (N_8409,N_8308,N_8269);
and U8410 (N_8410,N_8360,N_8257);
or U8411 (N_8411,N_8295,N_8393);
or U8412 (N_8412,N_8311,N_8247);
nand U8413 (N_8413,N_8371,N_8392);
nand U8414 (N_8414,N_8384,N_8217);
nand U8415 (N_8415,N_8201,N_8294);
and U8416 (N_8416,N_8376,N_8279);
and U8417 (N_8417,N_8227,N_8251);
or U8418 (N_8418,N_8272,N_8240);
nand U8419 (N_8419,N_8385,N_8256);
or U8420 (N_8420,N_8249,N_8318);
and U8421 (N_8421,N_8396,N_8323);
nand U8422 (N_8422,N_8369,N_8389);
nor U8423 (N_8423,N_8315,N_8304);
and U8424 (N_8424,N_8306,N_8309);
or U8425 (N_8425,N_8242,N_8341);
and U8426 (N_8426,N_8332,N_8348);
or U8427 (N_8427,N_8354,N_8300);
or U8428 (N_8428,N_8329,N_8244);
xor U8429 (N_8429,N_8322,N_8290);
nor U8430 (N_8430,N_8278,N_8394);
nand U8431 (N_8431,N_8381,N_8233);
nor U8432 (N_8432,N_8359,N_8250);
and U8433 (N_8433,N_8342,N_8337);
and U8434 (N_8434,N_8222,N_8386);
and U8435 (N_8435,N_8324,N_8355);
nand U8436 (N_8436,N_8303,N_8230);
xnor U8437 (N_8437,N_8204,N_8362);
or U8438 (N_8438,N_8237,N_8307);
and U8439 (N_8439,N_8320,N_8357);
and U8440 (N_8440,N_8245,N_8292);
or U8441 (N_8441,N_8350,N_8258);
nor U8442 (N_8442,N_8352,N_8356);
or U8443 (N_8443,N_8202,N_8338);
nor U8444 (N_8444,N_8297,N_8388);
nand U8445 (N_8445,N_8317,N_8313);
or U8446 (N_8446,N_8344,N_8213);
or U8447 (N_8447,N_8286,N_8312);
nand U8448 (N_8448,N_8273,N_8373);
xor U8449 (N_8449,N_8229,N_8235);
nor U8450 (N_8450,N_8366,N_8333);
or U8451 (N_8451,N_8364,N_8372);
nor U8452 (N_8452,N_8353,N_8200);
nand U8453 (N_8453,N_8289,N_8215);
and U8454 (N_8454,N_8228,N_8283);
nand U8455 (N_8455,N_8363,N_8383);
nand U8456 (N_8456,N_8301,N_8207);
or U8457 (N_8457,N_8276,N_8288);
and U8458 (N_8458,N_8238,N_8305);
nor U8459 (N_8459,N_8212,N_8263);
nor U8460 (N_8460,N_8375,N_8208);
nand U8461 (N_8461,N_8328,N_8211);
or U8462 (N_8462,N_8377,N_8260);
nand U8463 (N_8463,N_8214,N_8231);
and U8464 (N_8464,N_8280,N_8264);
and U8465 (N_8465,N_8236,N_8282);
and U8466 (N_8466,N_8205,N_8374);
or U8467 (N_8467,N_8335,N_8351);
nand U8468 (N_8468,N_8262,N_8285);
and U8469 (N_8469,N_8243,N_8334);
nand U8470 (N_8470,N_8296,N_8395);
nor U8471 (N_8471,N_8365,N_8234);
and U8472 (N_8472,N_8314,N_8261);
and U8473 (N_8473,N_8321,N_8382);
nor U8474 (N_8474,N_8203,N_8271);
and U8475 (N_8475,N_8339,N_8302);
nor U8476 (N_8476,N_8391,N_8325);
or U8477 (N_8477,N_8327,N_8379);
nand U8478 (N_8478,N_8293,N_8248);
nand U8479 (N_8479,N_8252,N_8291);
and U8480 (N_8480,N_8380,N_8218);
or U8481 (N_8481,N_8390,N_8299);
nand U8482 (N_8482,N_8310,N_8266);
and U8483 (N_8483,N_8370,N_8206);
xor U8484 (N_8484,N_8259,N_8253);
nor U8485 (N_8485,N_8284,N_8367);
and U8486 (N_8486,N_8209,N_8239);
xor U8487 (N_8487,N_8358,N_8225);
nor U8488 (N_8488,N_8224,N_8270);
nand U8489 (N_8489,N_8277,N_8343);
or U8490 (N_8490,N_8398,N_8347);
nand U8491 (N_8491,N_8281,N_8361);
or U8492 (N_8492,N_8287,N_8267);
xnor U8493 (N_8493,N_8378,N_8399);
nor U8494 (N_8494,N_8274,N_8319);
nand U8495 (N_8495,N_8340,N_8326);
nor U8496 (N_8496,N_8265,N_8210);
nor U8497 (N_8497,N_8246,N_8241);
or U8498 (N_8498,N_8316,N_8219);
nor U8499 (N_8499,N_8221,N_8223);
nand U8500 (N_8500,N_8316,N_8214);
or U8501 (N_8501,N_8200,N_8316);
nand U8502 (N_8502,N_8350,N_8293);
nor U8503 (N_8503,N_8257,N_8306);
and U8504 (N_8504,N_8347,N_8306);
or U8505 (N_8505,N_8385,N_8360);
or U8506 (N_8506,N_8298,N_8238);
and U8507 (N_8507,N_8393,N_8320);
nor U8508 (N_8508,N_8235,N_8344);
or U8509 (N_8509,N_8321,N_8376);
nor U8510 (N_8510,N_8273,N_8362);
nand U8511 (N_8511,N_8352,N_8276);
nand U8512 (N_8512,N_8210,N_8357);
and U8513 (N_8513,N_8356,N_8348);
nand U8514 (N_8514,N_8214,N_8237);
or U8515 (N_8515,N_8222,N_8287);
nor U8516 (N_8516,N_8232,N_8295);
nor U8517 (N_8517,N_8334,N_8375);
nand U8518 (N_8518,N_8209,N_8313);
and U8519 (N_8519,N_8344,N_8260);
or U8520 (N_8520,N_8307,N_8230);
and U8521 (N_8521,N_8289,N_8307);
nor U8522 (N_8522,N_8364,N_8212);
nand U8523 (N_8523,N_8217,N_8343);
nor U8524 (N_8524,N_8236,N_8230);
or U8525 (N_8525,N_8360,N_8377);
nor U8526 (N_8526,N_8282,N_8380);
or U8527 (N_8527,N_8396,N_8219);
nand U8528 (N_8528,N_8251,N_8329);
or U8529 (N_8529,N_8230,N_8219);
or U8530 (N_8530,N_8271,N_8387);
or U8531 (N_8531,N_8370,N_8331);
or U8532 (N_8532,N_8338,N_8236);
and U8533 (N_8533,N_8228,N_8323);
nor U8534 (N_8534,N_8362,N_8238);
nor U8535 (N_8535,N_8218,N_8263);
or U8536 (N_8536,N_8211,N_8395);
and U8537 (N_8537,N_8232,N_8284);
xor U8538 (N_8538,N_8278,N_8236);
and U8539 (N_8539,N_8273,N_8246);
nor U8540 (N_8540,N_8333,N_8369);
or U8541 (N_8541,N_8211,N_8225);
nand U8542 (N_8542,N_8284,N_8394);
nand U8543 (N_8543,N_8248,N_8259);
and U8544 (N_8544,N_8311,N_8336);
and U8545 (N_8545,N_8359,N_8200);
nand U8546 (N_8546,N_8246,N_8276);
and U8547 (N_8547,N_8270,N_8216);
or U8548 (N_8548,N_8392,N_8340);
or U8549 (N_8549,N_8226,N_8316);
nand U8550 (N_8550,N_8203,N_8353);
xor U8551 (N_8551,N_8362,N_8298);
nand U8552 (N_8552,N_8322,N_8393);
nand U8553 (N_8553,N_8211,N_8209);
nand U8554 (N_8554,N_8360,N_8388);
and U8555 (N_8555,N_8203,N_8390);
xor U8556 (N_8556,N_8262,N_8261);
nor U8557 (N_8557,N_8290,N_8277);
or U8558 (N_8558,N_8370,N_8219);
nand U8559 (N_8559,N_8368,N_8359);
xor U8560 (N_8560,N_8398,N_8300);
nand U8561 (N_8561,N_8247,N_8357);
xnor U8562 (N_8562,N_8399,N_8287);
and U8563 (N_8563,N_8225,N_8210);
and U8564 (N_8564,N_8256,N_8212);
or U8565 (N_8565,N_8240,N_8378);
and U8566 (N_8566,N_8291,N_8344);
and U8567 (N_8567,N_8240,N_8205);
nand U8568 (N_8568,N_8224,N_8317);
nand U8569 (N_8569,N_8371,N_8320);
or U8570 (N_8570,N_8344,N_8247);
or U8571 (N_8571,N_8234,N_8228);
nand U8572 (N_8572,N_8358,N_8327);
or U8573 (N_8573,N_8358,N_8329);
nor U8574 (N_8574,N_8298,N_8210);
and U8575 (N_8575,N_8240,N_8269);
nand U8576 (N_8576,N_8262,N_8267);
nand U8577 (N_8577,N_8387,N_8312);
and U8578 (N_8578,N_8326,N_8204);
and U8579 (N_8579,N_8244,N_8358);
nor U8580 (N_8580,N_8345,N_8290);
nand U8581 (N_8581,N_8201,N_8306);
nor U8582 (N_8582,N_8371,N_8291);
nor U8583 (N_8583,N_8385,N_8398);
nor U8584 (N_8584,N_8236,N_8284);
and U8585 (N_8585,N_8220,N_8276);
nand U8586 (N_8586,N_8272,N_8252);
or U8587 (N_8587,N_8336,N_8348);
or U8588 (N_8588,N_8330,N_8215);
and U8589 (N_8589,N_8276,N_8205);
nand U8590 (N_8590,N_8250,N_8343);
or U8591 (N_8591,N_8394,N_8395);
or U8592 (N_8592,N_8355,N_8286);
or U8593 (N_8593,N_8396,N_8226);
or U8594 (N_8594,N_8280,N_8314);
nand U8595 (N_8595,N_8248,N_8364);
nor U8596 (N_8596,N_8286,N_8320);
nor U8597 (N_8597,N_8384,N_8257);
and U8598 (N_8598,N_8250,N_8223);
or U8599 (N_8599,N_8391,N_8326);
or U8600 (N_8600,N_8586,N_8525);
nand U8601 (N_8601,N_8470,N_8543);
and U8602 (N_8602,N_8505,N_8423);
nand U8603 (N_8603,N_8424,N_8479);
nor U8604 (N_8604,N_8517,N_8437);
nand U8605 (N_8605,N_8575,N_8560);
nand U8606 (N_8606,N_8414,N_8589);
and U8607 (N_8607,N_8579,N_8478);
nor U8608 (N_8608,N_8494,N_8527);
and U8609 (N_8609,N_8540,N_8475);
or U8610 (N_8610,N_8521,N_8483);
nand U8611 (N_8611,N_8438,N_8440);
and U8612 (N_8612,N_8410,N_8569);
or U8613 (N_8613,N_8404,N_8509);
nand U8614 (N_8614,N_8556,N_8547);
or U8615 (N_8615,N_8412,N_8550);
and U8616 (N_8616,N_8476,N_8489);
and U8617 (N_8617,N_8598,N_8416);
nand U8618 (N_8618,N_8402,N_8587);
nand U8619 (N_8619,N_8452,N_8533);
and U8620 (N_8620,N_8458,N_8559);
and U8621 (N_8621,N_8595,N_8447);
or U8622 (N_8622,N_8488,N_8544);
nor U8623 (N_8623,N_8568,N_8405);
nor U8624 (N_8624,N_8585,N_8596);
and U8625 (N_8625,N_8464,N_8492);
and U8626 (N_8626,N_8431,N_8487);
or U8627 (N_8627,N_8512,N_8480);
nand U8628 (N_8628,N_8418,N_8549);
and U8629 (N_8629,N_8583,N_8571);
nand U8630 (N_8630,N_8481,N_8493);
nand U8631 (N_8631,N_8453,N_8457);
nand U8632 (N_8632,N_8584,N_8409);
nand U8633 (N_8633,N_8562,N_8523);
nor U8634 (N_8634,N_8461,N_8474);
nand U8635 (N_8635,N_8529,N_8422);
or U8636 (N_8636,N_8554,N_8473);
or U8637 (N_8637,N_8514,N_8430);
xor U8638 (N_8638,N_8506,N_8576);
or U8639 (N_8639,N_8518,N_8445);
or U8640 (N_8640,N_8566,N_8501);
nand U8641 (N_8641,N_8408,N_8495);
and U8642 (N_8642,N_8468,N_8439);
or U8643 (N_8643,N_8426,N_8420);
or U8644 (N_8644,N_8580,N_8551);
xor U8645 (N_8645,N_8526,N_8558);
xnor U8646 (N_8646,N_8538,N_8471);
nand U8647 (N_8647,N_8490,N_8515);
nand U8648 (N_8648,N_8441,N_8411);
or U8649 (N_8649,N_8401,N_8565);
or U8650 (N_8650,N_8511,N_8407);
nand U8651 (N_8651,N_8413,N_8536);
and U8652 (N_8652,N_8545,N_8444);
or U8653 (N_8653,N_8541,N_8588);
nor U8654 (N_8654,N_8593,N_8599);
or U8655 (N_8655,N_8557,N_8455);
or U8656 (N_8656,N_8561,N_8510);
or U8657 (N_8657,N_8532,N_8477);
nor U8658 (N_8658,N_8564,N_8432);
nor U8659 (N_8659,N_8429,N_8574);
and U8660 (N_8660,N_8552,N_8442);
nand U8661 (N_8661,N_8528,N_8482);
or U8662 (N_8662,N_8421,N_8415);
nor U8663 (N_8663,N_8594,N_8451);
nand U8664 (N_8664,N_8573,N_8400);
nor U8665 (N_8665,N_8572,N_8433);
and U8666 (N_8666,N_8472,N_8484);
and U8667 (N_8667,N_8443,N_8449);
nand U8668 (N_8668,N_8539,N_8555);
nor U8669 (N_8669,N_8570,N_8592);
or U8670 (N_8670,N_8534,N_8485);
and U8671 (N_8671,N_8446,N_8581);
xor U8672 (N_8672,N_8436,N_8582);
nor U8673 (N_8673,N_8537,N_8425);
or U8674 (N_8674,N_8535,N_8530);
nand U8675 (N_8675,N_8524,N_8591);
nand U8676 (N_8676,N_8520,N_8434);
and U8677 (N_8677,N_8597,N_8454);
nor U8678 (N_8678,N_8507,N_8553);
and U8679 (N_8679,N_8516,N_8450);
nand U8680 (N_8680,N_8519,N_8502);
nand U8681 (N_8681,N_8546,N_8513);
nor U8682 (N_8682,N_8428,N_8460);
nand U8683 (N_8683,N_8435,N_8497);
nand U8684 (N_8684,N_8448,N_8531);
nand U8685 (N_8685,N_8522,N_8496);
or U8686 (N_8686,N_8504,N_8463);
nor U8687 (N_8687,N_8427,N_8491);
or U8688 (N_8688,N_8469,N_8578);
nor U8689 (N_8689,N_8508,N_8486);
and U8690 (N_8690,N_8590,N_8466);
nor U8691 (N_8691,N_8499,N_8419);
or U8692 (N_8692,N_8403,N_8577);
and U8693 (N_8693,N_8467,N_8406);
nand U8694 (N_8694,N_8548,N_8456);
nand U8695 (N_8695,N_8542,N_8498);
or U8696 (N_8696,N_8417,N_8500);
and U8697 (N_8697,N_8459,N_8462);
nand U8698 (N_8698,N_8503,N_8563);
nand U8699 (N_8699,N_8465,N_8567);
and U8700 (N_8700,N_8577,N_8432);
or U8701 (N_8701,N_8426,N_8467);
or U8702 (N_8702,N_8567,N_8539);
or U8703 (N_8703,N_8532,N_8451);
xor U8704 (N_8704,N_8476,N_8529);
nor U8705 (N_8705,N_8533,N_8471);
and U8706 (N_8706,N_8452,N_8499);
and U8707 (N_8707,N_8404,N_8551);
or U8708 (N_8708,N_8456,N_8593);
or U8709 (N_8709,N_8571,N_8556);
nand U8710 (N_8710,N_8419,N_8403);
nor U8711 (N_8711,N_8549,N_8552);
or U8712 (N_8712,N_8448,N_8586);
nor U8713 (N_8713,N_8554,N_8556);
nand U8714 (N_8714,N_8403,N_8413);
nand U8715 (N_8715,N_8489,N_8538);
and U8716 (N_8716,N_8418,N_8559);
nor U8717 (N_8717,N_8527,N_8531);
nor U8718 (N_8718,N_8488,N_8444);
nor U8719 (N_8719,N_8530,N_8448);
nand U8720 (N_8720,N_8477,N_8439);
xor U8721 (N_8721,N_8494,N_8451);
and U8722 (N_8722,N_8524,N_8585);
and U8723 (N_8723,N_8534,N_8480);
and U8724 (N_8724,N_8514,N_8435);
nor U8725 (N_8725,N_8468,N_8444);
and U8726 (N_8726,N_8551,N_8503);
and U8727 (N_8727,N_8501,N_8449);
and U8728 (N_8728,N_8565,N_8440);
or U8729 (N_8729,N_8572,N_8594);
nor U8730 (N_8730,N_8483,N_8466);
or U8731 (N_8731,N_8443,N_8433);
nor U8732 (N_8732,N_8500,N_8563);
or U8733 (N_8733,N_8541,N_8515);
nand U8734 (N_8734,N_8486,N_8481);
nor U8735 (N_8735,N_8544,N_8553);
nand U8736 (N_8736,N_8558,N_8580);
or U8737 (N_8737,N_8588,N_8595);
nand U8738 (N_8738,N_8432,N_8463);
nand U8739 (N_8739,N_8440,N_8434);
or U8740 (N_8740,N_8506,N_8551);
nand U8741 (N_8741,N_8462,N_8421);
or U8742 (N_8742,N_8522,N_8576);
nand U8743 (N_8743,N_8519,N_8516);
or U8744 (N_8744,N_8400,N_8442);
and U8745 (N_8745,N_8517,N_8416);
nand U8746 (N_8746,N_8435,N_8500);
and U8747 (N_8747,N_8522,N_8554);
and U8748 (N_8748,N_8591,N_8497);
or U8749 (N_8749,N_8435,N_8553);
or U8750 (N_8750,N_8555,N_8501);
nand U8751 (N_8751,N_8439,N_8533);
xnor U8752 (N_8752,N_8422,N_8457);
nand U8753 (N_8753,N_8464,N_8531);
nand U8754 (N_8754,N_8404,N_8463);
and U8755 (N_8755,N_8562,N_8498);
nor U8756 (N_8756,N_8461,N_8432);
and U8757 (N_8757,N_8517,N_8490);
or U8758 (N_8758,N_8572,N_8573);
and U8759 (N_8759,N_8486,N_8504);
nor U8760 (N_8760,N_8456,N_8452);
nand U8761 (N_8761,N_8527,N_8499);
nor U8762 (N_8762,N_8579,N_8524);
and U8763 (N_8763,N_8578,N_8492);
and U8764 (N_8764,N_8444,N_8435);
nand U8765 (N_8765,N_8507,N_8577);
and U8766 (N_8766,N_8459,N_8476);
and U8767 (N_8767,N_8534,N_8532);
nor U8768 (N_8768,N_8561,N_8463);
nand U8769 (N_8769,N_8572,N_8535);
nor U8770 (N_8770,N_8404,N_8593);
nor U8771 (N_8771,N_8461,N_8492);
and U8772 (N_8772,N_8432,N_8411);
nand U8773 (N_8773,N_8493,N_8413);
nand U8774 (N_8774,N_8591,N_8578);
nor U8775 (N_8775,N_8438,N_8596);
or U8776 (N_8776,N_8568,N_8502);
and U8777 (N_8777,N_8405,N_8534);
nand U8778 (N_8778,N_8532,N_8493);
nand U8779 (N_8779,N_8486,N_8505);
nand U8780 (N_8780,N_8527,N_8472);
xor U8781 (N_8781,N_8506,N_8468);
nor U8782 (N_8782,N_8487,N_8555);
or U8783 (N_8783,N_8544,N_8499);
nor U8784 (N_8784,N_8457,N_8569);
nand U8785 (N_8785,N_8458,N_8413);
nor U8786 (N_8786,N_8482,N_8418);
and U8787 (N_8787,N_8576,N_8466);
nand U8788 (N_8788,N_8401,N_8487);
nand U8789 (N_8789,N_8427,N_8504);
nand U8790 (N_8790,N_8514,N_8581);
nor U8791 (N_8791,N_8487,N_8413);
and U8792 (N_8792,N_8410,N_8451);
nor U8793 (N_8793,N_8406,N_8435);
and U8794 (N_8794,N_8469,N_8497);
or U8795 (N_8795,N_8562,N_8437);
and U8796 (N_8796,N_8458,N_8499);
nor U8797 (N_8797,N_8434,N_8466);
and U8798 (N_8798,N_8445,N_8550);
and U8799 (N_8799,N_8469,N_8595);
nor U8800 (N_8800,N_8634,N_8748);
nand U8801 (N_8801,N_8743,N_8789);
nand U8802 (N_8802,N_8730,N_8760);
and U8803 (N_8803,N_8784,N_8605);
and U8804 (N_8804,N_8712,N_8621);
or U8805 (N_8805,N_8665,N_8600);
nor U8806 (N_8806,N_8669,N_8762);
or U8807 (N_8807,N_8617,N_8709);
and U8808 (N_8808,N_8662,N_8609);
and U8809 (N_8809,N_8719,N_8783);
nand U8810 (N_8810,N_8693,N_8771);
and U8811 (N_8811,N_8773,N_8657);
and U8812 (N_8812,N_8759,N_8641);
nand U8813 (N_8813,N_8765,N_8677);
nand U8814 (N_8814,N_8660,N_8684);
nor U8815 (N_8815,N_8650,N_8718);
nand U8816 (N_8816,N_8742,N_8739);
nor U8817 (N_8817,N_8612,N_8769);
nor U8818 (N_8818,N_8674,N_8735);
or U8819 (N_8819,N_8701,N_8686);
nand U8820 (N_8820,N_8694,N_8608);
xor U8821 (N_8821,N_8663,N_8607);
and U8822 (N_8822,N_8781,N_8724);
nand U8823 (N_8823,N_8623,N_8797);
or U8824 (N_8824,N_8697,N_8722);
nand U8825 (N_8825,N_8798,N_8792);
or U8826 (N_8826,N_8643,N_8714);
nand U8827 (N_8827,N_8729,N_8611);
and U8828 (N_8828,N_8782,N_8764);
or U8829 (N_8829,N_8645,N_8790);
xnor U8830 (N_8830,N_8635,N_8767);
nor U8831 (N_8831,N_8637,N_8658);
or U8832 (N_8832,N_8620,N_8689);
and U8833 (N_8833,N_8728,N_8750);
nand U8834 (N_8834,N_8647,N_8794);
nand U8835 (N_8835,N_8667,N_8648);
and U8836 (N_8836,N_8733,N_8675);
nand U8837 (N_8837,N_8616,N_8690);
and U8838 (N_8838,N_8779,N_8705);
or U8839 (N_8839,N_8630,N_8726);
nand U8840 (N_8840,N_8699,N_8651);
or U8841 (N_8841,N_8707,N_8668);
and U8842 (N_8842,N_8747,N_8664);
nand U8843 (N_8843,N_8796,N_8752);
nor U8844 (N_8844,N_8741,N_8632);
or U8845 (N_8845,N_8628,N_8780);
or U8846 (N_8846,N_8642,N_8755);
nand U8847 (N_8847,N_8622,N_8654);
nor U8848 (N_8848,N_8793,N_8703);
nand U8849 (N_8849,N_8644,N_8682);
or U8850 (N_8850,N_8702,N_8633);
nor U8851 (N_8851,N_8776,N_8695);
nor U8852 (N_8852,N_8672,N_8656);
or U8853 (N_8853,N_8614,N_8679);
nand U8854 (N_8854,N_8688,N_8626);
nand U8855 (N_8855,N_8671,N_8683);
nand U8856 (N_8856,N_8795,N_8710);
nand U8857 (N_8857,N_8661,N_8754);
or U8858 (N_8858,N_8676,N_8603);
and U8859 (N_8859,N_8638,N_8766);
nor U8860 (N_8860,N_8775,N_8770);
nor U8861 (N_8861,N_8720,N_8731);
and U8862 (N_8862,N_8787,N_8680);
nand U8863 (N_8863,N_8757,N_8799);
and U8864 (N_8864,N_8732,N_8649);
nand U8865 (N_8865,N_8691,N_8704);
or U8866 (N_8866,N_8716,N_8753);
and U8867 (N_8867,N_8713,N_8761);
or U8868 (N_8868,N_8768,N_8717);
and U8869 (N_8869,N_8746,N_8610);
nand U8870 (N_8870,N_8708,N_8618);
or U8871 (N_8871,N_8786,N_8778);
or U8872 (N_8872,N_8652,N_8624);
nor U8873 (N_8873,N_8791,N_8625);
nand U8874 (N_8874,N_8777,N_8758);
nor U8875 (N_8875,N_8745,N_8631);
nor U8876 (N_8876,N_8615,N_8736);
and U8877 (N_8877,N_8627,N_8737);
nor U8878 (N_8878,N_8772,N_8606);
nand U8879 (N_8879,N_8740,N_8687);
nand U8880 (N_8880,N_8619,N_8655);
or U8881 (N_8881,N_8763,N_8629);
and U8882 (N_8882,N_8749,N_8738);
nor U8883 (N_8883,N_8721,N_8604);
nand U8884 (N_8884,N_8715,N_8696);
xnor U8885 (N_8885,N_8636,N_8774);
or U8886 (N_8886,N_8639,N_8678);
and U8887 (N_8887,N_8727,N_8734);
nand U8888 (N_8888,N_8613,N_8756);
nand U8889 (N_8889,N_8700,N_8751);
nand U8890 (N_8890,N_8681,N_8744);
nor U8891 (N_8891,N_8698,N_8601);
nor U8892 (N_8892,N_8706,N_8725);
or U8893 (N_8893,N_8723,N_8711);
nor U8894 (N_8894,N_8692,N_8640);
nor U8895 (N_8895,N_8646,N_8653);
and U8896 (N_8896,N_8685,N_8666);
nand U8897 (N_8897,N_8602,N_8670);
and U8898 (N_8898,N_8659,N_8785);
or U8899 (N_8899,N_8788,N_8673);
nand U8900 (N_8900,N_8750,N_8770);
or U8901 (N_8901,N_8651,N_8628);
nand U8902 (N_8902,N_8679,N_8702);
nor U8903 (N_8903,N_8692,N_8719);
xor U8904 (N_8904,N_8661,N_8693);
and U8905 (N_8905,N_8660,N_8696);
nand U8906 (N_8906,N_8767,N_8671);
nor U8907 (N_8907,N_8618,N_8608);
nor U8908 (N_8908,N_8652,N_8665);
and U8909 (N_8909,N_8603,N_8722);
or U8910 (N_8910,N_8638,N_8640);
nand U8911 (N_8911,N_8762,N_8623);
and U8912 (N_8912,N_8765,N_8647);
and U8913 (N_8913,N_8771,N_8618);
or U8914 (N_8914,N_8633,N_8621);
nand U8915 (N_8915,N_8734,N_8780);
nand U8916 (N_8916,N_8762,N_8797);
and U8917 (N_8917,N_8617,N_8731);
and U8918 (N_8918,N_8697,N_8681);
nor U8919 (N_8919,N_8671,N_8649);
and U8920 (N_8920,N_8649,N_8610);
or U8921 (N_8921,N_8662,N_8675);
and U8922 (N_8922,N_8619,N_8797);
or U8923 (N_8923,N_8646,N_8654);
and U8924 (N_8924,N_8625,N_8672);
or U8925 (N_8925,N_8781,N_8643);
xor U8926 (N_8926,N_8778,N_8616);
nand U8927 (N_8927,N_8717,N_8661);
nand U8928 (N_8928,N_8766,N_8705);
or U8929 (N_8929,N_8626,N_8616);
and U8930 (N_8930,N_8724,N_8798);
xor U8931 (N_8931,N_8675,N_8695);
xnor U8932 (N_8932,N_8606,N_8615);
nand U8933 (N_8933,N_8666,N_8602);
xor U8934 (N_8934,N_8616,N_8714);
or U8935 (N_8935,N_8619,N_8613);
or U8936 (N_8936,N_8608,N_8692);
or U8937 (N_8937,N_8654,N_8603);
and U8938 (N_8938,N_8793,N_8754);
nand U8939 (N_8939,N_8739,N_8644);
or U8940 (N_8940,N_8677,N_8646);
and U8941 (N_8941,N_8618,N_8655);
and U8942 (N_8942,N_8603,N_8613);
nor U8943 (N_8943,N_8600,N_8669);
nor U8944 (N_8944,N_8767,N_8778);
xor U8945 (N_8945,N_8775,N_8638);
nand U8946 (N_8946,N_8612,N_8773);
and U8947 (N_8947,N_8665,N_8661);
nor U8948 (N_8948,N_8733,N_8604);
nand U8949 (N_8949,N_8700,N_8625);
nand U8950 (N_8950,N_8648,N_8615);
nand U8951 (N_8951,N_8735,N_8686);
and U8952 (N_8952,N_8702,N_8650);
nor U8953 (N_8953,N_8780,N_8637);
and U8954 (N_8954,N_8605,N_8783);
nand U8955 (N_8955,N_8652,N_8613);
and U8956 (N_8956,N_8738,N_8711);
nor U8957 (N_8957,N_8602,N_8635);
nand U8958 (N_8958,N_8719,N_8634);
nor U8959 (N_8959,N_8638,N_8610);
nor U8960 (N_8960,N_8766,N_8667);
or U8961 (N_8961,N_8641,N_8711);
nor U8962 (N_8962,N_8701,N_8795);
nand U8963 (N_8963,N_8686,N_8661);
nor U8964 (N_8964,N_8609,N_8713);
nand U8965 (N_8965,N_8735,N_8719);
nand U8966 (N_8966,N_8683,N_8625);
and U8967 (N_8967,N_8704,N_8717);
or U8968 (N_8968,N_8687,N_8615);
and U8969 (N_8969,N_8638,N_8765);
and U8970 (N_8970,N_8708,N_8684);
and U8971 (N_8971,N_8744,N_8687);
nor U8972 (N_8972,N_8666,N_8726);
or U8973 (N_8973,N_8786,N_8775);
or U8974 (N_8974,N_8762,N_8682);
and U8975 (N_8975,N_8679,N_8692);
and U8976 (N_8976,N_8679,N_8775);
nor U8977 (N_8977,N_8624,N_8732);
nor U8978 (N_8978,N_8668,N_8611);
nand U8979 (N_8979,N_8663,N_8678);
nand U8980 (N_8980,N_8659,N_8776);
and U8981 (N_8981,N_8683,N_8629);
or U8982 (N_8982,N_8688,N_8722);
nor U8983 (N_8983,N_8746,N_8772);
nor U8984 (N_8984,N_8750,N_8659);
nor U8985 (N_8985,N_8744,N_8768);
nand U8986 (N_8986,N_8782,N_8724);
and U8987 (N_8987,N_8771,N_8765);
nand U8988 (N_8988,N_8631,N_8721);
or U8989 (N_8989,N_8632,N_8749);
and U8990 (N_8990,N_8756,N_8627);
and U8991 (N_8991,N_8697,N_8688);
or U8992 (N_8992,N_8720,N_8706);
or U8993 (N_8993,N_8762,N_8730);
nand U8994 (N_8994,N_8675,N_8777);
or U8995 (N_8995,N_8791,N_8647);
and U8996 (N_8996,N_8696,N_8786);
and U8997 (N_8997,N_8671,N_8732);
nand U8998 (N_8998,N_8757,N_8614);
nand U8999 (N_8999,N_8697,N_8614);
nand U9000 (N_9000,N_8996,N_8899);
or U9001 (N_9001,N_8998,N_8986);
or U9002 (N_9002,N_8975,N_8909);
nor U9003 (N_9003,N_8843,N_8866);
or U9004 (N_9004,N_8857,N_8826);
or U9005 (N_9005,N_8898,N_8874);
or U9006 (N_9006,N_8905,N_8930);
nand U9007 (N_9007,N_8963,N_8868);
or U9008 (N_9008,N_8987,N_8838);
nor U9009 (N_9009,N_8992,N_8969);
nor U9010 (N_9010,N_8822,N_8994);
or U9011 (N_9011,N_8988,N_8985);
and U9012 (N_9012,N_8890,N_8984);
nand U9013 (N_9013,N_8973,N_8927);
and U9014 (N_9014,N_8958,N_8920);
nand U9015 (N_9015,N_8972,N_8901);
nand U9016 (N_9016,N_8907,N_8924);
or U9017 (N_9017,N_8879,N_8935);
nor U9018 (N_9018,N_8872,N_8944);
and U9019 (N_9019,N_8891,N_8810);
nand U9020 (N_9020,N_8928,N_8808);
nor U9021 (N_9021,N_8837,N_8933);
xor U9022 (N_9022,N_8895,N_8955);
nand U9023 (N_9023,N_8913,N_8981);
nor U9024 (N_9024,N_8851,N_8855);
and U9025 (N_9025,N_8802,N_8881);
or U9026 (N_9026,N_8814,N_8841);
or U9027 (N_9027,N_8856,N_8929);
nor U9028 (N_9028,N_8815,N_8902);
or U9029 (N_9029,N_8825,N_8803);
or U9030 (N_9030,N_8918,N_8806);
nand U9031 (N_9031,N_8862,N_8967);
xnor U9032 (N_9032,N_8961,N_8941);
nor U9033 (N_9033,N_8962,N_8940);
nor U9034 (N_9034,N_8942,N_8840);
nor U9035 (N_9035,N_8807,N_8811);
nand U9036 (N_9036,N_8816,N_8833);
nand U9037 (N_9037,N_8861,N_8812);
nor U9038 (N_9038,N_8974,N_8805);
nor U9039 (N_9039,N_8916,N_8859);
nand U9040 (N_9040,N_8893,N_8846);
xor U9041 (N_9041,N_8925,N_8950);
nor U9042 (N_9042,N_8850,N_8824);
or U9043 (N_9043,N_8858,N_8990);
or U9044 (N_9044,N_8892,N_8852);
nor U9045 (N_9045,N_8818,N_8813);
nand U9046 (N_9046,N_8835,N_8831);
nor U9047 (N_9047,N_8800,N_8820);
nor U9048 (N_9048,N_8885,N_8966);
nor U9049 (N_9049,N_8897,N_8936);
or U9050 (N_9050,N_8853,N_8964);
nand U9051 (N_9051,N_8884,N_8921);
nand U9052 (N_9052,N_8863,N_8948);
nor U9053 (N_9053,N_8980,N_8888);
or U9054 (N_9054,N_8943,N_8821);
or U9055 (N_9055,N_8977,N_8915);
xor U9056 (N_9056,N_8997,N_8968);
nand U9057 (N_9057,N_8991,N_8875);
and U9058 (N_9058,N_8983,N_8871);
and U9059 (N_9059,N_8959,N_8832);
nor U9060 (N_9060,N_8860,N_8819);
nor U9061 (N_9061,N_8900,N_8839);
nand U9062 (N_9062,N_8886,N_8842);
nand U9063 (N_9063,N_8829,N_8931);
nand U9064 (N_9064,N_8912,N_8823);
or U9065 (N_9065,N_8883,N_8878);
nand U9066 (N_9066,N_8946,N_8903);
nand U9067 (N_9067,N_8865,N_8923);
or U9068 (N_9068,N_8911,N_8982);
or U9069 (N_9069,N_8917,N_8922);
or U9070 (N_9070,N_8970,N_8828);
or U9071 (N_9071,N_8876,N_8834);
and U9072 (N_9072,N_8995,N_8926);
and U9073 (N_9073,N_8845,N_8947);
or U9074 (N_9074,N_8889,N_8873);
and U9075 (N_9075,N_8836,N_8801);
or U9076 (N_9076,N_8952,N_8867);
nor U9077 (N_9077,N_8827,N_8993);
and U9078 (N_9078,N_8880,N_8939);
nand U9079 (N_9079,N_8817,N_8934);
nor U9080 (N_9080,N_8847,N_8887);
or U9081 (N_9081,N_8904,N_8896);
nand U9082 (N_9082,N_8882,N_8957);
nor U9083 (N_9083,N_8877,N_8908);
and U9084 (N_9084,N_8804,N_8844);
or U9085 (N_9085,N_8910,N_8965);
nand U9086 (N_9086,N_8999,N_8809);
and U9087 (N_9087,N_8869,N_8932);
nor U9088 (N_9088,N_8864,N_8906);
or U9089 (N_9089,N_8989,N_8971);
nor U9090 (N_9090,N_8854,N_8945);
and U9091 (N_9091,N_8960,N_8938);
nand U9092 (N_9092,N_8848,N_8978);
and U9093 (N_9093,N_8976,N_8914);
and U9094 (N_9094,N_8949,N_8830);
nor U9095 (N_9095,N_8849,N_8956);
nand U9096 (N_9096,N_8870,N_8937);
nand U9097 (N_9097,N_8894,N_8951);
nand U9098 (N_9098,N_8953,N_8919);
or U9099 (N_9099,N_8954,N_8979);
nand U9100 (N_9100,N_8988,N_8850);
nor U9101 (N_9101,N_8837,N_8976);
or U9102 (N_9102,N_8999,N_8907);
and U9103 (N_9103,N_8813,N_8986);
or U9104 (N_9104,N_8956,N_8868);
or U9105 (N_9105,N_8816,N_8917);
nor U9106 (N_9106,N_8964,N_8978);
nand U9107 (N_9107,N_8968,N_8991);
and U9108 (N_9108,N_8875,N_8810);
or U9109 (N_9109,N_8946,N_8928);
nand U9110 (N_9110,N_8857,N_8979);
nand U9111 (N_9111,N_8885,N_8824);
nand U9112 (N_9112,N_8899,N_8875);
nand U9113 (N_9113,N_8824,N_8804);
nor U9114 (N_9114,N_8898,N_8840);
or U9115 (N_9115,N_8808,N_8872);
nor U9116 (N_9116,N_8887,N_8897);
or U9117 (N_9117,N_8903,N_8835);
nor U9118 (N_9118,N_8831,N_8946);
nand U9119 (N_9119,N_8943,N_8838);
nor U9120 (N_9120,N_8847,N_8849);
nor U9121 (N_9121,N_8832,N_8923);
nand U9122 (N_9122,N_8901,N_8961);
nor U9123 (N_9123,N_8859,N_8917);
nand U9124 (N_9124,N_8999,N_8997);
nand U9125 (N_9125,N_8886,N_8837);
nor U9126 (N_9126,N_8944,N_8819);
and U9127 (N_9127,N_8959,N_8855);
nor U9128 (N_9128,N_8997,N_8961);
or U9129 (N_9129,N_8832,N_8935);
and U9130 (N_9130,N_8880,N_8849);
nor U9131 (N_9131,N_8875,N_8928);
or U9132 (N_9132,N_8941,N_8887);
nand U9133 (N_9133,N_8982,N_8822);
or U9134 (N_9134,N_8848,N_8867);
and U9135 (N_9135,N_8829,N_8932);
nor U9136 (N_9136,N_8838,N_8897);
nor U9137 (N_9137,N_8858,N_8901);
and U9138 (N_9138,N_8913,N_8909);
nor U9139 (N_9139,N_8842,N_8807);
nand U9140 (N_9140,N_8895,N_8966);
nor U9141 (N_9141,N_8989,N_8899);
and U9142 (N_9142,N_8958,N_8882);
and U9143 (N_9143,N_8847,N_8850);
nand U9144 (N_9144,N_8914,N_8944);
and U9145 (N_9145,N_8844,N_8985);
nand U9146 (N_9146,N_8812,N_8848);
or U9147 (N_9147,N_8943,N_8855);
nand U9148 (N_9148,N_8894,N_8950);
nor U9149 (N_9149,N_8838,N_8860);
and U9150 (N_9150,N_8809,N_8920);
and U9151 (N_9151,N_8843,N_8961);
nor U9152 (N_9152,N_8860,N_8841);
and U9153 (N_9153,N_8927,N_8870);
nand U9154 (N_9154,N_8937,N_8854);
nand U9155 (N_9155,N_8883,N_8985);
nand U9156 (N_9156,N_8882,N_8977);
nand U9157 (N_9157,N_8900,N_8926);
or U9158 (N_9158,N_8879,N_8959);
or U9159 (N_9159,N_8959,N_8972);
or U9160 (N_9160,N_8957,N_8992);
and U9161 (N_9161,N_8931,N_8984);
or U9162 (N_9162,N_8901,N_8973);
and U9163 (N_9163,N_8928,N_8800);
and U9164 (N_9164,N_8982,N_8803);
nor U9165 (N_9165,N_8858,N_8873);
nor U9166 (N_9166,N_8957,N_8876);
nand U9167 (N_9167,N_8950,N_8895);
and U9168 (N_9168,N_8848,N_8900);
nor U9169 (N_9169,N_8963,N_8865);
nor U9170 (N_9170,N_8892,N_8912);
nand U9171 (N_9171,N_8897,N_8882);
and U9172 (N_9172,N_8893,N_8815);
nand U9173 (N_9173,N_8853,N_8913);
nor U9174 (N_9174,N_8998,N_8892);
and U9175 (N_9175,N_8828,N_8827);
nor U9176 (N_9176,N_8905,N_8864);
or U9177 (N_9177,N_8852,N_8897);
or U9178 (N_9178,N_8938,N_8827);
nor U9179 (N_9179,N_8933,N_8814);
xor U9180 (N_9180,N_8957,N_8987);
nand U9181 (N_9181,N_8897,N_8927);
nor U9182 (N_9182,N_8844,N_8879);
or U9183 (N_9183,N_8906,N_8811);
nand U9184 (N_9184,N_8971,N_8823);
or U9185 (N_9185,N_8938,N_8887);
nand U9186 (N_9186,N_8854,N_8849);
nor U9187 (N_9187,N_8829,N_8806);
nand U9188 (N_9188,N_8919,N_8874);
nand U9189 (N_9189,N_8999,N_8801);
nor U9190 (N_9190,N_8905,N_8992);
nand U9191 (N_9191,N_8852,N_8876);
and U9192 (N_9192,N_8806,N_8958);
nor U9193 (N_9193,N_8903,N_8924);
and U9194 (N_9194,N_8809,N_8926);
nand U9195 (N_9195,N_8810,N_8813);
and U9196 (N_9196,N_8838,N_8965);
xnor U9197 (N_9197,N_8969,N_8930);
and U9198 (N_9198,N_8966,N_8961);
nor U9199 (N_9199,N_8913,N_8851);
and U9200 (N_9200,N_9074,N_9100);
and U9201 (N_9201,N_9152,N_9159);
nand U9202 (N_9202,N_9103,N_9086);
nand U9203 (N_9203,N_9135,N_9003);
nor U9204 (N_9204,N_9094,N_9043);
nor U9205 (N_9205,N_9045,N_9155);
or U9206 (N_9206,N_9018,N_9198);
and U9207 (N_9207,N_9151,N_9013);
nor U9208 (N_9208,N_9049,N_9024);
nand U9209 (N_9209,N_9064,N_9133);
nor U9210 (N_9210,N_9029,N_9032);
nor U9211 (N_9211,N_9104,N_9089);
nand U9212 (N_9212,N_9191,N_9071);
or U9213 (N_9213,N_9118,N_9114);
nand U9214 (N_9214,N_9039,N_9107);
and U9215 (N_9215,N_9156,N_9096);
or U9216 (N_9216,N_9163,N_9053);
and U9217 (N_9217,N_9007,N_9019);
and U9218 (N_9218,N_9162,N_9161);
nand U9219 (N_9219,N_9176,N_9136);
xnor U9220 (N_9220,N_9088,N_9192);
and U9221 (N_9221,N_9066,N_9012);
nand U9222 (N_9222,N_9016,N_9183);
nor U9223 (N_9223,N_9142,N_9084);
nor U9224 (N_9224,N_9083,N_9079);
nor U9225 (N_9225,N_9120,N_9174);
nor U9226 (N_9226,N_9031,N_9122);
and U9227 (N_9227,N_9164,N_9126);
nor U9228 (N_9228,N_9052,N_9195);
and U9229 (N_9229,N_9048,N_9179);
or U9230 (N_9230,N_9129,N_9143);
nor U9231 (N_9231,N_9069,N_9020);
nand U9232 (N_9232,N_9115,N_9040);
xnor U9233 (N_9233,N_9193,N_9178);
nand U9234 (N_9234,N_9072,N_9025);
and U9235 (N_9235,N_9127,N_9093);
or U9236 (N_9236,N_9005,N_9116);
and U9237 (N_9237,N_9169,N_9060);
nand U9238 (N_9238,N_9121,N_9056);
or U9239 (N_9239,N_9008,N_9081);
nor U9240 (N_9240,N_9033,N_9187);
or U9241 (N_9241,N_9131,N_9036);
nor U9242 (N_9242,N_9124,N_9038);
nor U9243 (N_9243,N_9108,N_9180);
or U9244 (N_9244,N_9112,N_9001);
nand U9245 (N_9245,N_9030,N_9182);
or U9246 (N_9246,N_9184,N_9075);
nand U9247 (N_9247,N_9006,N_9128);
nor U9248 (N_9248,N_9197,N_9110);
nor U9249 (N_9249,N_9123,N_9145);
xnor U9250 (N_9250,N_9189,N_9141);
and U9251 (N_9251,N_9065,N_9028);
or U9252 (N_9252,N_9150,N_9000);
nor U9253 (N_9253,N_9011,N_9058);
nand U9254 (N_9254,N_9188,N_9021);
nor U9255 (N_9255,N_9067,N_9160);
nand U9256 (N_9256,N_9175,N_9090);
or U9257 (N_9257,N_9125,N_9144);
nand U9258 (N_9258,N_9185,N_9010);
nand U9259 (N_9259,N_9098,N_9015);
nor U9260 (N_9260,N_9023,N_9167);
and U9261 (N_9261,N_9130,N_9091);
nand U9262 (N_9262,N_9139,N_9014);
or U9263 (N_9263,N_9035,N_9170);
or U9264 (N_9264,N_9190,N_9099);
nor U9265 (N_9265,N_9051,N_9119);
nand U9266 (N_9266,N_9004,N_9148);
or U9267 (N_9267,N_9105,N_9199);
xor U9268 (N_9268,N_9082,N_9077);
or U9269 (N_9269,N_9153,N_9196);
nand U9270 (N_9270,N_9017,N_9073);
or U9271 (N_9271,N_9109,N_9181);
and U9272 (N_9272,N_9027,N_9194);
and U9273 (N_9273,N_9009,N_9050);
or U9274 (N_9274,N_9158,N_9026);
and U9275 (N_9275,N_9166,N_9106);
nor U9276 (N_9276,N_9146,N_9101);
and U9277 (N_9277,N_9168,N_9171);
nand U9278 (N_9278,N_9111,N_9149);
nand U9279 (N_9279,N_9173,N_9087);
or U9280 (N_9280,N_9022,N_9113);
xor U9281 (N_9281,N_9154,N_9002);
and U9282 (N_9282,N_9092,N_9042);
xor U9283 (N_9283,N_9046,N_9057);
nand U9284 (N_9284,N_9044,N_9117);
and U9285 (N_9285,N_9054,N_9165);
and U9286 (N_9286,N_9037,N_9172);
nand U9287 (N_9287,N_9095,N_9047);
nand U9288 (N_9288,N_9147,N_9132);
and U9289 (N_9289,N_9080,N_9140);
or U9290 (N_9290,N_9070,N_9134);
or U9291 (N_9291,N_9137,N_9034);
nand U9292 (N_9292,N_9102,N_9055);
nor U9293 (N_9293,N_9059,N_9078);
nand U9294 (N_9294,N_9068,N_9186);
or U9295 (N_9295,N_9138,N_9076);
and U9296 (N_9296,N_9097,N_9062);
or U9297 (N_9297,N_9085,N_9063);
and U9298 (N_9298,N_9157,N_9177);
nand U9299 (N_9299,N_9061,N_9041);
and U9300 (N_9300,N_9147,N_9188);
and U9301 (N_9301,N_9131,N_9188);
nor U9302 (N_9302,N_9174,N_9082);
and U9303 (N_9303,N_9083,N_9122);
and U9304 (N_9304,N_9099,N_9140);
and U9305 (N_9305,N_9016,N_9078);
or U9306 (N_9306,N_9112,N_9140);
nand U9307 (N_9307,N_9114,N_9152);
nor U9308 (N_9308,N_9027,N_9158);
nor U9309 (N_9309,N_9174,N_9107);
and U9310 (N_9310,N_9144,N_9191);
nand U9311 (N_9311,N_9172,N_9118);
or U9312 (N_9312,N_9005,N_9155);
xor U9313 (N_9313,N_9028,N_9062);
or U9314 (N_9314,N_9100,N_9015);
and U9315 (N_9315,N_9036,N_9129);
or U9316 (N_9316,N_9112,N_9150);
and U9317 (N_9317,N_9187,N_9054);
or U9318 (N_9318,N_9105,N_9031);
nor U9319 (N_9319,N_9030,N_9035);
or U9320 (N_9320,N_9132,N_9167);
and U9321 (N_9321,N_9148,N_9001);
nand U9322 (N_9322,N_9021,N_9193);
and U9323 (N_9323,N_9012,N_9097);
or U9324 (N_9324,N_9056,N_9064);
nor U9325 (N_9325,N_9059,N_9062);
and U9326 (N_9326,N_9125,N_9029);
or U9327 (N_9327,N_9113,N_9085);
nor U9328 (N_9328,N_9003,N_9124);
and U9329 (N_9329,N_9065,N_9010);
nor U9330 (N_9330,N_9156,N_9154);
or U9331 (N_9331,N_9151,N_9001);
or U9332 (N_9332,N_9137,N_9045);
nor U9333 (N_9333,N_9055,N_9112);
or U9334 (N_9334,N_9027,N_9079);
nor U9335 (N_9335,N_9003,N_9050);
nor U9336 (N_9336,N_9067,N_9078);
and U9337 (N_9337,N_9022,N_9097);
or U9338 (N_9338,N_9014,N_9023);
or U9339 (N_9339,N_9130,N_9098);
and U9340 (N_9340,N_9017,N_9180);
nand U9341 (N_9341,N_9015,N_9140);
and U9342 (N_9342,N_9052,N_9053);
nand U9343 (N_9343,N_9168,N_9082);
or U9344 (N_9344,N_9040,N_9149);
nor U9345 (N_9345,N_9155,N_9103);
and U9346 (N_9346,N_9121,N_9104);
and U9347 (N_9347,N_9026,N_9180);
and U9348 (N_9348,N_9053,N_9108);
nor U9349 (N_9349,N_9019,N_9016);
and U9350 (N_9350,N_9149,N_9075);
or U9351 (N_9351,N_9108,N_9035);
nor U9352 (N_9352,N_9111,N_9046);
nand U9353 (N_9353,N_9087,N_9051);
and U9354 (N_9354,N_9094,N_9033);
nand U9355 (N_9355,N_9027,N_9098);
nand U9356 (N_9356,N_9106,N_9013);
nand U9357 (N_9357,N_9015,N_9139);
nand U9358 (N_9358,N_9014,N_9191);
or U9359 (N_9359,N_9121,N_9015);
and U9360 (N_9360,N_9179,N_9030);
nand U9361 (N_9361,N_9012,N_9071);
nor U9362 (N_9362,N_9182,N_9029);
nor U9363 (N_9363,N_9134,N_9167);
or U9364 (N_9364,N_9163,N_9166);
nor U9365 (N_9365,N_9163,N_9112);
or U9366 (N_9366,N_9133,N_9023);
nand U9367 (N_9367,N_9034,N_9080);
or U9368 (N_9368,N_9121,N_9193);
nor U9369 (N_9369,N_9091,N_9063);
nand U9370 (N_9370,N_9111,N_9021);
nor U9371 (N_9371,N_9068,N_9162);
or U9372 (N_9372,N_9191,N_9108);
nor U9373 (N_9373,N_9059,N_9031);
and U9374 (N_9374,N_9106,N_9017);
nor U9375 (N_9375,N_9014,N_9013);
nor U9376 (N_9376,N_9016,N_9128);
nand U9377 (N_9377,N_9176,N_9132);
nor U9378 (N_9378,N_9078,N_9128);
or U9379 (N_9379,N_9090,N_9177);
nand U9380 (N_9380,N_9163,N_9090);
nor U9381 (N_9381,N_9172,N_9185);
nand U9382 (N_9382,N_9121,N_9069);
and U9383 (N_9383,N_9151,N_9174);
and U9384 (N_9384,N_9161,N_9008);
or U9385 (N_9385,N_9065,N_9057);
nor U9386 (N_9386,N_9120,N_9021);
nor U9387 (N_9387,N_9121,N_9034);
nor U9388 (N_9388,N_9102,N_9133);
or U9389 (N_9389,N_9131,N_9167);
nor U9390 (N_9390,N_9134,N_9180);
nor U9391 (N_9391,N_9000,N_9140);
and U9392 (N_9392,N_9054,N_9112);
or U9393 (N_9393,N_9199,N_9060);
nor U9394 (N_9394,N_9074,N_9174);
nor U9395 (N_9395,N_9164,N_9114);
and U9396 (N_9396,N_9043,N_9068);
nand U9397 (N_9397,N_9054,N_9126);
xnor U9398 (N_9398,N_9058,N_9045);
nor U9399 (N_9399,N_9047,N_9086);
xor U9400 (N_9400,N_9296,N_9307);
or U9401 (N_9401,N_9234,N_9326);
and U9402 (N_9402,N_9383,N_9317);
nor U9403 (N_9403,N_9302,N_9391);
nor U9404 (N_9404,N_9204,N_9252);
nand U9405 (N_9405,N_9247,N_9305);
nand U9406 (N_9406,N_9337,N_9268);
or U9407 (N_9407,N_9264,N_9309);
and U9408 (N_9408,N_9265,N_9368);
or U9409 (N_9409,N_9218,N_9333);
nand U9410 (N_9410,N_9294,N_9257);
and U9411 (N_9411,N_9269,N_9213);
or U9412 (N_9412,N_9358,N_9222);
nor U9413 (N_9413,N_9282,N_9224);
nor U9414 (N_9414,N_9350,N_9361);
nand U9415 (N_9415,N_9339,N_9279);
or U9416 (N_9416,N_9208,N_9322);
or U9417 (N_9417,N_9239,N_9342);
or U9418 (N_9418,N_9331,N_9344);
and U9419 (N_9419,N_9356,N_9386);
or U9420 (N_9420,N_9314,N_9238);
or U9421 (N_9421,N_9291,N_9332);
or U9422 (N_9422,N_9274,N_9263);
and U9423 (N_9423,N_9392,N_9364);
nand U9424 (N_9424,N_9323,N_9233);
nor U9425 (N_9425,N_9200,N_9280);
nor U9426 (N_9426,N_9262,N_9290);
nand U9427 (N_9427,N_9226,N_9243);
nor U9428 (N_9428,N_9343,N_9347);
and U9429 (N_9429,N_9345,N_9286);
nand U9430 (N_9430,N_9237,N_9285);
and U9431 (N_9431,N_9273,N_9380);
and U9432 (N_9432,N_9229,N_9308);
nand U9433 (N_9433,N_9271,N_9298);
and U9434 (N_9434,N_9212,N_9341);
nor U9435 (N_9435,N_9351,N_9381);
or U9436 (N_9436,N_9394,N_9359);
or U9437 (N_9437,N_9232,N_9276);
nor U9438 (N_9438,N_9375,N_9330);
nand U9439 (N_9439,N_9354,N_9256);
or U9440 (N_9440,N_9220,N_9369);
nor U9441 (N_9441,N_9312,N_9399);
or U9442 (N_9442,N_9242,N_9217);
and U9443 (N_9443,N_9227,N_9203);
nand U9444 (N_9444,N_9373,N_9367);
nor U9445 (N_9445,N_9251,N_9393);
nand U9446 (N_9446,N_9315,N_9254);
nor U9447 (N_9447,N_9365,N_9299);
nor U9448 (N_9448,N_9211,N_9201);
or U9449 (N_9449,N_9370,N_9230);
or U9450 (N_9450,N_9357,N_9219);
nand U9451 (N_9451,N_9248,N_9244);
or U9452 (N_9452,N_9202,N_9376);
and U9453 (N_9453,N_9398,N_9348);
and U9454 (N_9454,N_9295,N_9396);
nor U9455 (N_9455,N_9231,N_9382);
and U9456 (N_9456,N_9216,N_9306);
nor U9457 (N_9457,N_9260,N_9318);
or U9458 (N_9458,N_9310,N_9390);
nor U9459 (N_9459,N_9209,N_9275);
and U9460 (N_9460,N_9320,N_9215);
nand U9461 (N_9461,N_9372,N_9246);
nor U9462 (N_9462,N_9374,N_9205);
and U9463 (N_9463,N_9206,N_9258);
nand U9464 (N_9464,N_9272,N_9223);
xor U9465 (N_9465,N_9240,N_9384);
and U9466 (N_9466,N_9266,N_9324);
and U9467 (N_9467,N_9270,N_9336);
and U9468 (N_9468,N_9319,N_9207);
and U9469 (N_9469,N_9388,N_9346);
nor U9470 (N_9470,N_9245,N_9301);
nand U9471 (N_9471,N_9225,N_9387);
and U9472 (N_9472,N_9249,N_9250);
and U9473 (N_9473,N_9221,N_9377);
or U9474 (N_9474,N_9321,N_9327);
and U9475 (N_9475,N_9235,N_9255);
or U9476 (N_9476,N_9395,N_9277);
or U9477 (N_9477,N_9293,N_9304);
and U9478 (N_9478,N_9241,N_9397);
nor U9479 (N_9479,N_9385,N_9389);
xor U9480 (N_9480,N_9328,N_9284);
nand U9481 (N_9481,N_9289,N_9210);
or U9482 (N_9482,N_9236,N_9311);
nor U9483 (N_9483,N_9349,N_9228);
and U9484 (N_9484,N_9300,N_9288);
nand U9485 (N_9485,N_9353,N_9363);
nand U9486 (N_9486,N_9261,N_9303);
and U9487 (N_9487,N_9371,N_9338);
and U9488 (N_9488,N_9313,N_9362);
and U9489 (N_9489,N_9340,N_9335);
or U9490 (N_9490,N_9316,N_9366);
or U9491 (N_9491,N_9283,N_9292);
nor U9492 (N_9492,N_9297,N_9325);
nand U9493 (N_9493,N_9329,N_9253);
or U9494 (N_9494,N_9281,N_9278);
nor U9495 (N_9495,N_9287,N_9378);
or U9496 (N_9496,N_9259,N_9334);
and U9497 (N_9497,N_9355,N_9267);
and U9498 (N_9498,N_9214,N_9379);
nand U9499 (N_9499,N_9360,N_9352);
nor U9500 (N_9500,N_9308,N_9269);
nand U9501 (N_9501,N_9252,N_9289);
nor U9502 (N_9502,N_9302,N_9283);
xor U9503 (N_9503,N_9362,N_9292);
nand U9504 (N_9504,N_9381,N_9252);
nand U9505 (N_9505,N_9239,N_9301);
nand U9506 (N_9506,N_9312,N_9251);
nor U9507 (N_9507,N_9210,N_9344);
or U9508 (N_9508,N_9200,N_9221);
and U9509 (N_9509,N_9353,N_9218);
nand U9510 (N_9510,N_9317,N_9349);
or U9511 (N_9511,N_9278,N_9334);
nand U9512 (N_9512,N_9337,N_9232);
or U9513 (N_9513,N_9255,N_9316);
nand U9514 (N_9514,N_9216,N_9396);
nor U9515 (N_9515,N_9295,N_9366);
nor U9516 (N_9516,N_9217,N_9208);
nand U9517 (N_9517,N_9232,N_9201);
nand U9518 (N_9518,N_9297,N_9295);
nand U9519 (N_9519,N_9225,N_9222);
nand U9520 (N_9520,N_9301,N_9246);
or U9521 (N_9521,N_9365,N_9398);
and U9522 (N_9522,N_9238,N_9362);
and U9523 (N_9523,N_9300,N_9355);
and U9524 (N_9524,N_9314,N_9365);
nand U9525 (N_9525,N_9321,N_9298);
nor U9526 (N_9526,N_9381,N_9379);
nand U9527 (N_9527,N_9291,N_9234);
or U9528 (N_9528,N_9320,N_9235);
or U9529 (N_9529,N_9360,N_9301);
or U9530 (N_9530,N_9331,N_9302);
and U9531 (N_9531,N_9248,N_9263);
or U9532 (N_9532,N_9211,N_9358);
nor U9533 (N_9533,N_9317,N_9257);
nor U9534 (N_9534,N_9376,N_9243);
and U9535 (N_9535,N_9303,N_9316);
nand U9536 (N_9536,N_9202,N_9361);
nor U9537 (N_9537,N_9298,N_9327);
or U9538 (N_9538,N_9270,N_9272);
nor U9539 (N_9539,N_9357,N_9210);
nand U9540 (N_9540,N_9268,N_9376);
or U9541 (N_9541,N_9363,N_9271);
nand U9542 (N_9542,N_9306,N_9260);
nand U9543 (N_9543,N_9375,N_9363);
nand U9544 (N_9544,N_9246,N_9373);
nor U9545 (N_9545,N_9225,N_9243);
and U9546 (N_9546,N_9348,N_9212);
and U9547 (N_9547,N_9389,N_9387);
nand U9548 (N_9548,N_9289,N_9355);
and U9549 (N_9549,N_9358,N_9332);
nand U9550 (N_9550,N_9264,N_9209);
nand U9551 (N_9551,N_9236,N_9279);
nor U9552 (N_9552,N_9300,N_9210);
nand U9553 (N_9553,N_9327,N_9262);
or U9554 (N_9554,N_9398,N_9308);
and U9555 (N_9555,N_9376,N_9306);
nand U9556 (N_9556,N_9231,N_9341);
nor U9557 (N_9557,N_9313,N_9244);
and U9558 (N_9558,N_9317,N_9273);
and U9559 (N_9559,N_9296,N_9214);
nand U9560 (N_9560,N_9297,N_9275);
and U9561 (N_9561,N_9227,N_9252);
or U9562 (N_9562,N_9322,N_9373);
nand U9563 (N_9563,N_9218,N_9358);
nand U9564 (N_9564,N_9331,N_9266);
nand U9565 (N_9565,N_9240,N_9213);
nand U9566 (N_9566,N_9255,N_9378);
nand U9567 (N_9567,N_9227,N_9373);
nor U9568 (N_9568,N_9392,N_9215);
nand U9569 (N_9569,N_9323,N_9282);
nor U9570 (N_9570,N_9279,N_9357);
nor U9571 (N_9571,N_9299,N_9361);
nand U9572 (N_9572,N_9284,N_9373);
and U9573 (N_9573,N_9299,N_9236);
and U9574 (N_9574,N_9396,N_9265);
or U9575 (N_9575,N_9208,N_9201);
nor U9576 (N_9576,N_9233,N_9357);
or U9577 (N_9577,N_9228,N_9306);
and U9578 (N_9578,N_9208,N_9389);
or U9579 (N_9579,N_9253,N_9345);
and U9580 (N_9580,N_9338,N_9398);
nand U9581 (N_9581,N_9218,N_9211);
or U9582 (N_9582,N_9254,N_9276);
nand U9583 (N_9583,N_9318,N_9381);
nand U9584 (N_9584,N_9360,N_9394);
and U9585 (N_9585,N_9258,N_9291);
and U9586 (N_9586,N_9281,N_9265);
or U9587 (N_9587,N_9349,N_9251);
nand U9588 (N_9588,N_9345,N_9353);
nand U9589 (N_9589,N_9381,N_9212);
or U9590 (N_9590,N_9206,N_9275);
and U9591 (N_9591,N_9242,N_9386);
xor U9592 (N_9592,N_9270,N_9333);
nor U9593 (N_9593,N_9255,N_9225);
or U9594 (N_9594,N_9282,N_9366);
or U9595 (N_9595,N_9263,N_9284);
nand U9596 (N_9596,N_9267,N_9290);
and U9597 (N_9597,N_9228,N_9343);
or U9598 (N_9598,N_9241,N_9337);
xor U9599 (N_9599,N_9324,N_9379);
nor U9600 (N_9600,N_9489,N_9560);
or U9601 (N_9601,N_9483,N_9515);
nor U9602 (N_9602,N_9570,N_9541);
nand U9603 (N_9603,N_9456,N_9514);
nor U9604 (N_9604,N_9518,N_9440);
or U9605 (N_9605,N_9459,N_9471);
nand U9606 (N_9606,N_9400,N_9406);
nor U9607 (N_9607,N_9436,N_9485);
nand U9608 (N_9608,N_9506,N_9463);
and U9609 (N_9609,N_9487,N_9563);
and U9610 (N_9610,N_9408,N_9465);
nand U9611 (N_9611,N_9470,N_9493);
nor U9612 (N_9612,N_9451,N_9539);
nor U9613 (N_9613,N_9512,N_9543);
and U9614 (N_9614,N_9454,N_9547);
nand U9615 (N_9615,N_9409,N_9589);
or U9616 (N_9616,N_9519,N_9434);
nand U9617 (N_9617,N_9476,N_9484);
or U9618 (N_9618,N_9528,N_9402);
and U9619 (N_9619,N_9522,N_9486);
nor U9620 (N_9620,N_9510,N_9532);
nand U9621 (N_9621,N_9521,N_9533);
nor U9622 (N_9622,N_9420,N_9540);
nand U9623 (N_9623,N_9555,N_9500);
and U9624 (N_9624,N_9473,N_9588);
and U9625 (N_9625,N_9401,N_9417);
or U9626 (N_9626,N_9529,N_9558);
and U9627 (N_9627,N_9415,N_9536);
and U9628 (N_9628,N_9449,N_9425);
or U9629 (N_9629,N_9446,N_9504);
and U9630 (N_9630,N_9578,N_9579);
nand U9631 (N_9631,N_9403,N_9564);
nor U9632 (N_9632,N_9495,N_9534);
nand U9633 (N_9633,N_9468,N_9491);
or U9634 (N_9634,N_9404,N_9571);
or U9635 (N_9635,N_9542,N_9419);
nor U9636 (N_9636,N_9412,N_9479);
or U9637 (N_9637,N_9581,N_9430);
nor U9638 (N_9638,N_9592,N_9458);
nor U9639 (N_9639,N_9499,N_9494);
or U9640 (N_9640,N_9464,N_9525);
and U9641 (N_9641,N_9410,N_9552);
and U9642 (N_9642,N_9594,N_9573);
nor U9643 (N_9643,N_9439,N_9460);
and U9644 (N_9644,N_9452,N_9414);
xnor U9645 (N_9645,N_9482,N_9432);
nand U9646 (N_9646,N_9531,N_9523);
nand U9647 (N_9647,N_9561,N_9427);
and U9648 (N_9648,N_9527,N_9582);
nand U9649 (N_9649,N_9469,N_9587);
xnor U9650 (N_9650,N_9590,N_9435);
nor U9651 (N_9651,N_9447,N_9569);
nand U9652 (N_9652,N_9442,N_9443);
and U9653 (N_9653,N_9441,N_9405);
and U9654 (N_9654,N_9583,N_9545);
nand U9655 (N_9655,N_9538,N_9492);
nand U9656 (N_9656,N_9593,N_9407);
or U9657 (N_9657,N_9509,N_9575);
and U9658 (N_9658,N_9411,N_9537);
nand U9659 (N_9659,N_9576,N_9511);
nor U9660 (N_9660,N_9461,N_9503);
xor U9661 (N_9661,N_9466,N_9445);
or U9662 (N_9662,N_9429,N_9580);
nor U9663 (N_9663,N_9551,N_9549);
and U9664 (N_9664,N_9413,N_9548);
or U9665 (N_9665,N_9556,N_9572);
and U9666 (N_9666,N_9554,N_9457);
and U9667 (N_9667,N_9544,N_9584);
and U9668 (N_9668,N_9421,N_9565);
nand U9669 (N_9669,N_9497,N_9559);
nand U9670 (N_9670,N_9524,N_9422);
nor U9671 (N_9671,N_9508,N_9505);
or U9672 (N_9672,N_9574,N_9428);
and U9673 (N_9673,N_9513,N_9546);
nor U9674 (N_9674,N_9498,N_9475);
nand U9675 (N_9675,N_9530,N_9598);
and U9676 (N_9676,N_9520,N_9462);
nor U9677 (N_9677,N_9501,N_9535);
nor U9678 (N_9678,N_9431,N_9480);
nor U9679 (N_9679,N_9444,N_9478);
nand U9680 (N_9680,N_9453,N_9577);
or U9681 (N_9681,N_9490,N_9586);
or U9682 (N_9682,N_9416,N_9481);
xnor U9683 (N_9683,N_9448,N_9585);
and U9684 (N_9684,N_9557,N_9566);
nand U9685 (N_9685,N_9567,N_9516);
and U9686 (N_9686,N_9597,N_9418);
nor U9687 (N_9687,N_9450,N_9517);
nor U9688 (N_9688,N_9474,N_9507);
or U9689 (N_9689,N_9595,N_9472);
and U9690 (N_9690,N_9467,N_9568);
nor U9691 (N_9691,N_9502,N_9591);
or U9692 (N_9692,N_9437,N_9550);
xor U9693 (N_9693,N_9562,N_9553);
and U9694 (N_9694,N_9488,N_9455);
nor U9695 (N_9695,N_9496,N_9423);
or U9696 (N_9696,N_9426,N_9526);
nand U9697 (N_9697,N_9424,N_9599);
nor U9698 (N_9698,N_9477,N_9596);
or U9699 (N_9699,N_9433,N_9438);
and U9700 (N_9700,N_9564,N_9433);
or U9701 (N_9701,N_9418,N_9507);
or U9702 (N_9702,N_9493,N_9497);
nand U9703 (N_9703,N_9523,N_9459);
and U9704 (N_9704,N_9460,N_9469);
nor U9705 (N_9705,N_9521,N_9419);
or U9706 (N_9706,N_9408,N_9530);
or U9707 (N_9707,N_9442,N_9571);
xor U9708 (N_9708,N_9436,N_9479);
and U9709 (N_9709,N_9506,N_9404);
xnor U9710 (N_9710,N_9546,N_9598);
or U9711 (N_9711,N_9476,N_9563);
and U9712 (N_9712,N_9427,N_9568);
and U9713 (N_9713,N_9536,N_9413);
nor U9714 (N_9714,N_9473,N_9453);
nand U9715 (N_9715,N_9490,N_9542);
and U9716 (N_9716,N_9428,N_9511);
nand U9717 (N_9717,N_9556,N_9546);
nand U9718 (N_9718,N_9474,N_9553);
or U9719 (N_9719,N_9543,N_9473);
and U9720 (N_9720,N_9578,N_9415);
nor U9721 (N_9721,N_9566,N_9447);
and U9722 (N_9722,N_9545,N_9430);
nor U9723 (N_9723,N_9583,N_9428);
and U9724 (N_9724,N_9521,N_9441);
nor U9725 (N_9725,N_9414,N_9408);
and U9726 (N_9726,N_9430,N_9523);
and U9727 (N_9727,N_9557,N_9435);
nand U9728 (N_9728,N_9408,N_9491);
or U9729 (N_9729,N_9514,N_9401);
and U9730 (N_9730,N_9415,N_9552);
nand U9731 (N_9731,N_9530,N_9424);
and U9732 (N_9732,N_9450,N_9442);
nor U9733 (N_9733,N_9453,N_9428);
or U9734 (N_9734,N_9468,N_9419);
nor U9735 (N_9735,N_9502,N_9535);
nor U9736 (N_9736,N_9572,N_9467);
or U9737 (N_9737,N_9581,N_9516);
and U9738 (N_9738,N_9588,N_9529);
or U9739 (N_9739,N_9576,N_9484);
or U9740 (N_9740,N_9520,N_9566);
nor U9741 (N_9741,N_9481,N_9470);
or U9742 (N_9742,N_9457,N_9468);
nand U9743 (N_9743,N_9461,N_9429);
and U9744 (N_9744,N_9532,N_9587);
or U9745 (N_9745,N_9467,N_9515);
nor U9746 (N_9746,N_9545,N_9480);
nand U9747 (N_9747,N_9586,N_9554);
or U9748 (N_9748,N_9576,N_9400);
xnor U9749 (N_9749,N_9508,N_9439);
xor U9750 (N_9750,N_9584,N_9446);
xnor U9751 (N_9751,N_9471,N_9431);
and U9752 (N_9752,N_9521,N_9512);
and U9753 (N_9753,N_9565,N_9518);
nor U9754 (N_9754,N_9585,N_9502);
nand U9755 (N_9755,N_9524,N_9437);
or U9756 (N_9756,N_9522,N_9504);
nand U9757 (N_9757,N_9517,N_9412);
and U9758 (N_9758,N_9500,N_9459);
and U9759 (N_9759,N_9486,N_9406);
nand U9760 (N_9760,N_9550,N_9505);
nor U9761 (N_9761,N_9587,N_9435);
nand U9762 (N_9762,N_9503,N_9478);
nand U9763 (N_9763,N_9542,N_9497);
nor U9764 (N_9764,N_9462,N_9540);
nand U9765 (N_9765,N_9496,N_9539);
nand U9766 (N_9766,N_9588,N_9430);
xor U9767 (N_9767,N_9510,N_9526);
nand U9768 (N_9768,N_9466,N_9579);
nand U9769 (N_9769,N_9518,N_9597);
nand U9770 (N_9770,N_9440,N_9563);
and U9771 (N_9771,N_9427,N_9599);
or U9772 (N_9772,N_9438,N_9521);
nand U9773 (N_9773,N_9585,N_9512);
nand U9774 (N_9774,N_9496,N_9464);
nor U9775 (N_9775,N_9533,N_9587);
xor U9776 (N_9776,N_9534,N_9423);
nand U9777 (N_9777,N_9484,N_9545);
or U9778 (N_9778,N_9412,N_9502);
or U9779 (N_9779,N_9533,N_9570);
nor U9780 (N_9780,N_9453,N_9402);
or U9781 (N_9781,N_9504,N_9598);
nand U9782 (N_9782,N_9564,N_9519);
and U9783 (N_9783,N_9417,N_9407);
and U9784 (N_9784,N_9483,N_9563);
nand U9785 (N_9785,N_9417,N_9471);
and U9786 (N_9786,N_9552,N_9430);
or U9787 (N_9787,N_9486,N_9541);
nor U9788 (N_9788,N_9537,N_9573);
or U9789 (N_9789,N_9562,N_9580);
nor U9790 (N_9790,N_9554,N_9458);
and U9791 (N_9791,N_9544,N_9583);
nand U9792 (N_9792,N_9423,N_9439);
nand U9793 (N_9793,N_9478,N_9537);
nor U9794 (N_9794,N_9432,N_9474);
and U9795 (N_9795,N_9515,N_9434);
or U9796 (N_9796,N_9507,N_9459);
or U9797 (N_9797,N_9414,N_9529);
nor U9798 (N_9798,N_9419,N_9566);
and U9799 (N_9799,N_9560,N_9533);
nor U9800 (N_9800,N_9700,N_9743);
and U9801 (N_9801,N_9714,N_9744);
or U9802 (N_9802,N_9774,N_9654);
nand U9803 (N_9803,N_9685,N_9646);
nand U9804 (N_9804,N_9745,N_9695);
or U9805 (N_9805,N_9675,N_9606);
nand U9806 (N_9806,N_9756,N_9611);
nand U9807 (N_9807,N_9721,N_9698);
or U9808 (N_9808,N_9639,N_9788);
nand U9809 (N_9809,N_9794,N_9659);
and U9810 (N_9810,N_9795,N_9679);
and U9811 (N_9811,N_9682,N_9770);
nand U9812 (N_9812,N_9637,N_9783);
nand U9813 (N_9813,N_9663,N_9749);
nor U9814 (N_9814,N_9643,N_9723);
and U9815 (N_9815,N_9773,N_9716);
nor U9816 (N_9816,N_9612,N_9674);
and U9817 (N_9817,N_9705,N_9796);
and U9818 (N_9818,N_9656,N_9616);
nor U9819 (N_9819,N_9617,N_9691);
and U9820 (N_9820,N_9760,N_9621);
nor U9821 (N_9821,N_9687,N_9694);
or U9822 (N_9822,N_9733,N_9764);
nor U9823 (N_9823,N_9668,N_9603);
and U9824 (N_9824,N_9799,N_9672);
and U9825 (N_9825,N_9708,N_9759);
nand U9826 (N_9826,N_9734,N_9693);
nor U9827 (N_9827,N_9629,N_9625);
nand U9828 (N_9828,N_9701,N_9747);
nor U9829 (N_9829,N_9791,N_9624);
nand U9830 (N_9830,N_9785,N_9607);
nand U9831 (N_9831,N_9648,N_9667);
nor U9832 (N_9832,N_9697,N_9609);
nand U9833 (N_9833,N_9608,N_9720);
and U9834 (N_9834,N_9618,N_9731);
and U9835 (N_9835,N_9758,N_9664);
or U9836 (N_9836,N_9692,N_9657);
xor U9837 (N_9837,N_9626,N_9666);
or U9838 (N_9838,N_9623,N_9677);
xnor U9839 (N_9839,N_9752,N_9613);
nor U9840 (N_9840,N_9702,N_9600);
and U9841 (N_9841,N_9673,N_9620);
nand U9842 (N_9842,N_9653,N_9633);
and U9843 (N_9843,N_9670,N_9767);
nor U9844 (N_9844,N_9719,N_9661);
and U9845 (N_9845,N_9640,N_9790);
nor U9846 (N_9846,N_9736,N_9737);
or U9847 (N_9847,N_9746,N_9751);
and U9848 (N_9848,N_9699,N_9761);
xnor U9849 (N_9849,N_9614,N_9631);
nor U9850 (N_9850,N_9724,N_9615);
nor U9851 (N_9851,N_9688,N_9797);
nor U9852 (N_9852,N_9717,N_9622);
xor U9853 (N_9853,N_9722,N_9728);
and U9854 (N_9854,N_9781,N_9650);
and U9855 (N_9855,N_9610,N_9707);
nand U9856 (N_9856,N_9658,N_9776);
nand U9857 (N_9857,N_9642,N_9780);
nand U9858 (N_9858,N_9636,N_9712);
nand U9859 (N_9859,N_9789,N_9772);
or U9860 (N_9860,N_9740,N_9684);
or U9861 (N_9861,N_9604,N_9715);
and U9862 (N_9862,N_9676,N_9727);
or U9863 (N_9863,N_9696,N_9627);
or U9864 (N_9864,N_9634,N_9768);
nand U9865 (N_9865,N_9605,N_9638);
or U9866 (N_9866,N_9738,N_9711);
nor U9867 (N_9867,N_9678,N_9787);
nor U9868 (N_9868,N_9742,N_9644);
xor U9869 (N_9869,N_9645,N_9690);
nor U9870 (N_9870,N_9635,N_9769);
xnor U9871 (N_9871,N_9703,N_9725);
or U9872 (N_9872,N_9619,N_9706);
nor U9873 (N_9873,N_9748,N_9628);
nand U9874 (N_9874,N_9683,N_9753);
nor U9875 (N_9875,N_9689,N_9686);
nor U9876 (N_9876,N_9671,N_9778);
and U9877 (N_9877,N_9662,N_9632);
nor U9878 (N_9878,N_9730,N_9750);
or U9879 (N_9879,N_9775,N_9786);
nand U9880 (N_9880,N_9630,N_9680);
nor U9881 (N_9881,N_9601,N_9762);
nor U9882 (N_9882,N_9732,N_9718);
or U9883 (N_9883,N_9726,N_9709);
or U9884 (N_9884,N_9704,N_9765);
nor U9885 (N_9885,N_9602,N_9777);
nor U9886 (N_9886,N_9660,N_9655);
nand U9887 (N_9887,N_9729,N_9739);
nor U9888 (N_9888,N_9641,N_9766);
and U9889 (N_9889,N_9681,N_9647);
nand U9890 (N_9890,N_9782,N_9755);
nand U9891 (N_9891,N_9779,N_9757);
nor U9892 (N_9892,N_9784,N_9652);
nand U9893 (N_9893,N_9754,N_9735);
and U9894 (N_9894,N_9798,N_9792);
nor U9895 (N_9895,N_9713,N_9763);
or U9896 (N_9896,N_9651,N_9649);
nor U9897 (N_9897,N_9771,N_9669);
nand U9898 (N_9898,N_9741,N_9793);
or U9899 (N_9899,N_9710,N_9665);
and U9900 (N_9900,N_9648,N_9794);
or U9901 (N_9901,N_9677,N_9722);
nand U9902 (N_9902,N_9602,N_9723);
and U9903 (N_9903,N_9715,N_9702);
and U9904 (N_9904,N_9729,N_9605);
xor U9905 (N_9905,N_9741,N_9739);
nor U9906 (N_9906,N_9791,N_9613);
or U9907 (N_9907,N_9708,N_9624);
nand U9908 (N_9908,N_9602,N_9621);
nand U9909 (N_9909,N_9680,N_9694);
or U9910 (N_9910,N_9746,N_9632);
and U9911 (N_9911,N_9690,N_9671);
nor U9912 (N_9912,N_9683,N_9632);
nor U9913 (N_9913,N_9752,N_9726);
and U9914 (N_9914,N_9771,N_9611);
nor U9915 (N_9915,N_9735,N_9736);
nand U9916 (N_9916,N_9731,N_9659);
and U9917 (N_9917,N_9740,N_9780);
and U9918 (N_9918,N_9614,N_9679);
nand U9919 (N_9919,N_9744,N_9645);
nor U9920 (N_9920,N_9620,N_9751);
nor U9921 (N_9921,N_9768,N_9718);
nand U9922 (N_9922,N_9745,N_9706);
or U9923 (N_9923,N_9725,N_9653);
nor U9924 (N_9924,N_9716,N_9732);
or U9925 (N_9925,N_9786,N_9734);
nand U9926 (N_9926,N_9733,N_9640);
nand U9927 (N_9927,N_9757,N_9629);
xnor U9928 (N_9928,N_9646,N_9670);
nor U9929 (N_9929,N_9679,N_9733);
and U9930 (N_9930,N_9736,N_9664);
and U9931 (N_9931,N_9725,N_9635);
nand U9932 (N_9932,N_9750,N_9679);
nor U9933 (N_9933,N_9727,N_9799);
or U9934 (N_9934,N_9774,N_9735);
nor U9935 (N_9935,N_9705,N_9636);
nand U9936 (N_9936,N_9691,N_9696);
nor U9937 (N_9937,N_9711,N_9685);
nor U9938 (N_9938,N_9763,N_9755);
or U9939 (N_9939,N_9619,N_9646);
and U9940 (N_9940,N_9779,N_9613);
or U9941 (N_9941,N_9721,N_9752);
and U9942 (N_9942,N_9624,N_9785);
or U9943 (N_9943,N_9747,N_9785);
nand U9944 (N_9944,N_9600,N_9712);
or U9945 (N_9945,N_9685,N_9633);
nand U9946 (N_9946,N_9697,N_9796);
nand U9947 (N_9947,N_9652,N_9643);
nand U9948 (N_9948,N_9713,N_9777);
nand U9949 (N_9949,N_9711,N_9612);
and U9950 (N_9950,N_9776,N_9782);
and U9951 (N_9951,N_9754,N_9691);
and U9952 (N_9952,N_9636,N_9710);
xnor U9953 (N_9953,N_9686,N_9745);
or U9954 (N_9954,N_9735,N_9780);
and U9955 (N_9955,N_9706,N_9689);
or U9956 (N_9956,N_9746,N_9613);
nand U9957 (N_9957,N_9763,N_9626);
nand U9958 (N_9958,N_9705,N_9618);
and U9959 (N_9959,N_9723,N_9660);
nor U9960 (N_9960,N_9630,N_9671);
nand U9961 (N_9961,N_9796,N_9706);
or U9962 (N_9962,N_9613,N_9679);
nand U9963 (N_9963,N_9735,N_9728);
nand U9964 (N_9964,N_9716,N_9737);
and U9965 (N_9965,N_9745,N_9631);
and U9966 (N_9966,N_9788,N_9771);
or U9967 (N_9967,N_9637,N_9747);
and U9968 (N_9968,N_9689,N_9777);
or U9969 (N_9969,N_9664,N_9701);
xor U9970 (N_9970,N_9710,N_9644);
nand U9971 (N_9971,N_9751,N_9732);
nand U9972 (N_9972,N_9742,N_9613);
or U9973 (N_9973,N_9743,N_9633);
nor U9974 (N_9974,N_9695,N_9622);
nor U9975 (N_9975,N_9754,N_9685);
or U9976 (N_9976,N_9755,N_9709);
nand U9977 (N_9977,N_9786,N_9727);
and U9978 (N_9978,N_9680,N_9690);
nor U9979 (N_9979,N_9747,N_9765);
and U9980 (N_9980,N_9617,N_9701);
nor U9981 (N_9981,N_9782,N_9780);
or U9982 (N_9982,N_9754,N_9665);
or U9983 (N_9983,N_9631,N_9691);
nor U9984 (N_9984,N_9724,N_9707);
and U9985 (N_9985,N_9772,N_9619);
or U9986 (N_9986,N_9647,N_9687);
nor U9987 (N_9987,N_9700,N_9668);
or U9988 (N_9988,N_9671,N_9769);
and U9989 (N_9989,N_9605,N_9770);
or U9990 (N_9990,N_9760,N_9664);
nand U9991 (N_9991,N_9747,N_9673);
and U9992 (N_9992,N_9631,N_9744);
nand U9993 (N_9993,N_9694,N_9793);
nand U9994 (N_9994,N_9707,N_9681);
and U9995 (N_9995,N_9614,N_9772);
or U9996 (N_9996,N_9706,N_9697);
nand U9997 (N_9997,N_9617,N_9698);
nor U9998 (N_9998,N_9730,N_9721);
nand U9999 (N_9999,N_9664,N_9680);
nand U10000 (N_10000,N_9820,N_9815);
and U10001 (N_10001,N_9851,N_9891);
and U10002 (N_10002,N_9937,N_9987);
and U10003 (N_10003,N_9809,N_9860);
nand U10004 (N_10004,N_9900,N_9874);
nand U10005 (N_10005,N_9973,N_9837);
nand U10006 (N_10006,N_9804,N_9907);
nor U10007 (N_10007,N_9944,N_9818);
nand U10008 (N_10008,N_9908,N_9921);
xnor U10009 (N_10009,N_9914,N_9941);
or U10010 (N_10010,N_9835,N_9802);
nand U10011 (N_10011,N_9992,N_9883);
nor U10012 (N_10012,N_9866,N_9875);
or U10013 (N_10013,N_9884,N_9968);
nand U10014 (N_10014,N_9995,N_9857);
or U10015 (N_10015,N_9840,N_9810);
nor U10016 (N_10016,N_9825,N_9871);
or U10017 (N_10017,N_9890,N_9822);
nand U10018 (N_10018,N_9976,N_9811);
or U10019 (N_10019,N_9889,N_9915);
and U10020 (N_10020,N_9933,N_9988);
nor U10021 (N_10021,N_9909,N_9958);
and U10022 (N_10022,N_9967,N_9943);
nand U10023 (N_10023,N_9924,N_9852);
and U10024 (N_10024,N_9950,N_9865);
and U10025 (N_10025,N_9956,N_9942);
nor U10026 (N_10026,N_9990,N_9927);
nand U10027 (N_10027,N_9827,N_9954);
nor U10028 (N_10028,N_9910,N_9858);
nor U10029 (N_10029,N_9993,N_9952);
nand U10030 (N_10030,N_9962,N_9882);
or U10031 (N_10031,N_9917,N_9959);
or U10032 (N_10032,N_9980,N_9940);
xor U10033 (N_10033,N_9912,N_9977);
nor U10034 (N_10034,N_9894,N_9964);
or U10035 (N_10035,N_9824,N_9853);
nor U10036 (N_10036,N_9916,N_9850);
nor U10037 (N_10037,N_9949,N_9951);
nand U10038 (N_10038,N_9861,N_9862);
and U10039 (N_10039,N_9854,N_9945);
nor U10040 (N_10040,N_9832,N_9869);
xor U10041 (N_10041,N_9846,N_9981);
nand U10042 (N_10042,N_9946,N_9831);
or U10043 (N_10043,N_9934,N_9816);
nor U10044 (N_10044,N_9877,N_9885);
and U10045 (N_10045,N_9834,N_9975);
nand U10046 (N_10046,N_9955,N_9895);
xnor U10047 (N_10047,N_9925,N_9948);
and U10048 (N_10048,N_9872,N_9829);
and U10049 (N_10049,N_9984,N_9893);
nand U10050 (N_10050,N_9863,N_9898);
nor U10051 (N_10051,N_9978,N_9897);
nand U10052 (N_10052,N_9957,N_9803);
nor U10053 (N_10053,N_9807,N_9983);
or U10054 (N_10054,N_9801,N_9808);
and U10055 (N_10055,N_9918,N_9844);
and U10056 (N_10056,N_9888,N_9938);
and U10057 (N_10057,N_9930,N_9859);
or U10058 (N_10058,N_9974,N_9873);
nand U10059 (N_10059,N_9982,N_9848);
nor U10060 (N_10060,N_9991,N_9963);
or U10061 (N_10061,N_9979,N_9970);
nand U10062 (N_10062,N_9881,N_9901);
nand U10063 (N_10063,N_9969,N_9935);
and U10064 (N_10064,N_9986,N_9932);
and U10065 (N_10065,N_9887,N_9999);
nor U10066 (N_10066,N_9939,N_9806);
nor U10067 (N_10067,N_9870,N_9902);
and U10068 (N_10068,N_9886,N_9936);
or U10069 (N_10069,N_9998,N_9830);
nor U10070 (N_10070,N_9905,N_9826);
nor U10071 (N_10071,N_9828,N_9920);
or U10072 (N_10072,N_9855,N_9926);
or U10073 (N_10073,N_9814,N_9922);
nand U10074 (N_10074,N_9972,N_9997);
nand U10075 (N_10075,N_9896,N_9929);
or U10076 (N_10076,N_9817,N_9971);
or U10077 (N_10077,N_9845,N_9903);
nand U10078 (N_10078,N_9965,N_9994);
or U10079 (N_10079,N_9919,N_9812);
nand U10080 (N_10080,N_9843,N_9960);
nand U10081 (N_10081,N_9878,N_9868);
and U10082 (N_10082,N_9841,N_9842);
nand U10083 (N_10083,N_9856,N_9904);
or U10084 (N_10084,N_9800,N_9966);
and U10085 (N_10085,N_9996,N_9892);
or U10086 (N_10086,N_9928,N_9899);
or U10087 (N_10087,N_9985,N_9906);
and U10088 (N_10088,N_9847,N_9879);
nor U10089 (N_10089,N_9876,N_9836);
and U10090 (N_10090,N_9961,N_9989);
nand U10091 (N_10091,N_9805,N_9813);
or U10092 (N_10092,N_9911,N_9823);
and U10093 (N_10093,N_9923,N_9821);
and U10094 (N_10094,N_9913,N_9947);
or U10095 (N_10095,N_9838,N_9953);
or U10096 (N_10096,N_9839,N_9880);
or U10097 (N_10097,N_9864,N_9931);
nand U10098 (N_10098,N_9833,N_9849);
or U10099 (N_10099,N_9819,N_9867);
and U10100 (N_10100,N_9966,N_9995);
nor U10101 (N_10101,N_9902,N_9833);
nor U10102 (N_10102,N_9854,N_9875);
nand U10103 (N_10103,N_9802,N_9827);
nand U10104 (N_10104,N_9869,N_9942);
nand U10105 (N_10105,N_9883,N_9987);
or U10106 (N_10106,N_9916,N_9951);
nand U10107 (N_10107,N_9943,N_9957);
nor U10108 (N_10108,N_9806,N_9863);
nand U10109 (N_10109,N_9874,N_9985);
nor U10110 (N_10110,N_9908,N_9978);
nor U10111 (N_10111,N_9906,N_9907);
and U10112 (N_10112,N_9995,N_9812);
or U10113 (N_10113,N_9940,N_9902);
and U10114 (N_10114,N_9934,N_9946);
or U10115 (N_10115,N_9942,N_9814);
nor U10116 (N_10116,N_9874,N_9867);
nor U10117 (N_10117,N_9880,N_9943);
nor U10118 (N_10118,N_9918,N_9862);
nor U10119 (N_10119,N_9851,N_9823);
or U10120 (N_10120,N_9801,N_9991);
nor U10121 (N_10121,N_9903,N_9997);
and U10122 (N_10122,N_9951,N_9801);
and U10123 (N_10123,N_9821,N_9847);
or U10124 (N_10124,N_9895,N_9926);
nor U10125 (N_10125,N_9984,N_9972);
or U10126 (N_10126,N_9990,N_9928);
or U10127 (N_10127,N_9995,N_9915);
nand U10128 (N_10128,N_9883,N_9976);
or U10129 (N_10129,N_9894,N_9971);
or U10130 (N_10130,N_9864,N_9959);
nor U10131 (N_10131,N_9823,N_9828);
nor U10132 (N_10132,N_9804,N_9956);
or U10133 (N_10133,N_9890,N_9923);
and U10134 (N_10134,N_9849,N_9889);
nand U10135 (N_10135,N_9885,N_9992);
and U10136 (N_10136,N_9870,N_9862);
nor U10137 (N_10137,N_9996,N_9992);
nand U10138 (N_10138,N_9942,N_9897);
xor U10139 (N_10139,N_9948,N_9981);
and U10140 (N_10140,N_9988,N_9885);
or U10141 (N_10141,N_9985,N_9907);
and U10142 (N_10142,N_9861,N_9824);
or U10143 (N_10143,N_9859,N_9806);
nor U10144 (N_10144,N_9890,N_9981);
nor U10145 (N_10145,N_9933,N_9855);
nor U10146 (N_10146,N_9947,N_9953);
and U10147 (N_10147,N_9888,N_9832);
and U10148 (N_10148,N_9854,N_9887);
nand U10149 (N_10149,N_9904,N_9816);
and U10150 (N_10150,N_9880,N_9918);
nor U10151 (N_10151,N_9984,N_9934);
and U10152 (N_10152,N_9917,N_9879);
xor U10153 (N_10153,N_9905,N_9962);
nand U10154 (N_10154,N_9981,N_9817);
and U10155 (N_10155,N_9888,N_9890);
and U10156 (N_10156,N_9967,N_9890);
nor U10157 (N_10157,N_9913,N_9826);
nand U10158 (N_10158,N_9935,N_9887);
nor U10159 (N_10159,N_9802,N_9913);
nand U10160 (N_10160,N_9879,N_9945);
and U10161 (N_10161,N_9959,N_9956);
nand U10162 (N_10162,N_9877,N_9829);
nor U10163 (N_10163,N_9815,N_9816);
nand U10164 (N_10164,N_9860,N_9909);
nor U10165 (N_10165,N_9815,N_9940);
and U10166 (N_10166,N_9800,N_9928);
and U10167 (N_10167,N_9898,N_9866);
and U10168 (N_10168,N_9946,N_9941);
nand U10169 (N_10169,N_9820,N_9844);
nand U10170 (N_10170,N_9860,N_9918);
nor U10171 (N_10171,N_9974,N_9940);
or U10172 (N_10172,N_9877,N_9935);
or U10173 (N_10173,N_9802,N_9853);
or U10174 (N_10174,N_9985,N_9822);
and U10175 (N_10175,N_9903,N_9933);
nand U10176 (N_10176,N_9990,N_9904);
and U10177 (N_10177,N_9922,N_9851);
and U10178 (N_10178,N_9973,N_9919);
nor U10179 (N_10179,N_9896,N_9948);
or U10180 (N_10180,N_9840,N_9808);
and U10181 (N_10181,N_9933,N_9817);
nor U10182 (N_10182,N_9804,N_9929);
nand U10183 (N_10183,N_9941,N_9816);
nand U10184 (N_10184,N_9992,N_9938);
nand U10185 (N_10185,N_9993,N_9963);
or U10186 (N_10186,N_9936,N_9960);
nand U10187 (N_10187,N_9883,N_9945);
and U10188 (N_10188,N_9904,N_9935);
nand U10189 (N_10189,N_9863,N_9945);
nor U10190 (N_10190,N_9974,N_9890);
and U10191 (N_10191,N_9988,N_9900);
or U10192 (N_10192,N_9998,N_9947);
nand U10193 (N_10193,N_9870,N_9943);
nor U10194 (N_10194,N_9828,N_9922);
or U10195 (N_10195,N_9999,N_9949);
nand U10196 (N_10196,N_9844,N_9992);
or U10197 (N_10197,N_9858,N_9941);
xor U10198 (N_10198,N_9835,N_9885);
or U10199 (N_10199,N_9957,N_9888);
and U10200 (N_10200,N_10183,N_10176);
nand U10201 (N_10201,N_10088,N_10083);
nand U10202 (N_10202,N_10055,N_10085);
and U10203 (N_10203,N_10078,N_10033);
or U10204 (N_10204,N_10052,N_10080);
or U10205 (N_10205,N_10042,N_10061);
and U10206 (N_10206,N_10192,N_10063);
nor U10207 (N_10207,N_10199,N_10186);
nor U10208 (N_10208,N_10058,N_10056);
nor U10209 (N_10209,N_10006,N_10066);
or U10210 (N_10210,N_10030,N_10126);
or U10211 (N_10211,N_10004,N_10079);
and U10212 (N_10212,N_10068,N_10067);
nor U10213 (N_10213,N_10048,N_10188);
nor U10214 (N_10214,N_10040,N_10159);
nor U10215 (N_10215,N_10156,N_10144);
nor U10216 (N_10216,N_10106,N_10029);
and U10217 (N_10217,N_10115,N_10099);
nand U10218 (N_10218,N_10170,N_10046);
or U10219 (N_10219,N_10191,N_10023);
nand U10220 (N_10220,N_10034,N_10095);
nor U10221 (N_10221,N_10002,N_10054);
and U10222 (N_10222,N_10094,N_10032);
and U10223 (N_10223,N_10185,N_10158);
or U10224 (N_10224,N_10091,N_10049);
or U10225 (N_10225,N_10139,N_10116);
and U10226 (N_10226,N_10178,N_10124);
nor U10227 (N_10227,N_10028,N_10177);
or U10228 (N_10228,N_10018,N_10064);
or U10229 (N_10229,N_10130,N_10133);
or U10230 (N_10230,N_10117,N_10082);
and U10231 (N_10231,N_10003,N_10146);
nand U10232 (N_10232,N_10024,N_10044);
or U10233 (N_10233,N_10041,N_10057);
or U10234 (N_10234,N_10069,N_10093);
or U10235 (N_10235,N_10059,N_10107);
and U10236 (N_10236,N_10108,N_10123);
and U10237 (N_10237,N_10149,N_10071);
nor U10238 (N_10238,N_10167,N_10008);
nand U10239 (N_10239,N_10165,N_10189);
nand U10240 (N_10240,N_10171,N_10051);
and U10241 (N_10241,N_10053,N_10137);
and U10242 (N_10242,N_10136,N_10015);
nor U10243 (N_10243,N_10025,N_10169);
nand U10244 (N_10244,N_10087,N_10035);
nor U10245 (N_10245,N_10162,N_10145);
and U10246 (N_10246,N_10112,N_10160);
xor U10247 (N_10247,N_10007,N_10090);
or U10248 (N_10248,N_10072,N_10198);
nor U10249 (N_10249,N_10140,N_10077);
or U10250 (N_10250,N_10118,N_10001);
xnor U10251 (N_10251,N_10005,N_10122);
nor U10252 (N_10252,N_10142,N_10036);
nand U10253 (N_10253,N_10027,N_10075);
or U10254 (N_10254,N_10163,N_10148);
and U10255 (N_10255,N_10017,N_10179);
nand U10256 (N_10256,N_10070,N_10184);
nand U10257 (N_10257,N_10089,N_10104);
and U10258 (N_10258,N_10010,N_10153);
nor U10259 (N_10259,N_10060,N_10021);
or U10260 (N_10260,N_10138,N_10076);
and U10261 (N_10261,N_10012,N_10000);
nand U10262 (N_10262,N_10154,N_10196);
or U10263 (N_10263,N_10073,N_10098);
or U10264 (N_10264,N_10019,N_10097);
nand U10265 (N_10265,N_10150,N_10151);
or U10266 (N_10266,N_10141,N_10074);
nor U10267 (N_10267,N_10047,N_10043);
nand U10268 (N_10268,N_10172,N_10194);
or U10269 (N_10269,N_10180,N_10131);
and U10270 (N_10270,N_10084,N_10157);
nor U10271 (N_10271,N_10197,N_10020);
and U10272 (N_10272,N_10110,N_10164);
nand U10273 (N_10273,N_10038,N_10014);
or U10274 (N_10274,N_10190,N_10081);
nor U10275 (N_10275,N_10100,N_10135);
and U10276 (N_10276,N_10011,N_10101);
nor U10277 (N_10277,N_10120,N_10129);
or U10278 (N_10278,N_10013,N_10173);
or U10279 (N_10279,N_10121,N_10195);
and U10280 (N_10280,N_10187,N_10062);
or U10281 (N_10281,N_10125,N_10127);
nand U10282 (N_10282,N_10050,N_10119);
nand U10283 (N_10283,N_10147,N_10128);
nand U10284 (N_10284,N_10134,N_10182);
nor U10285 (N_10285,N_10175,N_10065);
or U10286 (N_10286,N_10166,N_10009);
nand U10287 (N_10287,N_10037,N_10109);
and U10288 (N_10288,N_10152,N_10031);
nand U10289 (N_10289,N_10096,N_10155);
and U10290 (N_10290,N_10045,N_10113);
nor U10291 (N_10291,N_10161,N_10039);
or U10292 (N_10292,N_10103,N_10181);
nor U10293 (N_10293,N_10022,N_10168);
or U10294 (N_10294,N_10105,N_10026);
and U10295 (N_10295,N_10111,N_10174);
nor U10296 (N_10296,N_10086,N_10132);
or U10297 (N_10297,N_10114,N_10092);
nor U10298 (N_10298,N_10016,N_10102);
nor U10299 (N_10299,N_10143,N_10193);
and U10300 (N_10300,N_10086,N_10166);
or U10301 (N_10301,N_10046,N_10007);
or U10302 (N_10302,N_10028,N_10031);
and U10303 (N_10303,N_10129,N_10107);
nor U10304 (N_10304,N_10059,N_10182);
nor U10305 (N_10305,N_10121,N_10018);
nand U10306 (N_10306,N_10049,N_10147);
nand U10307 (N_10307,N_10090,N_10171);
nor U10308 (N_10308,N_10052,N_10146);
and U10309 (N_10309,N_10125,N_10006);
and U10310 (N_10310,N_10064,N_10077);
and U10311 (N_10311,N_10174,N_10127);
and U10312 (N_10312,N_10096,N_10124);
nor U10313 (N_10313,N_10065,N_10106);
nand U10314 (N_10314,N_10152,N_10190);
and U10315 (N_10315,N_10170,N_10054);
and U10316 (N_10316,N_10137,N_10196);
nor U10317 (N_10317,N_10055,N_10187);
nand U10318 (N_10318,N_10193,N_10013);
nor U10319 (N_10319,N_10073,N_10102);
or U10320 (N_10320,N_10079,N_10002);
and U10321 (N_10321,N_10101,N_10149);
nand U10322 (N_10322,N_10152,N_10115);
or U10323 (N_10323,N_10017,N_10072);
nand U10324 (N_10324,N_10062,N_10039);
nand U10325 (N_10325,N_10026,N_10100);
nor U10326 (N_10326,N_10167,N_10043);
nand U10327 (N_10327,N_10102,N_10108);
or U10328 (N_10328,N_10092,N_10179);
and U10329 (N_10329,N_10043,N_10165);
nor U10330 (N_10330,N_10057,N_10085);
nor U10331 (N_10331,N_10021,N_10034);
or U10332 (N_10332,N_10166,N_10094);
nor U10333 (N_10333,N_10181,N_10153);
and U10334 (N_10334,N_10040,N_10160);
or U10335 (N_10335,N_10097,N_10067);
nor U10336 (N_10336,N_10180,N_10055);
nand U10337 (N_10337,N_10073,N_10112);
nor U10338 (N_10338,N_10199,N_10178);
xnor U10339 (N_10339,N_10014,N_10015);
xor U10340 (N_10340,N_10123,N_10112);
nand U10341 (N_10341,N_10168,N_10098);
nor U10342 (N_10342,N_10179,N_10068);
and U10343 (N_10343,N_10186,N_10022);
nor U10344 (N_10344,N_10055,N_10048);
or U10345 (N_10345,N_10188,N_10173);
and U10346 (N_10346,N_10085,N_10003);
and U10347 (N_10347,N_10082,N_10015);
xor U10348 (N_10348,N_10010,N_10150);
nand U10349 (N_10349,N_10133,N_10069);
nor U10350 (N_10350,N_10059,N_10027);
nor U10351 (N_10351,N_10179,N_10160);
nand U10352 (N_10352,N_10009,N_10143);
nor U10353 (N_10353,N_10014,N_10100);
nand U10354 (N_10354,N_10122,N_10194);
nand U10355 (N_10355,N_10040,N_10060);
nor U10356 (N_10356,N_10091,N_10116);
or U10357 (N_10357,N_10066,N_10104);
nor U10358 (N_10358,N_10137,N_10165);
or U10359 (N_10359,N_10079,N_10151);
and U10360 (N_10360,N_10188,N_10081);
nor U10361 (N_10361,N_10117,N_10035);
nand U10362 (N_10362,N_10079,N_10139);
xor U10363 (N_10363,N_10031,N_10082);
nor U10364 (N_10364,N_10050,N_10010);
or U10365 (N_10365,N_10150,N_10003);
nand U10366 (N_10366,N_10060,N_10165);
or U10367 (N_10367,N_10161,N_10095);
or U10368 (N_10368,N_10127,N_10151);
or U10369 (N_10369,N_10050,N_10177);
or U10370 (N_10370,N_10097,N_10070);
nor U10371 (N_10371,N_10084,N_10094);
and U10372 (N_10372,N_10008,N_10180);
or U10373 (N_10373,N_10088,N_10043);
or U10374 (N_10374,N_10193,N_10195);
nor U10375 (N_10375,N_10196,N_10041);
xnor U10376 (N_10376,N_10037,N_10024);
and U10377 (N_10377,N_10043,N_10046);
nor U10378 (N_10378,N_10133,N_10159);
nor U10379 (N_10379,N_10174,N_10160);
and U10380 (N_10380,N_10118,N_10141);
xnor U10381 (N_10381,N_10048,N_10025);
and U10382 (N_10382,N_10013,N_10052);
or U10383 (N_10383,N_10080,N_10179);
xor U10384 (N_10384,N_10078,N_10180);
nand U10385 (N_10385,N_10007,N_10001);
and U10386 (N_10386,N_10093,N_10025);
or U10387 (N_10387,N_10140,N_10130);
nor U10388 (N_10388,N_10156,N_10060);
or U10389 (N_10389,N_10026,N_10081);
nand U10390 (N_10390,N_10105,N_10113);
or U10391 (N_10391,N_10048,N_10177);
or U10392 (N_10392,N_10106,N_10150);
nand U10393 (N_10393,N_10008,N_10163);
or U10394 (N_10394,N_10059,N_10066);
nor U10395 (N_10395,N_10010,N_10177);
or U10396 (N_10396,N_10128,N_10198);
nand U10397 (N_10397,N_10177,N_10155);
and U10398 (N_10398,N_10104,N_10065);
and U10399 (N_10399,N_10024,N_10124);
and U10400 (N_10400,N_10287,N_10320);
nand U10401 (N_10401,N_10209,N_10351);
or U10402 (N_10402,N_10387,N_10348);
nand U10403 (N_10403,N_10262,N_10215);
nor U10404 (N_10404,N_10272,N_10370);
nor U10405 (N_10405,N_10278,N_10355);
and U10406 (N_10406,N_10396,N_10365);
and U10407 (N_10407,N_10301,N_10395);
nand U10408 (N_10408,N_10399,N_10205);
or U10409 (N_10409,N_10283,N_10288);
or U10410 (N_10410,N_10390,N_10362);
and U10411 (N_10411,N_10290,N_10207);
nor U10412 (N_10412,N_10391,N_10359);
nor U10413 (N_10413,N_10344,N_10393);
nand U10414 (N_10414,N_10200,N_10233);
or U10415 (N_10415,N_10254,N_10219);
nand U10416 (N_10416,N_10269,N_10389);
nand U10417 (N_10417,N_10237,N_10228);
nand U10418 (N_10418,N_10268,N_10230);
and U10419 (N_10419,N_10314,N_10336);
xor U10420 (N_10420,N_10379,N_10308);
or U10421 (N_10421,N_10236,N_10241);
nand U10422 (N_10422,N_10222,N_10211);
nand U10423 (N_10423,N_10274,N_10253);
nor U10424 (N_10424,N_10322,N_10339);
and U10425 (N_10425,N_10234,N_10243);
or U10426 (N_10426,N_10252,N_10276);
nor U10427 (N_10427,N_10358,N_10306);
nor U10428 (N_10428,N_10334,N_10335);
nor U10429 (N_10429,N_10353,N_10338);
or U10430 (N_10430,N_10307,N_10385);
or U10431 (N_10431,N_10225,N_10251);
and U10432 (N_10432,N_10261,N_10238);
nor U10433 (N_10433,N_10206,N_10388);
or U10434 (N_10434,N_10330,N_10375);
nand U10435 (N_10435,N_10323,N_10342);
nand U10436 (N_10436,N_10332,N_10352);
or U10437 (N_10437,N_10328,N_10369);
nand U10438 (N_10438,N_10394,N_10376);
xnor U10439 (N_10439,N_10216,N_10302);
nand U10440 (N_10440,N_10366,N_10231);
and U10441 (N_10441,N_10373,N_10380);
nand U10442 (N_10442,N_10255,N_10360);
or U10443 (N_10443,N_10232,N_10305);
nor U10444 (N_10444,N_10277,N_10291);
nor U10445 (N_10445,N_10368,N_10246);
nor U10446 (N_10446,N_10284,N_10245);
nor U10447 (N_10447,N_10208,N_10279);
or U10448 (N_10448,N_10235,N_10213);
nand U10449 (N_10449,N_10350,N_10220);
nand U10450 (N_10450,N_10265,N_10226);
nand U10451 (N_10451,N_10313,N_10247);
and U10452 (N_10452,N_10324,N_10367);
and U10453 (N_10453,N_10303,N_10217);
or U10454 (N_10454,N_10372,N_10240);
and U10455 (N_10455,N_10286,N_10341);
nor U10456 (N_10456,N_10212,N_10346);
nor U10457 (N_10457,N_10318,N_10383);
and U10458 (N_10458,N_10321,N_10386);
nand U10459 (N_10459,N_10271,N_10275);
and U10460 (N_10460,N_10343,N_10333);
and U10461 (N_10461,N_10382,N_10257);
or U10462 (N_10462,N_10293,N_10221);
and U10463 (N_10463,N_10239,N_10300);
nand U10464 (N_10464,N_10248,N_10292);
nor U10465 (N_10465,N_10317,N_10282);
and U10466 (N_10466,N_10256,N_10381);
and U10467 (N_10467,N_10357,N_10273);
and U10468 (N_10468,N_10250,N_10227);
nand U10469 (N_10469,N_10223,N_10263);
or U10470 (N_10470,N_10270,N_10326);
nand U10471 (N_10471,N_10378,N_10316);
or U10472 (N_10472,N_10363,N_10319);
and U10473 (N_10473,N_10364,N_10304);
and U10474 (N_10474,N_10202,N_10204);
and U10475 (N_10475,N_10224,N_10377);
or U10476 (N_10476,N_10214,N_10297);
nand U10477 (N_10477,N_10354,N_10285);
nand U10478 (N_10478,N_10249,N_10294);
nand U10479 (N_10479,N_10210,N_10258);
and U10480 (N_10480,N_10242,N_10259);
or U10481 (N_10481,N_10289,N_10356);
and U10482 (N_10482,N_10374,N_10311);
and U10483 (N_10483,N_10299,N_10203);
or U10484 (N_10484,N_10371,N_10296);
and U10485 (N_10485,N_10309,N_10312);
and U10486 (N_10486,N_10267,N_10340);
nor U10487 (N_10487,N_10345,N_10337);
nand U10488 (N_10488,N_10260,N_10331);
nand U10489 (N_10489,N_10264,N_10315);
nand U10490 (N_10490,N_10398,N_10201);
or U10491 (N_10491,N_10298,N_10397);
or U10492 (N_10492,N_10347,N_10295);
nand U10493 (N_10493,N_10266,N_10281);
and U10494 (N_10494,N_10361,N_10280);
or U10495 (N_10495,N_10349,N_10384);
or U10496 (N_10496,N_10218,N_10310);
nand U10497 (N_10497,N_10327,N_10325);
or U10498 (N_10498,N_10329,N_10244);
nor U10499 (N_10499,N_10229,N_10392);
nor U10500 (N_10500,N_10294,N_10261);
nand U10501 (N_10501,N_10341,N_10362);
or U10502 (N_10502,N_10368,N_10276);
and U10503 (N_10503,N_10315,N_10226);
or U10504 (N_10504,N_10340,N_10334);
nor U10505 (N_10505,N_10377,N_10308);
and U10506 (N_10506,N_10351,N_10288);
or U10507 (N_10507,N_10298,N_10288);
nand U10508 (N_10508,N_10235,N_10225);
and U10509 (N_10509,N_10344,N_10383);
nand U10510 (N_10510,N_10220,N_10259);
or U10511 (N_10511,N_10204,N_10357);
nor U10512 (N_10512,N_10339,N_10264);
nand U10513 (N_10513,N_10364,N_10328);
and U10514 (N_10514,N_10395,N_10321);
nor U10515 (N_10515,N_10334,N_10260);
or U10516 (N_10516,N_10345,N_10257);
and U10517 (N_10517,N_10242,N_10206);
or U10518 (N_10518,N_10218,N_10266);
or U10519 (N_10519,N_10245,N_10272);
and U10520 (N_10520,N_10370,N_10271);
nor U10521 (N_10521,N_10294,N_10347);
and U10522 (N_10522,N_10386,N_10303);
nor U10523 (N_10523,N_10212,N_10348);
nor U10524 (N_10524,N_10285,N_10210);
nand U10525 (N_10525,N_10339,N_10228);
and U10526 (N_10526,N_10249,N_10316);
and U10527 (N_10527,N_10247,N_10232);
nand U10528 (N_10528,N_10352,N_10206);
and U10529 (N_10529,N_10223,N_10347);
and U10530 (N_10530,N_10292,N_10378);
nand U10531 (N_10531,N_10273,N_10366);
and U10532 (N_10532,N_10204,N_10267);
nor U10533 (N_10533,N_10368,N_10295);
or U10534 (N_10534,N_10362,N_10219);
or U10535 (N_10535,N_10232,N_10231);
and U10536 (N_10536,N_10366,N_10286);
nor U10537 (N_10537,N_10391,N_10297);
or U10538 (N_10538,N_10303,N_10268);
nand U10539 (N_10539,N_10304,N_10260);
nor U10540 (N_10540,N_10332,N_10233);
or U10541 (N_10541,N_10389,N_10267);
nand U10542 (N_10542,N_10211,N_10322);
and U10543 (N_10543,N_10208,N_10302);
nand U10544 (N_10544,N_10335,N_10256);
nor U10545 (N_10545,N_10260,N_10253);
nor U10546 (N_10546,N_10206,N_10308);
or U10547 (N_10547,N_10270,N_10327);
or U10548 (N_10548,N_10268,N_10296);
xor U10549 (N_10549,N_10371,N_10220);
nor U10550 (N_10550,N_10367,N_10243);
and U10551 (N_10551,N_10206,N_10244);
or U10552 (N_10552,N_10224,N_10357);
nand U10553 (N_10553,N_10348,N_10272);
nor U10554 (N_10554,N_10294,N_10388);
or U10555 (N_10555,N_10206,N_10378);
xor U10556 (N_10556,N_10294,N_10221);
or U10557 (N_10557,N_10304,N_10243);
and U10558 (N_10558,N_10335,N_10227);
nor U10559 (N_10559,N_10209,N_10293);
nor U10560 (N_10560,N_10272,N_10262);
nand U10561 (N_10561,N_10247,N_10264);
or U10562 (N_10562,N_10280,N_10246);
and U10563 (N_10563,N_10360,N_10310);
nor U10564 (N_10564,N_10336,N_10328);
and U10565 (N_10565,N_10288,N_10239);
nor U10566 (N_10566,N_10240,N_10239);
nor U10567 (N_10567,N_10321,N_10293);
nand U10568 (N_10568,N_10300,N_10287);
and U10569 (N_10569,N_10346,N_10250);
and U10570 (N_10570,N_10203,N_10284);
nand U10571 (N_10571,N_10388,N_10218);
and U10572 (N_10572,N_10375,N_10353);
nor U10573 (N_10573,N_10311,N_10207);
nand U10574 (N_10574,N_10243,N_10263);
and U10575 (N_10575,N_10263,N_10209);
or U10576 (N_10576,N_10263,N_10233);
nand U10577 (N_10577,N_10353,N_10293);
or U10578 (N_10578,N_10387,N_10227);
nand U10579 (N_10579,N_10363,N_10322);
nor U10580 (N_10580,N_10202,N_10227);
or U10581 (N_10581,N_10228,N_10315);
nor U10582 (N_10582,N_10331,N_10350);
and U10583 (N_10583,N_10202,N_10393);
and U10584 (N_10584,N_10395,N_10305);
nand U10585 (N_10585,N_10236,N_10232);
nor U10586 (N_10586,N_10264,N_10242);
and U10587 (N_10587,N_10213,N_10374);
and U10588 (N_10588,N_10381,N_10230);
nand U10589 (N_10589,N_10292,N_10202);
or U10590 (N_10590,N_10336,N_10394);
nand U10591 (N_10591,N_10307,N_10311);
or U10592 (N_10592,N_10220,N_10359);
nand U10593 (N_10593,N_10207,N_10294);
nand U10594 (N_10594,N_10293,N_10206);
or U10595 (N_10595,N_10385,N_10306);
nand U10596 (N_10596,N_10203,N_10210);
or U10597 (N_10597,N_10355,N_10386);
and U10598 (N_10598,N_10357,N_10307);
nor U10599 (N_10599,N_10225,N_10210);
nand U10600 (N_10600,N_10518,N_10494);
xor U10601 (N_10601,N_10484,N_10568);
and U10602 (N_10602,N_10434,N_10403);
nand U10603 (N_10603,N_10407,N_10551);
nand U10604 (N_10604,N_10556,N_10510);
nand U10605 (N_10605,N_10445,N_10496);
nor U10606 (N_10606,N_10537,N_10454);
nand U10607 (N_10607,N_10536,N_10413);
nor U10608 (N_10608,N_10500,N_10583);
nor U10609 (N_10609,N_10559,N_10450);
nor U10610 (N_10610,N_10419,N_10433);
nand U10611 (N_10611,N_10520,N_10581);
nor U10612 (N_10612,N_10452,N_10401);
nor U10613 (N_10613,N_10589,N_10592);
and U10614 (N_10614,N_10491,N_10539);
nor U10615 (N_10615,N_10548,N_10572);
nor U10616 (N_10616,N_10406,N_10410);
and U10617 (N_10617,N_10471,N_10579);
or U10618 (N_10618,N_10501,N_10486);
nand U10619 (N_10619,N_10550,N_10545);
nor U10620 (N_10620,N_10405,N_10593);
nor U10621 (N_10621,N_10584,N_10522);
nor U10622 (N_10622,N_10553,N_10473);
or U10623 (N_10623,N_10586,N_10482);
or U10624 (N_10624,N_10570,N_10458);
and U10625 (N_10625,N_10532,N_10483);
xor U10626 (N_10626,N_10495,N_10465);
and U10627 (N_10627,N_10428,N_10513);
or U10628 (N_10628,N_10498,N_10489);
and U10629 (N_10629,N_10467,N_10426);
or U10630 (N_10630,N_10439,N_10488);
nor U10631 (N_10631,N_10567,N_10578);
and U10632 (N_10632,N_10460,N_10540);
nor U10633 (N_10633,N_10464,N_10590);
nor U10634 (N_10634,N_10475,N_10552);
or U10635 (N_10635,N_10427,N_10456);
and U10636 (N_10636,N_10443,N_10555);
xnor U10637 (N_10637,N_10577,N_10447);
and U10638 (N_10638,N_10431,N_10425);
nor U10639 (N_10639,N_10566,N_10504);
or U10640 (N_10640,N_10507,N_10526);
nor U10641 (N_10641,N_10565,N_10474);
or U10642 (N_10642,N_10525,N_10462);
nand U10643 (N_10643,N_10511,N_10476);
nand U10644 (N_10644,N_10595,N_10517);
nor U10645 (N_10645,N_10497,N_10446);
and U10646 (N_10646,N_10422,N_10492);
nor U10647 (N_10647,N_10530,N_10412);
or U10648 (N_10648,N_10562,N_10594);
and U10649 (N_10649,N_10499,N_10575);
nor U10650 (N_10650,N_10541,N_10527);
and U10651 (N_10651,N_10453,N_10466);
and U10652 (N_10652,N_10529,N_10506);
and U10653 (N_10653,N_10404,N_10429);
or U10654 (N_10654,N_10435,N_10535);
nor U10655 (N_10655,N_10569,N_10521);
nand U10656 (N_10656,N_10424,N_10547);
or U10657 (N_10657,N_10480,N_10432);
nand U10658 (N_10658,N_10418,N_10416);
xor U10659 (N_10659,N_10463,N_10417);
and U10660 (N_10660,N_10596,N_10508);
or U10661 (N_10661,N_10533,N_10534);
nor U10662 (N_10662,N_10469,N_10437);
or U10663 (N_10663,N_10414,N_10479);
nand U10664 (N_10664,N_10430,N_10451);
nor U10665 (N_10665,N_10523,N_10591);
xnor U10666 (N_10666,N_10524,N_10576);
or U10667 (N_10667,N_10438,N_10444);
nor U10668 (N_10668,N_10448,N_10481);
and U10669 (N_10669,N_10561,N_10485);
nor U10670 (N_10670,N_10538,N_10490);
and U10671 (N_10671,N_10516,N_10574);
nand U10672 (N_10672,N_10449,N_10509);
or U10673 (N_10673,N_10420,N_10477);
or U10674 (N_10674,N_10487,N_10571);
nand U10675 (N_10675,N_10441,N_10580);
or U10676 (N_10676,N_10546,N_10515);
and U10677 (N_10677,N_10436,N_10457);
nand U10678 (N_10678,N_10472,N_10470);
nor U10679 (N_10679,N_10599,N_10461);
nand U10680 (N_10680,N_10502,N_10543);
nor U10681 (N_10681,N_10531,N_10459);
nand U10682 (N_10682,N_10503,N_10585);
and U10683 (N_10683,N_10493,N_10442);
nor U10684 (N_10684,N_10421,N_10549);
nand U10685 (N_10685,N_10408,N_10588);
nor U10686 (N_10686,N_10542,N_10557);
and U10687 (N_10687,N_10587,N_10582);
and U10688 (N_10688,N_10400,N_10598);
nor U10689 (N_10689,N_10560,N_10519);
xnor U10690 (N_10690,N_10440,N_10564);
or U10691 (N_10691,N_10554,N_10528);
nand U10692 (N_10692,N_10402,N_10558);
or U10693 (N_10693,N_10415,N_10411);
nor U10694 (N_10694,N_10544,N_10409);
nor U10695 (N_10695,N_10478,N_10455);
and U10696 (N_10696,N_10505,N_10597);
or U10697 (N_10697,N_10573,N_10468);
nand U10698 (N_10698,N_10512,N_10514);
nor U10699 (N_10699,N_10563,N_10423);
nand U10700 (N_10700,N_10505,N_10464);
nor U10701 (N_10701,N_10430,N_10524);
or U10702 (N_10702,N_10599,N_10478);
nand U10703 (N_10703,N_10452,N_10543);
nand U10704 (N_10704,N_10582,N_10454);
and U10705 (N_10705,N_10434,N_10575);
nor U10706 (N_10706,N_10573,N_10561);
and U10707 (N_10707,N_10478,N_10486);
nor U10708 (N_10708,N_10443,N_10445);
nand U10709 (N_10709,N_10561,N_10482);
nand U10710 (N_10710,N_10511,N_10591);
and U10711 (N_10711,N_10534,N_10544);
or U10712 (N_10712,N_10544,N_10593);
nor U10713 (N_10713,N_10584,N_10512);
nor U10714 (N_10714,N_10432,N_10576);
nor U10715 (N_10715,N_10486,N_10477);
or U10716 (N_10716,N_10400,N_10425);
or U10717 (N_10717,N_10467,N_10506);
nand U10718 (N_10718,N_10556,N_10551);
or U10719 (N_10719,N_10404,N_10414);
or U10720 (N_10720,N_10457,N_10539);
and U10721 (N_10721,N_10434,N_10423);
xor U10722 (N_10722,N_10542,N_10420);
nand U10723 (N_10723,N_10450,N_10426);
or U10724 (N_10724,N_10584,N_10461);
nand U10725 (N_10725,N_10481,N_10422);
nor U10726 (N_10726,N_10401,N_10539);
and U10727 (N_10727,N_10480,N_10481);
nand U10728 (N_10728,N_10469,N_10473);
nand U10729 (N_10729,N_10552,N_10446);
and U10730 (N_10730,N_10483,N_10581);
nor U10731 (N_10731,N_10450,N_10471);
nand U10732 (N_10732,N_10487,N_10535);
nor U10733 (N_10733,N_10401,N_10540);
and U10734 (N_10734,N_10450,N_10451);
nor U10735 (N_10735,N_10571,N_10496);
and U10736 (N_10736,N_10592,N_10500);
and U10737 (N_10737,N_10570,N_10502);
and U10738 (N_10738,N_10597,N_10565);
and U10739 (N_10739,N_10456,N_10499);
nor U10740 (N_10740,N_10405,N_10433);
nor U10741 (N_10741,N_10549,N_10413);
and U10742 (N_10742,N_10507,N_10494);
nor U10743 (N_10743,N_10515,N_10564);
and U10744 (N_10744,N_10563,N_10531);
nand U10745 (N_10745,N_10451,N_10524);
nand U10746 (N_10746,N_10599,N_10417);
or U10747 (N_10747,N_10445,N_10562);
and U10748 (N_10748,N_10424,N_10508);
nand U10749 (N_10749,N_10547,N_10403);
nor U10750 (N_10750,N_10544,N_10581);
or U10751 (N_10751,N_10468,N_10459);
or U10752 (N_10752,N_10474,N_10480);
nor U10753 (N_10753,N_10482,N_10426);
nand U10754 (N_10754,N_10536,N_10423);
and U10755 (N_10755,N_10569,N_10527);
and U10756 (N_10756,N_10478,N_10546);
or U10757 (N_10757,N_10403,N_10489);
or U10758 (N_10758,N_10513,N_10522);
nand U10759 (N_10759,N_10433,N_10535);
nor U10760 (N_10760,N_10486,N_10548);
or U10761 (N_10761,N_10464,N_10496);
and U10762 (N_10762,N_10566,N_10544);
nor U10763 (N_10763,N_10560,N_10499);
or U10764 (N_10764,N_10532,N_10489);
and U10765 (N_10765,N_10431,N_10583);
and U10766 (N_10766,N_10473,N_10476);
nand U10767 (N_10767,N_10413,N_10466);
or U10768 (N_10768,N_10595,N_10555);
nand U10769 (N_10769,N_10599,N_10507);
or U10770 (N_10770,N_10500,N_10404);
and U10771 (N_10771,N_10486,N_10577);
nand U10772 (N_10772,N_10442,N_10531);
and U10773 (N_10773,N_10470,N_10428);
nand U10774 (N_10774,N_10470,N_10540);
or U10775 (N_10775,N_10445,N_10598);
and U10776 (N_10776,N_10583,N_10401);
or U10777 (N_10777,N_10427,N_10558);
nor U10778 (N_10778,N_10403,N_10549);
nand U10779 (N_10779,N_10523,N_10497);
and U10780 (N_10780,N_10592,N_10598);
nor U10781 (N_10781,N_10498,N_10499);
nand U10782 (N_10782,N_10477,N_10511);
nor U10783 (N_10783,N_10569,N_10485);
nor U10784 (N_10784,N_10577,N_10555);
nor U10785 (N_10785,N_10590,N_10450);
and U10786 (N_10786,N_10510,N_10444);
nand U10787 (N_10787,N_10462,N_10506);
and U10788 (N_10788,N_10570,N_10410);
nor U10789 (N_10789,N_10591,N_10468);
or U10790 (N_10790,N_10450,N_10594);
and U10791 (N_10791,N_10411,N_10568);
nor U10792 (N_10792,N_10503,N_10439);
and U10793 (N_10793,N_10595,N_10477);
and U10794 (N_10794,N_10412,N_10433);
and U10795 (N_10795,N_10498,N_10529);
or U10796 (N_10796,N_10472,N_10513);
or U10797 (N_10797,N_10466,N_10556);
or U10798 (N_10798,N_10533,N_10428);
nand U10799 (N_10799,N_10537,N_10503);
and U10800 (N_10800,N_10735,N_10630);
nor U10801 (N_10801,N_10673,N_10640);
or U10802 (N_10802,N_10760,N_10618);
nand U10803 (N_10803,N_10762,N_10773);
xnor U10804 (N_10804,N_10647,N_10662);
and U10805 (N_10805,N_10676,N_10753);
nand U10806 (N_10806,N_10686,N_10610);
and U10807 (N_10807,N_10786,N_10725);
or U10808 (N_10808,N_10653,N_10719);
or U10809 (N_10809,N_10732,N_10747);
and U10810 (N_10810,N_10778,N_10609);
and U10811 (N_10811,N_10720,N_10615);
and U10812 (N_10812,N_10613,N_10699);
or U10813 (N_10813,N_10777,N_10742);
nor U10814 (N_10814,N_10696,N_10632);
nor U10815 (N_10815,N_10757,N_10780);
nor U10816 (N_10816,N_10621,N_10769);
and U10817 (N_10817,N_10624,N_10741);
nor U10818 (N_10818,N_10669,N_10749);
nor U10819 (N_10819,N_10791,N_10694);
nand U10820 (N_10820,N_10603,N_10635);
nor U10821 (N_10821,N_10744,N_10756);
nand U10822 (N_10822,N_10681,N_10606);
nand U10823 (N_10823,N_10788,N_10770);
nor U10824 (N_10824,N_10767,N_10655);
nand U10825 (N_10825,N_10771,N_10710);
and U10826 (N_10826,N_10721,N_10690);
and U10827 (N_10827,N_10692,N_10759);
or U10828 (N_10828,N_10776,N_10703);
and U10829 (N_10829,N_10654,N_10712);
nor U10830 (N_10830,N_10600,N_10774);
nand U10831 (N_10831,N_10648,N_10665);
nor U10832 (N_10832,N_10693,N_10619);
and U10833 (N_10833,N_10734,N_10731);
nand U10834 (N_10834,N_10723,N_10738);
nand U10835 (N_10835,N_10628,N_10629);
nor U10836 (N_10836,N_10746,N_10718);
or U10837 (N_10837,N_10792,N_10722);
and U10838 (N_10838,N_10689,N_10781);
nand U10839 (N_10839,N_10709,N_10729);
nand U10840 (N_10840,N_10671,N_10768);
or U10841 (N_10841,N_10682,N_10638);
or U10842 (N_10842,N_10672,N_10684);
and U10843 (N_10843,N_10677,N_10795);
or U10844 (N_10844,N_10617,N_10737);
nor U10845 (N_10845,N_10755,N_10765);
or U10846 (N_10846,N_10704,N_10715);
or U10847 (N_10847,N_10761,N_10641);
nor U10848 (N_10848,N_10646,N_10797);
nor U10849 (N_10849,N_10724,N_10658);
xnor U10850 (N_10850,N_10775,N_10659);
and U10851 (N_10851,N_10651,N_10660);
and U10852 (N_10852,N_10740,N_10752);
or U10853 (N_10853,N_10708,N_10643);
nand U10854 (N_10854,N_10675,N_10796);
or U10855 (N_10855,N_10698,N_10697);
nor U10856 (N_10856,N_10605,N_10625);
and U10857 (N_10857,N_10645,N_10611);
nand U10858 (N_10858,N_10779,N_10656);
nand U10859 (N_10859,N_10649,N_10743);
or U10860 (N_10860,N_10644,N_10727);
nand U10861 (N_10861,N_10783,N_10639);
and U10862 (N_10862,N_10667,N_10631);
nand U10863 (N_10863,N_10634,N_10739);
nor U10864 (N_10864,N_10745,N_10763);
nand U10865 (N_10865,N_10793,N_10678);
nand U10866 (N_10866,N_10789,N_10730);
or U10867 (N_10867,N_10685,N_10716);
nand U10868 (N_10868,N_10754,N_10680);
nand U10869 (N_10869,N_10695,N_10706);
and U10870 (N_10870,N_10687,N_10799);
nand U10871 (N_10871,N_10620,N_10748);
and U10872 (N_10872,N_10612,N_10652);
nor U10873 (N_10873,N_10713,N_10794);
and U10874 (N_10874,N_10717,N_10764);
or U10875 (N_10875,N_10707,N_10758);
or U10876 (N_10876,N_10700,N_10627);
nor U10877 (N_10877,N_10782,N_10616);
and U10878 (N_10878,N_10601,N_10670);
or U10879 (N_10879,N_10679,N_10688);
nand U10880 (N_10880,N_10733,N_10657);
nand U10881 (N_10881,N_10608,N_10602);
and U10882 (N_10882,N_10728,N_10637);
nand U10883 (N_10883,N_10674,N_10623);
or U10884 (N_10884,N_10668,N_10772);
and U10885 (N_10885,N_10622,N_10750);
nand U10886 (N_10886,N_10798,N_10784);
nand U10887 (N_10887,N_10661,N_10691);
and U10888 (N_10888,N_10663,N_10702);
nor U10889 (N_10889,N_10705,N_10626);
and U10890 (N_10890,N_10650,N_10766);
and U10891 (N_10891,N_10790,N_10614);
and U10892 (N_10892,N_10664,N_10726);
or U10893 (N_10893,N_10736,N_10711);
or U10894 (N_10894,N_10666,N_10633);
nor U10895 (N_10895,N_10636,N_10607);
nand U10896 (N_10896,N_10642,N_10683);
or U10897 (N_10897,N_10785,N_10701);
nor U10898 (N_10898,N_10751,N_10787);
nor U10899 (N_10899,N_10714,N_10604);
and U10900 (N_10900,N_10717,N_10688);
and U10901 (N_10901,N_10633,N_10764);
nor U10902 (N_10902,N_10664,N_10634);
or U10903 (N_10903,N_10679,N_10749);
nor U10904 (N_10904,N_10708,N_10741);
nand U10905 (N_10905,N_10678,N_10642);
and U10906 (N_10906,N_10693,N_10712);
or U10907 (N_10907,N_10675,N_10755);
and U10908 (N_10908,N_10732,N_10671);
or U10909 (N_10909,N_10637,N_10780);
and U10910 (N_10910,N_10714,N_10727);
nor U10911 (N_10911,N_10641,N_10606);
nand U10912 (N_10912,N_10615,N_10750);
and U10913 (N_10913,N_10609,N_10610);
nor U10914 (N_10914,N_10755,N_10706);
or U10915 (N_10915,N_10747,N_10755);
nand U10916 (N_10916,N_10615,N_10634);
nand U10917 (N_10917,N_10710,N_10759);
and U10918 (N_10918,N_10707,N_10797);
nand U10919 (N_10919,N_10768,N_10636);
and U10920 (N_10920,N_10702,N_10693);
or U10921 (N_10921,N_10683,N_10664);
nand U10922 (N_10922,N_10753,N_10649);
nor U10923 (N_10923,N_10628,N_10799);
or U10924 (N_10924,N_10601,N_10785);
or U10925 (N_10925,N_10637,N_10783);
nand U10926 (N_10926,N_10798,N_10610);
or U10927 (N_10927,N_10642,N_10667);
xor U10928 (N_10928,N_10763,N_10681);
nand U10929 (N_10929,N_10700,N_10671);
or U10930 (N_10930,N_10652,N_10640);
or U10931 (N_10931,N_10668,N_10625);
and U10932 (N_10932,N_10681,N_10675);
nor U10933 (N_10933,N_10630,N_10733);
nor U10934 (N_10934,N_10669,N_10747);
or U10935 (N_10935,N_10759,N_10653);
and U10936 (N_10936,N_10749,N_10611);
or U10937 (N_10937,N_10794,N_10633);
and U10938 (N_10938,N_10684,N_10622);
or U10939 (N_10939,N_10781,N_10663);
and U10940 (N_10940,N_10677,N_10747);
and U10941 (N_10941,N_10697,N_10615);
and U10942 (N_10942,N_10612,N_10688);
nor U10943 (N_10943,N_10611,N_10633);
nor U10944 (N_10944,N_10625,N_10792);
or U10945 (N_10945,N_10730,N_10784);
nand U10946 (N_10946,N_10697,N_10621);
and U10947 (N_10947,N_10785,N_10758);
nor U10948 (N_10948,N_10631,N_10608);
and U10949 (N_10949,N_10601,N_10796);
or U10950 (N_10950,N_10704,N_10763);
and U10951 (N_10951,N_10625,N_10682);
nor U10952 (N_10952,N_10732,N_10621);
nor U10953 (N_10953,N_10680,N_10679);
or U10954 (N_10954,N_10735,N_10730);
or U10955 (N_10955,N_10728,N_10686);
nor U10956 (N_10956,N_10759,N_10736);
or U10957 (N_10957,N_10786,N_10676);
and U10958 (N_10958,N_10618,N_10619);
nand U10959 (N_10959,N_10743,N_10601);
or U10960 (N_10960,N_10717,N_10678);
and U10961 (N_10961,N_10690,N_10720);
and U10962 (N_10962,N_10665,N_10674);
nor U10963 (N_10963,N_10684,N_10654);
nor U10964 (N_10964,N_10760,N_10636);
or U10965 (N_10965,N_10667,N_10605);
or U10966 (N_10966,N_10759,N_10725);
or U10967 (N_10967,N_10718,N_10793);
and U10968 (N_10968,N_10677,N_10769);
and U10969 (N_10969,N_10618,N_10694);
nand U10970 (N_10970,N_10618,N_10631);
and U10971 (N_10971,N_10677,N_10755);
xnor U10972 (N_10972,N_10637,N_10719);
or U10973 (N_10973,N_10653,N_10710);
nand U10974 (N_10974,N_10737,N_10664);
nand U10975 (N_10975,N_10618,N_10673);
nor U10976 (N_10976,N_10693,N_10768);
or U10977 (N_10977,N_10726,N_10742);
and U10978 (N_10978,N_10735,N_10666);
or U10979 (N_10979,N_10766,N_10799);
nor U10980 (N_10980,N_10709,N_10688);
nand U10981 (N_10981,N_10749,N_10664);
nor U10982 (N_10982,N_10639,N_10659);
nand U10983 (N_10983,N_10693,N_10752);
nand U10984 (N_10984,N_10782,N_10730);
nor U10985 (N_10985,N_10715,N_10633);
xor U10986 (N_10986,N_10787,N_10747);
nor U10987 (N_10987,N_10664,N_10649);
or U10988 (N_10988,N_10660,N_10717);
or U10989 (N_10989,N_10646,N_10773);
and U10990 (N_10990,N_10747,N_10701);
or U10991 (N_10991,N_10701,N_10791);
nand U10992 (N_10992,N_10744,N_10609);
nand U10993 (N_10993,N_10725,N_10743);
and U10994 (N_10994,N_10682,N_10672);
or U10995 (N_10995,N_10695,N_10798);
or U10996 (N_10996,N_10707,N_10744);
or U10997 (N_10997,N_10678,N_10687);
and U10998 (N_10998,N_10711,N_10619);
nor U10999 (N_10999,N_10665,N_10609);
nand U11000 (N_11000,N_10990,N_10826);
or U11001 (N_11001,N_10930,N_10812);
nand U11002 (N_11002,N_10850,N_10925);
nand U11003 (N_11003,N_10848,N_10818);
nor U11004 (N_11004,N_10856,N_10940);
or U11005 (N_11005,N_10882,N_10912);
or U11006 (N_11006,N_10975,N_10891);
and U11007 (N_11007,N_10801,N_10811);
nor U11008 (N_11008,N_10987,N_10941);
xor U11009 (N_11009,N_10847,N_10837);
nor U11010 (N_11010,N_10867,N_10984);
and U11011 (N_11011,N_10851,N_10991);
and U11012 (N_11012,N_10905,N_10926);
nor U11013 (N_11013,N_10822,N_10995);
and U11014 (N_11014,N_10968,N_10982);
nor U11015 (N_11015,N_10932,N_10976);
and U11016 (N_11016,N_10810,N_10800);
nor U11017 (N_11017,N_10978,N_10808);
or U11018 (N_11018,N_10802,N_10960);
or U11019 (N_11019,N_10872,N_10832);
nand U11020 (N_11020,N_10804,N_10892);
and U11021 (N_11021,N_10927,N_10894);
nand U11022 (N_11022,N_10889,N_10883);
and U11023 (N_11023,N_10835,N_10899);
or U11024 (N_11024,N_10981,N_10942);
and U11025 (N_11025,N_10979,N_10996);
nand U11026 (N_11026,N_10859,N_10964);
nor U11027 (N_11027,N_10924,N_10920);
nor U11028 (N_11028,N_10913,N_10841);
xor U11029 (N_11029,N_10902,N_10819);
nand U11030 (N_11030,N_10877,N_10916);
nor U11031 (N_11031,N_10896,N_10852);
or U11032 (N_11032,N_10820,N_10962);
nand U11033 (N_11033,N_10831,N_10807);
nand U11034 (N_11034,N_10886,N_10988);
nand U11035 (N_11035,N_10961,N_10873);
or U11036 (N_11036,N_10907,N_10943);
nor U11037 (N_11037,N_10965,N_10885);
or U11038 (N_11038,N_10874,N_10897);
and U11039 (N_11039,N_10865,N_10842);
nand U11040 (N_11040,N_10906,N_10955);
and U11041 (N_11041,N_10983,N_10830);
or U11042 (N_11042,N_10838,N_10946);
nand U11043 (N_11043,N_10844,N_10898);
nand U11044 (N_11044,N_10936,N_10959);
or U11045 (N_11045,N_10803,N_10951);
nand U11046 (N_11046,N_10815,N_10845);
xnor U11047 (N_11047,N_10966,N_10824);
nor U11048 (N_11048,N_10862,N_10821);
nor U11049 (N_11049,N_10805,N_10895);
and U11050 (N_11050,N_10875,N_10993);
and U11051 (N_11051,N_10893,N_10997);
nor U11052 (N_11052,N_10828,N_10921);
and U11053 (N_11053,N_10937,N_10944);
nor U11054 (N_11054,N_10939,N_10958);
or U11055 (N_11055,N_10858,N_10827);
or U11056 (N_11056,N_10972,N_10854);
and U11057 (N_11057,N_10869,N_10910);
nor U11058 (N_11058,N_10911,N_10919);
and U11059 (N_11059,N_10881,N_10947);
nor U11060 (N_11060,N_10816,N_10908);
or U11061 (N_11061,N_10917,N_10934);
nor U11062 (N_11062,N_10878,N_10825);
and U11063 (N_11063,N_10949,N_10834);
or U11064 (N_11064,N_10853,N_10957);
and U11065 (N_11065,N_10971,N_10952);
nor U11066 (N_11066,N_10866,N_10863);
nor U11067 (N_11067,N_10823,N_10923);
nor U11068 (N_11068,N_10857,N_10843);
nand U11069 (N_11069,N_10948,N_10950);
nor U11070 (N_11070,N_10870,N_10829);
nand U11071 (N_11071,N_10840,N_10909);
and U11072 (N_11072,N_10806,N_10956);
nor U11073 (N_11073,N_10945,N_10880);
or U11074 (N_11074,N_10977,N_10900);
nor U11075 (N_11075,N_10914,N_10967);
nor U11076 (N_11076,N_10890,N_10922);
or U11077 (N_11077,N_10938,N_10985);
nand U11078 (N_11078,N_10833,N_10963);
or U11079 (N_11079,N_10836,N_10876);
nor U11080 (N_11080,N_10969,N_10999);
and U11081 (N_11081,N_10954,N_10970);
or U11082 (N_11082,N_10929,N_10980);
and U11083 (N_11083,N_10901,N_10868);
and U11084 (N_11084,N_10814,N_10974);
or U11085 (N_11085,N_10888,N_10903);
nand U11086 (N_11086,N_10933,N_10809);
nor U11087 (N_11087,N_10931,N_10864);
or U11088 (N_11088,N_10846,N_10855);
nand U11089 (N_11089,N_10871,N_10817);
nand U11090 (N_11090,N_10879,N_10992);
or U11091 (N_11091,N_10904,N_10973);
nor U11092 (N_11092,N_10849,N_10839);
nand U11093 (N_11093,N_10861,N_10887);
nand U11094 (N_11094,N_10953,N_10935);
or U11095 (N_11095,N_10884,N_10813);
nor U11096 (N_11096,N_10860,N_10986);
nor U11097 (N_11097,N_10989,N_10994);
or U11098 (N_11098,N_10915,N_10998);
nand U11099 (N_11099,N_10928,N_10918);
and U11100 (N_11100,N_10974,N_10800);
or U11101 (N_11101,N_10975,N_10915);
nor U11102 (N_11102,N_10929,N_10912);
nor U11103 (N_11103,N_10939,N_10940);
nor U11104 (N_11104,N_10828,N_10968);
nor U11105 (N_11105,N_10815,N_10854);
nand U11106 (N_11106,N_10816,N_10928);
or U11107 (N_11107,N_10944,N_10992);
and U11108 (N_11108,N_10837,N_10811);
or U11109 (N_11109,N_10821,N_10898);
or U11110 (N_11110,N_10841,N_10889);
or U11111 (N_11111,N_10820,N_10809);
or U11112 (N_11112,N_10920,N_10804);
nor U11113 (N_11113,N_10995,N_10800);
nand U11114 (N_11114,N_10893,N_10802);
nor U11115 (N_11115,N_10817,N_10984);
or U11116 (N_11116,N_10926,N_10850);
and U11117 (N_11117,N_10820,N_10841);
and U11118 (N_11118,N_10911,N_10802);
nand U11119 (N_11119,N_10896,N_10863);
or U11120 (N_11120,N_10959,N_10994);
and U11121 (N_11121,N_10969,N_10976);
or U11122 (N_11122,N_10963,N_10936);
nor U11123 (N_11123,N_10912,N_10957);
nand U11124 (N_11124,N_10909,N_10993);
xor U11125 (N_11125,N_10803,N_10812);
nor U11126 (N_11126,N_10806,N_10883);
nor U11127 (N_11127,N_10863,N_10977);
and U11128 (N_11128,N_10960,N_10920);
nand U11129 (N_11129,N_10877,N_10960);
nor U11130 (N_11130,N_10946,N_10897);
or U11131 (N_11131,N_10845,N_10990);
and U11132 (N_11132,N_10943,N_10920);
or U11133 (N_11133,N_10892,N_10942);
nor U11134 (N_11134,N_10897,N_10857);
nor U11135 (N_11135,N_10853,N_10998);
or U11136 (N_11136,N_10855,N_10875);
nor U11137 (N_11137,N_10841,N_10815);
and U11138 (N_11138,N_10968,N_10883);
nand U11139 (N_11139,N_10927,N_10986);
nor U11140 (N_11140,N_10944,N_10846);
or U11141 (N_11141,N_10821,N_10887);
or U11142 (N_11142,N_10996,N_10915);
or U11143 (N_11143,N_10986,N_10904);
or U11144 (N_11144,N_10986,N_10949);
and U11145 (N_11145,N_10924,N_10877);
nor U11146 (N_11146,N_10884,N_10832);
or U11147 (N_11147,N_10983,N_10895);
nand U11148 (N_11148,N_10804,N_10869);
and U11149 (N_11149,N_10955,N_10991);
nor U11150 (N_11150,N_10902,N_10963);
nand U11151 (N_11151,N_10831,N_10905);
nand U11152 (N_11152,N_10857,N_10823);
and U11153 (N_11153,N_10967,N_10913);
nand U11154 (N_11154,N_10903,N_10834);
or U11155 (N_11155,N_10864,N_10825);
nor U11156 (N_11156,N_10986,N_10831);
and U11157 (N_11157,N_10949,N_10895);
nor U11158 (N_11158,N_10951,N_10824);
and U11159 (N_11159,N_10809,N_10842);
nor U11160 (N_11160,N_10864,N_10885);
or U11161 (N_11161,N_10829,N_10804);
and U11162 (N_11162,N_10969,N_10820);
nor U11163 (N_11163,N_10895,N_10883);
nand U11164 (N_11164,N_10809,N_10993);
nand U11165 (N_11165,N_10996,N_10990);
nand U11166 (N_11166,N_10948,N_10986);
or U11167 (N_11167,N_10969,N_10913);
or U11168 (N_11168,N_10877,N_10861);
or U11169 (N_11169,N_10876,N_10980);
and U11170 (N_11170,N_10936,N_10983);
or U11171 (N_11171,N_10869,N_10984);
nand U11172 (N_11172,N_10976,N_10813);
and U11173 (N_11173,N_10876,N_10889);
or U11174 (N_11174,N_10922,N_10992);
nor U11175 (N_11175,N_10868,N_10969);
and U11176 (N_11176,N_10965,N_10871);
and U11177 (N_11177,N_10961,N_10807);
xnor U11178 (N_11178,N_10830,N_10902);
or U11179 (N_11179,N_10889,N_10976);
and U11180 (N_11180,N_10894,N_10960);
or U11181 (N_11181,N_10802,N_10923);
and U11182 (N_11182,N_10954,N_10842);
and U11183 (N_11183,N_10849,N_10898);
and U11184 (N_11184,N_10992,N_10915);
or U11185 (N_11185,N_10921,N_10812);
or U11186 (N_11186,N_10996,N_10886);
or U11187 (N_11187,N_10985,N_10837);
nand U11188 (N_11188,N_10949,N_10811);
nand U11189 (N_11189,N_10965,N_10817);
and U11190 (N_11190,N_10884,N_10985);
nor U11191 (N_11191,N_10989,N_10813);
nor U11192 (N_11192,N_10840,N_10926);
nand U11193 (N_11193,N_10948,N_10818);
or U11194 (N_11194,N_10831,N_10903);
nand U11195 (N_11195,N_10817,N_10819);
or U11196 (N_11196,N_10811,N_10991);
and U11197 (N_11197,N_10968,N_10808);
or U11198 (N_11198,N_10841,N_10927);
nor U11199 (N_11199,N_10828,N_10891);
nor U11200 (N_11200,N_11139,N_11054);
nand U11201 (N_11201,N_11153,N_11023);
and U11202 (N_11202,N_11081,N_11167);
nor U11203 (N_11203,N_11017,N_11003);
nand U11204 (N_11204,N_11118,N_11187);
nor U11205 (N_11205,N_11174,N_11095);
nor U11206 (N_11206,N_11058,N_11109);
nor U11207 (N_11207,N_11073,N_11159);
nor U11208 (N_11208,N_11063,N_11016);
nand U11209 (N_11209,N_11185,N_11028);
or U11210 (N_11210,N_11156,N_11101);
and U11211 (N_11211,N_11130,N_11088);
nand U11212 (N_11212,N_11078,N_11037);
and U11213 (N_11213,N_11050,N_11135);
nor U11214 (N_11214,N_11069,N_11123);
and U11215 (N_11215,N_11128,N_11131);
nor U11216 (N_11216,N_11198,N_11056);
and U11217 (N_11217,N_11029,N_11096);
or U11218 (N_11218,N_11090,N_11192);
or U11219 (N_11219,N_11154,N_11133);
and U11220 (N_11220,N_11002,N_11001);
nand U11221 (N_11221,N_11178,N_11147);
nand U11222 (N_11222,N_11195,N_11119);
and U11223 (N_11223,N_11146,N_11149);
or U11224 (N_11224,N_11022,N_11052);
nand U11225 (N_11225,N_11168,N_11074);
and U11226 (N_11226,N_11004,N_11160);
or U11227 (N_11227,N_11089,N_11100);
or U11228 (N_11228,N_11099,N_11181);
or U11229 (N_11229,N_11071,N_11025);
or U11230 (N_11230,N_11027,N_11068);
and U11231 (N_11231,N_11151,N_11102);
and U11232 (N_11232,N_11170,N_11018);
xor U11233 (N_11233,N_11110,N_11111);
or U11234 (N_11234,N_11083,N_11134);
and U11235 (N_11235,N_11082,N_11021);
and U11236 (N_11236,N_11136,N_11036);
nand U11237 (N_11237,N_11191,N_11094);
nor U11238 (N_11238,N_11152,N_11011);
or U11239 (N_11239,N_11010,N_11108);
nand U11240 (N_11240,N_11172,N_11044);
or U11241 (N_11241,N_11117,N_11049);
nand U11242 (N_11242,N_11066,N_11034);
nand U11243 (N_11243,N_11015,N_11144);
or U11244 (N_11244,N_11048,N_11196);
or U11245 (N_11245,N_11057,N_11105);
nand U11246 (N_11246,N_11177,N_11024);
or U11247 (N_11247,N_11114,N_11148);
or U11248 (N_11248,N_11098,N_11043);
nand U11249 (N_11249,N_11061,N_11039);
nand U11250 (N_11250,N_11051,N_11091);
and U11251 (N_11251,N_11155,N_11093);
or U11252 (N_11252,N_11047,N_11055);
and U11253 (N_11253,N_11169,N_11140);
and U11254 (N_11254,N_11121,N_11009);
nor U11255 (N_11255,N_11193,N_11179);
and U11256 (N_11256,N_11150,N_11086);
nor U11257 (N_11257,N_11182,N_11103);
nor U11258 (N_11258,N_11046,N_11040);
nand U11259 (N_11259,N_11012,N_11116);
nor U11260 (N_11260,N_11062,N_11180);
nor U11261 (N_11261,N_11158,N_11176);
and U11262 (N_11262,N_11013,N_11000);
nand U11263 (N_11263,N_11126,N_11127);
nor U11264 (N_11264,N_11107,N_11026);
or U11265 (N_11265,N_11077,N_11032);
nor U11266 (N_11266,N_11045,N_11197);
nor U11267 (N_11267,N_11041,N_11164);
and U11268 (N_11268,N_11053,N_11075);
nor U11269 (N_11269,N_11194,N_11161);
nand U11270 (N_11270,N_11184,N_11007);
nand U11271 (N_11271,N_11162,N_11163);
nand U11272 (N_11272,N_11064,N_11199);
or U11273 (N_11273,N_11190,N_11076);
and U11274 (N_11274,N_11188,N_11166);
nor U11275 (N_11275,N_11038,N_11145);
and U11276 (N_11276,N_11080,N_11186);
and U11277 (N_11277,N_11067,N_11124);
nor U11278 (N_11278,N_11020,N_11059);
nand U11279 (N_11279,N_11129,N_11183);
nor U11280 (N_11280,N_11092,N_11079);
nor U11281 (N_11281,N_11087,N_11120);
nand U11282 (N_11282,N_11165,N_11097);
nand U11283 (N_11283,N_11175,N_11112);
and U11284 (N_11284,N_11125,N_11142);
or U11285 (N_11285,N_11141,N_11171);
nor U11286 (N_11286,N_11005,N_11033);
and U11287 (N_11287,N_11173,N_11072);
and U11288 (N_11288,N_11042,N_11157);
and U11289 (N_11289,N_11008,N_11019);
or U11290 (N_11290,N_11132,N_11031);
or U11291 (N_11291,N_11104,N_11138);
and U11292 (N_11292,N_11014,N_11035);
nor U11293 (N_11293,N_11122,N_11085);
nand U11294 (N_11294,N_11106,N_11030);
nand U11295 (N_11295,N_11060,N_11084);
nand U11296 (N_11296,N_11115,N_11143);
xnor U11297 (N_11297,N_11113,N_11137);
nand U11298 (N_11298,N_11006,N_11189);
or U11299 (N_11299,N_11065,N_11070);
and U11300 (N_11300,N_11087,N_11159);
and U11301 (N_11301,N_11169,N_11047);
nand U11302 (N_11302,N_11056,N_11199);
or U11303 (N_11303,N_11090,N_11088);
or U11304 (N_11304,N_11120,N_11199);
or U11305 (N_11305,N_11196,N_11029);
xnor U11306 (N_11306,N_11154,N_11054);
or U11307 (N_11307,N_11097,N_11011);
and U11308 (N_11308,N_11018,N_11094);
nor U11309 (N_11309,N_11180,N_11075);
nand U11310 (N_11310,N_11130,N_11015);
nor U11311 (N_11311,N_11187,N_11184);
nand U11312 (N_11312,N_11026,N_11108);
nand U11313 (N_11313,N_11008,N_11011);
nor U11314 (N_11314,N_11102,N_11072);
and U11315 (N_11315,N_11046,N_11124);
and U11316 (N_11316,N_11020,N_11015);
and U11317 (N_11317,N_11190,N_11158);
nor U11318 (N_11318,N_11185,N_11153);
or U11319 (N_11319,N_11153,N_11090);
nand U11320 (N_11320,N_11122,N_11079);
nand U11321 (N_11321,N_11022,N_11143);
nor U11322 (N_11322,N_11006,N_11108);
or U11323 (N_11323,N_11165,N_11133);
nand U11324 (N_11324,N_11034,N_11147);
and U11325 (N_11325,N_11117,N_11037);
and U11326 (N_11326,N_11050,N_11144);
and U11327 (N_11327,N_11082,N_11135);
and U11328 (N_11328,N_11087,N_11071);
xnor U11329 (N_11329,N_11047,N_11180);
nor U11330 (N_11330,N_11174,N_11074);
or U11331 (N_11331,N_11156,N_11004);
and U11332 (N_11332,N_11061,N_11114);
and U11333 (N_11333,N_11171,N_11170);
nor U11334 (N_11334,N_11008,N_11179);
and U11335 (N_11335,N_11050,N_11038);
and U11336 (N_11336,N_11110,N_11036);
and U11337 (N_11337,N_11038,N_11183);
nor U11338 (N_11338,N_11046,N_11026);
or U11339 (N_11339,N_11137,N_11050);
nand U11340 (N_11340,N_11113,N_11154);
and U11341 (N_11341,N_11178,N_11174);
or U11342 (N_11342,N_11115,N_11027);
nand U11343 (N_11343,N_11148,N_11104);
and U11344 (N_11344,N_11009,N_11139);
and U11345 (N_11345,N_11051,N_11176);
nand U11346 (N_11346,N_11173,N_11164);
and U11347 (N_11347,N_11160,N_11186);
nand U11348 (N_11348,N_11089,N_11019);
and U11349 (N_11349,N_11018,N_11125);
nand U11350 (N_11350,N_11048,N_11031);
or U11351 (N_11351,N_11171,N_11043);
and U11352 (N_11352,N_11170,N_11004);
nand U11353 (N_11353,N_11069,N_11191);
or U11354 (N_11354,N_11186,N_11146);
nor U11355 (N_11355,N_11006,N_11149);
and U11356 (N_11356,N_11100,N_11158);
and U11357 (N_11357,N_11061,N_11081);
or U11358 (N_11358,N_11187,N_11054);
and U11359 (N_11359,N_11122,N_11167);
nand U11360 (N_11360,N_11122,N_11062);
or U11361 (N_11361,N_11079,N_11099);
nor U11362 (N_11362,N_11051,N_11026);
nand U11363 (N_11363,N_11118,N_11166);
nand U11364 (N_11364,N_11166,N_11124);
nor U11365 (N_11365,N_11098,N_11100);
nor U11366 (N_11366,N_11083,N_11018);
or U11367 (N_11367,N_11076,N_11160);
and U11368 (N_11368,N_11095,N_11043);
nor U11369 (N_11369,N_11003,N_11193);
and U11370 (N_11370,N_11056,N_11159);
nand U11371 (N_11371,N_11118,N_11044);
nand U11372 (N_11372,N_11192,N_11189);
nor U11373 (N_11373,N_11108,N_11111);
or U11374 (N_11374,N_11082,N_11168);
nor U11375 (N_11375,N_11055,N_11122);
nand U11376 (N_11376,N_11173,N_11129);
nor U11377 (N_11377,N_11151,N_11157);
and U11378 (N_11378,N_11177,N_11018);
or U11379 (N_11379,N_11054,N_11190);
and U11380 (N_11380,N_11066,N_11050);
nand U11381 (N_11381,N_11045,N_11141);
and U11382 (N_11382,N_11110,N_11082);
and U11383 (N_11383,N_11047,N_11044);
nand U11384 (N_11384,N_11138,N_11115);
nor U11385 (N_11385,N_11062,N_11112);
nor U11386 (N_11386,N_11101,N_11066);
or U11387 (N_11387,N_11164,N_11070);
nand U11388 (N_11388,N_11166,N_11127);
nor U11389 (N_11389,N_11012,N_11096);
and U11390 (N_11390,N_11138,N_11118);
nor U11391 (N_11391,N_11135,N_11010);
nand U11392 (N_11392,N_11103,N_11144);
nand U11393 (N_11393,N_11126,N_11196);
and U11394 (N_11394,N_11181,N_11078);
nor U11395 (N_11395,N_11167,N_11064);
or U11396 (N_11396,N_11153,N_11120);
or U11397 (N_11397,N_11164,N_11017);
and U11398 (N_11398,N_11078,N_11062);
or U11399 (N_11399,N_11100,N_11139);
nor U11400 (N_11400,N_11394,N_11364);
nand U11401 (N_11401,N_11244,N_11226);
or U11402 (N_11402,N_11238,N_11378);
xnor U11403 (N_11403,N_11269,N_11245);
nand U11404 (N_11404,N_11345,N_11361);
and U11405 (N_11405,N_11236,N_11205);
and U11406 (N_11406,N_11203,N_11386);
nand U11407 (N_11407,N_11330,N_11327);
nor U11408 (N_11408,N_11297,N_11301);
xor U11409 (N_11409,N_11232,N_11270);
or U11410 (N_11410,N_11304,N_11209);
and U11411 (N_11411,N_11337,N_11273);
and U11412 (N_11412,N_11279,N_11362);
nor U11413 (N_11413,N_11201,N_11287);
and U11414 (N_11414,N_11357,N_11384);
nor U11415 (N_11415,N_11370,N_11237);
and U11416 (N_11416,N_11217,N_11380);
xor U11417 (N_11417,N_11328,N_11289);
nand U11418 (N_11418,N_11381,N_11250);
nor U11419 (N_11419,N_11243,N_11341);
nand U11420 (N_11420,N_11314,N_11254);
nor U11421 (N_11421,N_11271,N_11216);
or U11422 (N_11422,N_11366,N_11343);
or U11423 (N_11423,N_11392,N_11240);
nor U11424 (N_11424,N_11223,N_11268);
and U11425 (N_11425,N_11204,N_11348);
nand U11426 (N_11426,N_11233,N_11280);
nand U11427 (N_11427,N_11372,N_11225);
and U11428 (N_11428,N_11339,N_11283);
nand U11429 (N_11429,N_11368,N_11340);
nand U11430 (N_11430,N_11231,N_11278);
and U11431 (N_11431,N_11334,N_11215);
nor U11432 (N_11432,N_11235,N_11256);
nor U11433 (N_11433,N_11376,N_11264);
and U11434 (N_11434,N_11352,N_11298);
xnor U11435 (N_11435,N_11285,N_11316);
nor U11436 (N_11436,N_11382,N_11311);
and U11437 (N_11437,N_11336,N_11275);
nor U11438 (N_11438,N_11212,N_11331);
nand U11439 (N_11439,N_11222,N_11211);
nor U11440 (N_11440,N_11207,N_11300);
xnor U11441 (N_11441,N_11208,N_11346);
and U11442 (N_11442,N_11385,N_11375);
nor U11443 (N_11443,N_11303,N_11379);
nand U11444 (N_11444,N_11306,N_11276);
or U11445 (N_11445,N_11224,N_11305);
nand U11446 (N_11446,N_11241,N_11326);
or U11447 (N_11447,N_11349,N_11324);
or U11448 (N_11448,N_11315,N_11296);
nand U11449 (N_11449,N_11329,N_11288);
xnor U11450 (N_11450,N_11277,N_11312);
and U11451 (N_11451,N_11387,N_11399);
nand U11452 (N_11452,N_11239,N_11246);
nor U11453 (N_11453,N_11320,N_11219);
or U11454 (N_11454,N_11318,N_11262);
nor U11455 (N_11455,N_11391,N_11388);
and U11456 (N_11456,N_11350,N_11309);
or U11457 (N_11457,N_11322,N_11397);
and U11458 (N_11458,N_11292,N_11286);
and U11459 (N_11459,N_11249,N_11367);
nand U11460 (N_11460,N_11265,N_11317);
nand U11461 (N_11461,N_11266,N_11354);
nand U11462 (N_11462,N_11206,N_11396);
and U11463 (N_11463,N_11313,N_11360);
nor U11464 (N_11464,N_11373,N_11323);
nand U11465 (N_11465,N_11247,N_11272);
or U11466 (N_11466,N_11351,N_11252);
or U11467 (N_11467,N_11259,N_11302);
nor U11468 (N_11468,N_11395,N_11325);
nand U11469 (N_11469,N_11200,N_11332);
or U11470 (N_11470,N_11213,N_11294);
nand U11471 (N_11471,N_11335,N_11261);
or U11472 (N_11472,N_11359,N_11202);
nor U11473 (N_11473,N_11338,N_11321);
nor U11474 (N_11474,N_11227,N_11347);
or U11475 (N_11475,N_11290,N_11358);
and U11476 (N_11476,N_11257,N_11398);
nand U11477 (N_11477,N_11295,N_11344);
and U11478 (N_11478,N_11234,N_11356);
xnor U11479 (N_11479,N_11218,N_11333);
nand U11480 (N_11480,N_11228,N_11374);
nand U11481 (N_11481,N_11282,N_11369);
and U11482 (N_11482,N_11260,N_11342);
xor U11483 (N_11483,N_11353,N_11293);
or U11484 (N_11484,N_11365,N_11221);
nand U11485 (N_11485,N_11310,N_11214);
or U11486 (N_11486,N_11230,N_11390);
and U11487 (N_11487,N_11393,N_11229);
and U11488 (N_11488,N_11377,N_11267);
xnor U11489 (N_11489,N_11371,N_11251);
and U11490 (N_11490,N_11210,N_11383);
and U11491 (N_11491,N_11242,N_11258);
nand U11492 (N_11492,N_11255,N_11307);
and U11493 (N_11493,N_11248,N_11389);
nor U11494 (N_11494,N_11220,N_11274);
or U11495 (N_11495,N_11355,N_11319);
and U11496 (N_11496,N_11281,N_11263);
or U11497 (N_11497,N_11363,N_11284);
and U11498 (N_11498,N_11308,N_11253);
nand U11499 (N_11499,N_11299,N_11291);
or U11500 (N_11500,N_11259,N_11294);
nand U11501 (N_11501,N_11347,N_11333);
or U11502 (N_11502,N_11321,N_11288);
or U11503 (N_11503,N_11268,N_11357);
nand U11504 (N_11504,N_11392,N_11397);
and U11505 (N_11505,N_11238,N_11357);
nor U11506 (N_11506,N_11215,N_11342);
nor U11507 (N_11507,N_11255,N_11342);
and U11508 (N_11508,N_11376,N_11204);
or U11509 (N_11509,N_11260,N_11213);
xnor U11510 (N_11510,N_11309,N_11315);
nor U11511 (N_11511,N_11348,N_11337);
and U11512 (N_11512,N_11322,N_11341);
nor U11513 (N_11513,N_11266,N_11353);
nand U11514 (N_11514,N_11207,N_11348);
and U11515 (N_11515,N_11303,N_11339);
and U11516 (N_11516,N_11297,N_11384);
and U11517 (N_11517,N_11242,N_11254);
nand U11518 (N_11518,N_11222,N_11359);
nand U11519 (N_11519,N_11241,N_11361);
and U11520 (N_11520,N_11379,N_11281);
nand U11521 (N_11521,N_11370,N_11263);
and U11522 (N_11522,N_11322,N_11248);
nor U11523 (N_11523,N_11354,N_11363);
nand U11524 (N_11524,N_11362,N_11226);
or U11525 (N_11525,N_11379,N_11296);
nor U11526 (N_11526,N_11298,N_11270);
and U11527 (N_11527,N_11248,N_11370);
nand U11528 (N_11528,N_11206,N_11366);
or U11529 (N_11529,N_11399,N_11220);
nor U11530 (N_11530,N_11371,N_11342);
nor U11531 (N_11531,N_11206,N_11324);
and U11532 (N_11532,N_11253,N_11239);
and U11533 (N_11533,N_11386,N_11248);
and U11534 (N_11534,N_11229,N_11334);
or U11535 (N_11535,N_11210,N_11251);
nor U11536 (N_11536,N_11216,N_11382);
nor U11537 (N_11537,N_11229,N_11220);
nand U11538 (N_11538,N_11292,N_11332);
nor U11539 (N_11539,N_11359,N_11271);
and U11540 (N_11540,N_11299,N_11356);
and U11541 (N_11541,N_11292,N_11326);
or U11542 (N_11542,N_11282,N_11328);
nand U11543 (N_11543,N_11212,N_11258);
nand U11544 (N_11544,N_11367,N_11250);
nor U11545 (N_11545,N_11335,N_11202);
and U11546 (N_11546,N_11294,N_11249);
nand U11547 (N_11547,N_11395,N_11291);
and U11548 (N_11548,N_11345,N_11299);
nand U11549 (N_11549,N_11329,N_11331);
nor U11550 (N_11550,N_11262,N_11325);
or U11551 (N_11551,N_11283,N_11327);
nor U11552 (N_11552,N_11355,N_11310);
or U11553 (N_11553,N_11266,N_11216);
or U11554 (N_11554,N_11293,N_11227);
nand U11555 (N_11555,N_11258,N_11356);
nand U11556 (N_11556,N_11283,N_11336);
or U11557 (N_11557,N_11287,N_11240);
and U11558 (N_11558,N_11330,N_11206);
or U11559 (N_11559,N_11347,N_11268);
and U11560 (N_11560,N_11337,N_11266);
nand U11561 (N_11561,N_11387,N_11375);
and U11562 (N_11562,N_11379,N_11364);
nor U11563 (N_11563,N_11352,N_11312);
nand U11564 (N_11564,N_11289,N_11217);
or U11565 (N_11565,N_11376,N_11200);
nor U11566 (N_11566,N_11372,N_11233);
nor U11567 (N_11567,N_11295,N_11362);
xor U11568 (N_11568,N_11321,N_11311);
nor U11569 (N_11569,N_11212,N_11240);
nor U11570 (N_11570,N_11282,N_11398);
nor U11571 (N_11571,N_11250,N_11200);
nor U11572 (N_11572,N_11215,N_11285);
and U11573 (N_11573,N_11251,N_11228);
or U11574 (N_11574,N_11206,N_11207);
and U11575 (N_11575,N_11238,N_11245);
or U11576 (N_11576,N_11237,N_11244);
nor U11577 (N_11577,N_11379,N_11338);
and U11578 (N_11578,N_11354,N_11383);
nor U11579 (N_11579,N_11270,N_11362);
nand U11580 (N_11580,N_11228,N_11282);
and U11581 (N_11581,N_11262,N_11338);
and U11582 (N_11582,N_11318,N_11331);
or U11583 (N_11583,N_11274,N_11200);
nand U11584 (N_11584,N_11382,N_11314);
and U11585 (N_11585,N_11391,N_11311);
xor U11586 (N_11586,N_11389,N_11285);
nor U11587 (N_11587,N_11314,N_11379);
nand U11588 (N_11588,N_11208,N_11315);
and U11589 (N_11589,N_11345,N_11396);
or U11590 (N_11590,N_11212,N_11383);
or U11591 (N_11591,N_11370,N_11231);
nor U11592 (N_11592,N_11233,N_11331);
and U11593 (N_11593,N_11214,N_11348);
or U11594 (N_11594,N_11209,N_11215);
nor U11595 (N_11595,N_11224,N_11203);
and U11596 (N_11596,N_11229,N_11216);
or U11597 (N_11597,N_11372,N_11312);
nand U11598 (N_11598,N_11386,N_11341);
nand U11599 (N_11599,N_11295,N_11261);
or U11600 (N_11600,N_11410,N_11409);
or U11601 (N_11601,N_11478,N_11578);
nand U11602 (N_11602,N_11564,N_11515);
nand U11603 (N_11603,N_11492,N_11594);
nand U11604 (N_11604,N_11416,N_11407);
nor U11605 (N_11605,N_11553,N_11475);
nand U11606 (N_11606,N_11504,N_11413);
nor U11607 (N_11607,N_11426,N_11435);
or U11608 (N_11608,N_11582,N_11574);
nand U11609 (N_11609,N_11599,N_11548);
nor U11610 (N_11610,N_11588,N_11489);
nand U11611 (N_11611,N_11495,N_11518);
or U11612 (N_11612,N_11436,N_11427);
and U11613 (N_11613,N_11437,N_11422);
or U11614 (N_11614,N_11482,N_11408);
and U11615 (N_11615,N_11540,N_11572);
nand U11616 (N_11616,N_11406,N_11464);
nand U11617 (N_11617,N_11595,N_11520);
and U11618 (N_11618,N_11587,N_11526);
nor U11619 (N_11619,N_11531,N_11494);
xnor U11620 (N_11620,N_11499,N_11506);
nor U11621 (N_11621,N_11431,N_11425);
nand U11622 (N_11622,N_11516,N_11446);
nand U11623 (N_11623,N_11598,N_11454);
or U11624 (N_11624,N_11428,N_11501);
and U11625 (N_11625,N_11462,N_11539);
nand U11626 (N_11626,N_11581,N_11415);
or U11627 (N_11627,N_11488,N_11584);
and U11628 (N_11628,N_11483,N_11403);
or U11629 (N_11629,N_11476,N_11512);
and U11630 (N_11630,N_11498,N_11565);
or U11631 (N_11631,N_11468,N_11466);
and U11632 (N_11632,N_11541,N_11493);
nor U11633 (N_11633,N_11438,N_11457);
or U11634 (N_11634,N_11513,N_11434);
or U11635 (N_11635,N_11502,N_11561);
or U11636 (N_11636,N_11538,N_11592);
or U11637 (N_11637,N_11485,N_11442);
or U11638 (N_11638,N_11544,N_11568);
or U11639 (N_11639,N_11432,N_11429);
or U11640 (N_11640,N_11577,N_11452);
and U11641 (N_11641,N_11490,N_11535);
and U11642 (N_11642,N_11563,N_11536);
and U11643 (N_11643,N_11511,N_11491);
or U11644 (N_11644,N_11527,N_11573);
and U11645 (N_11645,N_11579,N_11591);
nand U11646 (N_11646,N_11473,N_11542);
and U11647 (N_11647,N_11439,N_11585);
nand U11648 (N_11648,N_11401,N_11424);
xor U11649 (N_11649,N_11554,N_11400);
xor U11650 (N_11650,N_11458,N_11414);
and U11651 (N_11651,N_11529,N_11461);
nand U11652 (N_11652,N_11550,N_11508);
nand U11653 (N_11653,N_11433,N_11430);
or U11654 (N_11654,N_11593,N_11509);
or U11655 (N_11655,N_11590,N_11525);
or U11656 (N_11656,N_11523,N_11423);
and U11657 (N_11657,N_11552,N_11459);
or U11658 (N_11658,N_11505,N_11580);
or U11659 (N_11659,N_11558,N_11596);
and U11660 (N_11660,N_11421,N_11445);
nor U11661 (N_11661,N_11521,N_11453);
nor U11662 (N_11662,N_11532,N_11465);
nand U11663 (N_11663,N_11405,N_11460);
nor U11664 (N_11664,N_11545,N_11524);
nor U11665 (N_11665,N_11551,N_11507);
nand U11666 (N_11666,N_11455,N_11597);
nand U11667 (N_11667,N_11444,N_11575);
nor U11668 (N_11668,N_11522,N_11583);
or U11669 (N_11669,N_11569,N_11474);
nor U11670 (N_11670,N_11497,N_11486);
nor U11671 (N_11671,N_11419,N_11471);
nand U11672 (N_11672,N_11449,N_11571);
nand U11673 (N_11673,N_11472,N_11543);
nand U11674 (N_11674,N_11441,N_11562);
nand U11675 (N_11675,N_11510,N_11557);
nand U11676 (N_11676,N_11567,N_11469);
or U11677 (N_11677,N_11576,N_11418);
nand U11678 (N_11678,N_11479,N_11547);
nand U11679 (N_11679,N_11412,N_11484);
and U11680 (N_11680,N_11559,N_11530);
nor U11681 (N_11681,N_11519,N_11411);
or U11682 (N_11682,N_11500,N_11451);
or U11683 (N_11683,N_11496,N_11487);
or U11684 (N_11684,N_11443,N_11586);
or U11685 (N_11685,N_11549,N_11456);
and U11686 (N_11686,N_11534,N_11514);
nor U11687 (N_11687,N_11555,N_11440);
nor U11688 (N_11688,N_11570,N_11533);
or U11689 (N_11689,N_11589,N_11528);
and U11690 (N_11690,N_11481,N_11560);
or U11691 (N_11691,N_11467,N_11447);
nand U11692 (N_11692,N_11556,N_11402);
nand U11693 (N_11693,N_11450,N_11537);
nand U11694 (N_11694,N_11404,N_11420);
nand U11695 (N_11695,N_11480,N_11470);
and U11696 (N_11696,N_11448,N_11566);
nor U11697 (N_11697,N_11477,N_11417);
nor U11698 (N_11698,N_11546,N_11517);
nand U11699 (N_11699,N_11463,N_11503);
and U11700 (N_11700,N_11410,N_11448);
nand U11701 (N_11701,N_11530,N_11429);
nor U11702 (N_11702,N_11436,N_11457);
nand U11703 (N_11703,N_11571,N_11543);
and U11704 (N_11704,N_11560,N_11569);
nand U11705 (N_11705,N_11451,N_11406);
and U11706 (N_11706,N_11549,N_11545);
nor U11707 (N_11707,N_11423,N_11413);
and U11708 (N_11708,N_11416,N_11569);
and U11709 (N_11709,N_11544,N_11528);
nand U11710 (N_11710,N_11452,N_11549);
and U11711 (N_11711,N_11559,N_11465);
or U11712 (N_11712,N_11499,N_11579);
nor U11713 (N_11713,N_11497,N_11580);
or U11714 (N_11714,N_11589,N_11532);
nand U11715 (N_11715,N_11443,N_11546);
or U11716 (N_11716,N_11466,N_11406);
nand U11717 (N_11717,N_11510,N_11489);
nor U11718 (N_11718,N_11478,N_11404);
nor U11719 (N_11719,N_11520,N_11503);
or U11720 (N_11720,N_11435,N_11516);
nand U11721 (N_11721,N_11577,N_11424);
and U11722 (N_11722,N_11475,N_11596);
nor U11723 (N_11723,N_11429,N_11502);
or U11724 (N_11724,N_11527,N_11538);
nor U11725 (N_11725,N_11552,N_11584);
and U11726 (N_11726,N_11518,N_11550);
and U11727 (N_11727,N_11450,N_11463);
xor U11728 (N_11728,N_11500,N_11460);
nor U11729 (N_11729,N_11581,N_11597);
nand U11730 (N_11730,N_11553,N_11545);
nor U11731 (N_11731,N_11414,N_11531);
nand U11732 (N_11732,N_11466,N_11599);
and U11733 (N_11733,N_11415,N_11426);
nor U11734 (N_11734,N_11452,N_11415);
or U11735 (N_11735,N_11505,N_11592);
and U11736 (N_11736,N_11594,N_11505);
nor U11737 (N_11737,N_11483,N_11435);
and U11738 (N_11738,N_11599,N_11544);
nor U11739 (N_11739,N_11539,N_11541);
nor U11740 (N_11740,N_11534,N_11403);
nor U11741 (N_11741,N_11432,N_11520);
nand U11742 (N_11742,N_11576,N_11433);
nand U11743 (N_11743,N_11571,N_11477);
nand U11744 (N_11744,N_11560,N_11532);
nand U11745 (N_11745,N_11512,N_11524);
nand U11746 (N_11746,N_11481,N_11583);
and U11747 (N_11747,N_11597,N_11438);
nand U11748 (N_11748,N_11571,N_11509);
nor U11749 (N_11749,N_11452,N_11514);
xnor U11750 (N_11750,N_11540,N_11441);
nor U11751 (N_11751,N_11440,N_11439);
nand U11752 (N_11752,N_11513,N_11556);
nor U11753 (N_11753,N_11519,N_11479);
nor U11754 (N_11754,N_11567,N_11591);
or U11755 (N_11755,N_11418,N_11580);
or U11756 (N_11756,N_11426,N_11555);
or U11757 (N_11757,N_11592,N_11486);
nor U11758 (N_11758,N_11513,N_11462);
or U11759 (N_11759,N_11547,N_11543);
nand U11760 (N_11760,N_11441,N_11555);
and U11761 (N_11761,N_11531,N_11526);
nor U11762 (N_11762,N_11464,N_11484);
xor U11763 (N_11763,N_11559,N_11501);
or U11764 (N_11764,N_11521,N_11444);
nand U11765 (N_11765,N_11496,N_11555);
nor U11766 (N_11766,N_11591,N_11459);
or U11767 (N_11767,N_11539,N_11456);
nand U11768 (N_11768,N_11532,N_11500);
nand U11769 (N_11769,N_11515,N_11418);
nand U11770 (N_11770,N_11449,N_11568);
or U11771 (N_11771,N_11555,N_11442);
or U11772 (N_11772,N_11536,N_11525);
nand U11773 (N_11773,N_11561,N_11441);
nand U11774 (N_11774,N_11549,N_11537);
and U11775 (N_11775,N_11444,N_11579);
or U11776 (N_11776,N_11459,N_11465);
and U11777 (N_11777,N_11581,N_11506);
nor U11778 (N_11778,N_11591,N_11448);
nor U11779 (N_11779,N_11577,N_11544);
nor U11780 (N_11780,N_11571,N_11496);
nor U11781 (N_11781,N_11552,N_11546);
and U11782 (N_11782,N_11503,N_11401);
nand U11783 (N_11783,N_11589,N_11457);
nand U11784 (N_11784,N_11584,N_11412);
nand U11785 (N_11785,N_11530,N_11458);
nor U11786 (N_11786,N_11409,N_11525);
and U11787 (N_11787,N_11419,N_11538);
and U11788 (N_11788,N_11506,N_11504);
nor U11789 (N_11789,N_11585,N_11557);
or U11790 (N_11790,N_11536,N_11598);
and U11791 (N_11791,N_11513,N_11514);
nor U11792 (N_11792,N_11401,N_11460);
and U11793 (N_11793,N_11461,N_11580);
and U11794 (N_11794,N_11545,N_11422);
and U11795 (N_11795,N_11438,N_11408);
and U11796 (N_11796,N_11437,N_11523);
or U11797 (N_11797,N_11550,N_11459);
nor U11798 (N_11798,N_11591,N_11593);
nor U11799 (N_11799,N_11567,N_11433);
and U11800 (N_11800,N_11632,N_11606);
and U11801 (N_11801,N_11681,N_11628);
nand U11802 (N_11802,N_11702,N_11789);
and U11803 (N_11803,N_11629,N_11786);
or U11804 (N_11804,N_11647,N_11735);
nor U11805 (N_11805,N_11761,N_11602);
or U11806 (N_11806,N_11694,N_11620);
nand U11807 (N_11807,N_11668,N_11773);
and U11808 (N_11808,N_11762,N_11784);
nand U11809 (N_11809,N_11642,N_11715);
nor U11810 (N_11810,N_11664,N_11776);
nand U11811 (N_11811,N_11621,N_11712);
or U11812 (N_11812,N_11680,N_11682);
nor U11813 (N_11813,N_11779,N_11722);
and U11814 (N_11814,N_11794,N_11635);
and U11815 (N_11815,N_11766,N_11692);
nor U11816 (N_11816,N_11725,N_11674);
or U11817 (N_11817,N_11676,N_11609);
nand U11818 (N_11818,N_11751,N_11723);
nand U11819 (N_11819,N_11615,N_11636);
nor U11820 (N_11820,N_11749,N_11790);
nor U11821 (N_11821,N_11679,N_11771);
nor U11822 (N_11822,N_11795,N_11600);
nor U11823 (N_11823,N_11740,N_11660);
or U11824 (N_11824,N_11696,N_11703);
nor U11825 (N_11825,N_11764,N_11732);
and U11826 (N_11826,N_11788,N_11768);
or U11827 (N_11827,N_11633,N_11758);
or U11828 (N_11828,N_11730,N_11737);
nor U11829 (N_11829,N_11719,N_11688);
nor U11830 (N_11830,N_11641,N_11724);
nand U11831 (N_11831,N_11665,N_11753);
nand U11832 (N_11832,N_11663,N_11698);
and U11833 (N_11833,N_11716,N_11704);
nand U11834 (N_11834,N_11695,N_11608);
nor U11835 (N_11835,N_11685,N_11765);
nand U11836 (N_11836,N_11626,N_11739);
and U11837 (N_11837,N_11657,N_11745);
and U11838 (N_11838,N_11605,N_11623);
nand U11839 (N_11839,N_11700,N_11710);
and U11840 (N_11840,N_11783,N_11697);
nand U11841 (N_11841,N_11713,N_11701);
nor U11842 (N_11842,N_11686,N_11752);
or U11843 (N_11843,N_11661,N_11782);
and U11844 (N_11844,N_11747,N_11742);
or U11845 (N_11845,N_11616,N_11666);
nor U11846 (N_11846,N_11670,N_11748);
and U11847 (N_11847,N_11727,N_11675);
xnor U11848 (N_11848,N_11733,N_11774);
or U11849 (N_11849,N_11690,N_11678);
nand U11850 (N_11850,N_11652,N_11651);
nand U11851 (N_11851,N_11770,N_11691);
and U11852 (N_11852,N_11653,N_11622);
xnor U11853 (N_11853,N_11687,N_11777);
and U11854 (N_11854,N_11655,N_11799);
nor U11855 (N_11855,N_11650,N_11643);
nand U11856 (N_11856,N_11763,N_11717);
or U11857 (N_11857,N_11729,N_11707);
or U11858 (N_11858,N_11718,N_11772);
or U11859 (N_11859,N_11736,N_11614);
and U11860 (N_11860,N_11767,N_11798);
nand U11861 (N_11861,N_11607,N_11611);
nor U11862 (N_11862,N_11793,N_11734);
nand U11863 (N_11863,N_11673,N_11797);
nor U11864 (N_11864,N_11638,N_11644);
nand U11865 (N_11865,N_11744,N_11640);
nand U11866 (N_11866,N_11778,N_11754);
nor U11867 (N_11867,N_11603,N_11769);
nand U11868 (N_11868,N_11741,N_11617);
nand U11869 (N_11869,N_11684,N_11711);
nand U11870 (N_11870,N_11667,N_11625);
nand U11871 (N_11871,N_11728,N_11659);
nor U11872 (N_11872,N_11731,N_11743);
or U11873 (N_11873,N_11683,N_11662);
nand U11874 (N_11874,N_11760,N_11671);
nand U11875 (N_11875,N_11645,N_11709);
nor U11876 (N_11876,N_11738,N_11601);
or U11877 (N_11877,N_11726,N_11780);
and U11878 (N_11878,N_11634,N_11677);
or U11879 (N_11879,N_11759,N_11619);
nand U11880 (N_11880,N_11746,N_11699);
or U11881 (N_11881,N_11649,N_11791);
or U11882 (N_11882,N_11613,N_11631);
nand U11883 (N_11883,N_11787,N_11750);
and U11884 (N_11884,N_11669,N_11756);
nor U11885 (N_11885,N_11720,N_11672);
or U11886 (N_11886,N_11714,N_11624);
or U11887 (N_11887,N_11755,N_11721);
nor U11888 (N_11888,N_11693,N_11705);
and U11889 (N_11889,N_11757,N_11630);
nand U11890 (N_11890,N_11775,N_11781);
nand U11891 (N_11891,N_11658,N_11646);
and U11892 (N_11892,N_11656,N_11796);
nand U11893 (N_11893,N_11612,N_11648);
or U11894 (N_11894,N_11708,N_11792);
nor U11895 (N_11895,N_11637,N_11610);
and U11896 (N_11896,N_11785,N_11654);
nand U11897 (N_11897,N_11618,N_11706);
nand U11898 (N_11898,N_11639,N_11627);
nor U11899 (N_11899,N_11689,N_11604);
nor U11900 (N_11900,N_11772,N_11770);
and U11901 (N_11901,N_11612,N_11733);
and U11902 (N_11902,N_11680,N_11705);
xnor U11903 (N_11903,N_11626,N_11701);
nor U11904 (N_11904,N_11777,N_11662);
or U11905 (N_11905,N_11678,N_11682);
and U11906 (N_11906,N_11775,N_11632);
nand U11907 (N_11907,N_11681,N_11633);
or U11908 (N_11908,N_11724,N_11779);
and U11909 (N_11909,N_11702,N_11766);
nand U11910 (N_11910,N_11785,N_11740);
and U11911 (N_11911,N_11632,N_11609);
or U11912 (N_11912,N_11602,N_11688);
nor U11913 (N_11913,N_11662,N_11725);
or U11914 (N_11914,N_11744,N_11684);
xor U11915 (N_11915,N_11622,N_11657);
and U11916 (N_11916,N_11684,N_11758);
nor U11917 (N_11917,N_11678,N_11696);
nand U11918 (N_11918,N_11658,N_11794);
nand U11919 (N_11919,N_11791,N_11644);
nand U11920 (N_11920,N_11782,N_11773);
nor U11921 (N_11921,N_11727,N_11687);
and U11922 (N_11922,N_11678,N_11611);
and U11923 (N_11923,N_11782,N_11697);
nor U11924 (N_11924,N_11788,N_11639);
or U11925 (N_11925,N_11773,N_11793);
nand U11926 (N_11926,N_11672,N_11766);
and U11927 (N_11927,N_11775,N_11751);
nand U11928 (N_11928,N_11675,N_11629);
nand U11929 (N_11929,N_11777,N_11789);
or U11930 (N_11930,N_11628,N_11617);
nor U11931 (N_11931,N_11721,N_11626);
nand U11932 (N_11932,N_11715,N_11732);
nor U11933 (N_11933,N_11742,N_11682);
nor U11934 (N_11934,N_11708,N_11625);
nand U11935 (N_11935,N_11640,N_11754);
or U11936 (N_11936,N_11667,N_11638);
and U11937 (N_11937,N_11705,N_11683);
and U11938 (N_11938,N_11766,N_11612);
nor U11939 (N_11939,N_11666,N_11694);
or U11940 (N_11940,N_11661,N_11692);
nor U11941 (N_11941,N_11641,N_11620);
nand U11942 (N_11942,N_11621,N_11695);
or U11943 (N_11943,N_11656,N_11610);
xor U11944 (N_11944,N_11770,N_11769);
nor U11945 (N_11945,N_11601,N_11708);
or U11946 (N_11946,N_11615,N_11629);
nor U11947 (N_11947,N_11743,N_11636);
and U11948 (N_11948,N_11701,N_11747);
or U11949 (N_11949,N_11649,N_11795);
or U11950 (N_11950,N_11710,N_11645);
and U11951 (N_11951,N_11600,N_11759);
and U11952 (N_11952,N_11724,N_11695);
nand U11953 (N_11953,N_11746,N_11720);
nor U11954 (N_11954,N_11627,N_11633);
xor U11955 (N_11955,N_11739,N_11731);
nor U11956 (N_11956,N_11617,N_11738);
nor U11957 (N_11957,N_11662,N_11796);
nor U11958 (N_11958,N_11753,N_11666);
nor U11959 (N_11959,N_11695,N_11728);
nor U11960 (N_11960,N_11789,N_11697);
nand U11961 (N_11961,N_11648,N_11664);
and U11962 (N_11962,N_11737,N_11675);
and U11963 (N_11963,N_11669,N_11737);
and U11964 (N_11964,N_11615,N_11739);
nand U11965 (N_11965,N_11610,N_11717);
and U11966 (N_11966,N_11656,N_11659);
nor U11967 (N_11967,N_11765,N_11721);
nand U11968 (N_11968,N_11743,N_11711);
nor U11969 (N_11969,N_11700,N_11602);
or U11970 (N_11970,N_11610,N_11720);
and U11971 (N_11971,N_11641,N_11631);
xor U11972 (N_11972,N_11791,N_11684);
nand U11973 (N_11973,N_11709,N_11661);
and U11974 (N_11974,N_11680,N_11789);
or U11975 (N_11975,N_11667,N_11629);
nor U11976 (N_11976,N_11788,N_11628);
or U11977 (N_11977,N_11749,N_11748);
nand U11978 (N_11978,N_11750,N_11664);
and U11979 (N_11979,N_11720,N_11668);
or U11980 (N_11980,N_11654,N_11746);
and U11981 (N_11981,N_11652,N_11621);
nand U11982 (N_11982,N_11717,N_11680);
and U11983 (N_11983,N_11752,N_11622);
nand U11984 (N_11984,N_11645,N_11707);
xor U11985 (N_11985,N_11681,N_11720);
nand U11986 (N_11986,N_11752,N_11660);
nand U11987 (N_11987,N_11694,N_11722);
or U11988 (N_11988,N_11714,N_11782);
or U11989 (N_11989,N_11784,N_11606);
nor U11990 (N_11990,N_11758,N_11625);
and U11991 (N_11991,N_11600,N_11651);
and U11992 (N_11992,N_11710,N_11626);
nand U11993 (N_11993,N_11655,N_11729);
or U11994 (N_11994,N_11643,N_11668);
nand U11995 (N_11995,N_11745,N_11721);
nand U11996 (N_11996,N_11767,N_11719);
and U11997 (N_11997,N_11748,N_11706);
nor U11998 (N_11998,N_11746,N_11759);
or U11999 (N_11999,N_11694,N_11775);
or U12000 (N_12000,N_11911,N_11896);
and U12001 (N_12001,N_11860,N_11925);
nor U12002 (N_12002,N_11976,N_11894);
and U12003 (N_12003,N_11995,N_11877);
nor U12004 (N_12004,N_11891,N_11930);
nand U12005 (N_12005,N_11868,N_11953);
or U12006 (N_12006,N_11839,N_11916);
or U12007 (N_12007,N_11936,N_11947);
nand U12008 (N_12008,N_11988,N_11935);
nand U12009 (N_12009,N_11990,N_11972);
or U12010 (N_12010,N_11840,N_11897);
or U12011 (N_12011,N_11899,N_11890);
or U12012 (N_12012,N_11823,N_11801);
nand U12013 (N_12013,N_11973,N_11974);
or U12014 (N_12014,N_11817,N_11985);
or U12015 (N_12015,N_11956,N_11810);
nor U12016 (N_12016,N_11922,N_11955);
nand U12017 (N_12017,N_11999,N_11884);
nor U12018 (N_12018,N_11993,N_11926);
and U12019 (N_12019,N_11834,N_11883);
nor U12020 (N_12020,N_11886,N_11832);
or U12021 (N_12021,N_11917,N_11881);
or U12022 (N_12022,N_11994,N_11895);
and U12023 (N_12023,N_11984,N_11914);
and U12024 (N_12024,N_11904,N_11830);
nor U12025 (N_12025,N_11918,N_11991);
or U12026 (N_12026,N_11966,N_11802);
and U12027 (N_12027,N_11844,N_11932);
and U12028 (N_12028,N_11861,N_11855);
nand U12029 (N_12029,N_11815,N_11989);
nor U12030 (N_12030,N_11863,N_11825);
nand U12031 (N_12031,N_11983,N_11927);
or U12032 (N_12032,N_11905,N_11892);
nor U12033 (N_12033,N_11843,N_11921);
and U12034 (N_12034,N_11900,N_11866);
nor U12035 (N_12035,N_11813,N_11951);
xnor U12036 (N_12036,N_11806,N_11913);
nand U12037 (N_12037,N_11933,N_11814);
xor U12038 (N_12038,N_11804,N_11871);
or U12039 (N_12039,N_11878,N_11963);
or U12040 (N_12040,N_11812,N_11893);
or U12041 (N_12041,N_11977,N_11996);
and U12042 (N_12042,N_11885,N_11836);
nor U12043 (N_12043,N_11950,N_11987);
nand U12044 (N_12044,N_11888,N_11934);
and U12045 (N_12045,N_11901,N_11828);
nor U12046 (N_12046,N_11858,N_11915);
or U12047 (N_12047,N_11827,N_11969);
nand U12048 (N_12048,N_11962,N_11821);
and U12049 (N_12049,N_11873,N_11939);
and U12050 (N_12050,N_11808,N_11941);
and U12051 (N_12051,N_11853,N_11946);
nand U12052 (N_12052,N_11997,N_11923);
or U12053 (N_12053,N_11929,N_11875);
nor U12054 (N_12054,N_11979,N_11937);
and U12055 (N_12055,N_11906,N_11902);
nand U12056 (N_12056,N_11924,N_11903);
or U12057 (N_12057,N_11960,N_11958);
and U12058 (N_12058,N_11852,N_11998);
or U12059 (N_12059,N_11954,N_11818);
nand U12060 (N_12060,N_11908,N_11944);
nor U12061 (N_12061,N_11835,N_11838);
and U12062 (N_12062,N_11942,N_11851);
nor U12063 (N_12063,N_11874,N_11952);
or U12064 (N_12064,N_11879,N_11909);
or U12065 (N_12065,N_11826,N_11945);
nand U12066 (N_12066,N_11880,N_11889);
nor U12067 (N_12067,N_11845,N_11982);
nor U12068 (N_12068,N_11876,N_11943);
nor U12069 (N_12069,N_11959,N_11833);
or U12070 (N_12070,N_11846,N_11992);
nand U12071 (N_12071,N_11811,N_11865);
or U12072 (N_12072,N_11847,N_11967);
nand U12073 (N_12073,N_11986,N_11803);
and U12074 (N_12074,N_11820,N_11870);
and U12075 (N_12075,N_11822,N_11824);
nor U12076 (N_12076,N_11809,N_11961);
nand U12077 (N_12077,N_11978,N_11949);
nand U12078 (N_12078,N_11867,N_11842);
or U12079 (N_12079,N_11940,N_11862);
nand U12080 (N_12080,N_11857,N_11864);
and U12081 (N_12081,N_11859,N_11850);
nand U12082 (N_12082,N_11869,N_11841);
or U12083 (N_12083,N_11829,N_11912);
nand U12084 (N_12084,N_11965,N_11848);
nand U12085 (N_12085,N_11964,N_11854);
nor U12086 (N_12086,N_11980,N_11910);
nand U12087 (N_12087,N_11948,N_11928);
nand U12088 (N_12088,N_11931,N_11968);
nand U12089 (N_12089,N_11816,N_11856);
or U12090 (N_12090,N_11898,N_11887);
nor U12091 (N_12091,N_11819,N_11920);
nor U12092 (N_12092,N_11981,N_11919);
nor U12093 (N_12093,N_11837,N_11831);
nor U12094 (N_12094,N_11882,N_11907);
nand U12095 (N_12095,N_11807,N_11970);
and U12096 (N_12096,N_11938,N_11805);
nor U12097 (N_12097,N_11957,N_11975);
nor U12098 (N_12098,N_11872,N_11849);
nor U12099 (N_12099,N_11971,N_11800);
or U12100 (N_12100,N_11853,N_11969);
nand U12101 (N_12101,N_11837,N_11838);
and U12102 (N_12102,N_11979,N_11950);
xor U12103 (N_12103,N_11840,N_11827);
xnor U12104 (N_12104,N_11938,N_11959);
nand U12105 (N_12105,N_11879,N_11924);
nand U12106 (N_12106,N_11950,N_11996);
nor U12107 (N_12107,N_11852,N_11967);
nor U12108 (N_12108,N_11912,N_11979);
nor U12109 (N_12109,N_11840,N_11839);
or U12110 (N_12110,N_11895,N_11991);
nor U12111 (N_12111,N_11904,N_11999);
nand U12112 (N_12112,N_11994,N_11968);
nand U12113 (N_12113,N_11940,N_11854);
and U12114 (N_12114,N_11936,N_11939);
nor U12115 (N_12115,N_11969,N_11808);
or U12116 (N_12116,N_11849,N_11800);
nand U12117 (N_12117,N_11982,N_11936);
nand U12118 (N_12118,N_11977,N_11803);
nand U12119 (N_12119,N_11992,N_11852);
nand U12120 (N_12120,N_11931,N_11959);
nand U12121 (N_12121,N_11947,N_11835);
nor U12122 (N_12122,N_11828,N_11803);
nand U12123 (N_12123,N_11936,N_11930);
or U12124 (N_12124,N_11846,N_11955);
and U12125 (N_12125,N_11997,N_11960);
and U12126 (N_12126,N_11986,N_11934);
and U12127 (N_12127,N_11956,N_11828);
nand U12128 (N_12128,N_11929,N_11833);
nand U12129 (N_12129,N_11980,N_11895);
and U12130 (N_12130,N_11879,N_11870);
and U12131 (N_12131,N_11905,N_11937);
and U12132 (N_12132,N_11858,N_11814);
or U12133 (N_12133,N_11931,N_11906);
nor U12134 (N_12134,N_11992,N_11864);
or U12135 (N_12135,N_11817,N_11978);
and U12136 (N_12136,N_11880,N_11954);
or U12137 (N_12137,N_11965,N_11925);
nand U12138 (N_12138,N_11986,N_11951);
nand U12139 (N_12139,N_11893,N_11965);
nand U12140 (N_12140,N_11843,N_11876);
and U12141 (N_12141,N_11868,N_11843);
and U12142 (N_12142,N_11841,N_11837);
nor U12143 (N_12143,N_11835,N_11828);
or U12144 (N_12144,N_11962,N_11896);
nor U12145 (N_12145,N_11814,N_11915);
or U12146 (N_12146,N_11996,N_11921);
nor U12147 (N_12147,N_11807,N_11809);
nor U12148 (N_12148,N_11985,N_11886);
or U12149 (N_12149,N_11801,N_11868);
nor U12150 (N_12150,N_11801,N_11892);
and U12151 (N_12151,N_11814,N_11803);
nor U12152 (N_12152,N_11933,N_11867);
xor U12153 (N_12153,N_11987,N_11802);
or U12154 (N_12154,N_11802,N_11827);
or U12155 (N_12155,N_11931,N_11812);
or U12156 (N_12156,N_11896,N_11816);
or U12157 (N_12157,N_11999,N_11816);
nor U12158 (N_12158,N_11843,N_11963);
nand U12159 (N_12159,N_11903,N_11868);
nand U12160 (N_12160,N_11837,N_11803);
nand U12161 (N_12161,N_11912,N_11880);
nor U12162 (N_12162,N_11933,N_11835);
nor U12163 (N_12163,N_11897,N_11858);
nand U12164 (N_12164,N_11891,N_11815);
and U12165 (N_12165,N_11809,N_11815);
or U12166 (N_12166,N_11956,N_11875);
nor U12167 (N_12167,N_11915,N_11880);
xnor U12168 (N_12168,N_11972,N_11870);
and U12169 (N_12169,N_11917,N_11800);
and U12170 (N_12170,N_11913,N_11937);
nand U12171 (N_12171,N_11965,N_11975);
and U12172 (N_12172,N_11912,N_11864);
nor U12173 (N_12173,N_11816,N_11961);
nor U12174 (N_12174,N_11938,N_11977);
nor U12175 (N_12175,N_11811,N_11861);
and U12176 (N_12176,N_11804,N_11849);
or U12177 (N_12177,N_11901,N_11887);
and U12178 (N_12178,N_11807,N_11839);
and U12179 (N_12179,N_11969,N_11914);
and U12180 (N_12180,N_11951,N_11988);
nand U12181 (N_12181,N_11838,N_11926);
nor U12182 (N_12182,N_11924,N_11834);
nand U12183 (N_12183,N_11814,N_11821);
nor U12184 (N_12184,N_11980,N_11997);
or U12185 (N_12185,N_11885,N_11908);
or U12186 (N_12186,N_11982,N_11963);
and U12187 (N_12187,N_11831,N_11893);
or U12188 (N_12188,N_11877,N_11952);
nor U12189 (N_12189,N_11831,N_11830);
nand U12190 (N_12190,N_11867,N_11918);
and U12191 (N_12191,N_11919,N_11922);
or U12192 (N_12192,N_11817,N_11811);
nor U12193 (N_12193,N_11880,N_11846);
or U12194 (N_12194,N_11839,N_11854);
and U12195 (N_12195,N_11897,N_11871);
nor U12196 (N_12196,N_11977,N_11918);
or U12197 (N_12197,N_11847,N_11950);
nor U12198 (N_12198,N_11849,N_11850);
nor U12199 (N_12199,N_11826,N_11845);
and U12200 (N_12200,N_12090,N_12178);
nor U12201 (N_12201,N_12038,N_12144);
and U12202 (N_12202,N_12083,N_12124);
nor U12203 (N_12203,N_12074,N_12011);
or U12204 (N_12204,N_12128,N_12168);
and U12205 (N_12205,N_12098,N_12116);
nor U12206 (N_12206,N_12158,N_12054);
or U12207 (N_12207,N_12176,N_12031);
or U12208 (N_12208,N_12005,N_12096);
nor U12209 (N_12209,N_12131,N_12133);
nor U12210 (N_12210,N_12161,N_12013);
nor U12211 (N_12211,N_12071,N_12028);
or U12212 (N_12212,N_12137,N_12026);
and U12213 (N_12213,N_12153,N_12012);
or U12214 (N_12214,N_12094,N_12162);
and U12215 (N_12215,N_12042,N_12119);
nand U12216 (N_12216,N_12066,N_12198);
or U12217 (N_12217,N_12166,N_12065);
and U12218 (N_12218,N_12047,N_12018);
nor U12219 (N_12219,N_12089,N_12076);
nor U12220 (N_12220,N_12022,N_12113);
or U12221 (N_12221,N_12095,N_12175);
or U12222 (N_12222,N_12165,N_12025);
and U12223 (N_12223,N_12114,N_12030);
nor U12224 (N_12224,N_12062,N_12040);
nand U12225 (N_12225,N_12058,N_12180);
and U12226 (N_12226,N_12155,N_12021);
or U12227 (N_12227,N_12129,N_12057);
or U12228 (N_12228,N_12015,N_12164);
nand U12229 (N_12229,N_12147,N_12055);
and U12230 (N_12230,N_12050,N_12100);
nand U12231 (N_12231,N_12108,N_12138);
or U12232 (N_12232,N_12014,N_12084);
and U12233 (N_12233,N_12097,N_12061);
nand U12234 (N_12234,N_12056,N_12009);
or U12235 (N_12235,N_12002,N_12063);
or U12236 (N_12236,N_12051,N_12069);
and U12237 (N_12237,N_12188,N_12148);
nor U12238 (N_12238,N_12035,N_12078);
nand U12239 (N_12239,N_12199,N_12064);
or U12240 (N_12240,N_12104,N_12060);
and U12241 (N_12241,N_12163,N_12023);
or U12242 (N_12242,N_12016,N_12157);
and U12243 (N_12243,N_12192,N_12115);
and U12244 (N_12244,N_12149,N_12187);
nand U12245 (N_12245,N_12196,N_12190);
nand U12246 (N_12246,N_12156,N_12173);
nor U12247 (N_12247,N_12130,N_12117);
or U12248 (N_12248,N_12109,N_12032);
nor U12249 (N_12249,N_12179,N_12172);
and U12250 (N_12250,N_12101,N_12141);
nand U12251 (N_12251,N_12034,N_12185);
and U12252 (N_12252,N_12020,N_12082);
and U12253 (N_12253,N_12024,N_12154);
and U12254 (N_12254,N_12085,N_12017);
and U12255 (N_12255,N_12159,N_12046);
nand U12256 (N_12256,N_12122,N_12048);
and U12257 (N_12257,N_12044,N_12191);
nand U12258 (N_12258,N_12151,N_12105);
and U12259 (N_12259,N_12010,N_12160);
and U12260 (N_12260,N_12003,N_12093);
nand U12261 (N_12261,N_12077,N_12079);
and U12262 (N_12262,N_12184,N_12006);
or U12263 (N_12263,N_12174,N_12177);
nand U12264 (N_12264,N_12000,N_12103);
nand U12265 (N_12265,N_12036,N_12146);
xnor U12266 (N_12266,N_12150,N_12197);
nor U12267 (N_12267,N_12029,N_12033);
or U12268 (N_12268,N_12102,N_12106);
nand U12269 (N_12269,N_12067,N_12121);
and U12270 (N_12270,N_12134,N_12126);
nand U12271 (N_12271,N_12120,N_12193);
and U12272 (N_12272,N_12181,N_12059);
or U12273 (N_12273,N_12195,N_12001);
and U12274 (N_12274,N_12139,N_12142);
or U12275 (N_12275,N_12189,N_12073);
or U12276 (N_12276,N_12037,N_12136);
and U12277 (N_12277,N_12112,N_12182);
or U12278 (N_12278,N_12110,N_12019);
nand U12279 (N_12279,N_12111,N_12070);
nor U12280 (N_12280,N_12043,N_12099);
or U12281 (N_12281,N_12140,N_12004);
nor U12282 (N_12282,N_12087,N_12045);
nand U12283 (N_12283,N_12135,N_12183);
and U12284 (N_12284,N_12041,N_12170);
nor U12285 (N_12285,N_12092,N_12080);
or U12286 (N_12286,N_12075,N_12091);
or U12287 (N_12287,N_12027,N_12088);
nand U12288 (N_12288,N_12123,N_12152);
nor U12289 (N_12289,N_12052,N_12127);
and U12290 (N_12290,N_12118,N_12132);
nand U12291 (N_12291,N_12039,N_12068);
or U12292 (N_12292,N_12053,N_12186);
or U12293 (N_12293,N_12072,N_12008);
or U12294 (N_12294,N_12194,N_12145);
nand U12295 (N_12295,N_12086,N_12049);
nand U12296 (N_12296,N_12169,N_12125);
nand U12297 (N_12297,N_12107,N_12171);
nand U12298 (N_12298,N_12167,N_12143);
nor U12299 (N_12299,N_12007,N_12081);
nor U12300 (N_12300,N_12110,N_12159);
and U12301 (N_12301,N_12123,N_12048);
or U12302 (N_12302,N_12068,N_12157);
nand U12303 (N_12303,N_12106,N_12119);
and U12304 (N_12304,N_12185,N_12083);
nand U12305 (N_12305,N_12013,N_12104);
xor U12306 (N_12306,N_12092,N_12060);
nand U12307 (N_12307,N_12116,N_12017);
nand U12308 (N_12308,N_12089,N_12068);
and U12309 (N_12309,N_12180,N_12055);
or U12310 (N_12310,N_12017,N_12185);
nor U12311 (N_12311,N_12079,N_12039);
or U12312 (N_12312,N_12093,N_12138);
nand U12313 (N_12313,N_12070,N_12058);
or U12314 (N_12314,N_12138,N_12001);
nand U12315 (N_12315,N_12092,N_12074);
nor U12316 (N_12316,N_12062,N_12053);
nor U12317 (N_12317,N_12013,N_12075);
and U12318 (N_12318,N_12030,N_12161);
nand U12319 (N_12319,N_12159,N_12080);
nor U12320 (N_12320,N_12010,N_12113);
nor U12321 (N_12321,N_12134,N_12186);
and U12322 (N_12322,N_12075,N_12198);
nand U12323 (N_12323,N_12023,N_12128);
nor U12324 (N_12324,N_12081,N_12013);
or U12325 (N_12325,N_12090,N_12138);
and U12326 (N_12326,N_12038,N_12147);
nand U12327 (N_12327,N_12151,N_12187);
xnor U12328 (N_12328,N_12068,N_12070);
nor U12329 (N_12329,N_12060,N_12100);
and U12330 (N_12330,N_12165,N_12189);
nor U12331 (N_12331,N_12081,N_12185);
or U12332 (N_12332,N_12131,N_12099);
and U12333 (N_12333,N_12144,N_12066);
nor U12334 (N_12334,N_12182,N_12118);
nand U12335 (N_12335,N_12074,N_12067);
nor U12336 (N_12336,N_12095,N_12003);
or U12337 (N_12337,N_12122,N_12053);
nand U12338 (N_12338,N_12162,N_12164);
nand U12339 (N_12339,N_12058,N_12011);
or U12340 (N_12340,N_12133,N_12152);
nand U12341 (N_12341,N_12072,N_12181);
nand U12342 (N_12342,N_12035,N_12049);
xor U12343 (N_12343,N_12177,N_12108);
and U12344 (N_12344,N_12195,N_12097);
nor U12345 (N_12345,N_12002,N_12169);
or U12346 (N_12346,N_12006,N_12061);
xor U12347 (N_12347,N_12117,N_12003);
nor U12348 (N_12348,N_12135,N_12126);
and U12349 (N_12349,N_12031,N_12075);
nor U12350 (N_12350,N_12010,N_12171);
nand U12351 (N_12351,N_12171,N_12156);
and U12352 (N_12352,N_12048,N_12046);
nor U12353 (N_12353,N_12047,N_12119);
or U12354 (N_12354,N_12005,N_12095);
nand U12355 (N_12355,N_12117,N_12078);
nand U12356 (N_12356,N_12016,N_12043);
nor U12357 (N_12357,N_12000,N_12161);
nand U12358 (N_12358,N_12060,N_12014);
and U12359 (N_12359,N_12183,N_12179);
nand U12360 (N_12360,N_12127,N_12169);
nand U12361 (N_12361,N_12007,N_12135);
nor U12362 (N_12362,N_12123,N_12159);
and U12363 (N_12363,N_12017,N_12023);
nor U12364 (N_12364,N_12108,N_12028);
or U12365 (N_12365,N_12029,N_12054);
and U12366 (N_12366,N_12114,N_12098);
nor U12367 (N_12367,N_12035,N_12021);
and U12368 (N_12368,N_12165,N_12052);
and U12369 (N_12369,N_12004,N_12161);
and U12370 (N_12370,N_12177,N_12028);
nand U12371 (N_12371,N_12019,N_12039);
and U12372 (N_12372,N_12049,N_12057);
nand U12373 (N_12373,N_12027,N_12009);
nor U12374 (N_12374,N_12100,N_12139);
and U12375 (N_12375,N_12077,N_12049);
or U12376 (N_12376,N_12098,N_12020);
nand U12377 (N_12377,N_12078,N_12116);
or U12378 (N_12378,N_12009,N_12086);
or U12379 (N_12379,N_12082,N_12109);
or U12380 (N_12380,N_12046,N_12118);
or U12381 (N_12381,N_12112,N_12024);
nand U12382 (N_12382,N_12079,N_12167);
nor U12383 (N_12383,N_12068,N_12153);
nand U12384 (N_12384,N_12084,N_12013);
nor U12385 (N_12385,N_12111,N_12195);
nand U12386 (N_12386,N_12140,N_12044);
or U12387 (N_12387,N_12190,N_12090);
nand U12388 (N_12388,N_12161,N_12050);
and U12389 (N_12389,N_12066,N_12106);
and U12390 (N_12390,N_12027,N_12087);
nor U12391 (N_12391,N_12092,N_12072);
nor U12392 (N_12392,N_12129,N_12163);
or U12393 (N_12393,N_12125,N_12178);
and U12394 (N_12394,N_12069,N_12022);
nor U12395 (N_12395,N_12117,N_12011);
and U12396 (N_12396,N_12065,N_12142);
and U12397 (N_12397,N_12140,N_12174);
and U12398 (N_12398,N_12042,N_12022);
and U12399 (N_12399,N_12156,N_12007);
xnor U12400 (N_12400,N_12201,N_12378);
nand U12401 (N_12401,N_12271,N_12211);
and U12402 (N_12402,N_12339,N_12244);
and U12403 (N_12403,N_12368,N_12299);
nor U12404 (N_12404,N_12349,N_12372);
nand U12405 (N_12405,N_12386,N_12256);
nand U12406 (N_12406,N_12219,N_12303);
nand U12407 (N_12407,N_12379,N_12344);
nand U12408 (N_12408,N_12230,N_12311);
nor U12409 (N_12409,N_12218,N_12280);
or U12410 (N_12410,N_12321,N_12269);
or U12411 (N_12411,N_12340,N_12253);
nand U12412 (N_12412,N_12320,N_12291);
or U12413 (N_12413,N_12277,N_12364);
nor U12414 (N_12414,N_12210,N_12351);
nor U12415 (N_12415,N_12359,N_12394);
nor U12416 (N_12416,N_12264,N_12258);
nand U12417 (N_12417,N_12398,N_12318);
and U12418 (N_12418,N_12248,N_12384);
or U12419 (N_12419,N_12366,N_12262);
nand U12420 (N_12420,N_12371,N_12385);
nand U12421 (N_12421,N_12282,N_12236);
or U12422 (N_12422,N_12246,N_12273);
and U12423 (N_12423,N_12322,N_12206);
and U12424 (N_12424,N_12346,N_12239);
or U12425 (N_12425,N_12268,N_12361);
and U12426 (N_12426,N_12334,N_12250);
or U12427 (N_12427,N_12352,N_12267);
nand U12428 (N_12428,N_12216,N_12313);
nor U12429 (N_12429,N_12343,N_12284);
or U12430 (N_12430,N_12279,N_12336);
and U12431 (N_12431,N_12305,N_12209);
or U12432 (N_12432,N_12380,N_12274);
nor U12433 (N_12433,N_12254,N_12214);
or U12434 (N_12434,N_12288,N_12222);
nor U12435 (N_12435,N_12243,N_12393);
nand U12436 (N_12436,N_12332,N_12231);
and U12437 (N_12437,N_12247,N_12245);
nor U12438 (N_12438,N_12375,N_12241);
or U12439 (N_12439,N_12353,N_12221);
or U12440 (N_12440,N_12286,N_12227);
and U12441 (N_12441,N_12272,N_12345);
and U12442 (N_12442,N_12229,N_12381);
or U12443 (N_12443,N_12324,N_12217);
or U12444 (N_12444,N_12326,N_12342);
or U12445 (N_12445,N_12281,N_12377);
nand U12446 (N_12446,N_12213,N_12204);
nor U12447 (N_12447,N_12235,N_12337);
and U12448 (N_12448,N_12207,N_12355);
or U12449 (N_12449,N_12276,N_12360);
or U12450 (N_12450,N_12263,N_12370);
nand U12451 (N_12451,N_12260,N_12348);
nor U12452 (N_12452,N_12232,N_12327);
nor U12453 (N_12453,N_12323,N_12233);
or U12454 (N_12454,N_12301,N_12328);
or U12455 (N_12455,N_12293,N_12252);
nor U12456 (N_12456,N_12369,N_12338);
or U12457 (N_12457,N_12354,N_12285);
xor U12458 (N_12458,N_12283,N_12397);
or U12459 (N_12459,N_12240,N_12315);
xor U12460 (N_12460,N_12257,N_12396);
nand U12461 (N_12461,N_12391,N_12387);
and U12462 (N_12462,N_12278,N_12215);
and U12463 (N_12463,N_12316,N_12325);
nand U12464 (N_12464,N_12399,N_12202);
and U12465 (N_12465,N_12226,N_12295);
or U12466 (N_12466,N_12266,N_12304);
or U12467 (N_12467,N_12200,N_12358);
nand U12468 (N_12468,N_12298,N_12237);
or U12469 (N_12469,N_12389,N_12357);
nand U12470 (N_12470,N_12312,N_12297);
and U12471 (N_12471,N_12270,N_12212);
nor U12472 (N_12472,N_12350,N_12317);
xnor U12473 (N_12473,N_12294,N_12309);
xor U12474 (N_12474,N_12388,N_12225);
xnor U12475 (N_12475,N_12335,N_12392);
and U12476 (N_12476,N_12265,N_12234);
nor U12477 (N_12477,N_12255,N_12382);
or U12478 (N_12478,N_12296,N_12333);
and U12479 (N_12479,N_12356,N_12287);
nor U12480 (N_12480,N_12238,N_12292);
nor U12481 (N_12481,N_12205,N_12341);
and U12482 (N_12482,N_12362,N_12365);
or U12483 (N_12483,N_12224,N_12373);
nor U12484 (N_12484,N_12390,N_12314);
or U12485 (N_12485,N_12208,N_12363);
and U12486 (N_12486,N_12331,N_12374);
and U12487 (N_12487,N_12251,N_12395);
nand U12488 (N_12488,N_12347,N_12383);
nor U12489 (N_12489,N_12367,N_12249);
nor U12490 (N_12490,N_12319,N_12300);
nor U12491 (N_12491,N_12308,N_12259);
or U12492 (N_12492,N_12289,N_12302);
and U12493 (N_12493,N_12376,N_12223);
and U12494 (N_12494,N_12330,N_12307);
nand U12495 (N_12495,N_12220,N_12310);
and U12496 (N_12496,N_12329,N_12242);
nand U12497 (N_12497,N_12261,N_12290);
or U12498 (N_12498,N_12275,N_12306);
nor U12499 (N_12499,N_12203,N_12228);
nand U12500 (N_12500,N_12330,N_12324);
xor U12501 (N_12501,N_12284,N_12385);
or U12502 (N_12502,N_12299,N_12313);
nand U12503 (N_12503,N_12357,N_12385);
and U12504 (N_12504,N_12261,N_12216);
nand U12505 (N_12505,N_12261,N_12374);
nor U12506 (N_12506,N_12215,N_12259);
nand U12507 (N_12507,N_12321,N_12399);
or U12508 (N_12508,N_12292,N_12243);
nor U12509 (N_12509,N_12218,N_12314);
and U12510 (N_12510,N_12333,N_12367);
nor U12511 (N_12511,N_12286,N_12274);
nand U12512 (N_12512,N_12245,N_12222);
nand U12513 (N_12513,N_12341,N_12275);
and U12514 (N_12514,N_12285,N_12379);
or U12515 (N_12515,N_12213,N_12334);
or U12516 (N_12516,N_12254,N_12389);
nand U12517 (N_12517,N_12391,N_12342);
xor U12518 (N_12518,N_12208,N_12343);
or U12519 (N_12519,N_12260,N_12291);
nor U12520 (N_12520,N_12396,N_12264);
and U12521 (N_12521,N_12268,N_12221);
nor U12522 (N_12522,N_12300,N_12223);
nand U12523 (N_12523,N_12231,N_12352);
nand U12524 (N_12524,N_12259,N_12212);
nor U12525 (N_12525,N_12305,N_12287);
and U12526 (N_12526,N_12370,N_12228);
and U12527 (N_12527,N_12294,N_12202);
or U12528 (N_12528,N_12394,N_12236);
xor U12529 (N_12529,N_12226,N_12279);
or U12530 (N_12530,N_12229,N_12316);
nor U12531 (N_12531,N_12343,N_12378);
and U12532 (N_12532,N_12225,N_12209);
nor U12533 (N_12533,N_12380,N_12251);
nor U12534 (N_12534,N_12224,N_12388);
xor U12535 (N_12535,N_12313,N_12326);
nand U12536 (N_12536,N_12202,N_12314);
or U12537 (N_12537,N_12338,N_12278);
nand U12538 (N_12538,N_12311,N_12348);
or U12539 (N_12539,N_12372,N_12272);
or U12540 (N_12540,N_12327,N_12239);
nand U12541 (N_12541,N_12373,N_12377);
nand U12542 (N_12542,N_12383,N_12220);
and U12543 (N_12543,N_12312,N_12348);
and U12544 (N_12544,N_12329,N_12344);
and U12545 (N_12545,N_12348,N_12270);
xor U12546 (N_12546,N_12288,N_12361);
xor U12547 (N_12547,N_12340,N_12239);
nand U12548 (N_12548,N_12317,N_12214);
and U12549 (N_12549,N_12358,N_12332);
and U12550 (N_12550,N_12219,N_12261);
or U12551 (N_12551,N_12323,N_12263);
nand U12552 (N_12552,N_12338,N_12252);
and U12553 (N_12553,N_12204,N_12264);
or U12554 (N_12554,N_12204,N_12383);
and U12555 (N_12555,N_12307,N_12260);
or U12556 (N_12556,N_12227,N_12261);
nor U12557 (N_12557,N_12396,N_12235);
nand U12558 (N_12558,N_12362,N_12243);
nor U12559 (N_12559,N_12241,N_12296);
and U12560 (N_12560,N_12335,N_12210);
and U12561 (N_12561,N_12336,N_12204);
nor U12562 (N_12562,N_12268,N_12224);
nor U12563 (N_12563,N_12323,N_12311);
nand U12564 (N_12564,N_12224,N_12231);
and U12565 (N_12565,N_12278,N_12204);
nand U12566 (N_12566,N_12270,N_12246);
or U12567 (N_12567,N_12382,N_12379);
nor U12568 (N_12568,N_12317,N_12364);
or U12569 (N_12569,N_12234,N_12303);
xnor U12570 (N_12570,N_12252,N_12341);
nand U12571 (N_12571,N_12352,N_12377);
nor U12572 (N_12572,N_12243,N_12390);
and U12573 (N_12573,N_12374,N_12388);
nor U12574 (N_12574,N_12238,N_12291);
or U12575 (N_12575,N_12260,N_12253);
nor U12576 (N_12576,N_12272,N_12200);
and U12577 (N_12577,N_12265,N_12309);
nor U12578 (N_12578,N_12304,N_12380);
nand U12579 (N_12579,N_12325,N_12306);
nor U12580 (N_12580,N_12323,N_12258);
or U12581 (N_12581,N_12349,N_12325);
or U12582 (N_12582,N_12329,N_12314);
or U12583 (N_12583,N_12269,N_12237);
nor U12584 (N_12584,N_12280,N_12254);
or U12585 (N_12585,N_12346,N_12261);
nor U12586 (N_12586,N_12234,N_12393);
nand U12587 (N_12587,N_12232,N_12280);
nor U12588 (N_12588,N_12294,N_12207);
and U12589 (N_12589,N_12265,N_12257);
or U12590 (N_12590,N_12265,N_12335);
nand U12591 (N_12591,N_12264,N_12266);
nand U12592 (N_12592,N_12331,N_12321);
nor U12593 (N_12593,N_12255,N_12318);
or U12594 (N_12594,N_12240,N_12298);
and U12595 (N_12595,N_12279,N_12250);
and U12596 (N_12596,N_12349,N_12361);
nand U12597 (N_12597,N_12350,N_12291);
nand U12598 (N_12598,N_12392,N_12367);
or U12599 (N_12599,N_12353,N_12255);
or U12600 (N_12600,N_12419,N_12448);
nor U12601 (N_12601,N_12591,N_12589);
and U12602 (N_12602,N_12551,N_12532);
and U12603 (N_12603,N_12533,N_12476);
or U12604 (N_12604,N_12430,N_12574);
nand U12605 (N_12605,N_12545,N_12537);
or U12606 (N_12606,N_12525,N_12534);
nand U12607 (N_12607,N_12540,N_12413);
and U12608 (N_12608,N_12406,N_12546);
nand U12609 (N_12609,N_12426,N_12424);
and U12610 (N_12610,N_12513,N_12556);
nor U12611 (N_12611,N_12446,N_12455);
nand U12612 (N_12612,N_12434,N_12590);
nor U12613 (N_12613,N_12414,N_12437);
or U12614 (N_12614,N_12432,N_12599);
nor U12615 (N_12615,N_12529,N_12484);
nand U12616 (N_12616,N_12465,N_12597);
and U12617 (N_12617,N_12452,N_12527);
and U12618 (N_12618,N_12565,N_12412);
nor U12619 (N_12619,N_12548,N_12421);
and U12620 (N_12620,N_12415,N_12582);
or U12621 (N_12621,N_12555,N_12498);
and U12622 (N_12622,N_12468,N_12463);
or U12623 (N_12623,N_12439,N_12571);
xor U12624 (N_12624,N_12524,N_12487);
nand U12625 (N_12625,N_12445,N_12568);
nor U12626 (N_12626,N_12595,N_12536);
nand U12627 (N_12627,N_12442,N_12515);
nor U12628 (N_12628,N_12418,N_12499);
or U12629 (N_12629,N_12403,N_12497);
nand U12630 (N_12630,N_12443,N_12423);
or U12631 (N_12631,N_12526,N_12538);
and U12632 (N_12632,N_12504,N_12549);
or U12633 (N_12633,N_12454,N_12422);
and U12634 (N_12634,N_12411,N_12462);
nand U12635 (N_12635,N_12510,N_12508);
xor U12636 (N_12636,N_12501,N_12486);
nor U12637 (N_12637,N_12466,N_12552);
nor U12638 (N_12638,N_12559,N_12593);
nand U12639 (N_12639,N_12431,N_12461);
and U12640 (N_12640,N_12509,N_12436);
nor U12641 (N_12641,N_12428,N_12520);
or U12642 (N_12642,N_12457,N_12472);
and U12643 (N_12643,N_12459,N_12512);
and U12644 (N_12644,N_12456,N_12519);
and U12645 (N_12645,N_12410,N_12473);
nor U12646 (N_12646,N_12417,N_12514);
or U12647 (N_12647,N_12560,N_12596);
or U12648 (N_12648,N_12573,N_12507);
and U12649 (N_12649,N_12493,N_12592);
and U12650 (N_12650,N_12516,N_12429);
and U12651 (N_12651,N_12495,N_12469);
or U12652 (N_12652,N_12404,N_12594);
and U12653 (N_12653,N_12587,N_12492);
or U12654 (N_12654,N_12547,N_12542);
and U12655 (N_12655,N_12578,N_12488);
nand U12656 (N_12656,N_12440,N_12407);
and U12657 (N_12657,N_12543,N_12447);
or U12658 (N_12658,N_12577,N_12564);
nand U12659 (N_12659,N_12401,N_12598);
or U12660 (N_12660,N_12458,N_12505);
and U12661 (N_12661,N_12464,N_12531);
nand U12662 (N_12662,N_12474,N_12522);
nor U12663 (N_12663,N_12580,N_12579);
nand U12664 (N_12664,N_12584,N_12482);
nand U12665 (N_12665,N_12518,N_12544);
nand U12666 (N_12666,N_12517,N_12530);
nand U12667 (N_12667,N_12586,N_12450);
xor U12668 (N_12668,N_12427,N_12554);
and U12669 (N_12669,N_12563,N_12480);
and U12670 (N_12670,N_12500,N_12535);
and U12671 (N_12671,N_12471,N_12528);
or U12672 (N_12672,N_12503,N_12405);
nor U12673 (N_12673,N_12581,N_12477);
nand U12674 (N_12674,N_12569,N_12494);
or U12675 (N_12675,N_12402,N_12408);
and U12676 (N_12676,N_12441,N_12583);
nand U12677 (N_12677,N_12562,N_12572);
nand U12678 (N_12678,N_12425,N_12416);
and U12679 (N_12679,N_12485,N_12483);
xor U12680 (N_12680,N_12444,N_12511);
or U12681 (N_12681,N_12539,N_12478);
nor U12682 (N_12682,N_12470,N_12453);
nor U12683 (N_12683,N_12523,N_12550);
and U12684 (N_12684,N_12467,N_12420);
or U12685 (N_12685,N_12489,N_12576);
or U12686 (N_12686,N_12433,N_12491);
and U12687 (N_12687,N_12496,N_12575);
xor U12688 (N_12688,N_12567,N_12502);
and U12689 (N_12689,N_12481,N_12490);
or U12690 (N_12690,N_12570,N_12566);
nor U12691 (N_12691,N_12475,N_12460);
nor U12692 (N_12692,N_12409,N_12435);
and U12693 (N_12693,N_12400,N_12553);
and U12694 (N_12694,N_12506,N_12541);
nor U12695 (N_12695,N_12557,N_12561);
and U12696 (N_12696,N_12438,N_12585);
nand U12697 (N_12697,N_12479,N_12451);
nor U12698 (N_12698,N_12588,N_12449);
nor U12699 (N_12699,N_12521,N_12558);
nand U12700 (N_12700,N_12439,N_12570);
nor U12701 (N_12701,N_12478,N_12494);
or U12702 (N_12702,N_12492,N_12540);
nor U12703 (N_12703,N_12412,N_12518);
nand U12704 (N_12704,N_12490,N_12582);
nor U12705 (N_12705,N_12565,N_12486);
nand U12706 (N_12706,N_12426,N_12489);
or U12707 (N_12707,N_12484,N_12462);
and U12708 (N_12708,N_12411,N_12415);
nand U12709 (N_12709,N_12411,N_12586);
and U12710 (N_12710,N_12515,N_12416);
nand U12711 (N_12711,N_12584,N_12504);
or U12712 (N_12712,N_12589,N_12492);
or U12713 (N_12713,N_12587,N_12502);
nor U12714 (N_12714,N_12503,N_12594);
nand U12715 (N_12715,N_12443,N_12449);
nor U12716 (N_12716,N_12518,N_12540);
nor U12717 (N_12717,N_12422,N_12431);
and U12718 (N_12718,N_12570,N_12483);
or U12719 (N_12719,N_12551,N_12408);
nor U12720 (N_12720,N_12431,N_12502);
nor U12721 (N_12721,N_12560,N_12553);
or U12722 (N_12722,N_12533,N_12565);
or U12723 (N_12723,N_12574,N_12584);
or U12724 (N_12724,N_12456,N_12472);
or U12725 (N_12725,N_12404,N_12547);
and U12726 (N_12726,N_12513,N_12481);
or U12727 (N_12727,N_12406,N_12453);
xnor U12728 (N_12728,N_12485,N_12522);
and U12729 (N_12729,N_12571,N_12451);
and U12730 (N_12730,N_12582,N_12565);
nand U12731 (N_12731,N_12541,N_12454);
nand U12732 (N_12732,N_12428,N_12584);
nor U12733 (N_12733,N_12499,N_12509);
nand U12734 (N_12734,N_12418,N_12528);
and U12735 (N_12735,N_12420,N_12526);
or U12736 (N_12736,N_12518,N_12435);
or U12737 (N_12737,N_12567,N_12487);
and U12738 (N_12738,N_12427,N_12546);
xnor U12739 (N_12739,N_12414,N_12474);
or U12740 (N_12740,N_12562,N_12561);
and U12741 (N_12741,N_12587,N_12593);
nand U12742 (N_12742,N_12493,N_12470);
nand U12743 (N_12743,N_12491,N_12435);
or U12744 (N_12744,N_12519,N_12542);
or U12745 (N_12745,N_12565,N_12454);
or U12746 (N_12746,N_12481,N_12581);
or U12747 (N_12747,N_12440,N_12532);
nand U12748 (N_12748,N_12573,N_12560);
or U12749 (N_12749,N_12594,N_12521);
nor U12750 (N_12750,N_12558,N_12475);
nand U12751 (N_12751,N_12483,N_12466);
nor U12752 (N_12752,N_12589,N_12516);
or U12753 (N_12753,N_12565,N_12555);
or U12754 (N_12754,N_12533,N_12508);
or U12755 (N_12755,N_12480,N_12473);
or U12756 (N_12756,N_12505,N_12564);
xor U12757 (N_12757,N_12546,N_12593);
nand U12758 (N_12758,N_12545,N_12585);
and U12759 (N_12759,N_12422,N_12406);
and U12760 (N_12760,N_12564,N_12465);
nand U12761 (N_12761,N_12552,N_12599);
nor U12762 (N_12762,N_12472,N_12544);
nor U12763 (N_12763,N_12440,N_12467);
nand U12764 (N_12764,N_12550,N_12472);
and U12765 (N_12765,N_12421,N_12537);
and U12766 (N_12766,N_12566,N_12451);
nand U12767 (N_12767,N_12408,N_12528);
nand U12768 (N_12768,N_12548,N_12439);
nor U12769 (N_12769,N_12444,N_12469);
or U12770 (N_12770,N_12596,N_12587);
and U12771 (N_12771,N_12505,N_12551);
or U12772 (N_12772,N_12506,N_12591);
and U12773 (N_12773,N_12533,N_12442);
or U12774 (N_12774,N_12513,N_12486);
and U12775 (N_12775,N_12420,N_12524);
or U12776 (N_12776,N_12446,N_12401);
and U12777 (N_12777,N_12507,N_12514);
nor U12778 (N_12778,N_12472,N_12536);
or U12779 (N_12779,N_12530,N_12575);
and U12780 (N_12780,N_12569,N_12510);
and U12781 (N_12781,N_12426,N_12484);
and U12782 (N_12782,N_12573,N_12518);
nor U12783 (N_12783,N_12531,N_12592);
nor U12784 (N_12784,N_12546,N_12505);
and U12785 (N_12785,N_12463,N_12420);
nor U12786 (N_12786,N_12539,N_12472);
nand U12787 (N_12787,N_12573,N_12460);
or U12788 (N_12788,N_12563,N_12595);
and U12789 (N_12789,N_12449,N_12575);
or U12790 (N_12790,N_12540,N_12568);
or U12791 (N_12791,N_12578,N_12515);
and U12792 (N_12792,N_12588,N_12560);
and U12793 (N_12793,N_12593,N_12557);
nor U12794 (N_12794,N_12520,N_12431);
and U12795 (N_12795,N_12419,N_12481);
nor U12796 (N_12796,N_12429,N_12448);
nor U12797 (N_12797,N_12488,N_12520);
nor U12798 (N_12798,N_12543,N_12570);
nor U12799 (N_12799,N_12501,N_12417);
nand U12800 (N_12800,N_12748,N_12604);
or U12801 (N_12801,N_12657,N_12640);
nor U12802 (N_12802,N_12765,N_12625);
or U12803 (N_12803,N_12707,N_12697);
or U12804 (N_12804,N_12727,N_12614);
nor U12805 (N_12805,N_12655,N_12732);
nor U12806 (N_12806,N_12670,N_12767);
nand U12807 (N_12807,N_12665,N_12674);
or U12808 (N_12808,N_12624,N_12742);
and U12809 (N_12809,N_12631,N_12608);
or U12810 (N_12810,N_12743,N_12684);
and U12811 (N_12811,N_12620,N_12724);
nor U12812 (N_12812,N_12796,N_12781);
or U12813 (N_12813,N_12686,N_12760);
nand U12814 (N_12814,N_12616,N_12648);
or U12815 (N_12815,N_12696,N_12761);
nor U12816 (N_12816,N_12646,N_12744);
nand U12817 (N_12817,N_12641,N_12615);
or U12818 (N_12818,N_12714,N_12676);
nand U12819 (N_12819,N_12688,N_12662);
nor U12820 (N_12820,N_12692,N_12746);
or U12821 (N_12821,N_12764,N_12629);
nand U12822 (N_12822,N_12755,N_12651);
nand U12823 (N_12823,N_12789,N_12721);
and U12824 (N_12824,N_12605,N_12720);
nand U12825 (N_12825,N_12770,N_12647);
nand U12826 (N_12826,N_12689,N_12638);
nor U12827 (N_12827,N_12795,N_12787);
nand U12828 (N_12828,N_12705,N_12792);
or U12829 (N_12829,N_12741,N_12667);
nor U12830 (N_12830,N_12734,N_12610);
or U12831 (N_12831,N_12630,N_12680);
nor U12832 (N_12832,N_12603,N_12658);
or U12833 (N_12833,N_12611,N_12715);
nor U12834 (N_12834,N_12766,N_12784);
nor U12835 (N_12835,N_12683,N_12659);
nand U12836 (N_12836,N_12762,N_12699);
nor U12837 (N_12837,N_12704,N_12790);
nor U12838 (N_12838,N_12643,N_12606);
or U12839 (N_12839,N_12769,N_12799);
or U12840 (N_12840,N_12708,N_12702);
nand U12841 (N_12841,N_12717,N_12713);
nor U12842 (N_12842,N_12730,N_12709);
and U12843 (N_12843,N_12602,N_12642);
xor U12844 (N_12844,N_12750,N_12706);
or U12845 (N_12845,N_12726,N_12712);
nand U12846 (N_12846,N_12740,N_12664);
nand U12847 (N_12847,N_12645,N_12798);
or U12848 (N_12848,N_12666,N_12691);
and U12849 (N_12849,N_12749,N_12754);
nor U12850 (N_12850,N_12700,N_12785);
and U12851 (N_12851,N_12729,N_12679);
nand U12852 (N_12852,N_12780,N_12671);
or U12853 (N_12853,N_12622,N_12735);
or U12854 (N_12854,N_12627,N_12786);
nor U12855 (N_12855,N_12768,N_12653);
or U12856 (N_12856,N_12636,N_12621);
nor U12857 (N_12857,N_12772,N_12695);
nand U12858 (N_12858,N_12752,N_12633);
nor U12859 (N_12859,N_12600,N_12779);
and U12860 (N_12860,N_12723,N_12771);
nand U12861 (N_12861,N_12672,N_12678);
and U12862 (N_12862,N_12673,N_12736);
or U12863 (N_12863,N_12698,N_12701);
and U12864 (N_12864,N_12677,N_12751);
nand U12865 (N_12865,N_12618,N_12660);
or U12866 (N_12866,N_12797,N_12628);
or U12867 (N_12867,N_12711,N_12733);
nor U12868 (N_12868,N_12650,N_12632);
and U12869 (N_12869,N_12791,N_12668);
xnor U12870 (N_12870,N_12639,N_12681);
or U12871 (N_12871,N_12644,N_12617);
or U12872 (N_12872,N_12663,N_12775);
nor U12873 (N_12873,N_12793,N_12656);
nor U12874 (N_12874,N_12669,N_12778);
and U12875 (N_12875,N_12719,N_12685);
and U12876 (N_12876,N_12619,N_12693);
or U12877 (N_12877,N_12773,N_12687);
or U12878 (N_12878,N_12612,N_12782);
and U12879 (N_12879,N_12747,N_12753);
nand U12880 (N_12880,N_12783,N_12718);
nand U12881 (N_12881,N_12703,N_12613);
or U12882 (N_12882,N_12756,N_12637);
nand U12883 (N_12883,N_12728,N_12654);
and U12884 (N_12884,N_12788,N_12634);
or U12885 (N_12885,N_12758,N_12652);
nand U12886 (N_12886,N_12722,N_12738);
nor U12887 (N_12887,N_12649,N_12710);
nand U12888 (N_12888,N_12794,N_12626);
and U12889 (N_12889,N_12601,N_12661);
or U12890 (N_12890,N_12623,N_12609);
or U12891 (N_12891,N_12777,N_12745);
or U12892 (N_12892,N_12682,N_12607);
or U12893 (N_12893,N_12725,N_12716);
and U12894 (N_12894,N_12774,N_12759);
and U12895 (N_12895,N_12763,N_12739);
and U12896 (N_12896,N_12690,N_12635);
nor U12897 (N_12897,N_12757,N_12737);
and U12898 (N_12898,N_12776,N_12675);
nor U12899 (N_12899,N_12731,N_12694);
nand U12900 (N_12900,N_12678,N_12748);
nand U12901 (N_12901,N_12677,N_12782);
nor U12902 (N_12902,N_12715,N_12664);
xor U12903 (N_12903,N_12768,N_12738);
nor U12904 (N_12904,N_12727,N_12788);
nand U12905 (N_12905,N_12604,N_12768);
and U12906 (N_12906,N_12609,N_12663);
nand U12907 (N_12907,N_12640,N_12606);
or U12908 (N_12908,N_12696,N_12622);
nand U12909 (N_12909,N_12734,N_12695);
nor U12910 (N_12910,N_12615,N_12704);
or U12911 (N_12911,N_12695,N_12699);
nor U12912 (N_12912,N_12666,N_12725);
or U12913 (N_12913,N_12721,N_12746);
and U12914 (N_12914,N_12616,N_12664);
or U12915 (N_12915,N_12756,N_12792);
and U12916 (N_12916,N_12740,N_12787);
and U12917 (N_12917,N_12771,N_12679);
nand U12918 (N_12918,N_12664,N_12791);
nand U12919 (N_12919,N_12605,N_12699);
nand U12920 (N_12920,N_12704,N_12761);
or U12921 (N_12921,N_12632,N_12680);
or U12922 (N_12922,N_12712,N_12682);
nor U12923 (N_12923,N_12792,N_12612);
and U12924 (N_12924,N_12642,N_12600);
and U12925 (N_12925,N_12641,N_12604);
nor U12926 (N_12926,N_12635,N_12643);
nor U12927 (N_12927,N_12603,N_12732);
or U12928 (N_12928,N_12684,N_12658);
xnor U12929 (N_12929,N_12717,N_12751);
and U12930 (N_12930,N_12679,N_12637);
or U12931 (N_12931,N_12678,N_12755);
nand U12932 (N_12932,N_12614,N_12733);
or U12933 (N_12933,N_12647,N_12795);
or U12934 (N_12934,N_12663,N_12768);
nand U12935 (N_12935,N_12794,N_12795);
nand U12936 (N_12936,N_12728,N_12674);
nand U12937 (N_12937,N_12715,N_12740);
nor U12938 (N_12938,N_12626,N_12668);
nand U12939 (N_12939,N_12717,N_12740);
and U12940 (N_12940,N_12624,N_12666);
nor U12941 (N_12941,N_12606,N_12638);
nor U12942 (N_12942,N_12721,N_12661);
nand U12943 (N_12943,N_12704,N_12606);
nor U12944 (N_12944,N_12794,N_12674);
and U12945 (N_12945,N_12672,N_12795);
nand U12946 (N_12946,N_12637,N_12742);
nand U12947 (N_12947,N_12676,N_12777);
nor U12948 (N_12948,N_12759,N_12743);
or U12949 (N_12949,N_12765,N_12785);
nor U12950 (N_12950,N_12673,N_12675);
nand U12951 (N_12951,N_12688,N_12625);
and U12952 (N_12952,N_12636,N_12770);
nor U12953 (N_12953,N_12793,N_12742);
nor U12954 (N_12954,N_12736,N_12795);
xor U12955 (N_12955,N_12795,N_12724);
nor U12956 (N_12956,N_12790,N_12789);
or U12957 (N_12957,N_12741,N_12627);
or U12958 (N_12958,N_12679,N_12765);
and U12959 (N_12959,N_12714,N_12763);
or U12960 (N_12960,N_12608,N_12686);
nand U12961 (N_12961,N_12630,N_12757);
and U12962 (N_12962,N_12765,N_12667);
or U12963 (N_12963,N_12764,N_12693);
or U12964 (N_12964,N_12616,N_12736);
and U12965 (N_12965,N_12614,N_12764);
and U12966 (N_12966,N_12767,N_12784);
or U12967 (N_12967,N_12780,N_12698);
nand U12968 (N_12968,N_12728,N_12620);
nand U12969 (N_12969,N_12773,N_12643);
nor U12970 (N_12970,N_12663,N_12744);
nand U12971 (N_12971,N_12700,N_12726);
xnor U12972 (N_12972,N_12638,N_12769);
and U12973 (N_12973,N_12623,N_12740);
nor U12974 (N_12974,N_12676,N_12608);
and U12975 (N_12975,N_12786,N_12632);
or U12976 (N_12976,N_12678,N_12680);
nor U12977 (N_12977,N_12706,N_12627);
xor U12978 (N_12978,N_12662,N_12604);
nand U12979 (N_12979,N_12741,N_12735);
or U12980 (N_12980,N_12753,N_12755);
nand U12981 (N_12981,N_12755,N_12735);
nor U12982 (N_12982,N_12653,N_12787);
nor U12983 (N_12983,N_12665,N_12776);
nand U12984 (N_12984,N_12662,N_12634);
nand U12985 (N_12985,N_12758,N_12641);
nor U12986 (N_12986,N_12788,N_12669);
nand U12987 (N_12987,N_12678,N_12721);
and U12988 (N_12988,N_12708,N_12797);
or U12989 (N_12989,N_12650,N_12750);
nand U12990 (N_12990,N_12782,N_12714);
and U12991 (N_12991,N_12653,N_12771);
nor U12992 (N_12992,N_12696,N_12681);
nor U12993 (N_12993,N_12622,N_12785);
nor U12994 (N_12994,N_12658,N_12621);
nand U12995 (N_12995,N_12739,N_12704);
nand U12996 (N_12996,N_12759,N_12610);
nor U12997 (N_12997,N_12740,N_12655);
nand U12998 (N_12998,N_12758,N_12601);
and U12999 (N_12999,N_12722,N_12743);
nand U13000 (N_13000,N_12908,N_12976);
or U13001 (N_13001,N_12824,N_12887);
nand U13002 (N_13002,N_12919,N_12833);
nor U13003 (N_13003,N_12969,N_12975);
nor U13004 (N_13004,N_12958,N_12942);
or U13005 (N_13005,N_12854,N_12867);
xnor U13006 (N_13006,N_12986,N_12855);
and U13007 (N_13007,N_12924,N_12941);
or U13008 (N_13008,N_12966,N_12960);
and U13009 (N_13009,N_12868,N_12905);
or U13010 (N_13010,N_12999,N_12980);
or U13011 (N_13011,N_12995,N_12815);
or U13012 (N_13012,N_12982,N_12946);
xor U13013 (N_13013,N_12806,N_12820);
nor U13014 (N_13014,N_12923,N_12859);
nand U13015 (N_13015,N_12971,N_12954);
nand U13016 (N_13016,N_12807,N_12996);
and U13017 (N_13017,N_12852,N_12967);
nor U13018 (N_13018,N_12828,N_12907);
or U13019 (N_13019,N_12841,N_12836);
nor U13020 (N_13020,N_12922,N_12876);
nand U13021 (N_13021,N_12803,N_12873);
nand U13022 (N_13022,N_12963,N_12988);
and U13023 (N_13023,N_12962,N_12810);
nand U13024 (N_13024,N_12861,N_12952);
nand U13025 (N_13025,N_12898,N_12865);
nand U13026 (N_13026,N_12827,N_12968);
and U13027 (N_13027,N_12950,N_12929);
nand U13028 (N_13028,N_12818,N_12901);
and U13029 (N_13029,N_12826,N_12805);
and U13030 (N_13030,N_12956,N_12932);
nand U13031 (N_13031,N_12984,N_12850);
and U13032 (N_13032,N_12987,N_12981);
or U13033 (N_13033,N_12838,N_12825);
or U13034 (N_13034,N_12957,N_12910);
nor U13035 (N_13035,N_12893,N_12879);
and U13036 (N_13036,N_12877,N_12916);
nand U13037 (N_13037,N_12902,N_12993);
or U13038 (N_13038,N_12847,N_12939);
nor U13039 (N_13039,N_12851,N_12885);
and U13040 (N_13040,N_12886,N_12937);
nand U13041 (N_13041,N_12991,N_12899);
and U13042 (N_13042,N_12965,N_12953);
or U13043 (N_13043,N_12951,N_12849);
or U13044 (N_13044,N_12983,N_12931);
or U13045 (N_13045,N_12930,N_12881);
nand U13046 (N_13046,N_12871,N_12840);
and U13047 (N_13047,N_12874,N_12921);
or U13048 (N_13048,N_12915,N_12848);
and U13049 (N_13049,N_12853,N_12949);
and U13050 (N_13050,N_12823,N_12830);
nor U13051 (N_13051,N_12945,N_12998);
nor U13052 (N_13052,N_12911,N_12843);
or U13053 (N_13053,N_12977,N_12900);
or U13054 (N_13054,N_12903,N_12989);
nand U13055 (N_13055,N_12912,N_12882);
or U13056 (N_13056,N_12883,N_12846);
nor U13057 (N_13057,N_12940,N_12904);
nor U13058 (N_13058,N_12897,N_12816);
or U13059 (N_13059,N_12804,N_12819);
or U13060 (N_13060,N_12812,N_12866);
or U13061 (N_13061,N_12821,N_12834);
nor U13062 (N_13062,N_12896,N_12890);
nor U13063 (N_13063,N_12974,N_12813);
and U13064 (N_13064,N_12990,N_12891);
nor U13065 (N_13065,N_12884,N_12934);
nand U13066 (N_13066,N_12913,N_12808);
or U13067 (N_13067,N_12858,N_12928);
nand U13068 (N_13068,N_12837,N_12985);
nand U13069 (N_13069,N_12869,N_12800);
or U13070 (N_13070,N_12961,N_12918);
nand U13071 (N_13071,N_12856,N_12978);
nand U13072 (N_13072,N_12889,N_12822);
nor U13073 (N_13073,N_12809,N_12955);
and U13074 (N_13074,N_12863,N_12831);
or U13075 (N_13075,N_12917,N_12895);
nand U13076 (N_13076,N_12875,N_12835);
nor U13077 (N_13077,N_12906,N_12944);
and U13078 (N_13078,N_12914,N_12938);
and U13079 (N_13079,N_12878,N_12925);
nor U13080 (N_13080,N_12927,N_12970);
or U13081 (N_13081,N_12801,N_12964);
or U13082 (N_13082,N_12857,N_12839);
and U13083 (N_13083,N_12880,N_12926);
or U13084 (N_13084,N_12994,N_12844);
or U13085 (N_13085,N_12811,N_12845);
or U13086 (N_13086,N_12997,N_12973);
nand U13087 (N_13087,N_12972,N_12864);
or U13088 (N_13088,N_12959,N_12892);
and U13089 (N_13089,N_12948,N_12832);
or U13090 (N_13090,N_12936,N_12814);
nor U13091 (N_13091,N_12992,N_12872);
and U13092 (N_13092,N_12947,N_12933);
and U13093 (N_13093,N_12894,N_12842);
nand U13094 (N_13094,N_12802,N_12943);
and U13095 (N_13095,N_12979,N_12817);
or U13096 (N_13096,N_12888,N_12935);
or U13097 (N_13097,N_12862,N_12870);
or U13098 (N_13098,N_12860,N_12920);
nand U13099 (N_13099,N_12829,N_12909);
nor U13100 (N_13100,N_12931,N_12810);
nand U13101 (N_13101,N_12977,N_12965);
or U13102 (N_13102,N_12828,N_12856);
nand U13103 (N_13103,N_12807,N_12937);
and U13104 (N_13104,N_12877,N_12801);
nand U13105 (N_13105,N_12817,N_12961);
nand U13106 (N_13106,N_12920,N_12896);
xnor U13107 (N_13107,N_12933,N_12923);
or U13108 (N_13108,N_12933,N_12867);
nor U13109 (N_13109,N_12859,N_12805);
or U13110 (N_13110,N_12961,N_12980);
and U13111 (N_13111,N_12944,N_12883);
or U13112 (N_13112,N_12934,N_12962);
or U13113 (N_13113,N_12850,N_12952);
or U13114 (N_13114,N_12877,N_12936);
nor U13115 (N_13115,N_12951,N_12891);
and U13116 (N_13116,N_12951,N_12978);
nor U13117 (N_13117,N_12933,N_12937);
nor U13118 (N_13118,N_12828,N_12881);
or U13119 (N_13119,N_12972,N_12833);
nor U13120 (N_13120,N_12929,N_12925);
nor U13121 (N_13121,N_12840,N_12920);
or U13122 (N_13122,N_12810,N_12948);
nand U13123 (N_13123,N_12873,N_12975);
and U13124 (N_13124,N_12933,N_12927);
or U13125 (N_13125,N_12942,N_12924);
and U13126 (N_13126,N_12824,N_12945);
xor U13127 (N_13127,N_12896,N_12885);
nand U13128 (N_13128,N_12935,N_12869);
and U13129 (N_13129,N_12949,N_12838);
or U13130 (N_13130,N_12942,N_12928);
nor U13131 (N_13131,N_12916,N_12917);
nand U13132 (N_13132,N_12879,N_12810);
nor U13133 (N_13133,N_12924,N_12988);
and U13134 (N_13134,N_12913,N_12901);
or U13135 (N_13135,N_12851,N_12925);
xnor U13136 (N_13136,N_12895,N_12983);
or U13137 (N_13137,N_12947,N_12957);
nor U13138 (N_13138,N_12843,N_12805);
or U13139 (N_13139,N_12910,N_12935);
nand U13140 (N_13140,N_12805,N_12994);
nand U13141 (N_13141,N_12805,N_12850);
and U13142 (N_13142,N_12894,N_12913);
or U13143 (N_13143,N_12991,N_12919);
xnor U13144 (N_13144,N_12916,N_12872);
and U13145 (N_13145,N_12935,N_12989);
or U13146 (N_13146,N_12895,N_12888);
and U13147 (N_13147,N_12960,N_12910);
nand U13148 (N_13148,N_12947,N_12890);
or U13149 (N_13149,N_12849,N_12907);
and U13150 (N_13150,N_12885,N_12948);
and U13151 (N_13151,N_12804,N_12826);
nor U13152 (N_13152,N_12842,N_12929);
and U13153 (N_13153,N_12823,N_12996);
nor U13154 (N_13154,N_12922,N_12854);
nand U13155 (N_13155,N_12854,N_12965);
nand U13156 (N_13156,N_12961,N_12945);
or U13157 (N_13157,N_12862,N_12927);
nand U13158 (N_13158,N_12824,N_12949);
and U13159 (N_13159,N_12922,N_12821);
or U13160 (N_13160,N_12986,N_12994);
and U13161 (N_13161,N_12939,N_12838);
nand U13162 (N_13162,N_12875,N_12973);
xnor U13163 (N_13163,N_12834,N_12985);
nand U13164 (N_13164,N_12947,N_12958);
nor U13165 (N_13165,N_12914,N_12898);
or U13166 (N_13166,N_12875,N_12898);
nor U13167 (N_13167,N_12980,N_12968);
or U13168 (N_13168,N_12913,N_12848);
nor U13169 (N_13169,N_12863,N_12821);
nand U13170 (N_13170,N_12834,N_12805);
or U13171 (N_13171,N_12809,N_12880);
and U13172 (N_13172,N_12876,N_12829);
and U13173 (N_13173,N_12920,N_12831);
nor U13174 (N_13174,N_12939,N_12857);
or U13175 (N_13175,N_12866,N_12939);
nor U13176 (N_13176,N_12815,N_12864);
nor U13177 (N_13177,N_12905,N_12949);
or U13178 (N_13178,N_12920,N_12998);
nor U13179 (N_13179,N_12907,N_12900);
nor U13180 (N_13180,N_12938,N_12880);
or U13181 (N_13181,N_12959,N_12863);
nor U13182 (N_13182,N_12829,N_12877);
and U13183 (N_13183,N_12930,N_12876);
and U13184 (N_13184,N_12810,N_12909);
and U13185 (N_13185,N_12822,N_12948);
or U13186 (N_13186,N_12911,N_12889);
nand U13187 (N_13187,N_12907,N_12846);
nor U13188 (N_13188,N_12870,N_12954);
and U13189 (N_13189,N_12993,N_12824);
nor U13190 (N_13190,N_12834,N_12829);
and U13191 (N_13191,N_12958,N_12833);
or U13192 (N_13192,N_12949,N_12834);
nor U13193 (N_13193,N_12803,N_12874);
nand U13194 (N_13194,N_12982,N_12831);
or U13195 (N_13195,N_12986,N_12975);
nor U13196 (N_13196,N_12943,N_12935);
and U13197 (N_13197,N_12964,N_12864);
and U13198 (N_13198,N_12869,N_12836);
nand U13199 (N_13199,N_12985,N_12861);
and U13200 (N_13200,N_13136,N_13088);
nand U13201 (N_13201,N_13035,N_13070);
nand U13202 (N_13202,N_13069,N_13109);
nand U13203 (N_13203,N_13064,N_13146);
nor U13204 (N_13204,N_13032,N_13129);
nor U13205 (N_13205,N_13170,N_13186);
and U13206 (N_13206,N_13025,N_13125);
nor U13207 (N_13207,N_13149,N_13138);
and U13208 (N_13208,N_13062,N_13074);
and U13209 (N_13209,N_13050,N_13040);
nand U13210 (N_13210,N_13027,N_13181);
and U13211 (N_13211,N_13018,N_13199);
nor U13212 (N_13212,N_13141,N_13065);
and U13213 (N_13213,N_13108,N_13150);
or U13214 (N_13214,N_13084,N_13082);
nor U13215 (N_13215,N_13179,N_13028);
nand U13216 (N_13216,N_13154,N_13094);
nor U13217 (N_13217,N_13002,N_13176);
nor U13218 (N_13218,N_13111,N_13007);
and U13219 (N_13219,N_13024,N_13083);
or U13220 (N_13220,N_13010,N_13101);
and U13221 (N_13221,N_13049,N_13017);
or U13222 (N_13222,N_13004,N_13197);
and U13223 (N_13223,N_13068,N_13072);
nor U13224 (N_13224,N_13106,N_13080);
nand U13225 (N_13225,N_13172,N_13006);
xor U13226 (N_13226,N_13042,N_13066);
or U13227 (N_13227,N_13051,N_13016);
or U13228 (N_13228,N_13022,N_13081);
xnor U13229 (N_13229,N_13031,N_13118);
and U13230 (N_13230,N_13178,N_13053);
or U13231 (N_13231,N_13183,N_13001);
and U13232 (N_13232,N_13037,N_13063);
nor U13233 (N_13233,N_13153,N_13102);
and U13234 (N_13234,N_13000,N_13071);
nor U13235 (N_13235,N_13126,N_13085);
nand U13236 (N_13236,N_13099,N_13026);
nor U13237 (N_13237,N_13135,N_13029);
and U13238 (N_13238,N_13055,N_13113);
and U13239 (N_13239,N_13078,N_13134);
and U13240 (N_13240,N_13148,N_13090);
nand U13241 (N_13241,N_13155,N_13038);
nand U13242 (N_13242,N_13067,N_13142);
or U13243 (N_13243,N_13009,N_13039);
nand U13244 (N_13244,N_13145,N_13044);
nor U13245 (N_13245,N_13115,N_13046);
nor U13246 (N_13246,N_13097,N_13196);
or U13247 (N_13247,N_13117,N_13087);
and U13248 (N_13248,N_13008,N_13052);
nand U13249 (N_13249,N_13123,N_13079);
nor U13250 (N_13250,N_13048,N_13036);
nor U13251 (N_13251,N_13147,N_13120);
and U13252 (N_13252,N_13107,N_13171);
nor U13253 (N_13253,N_13177,N_13185);
nor U13254 (N_13254,N_13114,N_13015);
nand U13255 (N_13255,N_13021,N_13182);
xor U13256 (N_13256,N_13158,N_13054);
or U13257 (N_13257,N_13034,N_13077);
or U13258 (N_13258,N_13193,N_13165);
or U13259 (N_13259,N_13189,N_13012);
and U13260 (N_13260,N_13089,N_13103);
or U13261 (N_13261,N_13011,N_13169);
xor U13262 (N_13262,N_13093,N_13045);
nand U13263 (N_13263,N_13030,N_13061);
nand U13264 (N_13264,N_13131,N_13060);
or U13265 (N_13265,N_13105,N_13128);
or U13266 (N_13266,N_13163,N_13191);
and U13267 (N_13267,N_13047,N_13175);
and U13268 (N_13268,N_13152,N_13119);
and U13269 (N_13269,N_13073,N_13122);
nor U13270 (N_13270,N_13190,N_13164);
and U13271 (N_13271,N_13121,N_13192);
nand U13272 (N_13272,N_13143,N_13162);
and U13273 (N_13273,N_13058,N_13173);
nor U13274 (N_13274,N_13104,N_13095);
nand U13275 (N_13275,N_13014,N_13023);
and U13276 (N_13276,N_13161,N_13187);
and U13277 (N_13277,N_13166,N_13092);
nor U13278 (N_13278,N_13116,N_13140);
or U13279 (N_13279,N_13020,N_13188);
or U13280 (N_13280,N_13184,N_13096);
nand U13281 (N_13281,N_13156,N_13144);
nor U13282 (N_13282,N_13139,N_13098);
or U13283 (N_13283,N_13174,N_13157);
nor U13284 (N_13284,N_13059,N_13076);
and U13285 (N_13285,N_13159,N_13124);
nor U13286 (N_13286,N_13132,N_13110);
or U13287 (N_13287,N_13075,N_13056);
and U13288 (N_13288,N_13137,N_13151);
nand U13289 (N_13289,N_13133,N_13112);
nor U13290 (N_13290,N_13003,N_13194);
and U13291 (N_13291,N_13043,N_13041);
nand U13292 (N_13292,N_13160,N_13091);
nand U13293 (N_13293,N_13195,N_13057);
and U13294 (N_13294,N_13005,N_13167);
or U13295 (N_13295,N_13130,N_13086);
nand U13296 (N_13296,N_13168,N_13198);
or U13297 (N_13297,N_13019,N_13033);
nor U13298 (N_13298,N_13013,N_13180);
nor U13299 (N_13299,N_13100,N_13127);
and U13300 (N_13300,N_13039,N_13076);
nor U13301 (N_13301,N_13100,N_13082);
nor U13302 (N_13302,N_13048,N_13001);
and U13303 (N_13303,N_13156,N_13178);
or U13304 (N_13304,N_13100,N_13093);
nand U13305 (N_13305,N_13097,N_13142);
or U13306 (N_13306,N_13197,N_13102);
nor U13307 (N_13307,N_13170,N_13135);
and U13308 (N_13308,N_13091,N_13014);
nand U13309 (N_13309,N_13085,N_13150);
nand U13310 (N_13310,N_13189,N_13123);
xor U13311 (N_13311,N_13054,N_13075);
and U13312 (N_13312,N_13193,N_13079);
and U13313 (N_13313,N_13054,N_13065);
or U13314 (N_13314,N_13166,N_13134);
and U13315 (N_13315,N_13017,N_13142);
nand U13316 (N_13316,N_13108,N_13141);
nor U13317 (N_13317,N_13004,N_13120);
nor U13318 (N_13318,N_13107,N_13149);
xnor U13319 (N_13319,N_13071,N_13054);
nor U13320 (N_13320,N_13036,N_13097);
or U13321 (N_13321,N_13024,N_13087);
and U13322 (N_13322,N_13190,N_13077);
nand U13323 (N_13323,N_13168,N_13088);
nand U13324 (N_13324,N_13078,N_13196);
nor U13325 (N_13325,N_13012,N_13105);
or U13326 (N_13326,N_13191,N_13114);
or U13327 (N_13327,N_13193,N_13064);
and U13328 (N_13328,N_13023,N_13074);
nand U13329 (N_13329,N_13096,N_13170);
or U13330 (N_13330,N_13182,N_13172);
nand U13331 (N_13331,N_13097,N_13025);
and U13332 (N_13332,N_13120,N_13155);
nor U13333 (N_13333,N_13008,N_13197);
nand U13334 (N_13334,N_13088,N_13065);
or U13335 (N_13335,N_13059,N_13133);
or U13336 (N_13336,N_13038,N_13188);
xor U13337 (N_13337,N_13081,N_13099);
nor U13338 (N_13338,N_13160,N_13001);
nor U13339 (N_13339,N_13069,N_13153);
nand U13340 (N_13340,N_13184,N_13126);
or U13341 (N_13341,N_13196,N_13143);
or U13342 (N_13342,N_13131,N_13122);
xnor U13343 (N_13343,N_13027,N_13078);
nor U13344 (N_13344,N_13076,N_13137);
and U13345 (N_13345,N_13002,N_13190);
and U13346 (N_13346,N_13184,N_13111);
or U13347 (N_13347,N_13033,N_13037);
and U13348 (N_13348,N_13153,N_13114);
nand U13349 (N_13349,N_13035,N_13109);
xnor U13350 (N_13350,N_13008,N_13036);
nand U13351 (N_13351,N_13081,N_13015);
and U13352 (N_13352,N_13087,N_13157);
nand U13353 (N_13353,N_13122,N_13014);
or U13354 (N_13354,N_13049,N_13007);
nand U13355 (N_13355,N_13038,N_13156);
nand U13356 (N_13356,N_13168,N_13134);
nor U13357 (N_13357,N_13198,N_13151);
and U13358 (N_13358,N_13132,N_13066);
nor U13359 (N_13359,N_13127,N_13007);
nand U13360 (N_13360,N_13070,N_13076);
and U13361 (N_13361,N_13054,N_13122);
nand U13362 (N_13362,N_13062,N_13050);
nand U13363 (N_13363,N_13054,N_13048);
nand U13364 (N_13364,N_13063,N_13180);
nand U13365 (N_13365,N_13001,N_13129);
nor U13366 (N_13366,N_13131,N_13186);
nor U13367 (N_13367,N_13137,N_13089);
and U13368 (N_13368,N_13024,N_13050);
or U13369 (N_13369,N_13178,N_13111);
nor U13370 (N_13370,N_13145,N_13179);
and U13371 (N_13371,N_13003,N_13179);
and U13372 (N_13372,N_13189,N_13195);
or U13373 (N_13373,N_13003,N_13156);
nor U13374 (N_13374,N_13157,N_13066);
or U13375 (N_13375,N_13190,N_13055);
nor U13376 (N_13376,N_13032,N_13116);
nand U13377 (N_13377,N_13075,N_13100);
nor U13378 (N_13378,N_13135,N_13011);
or U13379 (N_13379,N_13186,N_13175);
nand U13380 (N_13380,N_13053,N_13045);
or U13381 (N_13381,N_13154,N_13017);
and U13382 (N_13382,N_13027,N_13117);
nor U13383 (N_13383,N_13120,N_13044);
and U13384 (N_13384,N_13127,N_13183);
or U13385 (N_13385,N_13134,N_13081);
and U13386 (N_13386,N_13189,N_13136);
and U13387 (N_13387,N_13127,N_13041);
or U13388 (N_13388,N_13094,N_13079);
or U13389 (N_13389,N_13179,N_13153);
nand U13390 (N_13390,N_13171,N_13003);
and U13391 (N_13391,N_13022,N_13026);
nor U13392 (N_13392,N_13128,N_13161);
or U13393 (N_13393,N_13199,N_13185);
nand U13394 (N_13394,N_13149,N_13013);
and U13395 (N_13395,N_13092,N_13188);
nor U13396 (N_13396,N_13048,N_13178);
nand U13397 (N_13397,N_13078,N_13142);
or U13398 (N_13398,N_13176,N_13117);
or U13399 (N_13399,N_13073,N_13074);
or U13400 (N_13400,N_13271,N_13397);
xnor U13401 (N_13401,N_13342,N_13236);
and U13402 (N_13402,N_13389,N_13285);
or U13403 (N_13403,N_13265,N_13233);
nor U13404 (N_13404,N_13266,N_13278);
or U13405 (N_13405,N_13373,N_13347);
or U13406 (N_13406,N_13311,N_13307);
and U13407 (N_13407,N_13344,N_13279);
nand U13408 (N_13408,N_13329,N_13354);
nor U13409 (N_13409,N_13201,N_13281);
or U13410 (N_13410,N_13372,N_13375);
or U13411 (N_13411,N_13391,N_13292);
nor U13412 (N_13412,N_13340,N_13222);
or U13413 (N_13413,N_13320,N_13240);
and U13414 (N_13414,N_13352,N_13243);
or U13415 (N_13415,N_13210,N_13386);
nand U13416 (N_13416,N_13218,N_13377);
nand U13417 (N_13417,N_13272,N_13356);
nand U13418 (N_13418,N_13263,N_13254);
nor U13419 (N_13419,N_13288,N_13219);
or U13420 (N_13420,N_13206,N_13255);
nor U13421 (N_13421,N_13246,N_13323);
or U13422 (N_13422,N_13363,N_13269);
and U13423 (N_13423,N_13298,N_13209);
nand U13424 (N_13424,N_13315,N_13286);
nor U13425 (N_13425,N_13290,N_13268);
nor U13426 (N_13426,N_13328,N_13317);
nand U13427 (N_13427,N_13249,N_13383);
nor U13428 (N_13428,N_13302,N_13361);
and U13429 (N_13429,N_13261,N_13225);
and U13430 (N_13430,N_13369,N_13299);
and U13431 (N_13431,N_13245,N_13264);
nor U13432 (N_13432,N_13313,N_13250);
nor U13433 (N_13433,N_13325,N_13384);
nor U13434 (N_13434,N_13208,N_13248);
nand U13435 (N_13435,N_13349,N_13385);
or U13436 (N_13436,N_13394,N_13327);
xor U13437 (N_13437,N_13395,N_13203);
nor U13438 (N_13438,N_13284,N_13223);
nand U13439 (N_13439,N_13220,N_13217);
and U13440 (N_13440,N_13357,N_13312);
and U13441 (N_13441,N_13216,N_13322);
xnor U13442 (N_13442,N_13341,N_13237);
nand U13443 (N_13443,N_13256,N_13213);
or U13444 (N_13444,N_13331,N_13260);
nor U13445 (N_13445,N_13362,N_13259);
nor U13446 (N_13446,N_13234,N_13310);
or U13447 (N_13447,N_13242,N_13300);
nand U13448 (N_13448,N_13293,N_13382);
nand U13449 (N_13449,N_13324,N_13318);
nor U13450 (N_13450,N_13258,N_13321);
nor U13451 (N_13451,N_13283,N_13371);
nor U13452 (N_13452,N_13277,N_13228);
or U13453 (N_13453,N_13304,N_13346);
and U13454 (N_13454,N_13238,N_13337);
nor U13455 (N_13455,N_13287,N_13200);
nand U13456 (N_13456,N_13274,N_13374);
nor U13457 (N_13457,N_13353,N_13332);
nor U13458 (N_13458,N_13244,N_13393);
nor U13459 (N_13459,N_13295,N_13365);
nor U13460 (N_13460,N_13221,N_13205);
and U13461 (N_13461,N_13398,N_13303);
and U13462 (N_13462,N_13229,N_13359);
nor U13463 (N_13463,N_13289,N_13336);
or U13464 (N_13464,N_13297,N_13379);
nand U13465 (N_13465,N_13291,N_13273);
nand U13466 (N_13466,N_13338,N_13276);
nand U13467 (N_13467,N_13360,N_13294);
and U13468 (N_13468,N_13282,N_13392);
nor U13469 (N_13469,N_13316,N_13335);
or U13470 (N_13470,N_13270,N_13326);
and U13471 (N_13471,N_13251,N_13309);
nand U13472 (N_13472,N_13358,N_13253);
or U13473 (N_13473,N_13364,N_13314);
or U13474 (N_13474,N_13224,N_13301);
or U13475 (N_13475,N_13296,N_13226);
nor U13476 (N_13476,N_13381,N_13267);
and U13477 (N_13477,N_13376,N_13239);
nand U13478 (N_13478,N_13252,N_13334);
nand U13479 (N_13479,N_13232,N_13319);
nor U13480 (N_13480,N_13345,N_13305);
xor U13481 (N_13481,N_13396,N_13366);
nand U13482 (N_13482,N_13348,N_13235);
nor U13483 (N_13483,N_13230,N_13231);
nor U13484 (N_13484,N_13399,N_13351);
nor U13485 (N_13485,N_13215,N_13350);
and U13486 (N_13486,N_13227,N_13330);
nand U13487 (N_13487,N_13204,N_13202);
nor U13488 (N_13488,N_13280,N_13257);
and U13489 (N_13489,N_13207,N_13380);
xor U13490 (N_13490,N_13308,N_13241);
nand U13491 (N_13491,N_13333,N_13275);
or U13492 (N_13492,N_13262,N_13390);
or U13493 (N_13493,N_13339,N_13355);
nor U13494 (N_13494,N_13388,N_13367);
and U13495 (N_13495,N_13343,N_13306);
and U13496 (N_13496,N_13378,N_13387);
nor U13497 (N_13497,N_13212,N_13211);
and U13498 (N_13498,N_13368,N_13247);
and U13499 (N_13499,N_13370,N_13214);
or U13500 (N_13500,N_13353,N_13200);
and U13501 (N_13501,N_13276,N_13301);
or U13502 (N_13502,N_13252,N_13359);
nor U13503 (N_13503,N_13303,N_13360);
or U13504 (N_13504,N_13328,N_13309);
xnor U13505 (N_13505,N_13273,N_13395);
or U13506 (N_13506,N_13324,N_13230);
nor U13507 (N_13507,N_13235,N_13296);
and U13508 (N_13508,N_13321,N_13390);
nor U13509 (N_13509,N_13372,N_13301);
nand U13510 (N_13510,N_13322,N_13347);
nor U13511 (N_13511,N_13377,N_13340);
nand U13512 (N_13512,N_13224,N_13311);
and U13513 (N_13513,N_13257,N_13221);
nand U13514 (N_13514,N_13223,N_13265);
nor U13515 (N_13515,N_13256,N_13350);
or U13516 (N_13516,N_13221,N_13247);
or U13517 (N_13517,N_13249,N_13229);
nand U13518 (N_13518,N_13270,N_13241);
nand U13519 (N_13519,N_13294,N_13339);
and U13520 (N_13520,N_13328,N_13344);
or U13521 (N_13521,N_13388,N_13257);
nor U13522 (N_13522,N_13225,N_13393);
nand U13523 (N_13523,N_13346,N_13326);
and U13524 (N_13524,N_13278,N_13279);
and U13525 (N_13525,N_13226,N_13207);
nor U13526 (N_13526,N_13284,N_13202);
and U13527 (N_13527,N_13290,N_13277);
nand U13528 (N_13528,N_13387,N_13245);
or U13529 (N_13529,N_13247,N_13366);
nand U13530 (N_13530,N_13379,N_13345);
or U13531 (N_13531,N_13303,N_13335);
or U13532 (N_13532,N_13362,N_13214);
xor U13533 (N_13533,N_13370,N_13255);
nand U13534 (N_13534,N_13305,N_13332);
xor U13535 (N_13535,N_13365,N_13356);
or U13536 (N_13536,N_13365,N_13236);
nand U13537 (N_13537,N_13328,N_13336);
nand U13538 (N_13538,N_13377,N_13273);
nand U13539 (N_13539,N_13341,N_13287);
nand U13540 (N_13540,N_13337,N_13361);
nand U13541 (N_13541,N_13204,N_13365);
nand U13542 (N_13542,N_13230,N_13248);
and U13543 (N_13543,N_13259,N_13273);
nand U13544 (N_13544,N_13326,N_13347);
nor U13545 (N_13545,N_13355,N_13315);
or U13546 (N_13546,N_13226,N_13366);
and U13547 (N_13547,N_13346,N_13267);
or U13548 (N_13548,N_13226,N_13371);
and U13549 (N_13549,N_13200,N_13351);
nor U13550 (N_13550,N_13346,N_13300);
nand U13551 (N_13551,N_13264,N_13213);
nor U13552 (N_13552,N_13346,N_13274);
nand U13553 (N_13553,N_13238,N_13303);
xnor U13554 (N_13554,N_13348,N_13249);
nand U13555 (N_13555,N_13248,N_13226);
nor U13556 (N_13556,N_13349,N_13309);
nand U13557 (N_13557,N_13226,N_13317);
or U13558 (N_13558,N_13329,N_13281);
nand U13559 (N_13559,N_13303,N_13229);
xor U13560 (N_13560,N_13294,N_13269);
and U13561 (N_13561,N_13324,N_13316);
nand U13562 (N_13562,N_13325,N_13214);
and U13563 (N_13563,N_13397,N_13206);
and U13564 (N_13564,N_13283,N_13391);
nand U13565 (N_13565,N_13228,N_13265);
nand U13566 (N_13566,N_13260,N_13293);
nor U13567 (N_13567,N_13273,N_13217);
or U13568 (N_13568,N_13376,N_13273);
and U13569 (N_13569,N_13241,N_13348);
nor U13570 (N_13570,N_13367,N_13244);
nor U13571 (N_13571,N_13328,N_13233);
nand U13572 (N_13572,N_13213,N_13383);
and U13573 (N_13573,N_13268,N_13323);
nand U13574 (N_13574,N_13269,N_13327);
nor U13575 (N_13575,N_13328,N_13341);
and U13576 (N_13576,N_13248,N_13277);
or U13577 (N_13577,N_13354,N_13265);
or U13578 (N_13578,N_13362,N_13220);
nand U13579 (N_13579,N_13314,N_13393);
or U13580 (N_13580,N_13361,N_13353);
nand U13581 (N_13581,N_13316,N_13397);
or U13582 (N_13582,N_13214,N_13202);
nor U13583 (N_13583,N_13208,N_13330);
nand U13584 (N_13584,N_13328,N_13277);
and U13585 (N_13585,N_13253,N_13361);
or U13586 (N_13586,N_13230,N_13322);
nand U13587 (N_13587,N_13224,N_13201);
or U13588 (N_13588,N_13218,N_13368);
and U13589 (N_13589,N_13340,N_13296);
or U13590 (N_13590,N_13351,N_13233);
or U13591 (N_13591,N_13221,N_13241);
or U13592 (N_13592,N_13356,N_13388);
nor U13593 (N_13593,N_13237,N_13267);
and U13594 (N_13594,N_13298,N_13335);
or U13595 (N_13595,N_13214,N_13232);
nand U13596 (N_13596,N_13354,N_13244);
or U13597 (N_13597,N_13255,N_13395);
and U13598 (N_13598,N_13391,N_13304);
or U13599 (N_13599,N_13345,N_13351);
and U13600 (N_13600,N_13410,N_13580);
and U13601 (N_13601,N_13549,N_13500);
or U13602 (N_13602,N_13510,N_13586);
and U13603 (N_13603,N_13540,N_13467);
nand U13604 (N_13604,N_13502,N_13424);
nor U13605 (N_13605,N_13523,N_13584);
or U13606 (N_13606,N_13558,N_13568);
or U13607 (N_13607,N_13536,N_13539);
nor U13608 (N_13608,N_13454,N_13594);
xnor U13609 (N_13609,N_13447,N_13453);
and U13610 (N_13610,N_13517,N_13498);
nand U13611 (N_13611,N_13521,N_13529);
or U13612 (N_13612,N_13463,N_13570);
or U13613 (N_13613,N_13501,N_13435);
nor U13614 (N_13614,N_13417,N_13518);
nand U13615 (N_13615,N_13461,N_13491);
nor U13616 (N_13616,N_13566,N_13581);
nand U13617 (N_13617,N_13579,N_13413);
or U13618 (N_13618,N_13489,N_13555);
nor U13619 (N_13619,N_13451,N_13483);
and U13620 (N_13620,N_13543,N_13565);
or U13621 (N_13621,N_13578,N_13478);
nand U13622 (N_13622,N_13577,N_13462);
nor U13623 (N_13623,N_13468,N_13469);
nand U13624 (N_13624,N_13403,N_13457);
nand U13625 (N_13625,N_13430,N_13431);
and U13626 (N_13626,N_13547,N_13401);
nor U13627 (N_13627,N_13575,N_13573);
and U13628 (N_13628,N_13554,N_13438);
nor U13629 (N_13629,N_13595,N_13567);
xnor U13630 (N_13630,N_13422,N_13522);
nor U13631 (N_13631,N_13509,N_13599);
and U13632 (N_13632,N_13545,N_13429);
nor U13633 (N_13633,N_13512,N_13443);
nor U13634 (N_13634,N_13433,N_13464);
or U13635 (N_13635,N_13414,N_13562);
nand U13636 (N_13636,N_13470,N_13556);
and U13637 (N_13637,N_13592,N_13436);
nor U13638 (N_13638,N_13564,N_13425);
and U13639 (N_13639,N_13471,N_13546);
nand U13640 (N_13640,N_13484,N_13513);
or U13641 (N_13641,N_13588,N_13511);
nand U13642 (N_13642,N_13458,N_13475);
or U13643 (N_13643,N_13412,N_13585);
nand U13644 (N_13644,N_13507,N_13526);
nor U13645 (N_13645,N_13550,N_13520);
nand U13646 (N_13646,N_13593,N_13452);
or U13647 (N_13647,N_13477,N_13466);
nand U13648 (N_13648,N_13418,N_13450);
and U13649 (N_13649,N_13559,N_13419);
and U13650 (N_13650,N_13537,N_13408);
and U13651 (N_13651,N_13428,N_13449);
or U13652 (N_13652,N_13538,N_13440);
or U13653 (N_13653,N_13508,N_13544);
and U13654 (N_13654,N_13404,N_13542);
nor U13655 (N_13655,N_13494,N_13527);
nor U13656 (N_13656,N_13590,N_13506);
nand U13657 (N_13657,N_13474,N_13492);
nor U13658 (N_13658,N_13446,N_13548);
nand U13659 (N_13659,N_13591,N_13530);
nor U13660 (N_13660,N_13488,N_13514);
nor U13661 (N_13661,N_13407,N_13426);
nand U13662 (N_13662,N_13456,N_13485);
nand U13663 (N_13663,N_13486,N_13533);
nor U13664 (N_13664,N_13532,N_13515);
and U13665 (N_13665,N_13531,N_13441);
nand U13666 (N_13666,N_13445,N_13495);
nand U13667 (N_13667,N_13434,N_13437);
or U13668 (N_13668,N_13561,N_13493);
or U13669 (N_13669,N_13504,N_13465);
and U13670 (N_13670,N_13596,N_13420);
nor U13671 (N_13671,N_13423,N_13519);
nor U13672 (N_13672,N_13598,N_13442);
nand U13673 (N_13673,N_13490,N_13439);
nand U13674 (N_13674,N_13560,N_13503);
nand U13675 (N_13675,N_13473,N_13482);
or U13676 (N_13676,N_13553,N_13541);
or U13677 (N_13677,N_13444,N_13405);
nor U13678 (N_13678,N_13597,N_13576);
nand U13679 (N_13679,N_13557,N_13582);
nor U13680 (N_13680,N_13416,N_13497);
or U13681 (N_13681,N_13402,N_13583);
nor U13682 (N_13682,N_13552,N_13551);
nor U13683 (N_13683,N_13460,N_13528);
nand U13684 (N_13684,N_13487,N_13459);
or U13685 (N_13685,N_13448,N_13505);
nor U13686 (N_13686,N_13496,N_13525);
nand U13687 (N_13687,N_13535,N_13406);
nand U13688 (N_13688,N_13589,N_13571);
nand U13689 (N_13689,N_13455,N_13499);
nand U13690 (N_13690,N_13587,N_13476);
and U13691 (N_13691,N_13479,N_13563);
nor U13692 (N_13692,N_13572,N_13574);
and U13693 (N_13693,N_13432,N_13516);
nor U13694 (N_13694,N_13411,N_13481);
and U13695 (N_13695,N_13472,N_13524);
and U13696 (N_13696,N_13534,N_13569);
nand U13697 (N_13697,N_13480,N_13400);
nand U13698 (N_13698,N_13427,N_13409);
and U13699 (N_13699,N_13421,N_13415);
and U13700 (N_13700,N_13548,N_13524);
nand U13701 (N_13701,N_13531,N_13413);
or U13702 (N_13702,N_13451,N_13419);
and U13703 (N_13703,N_13517,N_13519);
and U13704 (N_13704,N_13586,N_13530);
and U13705 (N_13705,N_13404,N_13532);
and U13706 (N_13706,N_13430,N_13524);
nor U13707 (N_13707,N_13516,N_13400);
nor U13708 (N_13708,N_13529,N_13415);
and U13709 (N_13709,N_13520,N_13435);
nand U13710 (N_13710,N_13406,N_13581);
nand U13711 (N_13711,N_13536,N_13476);
or U13712 (N_13712,N_13574,N_13583);
nor U13713 (N_13713,N_13505,N_13517);
nand U13714 (N_13714,N_13491,N_13462);
nor U13715 (N_13715,N_13404,N_13423);
and U13716 (N_13716,N_13426,N_13529);
and U13717 (N_13717,N_13572,N_13494);
and U13718 (N_13718,N_13459,N_13476);
nand U13719 (N_13719,N_13504,N_13502);
nand U13720 (N_13720,N_13475,N_13416);
and U13721 (N_13721,N_13484,N_13517);
nand U13722 (N_13722,N_13560,N_13492);
and U13723 (N_13723,N_13572,N_13544);
or U13724 (N_13724,N_13500,N_13597);
and U13725 (N_13725,N_13437,N_13518);
nand U13726 (N_13726,N_13445,N_13598);
nand U13727 (N_13727,N_13562,N_13546);
and U13728 (N_13728,N_13405,N_13509);
nor U13729 (N_13729,N_13425,N_13419);
nor U13730 (N_13730,N_13474,N_13527);
or U13731 (N_13731,N_13439,N_13569);
and U13732 (N_13732,N_13454,N_13470);
nor U13733 (N_13733,N_13533,N_13443);
xnor U13734 (N_13734,N_13410,N_13417);
nand U13735 (N_13735,N_13479,N_13532);
nand U13736 (N_13736,N_13489,N_13511);
nor U13737 (N_13737,N_13582,N_13427);
nand U13738 (N_13738,N_13511,N_13540);
and U13739 (N_13739,N_13441,N_13494);
nor U13740 (N_13740,N_13498,N_13526);
or U13741 (N_13741,N_13413,N_13562);
xnor U13742 (N_13742,N_13400,N_13556);
and U13743 (N_13743,N_13564,N_13467);
and U13744 (N_13744,N_13576,N_13524);
and U13745 (N_13745,N_13489,N_13563);
nand U13746 (N_13746,N_13421,N_13533);
and U13747 (N_13747,N_13530,N_13412);
or U13748 (N_13748,N_13448,N_13512);
or U13749 (N_13749,N_13498,N_13519);
nor U13750 (N_13750,N_13493,N_13550);
nor U13751 (N_13751,N_13429,N_13401);
nor U13752 (N_13752,N_13407,N_13575);
and U13753 (N_13753,N_13578,N_13424);
and U13754 (N_13754,N_13492,N_13592);
and U13755 (N_13755,N_13537,N_13500);
and U13756 (N_13756,N_13548,N_13552);
and U13757 (N_13757,N_13558,N_13436);
nor U13758 (N_13758,N_13570,N_13583);
or U13759 (N_13759,N_13556,N_13482);
and U13760 (N_13760,N_13446,N_13549);
nor U13761 (N_13761,N_13441,N_13416);
nand U13762 (N_13762,N_13449,N_13519);
and U13763 (N_13763,N_13467,N_13476);
nor U13764 (N_13764,N_13487,N_13479);
or U13765 (N_13765,N_13531,N_13426);
nand U13766 (N_13766,N_13515,N_13441);
nor U13767 (N_13767,N_13463,N_13423);
and U13768 (N_13768,N_13537,N_13481);
nand U13769 (N_13769,N_13554,N_13584);
nor U13770 (N_13770,N_13558,N_13438);
nand U13771 (N_13771,N_13449,N_13573);
nand U13772 (N_13772,N_13404,N_13449);
and U13773 (N_13773,N_13524,N_13404);
or U13774 (N_13774,N_13579,N_13483);
nor U13775 (N_13775,N_13437,N_13590);
and U13776 (N_13776,N_13521,N_13438);
or U13777 (N_13777,N_13556,N_13451);
and U13778 (N_13778,N_13481,N_13534);
nand U13779 (N_13779,N_13451,N_13586);
and U13780 (N_13780,N_13560,N_13522);
nor U13781 (N_13781,N_13497,N_13400);
nor U13782 (N_13782,N_13474,N_13595);
or U13783 (N_13783,N_13437,N_13482);
or U13784 (N_13784,N_13403,N_13452);
nor U13785 (N_13785,N_13456,N_13591);
and U13786 (N_13786,N_13568,N_13403);
or U13787 (N_13787,N_13434,N_13421);
nor U13788 (N_13788,N_13465,N_13457);
and U13789 (N_13789,N_13468,N_13522);
nand U13790 (N_13790,N_13539,N_13532);
and U13791 (N_13791,N_13450,N_13511);
and U13792 (N_13792,N_13492,N_13527);
and U13793 (N_13793,N_13580,N_13449);
and U13794 (N_13794,N_13452,N_13462);
nor U13795 (N_13795,N_13514,N_13417);
nand U13796 (N_13796,N_13545,N_13509);
nor U13797 (N_13797,N_13584,N_13405);
nor U13798 (N_13798,N_13596,N_13489);
nor U13799 (N_13799,N_13474,N_13475);
nor U13800 (N_13800,N_13764,N_13660);
or U13801 (N_13801,N_13752,N_13699);
nand U13802 (N_13802,N_13748,N_13630);
nand U13803 (N_13803,N_13626,N_13682);
and U13804 (N_13804,N_13724,N_13762);
or U13805 (N_13805,N_13749,N_13687);
nand U13806 (N_13806,N_13732,N_13665);
or U13807 (N_13807,N_13627,N_13781);
and U13808 (N_13808,N_13712,N_13641);
nor U13809 (N_13809,N_13685,N_13717);
nand U13810 (N_13810,N_13667,N_13628);
and U13811 (N_13811,N_13737,N_13734);
nand U13812 (N_13812,N_13671,N_13694);
nand U13813 (N_13813,N_13600,N_13650);
and U13814 (N_13814,N_13690,N_13646);
and U13815 (N_13815,N_13735,N_13775);
or U13816 (N_13816,N_13779,N_13635);
nand U13817 (N_13817,N_13746,N_13788);
nor U13818 (N_13818,N_13686,N_13701);
nor U13819 (N_13819,N_13725,N_13758);
nand U13820 (N_13820,N_13745,N_13778);
or U13821 (N_13821,N_13772,N_13692);
nor U13822 (N_13822,N_13704,N_13607);
nor U13823 (N_13823,N_13615,N_13765);
nand U13824 (N_13824,N_13611,N_13657);
nor U13825 (N_13825,N_13661,N_13766);
nor U13826 (N_13826,N_13640,N_13643);
nand U13827 (N_13827,N_13654,N_13681);
nand U13828 (N_13828,N_13776,N_13777);
nor U13829 (N_13829,N_13696,N_13618);
or U13830 (N_13830,N_13614,N_13794);
or U13831 (N_13831,N_13786,N_13689);
nand U13832 (N_13832,N_13683,N_13706);
nand U13833 (N_13833,N_13715,N_13609);
nor U13834 (N_13834,N_13602,N_13638);
nand U13835 (N_13835,N_13739,N_13782);
or U13836 (N_13836,N_13798,N_13670);
or U13837 (N_13837,N_13768,N_13714);
nor U13838 (N_13838,N_13727,N_13708);
and U13839 (N_13839,N_13709,N_13723);
nor U13840 (N_13840,N_13639,N_13738);
xnor U13841 (N_13841,N_13610,N_13722);
nand U13842 (N_13842,N_13617,N_13783);
nor U13843 (N_13843,N_13744,N_13637);
or U13844 (N_13844,N_13642,N_13678);
nand U13845 (N_13845,N_13759,N_13625);
nand U13846 (N_13846,N_13655,N_13733);
nor U13847 (N_13847,N_13698,N_13791);
and U13848 (N_13848,N_13726,N_13785);
nor U13849 (N_13849,N_13741,N_13713);
xnor U13850 (N_13850,N_13619,N_13750);
and U13851 (N_13851,N_13796,N_13623);
nand U13852 (N_13852,N_13774,N_13771);
or U13853 (N_13853,N_13649,N_13684);
and U13854 (N_13854,N_13621,N_13616);
or U13855 (N_13855,N_13674,N_13658);
xor U13856 (N_13856,N_13664,N_13624);
nor U13857 (N_13857,N_13608,N_13760);
nand U13858 (N_13858,N_13730,N_13799);
nand U13859 (N_13859,N_13718,N_13677);
xnor U13860 (N_13860,N_13620,N_13672);
nor U13861 (N_13861,N_13691,N_13613);
nor U13862 (N_13862,N_13731,N_13755);
nor U13863 (N_13863,N_13612,N_13663);
nor U13864 (N_13864,N_13675,N_13622);
nor U13865 (N_13865,N_13688,N_13652);
nand U13866 (N_13866,N_13700,N_13740);
nor U13867 (N_13867,N_13716,N_13710);
nor U13868 (N_13868,N_13656,N_13721);
nor U13869 (N_13869,N_13728,N_13659);
nand U13870 (N_13870,N_13797,N_13756);
nor U13871 (N_13871,N_13780,N_13648);
or U13872 (N_13872,N_13754,N_13662);
nor U13873 (N_13873,N_13753,N_13720);
nand U13874 (N_13874,N_13742,N_13784);
and U13875 (N_13875,N_13601,N_13787);
nor U13876 (N_13876,N_13633,N_13634);
nand U13877 (N_13877,N_13651,N_13673);
and U13878 (N_13878,N_13680,N_13631);
and U13879 (N_13879,N_13757,N_13793);
nor U13880 (N_13880,N_13763,N_13789);
or U13881 (N_13881,N_13604,N_13603);
nand U13882 (N_13882,N_13773,N_13795);
or U13883 (N_13883,N_13751,N_13743);
or U13884 (N_13884,N_13697,N_13605);
nor U13885 (N_13885,N_13747,N_13705);
and U13886 (N_13886,N_13790,N_13669);
nand U13887 (N_13887,N_13676,N_13792);
or U13888 (N_13888,N_13702,N_13606);
nor U13889 (N_13889,N_13679,N_13644);
or U13890 (N_13890,N_13769,N_13647);
and U13891 (N_13891,N_13729,N_13767);
and U13892 (N_13892,N_13695,N_13703);
nand U13893 (N_13893,N_13693,N_13636);
and U13894 (N_13894,N_13666,N_13719);
or U13895 (N_13895,N_13668,N_13645);
nand U13896 (N_13896,N_13711,N_13761);
or U13897 (N_13897,N_13629,N_13707);
nand U13898 (N_13898,N_13653,N_13632);
nand U13899 (N_13899,N_13736,N_13770);
nor U13900 (N_13900,N_13649,N_13693);
or U13901 (N_13901,N_13768,N_13658);
nor U13902 (N_13902,N_13705,N_13778);
nand U13903 (N_13903,N_13687,N_13658);
and U13904 (N_13904,N_13719,N_13662);
or U13905 (N_13905,N_13627,N_13651);
nand U13906 (N_13906,N_13707,N_13678);
and U13907 (N_13907,N_13798,N_13646);
or U13908 (N_13908,N_13782,N_13733);
or U13909 (N_13909,N_13797,N_13785);
or U13910 (N_13910,N_13706,N_13781);
xnor U13911 (N_13911,N_13761,N_13709);
nand U13912 (N_13912,N_13661,N_13730);
and U13913 (N_13913,N_13634,N_13672);
and U13914 (N_13914,N_13735,N_13601);
and U13915 (N_13915,N_13639,N_13654);
nor U13916 (N_13916,N_13738,N_13689);
and U13917 (N_13917,N_13707,N_13762);
nor U13918 (N_13918,N_13742,N_13780);
nor U13919 (N_13919,N_13782,N_13735);
nand U13920 (N_13920,N_13754,N_13674);
and U13921 (N_13921,N_13653,N_13772);
nand U13922 (N_13922,N_13602,N_13729);
and U13923 (N_13923,N_13746,N_13764);
or U13924 (N_13924,N_13673,N_13723);
nand U13925 (N_13925,N_13787,N_13655);
nor U13926 (N_13926,N_13722,N_13656);
nand U13927 (N_13927,N_13605,N_13613);
and U13928 (N_13928,N_13753,N_13716);
nand U13929 (N_13929,N_13715,N_13633);
nand U13930 (N_13930,N_13603,N_13631);
and U13931 (N_13931,N_13779,N_13657);
nor U13932 (N_13932,N_13616,N_13635);
and U13933 (N_13933,N_13773,N_13631);
nor U13934 (N_13934,N_13792,N_13755);
nor U13935 (N_13935,N_13604,N_13627);
nand U13936 (N_13936,N_13624,N_13768);
and U13937 (N_13937,N_13709,N_13615);
or U13938 (N_13938,N_13608,N_13601);
or U13939 (N_13939,N_13722,N_13663);
and U13940 (N_13940,N_13698,N_13652);
nand U13941 (N_13941,N_13736,N_13710);
nor U13942 (N_13942,N_13736,N_13684);
or U13943 (N_13943,N_13666,N_13773);
and U13944 (N_13944,N_13690,N_13714);
xnor U13945 (N_13945,N_13704,N_13771);
and U13946 (N_13946,N_13635,N_13777);
nand U13947 (N_13947,N_13754,N_13701);
nor U13948 (N_13948,N_13741,N_13600);
and U13949 (N_13949,N_13714,N_13695);
nor U13950 (N_13950,N_13676,N_13701);
nor U13951 (N_13951,N_13796,N_13787);
nor U13952 (N_13952,N_13678,N_13784);
nor U13953 (N_13953,N_13602,N_13634);
and U13954 (N_13954,N_13725,N_13717);
nor U13955 (N_13955,N_13636,N_13795);
and U13956 (N_13956,N_13620,N_13651);
nor U13957 (N_13957,N_13737,N_13703);
nor U13958 (N_13958,N_13739,N_13696);
nor U13959 (N_13959,N_13692,N_13779);
or U13960 (N_13960,N_13709,N_13685);
and U13961 (N_13961,N_13729,N_13645);
nor U13962 (N_13962,N_13678,N_13789);
and U13963 (N_13963,N_13725,N_13663);
nor U13964 (N_13964,N_13627,N_13792);
or U13965 (N_13965,N_13646,N_13778);
nor U13966 (N_13966,N_13692,N_13778);
or U13967 (N_13967,N_13799,N_13766);
nor U13968 (N_13968,N_13730,N_13670);
or U13969 (N_13969,N_13643,N_13668);
nand U13970 (N_13970,N_13645,N_13763);
or U13971 (N_13971,N_13710,N_13720);
nor U13972 (N_13972,N_13778,N_13731);
or U13973 (N_13973,N_13672,N_13752);
nor U13974 (N_13974,N_13630,N_13742);
and U13975 (N_13975,N_13719,N_13612);
or U13976 (N_13976,N_13712,N_13606);
and U13977 (N_13977,N_13722,N_13619);
or U13978 (N_13978,N_13725,N_13658);
and U13979 (N_13979,N_13732,N_13710);
nor U13980 (N_13980,N_13783,N_13712);
or U13981 (N_13981,N_13606,N_13771);
and U13982 (N_13982,N_13661,N_13639);
nand U13983 (N_13983,N_13723,N_13698);
and U13984 (N_13984,N_13662,N_13749);
nand U13985 (N_13985,N_13774,N_13617);
nand U13986 (N_13986,N_13747,N_13760);
or U13987 (N_13987,N_13711,N_13734);
nor U13988 (N_13988,N_13649,N_13695);
and U13989 (N_13989,N_13603,N_13777);
or U13990 (N_13990,N_13621,N_13738);
and U13991 (N_13991,N_13687,N_13759);
nand U13992 (N_13992,N_13695,N_13788);
and U13993 (N_13993,N_13693,N_13718);
nor U13994 (N_13994,N_13740,N_13600);
and U13995 (N_13995,N_13676,N_13770);
and U13996 (N_13996,N_13777,N_13770);
or U13997 (N_13997,N_13731,N_13743);
or U13998 (N_13998,N_13676,N_13716);
nand U13999 (N_13999,N_13712,N_13781);
and U14000 (N_14000,N_13889,N_13844);
or U14001 (N_14001,N_13820,N_13807);
nor U14002 (N_14002,N_13813,N_13929);
nor U14003 (N_14003,N_13890,N_13946);
nand U14004 (N_14004,N_13804,N_13836);
xnor U14005 (N_14005,N_13920,N_13816);
nor U14006 (N_14006,N_13870,N_13909);
nand U14007 (N_14007,N_13961,N_13885);
nand U14008 (N_14008,N_13990,N_13956);
or U14009 (N_14009,N_13966,N_13965);
and U14010 (N_14010,N_13864,N_13896);
nand U14011 (N_14011,N_13975,N_13922);
and U14012 (N_14012,N_13959,N_13850);
nor U14013 (N_14013,N_13888,N_13993);
or U14014 (N_14014,N_13949,N_13884);
nand U14015 (N_14015,N_13863,N_13833);
nor U14016 (N_14016,N_13845,N_13998);
nor U14017 (N_14017,N_13932,N_13962);
nor U14018 (N_14018,N_13916,N_13950);
or U14019 (N_14019,N_13802,N_13840);
nor U14020 (N_14020,N_13823,N_13847);
nand U14021 (N_14021,N_13900,N_13851);
nor U14022 (N_14022,N_13968,N_13999);
or U14023 (N_14023,N_13967,N_13817);
and U14024 (N_14024,N_13919,N_13924);
or U14025 (N_14025,N_13992,N_13879);
nand U14026 (N_14026,N_13953,N_13986);
nor U14027 (N_14027,N_13877,N_13859);
nand U14028 (N_14028,N_13891,N_13837);
nand U14029 (N_14029,N_13893,N_13939);
xnor U14030 (N_14030,N_13857,N_13810);
nor U14031 (N_14031,N_13908,N_13855);
nand U14032 (N_14032,N_13971,N_13963);
and U14033 (N_14033,N_13806,N_13865);
nor U14034 (N_14034,N_13812,N_13832);
nor U14035 (N_14035,N_13991,N_13871);
nor U14036 (N_14036,N_13977,N_13936);
nand U14037 (N_14037,N_13982,N_13839);
nand U14038 (N_14038,N_13997,N_13876);
and U14039 (N_14039,N_13921,N_13996);
or U14040 (N_14040,N_13853,N_13869);
or U14041 (N_14041,N_13803,N_13886);
nor U14042 (N_14042,N_13834,N_13866);
nand U14043 (N_14043,N_13994,N_13911);
nor U14044 (N_14044,N_13913,N_13948);
nand U14045 (N_14045,N_13987,N_13973);
nand U14046 (N_14046,N_13821,N_13860);
nand U14047 (N_14047,N_13960,N_13905);
nor U14048 (N_14048,N_13856,N_13852);
or U14049 (N_14049,N_13835,N_13849);
nand U14050 (N_14050,N_13831,N_13874);
nand U14051 (N_14051,N_13944,N_13880);
nor U14052 (N_14052,N_13969,N_13901);
and U14053 (N_14053,N_13827,N_13898);
or U14054 (N_14054,N_13981,N_13897);
nor U14055 (N_14055,N_13941,N_13964);
nor U14056 (N_14056,N_13976,N_13927);
and U14057 (N_14057,N_13995,N_13972);
nand U14058 (N_14058,N_13811,N_13970);
and U14059 (N_14059,N_13930,N_13979);
nor U14060 (N_14060,N_13808,N_13826);
or U14061 (N_14061,N_13819,N_13825);
and U14062 (N_14062,N_13828,N_13937);
or U14063 (N_14063,N_13923,N_13934);
and U14064 (N_14064,N_13824,N_13952);
nand U14065 (N_14065,N_13988,N_13872);
or U14066 (N_14066,N_13894,N_13938);
xor U14067 (N_14067,N_13903,N_13892);
or U14068 (N_14068,N_13805,N_13830);
nand U14069 (N_14069,N_13935,N_13809);
nand U14070 (N_14070,N_13822,N_13984);
nand U14071 (N_14071,N_13926,N_13883);
or U14072 (N_14072,N_13904,N_13842);
or U14073 (N_14073,N_13933,N_13887);
nor U14074 (N_14074,N_13868,N_13931);
or U14075 (N_14075,N_13875,N_13917);
nand U14076 (N_14076,N_13951,N_13943);
nand U14077 (N_14077,N_13862,N_13907);
nor U14078 (N_14078,N_13940,N_13985);
nand U14079 (N_14079,N_13846,N_13801);
or U14080 (N_14080,N_13899,N_13947);
or U14081 (N_14081,N_13910,N_13848);
and U14082 (N_14082,N_13914,N_13980);
and U14083 (N_14083,N_13925,N_13912);
or U14084 (N_14084,N_13928,N_13878);
or U14085 (N_14085,N_13882,N_13818);
and U14086 (N_14086,N_13814,N_13902);
and U14087 (N_14087,N_13983,N_13854);
nand U14088 (N_14088,N_13942,N_13867);
and U14089 (N_14089,N_13873,N_13918);
nor U14090 (N_14090,N_13957,N_13974);
xor U14091 (N_14091,N_13955,N_13843);
nand U14092 (N_14092,N_13841,N_13945);
and U14093 (N_14093,N_13881,N_13954);
or U14094 (N_14094,N_13815,N_13989);
or U14095 (N_14095,N_13861,N_13829);
nor U14096 (N_14096,N_13915,N_13906);
nor U14097 (N_14097,N_13800,N_13958);
or U14098 (N_14098,N_13858,N_13838);
nand U14099 (N_14099,N_13895,N_13978);
or U14100 (N_14100,N_13813,N_13969);
and U14101 (N_14101,N_13890,N_13823);
nor U14102 (N_14102,N_13955,N_13890);
nand U14103 (N_14103,N_13920,N_13878);
nand U14104 (N_14104,N_13993,N_13900);
or U14105 (N_14105,N_13831,N_13811);
nor U14106 (N_14106,N_13889,N_13900);
and U14107 (N_14107,N_13911,N_13863);
nand U14108 (N_14108,N_13983,N_13801);
and U14109 (N_14109,N_13825,N_13921);
nand U14110 (N_14110,N_13880,N_13987);
or U14111 (N_14111,N_13918,N_13946);
nor U14112 (N_14112,N_13822,N_13957);
and U14113 (N_14113,N_13844,N_13803);
or U14114 (N_14114,N_13834,N_13858);
and U14115 (N_14115,N_13978,N_13897);
nand U14116 (N_14116,N_13885,N_13903);
nor U14117 (N_14117,N_13988,N_13890);
or U14118 (N_14118,N_13901,N_13935);
or U14119 (N_14119,N_13820,N_13877);
nor U14120 (N_14120,N_13823,N_13944);
or U14121 (N_14121,N_13982,N_13824);
nand U14122 (N_14122,N_13972,N_13832);
nand U14123 (N_14123,N_13892,N_13850);
nand U14124 (N_14124,N_13965,N_13956);
and U14125 (N_14125,N_13967,N_13920);
nor U14126 (N_14126,N_13807,N_13812);
xnor U14127 (N_14127,N_13937,N_13843);
or U14128 (N_14128,N_13833,N_13957);
nor U14129 (N_14129,N_13976,N_13986);
nand U14130 (N_14130,N_13958,N_13879);
nor U14131 (N_14131,N_13849,N_13971);
or U14132 (N_14132,N_13967,N_13803);
and U14133 (N_14133,N_13814,N_13947);
or U14134 (N_14134,N_13952,N_13891);
nor U14135 (N_14135,N_13913,N_13838);
xnor U14136 (N_14136,N_13808,N_13841);
nor U14137 (N_14137,N_13960,N_13938);
xnor U14138 (N_14138,N_13887,N_13836);
or U14139 (N_14139,N_13949,N_13885);
nor U14140 (N_14140,N_13908,N_13955);
nand U14141 (N_14141,N_13806,N_13867);
nor U14142 (N_14142,N_13861,N_13922);
nand U14143 (N_14143,N_13943,N_13927);
or U14144 (N_14144,N_13957,N_13875);
and U14145 (N_14145,N_13974,N_13987);
and U14146 (N_14146,N_13863,N_13922);
or U14147 (N_14147,N_13955,N_13827);
or U14148 (N_14148,N_13890,N_13900);
xor U14149 (N_14149,N_13824,N_13830);
nand U14150 (N_14150,N_13845,N_13944);
or U14151 (N_14151,N_13840,N_13869);
nand U14152 (N_14152,N_13854,N_13853);
nand U14153 (N_14153,N_13864,N_13874);
and U14154 (N_14154,N_13911,N_13917);
and U14155 (N_14155,N_13802,N_13907);
nand U14156 (N_14156,N_13805,N_13923);
nand U14157 (N_14157,N_13805,N_13823);
nand U14158 (N_14158,N_13944,N_13930);
nor U14159 (N_14159,N_13844,N_13906);
or U14160 (N_14160,N_13818,N_13888);
or U14161 (N_14161,N_13961,N_13865);
and U14162 (N_14162,N_13879,N_13856);
nand U14163 (N_14163,N_13942,N_13892);
and U14164 (N_14164,N_13863,N_13995);
or U14165 (N_14165,N_13993,N_13940);
nor U14166 (N_14166,N_13983,N_13873);
nor U14167 (N_14167,N_13899,N_13916);
nor U14168 (N_14168,N_13891,N_13836);
or U14169 (N_14169,N_13973,N_13931);
nand U14170 (N_14170,N_13971,N_13894);
nor U14171 (N_14171,N_13924,N_13965);
or U14172 (N_14172,N_13884,N_13960);
nand U14173 (N_14173,N_13876,N_13862);
nand U14174 (N_14174,N_13942,N_13930);
and U14175 (N_14175,N_13875,N_13954);
nand U14176 (N_14176,N_13832,N_13866);
and U14177 (N_14177,N_13825,N_13901);
and U14178 (N_14178,N_13954,N_13963);
nand U14179 (N_14179,N_13996,N_13809);
nor U14180 (N_14180,N_13921,N_13873);
xor U14181 (N_14181,N_13830,N_13932);
or U14182 (N_14182,N_13901,N_13810);
nor U14183 (N_14183,N_13839,N_13896);
nor U14184 (N_14184,N_13861,N_13998);
nor U14185 (N_14185,N_13810,N_13872);
xnor U14186 (N_14186,N_13906,N_13917);
nor U14187 (N_14187,N_13802,N_13834);
and U14188 (N_14188,N_13958,N_13826);
or U14189 (N_14189,N_13870,N_13991);
or U14190 (N_14190,N_13842,N_13929);
or U14191 (N_14191,N_13820,N_13868);
nor U14192 (N_14192,N_13832,N_13816);
and U14193 (N_14193,N_13900,N_13843);
and U14194 (N_14194,N_13981,N_13990);
nand U14195 (N_14195,N_13889,N_13890);
nand U14196 (N_14196,N_13874,N_13840);
nor U14197 (N_14197,N_13824,N_13803);
nand U14198 (N_14198,N_13938,N_13812);
nor U14199 (N_14199,N_13822,N_13859);
or U14200 (N_14200,N_14092,N_14169);
nor U14201 (N_14201,N_14004,N_14052);
nand U14202 (N_14202,N_14174,N_14139);
nand U14203 (N_14203,N_14172,N_14003);
nand U14204 (N_14204,N_14187,N_14019);
and U14205 (N_14205,N_14170,N_14072);
nand U14206 (N_14206,N_14165,N_14021);
and U14207 (N_14207,N_14007,N_14060);
nand U14208 (N_14208,N_14142,N_14050);
and U14209 (N_14209,N_14127,N_14132);
nor U14210 (N_14210,N_14159,N_14062);
or U14211 (N_14211,N_14158,N_14084);
or U14212 (N_14212,N_14186,N_14009);
nor U14213 (N_14213,N_14001,N_14031);
nand U14214 (N_14214,N_14155,N_14051);
and U14215 (N_14215,N_14049,N_14033);
nor U14216 (N_14216,N_14077,N_14199);
or U14217 (N_14217,N_14163,N_14128);
or U14218 (N_14218,N_14067,N_14055);
nand U14219 (N_14219,N_14103,N_14089);
nor U14220 (N_14220,N_14056,N_14039);
or U14221 (N_14221,N_14016,N_14150);
nor U14222 (N_14222,N_14015,N_14063);
and U14223 (N_14223,N_14164,N_14090);
and U14224 (N_14224,N_14087,N_14102);
nand U14225 (N_14225,N_14178,N_14119);
nor U14226 (N_14226,N_14010,N_14146);
nor U14227 (N_14227,N_14101,N_14027);
and U14228 (N_14228,N_14040,N_14037);
and U14229 (N_14229,N_14195,N_14153);
nand U14230 (N_14230,N_14093,N_14097);
or U14231 (N_14231,N_14191,N_14141);
nor U14232 (N_14232,N_14036,N_14152);
and U14233 (N_14233,N_14129,N_14130);
nand U14234 (N_14234,N_14022,N_14065);
and U14235 (N_14235,N_14059,N_14176);
nand U14236 (N_14236,N_14110,N_14151);
or U14237 (N_14237,N_14184,N_14198);
nor U14238 (N_14238,N_14156,N_14014);
and U14239 (N_14239,N_14100,N_14166);
or U14240 (N_14240,N_14123,N_14053);
nor U14241 (N_14241,N_14182,N_14085);
nand U14242 (N_14242,N_14026,N_14017);
or U14243 (N_14243,N_14035,N_14098);
and U14244 (N_14244,N_14108,N_14183);
nor U14245 (N_14245,N_14185,N_14066);
and U14246 (N_14246,N_14112,N_14088);
or U14247 (N_14247,N_14121,N_14116);
and U14248 (N_14248,N_14061,N_14073);
nor U14249 (N_14249,N_14173,N_14058);
and U14250 (N_14250,N_14136,N_14011);
or U14251 (N_14251,N_14125,N_14189);
or U14252 (N_14252,N_14041,N_14030);
or U14253 (N_14253,N_14157,N_14194);
nor U14254 (N_14254,N_14042,N_14095);
nand U14255 (N_14255,N_14000,N_14024);
or U14256 (N_14256,N_14074,N_14149);
and U14257 (N_14257,N_14109,N_14181);
or U14258 (N_14258,N_14029,N_14147);
nor U14259 (N_14259,N_14079,N_14005);
nand U14260 (N_14260,N_14081,N_14020);
and U14261 (N_14261,N_14190,N_14122);
nor U14262 (N_14262,N_14076,N_14078);
nand U14263 (N_14263,N_14038,N_14161);
and U14264 (N_14264,N_14025,N_14126);
and U14265 (N_14265,N_14044,N_14143);
nor U14266 (N_14266,N_14080,N_14034);
and U14267 (N_14267,N_14032,N_14086);
or U14268 (N_14268,N_14046,N_14105);
nor U14269 (N_14269,N_14018,N_14107);
nor U14270 (N_14270,N_14138,N_14197);
or U14271 (N_14271,N_14168,N_14002);
xor U14272 (N_14272,N_14140,N_14193);
or U14273 (N_14273,N_14054,N_14012);
or U14274 (N_14274,N_14008,N_14069);
xnor U14275 (N_14275,N_14162,N_14144);
or U14276 (N_14276,N_14192,N_14048);
and U14277 (N_14277,N_14099,N_14023);
nand U14278 (N_14278,N_14045,N_14177);
and U14279 (N_14279,N_14148,N_14160);
and U14280 (N_14280,N_14013,N_14047);
or U14281 (N_14281,N_14131,N_14114);
or U14282 (N_14282,N_14064,N_14133);
nor U14283 (N_14283,N_14043,N_14124);
or U14284 (N_14284,N_14188,N_14106);
and U14285 (N_14285,N_14068,N_14145);
nor U14286 (N_14286,N_14117,N_14175);
nor U14287 (N_14287,N_14118,N_14137);
nand U14288 (N_14288,N_14115,N_14179);
nand U14289 (N_14289,N_14167,N_14071);
or U14290 (N_14290,N_14070,N_14083);
nor U14291 (N_14291,N_14111,N_14075);
or U14292 (N_14292,N_14091,N_14171);
nor U14293 (N_14293,N_14028,N_14057);
nand U14294 (N_14294,N_14082,N_14094);
nand U14295 (N_14295,N_14196,N_14006);
nand U14296 (N_14296,N_14180,N_14120);
nor U14297 (N_14297,N_14134,N_14104);
nor U14298 (N_14298,N_14096,N_14135);
and U14299 (N_14299,N_14113,N_14154);
or U14300 (N_14300,N_14030,N_14052);
nand U14301 (N_14301,N_14024,N_14007);
or U14302 (N_14302,N_14168,N_14086);
and U14303 (N_14303,N_14110,N_14041);
nor U14304 (N_14304,N_14039,N_14068);
nand U14305 (N_14305,N_14087,N_14143);
nor U14306 (N_14306,N_14183,N_14184);
or U14307 (N_14307,N_14095,N_14031);
and U14308 (N_14308,N_14064,N_14105);
nand U14309 (N_14309,N_14024,N_14094);
nand U14310 (N_14310,N_14164,N_14046);
nand U14311 (N_14311,N_14122,N_14008);
nand U14312 (N_14312,N_14151,N_14084);
nand U14313 (N_14313,N_14101,N_14064);
nor U14314 (N_14314,N_14082,N_14122);
and U14315 (N_14315,N_14190,N_14117);
or U14316 (N_14316,N_14069,N_14133);
or U14317 (N_14317,N_14025,N_14162);
and U14318 (N_14318,N_14165,N_14011);
nand U14319 (N_14319,N_14198,N_14128);
or U14320 (N_14320,N_14189,N_14115);
or U14321 (N_14321,N_14111,N_14013);
nor U14322 (N_14322,N_14045,N_14030);
and U14323 (N_14323,N_14137,N_14064);
nor U14324 (N_14324,N_14159,N_14181);
and U14325 (N_14325,N_14050,N_14185);
and U14326 (N_14326,N_14062,N_14193);
nand U14327 (N_14327,N_14182,N_14042);
nand U14328 (N_14328,N_14190,N_14076);
or U14329 (N_14329,N_14022,N_14031);
or U14330 (N_14330,N_14022,N_14140);
and U14331 (N_14331,N_14153,N_14184);
or U14332 (N_14332,N_14174,N_14156);
and U14333 (N_14333,N_14134,N_14075);
and U14334 (N_14334,N_14099,N_14112);
nor U14335 (N_14335,N_14067,N_14174);
or U14336 (N_14336,N_14112,N_14147);
nor U14337 (N_14337,N_14139,N_14199);
xnor U14338 (N_14338,N_14103,N_14157);
or U14339 (N_14339,N_14124,N_14035);
or U14340 (N_14340,N_14000,N_14044);
nand U14341 (N_14341,N_14021,N_14046);
nand U14342 (N_14342,N_14052,N_14086);
or U14343 (N_14343,N_14191,N_14180);
nor U14344 (N_14344,N_14185,N_14150);
or U14345 (N_14345,N_14199,N_14078);
nand U14346 (N_14346,N_14153,N_14155);
nor U14347 (N_14347,N_14112,N_14140);
and U14348 (N_14348,N_14119,N_14153);
and U14349 (N_14349,N_14001,N_14199);
nand U14350 (N_14350,N_14073,N_14112);
and U14351 (N_14351,N_14124,N_14123);
nor U14352 (N_14352,N_14189,N_14051);
or U14353 (N_14353,N_14173,N_14009);
or U14354 (N_14354,N_14078,N_14127);
or U14355 (N_14355,N_14105,N_14180);
and U14356 (N_14356,N_14065,N_14014);
or U14357 (N_14357,N_14128,N_14059);
nand U14358 (N_14358,N_14106,N_14103);
nand U14359 (N_14359,N_14191,N_14134);
or U14360 (N_14360,N_14049,N_14014);
nand U14361 (N_14361,N_14040,N_14168);
and U14362 (N_14362,N_14175,N_14169);
nand U14363 (N_14363,N_14141,N_14085);
or U14364 (N_14364,N_14114,N_14034);
or U14365 (N_14365,N_14115,N_14012);
nor U14366 (N_14366,N_14112,N_14153);
or U14367 (N_14367,N_14018,N_14106);
or U14368 (N_14368,N_14190,N_14002);
and U14369 (N_14369,N_14189,N_14063);
or U14370 (N_14370,N_14023,N_14195);
and U14371 (N_14371,N_14045,N_14060);
nand U14372 (N_14372,N_14053,N_14144);
nor U14373 (N_14373,N_14122,N_14101);
or U14374 (N_14374,N_14183,N_14048);
nor U14375 (N_14375,N_14128,N_14174);
xor U14376 (N_14376,N_14051,N_14163);
and U14377 (N_14377,N_14092,N_14166);
nand U14378 (N_14378,N_14036,N_14146);
nor U14379 (N_14379,N_14064,N_14041);
and U14380 (N_14380,N_14067,N_14025);
or U14381 (N_14381,N_14157,N_14114);
nand U14382 (N_14382,N_14116,N_14023);
or U14383 (N_14383,N_14134,N_14125);
nor U14384 (N_14384,N_14006,N_14150);
and U14385 (N_14385,N_14022,N_14147);
and U14386 (N_14386,N_14035,N_14037);
nor U14387 (N_14387,N_14184,N_14095);
or U14388 (N_14388,N_14074,N_14051);
and U14389 (N_14389,N_14178,N_14159);
nor U14390 (N_14390,N_14069,N_14001);
and U14391 (N_14391,N_14170,N_14049);
and U14392 (N_14392,N_14030,N_14043);
nand U14393 (N_14393,N_14124,N_14107);
nand U14394 (N_14394,N_14009,N_14046);
nand U14395 (N_14395,N_14192,N_14176);
or U14396 (N_14396,N_14083,N_14138);
or U14397 (N_14397,N_14108,N_14100);
nand U14398 (N_14398,N_14170,N_14126);
xor U14399 (N_14399,N_14061,N_14002);
nor U14400 (N_14400,N_14337,N_14287);
nor U14401 (N_14401,N_14214,N_14275);
nand U14402 (N_14402,N_14314,N_14347);
or U14403 (N_14403,N_14306,N_14340);
and U14404 (N_14404,N_14398,N_14213);
and U14405 (N_14405,N_14239,N_14290);
or U14406 (N_14406,N_14203,N_14258);
or U14407 (N_14407,N_14349,N_14238);
and U14408 (N_14408,N_14270,N_14206);
and U14409 (N_14409,N_14378,N_14274);
nand U14410 (N_14410,N_14388,N_14233);
and U14411 (N_14411,N_14363,N_14295);
or U14412 (N_14412,N_14226,N_14269);
nand U14413 (N_14413,N_14305,N_14297);
and U14414 (N_14414,N_14389,N_14261);
and U14415 (N_14415,N_14367,N_14382);
nand U14416 (N_14416,N_14322,N_14205);
and U14417 (N_14417,N_14257,N_14312);
or U14418 (N_14418,N_14341,N_14323);
and U14419 (N_14419,N_14212,N_14384);
or U14420 (N_14420,N_14316,N_14273);
nor U14421 (N_14421,N_14250,N_14379);
nor U14422 (N_14422,N_14211,N_14210);
xnor U14423 (N_14423,N_14240,N_14373);
or U14424 (N_14424,N_14393,N_14215);
or U14425 (N_14425,N_14292,N_14286);
nor U14426 (N_14426,N_14247,N_14326);
nor U14427 (N_14427,N_14396,N_14390);
and U14428 (N_14428,N_14294,N_14264);
and U14429 (N_14429,N_14299,N_14332);
nor U14430 (N_14430,N_14364,N_14344);
nand U14431 (N_14431,N_14317,N_14267);
and U14432 (N_14432,N_14370,N_14200);
and U14433 (N_14433,N_14204,N_14350);
and U14434 (N_14434,N_14217,N_14228);
nand U14435 (N_14435,N_14324,N_14331);
and U14436 (N_14436,N_14333,N_14361);
and U14437 (N_14437,N_14289,N_14220);
or U14438 (N_14438,N_14381,N_14319);
nand U14439 (N_14439,N_14293,N_14309);
or U14440 (N_14440,N_14207,N_14387);
nor U14441 (N_14441,N_14300,N_14249);
nand U14442 (N_14442,N_14385,N_14298);
nand U14443 (N_14443,N_14236,N_14260);
and U14444 (N_14444,N_14235,N_14377);
nor U14445 (N_14445,N_14234,N_14345);
nor U14446 (N_14446,N_14380,N_14291);
or U14447 (N_14447,N_14343,N_14328);
and U14448 (N_14448,N_14383,N_14315);
or U14449 (N_14449,N_14329,N_14266);
or U14450 (N_14450,N_14359,N_14218);
nand U14451 (N_14451,N_14395,N_14368);
nand U14452 (N_14452,N_14375,N_14366);
nor U14453 (N_14453,N_14357,N_14369);
xor U14454 (N_14454,N_14285,N_14253);
nand U14455 (N_14455,N_14334,N_14224);
or U14456 (N_14456,N_14254,N_14356);
nor U14457 (N_14457,N_14263,N_14372);
or U14458 (N_14458,N_14321,N_14320);
nand U14459 (N_14459,N_14346,N_14245);
or U14460 (N_14460,N_14342,N_14313);
nand U14461 (N_14461,N_14251,N_14242);
and U14462 (N_14462,N_14386,N_14376);
nor U14463 (N_14463,N_14283,N_14237);
and U14464 (N_14464,N_14255,N_14256);
nand U14465 (N_14465,N_14311,N_14248);
nor U14466 (N_14466,N_14252,N_14307);
or U14467 (N_14467,N_14353,N_14310);
xor U14468 (N_14468,N_14223,N_14230);
or U14469 (N_14469,N_14338,N_14371);
or U14470 (N_14470,N_14277,N_14243);
and U14471 (N_14471,N_14259,N_14244);
nand U14472 (N_14472,N_14339,N_14348);
nor U14473 (N_14473,N_14351,N_14282);
or U14474 (N_14474,N_14335,N_14365);
and U14475 (N_14475,N_14330,N_14280);
nor U14476 (N_14476,N_14231,N_14272);
or U14477 (N_14477,N_14318,N_14394);
nor U14478 (N_14478,N_14225,N_14281);
nor U14479 (N_14479,N_14209,N_14278);
nor U14480 (N_14480,N_14219,N_14221);
nor U14481 (N_14481,N_14284,N_14288);
and U14482 (N_14482,N_14303,N_14279);
xnor U14483 (N_14483,N_14399,N_14268);
nor U14484 (N_14484,N_14355,N_14336);
nand U14485 (N_14485,N_14302,N_14229);
and U14486 (N_14486,N_14208,N_14301);
or U14487 (N_14487,N_14202,N_14232);
nor U14488 (N_14488,N_14391,N_14362);
and U14489 (N_14489,N_14358,N_14308);
and U14490 (N_14490,N_14360,N_14216);
and U14491 (N_14491,N_14227,N_14296);
nand U14492 (N_14492,N_14201,N_14222);
and U14493 (N_14493,N_14352,N_14354);
nand U14494 (N_14494,N_14397,N_14271);
or U14495 (N_14495,N_14262,N_14327);
nand U14496 (N_14496,N_14304,N_14241);
nand U14497 (N_14497,N_14392,N_14265);
nand U14498 (N_14498,N_14374,N_14276);
or U14499 (N_14499,N_14246,N_14325);
and U14500 (N_14500,N_14309,N_14351);
nor U14501 (N_14501,N_14284,N_14331);
or U14502 (N_14502,N_14313,N_14378);
xnor U14503 (N_14503,N_14394,N_14240);
xor U14504 (N_14504,N_14374,N_14359);
or U14505 (N_14505,N_14211,N_14200);
and U14506 (N_14506,N_14276,N_14347);
and U14507 (N_14507,N_14284,N_14327);
nand U14508 (N_14508,N_14344,N_14219);
nand U14509 (N_14509,N_14295,N_14339);
or U14510 (N_14510,N_14247,N_14316);
and U14511 (N_14511,N_14343,N_14381);
and U14512 (N_14512,N_14292,N_14218);
and U14513 (N_14513,N_14231,N_14204);
or U14514 (N_14514,N_14331,N_14352);
nor U14515 (N_14515,N_14316,N_14325);
and U14516 (N_14516,N_14326,N_14379);
nand U14517 (N_14517,N_14241,N_14383);
xnor U14518 (N_14518,N_14333,N_14200);
or U14519 (N_14519,N_14363,N_14323);
and U14520 (N_14520,N_14347,N_14288);
nor U14521 (N_14521,N_14344,N_14378);
or U14522 (N_14522,N_14364,N_14231);
and U14523 (N_14523,N_14227,N_14396);
and U14524 (N_14524,N_14258,N_14248);
xor U14525 (N_14525,N_14254,N_14324);
nand U14526 (N_14526,N_14202,N_14223);
nand U14527 (N_14527,N_14263,N_14370);
or U14528 (N_14528,N_14295,N_14332);
nor U14529 (N_14529,N_14201,N_14230);
or U14530 (N_14530,N_14294,N_14304);
nor U14531 (N_14531,N_14217,N_14286);
nand U14532 (N_14532,N_14376,N_14280);
nor U14533 (N_14533,N_14313,N_14348);
nand U14534 (N_14534,N_14233,N_14332);
and U14535 (N_14535,N_14251,N_14342);
nor U14536 (N_14536,N_14275,N_14240);
and U14537 (N_14537,N_14226,N_14360);
nand U14538 (N_14538,N_14220,N_14329);
or U14539 (N_14539,N_14370,N_14394);
nor U14540 (N_14540,N_14305,N_14250);
or U14541 (N_14541,N_14250,N_14316);
and U14542 (N_14542,N_14393,N_14256);
nor U14543 (N_14543,N_14341,N_14272);
and U14544 (N_14544,N_14263,N_14397);
nand U14545 (N_14545,N_14261,N_14234);
or U14546 (N_14546,N_14331,N_14294);
or U14547 (N_14547,N_14221,N_14318);
nand U14548 (N_14548,N_14326,N_14321);
nand U14549 (N_14549,N_14377,N_14386);
nand U14550 (N_14550,N_14269,N_14316);
xor U14551 (N_14551,N_14231,N_14314);
nor U14552 (N_14552,N_14337,N_14279);
nand U14553 (N_14553,N_14268,N_14395);
xor U14554 (N_14554,N_14305,N_14213);
nor U14555 (N_14555,N_14245,N_14237);
nand U14556 (N_14556,N_14389,N_14398);
and U14557 (N_14557,N_14293,N_14220);
nor U14558 (N_14558,N_14333,N_14287);
nand U14559 (N_14559,N_14299,N_14206);
and U14560 (N_14560,N_14358,N_14318);
or U14561 (N_14561,N_14308,N_14335);
nor U14562 (N_14562,N_14242,N_14347);
or U14563 (N_14563,N_14257,N_14295);
or U14564 (N_14564,N_14235,N_14364);
nor U14565 (N_14565,N_14338,N_14348);
nand U14566 (N_14566,N_14361,N_14366);
or U14567 (N_14567,N_14398,N_14287);
or U14568 (N_14568,N_14245,N_14254);
nand U14569 (N_14569,N_14211,N_14238);
nor U14570 (N_14570,N_14239,N_14202);
nor U14571 (N_14571,N_14344,N_14301);
nand U14572 (N_14572,N_14240,N_14215);
or U14573 (N_14573,N_14363,N_14395);
or U14574 (N_14574,N_14356,N_14299);
nand U14575 (N_14575,N_14321,N_14208);
nor U14576 (N_14576,N_14314,N_14310);
nor U14577 (N_14577,N_14300,N_14279);
or U14578 (N_14578,N_14256,N_14237);
nor U14579 (N_14579,N_14280,N_14224);
or U14580 (N_14580,N_14349,N_14397);
and U14581 (N_14581,N_14269,N_14295);
nand U14582 (N_14582,N_14305,N_14236);
and U14583 (N_14583,N_14222,N_14354);
nor U14584 (N_14584,N_14265,N_14238);
nand U14585 (N_14585,N_14280,N_14234);
or U14586 (N_14586,N_14353,N_14385);
and U14587 (N_14587,N_14364,N_14336);
nand U14588 (N_14588,N_14350,N_14389);
nor U14589 (N_14589,N_14272,N_14218);
or U14590 (N_14590,N_14395,N_14359);
or U14591 (N_14591,N_14334,N_14299);
nor U14592 (N_14592,N_14339,N_14376);
or U14593 (N_14593,N_14366,N_14204);
nor U14594 (N_14594,N_14380,N_14329);
nor U14595 (N_14595,N_14358,N_14217);
and U14596 (N_14596,N_14266,N_14243);
or U14597 (N_14597,N_14271,N_14366);
and U14598 (N_14598,N_14361,N_14319);
nor U14599 (N_14599,N_14363,N_14296);
nand U14600 (N_14600,N_14496,N_14519);
nor U14601 (N_14601,N_14597,N_14404);
nand U14602 (N_14602,N_14579,N_14440);
nand U14603 (N_14603,N_14569,N_14598);
nor U14604 (N_14604,N_14526,N_14459);
nor U14605 (N_14605,N_14448,N_14441);
nor U14606 (N_14606,N_14456,N_14555);
or U14607 (N_14607,N_14577,N_14430);
nor U14608 (N_14608,N_14432,N_14501);
and U14609 (N_14609,N_14450,N_14524);
or U14610 (N_14610,N_14495,N_14537);
or U14611 (N_14611,N_14434,N_14594);
nand U14612 (N_14612,N_14575,N_14509);
nor U14613 (N_14613,N_14408,N_14467);
nand U14614 (N_14614,N_14489,N_14446);
or U14615 (N_14615,N_14425,N_14527);
or U14616 (N_14616,N_14589,N_14436);
nand U14617 (N_14617,N_14560,N_14574);
or U14618 (N_14618,N_14426,N_14571);
nand U14619 (N_14619,N_14549,N_14592);
nor U14620 (N_14620,N_14573,N_14559);
nor U14621 (N_14621,N_14578,N_14492);
xnor U14622 (N_14622,N_14523,N_14444);
nand U14623 (N_14623,N_14529,N_14503);
nand U14624 (N_14624,N_14542,N_14435);
and U14625 (N_14625,N_14507,N_14505);
nand U14626 (N_14626,N_14593,N_14469);
and U14627 (N_14627,N_14514,N_14530);
or U14628 (N_14628,N_14554,N_14424);
nand U14629 (N_14629,N_14468,N_14499);
nor U14630 (N_14630,N_14451,N_14536);
nor U14631 (N_14631,N_14419,N_14453);
xor U14632 (N_14632,N_14525,N_14403);
and U14633 (N_14633,N_14420,N_14457);
and U14634 (N_14634,N_14515,N_14433);
and U14635 (N_14635,N_14556,N_14476);
nor U14636 (N_14636,N_14405,N_14557);
and U14637 (N_14637,N_14564,N_14413);
or U14638 (N_14638,N_14570,N_14493);
or U14639 (N_14639,N_14502,N_14581);
and U14640 (N_14640,N_14548,N_14479);
or U14641 (N_14641,N_14544,N_14498);
nor U14642 (N_14642,N_14506,N_14484);
or U14643 (N_14643,N_14587,N_14416);
nor U14644 (N_14644,N_14494,N_14483);
nand U14645 (N_14645,N_14504,N_14552);
nand U14646 (N_14646,N_14562,N_14533);
nand U14647 (N_14647,N_14462,N_14547);
nand U14648 (N_14648,N_14568,N_14541);
and U14649 (N_14649,N_14422,N_14497);
nand U14650 (N_14650,N_14461,N_14539);
and U14651 (N_14651,N_14463,N_14521);
and U14652 (N_14652,N_14400,N_14576);
nor U14653 (N_14653,N_14500,N_14595);
xor U14654 (N_14654,N_14517,N_14565);
and U14655 (N_14655,N_14474,N_14510);
and U14656 (N_14656,N_14477,N_14466);
nor U14657 (N_14657,N_14478,N_14572);
or U14658 (N_14658,N_14508,N_14402);
nor U14659 (N_14659,N_14580,N_14485);
or U14660 (N_14660,N_14550,N_14567);
and U14661 (N_14661,N_14518,N_14584);
or U14662 (N_14662,N_14472,N_14455);
and U14663 (N_14663,N_14561,N_14428);
nand U14664 (N_14664,N_14558,N_14540);
and U14665 (N_14665,N_14454,N_14599);
or U14666 (N_14666,N_14427,N_14487);
nor U14667 (N_14667,N_14417,N_14407);
and U14668 (N_14668,N_14591,N_14482);
and U14669 (N_14669,N_14583,N_14488);
nor U14670 (N_14670,N_14409,N_14532);
or U14671 (N_14671,N_14406,N_14520);
nand U14672 (N_14672,N_14442,N_14538);
nand U14673 (N_14673,N_14438,N_14473);
nand U14674 (N_14674,N_14491,N_14423);
nor U14675 (N_14675,N_14534,N_14411);
nor U14676 (N_14676,N_14588,N_14415);
nor U14677 (N_14677,N_14543,N_14585);
nand U14678 (N_14678,N_14590,N_14464);
or U14679 (N_14679,N_14445,N_14437);
and U14680 (N_14680,N_14586,N_14401);
nor U14681 (N_14681,N_14460,N_14596);
and U14682 (N_14682,N_14452,N_14481);
or U14683 (N_14683,N_14414,N_14513);
or U14684 (N_14684,N_14418,N_14553);
and U14685 (N_14685,N_14470,N_14421);
nor U14686 (N_14686,N_14522,N_14475);
or U14687 (N_14687,N_14447,N_14449);
nor U14688 (N_14688,N_14471,N_14516);
nand U14689 (N_14689,N_14511,N_14582);
and U14690 (N_14690,N_14566,N_14443);
and U14691 (N_14691,N_14546,N_14545);
nand U14692 (N_14692,N_14490,N_14458);
and U14693 (N_14693,N_14410,N_14431);
nor U14694 (N_14694,N_14412,N_14486);
nand U14695 (N_14695,N_14512,N_14480);
nand U14696 (N_14696,N_14528,N_14429);
and U14697 (N_14697,N_14465,N_14531);
nor U14698 (N_14698,N_14551,N_14535);
or U14699 (N_14699,N_14439,N_14563);
or U14700 (N_14700,N_14553,N_14510);
and U14701 (N_14701,N_14492,N_14530);
nor U14702 (N_14702,N_14525,N_14504);
nand U14703 (N_14703,N_14583,N_14522);
nand U14704 (N_14704,N_14434,N_14567);
nand U14705 (N_14705,N_14453,N_14517);
and U14706 (N_14706,N_14545,N_14557);
or U14707 (N_14707,N_14407,N_14537);
nor U14708 (N_14708,N_14519,N_14528);
nor U14709 (N_14709,N_14433,N_14599);
or U14710 (N_14710,N_14491,N_14479);
and U14711 (N_14711,N_14528,N_14576);
and U14712 (N_14712,N_14560,N_14593);
nand U14713 (N_14713,N_14596,N_14405);
nand U14714 (N_14714,N_14449,N_14550);
or U14715 (N_14715,N_14524,N_14511);
or U14716 (N_14716,N_14482,N_14547);
nor U14717 (N_14717,N_14586,N_14453);
or U14718 (N_14718,N_14418,N_14454);
or U14719 (N_14719,N_14524,N_14543);
nor U14720 (N_14720,N_14598,N_14579);
nor U14721 (N_14721,N_14481,N_14526);
nand U14722 (N_14722,N_14475,N_14480);
or U14723 (N_14723,N_14561,N_14440);
or U14724 (N_14724,N_14546,N_14403);
or U14725 (N_14725,N_14408,N_14510);
or U14726 (N_14726,N_14469,N_14545);
or U14727 (N_14727,N_14428,N_14533);
or U14728 (N_14728,N_14598,N_14543);
nand U14729 (N_14729,N_14457,N_14559);
and U14730 (N_14730,N_14438,N_14456);
and U14731 (N_14731,N_14487,N_14584);
and U14732 (N_14732,N_14433,N_14533);
and U14733 (N_14733,N_14590,N_14589);
and U14734 (N_14734,N_14478,N_14455);
nand U14735 (N_14735,N_14435,N_14515);
nand U14736 (N_14736,N_14521,N_14480);
nand U14737 (N_14737,N_14467,N_14584);
nand U14738 (N_14738,N_14417,N_14554);
or U14739 (N_14739,N_14529,N_14443);
and U14740 (N_14740,N_14562,N_14515);
nor U14741 (N_14741,N_14521,N_14475);
nand U14742 (N_14742,N_14481,N_14573);
or U14743 (N_14743,N_14408,N_14493);
nor U14744 (N_14744,N_14556,N_14450);
xor U14745 (N_14745,N_14584,N_14594);
and U14746 (N_14746,N_14523,N_14547);
nand U14747 (N_14747,N_14470,N_14458);
or U14748 (N_14748,N_14537,N_14430);
nor U14749 (N_14749,N_14485,N_14590);
nor U14750 (N_14750,N_14565,N_14440);
or U14751 (N_14751,N_14551,N_14420);
nand U14752 (N_14752,N_14441,N_14430);
and U14753 (N_14753,N_14524,N_14576);
nand U14754 (N_14754,N_14522,N_14488);
xnor U14755 (N_14755,N_14574,N_14426);
and U14756 (N_14756,N_14448,N_14419);
and U14757 (N_14757,N_14418,N_14416);
nand U14758 (N_14758,N_14493,N_14585);
xor U14759 (N_14759,N_14551,N_14548);
nor U14760 (N_14760,N_14403,N_14581);
and U14761 (N_14761,N_14462,N_14542);
nor U14762 (N_14762,N_14469,N_14467);
and U14763 (N_14763,N_14414,N_14573);
and U14764 (N_14764,N_14427,N_14418);
and U14765 (N_14765,N_14531,N_14501);
nor U14766 (N_14766,N_14596,N_14454);
and U14767 (N_14767,N_14539,N_14447);
nand U14768 (N_14768,N_14476,N_14400);
or U14769 (N_14769,N_14512,N_14564);
and U14770 (N_14770,N_14544,N_14509);
nor U14771 (N_14771,N_14431,N_14479);
xor U14772 (N_14772,N_14401,N_14534);
or U14773 (N_14773,N_14488,N_14587);
nor U14774 (N_14774,N_14565,N_14455);
nor U14775 (N_14775,N_14531,N_14549);
and U14776 (N_14776,N_14495,N_14471);
xor U14777 (N_14777,N_14534,N_14548);
and U14778 (N_14778,N_14473,N_14414);
nand U14779 (N_14779,N_14414,N_14588);
or U14780 (N_14780,N_14430,N_14510);
nor U14781 (N_14781,N_14574,N_14485);
nand U14782 (N_14782,N_14539,N_14560);
and U14783 (N_14783,N_14550,N_14597);
or U14784 (N_14784,N_14592,N_14526);
nand U14785 (N_14785,N_14485,N_14569);
nor U14786 (N_14786,N_14501,N_14594);
and U14787 (N_14787,N_14564,N_14502);
nor U14788 (N_14788,N_14483,N_14474);
nand U14789 (N_14789,N_14491,N_14512);
or U14790 (N_14790,N_14532,N_14428);
or U14791 (N_14791,N_14592,N_14530);
or U14792 (N_14792,N_14537,N_14424);
nand U14793 (N_14793,N_14493,N_14582);
and U14794 (N_14794,N_14437,N_14589);
or U14795 (N_14795,N_14532,N_14407);
or U14796 (N_14796,N_14491,N_14485);
and U14797 (N_14797,N_14498,N_14504);
xor U14798 (N_14798,N_14403,N_14597);
nand U14799 (N_14799,N_14554,N_14443);
nand U14800 (N_14800,N_14777,N_14794);
and U14801 (N_14801,N_14733,N_14782);
nand U14802 (N_14802,N_14750,N_14604);
nor U14803 (N_14803,N_14679,N_14779);
nand U14804 (N_14804,N_14764,N_14703);
xor U14805 (N_14805,N_14690,N_14674);
and U14806 (N_14806,N_14633,N_14704);
nor U14807 (N_14807,N_14728,N_14644);
nand U14808 (N_14808,N_14743,N_14762);
and U14809 (N_14809,N_14744,N_14615);
and U14810 (N_14810,N_14659,N_14793);
nor U14811 (N_14811,N_14612,N_14607);
and U14812 (N_14812,N_14675,N_14647);
or U14813 (N_14813,N_14742,N_14732);
nand U14814 (N_14814,N_14713,N_14684);
or U14815 (N_14815,N_14619,N_14668);
nor U14816 (N_14816,N_14747,N_14796);
nand U14817 (N_14817,N_14707,N_14798);
nand U14818 (N_14818,N_14755,N_14697);
nand U14819 (N_14819,N_14759,N_14631);
or U14820 (N_14820,N_14771,N_14624);
nand U14821 (N_14821,N_14692,N_14613);
or U14822 (N_14822,N_14652,N_14716);
or U14823 (N_14823,N_14726,N_14712);
and U14824 (N_14824,N_14710,N_14786);
xnor U14825 (N_14825,N_14635,N_14775);
or U14826 (N_14826,N_14736,N_14671);
nor U14827 (N_14827,N_14702,N_14686);
nand U14828 (N_14828,N_14774,N_14749);
and U14829 (N_14829,N_14791,N_14795);
nor U14830 (N_14830,N_14719,N_14783);
or U14831 (N_14831,N_14642,N_14694);
and U14832 (N_14832,N_14722,N_14617);
nand U14833 (N_14833,N_14641,N_14706);
nor U14834 (N_14834,N_14632,N_14741);
nor U14835 (N_14835,N_14745,N_14663);
nand U14836 (N_14836,N_14614,N_14778);
and U14837 (N_14837,N_14609,N_14622);
nand U14838 (N_14838,N_14754,N_14653);
and U14839 (N_14839,N_14691,N_14763);
or U14840 (N_14840,N_14689,N_14621);
nor U14841 (N_14841,N_14758,N_14651);
nand U14842 (N_14842,N_14780,N_14799);
nor U14843 (N_14843,N_14715,N_14648);
nand U14844 (N_14844,N_14616,N_14623);
and U14845 (N_14845,N_14753,N_14611);
nor U14846 (N_14846,N_14629,N_14752);
nor U14847 (N_14847,N_14678,N_14693);
nand U14848 (N_14848,N_14731,N_14768);
or U14849 (N_14849,N_14602,N_14725);
or U14850 (N_14850,N_14717,N_14682);
and U14851 (N_14851,N_14688,N_14746);
nand U14852 (N_14852,N_14672,N_14676);
nor U14853 (N_14853,N_14767,N_14657);
and U14854 (N_14854,N_14681,N_14637);
and U14855 (N_14855,N_14720,N_14721);
and U14856 (N_14856,N_14660,N_14698);
xnor U14857 (N_14857,N_14656,N_14711);
nand U14858 (N_14858,N_14639,N_14792);
or U14859 (N_14859,N_14789,N_14603);
nor U14860 (N_14860,N_14646,N_14634);
nand U14861 (N_14861,N_14640,N_14667);
and U14862 (N_14862,N_14709,N_14649);
and U14863 (N_14863,N_14769,N_14654);
nor U14864 (N_14864,N_14655,N_14738);
nand U14865 (N_14865,N_14636,N_14626);
and U14866 (N_14866,N_14628,N_14605);
or U14867 (N_14867,N_14724,N_14670);
or U14868 (N_14868,N_14773,N_14797);
and U14869 (N_14869,N_14708,N_14705);
and U14870 (N_14870,N_14790,N_14665);
nor U14871 (N_14871,N_14739,N_14601);
or U14872 (N_14872,N_14608,N_14645);
nor U14873 (N_14873,N_14620,N_14756);
or U14874 (N_14874,N_14638,N_14760);
and U14875 (N_14875,N_14664,N_14680);
or U14876 (N_14876,N_14781,N_14748);
or U14877 (N_14877,N_14772,N_14699);
and U14878 (N_14878,N_14625,N_14701);
or U14879 (N_14879,N_14788,N_14770);
nand U14880 (N_14880,N_14661,N_14666);
or U14881 (N_14881,N_14696,N_14730);
nand U14882 (N_14882,N_14761,N_14662);
or U14883 (N_14883,N_14729,N_14751);
or U14884 (N_14884,N_14723,N_14785);
or U14885 (N_14885,N_14734,N_14683);
nor U14886 (N_14886,N_14776,N_14757);
nor U14887 (N_14887,N_14784,N_14766);
nand U14888 (N_14888,N_14695,N_14727);
and U14889 (N_14889,N_14765,N_14643);
or U14890 (N_14890,N_14658,N_14606);
nand U14891 (N_14891,N_14677,N_14669);
and U14892 (N_14892,N_14735,N_14718);
nand U14893 (N_14893,N_14610,N_14630);
or U14894 (N_14894,N_14627,N_14787);
nor U14895 (N_14895,N_14687,N_14600);
and U14896 (N_14896,N_14685,N_14740);
and U14897 (N_14897,N_14673,N_14650);
nor U14898 (N_14898,N_14700,N_14737);
or U14899 (N_14899,N_14618,N_14714);
and U14900 (N_14900,N_14699,N_14786);
and U14901 (N_14901,N_14734,N_14666);
or U14902 (N_14902,N_14707,N_14701);
nor U14903 (N_14903,N_14682,N_14642);
or U14904 (N_14904,N_14633,N_14785);
or U14905 (N_14905,N_14664,N_14688);
nand U14906 (N_14906,N_14794,N_14653);
nand U14907 (N_14907,N_14625,N_14698);
xor U14908 (N_14908,N_14789,N_14674);
nor U14909 (N_14909,N_14780,N_14744);
nand U14910 (N_14910,N_14619,N_14600);
nor U14911 (N_14911,N_14601,N_14691);
and U14912 (N_14912,N_14715,N_14659);
nor U14913 (N_14913,N_14615,N_14794);
and U14914 (N_14914,N_14781,N_14653);
or U14915 (N_14915,N_14645,N_14604);
nand U14916 (N_14916,N_14652,N_14722);
or U14917 (N_14917,N_14658,N_14688);
and U14918 (N_14918,N_14738,N_14613);
nand U14919 (N_14919,N_14650,N_14623);
nand U14920 (N_14920,N_14656,N_14686);
nand U14921 (N_14921,N_14637,N_14633);
or U14922 (N_14922,N_14641,N_14676);
nor U14923 (N_14923,N_14727,N_14772);
nand U14924 (N_14924,N_14732,N_14681);
or U14925 (N_14925,N_14781,N_14637);
nor U14926 (N_14926,N_14780,N_14724);
nand U14927 (N_14927,N_14750,N_14652);
and U14928 (N_14928,N_14764,N_14607);
or U14929 (N_14929,N_14641,N_14691);
nand U14930 (N_14930,N_14748,N_14797);
nand U14931 (N_14931,N_14794,N_14745);
nand U14932 (N_14932,N_14613,N_14666);
or U14933 (N_14933,N_14622,N_14686);
nor U14934 (N_14934,N_14722,N_14762);
and U14935 (N_14935,N_14753,N_14609);
nor U14936 (N_14936,N_14620,N_14625);
nand U14937 (N_14937,N_14664,N_14656);
and U14938 (N_14938,N_14676,N_14632);
nor U14939 (N_14939,N_14780,N_14711);
nor U14940 (N_14940,N_14623,N_14777);
nand U14941 (N_14941,N_14790,N_14735);
xor U14942 (N_14942,N_14632,N_14767);
xor U14943 (N_14943,N_14709,N_14753);
and U14944 (N_14944,N_14624,N_14614);
or U14945 (N_14945,N_14758,N_14626);
nor U14946 (N_14946,N_14673,N_14783);
nand U14947 (N_14947,N_14740,N_14764);
and U14948 (N_14948,N_14778,N_14665);
nor U14949 (N_14949,N_14686,N_14790);
xor U14950 (N_14950,N_14795,N_14720);
nand U14951 (N_14951,N_14751,N_14774);
or U14952 (N_14952,N_14728,N_14669);
or U14953 (N_14953,N_14717,N_14666);
or U14954 (N_14954,N_14794,N_14684);
or U14955 (N_14955,N_14614,N_14713);
or U14956 (N_14956,N_14615,N_14617);
nor U14957 (N_14957,N_14763,N_14754);
nor U14958 (N_14958,N_14611,N_14745);
nor U14959 (N_14959,N_14797,N_14693);
and U14960 (N_14960,N_14740,N_14678);
nor U14961 (N_14961,N_14773,N_14726);
and U14962 (N_14962,N_14670,N_14763);
xnor U14963 (N_14963,N_14739,N_14639);
or U14964 (N_14964,N_14650,N_14701);
and U14965 (N_14965,N_14763,N_14612);
nand U14966 (N_14966,N_14712,N_14600);
and U14967 (N_14967,N_14785,N_14766);
nand U14968 (N_14968,N_14764,N_14616);
and U14969 (N_14969,N_14689,N_14734);
and U14970 (N_14970,N_14619,N_14793);
or U14971 (N_14971,N_14644,N_14738);
xor U14972 (N_14972,N_14707,N_14704);
and U14973 (N_14973,N_14728,N_14764);
nor U14974 (N_14974,N_14614,N_14685);
or U14975 (N_14975,N_14688,N_14608);
and U14976 (N_14976,N_14720,N_14778);
and U14977 (N_14977,N_14751,N_14675);
and U14978 (N_14978,N_14626,N_14625);
or U14979 (N_14979,N_14743,N_14672);
xnor U14980 (N_14980,N_14797,N_14784);
nor U14981 (N_14981,N_14699,N_14751);
or U14982 (N_14982,N_14707,N_14732);
nor U14983 (N_14983,N_14602,N_14671);
and U14984 (N_14984,N_14620,N_14668);
or U14985 (N_14985,N_14643,N_14729);
nor U14986 (N_14986,N_14761,N_14683);
nand U14987 (N_14987,N_14672,N_14606);
nor U14988 (N_14988,N_14660,N_14683);
and U14989 (N_14989,N_14645,N_14696);
or U14990 (N_14990,N_14782,N_14723);
or U14991 (N_14991,N_14613,N_14707);
and U14992 (N_14992,N_14728,N_14735);
and U14993 (N_14993,N_14654,N_14621);
or U14994 (N_14994,N_14727,N_14616);
nor U14995 (N_14995,N_14659,N_14633);
nor U14996 (N_14996,N_14704,N_14648);
and U14997 (N_14997,N_14615,N_14755);
and U14998 (N_14998,N_14736,N_14721);
and U14999 (N_14999,N_14715,N_14780);
nor U15000 (N_15000,N_14917,N_14924);
nand U15001 (N_15001,N_14854,N_14839);
or U15002 (N_15002,N_14887,N_14956);
or U15003 (N_15003,N_14965,N_14810);
and U15004 (N_15004,N_14837,N_14934);
and U15005 (N_15005,N_14981,N_14951);
nand U15006 (N_15006,N_14930,N_14911);
and U15007 (N_15007,N_14952,N_14967);
xnor U15008 (N_15008,N_14989,N_14844);
nor U15009 (N_15009,N_14853,N_14868);
or U15010 (N_15010,N_14800,N_14835);
nor U15011 (N_15011,N_14976,N_14852);
nor U15012 (N_15012,N_14836,N_14914);
and U15013 (N_15013,N_14906,N_14802);
nand U15014 (N_15014,N_14954,N_14961);
nor U15015 (N_15015,N_14859,N_14849);
or U15016 (N_15016,N_14824,N_14979);
or U15017 (N_15017,N_14933,N_14960);
or U15018 (N_15018,N_14832,N_14807);
and U15019 (N_15019,N_14826,N_14827);
nor U15020 (N_15020,N_14829,N_14994);
or U15021 (N_15021,N_14897,N_14805);
nand U15022 (N_15022,N_14817,N_14885);
nand U15023 (N_15023,N_14957,N_14905);
and U15024 (N_15024,N_14898,N_14922);
nand U15025 (N_15025,N_14867,N_14937);
xor U15026 (N_15026,N_14808,N_14822);
nand U15027 (N_15027,N_14980,N_14935);
nand U15028 (N_15028,N_14964,N_14928);
nand U15029 (N_15029,N_14971,N_14975);
nand U15030 (N_15030,N_14955,N_14865);
and U15031 (N_15031,N_14878,N_14988);
nand U15032 (N_15032,N_14889,N_14936);
nand U15033 (N_15033,N_14846,N_14995);
or U15034 (N_15034,N_14904,N_14876);
or U15035 (N_15035,N_14909,N_14823);
nand U15036 (N_15036,N_14803,N_14863);
nand U15037 (N_15037,N_14931,N_14915);
or U15038 (N_15038,N_14834,N_14891);
nand U15039 (N_15039,N_14886,N_14926);
nor U15040 (N_15040,N_14820,N_14938);
nor U15041 (N_15041,N_14860,N_14812);
nand U15042 (N_15042,N_14929,N_14992);
and U15043 (N_15043,N_14809,N_14958);
nand U15044 (N_15044,N_14825,N_14972);
nand U15045 (N_15045,N_14841,N_14977);
nand U15046 (N_15046,N_14946,N_14959);
or U15047 (N_15047,N_14828,N_14923);
and U15048 (N_15048,N_14847,N_14850);
or U15049 (N_15049,N_14899,N_14881);
nand U15050 (N_15050,N_14996,N_14902);
or U15051 (N_15051,N_14893,N_14900);
or U15052 (N_15052,N_14940,N_14845);
nand U15053 (N_15053,N_14999,N_14816);
nor U15054 (N_15054,N_14920,N_14877);
nand U15055 (N_15055,N_14806,N_14963);
and U15056 (N_15056,N_14990,N_14895);
and U15057 (N_15057,N_14927,N_14862);
nor U15058 (N_15058,N_14883,N_14840);
or U15059 (N_15059,N_14998,N_14872);
nor U15060 (N_15060,N_14908,N_14821);
and U15061 (N_15061,N_14987,N_14871);
nand U15062 (N_15062,N_14907,N_14875);
nor U15063 (N_15063,N_14997,N_14811);
nor U15064 (N_15064,N_14813,N_14983);
nor U15065 (N_15065,N_14944,N_14966);
and U15066 (N_15066,N_14831,N_14892);
nand U15067 (N_15067,N_14901,N_14953);
nand U15068 (N_15068,N_14861,N_14888);
and U15069 (N_15069,N_14879,N_14857);
or U15070 (N_15070,N_14848,N_14880);
or U15071 (N_15071,N_14864,N_14945);
or U15072 (N_15072,N_14869,N_14921);
and U15073 (N_15073,N_14947,N_14939);
and U15074 (N_15074,N_14912,N_14974);
nor U15075 (N_15075,N_14882,N_14970);
nor U15076 (N_15076,N_14925,N_14910);
nor U15077 (N_15077,N_14818,N_14896);
nand U15078 (N_15078,N_14943,N_14833);
nand U15079 (N_15079,N_14903,N_14866);
or U15080 (N_15080,N_14843,N_14973);
or U15081 (N_15081,N_14819,N_14894);
or U15082 (N_15082,N_14949,N_14968);
and U15083 (N_15083,N_14948,N_14913);
or U15084 (N_15084,N_14858,N_14916);
and U15085 (N_15085,N_14842,N_14969);
nand U15086 (N_15086,N_14870,N_14985);
or U15087 (N_15087,N_14830,N_14838);
nor U15088 (N_15088,N_14993,N_14814);
nand U15089 (N_15089,N_14986,N_14962);
or U15090 (N_15090,N_14950,N_14855);
and U15091 (N_15091,N_14890,N_14932);
or U15092 (N_15092,N_14804,N_14984);
and U15093 (N_15093,N_14918,N_14874);
nor U15094 (N_15094,N_14851,N_14815);
nor U15095 (N_15095,N_14991,N_14884);
nand U15096 (N_15096,N_14856,N_14873);
or U15097 (N_15097,N_14919,N_14982);
or U15098 (N_15098,N_14942,N_14978);
nand U15099 (N_15099,N_14801,N_14941);
or U15100 (N_15100,N_14965,N_14819);
and U15101 (N_15101,N_14834,N_14869);
nor U15102 (N_15102,N_14826,N_14921);
or U15103 (N_15103,N_14885,N_14955);
nor U15104 (N_15104,N_14823,N_14944);
or U15105 (N_15105,N_14993,N_14804);
nor U15106 (N_15106,N_14849,N_14867);
or U15107 (N_15107,N_14871,N_14913);
or U15108 (N_15108,N_14987,N_14804);
and U15109 (N_15109,N_14933,N_14955);
or U15110 (N_15110,N_14990,N_14823);
nor U15111 (N_15111,N_14897,N_14862);
nand U15112 (N_15112,N_14926,N_14884);
nand U15113 (N_15113,N_14932,N_14833);
nor U15114 (N_15114,N_14958,N_14816);
or U15115 (N_15115,N_14885,N_14882);
nor U15116 (N_15116,N_14880,N_14852);
nand U15117 (N_15117,N_14924,N_14884);
nand U15118 (N_15118,N_14864,N_14976);
and U15119 (N_15119,N_14940,N_14956);
nand U15120 (N_15120,N_14835,N_14941);
xnor U15121 (N_15121,N_14931,N_14917);
and U15122 (N_15122,N_14926,N_14870);
nand U15123 (N_15123,N_14860,N_14879);
nand U15124 (N_15124,N_14901,N_14810);
and U15125 (N_15125,N_14904,N_14966);
or U15126 (N_15126,N_14945,N_14978);
or U15127 (N_15127,N_14968,N_14915);
nand U15128 (N_15128,N_14906,N_14860);
and U15129 (N_15129,N_14842,N_14800);
nand U15130 (N_15130,N_14909,N_14835);
nand U15131 (N_15131,N_14911,N_14896);
nor U15132 (N_15132,N_14922,N_14807);
xor U15133 (N_15133,N_14838,N_14857);
nand U15134 (N_15134,N_14965,N_14825);
and U15135 (N_15135,N_14999,N_14872);
or U15136 (N_15136,N_14847,N_14931);
or U15137 (N_15137,N_14888,N_14934);
nor U15138 (N_15138,N_14953,N_14890);
and U15139 (N_15139,N_14856,N_14949);
nand U15140 (N_15140,N_14876,N_14911);
nand U15141 (N_15141,N_14850,N_14914);
or U15142 (N_15142,N_14960,N_14883);
and U15143 (N_15143,N_14814,N_14959);
or U15144 (N_15144,N_14865,N_14914);
nor U15145 (N_15145,N_14873,N_14857);
nand U15146 (N_15146,N_14960,N_14921);
nor U15147 (N_15147,N_14834,N_14884);
or U15148 (N_15148,N_14839,N_14910);
and U15149 (N_15149,N_14936,N_14970);
xnor U15150 (N_15150,N_14891,N_14978);
or U15151 (N_15151,N_14975,N_14830);
nand U15152 (N_15152,N_14863,N_14843);
or U15153 (N_15153,N_14815,N_14920);
and U15154 (N_15154,N_14931,N_14839);
or U15155 (N_15155,N_14811,N_14900);
or U15156 (N_15156,N_14863,N_14828);
or U15157 (N_15157,N_14932,N_14828);
nor U15158 (N_15158,N_14913,N_14949);
and U15159 (N_15159,N_14910,N_14918);
nand U15160 (N_15160,N_14889,N_14973);
nand U15161 (N_15161,N_14879,N_14846);
or U15162 (N_15162,N_14900,N_14864);
and U15163 (N_15163,N_14841,N_14948);
and U15164 (N_15164,N_14818,N_14923);
nor U15165 (N_15165,N_14949,N_14899);
nor U15166 (N_15166,N_14938,N_14843);
or U15167 (N_15167,N_14804,N_14836);
nand U15168 (N_15168,N_14894,N_14988);
or U15169 (N_15169,N_14887,N_14914);
nor U15170 (N_15170,N_14829,N_14993);
xor U15171 (N_15171,N_14980,N_14910);
or U15172 (N_15172,N_14906,N_14937);
nand U15173 (N_15173,N_14831,N_14992);
and U15174 (N_15174,N_14950,N_14969);
or U15175 (N_15175,N_14820,N_14952);
or U15176 (N_15176,N_14879,N_14885);
nor U15177 (N_15177,N_14899,N_14825);
or U15178 (N_15178,N_14910,N_14901);
and U15179 (N_15179,N_14851,N_14829);
or U15180 (N_15180,N_14863,N_14810);
nor U15181 (N_15181,N_14870,N_14816);
and U15182 (N_15182,N_14997,N_14812);
and U15183 (N_15183,N_14921,N_14866);
nor U15184 (N_15184,N_14905,N_14956);
nor U15185 (N_15185,N_14912,N_14815);
nand U15186 (N_15186,N_14945,N_14870);
nor U15187 (N_15187,N_14918,N_14937);
nor U15188 (N_15188,N_14841,N_14844);
nor U15189 (N_15189,N_14841,N_14989);
xnor U15190 (N_15190,N_14896,N_14802);
or U15191 (N_15191,N_14908,N_14969);
nand U15192 (N_15192,N_14923,N_14853);
nor U15193 (N_15193,N_14969,N_14848);
and U15194 (N_15194,N_14973,N_14911);
nor U15195 (N_15195,N_14813,N_14839);
nand U15196 (N_15196,N_14833,N_14888);
nand U15197 (N_15197,N_14954,N_14970);
or U15198 (N_15198,N_14919,N_14800);
nor U15199 (N_15199,N_14830,N_14803);
nor U15200 (N_15200,N_15128,N_15097);
nand U15201 (N_15201,N_15112,N_15003);
and U15202 (N_15202,N_15163,N_15186);
and U15203 (N_15203,N_15007,N_15054);
or U15204 (N_15204,N_15087,N_15149);
and U15205 (N_15205,N_15002,N_15019);
nand U15206 (N_15206,N_15071,N_15173);
and U15207 (N_15207,N_15113,N_15062);
nor U15208 (N_15208,N_15165,N_15020);
nor U15209 (N_15209,N_15065,N_15042);
nand U15210 (N_15210,N_15194,N_15089);
or U15211 (N_15211,N_15157,N_15013);
nor U15212 (N_15212,N_15198,N_15080);
nor U15213 (N_15213,N_15055,N_15048);
or U15214 (N_15214,N_15075,N_15061);
and U15215 (N_15215,N_15144,N_15159);
nand U15216 (N_15216,N_15076,N_15098);
nand U15217 (N_15217,N_15074,N_15132);
or U15218 (N_15218,N_15050,N_15160);
nor U15219 (N_15219,N_15183,N_15170);
nor U15220 (N_15220,N_15116,N_15038);
and U15221 (N_15221,N_15179,N_15049);
nand U15222 (N_15222,N_15109,N_15090);
and U15223 (N_15223,N_15051,N_15127);
nand U15224 (N_15224,N_15084,N_15135);
or U15225 (N_15225,N_15063,N_15047);
or U15226 (N_15226,N_15091,N_15199);
nor U15227 (N_15227,N_15122,N_15012);
or U15228 (N_15228,N_15083,N_15150);
nand U15229 (N_15229,N_15192,N_15162);
nor U15230 (N_15230,N_15129,N_15161);
or U15231 (N_15231,N_15156,N_15033);
or U15232 (N_15232,N_15008,N_15147);
nor U15233 (N_15233,N_15145,N_15169);
and U15234 (N_15234,N_15015,N_15175);
and U15235 (N_15235,N_15124,N_15140);
and U15236 (N_15236,N_15028,N_15040);
nand U15237 (N_15237,N_15014,N_15103);
and U15238 (N_15238,N_15036,N_15184);
and U15239 (N_15239,N_15121,N_15011);
nor U15240 (N_15240,N_15096,N_15110);
nor U15241 (N_15241,N_15185,N_15095);
or U15242 (N_15242,N_15056,N_15106);
or U15243 (N_15243,N_15044,N_15088);
or U15244 (N_15244,N_15118,N_15093);
nand U15245 (N_15245,N_15025,N_15153);
and U15246 (N_15246,N_15057,N_15060);
and U15247 (N_15247,N_15041,N_15154);
nand U15248 (N_15248,N_15176,N_15142);
xnor U15249 (N_15249,N_15077,N_15148);
nand U15250 (N_15250,N_15059,N_15182);
nor U15251 (N_15251,N_15026,N_15034);
and U15252 (N_15252,N_15081,N_15125);
or U15253 (N_15253,N_15187,N_15123);
nand U15254 (N_15254,N_15174,N_15104);
nand U15255 (N_15255,N_15195,N_15067);
nor U15256 (N_15256,N_15111,N_15130);
or U15257 (N_15257,N_15043,N_15004);
nand U15258 (N_15258,N_15178,N_15133);
or U15259 (N_15259,N_15092,N_15101);
or U15260 (N_15260,N_15181,N_15085);
or U15261 (N_15261,N_15068,N_15039);
nand U15262 (N_15262,N_15191,N_15006);
nand U15263 (N_15263,N_15079,N_15190);
or U15264 (N_15264,N_15022,N_15164);
nor U15265 (N_15265,N_15146,N_15070);
and U15266 (N_15266,N_15053,N_15086);
xnor U15267 (N_15267,N_15045,N_15143);
nand U15268 (N_15268,N_15027,N_15167);
nor U15269 (N_15269,N_15115,N_15134);
and U15270 (N_15270,N_15177,N_15108);
xor U15271 (N_15271,N_15107,N_15126);
and U15272 (N_15272,N_15171,N_15035);
or U15273 (N_15273,N_15131,N_15046);
or U15274 (N_15274,N_15094,N_15189);
and U15275 (N_15275,N_15117,N_15155);
or U15276 (N_15276,N_15137,N_15100);
or U15277 (N_15277,N_15172,N_15166);
xor U15278 (N_15278,N_15037,N_15193);
nor U15279 (N_15279,N_15024,N_15066);
nor U15280 (N_15280,N_15064,N_15139);
and U15281 (N_15281,N_15120,N_15138);
nor U15282 (N_15282,N_15082,N_15018);
or U15283 (N_15283,N_15023,N_15119);
nand U15284 (N_15284,N_15197,N_15016);
or U15285 (N_15285,N_15152,N_15099);
and U15286 (N_15286,N_15005,N_15009);
nand U15287 (N_15287,N_15141,N_15151);
and U15288 (N_15288,N_15000,N_15105);
or U15289 (N_15289,N_15069,N_15052);
and U15290 (N_15290,N_15168,N_15188);
and U15291 (N_15291,N_15073,N_15021);
nor U15292 (N_15292,N_15029,N_15072);
nand U15293 (N_15293,N_15017,N_15078);
nand U15294 (N_15294,N_15158,N_15136);
nor U15295 (N_15295,N_15031,N_15114);
nand U15296 (N_15296,N_15010,N_15030);
nand U15297 (N_15297,N_15058,N_15102);
nand U15298 (N_15298,N_15196,N_15180);
nand U15299 (N_15299,N_15001,N_15032);
nor U15300 (N_15300,N_15157,N_15162);
nor U15301 (N_15301,N_15108,N_15112);
and U15302 (N_15302,N_15167,N_15021);
nand U15303 (N_15303,N_15062,N_15103);
or U15304 (N_15304,N_15024,N_15110);
nor U15305 (N_15305,N_15074,N_15117);
nor U15306 (N_15306,N_15091,N_15022);
nor U15307 (N_15307,N_15030,N_15165);
nor U15308 (N_15308,N_15082,N_15042);
nand U15309 (N_15309,N_15036,N_15173);
or U15310 (N_15310,N_15146,N_15074);
or U15311 (N_15311,N_15190,N_15081);
or U15312 (N_15312,N_15036,N_15129);
nand U15313 (N_15313,N_15102,N_15025);
xor U15314 (N_15314,N_15104,N_15012);
or U15315 (N_15315,N_15055,N_15187);
nand U15316 (N_15316,N_15090,N_15001);
and U15317 (N_15317,N_15140,N_15126);
nand U15318 (N_15318,N_15156,N_15088);
and U15319 (N_15319,N_15094,N_15068);
nand U15320 (N_15320,N_15012,N_15148);
or U15321 (N_15321,N_15054,N_15048);
and U15322 (N_15322,N_15128,N_15162);
nor U15323 (N_15323,N_15149,N_15002);
nor U15324 (N_15324,N_15091,N_15151);
and U15325 (N_15325,N_15032,N_15009);
and U15326 (N_15326,N_15149,N_15031);
nand U15327 (N_15327,N_15091,N_15117);
nand U15328 (N_15328,N_15190,N_15123);
nand U15329 (N_15329,N_15061,N_15167);
and U15330 (N_15330,N_15199,N_15136);
nand U15331 (N_15331,N_15161,N_15122);
or U15332 (N_15332,N_15150,N_15054);
and U15333 (N_15333,N_15163,N_15134);
or U15334 (N_15334,N_15083,N_15142);
or U15335 (N_15335,N_15163,N_15178);
nand U15336 (N_15336,N_15093,N_15043);
nand U15337 (N_15337,N_15128,N_15108);
or U15338 (N_15338,N_15100,N_15060);
or U15339 (N_15339,N_15078,N_15111);
and U15340 (N_15340,N_15149,N_15062);
or U15341 (N_15341,N_15085,N_15092);
or U15342 (N_15342,N_15041,N_15118);
and U15343 (N_15343,N_15002,N_15055);
nor U15344 (N_15344,N_15026,N_15054);
and U15345 (N_15345,N_15180,N_15156);
or U15346 (N_15346,N_15142,N_15141);
or U15347 (N_15347,N_15141,N_15130);
nor U15348 (N_15348,N_15111,N_15042);
nand U15349 (N_15349,N_15021,N_15097);
nand U15350 (N_15350,N_15189,N_15018);
and U15351 (N_15351,N_15156,N_15087);
or U15352 (N_15352,N_15125,N_15045);
nor U15353 (N_15353,N_15003,N_15114);
and U15354 (N_15354,N_15177,N_15031);
nand U15355 (N_15355,N_15184,N_15052);
nor U15356 (N_15356,N_15018,N_15014);
nand U15357 (N_15357,N_15147,N_15084);
nand U15358 (N_15358,N_15001,N_15138);
nand U15359 (N_15359,N_15083,N_15075);
nand U15360 (N_15360,N_15161,N_15176);
or U15361 (N_15361,N_15175,N_15126);
nand U15362 (N_15362,N_15103,N_15093);
nand U15363 (N_15363,N_15170,N_15193);
and U15364 (N_15364,N_15033,N_15146);
or U15365 (N_15365,N_15175,N_15083);
or U15366 (N_15366,N_15126,N_15170);
nand U15367 (N_15367,N_15110,N_15176);
and U15368 (N_15368,N_15020,N_15111);
or U15369 (N_15369,N_15070,N_15147);
and U15370 (N_15370,N_15058,N_15001);
or U15371 (N_15371,N_15007,N_15024);
nand U15372 (N_15372,N_15143,N_15006);
nor U15373 (N_15373,N_15154,N_15167);
xnor U15374 (N_15374,N_15024,N_15107);
nor U15375 (N_15375,N_15179,N_15162);
and U15376 (N_15376,N_15003,N_15097);
xor U15377 (N_15377,N_15106,N_15095);
nor U15378 (N_15378,N_15045,N_15133);
and U15379 (N_15379,N_15028,N_15103);
or U15380 (N_15380,N_15109,N_15025);
nor U15381 (N_15381,N_15190,N_15090);
and U15382 (N_15382,N_15129,N_15187);
nand U15383 (N_15383,N_15046,N_15007);
nor U15384 (N_15384,N_15032,N_15183);
and U15385 (N_15385,N_15002,N_15075);
nand U15386 (N_15386,N_15133,N_15110);
and U15387 (N_15387,N_15067,N_15165);
nor U15388 (N_15388,N_15024,N_15148);
or U15389 (N_15389,N_15164,N_15148);
or U15390 (N_15390,N_15199,N_15093);
nand U15391 (N_15391,N_15025,N_15052);
and U15392 (N_15392,N_15056,N_15045);
or U15393 (N_15393,N_15172,N_15179);
nor U15394 (N_15394,N_15026,N_15082);
or U15395 (N_15395,N_15083,N_15015);
nand U15396 (N_15396,N_15168,N_15066);
or U15397 (N_15397,N_15171,N_15009);
nor U15398 (N_15398,N_15147,N_15122);
and U15399 (N_15399,N_15139,N_15158);
nand U15400 (N_15400,N_15346,N_15263);
nor U15401 (N_15401,N_15364,N_15215);
nand U15402 (N_15402,N_15200,N_15274);
or U15403 (N_15403,N_15305,N_15240);
nand U15404 (N_15404,N_15341,N_15242);
nor U15405 (N_15405,N_15219,N_15291);
or U15406 (N_15406,N_15233,N_15298);
nand U15407 (N_15407,N_15326,N_15335);
nand U15408 (N_15408,N_15210,N_15258);
nand U15409 (N_15409,N_15336,N_15322);
or U15410 (N_15410,N_15338,N_15262);
and U15411 (N_15411,N_15317,N_15371);
nand U15412 (N_15412,N_15390,N_15362);
nand U15413 (N_15413,N_15286,N_15299);
nand U15414 (N_15414,N_15208,N_15300);
and U15415 (N_15415,N_15348,N_15380);
or U15416 (N_15416,N_15321,N_15368);
nand U15417 (N_15417,N_15257,N_15279);
and U15418 (N_15418,N_15393,N_15352);
and U15419 (N_15419,N_15293,N_15342);
or U15420 (N_15420,N_15244,N_15354);
or U15421 (N_15421,N_15289,N_15343);
nor U15422 (N_15422,N_15246,N_15217);
nand U15423 (N_15423,N_15334,N_15234);
nor U15424 (N_15424,N_15382,N_15224);
or U15425 (N_15425,N_15302,N_15369);
nor U15426 (N_15426,N_15308,N_15271);
nand U15427 (N_15427,N_15238,N_15301);
and U15428 (N_15428,N_15207,N_15331);
and U15429 (N_15429,N_15222,N_15248);
or U15430 (N_15430,N_15282,N_15243);
and U15431 (N_15431,N_15265,N_15225);
and U15432 (N_15432,N_15391,N_15333);
or U15433 (N_15433,N_15351,N_15385);
nand U15434 (N_15434,N_15296,N_15350);
or U15435 (N_15435,N_15277,N_15211);
or U15436 (N_15436,N_15231,N_15314);
or U15437 (N_15437,N_15278,N_15344);
nand U15438 (N_15438,N_15376,N_15209);
nand U15439 (N_15439,N_15313,N_15239);
and U15440 (N_15440,N_15294,N_15212);
and U15441 (N_15441,N_15221,N_15230);
or U15442 (N_15442,N_15315,N_15259);
nand U15443 (N_15443,N_15247,N_15363);
nand U15444 (N_15444,N_15395,N_15310);
or U15445 (N_15445,N_15204,N_15353);
or U15446 (N_15446,N_15396,N_15304);
nor U15447 (N_15447,N_15366,N_15281);
or U15448 (N_15448,N_15307,N_15252);
nor U15449 (N_15449,N_15254,N_15276);
nand U15450 (N_15450,N_15398,N_15241);
or U15451 (N_15451,N_15303,N_15374);
nand U15452 (N_15452,N_15386,N_15378);
and U15453 (N_15453,N_15251,N_15201);
nor U15454 (N_15454,N_15202,N_15280);
nand U15455 (N_15455,N_15226,N_15216);
xor U15456 (N_15456,N_15250,N_15236);
nor U15457 (N_15457,N_15228,N_15345);
and U15458 (N_15458,N_15261,N_15397);
nor U15459 (N_15459,N_15218,N_15379);
nand U15460 (N_15460,N_15394,N_15266);
and U15461 (N_15461,N_15316,N_15339);
nor U15462 (N_15462,N_15381,N_15358);
nor U15463 (N_15463,N_15290,N_15332);
nand U15464 (N_15464,N_15213,N_15399);
xnor U15465 (N_15465,N_15311,N_15288);
nand U15466 (N_15466,N_15232,N_15355);
and U15467 (N_15467,N_15347,N_15267);
nor U15468 (N_15468,N_15206,N_15270);
and U15469 (N_15469,N_15273,N_15365);
nand U15470 (N_15470,N_15329,N_15235);
or U15471 (N_15471,N_15387,N_15327);
xnor U15472 (N_15472,N_15284,N_15330);
nand U15473 (N_15473,N_15367,N_15375);
and U15474 (N_15474,N_15320,N_15377);
nand U15475 (N_15475,N_15214,N_15260);
or U15476 (N_15476,N_15388,N_15323);
nand U15477 (N_15477,N_15357,N_15349);
or U15478 (N_15478,N_15227,N_15328);
or U15479 (N_15479,N_15384,N_15389);
nand U15480 (N_15480,N_15285,N_15253);
nor U15481 (N_15481,N_15361,N_15370);
nand U15482 (N_15482,N_15383,N_15372);
and U15483 (N_15483,N_15318,N_15295);
or U15484 (N_15484,N_15373,N_15268);
and U15485 (N_15485,N_15203,N_15287);
and U15486 (N_15486,N_15324,N_15360);
and U15487 (N_15487,N_15297,N_15337);
nor U15488 (N_15488,N_15256,N_15269);
nand U15489 (N_15489,N_15249,N_15319);
and U15490 (N_15490,N_15325,N_15283);
or U15491 (N_15491,N_15275,N_15264);
nor U15492 (N_15492,N_15392,N_15255);
or U15493 (N_15493,N_15356,N_15229);
and U15494 (N_15494,N_15359,N_15205);
or U15495 (N_15495,N_15312,N_15309);
and U15496 (N_15496,N_15245,N_15220);
or U15497 (N_15497,N_15223,N_15306);
and U15498 (N_15498,N_15237,N_15272);
nand U15499 (N_15499,N_15292,N_15340);
and U15500 (N_15500,N_15264,N_15278);
nor U15501 (N_15501,N_15212,N_15289);
or U15502 (N_15502,N_15367,N_15255);
nand U15503 (N_15503,N_15214,N_15268);
nor U15504 (N_15504,N_15249,N_15205);
and U15505 (N_15505,N_15265,N_15331);
nand U15506 (N_15506,N_15335,N_15301);
and U15507 (N_15507,N_15302,N_15220);
or U15508 (N_15508,N_15254,N_15327);
or U15509 (N_15509,N_15315,N_15370);
nand U15510 (N_15510,N_15298,N_15302);
nor U15511 (N_15511,N_15215,N_15243);
nor U15512 (N_15512,N_15390,N_15281);
nor U15513 (N_15513,N_15201,N_15317);
nand U15514 (N_15514,N_15285,N_15216);
or U15515 (N_15515,N_15365,N_15327);
nand U15516 (N_15516,N_15328,N_15393);
nor U15517 (N_15517,N_15300,N_15284);
or U15518 (N_15518,N_15212,N_15264);
nand U15519 (N_15519,N_15216,N_15234);
nor U15520 (N_15520,N_15309,N_15289);
nand U15521 (N_15521,N_15264,N_15310);
nand U15522 (N_15522,N_15243,N_15203);
nor U15523 (N_15523,N_15398,N_15387);
or U15524 (N_15524,N_15201,N_15316);
or U15525 (N_15525,N_15295,N_15307);
nand U15526 (N_15526,N_15208,N_15224);
and U15527 (N_15527,N_15259,N_15244);
nand U15528 (N_15528,N_15395,N_15222);
and U15529 (N_15529,N_15286,N_15337);
or U15530 (N_15530,N_15210,N_15222);
nor U15531 (N_15531,N_15250,N_15213);
or U15532 (N_15532,N_15325,N_15242);
nand U15533 (N_15533,N_15387,N_15309);
nand U15534 (N_15534,N_15371,N_15236);
and U15535 (N_15535,N_15309,N_15258);
and U15536 (N_15536,N_15364,N_15381);
nor U15537 (N_15537,N_15269,N_15234);
and U15538 (N_15538,N_15207,N_15387);
and U15539 (N_15539,N_15234,N_15301);
xnor U15540 (N_15540,N_15249,N_15209);
nand U15541 (N_15541,N_15206,N_15219);
or U15542 (N_15542,N_15283,N_15303);
and U15543 (N_15543,N_15338,N_15342);
nand U15544 (N_15544,N_15310,N_15311);
and U15545 (N_15545,N_15220,N_15390);
and U15546 (N_15546,N_15359,N_15256);
nor U15547 (N_15547,N_15219,N_15276);
and U15548 (N_15548,N_15237,N_15238);
or U15549 (N_15549,N_15392,N_15351);
nand U15550 (N_15550,N_15363,N_15203);
nand U15551 (N_15551,N_15225,N_15232);
or U15552 (N_15552,N_15206,N_15350);
xor U15553 (N_15553,N_15312,N_15321);
xor U15554 (N_15554,N_15204,N_15350);
and U15555 (N_15555,N_15205,N_15229);
nand U15556 (N_15556,N_15377,N_15364);
and U15557 (N_15557,N_15341,N_15352);
nand U15558 (N_15558,N_15357,N_15376);
or U15559 (N_15559,N_15332,N_15262);
nor U15560 (N_15560,N_15229,N_15348);
nand U15561 (N_15561,N_15347,N_15204);
nand U15562 (N_15562,N_15387,N_15316);
nor U15563 (N_15563,N_15334,N_15206);
or U15564 (N_15564,N_15226,N_15301);
nand U15565 (N_15565,N_15339,N_15369);
or U15566 (N_15566,N_15210,N_15233);
and U15567 (N_15567,N_15289,N_15241);
or U15568 (N_15568,N_15260,N_15321);
or U15569 (N_15569,N_15384,N_15231);
nand U15570 (N_15570,N_15316,N_15399);
and U15571 (N_15571,N_15296,N_15377);
and U15572 (N_15572,N_15280,N_15398);
nor U15573 (N_15573,N_15378,N_15353);
or U15574 (N_15574,N_15294,N_15304);
nand U15575 (N_15575,N_15365,N_15352);
nand U15576 (N_15576,N_15373,N_15282);
nor U15577 (N_15577,N_15207,N_15310);
nor U15578 (N_15578,N_15240,N_15276);
nor U15579 (N_15579,N_15249,N_15374);
nand U15580 (N_15580,N_15367,N_15361);
nand U15581 (N_15581,N_15282,N_15208);
nand U15582 (N_15582,N_15328,N_15356);
xor U15583 (N_15583,N_15391,N_15266);
nor U15584 (N_15584,N_15373,N_15228);
or U15585 (N_15585,N_15379,N_15393);
nor U15586 (N_15586,N_15299,N_15220);
or U15587 (N_15587,N_15238,N_15282);
xor U15588 (N_15588,N_15349,N_15218);
and U15589 (N_15589,N_15358,N_15329);
nor U15590 (N_15590,N_15346,N_15241);
nand U15591 (N_15591,N_15249,N_15336);
nor U15592 (N_15592,N_15211,N_15301);
nor U15593 (N_15593,N_15273,N_15217);
nor U15594 (N_15594,N_15325,N_15258);
nor U15595 (N_15595,N_15313,N_15304);
nor U15596 (N_15596,N_15375,N_15372);
and U15597 (N_15597,N_15386,N_15262);
nor U15598 (N_15598,N_15293,N_15382);
nand U15599 (N_15599,N_15320,N_15277);
or U15600 (N_15600,N_15540,N_15442);
or U15601 (N_15601,N_15534,N_15502);
and U15602 (N_15602,N_15424,N_15452);
or U15603 (N_15603,N_15454,N_15523);
and U15604 (N_15604,N_15538,N_15473);
or U15605 (N_15605,N_15478,N_15574);
or U15606 (N_15606,N_15597,N_15494);
nor U15607 (N_15607,N_15592,N_15566);
nand U15608 (N_15608,N_15510,N_15584);
nor U15609 (N_15609,N_15599,N_15436);
and U15610 (N_15610,N_15570,N_15556);
nor U15611 (N_15611,N_15497,N_15575);
and U15612 (N_15612,N_15480,N_15484);
or U15613 (N_15613,N_15503,N_15524);
nor U15614 (N_15614,N_15460,N_15462);
xnor U15615 (N_15615,N_15578,N_15589);
nor U15616 (N_15616,N_15505,N_15428);
or U15617 (N_15617,N_15451,N_15545);
and U15618 (N_15618,N_15542,N_15509);
nand U15619 (N_15619,N_15506,N_15457);
or U15620 (N_15620,N_15521,N_15400);
nand U15621 (N_15621,N_15409,N_15455);
and U15622 (N_15622,N_15475,N_15583);
or U15623 (N_15623,N_15554,N_15437);
or U15624 (N_15624,N_15486,N_15560);
or U15625 (N_15625,N_15474,N_15432);
and U15626 (N_15626,N_15543,N_15579);
and U15627 (N_15627,N_15552,N_15466);
and U15628 (N_15628,N_15412,N_15580);
and U15629 (N_15629,N_15450,N_15498);
and U15630 (N_15630,N_15553,N_15529);
nand U15631 (N_15631,N_15551,N_15563);
and U15632 (N_15632,N_15535,N_15422);
nor U15633 (N_15633,N_15469,N_15504);
and U15634 (N_15634,N_15585,N_15572);
or U15635 (N_15635,N_15470,N_15407);
and U15636 (N_15636,N_15472,N_15547);
or U15637 (N_15637,N_15453,N_15487);
and U15638 (N_15638,N_15587,N_15573);
nor U15639 (N_15639,N_15515,N_15403);
nor U15640 (N_15640,N_15488,N_15447);
nand U15641 (N_15641,N_15439,N_15448);
nor U15642 (N_15642,N_15525,N_15561);
or U15643 (N_15643,N_15458,N_15519);
and U15644 (N_15644,N_15490,N_15401);
and U15645 (N_15645,N_15415,N_15511);
or U15646 (N_15646,N_15402,N_15500);
nand U15647 (N_15647,N_15434,N_15404);
nand U15648 (N_15648,N_15418,N_15406);
and U15649 (N_15649,N_15531,N_15483);
nand U15650 (N_15650,N_15533,N_15445);
or U15651 (N_15651,N_15517,N_15408);
nor U15652 (N_15652,N_15588,N_15438);
or U15653 (N_15653,N_15586,N_15507);
nand U15654 (N_15654,N_15539,N_15405);
or U15655 (N_15655,N_15512,N_15594);
nand U15656 (N_15656,N_15493,N_15420);
or U15657 (N_15657,N_15444,N_15431);
nand U15658 (N_15658,N_15532,N_15421);
nand U15659 (N_15659,N_15590,N_15443);
xor U15660 (N_15660,N_15426,N_15546);
xnor U15661 (N_15661,N_15598,N_15482);
xor U15662 (N_15662,N_15427,N_15576);
nor U15663 (N_15663,N_15548,N_15537);
nor U15664 (N_15664,N_15564,N_15465);
nor U15665 (N_15665,N_15481,N_15514);
nand U15666 (N_15666,N_15461,N_15430);
nand U15667 (N_15667,N_15520,N_15467);
or U15668 (N_15668,N_15591,N_15558);
and U15669 (N_15669,N_15459,N_15508);
nor U15670 (N_15670,N_15423,N_15516);
or U15671 (N_15671,N_15577,N_15433);
and U15672 (N_15672,N_15562,N_15499);
or U15673 (N_15673,N_15565,N_15569);
nand U15674 (N_15674,N_15571,N_15491);
nor U15675 (N_15675,N_15485,N_15477);
and U15676 (N_15676,N_15446,N_15410);
and U15677 (N_15677,N_15568,N_15581);
and U15678 (N_15678,N_15518,N_15449);
nand U15679 (N_15679,N_15417,N_15522);
nor U15680 (N_15680,N_15567,N_15413);
and U15681 (N_15681,N_15414,N_15550);
or U15682 (N_15682,N_15526,N_15596);
nor U15683 (N_15683,N_15463,N_15527);
nor U15684 (N_15684,N_15440,N_15501);
nand U15685 (N_15685,N_15411,N_15464);
or U15686 (N_15686,N_15513,N_15441);
nand U15687 (N_15687,N_15489,N_15582);
nor U15688 (N_15688,N_15456,N_15496);
nor U15689 (N_15689,N_15541,N_15544);
nor U15690 (N_15690,N_15468,N_15435);
or U15691 (N_15691,N_15479,N_15416);
nor U15692 (N_15692,N_15559,N_15530);
nand U15693 (N_15693,N_15492,N_15476);
nor U15694 (N_15694,N_15536,N_15557);
and U15695 (N_15695,N_15593,N_15549);
nor U15696 (N_15696,N_15471,N_15495);
nand U15697 (N_15697,N_15429,N_15555);
and U15698 (N_15698,N_15528,N_15419);
or U15699 (N_15699,N_15595,N_15425);
nand U15700 (N_15700,N_15561,N_15586);
nand U15701 (N_15701,N_15499,N_15502);
and U15702 (N_15702,N_15453,N_15413);
and U15703 (N_15703,N_15412,N_15509);
nor U15704 (N_15704,N_15521,N_15541);
xor U15705 (N_15705,N_15456,N_15579);
nand U15706 (N_15706,N_15409,N_15458);
nor U15707 (N_15707,N_15468,N_15459);
and U15708 (N_15708,N_15443,N_15515);
nor U15709 (N_15709,N_15463,N_15423);
nor U15710 (N_15710,N_15400,N_15449);
or U15711 (N_15711,N_15559,N_15528);
nand U15712 (N_15712,N_15412,N_15456);
or U15713 (N_15713,N_15499,N_15598);
or U15714 (N_15714,N_15500,N_15497);
nor U15715 (N_15715,N_15447,N_15516);
and U15716 (N_15716,N_15539,N_15484);
nor U15717 (N_15717,N_15480,N_15434);
or U15718 (N_15718,N_15561,N_15456);
xor U15719 (N_15719,N_15458,N_15413);
nand U15720 (N_15720,N_15438,N_15466);
nand U15721 (N_15721,N_15557,N_15457);
nor U15722 (N_15722,N_15518,N_15421);
nand U15723 (N_15723,N_15585,N_15528);
or U15724 (N_15724,N_15576,N_15598);
and U15725 (N_15725,N_15473,N_15544);
and U15726 (N_15726,N_15575,N_15528);
nand U15727 (N_15727,N_15427,N_15450);
or U15728 (N_15728,N_15503,N_15472);
nand U15729 (N_15729,N_15414,N_15470);
or U15730 (N_15730,N_15522,N_15483);
and U15731 (N_15731,N_15588,N_15526);
nor U15732 (N_15732,N_15523,N_15598);
and U15733 (N_15733,N_15557,N_15498);
or U15734 (N_15734,N_15518,N_15459);
or U15735 (N_15735,N_15423,N_15580);
or U15736 (N_15736,N_15535,N_15454);
nor U15737 (N_15737,N_15491,N_15498);
and U15738 (N_15738,N_15434,N_15424);
nand U15739 (N_15739,N_15569,N_15578);
or U15740 (N_15740,N_15595,N_15474);
nand U15741 (N_15741,N_15424,N_15513);
and U15742 (N_15742,N_15411,N_15500);
nand U15743 (N_15743,N_15479,N_15422);
nand U15744 (N_15744,N_15567,N_15425);
or U15745 (N_15745,N_15572,N_15435);
xor U15746 (N_15746,N_15556,N_15525);
and U15747 (N_15747,N_15571,N_15553);
nand U15748 (N_15748,N_15425,N_15452);
or U15749 (N_15749,N_15405,N_15426);
and U15750 (N_15750,N_15588,N_15525);
nand U15751 (N_15751,N_15518,N_15574);
nor U15752 (N_15752,N_15527,N_15477);
nand U15753 (N_15753,N_15522,N_15593);
xnor U15754 (N_15754,N_15564,N_15403);
or U15755 (N_15755,N_15427,N_15433);
or U15756 (N_15756,N_15416,N_15420);
nor U15757 (N_15757,N_15470,N_15406);
and U15758 (N_15758,N_15585,N_15523);
and U15759 (N_15759,N_15453,N_15538);
nor U15760 (N_15760,N_15532,N_15551);
nor U15761 (N_15761,N_15482,N_15589);
nor U15762 (N_15762,N_15430,N_15517);
and U15763 (N_15763,N_15468,N_15575);
nor U15764 (N_15764,N_15527,N_15416);
or U15765 (N_15765,N_15582,N_15552);
and U15766 (N_15766,N_15473,N_15579);
nor U15767 (N_15767,N_15453,N_15435);
nor U15768 (N_15768,N_15592,N_15571);
and U15769 (N_15769,N_15413,N_15533);
or U15770 (N_15770,N_15436,N_15594);
xnor U15771 (N_15771,N_15492,N_15502);
xor U15772 (N_15772,N_15540,N_15515);
nor U15773 (N_15773,N_15570,N_15512);
xnor U15774 (N_15774,N_15530,N_15490);
or U15775 (N_15775,N_15589,N_15549);
or U15776 (N_15776,N_15573,N_15491);
or U15777 (N_15777,N_15476,N_15560);
nor U15778 (N_15778,N_15593,N_15480);
nor U15779 (N_15779,N_15596,N_15423);
nand U15780 (N_15780,N_15444,N_15518);
and U15781 (N_15781,N_15468,N_15471);
or U15782 (N_15782,N_15498,N_15434);
nor U15783 (N_15783,N_15518,N_15587);
nor U15784 (N_15784,N_15549,N_15571);
or U15785 (N_15785,N_15424,N_15462);
and U15786 (N_15786,N_15548,N_15509);
nand U15787 (N_15787,N_15449,N_15450);
nand U15788 (N_15788,N_15574,N_15519);
nand U15789 (N_15789,N_15463,N_15578);
or U15790 (N_15790,N_15424,N_15522);
nor U15791 (N_15791,N_15426,N_15464);
xnor U15792 (N_15792,N_15595,N_15508);
nor U15793 (N_15793,N_15519,N_15553);
nand U15794 (N_15794,N_15482,N_15464);
nor U15795 (N_15795,N_15421,N_15465);
or U15796 (N_15796,N_15518,N_15468);
nor U15797 (N_15797,N_15591,N_15410);
nand U15798 (N_15798,N_15456,N_15452);
and U15799 (N_15799,N_15565,N_15461);
nand U15800 (N_15800,N_15731,N_15671);
nand U15801 (N_15801,N_15786,N_15604);
and U15802 (N_15802,N_15748,N_15762);
nor U15803 (N_15803,N_15780,N_15634);
nand U15804 (N_15804,N_15721,N_15703);
or U15805 (N_15805,N_15701,N_15720);
nor U15806 (N_15806,N_15694,N_15625);
or U15807 (N_15807,N_15702,N_15754);
or U15808 (N_15808,N_15610,N_15718);
nor U15809 (N_15809,N_15799,N_15618);
nand U15810 (N_15810,N_15645,N_15647);
nand U15811 (N_15811,N_15750,N_15656);
nor U15812 (N_15812,N_15752,N_15622);
and U15813 (N_15813,N_15785,N_15707);
or U15814 (N_15814,N_15741,N_15773);
nand U15815 (N_15815,N_15724,N_15766);
nand U15816 (N_15816,N_15690,N_15660);
nor U15817 (N_15817,N_15782,N_15661);
or U15818 (N_15818,N_15640,N_15646);
and U15819 (N_15819,N_15715,N_15742);
and U15820 (N_15820,N_15744,N_15617);
nand U15821 (N_15821,N_15717,N_15793);
nand U15822 (N_15822,N_15686,N_15629);
nor U15823 (N_15823,N_15619,N_15781);
nor U15824 (N_15824,N_15749,N_15601);
and U15825 (N_15825,N_15740,N_15708);
nand U15826 (N_15826,N_15732,N_15638);
nor U15827 (N_15827,N_15735,N_15607);
and U15828 (N_15828,N_15736,N_15776);
and U15829 (N_15829,N_15746,N_15630);
and U15830 (N_15830,N_15758,N_15756);
nand U15831 (N_15831,N_15649,N_15669);
nand U15832 (N_15832,N_15730,N_15757);
or U15833 (N_15833,N_15655,N_15613);
nand U15834 (N_15834,N_15689,N_15612);
and U15835 (N_15835,N_15668,N_15697);
nand U15836 (N_15836,N_15795,N_15695);
nand U15837 (N_15837,N_15779,N_15792);
nor U15838 (N_15838,N_15631,N_15751);
or U15839 (N_15839,N_15719,N_15600);
and U15840 (N_15840,N_15706,N_15674);
xnor U15841 (N_15841,N_15672,N_15771);
and U15842 (N_15842,N_15683,N_15652);
nor U15843 (N_15843,N_15775,N_15783);
nand U15844 (N_15844,N_15737,N_15784);
or U15845 (N_15845,N_15609,N_15624);
nand U15846 (N_15846,N_15699,N_15768);
and U15847 (N_15847,N_15787,N_15663);
or U15848 (N_15848,N_15725,N_15675);
and U15849 (N_15849,N_15658,N_15621);
or U15850 (N_15850,N_15602,N_15777);
nand U15851 (N_15851,N_15769,N_15774);
or U15852 (N_15852,N_15636,N_15680);
or U15853 (N_15853,N_15677,N_15615);
nand U15854 (N_15854,N_15760,N_15653);
or U15855 (N_15855,N_15798,N_15722);
or U15856 (N_15856,N_15767,N_15673);
nor U15857 (N_15857,N_15712,N_15691);
nand U15858 (N_15858,N_15763,N_15778);
nand U15859 (N_15859,N_15709,N_15666);
and U15860 (N_15860,N_15794,N_15791);
or U15861 (N_15861,N_15692,N_15606);
or U15862 (N_15862,N_15698,N_15772);
nor U15863 (N_15863,N_15633,N_15761);
or U15864 (N_15864,N_15679,N_15710);
nor U15865 (N_15865,N_15693,N_15650);
and U15866 (N_15866,N_15665,N_15696);
nand U15867 (N_15867,N_15662,N_15605);
and U15868 (N_15868,N_15685,N_15700);
or U15869 (N_15869,N_15632,N_15644);
nand U15870 (N_15870,N_15733,N_15648);
nand U15871 (N_15871,N_15727,N_15765);
nor U15872 (N_15872,N_15628,N_15635);
and U15873 (N_15873,N_15705,N_15654);
and U15874 (N_15874,N_15711,N_15729);
nor U15875 (N_15875,N_15714,N_15620);
nand U15876 (N_15876,N_15637,N_15688);
nand U15877 (N_15877,N_15678,N_15716);
or U15878 (N_15878,N_15651,N_15726);
nor U15879 (N_15879,N_15639,N_15738);
and U15880 (N_15880,N_15676,N_15614);
nor U15881 (N_15881,N_15684,N_15747);
and U15882 (N_15882,N_15627,N_15641);
nand U15883 (N_15883,N_15704,N_15603);
nand U15884 (N_15884,N_15739,N_15743);
and U15885 (N_15885,N_15659,N_15789);
nand U15886 (N_15886,N_15626,N_15657);
or U15887 (N_15887,N_15797,N_15796);
nor U15888 (N_15888,N_15687,N_15664);
nand U15889 (N_15889,N_15681,N_15790);
nor U15890 (N_15890,N_15788,N_15667);
nor U15891 (N_15891,N_15608,N_15755);
nor U15892 (N_15892,N_15670,N_15611);
nor U15893 (N_15893,N_15642,N_15759);
or U15894 (N_15894,N_15643,N_15723);
and U15895 (N_15895,N_15616,N_15682);
or U15896 (N_15896,N_15764,N_15623);
and U15897 (N_15897,N_15728,N_15734);
nor U15898 (N_15898,N_15770,N_15713);
nor U15899 (N_15899,N_15745,N_15753);
nor U15900 (N_15900,N_15731,N_15747);
or U15901 (N_15901,N_15743,N_15654);
xor U15902 (N_15902,N_15721,N_15657);
nor U15903 (N_15903,N_15613,N_15721);
nand U15904 (N_15904,N_15695,N_15721);
nor U15905 (N_15905,N_15623,N_15711);
nand U15906 (N_15906,N_15637,N_15760);
nand U15907 (N_15907,N_15710,N_15740);
nand U15908 (N_15908,N_15662,N_15627);
or U15909 (N_15909,N_15747,N_15703);
or U15910 (N_15910,N_15682,N_15755);
or U15911 (N_15911,N_15638,N_15686);
nand U15912 (N_15912,N_15772,N_15611);
and U15913 (N_15913,N_15770,N_15644);
or U15914 (N_15914,N_15690,N_15777);
or U15915 (N_15915,N_15675,N_15621);
and U15916 (N_15916,N_15626,N_15715);
nand U15917 (N_15917,N_15703,N_15753);
nor U15918 (N_15918,N_15644,N_15643);
nand U15919 (N_15919,N_15707,N_15694);
and U15920 (N_15920,N_15604,N_15671);
or U15921 (N_15921,N_15684,N_15765);
xnor U15922 (N_15922,N_15614,N_15633);
and U15923 (N_15923,N_15661,N_15670);
nor U15924 (N_15924,N_15704,N_15717);
and U15925 (N_15925,N_15657,N_15740);
or U15926 (N_15926,N_15729,N_15741);
nand U15927 (N_15927,N_15662,N_15609);
or U15928 (N_15928,N_15793,N_15758);
nand U15929 (N_15929,N_15793,N_15786);
nand U15930 (N_15930,N_15774,N_15676);
nor U15931 (N_15931,N_15609,N_15668);
and U15932 (N_15932,N_15637,N_15681);
or U15933 (N_15933,N_15770,N_15668);
and U15934 (N_15934,N_15704,N_15642);
and U15935 (N_15935,N_15627,N_15677);
nand U15936 (N_15936,N_15759,N_15783);
and U15937 (N_15937,N_15670,N_15601);
and U15938 (N_15938,N_15724,N_15628);
nor U15939 (N_15939,N_15761,N_15613);
nand U15940 (N_15940,N_15742,N_15758);
nand U15941 (N_15941,N_15793,N_15773);
and U15942 (N_15942,N_15614,N_15735);
nand U15943 (N_15943,N_15792,N_15703);
or U15944 (N_15944,N_15784,N_15713);
and U15945 (N_15945,N_15655,N_15752);
and U15946 (N_15946,N_15665,N_15662);
or U15947 (N_15947,N_15721,N_15658);
or U15948 (N_15948,N_15658,N_15668);
and U15949 (N_15949,N_15690,N_15630);
nand U15950 (N_15950,N_15617,N_15722);
and U15951 (N_15951,N_15715,N_15675);
xor U15952 (N_15952,N_15617,N_15619);
and U15953 (N_15953,N_15798,N_15795);
nor U15954 (N_15954,N_15656,N_15789);
nor U15955 (N_15955,N_15788,N_15797);
nor U15956 (N_15956,N_15695,N_15746);
or U15957 (N_15957,N_15681,N_15759);
nand U15958 (N_15958,N_15757,N_15657);
nor U15959 (N_15959,N_15729,N_15726);
or U15960 (N_15960,N_15618,N_15792);
nand U15961 (N_15961,N_15725,N_15701);
or U15962 (N_15962,N_15792,N_15629);
and U15963 (N_15963,N_15756,N_15709);
and U15964 (N_15964,N_15613,N_15775);
or U15965 (N_15965,N_15703,N_15659);
and U15966 (N_15966,N_15613,N_15717);
nor U15967 (N_15967,N_15717,N_15685);
nor U15968 (N_15968,N_15664,N_15741);
or U15969 (N_15969,N_15647,N_15768);
or U15970 (N_15970,N_15725,N_15696);
nand U15971 (N_15971,N_15749,N_15605);
and U15972 (N_15972,N_15676,N_15779);
or U15973 (N_15973,N_15666,N_15772);
or U15974 (N_15974,N_15617,N_15775);
nor U15975 (N_15975,N_15688,N_15766);
nor U15976 (N_15976,N_15689,N_15734);
nor U15977 (N_15977,N_15674,N_15724);
and U15978 (N_15978,N_15681,N_15735);
or U15979 (N_15979,N_15671,N_15608);
nand U15980 (N_15980,N_15791,N_15707);
and U15981 (N_15981,N_15782,N_15632);
and U15982 (N_15982,N_15605,N_15797);
or U15983 (N_15983,N_15662,N_15641);
or U15984 (N_15984,N_15798,N_15654);
and U15985 (N_15985,N_15706,N_15630);
nor U15986 (N_15986,N_15640,N_15697);
nand U15987 (N_15987,N_15740,N_15662);
nand U15988 (N_15988,N_15725,N_15740);
nand U15989 (N_15989,N_15673,N_15688);
nor U15990 (N_15990,N_15659,N_15716);
nor U15991 (N_15991,N_15607,N_15642);
and U15992 (N_15992,N_15722,N_15739);
nor U15993 (N_15993,N_15643,N_15703);
and U15994 (N_15994,N_15681,N_15636);
and U15995 (N_15995,N_15652,N_15631);
and U15996 (N_15996,N_15745,N_15640);
nand U15997 (N_15997,N_15765,N_15721);
nor U15998 (N_15998,N_15668,N_15655);
nor U15999 (N_15999,N_15619,N_15761);
and U16000 (N_16000,N_15961,N_15840);
and U16001 (N_16001,N_15920,N_15894);
nor U16002 (N_16002,N_15898,N_15856);
nor U16003 (N_16003,N_15860,N_15835);
nand U16004 (N_16004,N_15883,N_15870);
and U16005 (N_16005,N_15848,N_15949);
or U16006 (N_16006,N_15943,N_15804);
xor U16007 (N_16007,N_15864,N_15983);
nand U16008 (N_16008,N_15993,N_15915);
nor U16009 (N_16009,N_15982,N_15812);
nand U16010 (N_16010,N_15990,N_15985);
or U16011 (N_16011,N_15893,N_15934);
or U16012 (N_16012,N_15865,N_15878);
nor U16013 (N_16013,N_15815,N_15922);
nor U16014 (N_16014,N_15939,N_15823);
nor U16015 (N_16015,N_15813,N_15834);
nor U16016 (N_16016,N_15897,N_15832);
or U16017 (N_16017,N_15821,N_15891);
or U16018 (N_16018,N_15937,N_15968);
and U16019 (N_16019,N_15808,N_15841);
nor U16020 (N_16020,N_15988,N_15839);
nor U16021 (N_16021,N_15805,N_15825);
nand U16022 (N_16022,N_15852,N_15923);
nand U16023 (N_16023,N_15946,N_15999);
xnor U16024 (N_16024,N_15964,N_15828);
or U16025 (N_16025,N_15887,N_15912);
nor U16026 (N_16026,N_15882,N_15998);
or U16027 (N_16027,N_15827,N_15970);
nand U16028 (N_16028,N_15904,N_15969);
nor U16029 (N_16029,N_15986,N_15824);
nor U16030 (N_16030,N_15822,N_15959);
and U16031 (N_16031,N_15933,N_15967);
nand U16032 (N_16032,N_15927,N_15910);
nor U16033 (N_16033,N_15890,N_15908);
nor U16034 (N_16034,N_15972,N_15957);
and U16035 (N_16035,N_15849,N_15948);
nor U16036 (N_16036,N_15863,N_15888);
and U16037 (N_16037,N_15979,N_15976);
or U16038 (N_16038,N_15899,N_15845);
or U16039 (N_16039,N_15900,N_15811);
or U16040 (N_16040,N_15944,N_15809);
nor U16041 (N_16041,N_15886,N_15962);
or U16042 (N_16042,N_15877,N_15911);
and U16043 (N_16043,N_15913,N_15858);
nand U16044 (N_16044,N_15992,N_15838);
and U16045 (N_16045,N_15855,N_15928);
and U16046 (N_16046,N_15989,N_15879);
nand U16047 (N_16047,N_15942,N_15866);
nand U16048 (N_16048,N_15902,N_15956);
or U16049 (N_16049,N_15916,N_15803);
nand U16050 (N_16050,N_15954,N_15884);
nand U16051 (N_16051,N_15874,N_15867);
nor U16052 (N_16052,N_15929,N_15826);
nand U16053 (N_16053,N_15971,N_15925);
xnor U16054 (N_16054,N_15991,N_15862);
nand U16055 (N_16055,N_15966,N_15950);
nand U16056 (N_16056,N_15987,N_15857);
and U16057 (N_16057,N_15918,N_15806);
nor U16058 (N_16058,N_15947,N_15994);
or U16059 (N_16059,N_15958,N_15936);
nor U16060 (N_16060,N_15926,N_15873);
or U16061 (N_16061,N_15802,N_15940);
and U16062 (N_16062,N_15833,N_15901);
or U16063 (N_16063,N_15931,N_15980);
nand U16064 (N_16064,N_15816,N_15847);
and U16065 (N_16065,N_15871,N_15881);
nor U16066 (N_16066,N_15850,N_15817);
nor U16067 (N_16067,N_15820,N_15896);
nand U16068 (N_16068,N_15963,N_15861);
and U16069 (N_16069,N_15975,N_15889);
nand U16070 (N_16070,N_15875,N_15914);
or U16071 (N_16071,N_15917,N_15938);
and U16072 (N_16072,N_15869,N_15810);
or U16073 (N_16073,N_15844,N_15930);
nor U16074 (N_16074,N_15932,N_15924);
nand U16075 (N_16075,N_15831,N_15995);
or U16076 (N_16076,N_15872,N_15801);
or U16077 (N_16077,N_15996,N_15903);
nor U16078 (N_16078,N_15907,N_15905);
and U16079 (N_16079,N_15868,N_15851);
nand U16080 (N_16080,N_15814,N_15830);
and U16081 (N_16081,N_15836,N_15941);
or U16082 (N_16082,N_15977,N_15895);
nor U16083 (N_16083,N_15965,N_15921);
nand U16084 (N_16084,N_15997,N_15974);
or U16085 (N_16085,N_15906,N_15955);
nor U16086 (N_16086,N_15978,N_15885);
nand U16087 (N_16087,N_15945,N_15837);
or U16088 (N_16088,N_15973,N_15818);
xnor U16089 (N_16089,N_15880,N_15807);
or U16090 (N_16090,N_15951,N_15919);
nor U16091 (N_16091,N_15952,N_15859);
and U16092 (N_16092,N_15876,N_15960);
or U16093 (N_16093,N_15984,N_15854);
and U16094 (N_16094,N_15892,N_15981);
or U16095 (N_16095,N_15953,N_15842);
or U16096 (N_16096,N_15843,N_15800);
or U16097 (N_16097,N_15819,N_15853);
or U16098 (N_16098,N_15909,N_15846);
nor U16099 (N_16099,N_15829,N_15935);
nand U16100 (N_16100,N_15823,N_15947);
or U16101 (N_16101,N_15958,N_15872);
nor U16102 (N_16102,N_15979,N_15800);
or U16103 (N_16103,N_15920,N_15838);
and U16104 (N_16104,N_15953,N_15827);
or U16105 (N_16105,N_15868,N_15937);
nor U16106 (N_16106,N_15821,N_15857);
nor U16107 (N_16107,N_15877,N_15867);
and U16108 (N_16108,N_15915,N_15982);
or U16109 (N_16109,N_15973,N_15952);
nand U16110 (N_16110,N_15827,N_15877);
nor U16111 (N_16111,N_15933,N_15961);
nand U16112 (N_16112,N_15935,N_15802);
or U16113 (N_16113,N_15872,N_15834);
and U16114 (N_16114,N_15880,N_15908);
nor U16115 (N_16115,N_15951,N_15870);
or U16116 (N_16116,N_15927,N_15963);
and U16117 (N_16117,N_15847,N_15877);
and U16118 (N_16118,N_15877,N_15849);
xnor U16119 (N_16119,N_15802,N_15803);
and U16120 (N_16120,N_15914,N_15973);
and U16121 (N_16121,N_15864,N_15973);
nand U16122 (N_16122,N_15844,N_15819);
xor U16123 (N_16123,N_15850,N_15845);
nand U16124 (N_16124,N_15843,N_15938);
or U16125 (N_16125,N_15850,N_15980);
xnor U16126 (N_16126,N_15964,N_15960);
nand U16127 (N_16127,N_15808,N_15845);
and U16128 (N_16128,N_15858,N_15827);
xnor U16129 (N_16129,N_15845,N_15971);
and U16130 (N_16130,N_15873,N_15885);
nor U16131 (N_16131,N_15996,N_15989);
or U16132 (N_16132,N_15944,N_15841);
nand U16133 (N_16133,N_15858,N_15840);
nand U16134 (N_16134,N_15966,N_15868);
or U16135 (N_16135,N_15870,N_15899);
nor U16136 (N_16136,N_15865,N_15807);
nand U16137 (N_16137,N_15988,N_15941);
nand U16138 (N_16138,N_15980,N_15893);
or U16139 (N_16139,N_15862,N_15830);
nand U16140 (N_16140,N_15924,N_15861);
xor U16141 (N_16141,N_15848,N_15920);
or U16142 (N_16142,N_15837,N_15976);
nand U16143 (N_16143,N_15998,N_15917);
or U16144 (N_16144,N_15848,N_15842);
nor U16145 (N_16145,N_15978,N_15907);
nand U16146 (N_16146,N_15912,N_15957);
nand U16147 (N_16147,N_15807,N_15889);
or U16148 (N_16148,N_15966,N_15805);
nor U16149 (N_16149,N_15827,N_15874);
or U16150 (N_16150,N_15989,N_15807);
and U16151 (N_16151,N_15879,N_15830);
and U16152 (N_16152,N_15839,N_15928);
nor U16153 (N_16153,N_15825,N_15928);
or U16154 (N_16154,N_15872,N_15922);
nor U16155 (N_16155,N_15858,N_15940);
or U16156 (N_16156,N_15925,N_15852);
and U16157 (N_16157,N_15862,N_15805);
or U16158 (N_16158,N_15970,N_15853);
or U16159 (N_16159,N_15899,N_15800);
and U16160 (N_16160,N_15943,N_15839);
nand U16161 (N_16161,N_15823,N_15840);
nand U16162 (N_16162,N_15962,N_15929);
or U16163 (N_16163,N_15859,N_15899);
and U16164 (N_16164,N_15811,N_15809);
and U16165 (N_16165,N_15935,N_15800);
nand U16166 (N_16166,N_15961,N_15834);
nor U16167 (N_16167,N_15995,N_15955);
nor U16168 (N_16168,N_15821,N_15983);
nor U16169 (N_16169,N_15871,N_15873);
nor U16170 (N_16170,N_15824,N_15906);
nor U16171 (N_16171,N_15880,N_15848);
nand U16172 (N_16172,N_15979,N_15813);
or U16173 (N_16173,N_15900,N_15931);
or U16174 (N_16174,N_15984,N_15880);
and U16175 (N_16175,N_15909,N_15897);
nand U16176 (N_16176,N_15805,N_15998);
xnor U16177 (N_16177,N_15819,N_15964);
nor U16178 (N_16178,N_15983,N_15860);
xor U16179 (N_16179,N_15930,N_15842);
or U16180 (N_16180,N_15975,N_15827);
and U16181 (N_16181,N_15974,N_15840);
or U16182 (N_16182,N_15897,N_15953);
or U16183 (N_16183,N_15870,N_15864);
and U16184 (N_16184,N_15855,N_15879);
nand U16185 (N_16185,N_15985,N_15861);
nand U16186 (N_16186,N_15966,N_15876);
nand U16187 (N_16187,N_15896,N_15818);
nand U16188 (N_16188,N_15873,N_15929);
and U16189 (N_16189,N_15912,N_15888);
or U16190 (N_16190,N_15887,N_15813);
and U16191 (N_16191,N_15910,N_15978);
and U16192 (N_16192,N_15825,N_15803);
nand U16193 (N_16193,N_15806,N_15821);
nand U16194 (N_16194,N_15967,N_15953);
nor U16195 (N_16195,N_15996,N_15962);
nor U16196 (N_16196,N_15901,N_15844);
nand U16197 (N_16197,N_15942,N_15828);
or U16198 (N_16198,N_15851,N_15830);
nor U16199 (N_16199,N_15960,N_15968);
or U16200 (N_16200,N_16147,N_16089);
and U16201 (N_16201,N_16059,N_16071);
and U16202 (N_16202,N_16024,N_16053);
or U16203 (N_16203,N_16061,N_16079);
and U16204 (N_16204,N_16066,N_16078);
and U16205 (N_16205,N_16149,N_16070);
nand U16206 (N_16206,N_16092,N_16174);
or U16207 (N_16207,N_16158,N_16123);
or U16208 (N_16208,N_16075,N_16102);
nand U16209 (N_16209,N_16140,N_16197);
and U16210 (N_16210,N_16035,N_16036);
and U16211 (N_16211,N_16116,N_16108);
and U16212 (N_16212,N_16050,N_16088);
nand U16213 (N_16213,N_16172,N_16192);
nand U16214 (N_16214,N_16196,N_16187);
or U16215 (N_16215,N_16160,N_16083);
nand U16216 (N_16216,N_16132,N_16150);
or U16217 (N_16217,N_16073,N_16182);
xnor U16218 (N_16218,N_16011,N_16098);
and U16219 (N_16219,N_16085,N_16032);
and U16220 (N_16220,N_16020,N_16183);
nor U16221 (N_16221,N_16159,N_16090);
or U16222 (N_16222,N_16166,N_16042);
or U16223 (N_16223,N_16016,N_16003);
nand U16224 (N_16224,N_16169,N_16189);
or U16225 (N_16225,N_16179,N_16076);
nand U16226 (N_16226,N_16163,N_16162);
nor U16227 (N_16227,N_16046,N_16057);
and U16228 (N_16228,N_16062,N_16007);
nand U16229 (N_16229,N_16101,N_16081);
and U16230 (N_16230,N_16063,N_16038);
or U16231 (N_16231,N_16154,N_16068);
or U16232 (N_16232,N_16039,N_16188);
or U16233 (N_16233,N_16137,N_16195);
or U16234 (N_16234,N_16190,N_16069);
nor U16235 (N_16235,N_16018,N_16129);
nor U16236 (N_16236,N_16049,N_16152);
and U16237 (N_16237,N_16146,N_16009);
xnor U16238 (N_16238,N_16047,N_16131);
and U16239 (N_16239,N_16161,N_16110);
or U16240 (N_16240,N_16151,N_16033);
or U16241 (N_16241,N_16013,N_16012);
or U16242 (N_16242,N_16103,N_16014);
nor U16243 (N_16243,N_16099,N_16074);
nor U16244 (N_16244,N_16043,N_16128);
nand U16245 (N_16245,N_16113,N_16023);
nor U16246 (N_16246,N_16127,N_16026);
and U16247 (N_16247,N_16028,N_16055);
nand U16248 (N_16248,N_16142,N_16115);
or U16249 (N_16249,N_16177,N_16109);
or U16250 (N_16250,N_16048,N_16082);
and U16251 (N_16251,N_16040,N_16126);
xor U16252 (N_16252,N_16100,N_16145);
or U16253 (N_16253,N_16155,N_16120);
nand U16254 (N_16254,N_16060,N_16045);
nand U16255 (N_16255,N_16135,N_16095);
or U16256 (N_16256,N_16105,N_16119);
nand U16257 (N_16257,N_16117,N_16176);
nand U16258 (N_16258,N_16054,N_16025);
or U16259 (N_16259,N_16017,N_16037);
nand U16260 (N_16260,N_16136,N_16121);
nor U16261 (N_16261,N_16198,N_16193);
or U16262 (N_16262,N_16164,N_16156);
nand U16263 (N_16263,N_16093,N_16171);
and U16264 (N_16264,N_16141,N_16134);
nand U16265 (N_16265,N_16001,N_16157);
or U16266 (N_16266,N_16096,N_16000);
nor U16267 (N_16267,N_16087,N_16165);
nand U16268 (N_16268,N_16084,N_16153);
and U16269 (N_16269,N_16184,N_16006);
nor U16270 (N_16270,N_16072,N_16168);
and U16271 (N_16271,N_16077,N_16138);
and U16272 (N_16272,N_16029,N_16091);
or U16273 (N_16273,N_16104,N_16064);
or U16274 (N_16274,N_16031,N_16086);
nand U16275 (N_16275,N_16094,N_16056);
nor U16276 (N_16276,N_16170,N_16005);
nor U16277 (N_16277,N_16058,N_16139);
nor U16278 (N_16278,N_16122,N_16180);
nand U16279 (N_16279,N_16178,N_16044);
or U16280 (N_16280,N_16027,N_16041);
nor U16281 (N_16281,N_16052,N_16004);
or U16282 (N_16282,N_16065,N_16124);
nand U16283 (N_16283,N_16191,N_16010);
nand U16284 (N_16284,N_16051,N_16002);
nand U16285 (N_16285,N_16067,N_16143);
and U16286 (N_16286,N_16106,N_16022);
nor U16287 (N_16287,N_16080,N_16173);
or U16288 (N_16288,N_16097,N_16034);
and U16289 (N_16289,N_16186,N_16008);
nor U16290 (N_16290,N_16015,N_16185);
nand U16291 (N_16291,N_16167,N_16130);
nor U16292 (N_16292,N_16107,N_16114);
nor U16293 (N_16293,N_16111,N_16112);
and U16294 (N_16294,N_16181,N_16133);
nor U16295 (N_16295,N_16199,N_16118);
and U16296 (N_16296,N_16030,N_16125);
and U16297 (N_16297,N_16021,N_16144);
nor U16298 (N_16298,N_16148,N_16194);
or U16299 (N_16299,N_16175,N_16019);
and U16300 (N_16300,N_16037,N_16028);
or U16301 (N_16301,N_16129,N_16191);
and U16302 (N_16302,N_16083,N_16119);
nand U16303 (N_16303,N_16144,N_16067);
nand U16304 (N_16304,N_16174,N_16000);
and U16305 (N_16305,N_16035,N_16153);
or U16306 (N_16306,N_16104,N_16157);
and U16307 (N_16307,N_16176,N_16009);
nor U16308 (N_16308,N_16124,N_16014);
or U16309 (N_16309,N_16057,N_16151);
or U16310 (N_16310,N_16074,N_16039);
nand U16311 (N_16311,N_16135,N_16100);
or U16312 (N_16312,N_16005,N_16003);
nand U16313 (N_16313,N_16110,N_16073);
and U16314 (N_16314,N_16012,N_16067);
or U16315 (N_16315,N_16045,N_16199);
and U16316 (N_16316,N_16069,N_16181);
nand U16317 (N_16317,N_16111,N_16002);
and U16318 (N_16318,N_16091,N_16001);
and U16319 (N_16319,N_16176,N_16161);
and U16320 (N_16320,N_16133,N_16139);
and U16321 (N_16321,N_16108,N_16122);
xnor U16322 (N_16322,N_16145,N_16143);
nor U16323 (N_16323,N_16025,N_16111);
nor U16324 (N_16324,N_16056,N_16006);
or U16325 (N_16325,N_16039,N_16114);
nand U16326 (N_16326,N_16156,N_16170);
and U16327 (N_16327,N_16171,N_16004);
and U16328 (N_16328,N_16041,N_16091);
or U16329 (N_16329,N_16081,N_16108);
nor U16330 (N_16330,N_16166,N_16087);
or U16331 (N_16331,N_16092,N_16190);
nand U16332 (N_16332,N_16054,N_16111);
and U16333 (N_16333,N_16120,N_16122);
nand U16334 (N_16334,N_16171,N_16140);
or U16335 (N_16335,N_16008,N_16058);
nor U16336 (N_16336,N_16098,N_16039);
nand U16337 (N_16337,N_16075,N_16107);
or U16338 (N_16338,N_16146,N_16025);
nand U16339 (N_16339,N_16070,N_16058);
nor U16340 (N_16340,N_16006,N_16093);
or U16341 (N_16341,N_16051,N_16153);
and U16342 (N_16342,N_16183,N_16152);
or U16343 (N_16343,N_16050,N_16119);
or U16344 (N_16344,N_16087,N_16041);
nand U16345 (N_16345,N_16196,N_16170);
and U16346 (N_16346,N_16185,N_16172);
and U16347 (N_16347,N_16189,N_16185);
nand U16348 (N_16348,N_16190,N_16009);
nor U16349 (N_16349,N_16094,N_16009);
or U16350 (N_16350,N_16188,N_16100);
nand U16351 (N_16351,N_16166,N_16099);
nor U16352 (N_16352,N_16133,N_16164);
or U16353 (N_16353,N_16017,N_16143);
nor U16354 (N_16354,N_16036,N_16187);
and U16355 (N_16355,N_16058,N_16180);
and U16356 (N_16356,N_16174,N_16182);
nand U16357 (N_16357,N_16001,N_16150);
and U16358 (N_16358,N_16165,N_16190);
or U16359 (N_16359,N_16170,N_16127);
and U16360 (N_16360,N_16081,N_16116);
and U16361 (N_16361,N_16137,N_16154);
nor U16362 (N_16362,N_16015,N_16190);
or U16363 (N_16363,N_16120,N_16066);
or U16364 (N_16364,N_16065,N_16087);
nand U16365 (N_16365,N_16197,N_16061);
or U16366 (N_16366,N_16034,N_16179);
nand U16367 (N_16367,N_16150,N_16153);
or U16368 (N_16368,N_16197,N_16074);
or U16369 (N_16369,N_16178,N_16184);
and U16370 (N_16370,N_16026,N_16007);
and U16371 (N_16371,N_16043,N_16007);
and U16372 (N_16372,N_16056,N_16180);
or U16373 (N_16373,N_16117,N_16081);
and U16374 (N_16374,N_16141,N_16008);
nor U16375 (N_16375,N_16098,N_16091);
or U16376 (N_16376,N_16136,N_16127);
or U16377 (N_16377,N_16010,N_16130);
and U16378 (N_16378,N_16059,N_16190);
and U16379 (N_16379,N_16174,N_16169);
nor U16380 (N_16380,N_16087,N_16167);
nand U16381 (N_16381,N_16174,N_16101);
nor U16382 (N_16382,N_16165,N_16065);
or U16383 (N_16383,N_16090,N_16055);
nor U16384 (N_16384,N_16054,N_16192);
nor U16385 (N_16385,N_16174,N_16115);
xor U16386 (N_16386,N_16115,N_16013);
nor U16387 (N_16387,N_16047,N_16012);
and U16388 (N_16388,N_16018,N_16033);
nand U16389 (N_16389,N_16149,N_16047);
and U16390 (N_16390,N_16045,N_16034);
and U16391 (N_16391,N_16047,N_16104);
nand U16392 (N_16392,N_16122,N_16119);
and U16393 (N_16393,N_16064,N_16126);
xor U16394 (N_16394,N_16119,N_16062);
nor U16395 (N_16395,N_16021,N_16029);
nor U16396 (N_16396,N_16173,N_16047);
nand U16397 (N_16397,N_16154,N_16151);
or U16398 (N_16398,N_16011,N_16185);
or U16399 (N_16399,N_16185,N_16068);
and U16400 (N_16400,N_16202,N_16373);
or U16401 (N_16401,N_16279,N_16245);
nor U16402 (N_16402,N_16285,N_16203);
nor U16403 (N_16403,N_16378,N_16208);
and U16404 (N_16404,N_16253,N_16316);
nand U16405 (N_16405,N_16352,N_16290);
or U16406 (N_16406,N_16367,N_16201);
nor U16407 (N_16407,N_16219,N_16206);
nand U16408 (N_16408,N_16260,N_16377);
nand U16409 (N_16409,N_16358,N_16235);
nand U16410 (N_16410,N_16293,N_16212);
or U16411 (N_16411,N_16281,N_16226);
nand U16412 (N_16412,N_16356,N_16240);
nand U16413 (N_16413,N_16259,N_16372);
nand U16414 (N_16414,N_16343,N_16286);
or U16415 (N_16415,N_16315,N_16318);
nor U16416 (N_16416,N_16241,N_16230);
nand U16417 (N_16417,N_16351,N_16247);
nor U16418 (N_16418,N_16228,N_16232);
nor U16419 (N_16419,N_16234,N_16225);
and U16420 (N_16420,N_16283,N_16313);
and U16421 (N_16421,N_16252,N_16256);
nand U16422 (N_16422,N_16340,N_16391);
or U16423 (N_16423,N_16324,N_16380);
nand U16424 (N_16424,N_16217,N_16389);
and U16425 (N_16425,N_16331,N_16242);
and U16426 (N_16426,N_16332,N_16221);
nand U16427 (N_16427,N_16271,N_16238);
and U16428 (N_16428,N_16334,N_16394);
and U16429 (N_16429,N_16254,N_16353);
or U16430 (N_16430,N_16268,N_16323);
and U16431 (N_16431,N_16326,N_16295);
and U16432 (N_16432,N_16258,N_16213);
or U16433 (N_16433,N_16303,N_16248);
nor U16434 (N_16434,N_16220,N_16388);
and U16435 (N_16435,N_16306,N_16250);
nor U16436 (N_16436,N_16344,N_16282);
and U16437 (N_16437,N_16223,N_16210);
or U16438 (N_16438,N_16320,N_16297);
nor U16439 (N_16439,N_16347,N_16349);
and U16440 (N_16440,N_16298,N_16299);
or U16441 (N_16441,N_16305,N_16255);
nor U16442 (N_16442,N_16335,N_16207);
nor U16443 (N_16443,N_16276,N_16222);
nor U16444 (N_16444,N_16392,N_16257);
or U16445 (N_16445,N_16355,N_16224);
nor U16446 (N_16446,N_16327,N_16251);
nand U16447 (N_16447,N_16287,N_16288);
and U16448 (N_16448,N_16272,N_16277);
nor U16449 (N_16449,N_16379,N_16244);
nand U16450 (N_16450,N_16291,N_16311);
or U16451 (N_16451,N_16322,N_16381);
and U16452 (N_16452,N_16264,N_16270);
nand U16453 (N_16453,N_16375,N_16374);
and U16454 (N_16454,N_16399,N_16205);
nand U16455 (N_16455,N_16227,N_16312);
xnor U16456 (N_16456,N_16246,N_16273);
and U16457 (N_16457,N_16300,N_16229);
nand U16458 (N_16458,N_16302,N_16215);
and U16459 (N_16459,N_16301,N_16216);
or U16460 (N_16460,N_16289,N_16231);
or U16461 (N_16461,N_16393,N_16341);
nand U16462 (N_16462,N_16274,N_16346);
nand U16463 (N_16463,N_16348,N_16280);
and U16464 (N_16464,N_16370,N_16304);
nand U16465 (N_16465,N_16266,N_16360);
nor U16466 (N_16466,N_16292,N_16368);
nor U16467 (N_16467,N_16396,N_16328);
nor U16468 (N_16468,N_16321,N_16294);
and U16469 (N_16469,N_16211,N_16239);
or U16470 (N_16470,N_16317,N_16267);
xnor U16471 (N_16471,N_16329,N_16354);
nor U16472 (N_16472,N_16269,N_16383);
and U16473 (N_16473,N_16345,N_16233);
or U16474 (N_16474,N_16236,N_16218);
xnor U16475 (N_16475,N_16390,N_16386);
nor U16476 (N_16476,N_16309,N_16308);
or U16477 (N_16477,N_16278,N_16371);
and U16478 (N_16478,N_16366,N_16249);
nor U16479 (N_16479,N_16284,N_16263);
nand U16480 (N_16480,N_16314,N_16369);
or U16481 (N_16481,N_16200,N_16397);
nand U16482 (N_16482,N_16376,N_16204);
nor U16483 (N_16483,N_16243,N_16319);
or U16484 (N_16484,N_16330,N_16307);
nand U16485 (N_16485,N_16395,N_16336);
and U16486 (N_16486,N_16361,N_16364);
nor U16487 (N_16487,N_16333,N_16398);
xnor U16488 (N_16488,N_16296,N_16363);
nor U16489 (N_16489,N_16357,N_16382);
nand U16490 (N_16490,N_16337,N_16342);
nand U16491 (N_16491,N_16384,N_16275);
nand U16492 (N_16492,N_16214,N_16310);
xnor U16493 (N_16493,N_16385,N_16265);
or U16494 (N_16494,N_16237,N_16350);
nor U16495 (N_16495,N_16325,N_16359);
or U16496 (N_16496,N_16261,N_16339);
nor U16497 (N_16497,N_16209,N_16362);
nand U16498 (N_16498,N_16262,N_16387);
and U16499 (N_16499,N_16338,N_16365);
nand U16500 (N_16500,N_16325,N_16218);
and U16501 (N_16501,N_16321,N_16201);
xor U16502 (N_16502,N_16308,N_16377);
nor U16503 (N_16503,N_16260,N_16348);
or U16504 (N_16504,N_16385,N_16353);
or U16505 (N_16505,N_16343,N_16296);
or U16506 (N_16506,N_16276,N_16363);
nand U16507 (N_16507,N_16398,N_16259);
or U16508 (N_16508,N_16206,N_16205);
and U16509 (N_16509,N_16279,N_16261);
nor U16510 (N_16510,N_16263,N_16281);
nand U16511 (N_16511,N_16235,N_16292);
nor U16512 (N_16512,N_16271,N_16281);
nand U16513 (N_16513,N_16306,N_16249);
nor U16514 (N_16514,N_16286,N_16346);
nor U16515 (N_16515,N_16305,N_16225);
and U16516 (N_16516,N_16292,N_16342);
nand U16517 (N_16517,N_16223,N_16392);
or U16518 (N_16518,N_16382,N_16291);
nand U16519 (N_16519,N_16295,N_16331);
nor U16520 (N_16520,N_16357,N_16244);
and U16521 (N_16521,N_16211,N_16351);
or U16522 (N_16522,N_16297,N_16334);
and U16523 (N_16523,N_16359,N_16399);
nand U16524 (N_16524,N_16211,N_16299);
nand U16525 (N_16525,N_16243,N_16233);
or U16526 (N_16526,N_16387,N_16358);
nor U16527 (N_16527,N_16203,N_16310);
or U16528 (N_16528,N_16218,N_16372);
xnor U16529 (N_16529,N_16304,N_16390);
or U16530 (N_16530,N_16321,N_16208);
nor U16531 (N_16531,N_16217,N_16258);
or U16532 (N_16532,N_16381,N_16284);
nand U16533 (N_16533,N_16247,N_16385);
nand U16534 (N_16534,N_16287,N_16277);
or U16535 (N_16535,N_16352,N_16258);
nand U16536 (N_16536,N_16268,N_16259);
nand U16537 (N_16537,N_16209,N_16222);
or U16538 (N_16538,N_16239,N_16225);
nor U16539 (N_16539,N_16279,N_16366);
nand U16540 (N_16540,N_16382,N_16385);
and U16541 (N_16541,N_16256,N_16248);
nor U16542 (N_16542,N_16242,N_16266);
nand U16543 (N_16543,N_16284,N_16252);
or U16544 (N_16544,N_16292,N_16328);
nor U16545 (N_16545,N_16210,N_16238);
nor U16546 (N_16546,N_16315,N_16214);
nor U16547 (N_16547,N_16327,N_16205);
nor U16548 (N_16548,N_16232,N_16352);
nor U16549 (N_16549,N_16372,N_16264);
and U16550 (N_16550,N_16204,N_16371);
nand U16551 (N_16551,N_16233,N_16289);
nand U16552 (N_16552,N_16317,N_16351);
and U16553 (N_16553,N_16313,N_16235);
nor U16554 (N_16554,N_16298,N_16386);
and U16555 (N_16555,N_16210,N_16349);
or U16556 (N_16556,N_16222,N_16233);
and U16557 (N_16557,N_16308,N_16284);
or U16558 (N_16558,N_16214,N_16286);
and U16559 (N_16559,N_16308,N_16399);
or U16560 (N_16560,N_16380,N_16201);
nand U16561 (N_16561,N_16242,N_16396);
nor U16562 (N_16562,N_16271,N_16351);
or U16563 (N_16563,N_16245,N_16217);
nor U16564 (N_16564,N_16290,N_16216);
nor U16565 (N_16565,N_16390,N_16291);
nand U16566 (N_16566,N_16337,N_16399);
and U16567 (N_16567,N_16240,N_16385);
or U16568 (N_16568,N_16340,N_16384);
or U16569 (N_16569,N_16284,N_16343);
or U16570 (N_16570,N_16360,N_16361);
and U16571 (N_16571,N_16340,N_16326);
nand U16572 (N_16572,N_16390,N_16350);
nand U16573 (N_16573,N_16346,N_16225);
and U16574 (N_16574,N_16217,N_16220);
nor U16575 (N_16575,N_16385,N_16386);
nand U16576 (N_16576,N_16227,N_16325);
nor U16577 (N_16577,N_16313,N_16286);
xnor U16578 (N_16578,N_16342,N_16329);
nand U16579 (N_16579,N_16327,N_16238);
nand U16580 (N_16580,N_16291,N_16375);
and U16581 (N_16581,N_16236,N_16373);
nor U16582 (N_16582,N_16372,N_16393);
or U16583 (N_16583,N_16389,N_16351);
or U16584 (N_16584,N_16278,N_16204);
and U16585 (N_16585,N_16211,N_16274);
or U16586 (N_16586,N_16262,N_16331);
nor U16587 (N_16587,N_16303,N_16301);
or U16588 (N_16588,N_16235,N_16237);
and U16589 (N_16589,N_16299,N_16350);
or U16590 (N_16590,N_16318,N_16248);
nand U16591 (N_16591,N_16335,N_16328);
and U16592 (N_16592,N_16300,N_16385);
and U16593 (N_16593,N_16397,N_16380);
or U16594 (N_16594,N_16341,N_16306);
or U16595 (N_16595,N_16272,N_16240);
nand U16596 (N_16596,N_16364,N_16308);
nor U16597 (N_16597,N_16313,N_16259);
nor U16598 (N_16598,N_16285,N_16296);
or U16599 (N_16599,N_16336,N_16249);
and U16600 (N_16600,N_16590,N_16477);
nand U16601 (N_16601,N_16456,N_16445);
or U16602 (N_16602,N_16546,N_16582);
or U16603 (N_16603,N_16431,N_16522);
nand U16604 (N_16604,N_16547,N_16491);
nand U16605 (N_16605,N_16432,N_16427);
nand U16606 (N_16606,N_16455,N_16468);
nor U16607 (N_16607,N_16458,N_16441);
or U16608 (N_16608,N_16406,N_16413);
or U16609 (N_16609,N_16443,N_16426);
and U16610 (N_16610,N_16503,N_16478);
and U16611 (N_16611,N_16452,N_16595);
nor U16612 (N_16612,N_16552,N_16417);
nor U16613 (N_16613,N_16531,N_16580);
or U16614 (N_16614,N_16402,N_16557);
nor U16615 (N_16615,N_16558,N_16579);
or U16616 (N_16616,N_16492,N_16533);
or U16617 (N_16617,N_16471,N_16520);
nand U16618 (N_16618,N_16586,N_16514);
nor U16619 (N_16619,N_16424,N_16448);
or U16620 (N_16620,N_16501,N_16504);
nor U16621 (N_16621,N_16559,N_16566);
and U16622 (N_16622,N_16457,N_16493);
nand U16623 (N_16623,N_16572,N_16551);
and U16624 (N_16624,N_16485,N_16447);
and U16625 (N_16625,N_16555,N_16506);
and U16626 (N_16626,N_16470,N_16516);
and U16627 (N_16627,N_16488,N_16513);
nand U16628 (N_16628,N_16562,N_16460);
or U16629 (N_16629,N_16404,N_16518);
nor U16630 (N_16630,N_16573,N_16553);
and U16631 (N_16631,N_16400,N_16544);
nor U16632 (N_16632,N_16484,N_16490);
nand U16633 (N_16633,N_16411,N_16405);
nand U16634 (N_16634,N_16463,N_16569);
and U16635 (N_16635,N_16494,N_16565);
nor U16636 (N_16636,N_16592,N_16540);
nand U16637 (N_16637,N_16534,N_16473);
nand U16638 (N_16638,N_16549,N_16451);
or U16639 (N_16639,N_16548,N_16422);
and U16640 (N_16640,N_16521,N_16560);
or U16641 (N_16641,N_16510,N_16556);
or U16642 (N_16642,N_16438,N_16433);
and U16643 (N_16643,N_16482,N_16483);
and U16644 (N_16644,N_16589,N_16428);
and U16645 (N_16645,N_16597,N_16571);
or U16646 (N_16646,N_16583,N_16529);
xor U16647 (N_16647,N_16416,N_16541);
nand U16648 (N_16648,N_16496,N_16511);
and U16649 (N_16649,N_16576,N_16436);
and U16650 (N_16650,N_16498,N_16434);
nor U16651 (N_16651,N_16591,N_16430);
or U16652 (N_16652,N_16593,N_16536);
or U16653 (N_16653,N_16495,N_16554);
nand U16654 (N_16654,N_16542,N_16585);
nor U16655 (N_16655,N_16418,N_16538);
and U16656 (N_16656,N_16412,N_16587);
or U16657 (N_16657,N_16479,N_16570);
nand U16658 (N_16658,N_16505,N_16440);
nor U16659 (N_16659,N_16454,N_16599);
or U16660 (N_16660,N_16453,N_16575);
and U16661 (N_16661,N_16588,N_16469);
nand U16662 (N_16662,N_16528,N_16466);
nor U16663 (N_16663,N_16461,N_16439);
nor U16664 (N_16664,N_16499,N_16574);
or U16665 (N_16665,N_16497,N_16474);
nand U16666 (N_16666,N_16450,N_16435);
or U16667 (N_16667,N_16421,N_16480);
and U16668 (N_16668,N_16486,N_16446);
nor U16669 (N_16669,N_16408,N_16517);
and U16670 (N_16670,N_16596,N_16410);
and U16671 (N_16671,N_16442,N_16415);
or U16672 (N_16672,N_16507,N_16568);
or U16673 (N_16673,N_16459,N_16532);
and U16674 (N_16674,N_16567,N_16509);
or U16675 (N_16675,N_16444,N_16578);
nand U16676 (N_16676,N_16425,N_16437);
nand U16677 (N_16677,N_16563,N_16526);
nand U16678 (N_16678,N_16512,N_16407);
or U16679 (N_16679,N_16481,N_16423);
and U16680 (N_16680,N_16527,N_16598);
nor U16681 (N_16681,N_16476,N_16594);
nand U16682 (N_16682,N_16414,N_16543);
nand U16683 (N_16683,N_16524,N_16401);
nor U16684 (N_16684,N_16584,N_16561);
nor U16685 (N_16685,N_16472,N_16409);
and U16686 (N_16686,N_16465,N_16564);
and U16687 (N_16687,N_16467,N_16539);
nor U16688 (N_16688,N_16535,N_16487);
nand U16689 (N_16689,N_16449,N_16419);
or U16690 (N_16690,N_16429,N_16537);
nor U16691 (N_16691,N_16525,N_16508);
or U16692 (N_16692,N_16515,N_16519);
and U16693 (N_16693,N_16464,N_16581);
and U16694 (N_16694,N_16530,N_16500);
xor U16695 (N_16695,N_16420,N_16550);
nor U16696 (N_16696,N_16489,N_16523);
nand U16697 (N_16697,N_16545,N_16475);
nor U16698 (N_16698,N_16577,N_16502);
and U16699 (N_16699,N_16403,N_16462);
nor U16700 (N_16700,N_16411,N_16557);
nor U16701 (N_16701,N_16536,N_16414);
nor U16702 (N_16702,N_16463,N_16573);
nand U16703 (N_16703,N_16436,N_16429);
and U16704 (N_16704,N_16497,N_16507);
nand U16705 (N_16705,N_16508,N_16556);
and U16706 (N_16706,N_16401,N_16574);
nor U16707 (N_16707,N_16423,N_16542);
or U16708 (N_16708,N_16478,N_16468);
nand U16709 (N_16709,N_16425,N_16596);
xnor U16710 (N_16710,N_16585,N_16424);
or U16711 (N_16711,N_16498,N_16444);
and U16712 (N_16712,N_16499,N_16471);
nor U16713 (N_16713,N_16427,N_16440);
xor U16714 (N_16714,N_16462,N_16417);
nor U16715 (N_16715,N_16496,N_16581);
and U16716 (N_16716,N_16456,N_16503);
or U16717 (N_16717,N_16566,N_16474);
or U16718 (N_16718,N_16444,N_16587);
and U16719 (N_16719,N_16524,N_16457);
or U16720 (N_16720,N_16406,N_16459);
or U16721 (N_16721,N_16519,N_16578);
nand U16722 (N_16722,N_16460,N_16466);
or U16723 (N_16723,N_16404,N_16587);
nor U16724 (N_16724,N_16560,N_16455);
nand U16725 (N_16725,N_16556,N_16516);
nor U16726 (N_16726,N_16430,N_16502);
nand U16727 (N_16727,N_16418,N_16543);
nand U16728 (N_16728,N_16590,N_16407);
nor U16729 (N_16729,N_16488,N_16401);
and U16730 (N_16730,N_16509,N_16566);
nor U16731 (N_16731,N_16572,N_16533);
nor U16732 (N_16732,N_16541,N_16446);
nor U16733 (N_16733,N_16544,N_16516);
and U16734 (N_16734,N_16501,N_16492);
or U16735 (N_16735,N_16555,N_16444);
nand U16736 (N_16736,N_16433,N_16575);
nor U16737 (N_16737,N_16588,N_16489);
nand U16738 (N_16738,N_16426,N_16592);
and U16739 (N_16739,N_16557,N_16459);
xor U16740 (N_16740,N_16549,N_16408);
and U16741 (N_16741,N_16545,N_16444);
or U16742 (N_16742,N_16487,N_16508);
nand U16743 (N_16743,N_16543,N_16506);
or U16744 (N_16744,N_16540,N_16570);
and U16745 (N_16745,N_16506,N_16435);
and U16746 (N_16746,N_16569,N_16486);
or U16747 (N_16747,N_16583,N_16517);
nand U16748 (N_16748,N_16501,N_16433);
or U16749 (N_16749,N_16444,N_16442);
and U16750 (N_16750,N_16488,N_16484);
nor U16751 (N_16751,N_16402,N_16499);
nor U16752 (N_16752,N_16573,N_16578);
nor U16753 (N_16753,N_16529,N_16555);
nand U16754 (N_16754,N_16501,N_16469);
nand U16755 (N_16755,N_16543,N_16417);
and U16756 (N_16756,N_16456,N_16544);
nand U16757 (N_16757,N_16475,N_16565);
nor U16758 (N_16758,N_16531,N_16417);
nand U16759 (N_16759,N_16538,N_16579);
or U16760 (N_16760,N_16404,N_16453);
xnor U16761 (N_16761,N_16412,N_16419);
nor U16762 (N_16762,N_16526,N_16406);
nor U16763 (N_16763,N_16538,N_16582);
nand U16764 (N_16764,N_16572,N_16556);
nand U16765 (N_16765,N_16419,N_16484);
nand U16766 (N_16766,N_16513,N_16486);
nor U16767 (N_16767,N_16416,N_16461);
nand U16768 (N_16768,N_16421,N_16497);
nor U16769 (N_16769,N_16471,N_16405);
or U16770 (N_16770,N_16533,N_16505);
nand U16771 (N_16771,N_16599,N_16548);
nand U16772 (N_16772,N_16506,N_16493);
and U16773 (N_16773,N_16554,N_16491);
or U16774 (N_16774,N_16518,N_16579);
nor U16775 (N_16775,N_16412,N_16460);
and U16776 (N_16776,N_16584,N_16459);
or U16777 (N_16777,N_16529,N_16476);
nand U16778 (N_16778,N_16580,N_16507);
and U16779 (N_16779,N_16578,N_16581);
nand U16780 (N_16780,N_16474,N_16537);
nand U16781 (N_16781,N_16405,N_16412);
and U16782 (N_16782,N_16535,N_16547);
nor U16783 (N_16783,N_16592,N_16503);
nor U16784 (N_16784,N_16516,N_16459);
and U16785 (N_16785,N_16449,N_16452);
nor U16786 (N_16786,N_16407,N_16415);
and U16787 (N_16787,N_16413,N_16445);
nor U16788 (N_16788,N_16410,N_16521);
or U16789 (N_16789,N_16591,N_16497);
nand U16790 (N_16790,N_16550,N_16435);
nand U16791 (N_16791,N_16451,N_16432);
nand U16792 (N_16792,N_16482,N_16537);
nor U16793 (N_16793,N_16494,N_16450);
or U16794 (N_16794,N_16468,N_16483);
xnor U16795 (N_16795,N_16429,N_16442);
nor U16796 (N_16796,N_16567,N_16545);
nand U16797 (N_16797,N_16455,N_16506);
nand U16798 (N_16798,N_16413,N_16474);
nand U16799 (N_16799,N_16428,N_16497);
or U16800 (N_16800,N_16735,N_16608);
and U16801 (N_16801,N_16633,N_16706);
or U16802 (N_16802,N_16799,N_16687);
nor U16803 (N_16803,N_16770,N_16725);
and U16804 (N_16804,N_16632,N_16626);
or U16805 (N_16805,N_16617,N_16756);
xnor U16806 (N_16806,N_16700,N_16786);
nand U16807 (N_16807,N_16602,N_16755);
nor U16808 (N_16808,N_16657,N_16665);
nand U16809 (N_16809,N_16722,N_16792);
and U16810 (N_16810,N_16682,N_16796);
nand U16811 (N_16811,N_16738,N_16708);
and U16812 (N_16812,N_16754,N_16763);
and U16813 (N_16813,N_16788,N_16628);
xnor U16814 (N_16814,N_16787,N_16653);
nor U16815 (N_16815,N_16724,N_16669);
and U16816 (N_16816,N_16666,N_16723);
or U16817 (N_16817,N_16643,N_16703);
or U16818 (N_16818,N_16721,N_16651);
or U16819 (N_16819,N_16603,N_16690);
and U16820 (N_16820,N_16622,N_16672);
nor U16821 (N_16821,N_16764,N_16733);
nand U16822 (N_16822,N_16782,N_16776);
nand U16823 (N_16823,N_16771,N_16716);
nand U16824 (N_16824,N_16613,N_16798);
nand U16825 (N_16825,N_16652,N_16696);
nor U16826 (N_16826,N_16650,N_16619);
and U16827 (N_16827,N_16660,N_16697);
nand U16828 (N_16828,N_16752,N_16714);
or U16829 (N_16829,N_16728,N_16689);
xor U16830 (N_16830,N_16790,N_16719);
nor U16831 (N_16831,N_16670,N_16709);
and U16832 (N_16832,N_16795,N_16627);
nor U16833 (N_16833,N_16664,N_16705);
and U16834 (N_16834,N_16750,N_16695);
nor U16835 (N_16835,N_16692,N_16784);
and U16836 (N_16836,N_16760,N_16618);
nand U16837 (N_16837,N_16717,N_16640);
nor U16838 (N_16838,N_16704,N_16772);
or U16839 (N_16839,N_16773,N_16747);
or U16840 (N_16840,N_16641,N_16785);
or U16841 (N_16841,N_16688,N_16767);
nand U16842 (N_16842,N_16631,N_16729);
and U16843 (N_16843,N_16793,N_16607);
nand U16844 (N_16844,N_16600,N_16783);
nand U16845 (N_16845,N_16759,N_16727);
nand U16846 (N_16846,N_16761,N_16685);
nand U16847 (N_16847,N_16615,N_16610);
nor U16848 (N_16848,N_16702,N_16625);
and U16849 (N_16849,N_16791,N_16646);
and U16850 (N_16850,N_16720,N_16768);
or U16851 (N_16851,N_16779,N_16609);
nor U16852 (N_16852,N_16671,N_16736);
and U16853 (N_16853,N_16741,N_16656);
and U16854 (N_16854,N_16693,N_16744);
and U16855 (N_16855,N_16637,N_16616);
or U16856 (N_16856,N_16661,N_16635);
or U16857 (N_16857,N_16730,N_16758);
or U16858 (N_16858,N_16731,N_16691);
or U16859 (N_16859,N_16745,N_16746);
nand U16860 (N_16860,N_16781,N_16683);
or U16861 (N_16861,N_16734,N_16663);
xnor U16862 (N_16862,N_16680,N_16645);
nand U16863 (N_16863,N_16658,N_16612);
or U16864 (N_16864,N_16620,N_16679);
nand U16865 (N_16865,N_16748,N_16606);
nor U16866 (N_16866,N_16777,N_16667);
nor U16867 (N_16867,N_16739,N_16762);
and U16868 (N_16868,N_16737,N_16638);
and U16869 (N_16869,N_16636,N_16673);
nand U16870 (N_16870,N_16751,N_16774);
nor U16871 (N_16871,N_16644,N_16654);
nor U16872 (N_16872,N_16769,N_16699);
nand U16873 (N_16873,N_16611,N_16647);
nor U16874 (N_16874,N_16710,N_16732);
nor U16875 (N_16875,N_16698,N_16639);
or U16876 (N_16876,N_16630,N_16648);
or U16877 (N_16877,N_16707,N_16743);
xor U16878 (N_16878,N_16742,N_16749);
or U16879 (N_16879,N_16649,N_16621);
and U16880 (N_16880,N_16753,N_16624);
nand U16881 (N_16881,N_16684,N_16794);
nor U16882 (N_16882,N_16712,N_16726);
nand U16883 (N_16883,N_16677,N_16789);
and U16884 (N_16884,N_16674,N_16757);
nor U16885 (N_16885,N_16797,N_16662);
xor U16886 (N_16886,N_16694,N_16686);
and U16887 (N_16887,N_16778,N_16605);
nand U16888 (N_16888,N_16718,N_16676);
nor U16889 (N_16889,N_16659,N_16713);
and U16890 (N_16890,N_16715,N_16701);
nand U16891 (N_16891,N_16614,N_16629);
nor U16892 (N_16892,N_16740,N_16601);
and U16893 (N_16893,N_16623,N_16678);
and U16894 (N_16894,N_16711,N_16604);
nor U16895 (N_16895,N_16634,N_16681);
nor U16896 (N_16896,N_16765,N_16642);
or U16897 (N_16897,N_16668,N_16655);
or U16898 (N_16898,N_16775,N_16780);
or U16899 (N_16899,N_16766,N_16675);
and U16900 (N_16900,N_16728,N_16699);
or U16901 (N_16901,N_16627,N_16775);
or U16902 (N_16902,N_16662,N_16643);
or U16903 (N_16903,N_16779,N_16786);
or U16904 (N_16904,N_16738,N_16734);
and U16905 (N_16905,N_16729,N_16742);
and U16906 (N_16906,N_16670,N_16657);
nor U16907 (N_16907,N_16779,N_16623);
or U16908 (N_16908,N_16639,N_16742);
and U16909 (N_16909,N_16620,N_16669);
or U16910 (N_16910,N_16671,N_16653);
and U16911 (N_16911,N_16665,N_16728);
or U16912 (N_16912,N_16687,N_16712);
or U16913 (N_16913,N_16799,N_16653);
nand U16914 (N_16914,N_16633,N_16676);
or U16915 (N_16915,N_16664,N_16626);
and U16916 (N_16916,N_16738,N_16608);
nand U16917 (N_16917,N_16693,N_16792);
nor U16918 (N_16918,N_16773,N_16644);
or U16919 (N_16919,N_16796,N_16780);
nand U16920 (N_16920,N_16607,N_16717);
and U16921 (N_16921,N_16749,N_16750);
and U16922 (N_16922,N_16680,N_16785);
nand U16923 (N_16923,N_16643,N_16623);
or U16924 (N_16924,N_16733,N_16719);
or U16925 (N_16925,N_16675,N_16673);
nor U16926 (N_16926,N_16794,N_16752);
nor U16927 (N_16927,N_16703,N_16751);
or U16928 (N_16928,N_16751,N_16658);
and U16929 (N_16929,N_16619,N_16637);
or U16930 (N_16930,N_16630,N_16712);
or U16931 (N_16931,N_16630,N_16735);
or U16932 (N_16932,N_16710,N_16795);
nor U16933 (N_16933,N_16653,N_16699);
and U16934 (N_16934,N_16629,N_16769);
nand U16935 (N_16935,N_16601,N_16767);
nand U16936 (N_16936,N_16621,N_16743);
and U16937 (N_16937,N_16715,N_16784);
xnor U16938 (N_16938,N_16640,N_16708);
nand U16939 (N_16939,N_16604,N_16646);
or U16940 (N_16940,N_16623,N_16693);
or U16941 (N_16941,N_16732,N_16730);
or U16942 (N_16942,N_16740,N_16719);
nor U16943 (N_16943,N_16727,N_16728);
and U16944 (N_16944,N_16609,N_16690);
or U16945 (N_16945,N_16628,N_16787);
and U16946 (N_16946,N_16769,N_16691);
nor U16947 (N_16947,N_16626,N_16669);
and U16948 (N_16948,N_16727,N_16791);
or U16949 (N_16949,N_16656,N_16783);
nor U16950 (N_16950,N_16769,N_16730);
or U16951 (N_16951,N_16777,N_16736);
or U16952 (N_16952,N_16688,N_16756);
nor U16953 (N_16953,N_16765,N_16795);
and U16954 (N_16954,N_16766,N_16764);
nor U16955 (N_16955,N_16792,N_16637);
nand U16956 (N_16956,N_16711,N_16750);
and U16957 (N_16957,N_16665,N_16642);
nand U16958 (N_16958,N_16644,N_16612);
nor U16959 (N_16959,N_16780,N_16617);
nand U16960 (N_16960,N_16650,N_16797);
or U16961 (N_16961,N_16612,N_16695);
or U16962 (N_16962,N_16681,N_16703);
nor U16963 (N_16963,N_16646,N_16757);
or U16964 (N_16964,N_16726,N_16627);
nand U16965 (N_16965,N_16645,N_16618);
nand U16966 (N_16966,N_16637,N_16632);
nand U16967 (N_16967,N_16722,N_16695);
nand U16968 (N_16968,N_16664,N_16606);
or U16969 (N_16969,N_16785,N_16737);
and U16970 (N_16970,N_16778,N_16661);
nor U16971 (N_16971,N_16745,N_16634);
nor U16972 (N_16972,N_16775,N_16770);
nand U16973 (N_16973,N_16771,N_16654);
and U16974 (N_16974,N_16781,N_16736);
nand U16975 (N_16975,N_16678,N_16773);
nand U16976 (N_16976,N_16768,N_16756);
or U16977 (N_16977,N_16791,N_16753);
and U16978 (N_16978,N_16680,N_16776);
nand U16979 (N_16979,N_16700,N_16790);
nor U16980 (N_16980,N_16763,N_16781);
or U16981 (N_16981,N_16779,N_16790);
nor U16982 (N_16982,N_16671,N_16752);
or U16983 (N_16983,N_16738,N_16753);
nand U16984 (N_16984,N_16618,N_16750);
and U16985 (N_16985,N_16797,N_16796);
nand U16986 (N_16986,N_16763,N_16678);
nand U16987 (N_16987,N_16780,N_16677);
or U16988 (N_16988,N_16710,N_16723);
and U16989 (N_16989,N_16640,N_16677);
or U16990 (N_16990,N_16764,N_16650);
and U16991 (N_16991,N_16747,N_16710);
and U16992 (N_16992,N_16699,N_16600);
nor U16993 (N_16993,N_16696,N_16612);
or U16994 (N_16994,N_16694,N_16685);
nor U16995 (N_16995,N_16735,N_16724);
or U16996 (N_16996,N_16709,N_16741);
and U16997 (N_16997,N_16623,N_16786);
or U16998 (N_16998,N_16721,N_16686);
nor U16999 (N_16999,N_16623,N_16761);
xnor U17000 (N_17000,N_16868,N_16847);
nor U17001 (N_17001,N_16909,N_16993);
nand U17002 (N_17002,N_16984,N_16999);
nand U17003 (N_17003,N_16818,N_16962);
nand U17004 (N_17004,N_16820,N_16878);
or U17005 (N_17005,N_16947,N_16848);
nand U17006 (N_17006,N_16900,N_16828);
nor U17007 (N_17007,N_16985,N_16824);
or U17008 (N_17008,N_16854,N_16932);
or U17009 (N_17009,N_16905,N_16930);
and U17010 (N_17010,N_16906,N_16800);
or U17011 (N_17011,N_16831,N_16889);
nand U17012 (N_17012,N_16966,N_16978);
nand U17013 (N_17013,N_16840,N_16986);
nand U17014 (N_17014,N_16870,N_16945);
nor U17015 (N_17015,N_16917,N_16901);
xnor U17016 (N_17016,N_16876,N_16821);
nor U17017 (N_17017,N_16975,N_16851);
or U17018 (N_17018,N_16886,N_16974);
nor U17019 (N_17019,N_16817,N_16941);
nand U17020 (N_17020,N_16861,N_16931);
nor U17021 (N_17021,N_16850,N_16977);
or U17022 (N_17022,N_16896,N_16895);
nor U17023 (N_17023,N_16921,N_16804);
nand U17024 (N_17024,N_16825,N_16997);
and U17025 (N_17025,N_16926,N_16858);
nand U17026 (N_17026,N_16910,N_16830);
and U17027 (N_17027,N_16834,N_16855);
and U17028 (N_17028,N_16822,N_16898);
or U17029 (N_17029,N_16991,N_16934);
nand U17030 (N_17030,N_16839,N_16836);
nor U17031 (N_17031,N_16862,N_16807);
or U17032 (N_17032,N_16912,N_16942);
nand U17033 (N_17033,N_16965,N_16856);
and U17034 (N_17034,N_16819,N_16960);
or U17035 (N_17035,N_16990,N_16995);
or U17036 (N_17036,N_16994,N_16950);
and U17037 (N_17037,N_16955,N_16815);
and U17038 (N_17038,N_16863,N_16964);
nand U17039 (N_17039,N_16814,N_16860);
nor U17040 (N_17040,N_16838,N_16865);
nand U17041 (N_17041,N_16810,N_16989);
and U17042 (N_17042,N_16888,N_16951);
nor U17043 (N_17043,N_16826,N_16943);
nand U17044 (N_17044,N_16933,N_16922);
or U17045 (N_17045,N_16976,N_16899);
and U17046 (N_17046,N_16812,N_16927);
or U17047 (N_17047,N_16925,N_16969);
and U17048 (N_17048,N_16938,N_16988);
nor U17049 (N_17049,N_16940,N_16992);
nand U17050 (N_17050,N_16967,N_16894);
and U17051 (N_17051,N_16890,N_16983);
and U17052 (N_17052,N_16875,N_16843);
and U17053 (N_17053,N_16880,N_16903);
or U17054 (N_17054,N_16996,N_16884);
nand U17055 (N_17055,N_16844,N_16904);
or U17056 (N_17056,N_16841,N_16857);
nor U17057 (N_17057,N_16832,N_16902);
nand U17058 (N_17058,N_16956,N_16873);
or U17059 (N_17059,N_16893,N_16852);
nand U17060 (N_17060,N_16939,N_16864);
or U17061 (N_17061,N_16916,N_16929);
nand U17062 (N_17062,N_16846,N_16802);
nor U17063 (N_17063,N_16919,N_16979);
nor U17064 (N_17064,N_16891,N_16970);
nand U17065 (N_17065,N_16803,N_16954);
nand U17066 (N_17066,N_16801,N_16914);
nand U17067 (N_17067,N_16998,N_16920);
or U17068 (N_17068,N_16882,N_16944);
and U17069 (N_17069,N_16952,N_16879);
nor U17070 (N_17070,N_16827,N_16874);
nor U17071 (N_17071,N_16935,N_16971);
or U17072 (N_17072,N_16829,N_16936);
and U17073 (N_17073,N_16877,N_16937);
or U17074 (N_17074,N_16913,N_16968);
nand U17075 (N_17075,N_16959,N_16845);
nand U17076 (N_17076,N_16949,N_16958);
nand U17077 (N_17077,N_16881,N_16982);
and U17078 (N_17078,N_16887,N_16918);
and U17079 (N_17079,N_16835,N_16908);
and U17080 (N_17080,N_16961,N_16842);
xnor U17081 (N_17081,N_16811,N_16923);
nand U17082 (N_17082,N_16823,N_16859);
and U17083 (N_17083,N_16892,N_16928);
nor U17084 (N_17084,N_16853,N_16806);
xnor U17085 (N_17085,N_16869,N_16897);
nand U17086 (N_17086,N_16805,N_16867);
nor U17087 (N_17087,N_16813,N_16924);
or U17088 (N_17088,N_16883,N_16871);
and U17089 (N_17089,N_16816,N_16849);
and U17090 (N_17090,N_16837,N_16808);
nand U17091 (N_17091,N_16973,N_16866);
nand U17092 (N_17092,N_16809,N_16946);
or U17093 (N_17093,N_16833,N_16972);
and U17094 (N_17094,N_16915,N_16872);
nand U17095 (N_17095,N_16885,N_16963);
or U17096 (N_17096,N_16957,N_16987);
nor U17097 (N_17097,N_16980,N_16911);
nand U17098 (N_17098,N_16907,N_16953);
or U17099 (N_17099,N_16981,N_16948);
or U17100 (N_17100,N_16872,N_16932);
nor U17101 (N_17101,N_16951,N_16805);
and U17102 (N_17102,N_16870,N_16955);
and U17103 (N_17103,N_16860,N_16901);
and U17104 (N_17104,N_16876,N_16944);
nand U17105 (N_17105,N_16980,N_16904);
or U17106 (N_17106,N_16820,N_16877);
nor U17107 (N_17107,N_16996,N_16858);
nor U17108 (N_17108,N_16933,N_16809);
nand U17109 (N_17109,N_16906,N_16913);
nand U17110 (N_17110,N_16902,N_16882);
or U17111 (N_17111,N_16962,N_16953);
or U17112 (N_17112,N_16834,N_16830);
and U17113 (N_17113,N_16814,N_16986);
nand U17114 (N_17114,N_16859,N_16858);
or U17115 (N_17115,N_16913,N_16851);
nor U17116 (N_17116,N_16804,N_16960);
nor U17117 (N_17117,N_16851,N_16901);
xnor U17118 (N_17118,N_16921,N_16897);
or U17119 (N_17119,N_16950,N_16838);
nor U17120 (N_17120,N_16940,N_16954);
and U17121 (N_17121,N_16959,N_16917);
nand U17122 (N_17122,N_16963,N_16896);
and U17123 (N_17123,N_16826,N_16816);
nor U17124 (N_17124,N_16850,N_16820);
nor U17125 (N_17125,N_16829,N_16987);
and U17126 (N_17126,N_16807,N_16888);
and U17127 (N_17127,N_16906,N_16921);
or U17128 (N_17128,N_16913,N_16958);
nand U17129 (N_17129,N_16962,N_16910);
nor U17130 (N_17130,N_16939,N_16836);
nand U17131 (N_17131,N_16988,N_16877);
nand U17132 (N_17132,N_16929,N_16965);
xor U17133 (N_17133,N_16889,N_16901);
and U17134 (N_17134,N_16860,N_16822);
or U17135 (N_17135,N_16805,N_16910);
nor U17136 (N_17136,N_16986,N_16929);
nand U17137 (N_17137,N_16995,N_16905);
or U17138 (N_17138,N_16852,N_16970);
nand U17139 (N_17139,N_16924,N_16803);
nor U17140 (N_17140,N_16959,N_16982);
nand U17141 (N_17141,N_16969,N_16917);
or U17142 (N_17142,N_16884,N_16888);
or U17143 (N_17143,N_16952,N_16918);
or U17144 (N_17144,N_16976,N_16966);
nor U17145 (N_17145,N_16921,N_16901);
and U17146 (N_17146,N_16866,N_16936);
or U17147 (N_17147,N_16883,N_16984);
nand U17148 (N_17148,N_16964,N_16832);
nor U17149 (N_17149,N_16910,N_16964);
and U17150 (N_17150,N_16814,N_16900);
and U17151 (N_17151,N_16973,N_16975);
nand U17152 (N_17152,N_16822,N_16911);
nand U17153 (N_17153,N_16969,N_16920);
and U17154 (N_17154,N_16986,N_16805);
and U17155 (N_17155,N_16854,N_16968);
and U17156 (N_17156,N_16900,N_16816);
or U17157 (N_17157,N_16849,N_16839);
nand U17158 (N_17158,N_16864,N_16800);
nand U17159 (N_17159,N_16957,N_16893);
nand U17160 (N_17160,N_16984,N_16964);
nand U17161 (N_17161,N_16879,N_16963);
and U17162 (N_17162,N_16972,N_16965);
and U17163 (N_17163,N_16877,N_16987);
nor U17164 (N_17164,N_16960,N_16886);
and U17165 (N_17165,N_16938,N_16942);
and U17166 (N_17166,N_16835,N_16916);
nand U17167 (N_17167,N_16809,N_16853);
and U17168 (N_17168,N_16826,N_16820);
or U17169 (N_17169,N_16891,N_16834);
and U17170 (N_17170,N_16917,N_16932);
nor U17171 (N_17171,N_16896,N_16981);
or U17172 (N_17172,N_16827,N_16934);
nor U17173 (N_17173,N_16825,N_16946);
nand U17174 (N_17174,N_16974,N_16878);
or U17175 (N_17175,N_16921,N_16843);
nand U17176 (N_17176,N_16924,N_16807);
and U17177 (N_17177,N_16907,N_16983);
and U17178 (N_17178,N_16870,N_16896);
nand U17179 (N_17179,N_16989,N_16873);
nand U17180 (N_17180,N_16865,N_16976);
or U17181 (N_17181,N_16826,N_16866);
nor U17182 (N_17182,N_16916,N_16953);
nand U17183 (N_17183,N_16834,N_16904);
or U17184 (N_17184,N_16808,N_16940);
nand U17185 (N_17185,N_16912,N_16908);
nand U17186 (N_17186,N_16846,N_16970);
and U17187 (N_17187,N_16836,N_16915);
and U17188 (N_17188,N_16940,N_16924);
or U17189 (N_17189,N_16839,N_16844);
or U17190 (N_17190,N_16834,N_16956);
or U17191 (N_17191,N_16907,N_16943);
or U17192 (N_17192,N_16914,N_16988);
or U17193 (N_17193,N_16982,N_16927);
or U17194 (N_17194,N_16986,N_16872);
nand U17195 (N_17195,N_16875,N_16908);
nand U17196 (N_17196,N_16841,N_16929);
and U17197 (N_17197,N_16904,N_16820);
nand U17198 (N_17198,N_16966,N_16881);
or U17199 (N_17199,N_16892,N_16800);
nor U17200 (N_17200,N_17139,N_17199);
and U17201 (N_17201,N_17115,N_17014);
nor U17202 (N_17202,N_17168,N_17042);
and U17203 (N_17203,N_17100,N_17015);
or U17204 (N_17204,N_17138,N_17072);
and U17205 (N_17205,N_17029,N_17060);
and U17206 (N_17206,N_17119,N_17126);
nor U17207 (N_17207,N_17067,N_17163);
or U17208 (N_17208,N_17046,N_17169);
nand U17209 (N_17209,N_17142,N_17098);
or U17210 (N_17210,N_17088,N_17122);
nand U17211 (N_17211,N_17141,N_17040);
nand U17212 (N_17212,N_17077,N_17125);
or U17213 (N_17213,N_17034,N_17021);
and U17214 (N_17214,N_17105,N_17028);
and U17215 (N_17215,N_17073,N_17045);
nand U17216 (N_17216,N_17024,N_17195);
and U17217 (N_17217,N_17056,N_17026);
nand U17218 (N_17218,N_17117,N_17071);
nand U17219 (N_17219,N_17008,N_17143);
and U17220 (N_17220,N_17104,N_17121);
or U17221 (N_17221,N_17118,N_17180);
nor U17222 (N_17222,N_17110,N_17131);
and U17223 (N_17223,N_17062,N_17010);
nor U17224 (N_17224,N_17137,N_17091);
or U17225 (N_17225,N_17149,N_17099);
or U17226 (N_17226,N_17147,N_17055);
or U17227 (N_17227,N_17124,N_17038);
nand U17228 (N_17228,N_17170,N_17171);
and U17229 (N_17229,N_17150,N_17123);
or U17230 (N_17230,N_17096,N_17069);
nor U17231 (N_17231,N_17101,N_17114);
and U17232 (N_17232,N_17127,N_17039);
nand U17233 (N_17233,N_17043,N_17068);
or U17234 (N_17234,N_17074,N_17094);
nor U17235 (N_17235,N_17061,N_17189);
or U17236 (N_17236,N_17035,N_17063);
or U17237 (N_17237,N_17174,N_17113);
nand U17238 (N_17238,N_17109,N_17082);
nand U17239 (N_17239,N_17019,N_17191);
nand U17240 (N_17240,N_17044,N_17197);
nor U17241 (N_17241,N_17106,N_17182);
or U17242 (N_17242,N_17116,N_17185);
or U17243 (N_17243,N_17097,N_17187);
or U17244 (N_17244,N_17000,N_17081);
and U17245 (N_17245,N_17192,N_17186);
nand U17246 (N_17246,N_17162,N_17166);
or U17247 (N_17247,N_17005,N_17002);
nor U17248 (N_17248,N_17037,N_17193);
nor U17249 (N_17249,N_17135,N_17066);
nor U17250 (N_17250,N_17012,N_17001);
or U17251 (N_17251,N_17181,N_17048);
or U17252 (N_17252,N_17058,N_17052);
or U17253 (N_17253,N_17030,N_17032);
nand U17254 (N_17254,N_17017,N_17031);
and U17255 (N_17255,N_17049,N_17151);
nor U17256 (N_17256,N_17018,N_17053);
and U17257 (N_17257,N_17190,N_17188);
nor U17258 (N_17258,N_17136,N_17004);
nand U17259 (N_17259,N_17112,N_17089);
or U17260 (N_17260,N_17183,N_17103);
nor U17261 (N_17261,N_17178,N_17108);
or U17262 (N_17262,N_17157,N_17054);
or U17263 (N_17263,N_17173,N_17175);
nand U17264 (N_17264,N_17003,N_17172);
nand U17265 (N_17265,N_17007,N_17176);
or U17266 (N_17266,N_17194,N_17095);
nand U17267 (N_17267,N_17047,N_17020);
xnor U17268 (N_17268,N_17084,N_17158);
nor U17269 (N_17269,N_17041,N_17177);
and U17270 (N_17270,N_17144,N_17198);
nand U17271 (N_17271,N_17064,N_17080);
nand U17272 (N_17272,N_17057,N_17152);
nor U17273 (N_17273,N_17165,N_17065);
and U17274 (N_17274,N_17033,N_17079);
or U17275 (N_17275,N_17128,N_17120);
nor U17276 (N_17276,N_17184,N_17006);
or U17277 (N_17277,N_17140,N_17161);
nand U17278 (N_17278,N_17167,N_17051);
nand U17279 (N_17279,N_17085,N_17179);
xor U17280 (N_17280,N_17092,N_17090);
or U17281 (N_17281,N_17155,N_17146);
nand U17282 (N_17282,N_17076,N_17025);
nand U17283 (N_17283,N_17023,N_17107);
or U17284 (N_17284,N_17111,N_17133);
nor U17285 (N_17285,N_17153,N_17164);
and U17286 (N_17286,N_17145,N_17075);
or U17287 (N_17287,N_17134,N_17154);
nor U17288 (N_17288,N_17059,N_17156);
or U17289 (N_17289,N_17016,N_17009);
xnor U17290 (N_17290,N_17078,N_17070);
nor U17291 (N_17291,N_17087,N_17050);
nor U17292 (N_17292,N_17022,N_17102);
nand U17293 (N_17293,N_17013,N_17130);
nand U17294 (N_17294,N_17129,N_17159);
nor U17295 (N_17295,N_17027,N_17011);
or U17296 (N_17296,N_17160,N_17196);
nand U17297 (N_17297,N_17132,N_17148);
nor U17298 (N_17298,N_17086,N_17036);
or U17299 (N_17299,N_17083,N_17093);
nand U17300 (N_17300,N_17191,N_17141);
nor U17301 (N_17301,N_17145,N_17097);
nor U17302 (N_17302,N_17052,N_17167);
nand U17303 (N_17303,N_17168,N_17180);
and U17304 (N_17304,N_17084,N_17092);
or U17305 (N_17305,N_17049,N_17109);
and U17306 (N_17306,N_17047,N_17018);
nor U17307 (N_17307,N_17107,N_17145);
or U17308 (N_17308,N_17199,N_17095);
or U17309 (N_17309,N_17166,N_17058);
or U17310 (N_17310,N_17023,N_17020);
nand U17311 (N_17311,N_17073,N_17126);
and U17312 (N_17312,N_17033,N_17108);
nor U17313 (N_17313,N_17074,N_17066);
nand U17314 (N_17314,N_17183,N_17140);
or U17315 (N_17315,N_17156,N_17104);
and U17316 (N_17316,N_17021,N_17111);
and U17317 (N_17317,N_17164,N_17151);
nand U17318 (N_17318,N_17160,N_17062);
and U17319 (N_17319,N_17162,N_17149);
nor U17320 (N_17320,N_17029,N_17161);
nand U17321 (N_17321,N_17010,N_17154);
or U17322 (N_17322,N_17072,N_17012);
and U17323 (N_17323,N_17055,N_17029);
and U17324 (N_17324,N_17001,N_17047);
nor U17325 (N_17325,N_17175,N_17065);
and U17326 (N_17326,N_17099,N_17194);
nor U17327 (N_17327,N_17028,N_17085);
or U17328 (N_17328,N_17123,N_17186);
nor U17329 (N_17329,N_17149,N_17169);
nand U17330 (N_17330,N_17010,N_17038);
nor U17331 (N_17331,N_17078,N_17135);
and U17332 (N_17332,N_17153,N_17075);
nor U17333 (N_17333,N_17028,N_17129);
nor U17334 (N_17334,N_17083,N_17098);
and U17335 (N_17335,N_17162,N_17182);
and U17336 (N_17336,N_17112,N_17091);
nor U17337 (N_17337,N_17012,N_17137);
nor U17338 (N_17338,N_17067,N_17133);
nor U17339 (N_17339,N_17163,N_17078);
nand U17340 (N_17340,N_17079,N_17165);
or U17341 (N_17341,N_17020,N_17106);
and U17342 (N_17342,N_17063,N_17040);
nand U17343 (N_17343,N_17144,N_17119);
and U17344 (N_17344,N_17177,N_17058);
nor U17345 (N_17345,N_17134,N_17045);
nor U17346 (N_17346,N_17124,N_17197);
nand U17347 (N_17347,N_17075,N_17183);
or U17348 (N_17348,N_17009,N_17161);
and U17349 (N_17349,N_17083,N_17024);
nor U17350 (N_17350,N_17011,N_17120);
nor U17351 (N_17351,N_17034,N_17124);
nand U17352 (N_17352,N_17017,N_17088);
nor U17353 (N_17353,N_17177,N_17141);
and U17354 (N_17354,N_17194,N_17033);
or U17355 (N_17355,N_17011,N_17069);
nor U17356 (N_17356,N_17145,N_17165);
and U17357 (N_17357,N_17035,N_17102);
nand U17358 (N_17358,N_17090,N_17135);
and U17359 (N_17359,N_17009,N_17044);
or U17360 (N_17360,N_17191,N_17002);
nor U17361 (N_17361,N_17014,N_17075);
and U17362 (N_17362,N_17032,N_17111);
or U17363 (N_17363,N_17042,N_17066);
nor U17364 (N_17364,N_17029,N_17018);
or U17365 (N_17365,N_17039,N_17038);
nand U17366 (N_17366,N_17025,N_17164);
nor U17367 (N_17367,N_17003,N_17054);
or U17368 (N_17368,N_17000,N_17107);
nand U17369 (N_17369,N_17078,N_17097);
nor U17370 (N_17370,N_17192,N_17141);
and U17371 (N_17371,N_17176,N_17025);
nor U17372 (N_17372,N_17140,N_17057);
and U17373 (N_17373,N_17004,N_17082);
or U17374 (N_17374,N_17003,N_17151);
nor U17375 (N_17375,N_17171,N_17094);
xnor U17376 (N_17376,N_17011,N_17132);
and U17377 (N_17377,N_17091,N_17169);
nor U17378 (N_17378,N_17129,N_17096);
nor U17379 (N_17379,N_17146,N_17066);
and U17380 (N_17380,N_17031,N_17195);
nor U17381 (N_17381,N_17092,N_17170);
or U17382 (N_17382,N_17164,N_17146);
or U17383 (N_17383,N_17162,N_17151);
or U17384 (N_17384,N_17092,N_17163);
nor U17385 (N_17385,N_17079,N_17008);
nor U17386 (N_17386,N_17191,N_17006);
nor U17387 (N_17387,N_17199,N_17127);
nor U17388 (N_17388,N_17190,N_17070);
nor U17389 (N_17389,N_17078,N_17107);
or U17390 (N_17390,N_17096,N_17050);
nand U17391 (N_17391,N_17199,N_17075);
and U17392 (N_17392,N_17130,N_17184);
and U17393 (N_17393,N_17178,N_17177);
nand U17394 (N_17394,N_17040,N_17012);
or U17395 (N_17395,N_17163,N_17002);
nand U17396 (N_17396,N_17040,N_17127);
or U17397 (N_17397,N_17135,N_17070);
nor U17398 (N_17398,N_17106,N_17129);
or U17399 (N_17399,N_17144,N_17196);
nand U17400 (N_17400,N_17285,N_17370);
nor U17401 (N_17401,N_17304,N_17308);
nand U17402 (N_17402,N_17367,N_17207);
xnor U17403 (N_17403,N_17244,N_17263);
nand U17404 (N_17404,N_17346,N_17216);
nor U17405 (N_17405,N_17347,N_17268);
nand U17406 (N_17406,N_17355,N_17351);
nand U17407 (N_17407,N_17239,N_17302);
or U17408 (N_17408,N_17327,N_17376);
nor U17409 (N_17409,N_17241,N_17318);
nand U17410 (N_17410,N_17253,N_17298);
or U17411 (N_17411,N_17294,N_17372);
nor U17412 (N_17412,N_17356,N_17309);
nand U17413 (N_17413,N_17303,N_17206);
nand U17414 (N_17414,N_17387,N_17229);
or U17415 (N_17415,N_17366,N_17301);
nor U17416 (N_17416,N_17250,N_17369);
or U17417 (N_17417,N_17320,N_17329);
and U17418 (N_17418,N_17277,N_17278);
nand U17419 (N_17419,N_17251,N_17214);
nand U17420 (N_17420,N_17340,N_17295);
nor U17421 (N_17421,N_17338,N_17392);
nor U17422 (N_17422,N_17322,N_17345);
and U17423 (N_17423,N_17380,N_17328);
and U17424 (N_17424,N_17281,N_17326);
and U17425 (N_17425,N_17260,N_17249);
nor U17426 (N_17426,N_17323,N_17381);
nand U17427 (N_17427,N_17266,N_17385);
or U17428 (N_17428,N_17225,N_17292);
and U17429 (N_17429,N_17352,N_17297);
or U17430 (N_17430,N_17362,N_17264);
nor U17431 (N_17431,N_17371,N_17288);
or U17432 (N_17432,N_17291,N_17311);
or U17433 (N_17433,N_17348,N_17286);
nor U17434 (N_17434,N_17389,N_17396);
and U17435 (N_17435,N_17221,N_17330);
nand U17436 (N_17436,N_17365,N_17236);
nor U17437 (N_17437,N_17240,N_17305);
nand U17438 (N_17438,N_17200,N_17350);
and U17439 (N_17439,N_17339,N_17373);
or U17440 (N_17440,N_17276,N_17315);
nand U17441 (N_17441,N_17242,N_17296);
or U17442 (N_17442,N_17306,N_17254);
nor U17443 (N_17443,N_17210,N_17270);
or U17444 (N_17444,N_17272,N_17220);
and U17445 (N_17445,N_17235,N_17314);
and U17446 (N_17446,N_17324,N_17223);
nand U17447 (N_17447,N_17289,N_17222);
and U17448 (N_17448,N_17265,N_17247);
nand U17449 (N_17449,N_17357,N_17273);
nor U17450 (N_17450,N_17243,N_17349);
nand U17451 (N_17451,N_17290,N_17237);
nand U17452 (N_17452,N_17246,N_17397);
and U17453 (N_17453,N_17258,N_17252);
and U17454 (N_17454,N_17230,N_17337);
or U17455 (N_17455,N_17218,N_17382);
or U17456 (N_17456,N_17307,N_17211);
and U17457 (N_17457,N_17300,N_17361);
and U17458 (N_17458,N_17398,N_17394);
nand U17459 (N_17459,N_17359,N_17209);
nand U17460 (N_17460,N_17299,N_17375);
nor U17461 (N_17461,N_17201,N_17317);
or U17462 (N_17462,N_17377,N_17293);
nor U17463 (N_17463,N_17231,N_17257);
nor U17464 (N_17464,N_17334,N_17259);
nor U17465 (N_17465,N_17202,N_17378);
nand U17466 (N_17466,N_17232,N_17219);
nor U17467 (N_17467,N_17208,N_17227);
nand U17468 (N_17468,N_17245,N_17332);
nor U17469 (N_17469,N_17333,N_17312);
nand U17470 (N_17470,N_17379,N_17212);
nor U17471 (N_17471,N_17364,N_17336);
nor U17472 (N_17472,N_17284,N_17269);
nor U17473 (N_17473,N_17287,N_17331);
and U17474 (N_17474,N_17280,N_17233);
nand U17475 (N_17475,N_17255,N_17213);
or U17476 (N_17476,N_17313,N_17321);
or U17477 (N_17477,N_17399,N_17234);
nor U17478 (N_17478,N_17261,N_17360);
nand U17479 (N_17479,N_17391,N_17368);
xor U17480 (N_17480,N_17395,N_17325);
and U17481 (N_17481,N_17262,N_17274);
nor U17482 (N_17482,N_17386,N_17343);
nor U17483 (N_17483,N_17238,N_17342);
nor U17484 (N_17484,N_17335,N_17374);
nand U17485 (N_17485,N_17310,N_17256);
and U17486 (N_17486,N_17226,N_17363);
nor U17487 (N_17487,N_17388,N_17393);
nor U17488 (N_17488,N_17316,N_17204);
nand U17489 (N_17489,N_17271,N_17228);
nor U17490 (N_17490,N_17354,N_17353);
nand U17491 (N_17491,N_17341,N_17275);
xnor U17492 (N_17492,N_17224,N_17267);
and U17493 (N_17493,N_17203,N_17217);
or U17494 (N_17494,N_17282,N_17383);
and U17495 (N_17495,N_17358,N_17390);
nand U17496 (N_17496,N_17319,N_17384);
or U17497 (N_17497,N_17248,N_17344);
nor U17498 (N_17498,N_17279,N_17215);
xor U17499 (N_17499,N_17283,N_17205);
or U17500 (N_17500,N_17210,N_17393);
or U17501 (N_17501,N_17261,N_17241);
nor U17502 (N_17502,N_17206,N_17234);
or U17503 (N_17503,N_17244,N_17357);
nand U17504 (N_17504,N_17347,N_17358);
nand U17505 (N_17505,N_17211,N_17295);
or U17506 (N_17506,N_17322,N_17384);
and U17507 (N_17507,N_17374,N_17307);
nor U17508 (N_17508,N_17249,N_17366);
nand U17509 (N_17509,N_17247,N_17353);
nand U17510 (N_17510,N_17364,N_17262);
or U17511 (N_17511,N_17297,N_17316);
nor U17512 (N_17512,N_17231,N_17294);
and U17513 (N_17513,N_17213,N_17318);
nor U17514 (N_17514,N_17316,N_17345);
xnor U17515 (N_17515,N_17213,N_17243);
nand U17516 (N_17516,N_17267,N_17252);
and U17517 (N_17517,N_17280,N_17262);
nand U17518 (N_17518,N_17394,N_17264);
nand U17519 (N_17519,N_17345,N_17398);
nor U17520 (N_17520,N_17322,N_17306);
nand U17521 (N_17521,N_17281,N_17396);
nor U17522 (N_17522,N_17375,N_17271);
and U17523 (N_17523,N_17324,N_17387);
nor U17524 (N_17524,N_17288,N_17227);
nand U17525 (N_17525,N_17345,N_17320);
nor U17526 (N_17526,N_17216,N_17369);
or U17527 (N_17527,N_17398,N_17309);
nor U17528 (N_17528,N_17361,N_17202);
or U17529 (N_17529,N_17375,N_17254);
nand U17530 (N_17530,N_17308,N_17357);
nand U17531 (N_17531,N_17370,N_17247);
or U17532 (N_17532,N_17226,N_17360);
or U17533 (N_17533,N_17227,N_17297);
nor U17534 (N_17534,N_17381,N_17243);
nand U17535 (N_17535,N_17300,N_17293);
nand U17536 (N_17536,N_17341,N_17355);
and U17537 (N_17537,N_17379,N_17269);
nand U17538 (N_17538,N_17286,N_17241);
or U17539 (N_17539,N_17206,N_17207);
nand U17540 (N_17540,N_17298,N_17353);
and U17541 (N_17541,N_17219,N_17348);
nand U17542 (N_17542,N_17256,N_17340);
or U17543 (N_17543,N_17363,N_17277);
or U17544 (N_17544,N_17233,N_17352);
nor U17545 (N_17545,N_17388,N_17267);
and U17546 (N_17546,N_17229,N_17347);
nor U17547 (N_17547,N_17330,N_17235);
nand U17548 (N_17548,N_17374,N_17372);
nor U17549 (N_17549,N_17245,N_17200);
or U17550 (N_17550,N_17344,N_17293);
and U17551 (N_17551,N_17365,N_17206);
nor U17552 (N_17552,N_17348,N_17333);
xor U17553 (N_17553,N_17393,N_17341);
or U17554 (N_17554,N_17215,N_17272);
and U17555 (N_17555,N_17383,N_17396);
nor U17556 (N_17556,N_17311,N_17334);
and U17557 (N_17557,N_17395,N_17383);
and U17558 (N_17558,N_17278,N_17345);
or U17559 (N_17559,N_17277,N_17356);
or U17560 (N_17560,N_17237,N_17343);
and U17561 (N_17561,N_17213,N_17336);
or U17562 (N_17562,N_17354,N_17314);
and U17563 (N_17563,N_17212,N_17221);
xor U17564 (N_17564,N_17396,N_17330);
nand U17565 (N_17565,N_17220,N_17254);
nor U17566 (N_17566,N_17263,N_17251);
nor U17567 (N_17567,N_17389,N_17286);
xnor U17568 (N_17568,N_17222,N_17263);
nand U17569 (N_17569,N_17205,N_17308);
or U17570 (N_17570,N_17231,N_17352);
or U17571 (N_17571,N_17354,N_17317);
or U17572 (N_17572,N_17291,N_17277);
nor U17573 (N_17573,N_17304,N_17246);
nand U17574 (N_17574,N_17378,N_17264);
xor U17575 (N_17575,N_17204,N_17266);
and U17576 (N_17576,N_17352,N_17382);
or U17577 (N_17577,N_17382,N_17294);
nor U17578 (N_17578,N_17255,N_17295);
or U17579 (N_17579,N_17384,N_17200);
nor U17580 (N_17580,N_17298,N_17336);
or U17581 (N_17581,N_17318,N_17255);
or U17582 (N_17582,N_17242,N_17226);
and U17583 (N_17583,N_17287,N_17342);
and U17584 (N_17584,N_17209,N_17250);
nand U17585 (N_17585,N_17362,N_17202);
nand U17586 (N_17586,N_17258,N_17220);
nor U17587 (N_17587,N_17268,N_17211);
and U17588 (N_17588,N_17254,N_17335);
nand U17589 (N_17589,N_17201,N_17232);
xnor U17590 (N_17590,N_17349,N_17308);
or U17591 (N_17591,N_17282,N_17293);
nor U17592 (N_17592,N_17394,N_17321);
nor U17593 (N_17593,N_17287,N_17279);
nand U17594 (N_17594,N_17278,N_17266);
nor U17595 (N_17595,N_17204,N_17232);
nor U17596 (N_17596,N_17231,N_17219);
nand U17597 (N_17597,N_17266,N_17233);
and U17598 (N_17598,N_17266,N_17286);
nor U17599 (N_17599,N_17314,N_17392);
nand U17600 (N_17600,N_17403,N_17441);
nor U17601 (N_17601,N_17465,N_17519);
nor U17602 (N_17602,N_17596,N_17520);
nand U17603 (N_17603,N_17434,N_17572);
and U17604 (N_17604,N_17530,N_17451);
nand U17605 (N_17605,N_17540,N_17553);
or U17606 (N_17606,N_17427,N_17505);
or U17607 (N_17607,N_17438,N_17576);
or U17608 (N_17608,N_17457,N_17518);
and U17609 (N_17609,N_17580,N_17581);
and U17610 (N_17610,N_17545,N_17516);
or U17611 (N_17611,N_17532,N_17582);
nor U17612 (N_17612,N_17436,N_17578);
xnor U17613 (N_17613,N_17497,N_17543);
nor U17614 (N_17614,N_17423,N_17536);
or U17615 (N_17615,N_17432,N_17597);
nand U17616 (N_17616,N_17498,N_17531);
or U17617 (N_17617,N_17546,N_17430);
or U17618 (N_17618,N_17431,N_17420);
nand U17619 (N_17619,N_17405,N_17475);
nand U17620 (N_17620,N_17538,N_17474);
nor U17621 (N_17621,N_17489,N_17586);
or U17622 (N_17622,N_17426,N_17537);
and U17623 (N_17623,N_17407,N_17483);
nor U17624 (N_17624,N_17473,N_17484);
and U17625 (N_17625,N_17452,N_17523);
nand U17626 (N_17626,N_17535,N_17588);
nand U17627 (N_17627,N_17554,N_17468);
nor U17628 (N_17628,N_17459,N_17443);
nor U17629 (N_17629,N_17563,N_17401);
nand U17630 (N_17630,N_17534,N_17555);
or U17631 (N_17631,N_17560,N_17525);
or U17632 (N_17632,N_17562,N_17558);
and U17633 (N_17633,N_17450,N_17585);
nand U17634 (N_17634,N_17491,N_17404);
nor U17635 (N_17635,N_17466,N_17564);
nor U17636 (N_17636,N_17449,N_17512);
nand U17637 (N_17637,N_17589,N_17527);
nand U17638 (N_17638,N_17460,N_17458);
or U17639 (N_17639,N_17476,N_17501);
and U17640 (N_17640,N_17469,N_17444);
and U17641 (N_17641,N_17570,N_17446);
nor U17642 (N_17642,N_17524,N_17425);
or U17643 (N_17643,N_17481,N_17488);
nor U17644 (N_17644,N_17511,N_17528);
nand U17645 (N_17645,N_17565,N_17499);
or U17646 (N_17646,N_17593,N_17418);
xnor U17647 (N_17647,N_17406,N_17400);
or U17648 (N_17648,N_17504,N_17573);
nor U17649 (N_17649,N_17591,N_17409);
or U17650 (N_17650,N_17548,N_17453);
nor U17651 (N_17651,N_17502,N_17567);
nand U17652 (N_17652,N_17470,N_17419);
nand U17653 (N_17653,N_17503,N_17556);
or U17654 (N_17654,N_17542,N_17428);
or U17655 (N_17655,N_17541,N_17472);
nand U17656 (N_17656,N_17482,N_17408);
nand U17657 (N_17657,N_17583,N_17549);
nor U17658 (N_17658,N_17594,N_17508);
or U17659 (N_17659,N_17415,N_17526);
nand U17660 (N_17660,N_17485,N_17456);
nor U17661 (N_17661,N_17447,N_17575);
and U17662 (N_17662,N_17552,N_17467);
or U17663 (N_17663,N_17595,N_17584);
nor U17664 (N_17664,N_17429,N_17442);
or U17665 (N_17665,N_17529,N_17463);
or U17666 (N_17666,N_17507,N_17510);
nand U17667 (N_17667,N_17454,N_17577);
nand U17668 (N_17668,N_17551,N_17592);
nand U17669 (N_17669,N_17550,N_17533);
or U17670 (N_17670,N_17496,N_17471);
nor U17671 (N_17671,N_17437,N_17410);
nor U17672 (N_17672,N_17506,N_17490);
nand U17673 (N_17673,N_17413,N_17433);
and U17674 (N_17674,N_17515,N_17574);
or U17675 (N_17675,N_17464,N_17412);
and U17676 (N_17676,N_17539,N_17487);
nand U17677 (N_17677,N_17522,N_17402);
nor U17678 (N_17678,N_17455,N_17416);
and U17679 (N_17679,N_17559,N_17599);
or U17680 (N_17680,N_17486,N_17561);
or U17681 (N_17681,N_17435,N_17571);
nor U17682 (N_17682,N_17514,N_17422);
xor U17683 (N_17683,N_17557,N_17569);
nand U17684 (N_17684,N_17598,N_17568);
nor U17685 (N_17685,N_17513,N_17500);
and U17686 (N_17686,N_17448,N_17544);
and U17687 (N_17687,N_17439,N_17477);
or U17688 (N_17688,N_17461,N_17440);
or U17689 (N_17689,N_17587,N_17462);
xnor U17690 (N_17690,N_17417,N_17579);
nor U17691 (N_17691,N_17421,N_17492);
and U17692 (N_17692,N_17424,N_17495);
nor U17693 (N_17693,N_17445,N_17479);
and U17694 (N_17694,N_17414,N_17493);
nand U17695 (N_17695,N_17590,N_17547);
nor U17696 (N_17696,N_17494,N_17517);
and U17697 (N_17697,N_17509,N_17480);
and U17698 (N_17698,N_17566,N_17521);
and U17699 (N_17699,N_17478,N_17411);
nand U17700 (N_17700,N_17402,N_17418);
nor U17701 (N_17701,N_17431,N_17471);
nor U17702 (N_17702,N_17419,N_17557);
or U17703 (N_17703,N_17504,N_17517);
and U17704 (N_17704,N_17569,N_17445);
or U17705 (N_17705,N_17432,N_17471);
and U17706 (N_17706,N_17410,N_17461);
or U17707 (N_17707,N_17492,N_17453);
or U17708 (N_17708,N_17527,N_17448);
nor U17709 (N_17709,N_17406,N_17516);
nand U17710 (N_17710,N_17559,N_17463);
nand U17711 (N_17711,N_17522,N_17515);
and U17712 (N_17712,N_17494,N_17589);
or U17713 (N_17713,N_17502,N_17444);
nor U17714 (N_17714,N_17524,N_17584);
nor U17715 (N_17715,N_17537,N_17476);
or U17716 (N_17716,N_17471,N_17508);
and U17717 (N_17717,N_17513,N_17482);
or U17718 (N_17718,N_17585,N_17554);
nand U17719 (N_17719,N_17508,N_17433);
or U17720 (N_17720,N_17596,N_17555);
xnor U17721 (N_17721,N_17515,N_17590);
or U17722 (N_17722,N_17487,N_17458);
nand U17723 (N_17723,N_17521,N_17409);
nor U17724 (N_17724,N_17592,N_17597);
nor U17725 (N_17725,N_17440,N_17521);
nand U17726 (N_17726,N_17593,N_17531);
nor U17727 (N_17727,N_17543,N_17454);
or U17728 (N_17728,N_17568,N_17559);
nand U17729 (N_17729,N_17467,N_17412);
nand U17730 (N_17730,N_17449,N_17455);
and U17731 (N_17731,N_17528,N_17556);
or U17732 (N_17732,N_17406,N_17422);
nor U17733 (N_17733,N_17469,N_17512);
or U17734 (N_17734,N_17421,N_17597);
or U17735 (N_17735,N_17415,N_17563);
and U17736 (N_17736,N_17456,N_17486);
or U17737 (N_17737,N_17501,N_17401);
nand U17738 (N_17738,N_17539,N_17518);
or U17739 (N_17739,N_17423,N_17556);
nor U17740 (N_17740,N_17584,N_17476);
nor U17741 (N_17741,N_17500,N_17494);
or U17742 (N_17742,N_17549,N_17473);
xnor U17743 (N_17743,N_17594,N_17440);
and U17744 (N_17744,N_17490,N_17456);
or U17745 (N_17745,N_17508,N_17540);
nand U17746 (N_17746,N_17507,N_17477);
and U17747 (N_17747,N_17494,N_17449);
or U17748 (N_17748,N_17464,N_17527);
and U17749 (N_17749,N_17545,N_17587);
nor U17750 (N_17750,N_17580,N_17573);
and U17751 (N_17751,N_17516,N_17425);
nand U17752 (N_17752,N_17474,N_17408);
nor U17753 (N_17753,N_17454,N_17496);
nor U17754 (N_17754,N_17569,N_17410);
nor U17755 (N_17755,N_17468,N_17552);
nor U17756 (N_17756,N_17429,N_17543);
nand U17757 (N_17757,N_17572,N_17508);
and U17758 (N_17758,N_17406,N_17456);
nor U17759 (N_17759,N_17453,N_17580);
and U17760 (N_17760,N_17452,N_17592);
or U17761 (N_17761,N_17449,N_17594);
nor U17762 (N_17762,N_17452,N_17462);
nor U17763 (N_17763,N_17493,N_17580);
and U17764 (N_17764,N_17403,N_17478);
and U17765 (N_17765,N_17488,N_17431);
or U17766 (N_17766,N_17589,N_17587);
or U17767 (N_17767,N_17593,N_17482);
nand U17768 (N_17768,N_17594,N_17488);
nand U17769 (N_17769,N_17424,N_17481);
nand U17770 (N_17770,N_17422,N_17591);
nor U17771 (N_17771,N_17591,N_17434);
nor U17772 (N_17772,N_17553,N_17552);
nor U17773 (N_17773,N_17424,N_17595);
nand U17774 (N_17774,N_17486,N_17427);
nor U17775 (N_17775,N_17404,N_17569);
nand U17776 (N_17776,N_17425,N_17474);
nor U17777 (N_17777,N_17484,N_17553);
nor U17778 (N_17778,N_17419,N_17434);
or U17779 (N_17779,N_17562,N_17524);
nor U17780 (N_17780,N_17529,N_17556);
and U17781 (N_17781,N_17586,N_17536);
nor U17782 (N_17782,N_17446,N_17499);
nand U17783 (N_17783,N_17564,N_17470);
nand U17784 (N_17784,N_17573,N_17417);
and U17785 (N_17785,N_17541,N_17599);
nor U17786 (N_17786,N_17476,N_17466);
nand U17787 (N_17787,N_17590,N_17534);
or U17788 (N_17788,N_17454,N_17491);
nor U17789 (N_17789,N_17436,N_17421);
nand U17790 (N_17790,N_17596,N_17517);
nor U17791 (N_17791,N_17577,N_17410);
nor U17792 (N_17792,N_17515,N_17552);
nand U17793 (N_17793,N_17453,N_17456);
nand U17794 (N_17794,N_17471,N_17571);
or U17795 (N_17795,N_17422,N_17537);
nand U17796 (N_17796,N_17487,N_17594);
xnor U17797 (N_17797,N_17551,N_17527);
or U17798 (N_17798,N_17471,N_17400);
nand U17799 (N_17799,N_17512,N_17511);
and U17800 (N_17800,N_17791,N_17656);
or U17801 (N_17801,N_17754,N_17614);
and U17802 (N_17802,N_17618,N_17743);
or U17803 (N_17803,N_17790,N_17767);
or U17804 (N_17804,N_17724,N_17745);
nand U17805 (N_17805,N_17608,N_17646);
and U17806 (N_17806,N_17648,N_17616);
or U17807 (N_17807,N_17633,N_17717);
or U17808 (N_17808,N_17692,N_17715);
xor U17809 (N_17809,N_17652,N_17786);
nand U17810 (N_17810,N_17749,N_17739);
and U17811 (N_17811,N_17613,N_17702);
or U17812 (N_17812,N_17683,N_17611);
nand U17813 (N_17813,N_17780,N_17621);
or U17814 (N_17814,N_17678,N_17769);
xnor U17815 (N_17815,N_17689,N_17615);
and U17816 (N_17816,N_17737,N_17667);
or U17817 (N_17817,N_17766,N_17744);
nand U17818 (N_17818,N_17604,N_17777);
or U17819 (N_17819,N_17626,N_17703);
and U17820 (N_17820,N_17783,N_17636);
nor U17821 (N_17821,N_17758,N_17684);
nand U17822 (N_17822,N_17710,N_17778);
nand U17823 (N_17823,N_17741,N_17666);
or U17824 (N_17824,N_17610,N_17617);
or U17825 (N_17825,N_17771,N_17774);
or U17826 (N_17826,N_17619,N_17728);
nand U17827 (N_17827,N_17671,N_17627);
nor U17828 (N_17828,N_17788,N_17709);
nand U17829 (N_17829,N_17712,N_17779);
nor U17830 (N_17830,N_17696,N_17606);
nand U17831 (N_17831,N_17609,N_17649);
nand U17832 (N_17832,N_17795,N_17731);
nand U17833 (N_17833,N_17630,N_17693);
and U17834 (N_17834,N_17650,N_17768);
and U17835 (N_17835,N_17781,N_17670);
nand U17836 (N_17836,N_17668,N_17644);
xnor U17837 (N_17837,N_17775,N_17740);
and U17838 (N_17838,N_17665,N_17723);
nor U17839 (N_17839,N_17755,N_17752);
and U17840 (N_17840,N_17794,N_17759);
or U17841 (N_17841,N_17705,N_17645);
or U17842 (N_17842,N_17789,N_17699);
nor U17843 (N_17843,N_17708,N_17625);
nand U17844 (N_17844,N_17729,N_17694);
nand U17845 (N_17845,N_17716,N_17719);
nand U17846 (N_17846,N_17757,N_17772);
nor U17847 (N_17847,N_17776,N_17727);
or U17848 (N_17848,N_17661,N_17798);
and U17849 (N_17849,N_17605,N_17675);
and U17850 (N_17850,N_17647,N_17713);
nor U17851 (N_17851,N_17761,N_17762);
nand U17852 (N_17852,N_17628,N_17722);
nor U17853 (N_17853,N_17711,N_17607);
and U17854 (N_17854,N_17796,N_17688);
or U17855 (N_17855,N_17742,N_17721);
and U17856 (N_17856,N_17679,N_17706);
nand U17857 (N_17857,N_17651,N_17787);
nand U17858 (N_17858,N_17736,N_17746);
xor U17859 (N_17859,N_17756,N_17750);
or U17860 (N_17860,N_17681,N_17635);
and U17861 (N_17861,N_17748,N_17691);
or U17862 (N_17862,N_17733,N_17634);
nor U17863 (N_17863,N_17700,N_17640);
and U17864 (N_17864,N_17660,N_17738);
or U17865 (N_17865,N_17687,N_17793);
nand U17866 (N_17866,N_17674,N_17701);
nand U17867 (N_17867,N_17765,N_17718);
and U17868 (N_17868,N_17697,N_17676);
nand U17869 (N_17869,N_17695,N_17664);
and U17870 (N_17870,N_17638,N_17732);
and U17871 (N_17871,N_17654,N_17641);
xor U17872 (N_17872,N_17792,N_17799);
nor U17873 (N_17873,N_17773,N_17760);
and U17874 (N_17874,N_17631,N_17704);
or U17875 (N_17875,N_17612,N_17707);
nor U17876 (N_17876,N_17734,N_17690);
or U17877 (N_17877,N_17763,N_17686);
nand U17878 (N_17878,N_17653,N_17751);
nor U17879 (N_17879,N_17725,N_17622);
and U17880 (N_17880,N_17643,N_17632);
nand U17881 (N_17881,N_17698,N_17730);
nor U17882 (N_17882,N_17642,N_17682);
nand U17883 (N_17883,N_17669,N_17672);
nand U17884 (N_17884,N_17677,N_17714);
and U17885 (N_17885,N_17720,N_17770);
and U17886 (N_17886,N_17782,N_17680);
nand U17887 (N_17887,N_17797,N_17662);
nand U17888 (N_17888,N_17673,N_17764);
nand U17889 (N_17889,N_17639,N_17726);
nand U17890 (N_17890,N_17747,N_17753);
and U17891 (N_17891,N_17602,N_17785);
nor U17892 (N_17892,N_17735,N_17601);
nor U17893 (N_17893,N_17659,N_17685);
nor U17894 (N_17894,N_17624,N_17629);
and U17895 (N_17895,N_17655,N_17600);
nor U17896 (N_17896,N_17663,N_17623);
nor U17897 (N_17897,N_17784,N_17637);
or U17898 (N_17898,N_17658,N_17657);
nor U17899 (N_17899,N_17620,N_17603);
and U17900 (N_17900,N_17635,N_17616);
and U17901 (N_17901,N_17776,N_17721);
nor U17902 (N_17902,N_17785,N_17639);
and U17903 (N_17903,N_17615,N_17748);
xor U17904 (N_17904,N_17750,N_17700);
nor U17905 (N_17905,N_17718,N_17773);
nand U17906 (N_17906,N_17740,N_17608);
nand U17907 (N_17907,N_17705,N_17723);
and U17908 (N_17908,N_17603,N_17633);
nor U17909 (N_17909,N_17766,N_17619);
nand U17910 (N_17910,N_17605,N_17681);
nor U17911 (N_17911,N_17719,N_17602);
nand U17912 (N_17912,N_17686,N_17794);
or U17913 (N_17913,N_17794,N_17750);
and U17914 (N_17914,N_17759,N_17738);
nor U17915 (N_17915,N_17710,N_17651);
and U17916 (N_17916,N_17680,N_17761);
nand U17917 (N_17917,N_17772,N_17752);
nand U17918 (N_17918,N_17614,N_17643);
and U17919 (N_17919,N_17774,N_17605);
and U17920 (N_17920,N_17732,N_17796);
nand U17921 (N_17921,N_17717,N_17781);
nor U17922 (N_17922,N_17672,N_17630);
nor U17923 (N_17923,N_17666,N_17658);
nand U17924 (N_17924,N_17776,N_17792);
or U17925 (N_17925,N_17606,N_17749);
and U17926 (N_17926,N_17728,N_17682);
nor U17927 (N_17927,N_17761,N_17608);
nand U17928 (N_17928,N_17617,N_17651);
and U17929 (N_17929,N_17601,N_17668);
and U17930 (N_17930,N_17675,N_17699);
nand U17931 (N_17931,N_17789,N_17672);
nand U17932 (N_17932,N_17760,N_17609);
nor U17933 (N_17933,N_17708,N_17686);
or U17934 (N_17934,N_17645,N_17686);
and U17935 (N_17935,N_17623,N_17774);
or U17936 (N_17936,N_17615,N_17774);
nand U17937 (N_17937,N_17796,N_17758);
nor U17938 (N_17938,N_17664,N_17726);
nor U17939 (N_17939,N_17605,N_17642);
xor U17940 (N_17940,N_17776,N_17675);
nor U17941 (N_17941,N_17730,N_17619);
nor U17942 (N_17942,N_17770,N_17600);
or U17943 (N_17943,N_17730,N_17738);
and U17944 (N_17944,N_17770,N_17616);
xor U17945 (N_17945,N_17772,N_17711);
nor U17946 (N_17946,N_17703,N_17620);
nor U17947 (N_17947,N_17794,N_17658);
or U17948 (N_17948,N_17739,N_17627);
and U17949 (N_17949,N_17713,N_17759);
and U17950 (N_17950,N_17701,N_17770);
or U17951 (N_17951,N_17670,N_17601);
or U17952 (N_17952,N_17728,N_17641);
nor U17953 (N_17953,N_17771,N_17720);
nand U17954 (N_17954,N_17750,N_17782);
nor U17955 (N_17955,N_17695,N_17779);
nand U17956 (N_17956,N_17789,N_17681);
nand U17957 (N_17957,N_17615,N_17775);
nor U17958 (N_17958,N_17746,N_17795);
nor U17959 (N_17959,N_17755,N_17669);
and U17960 (N_17960,N_17791,N_17604);
and U17961 (N_17961,N_17786,N_17727);
nor U17962 (N_17962,N_17671,N_17615);
nor U17963 (N_17963,N_17723,N_17768);
or U17964 (N_17964,N_17717,N_17764);
nand U17965 (N_17965,N_17716,N_17635);
and U17966 (N_17966,N_17695,N_17689);
nand U17967 (N_17967,N_17699,N_17634);
or U17968 (N_17968,N_17620,N_17604);
nand U17969 (N_17969,N_17688,N_17763);
or U17970 (N_17970,N_17643,N_17762);
and U17971 (N_17971,N_17712,N_17728);
and U17972 (N_17972,N_17711,N_17635);
or U17973 (N_17973,N_17647,N_17769);
nor U17974 (N_17974,N_17751,N_17788);
or U17975 (N_17975,N_17646,N_17782);
nand U17976 (N_17976,N_17646,N_17638);
and U17977 (N_17977,N_17652,N_17690);
and U17978 (N_17978,N_17731,N_17732);
or U17979 (N_17979,N_17740,N_17727);
nand U17980 (N_17980,N_17623,N_17794);
nand U17981 (N_17981,N_17704,N_17636);
nor U17982 (N_17982,N_17711,N_17771);
nor U17983 (N_17983,N_17751,N_17676);
nor U17984 (N_17984,N_17754,N_17654);
or U17985 (N_17985,N_17623,N_17772);
nand U17986 (N_17986,N_17694,N_17681);
nor U17987 (N_17987,N_17785,N_17622);
nor U17988 (N_17988,N_17788,N_17706);
nand U17989 (N_17989,N_17747,N_17749);
nand U17990 (N_17990,N_17668,N_17740);
nand U17991 (N_17991,N_17797,N_17716);
and U17992 (N_17992,N_17699,N_17638);
and U17993 (N_17993,N_17698,N_17797);
nand U17994 (N_17994,N_17772,N_17675);
nor U17995 (N_17995,N_17615,N_17785);
nand U17996 (N_17996,N_17678,N_17633);
or U17997 (N_17997,N_17717,N_17709);
and U17998 (N_17998,N_17781,N_17793);
nor U17999 (N_17999,N_17683,N_17691);
nand U18000 (N_18000,N_17905,N_17922);
nor U18001 (N_18001,N_17947,N_17871);
nor U18002 (N_18002,N_17962,N_17920);
nand U18003 (N_18003,N_17921,N_17973);
nand U18004 (N_18004,N_17887,N_17810);
nor U18005 (N_18005,N_17833,N_17919);
nor U18006 (N_18006,N_17906,N_17896);
or U18007 (N_18007,N_17937,N_17945);
or U18008 (N_18008,N_17959,N_17889);
or U18009 (N_18009,N_17949,N_17878);
or U18010 (N_18010,N_17900,N_17943);
and U18011 (N_18011,N_17916,N_17899);
or U18012 (N_18012,N_17820,N_17873);
nor U18013 (N_18013,N_17952,N_17848);
nand U18014 (N_18014,N_17941,N_17968);
nand U18015 (N_18015,N_17998,N_17917);
nor U18016 (N_18016,N_17961,N_17802);
or U18017 (N_18017,N_17805,N_17809);
nor U18018 (N_18018,N_17825,N_17827);
nand U18019 (N_18019,N_17874,N_17865);
and U18020 (N_18020,N_17929,N_17958);
or U18021 (N_18021,N_17985,N_17880);
nand U18022 (N_18022,N_17861,N_17845);
and U18023 (N_18023,N_17898,N_17924);
and U18024 (N_18024,N_17829,N_17815);
and U18025 (N_18025,N_17976,N_17844);
or U18026 (N_18026,N_17938,N_17955);
or U18027 (N_18027,N_17866,N_17875);
and U18028 (N_18028,N_17864,N_17930);
xnor U18029 (N_18029,N_17821,N_17852);
nor U18030 (N_18030,N_17808,N_17855);
and U18031 (N_18031,N_17847,N_17860);
nor U18032 (N_18032,N_17902,N_17895);
nor U18033 (N_18033,N_17823,N_17980);
nand U18034 (N_18034,N_17806,N_17960);
nand U18035 (N_18035,N_17869,N_17926);
nand U18036 (N_18036,N_17863,N_17927);
and U18037 (N_18037,N_17867,N_17837);
nand U18038 (N_18038,N_17840,N_17939);
or U18039 (N_18039,N_17982,N_17835);
nand U18040 (N_18040,N_17836,N_17911);
nor U18041 (N_18041,N_17842,N_17963);
nand U18042 (N_18042,N_17993,N_17817);
or U18043 (N_18043,N_17944,N_17931);
nand U18044 (N_18044,N_17913,N_17872);
and U18045 (N_18045,N_17850,N_17935);
nor U18046 (N_18046,N_17977,N_17942);
and U18047 (N_18047,N_17992,N_17908);
nor U18048 (N_18048,N_17828,N_17886);
nor U18049 (N_18049,N_17834,N_17818);
or U18050 (N_18050,N_17890,N_17954);
nand U18051 (N_18051,N_17965,N_17813);
nor U18052 (N_18052,N_17975,N_17923);
nor U18053 (N_18053,N_17995,N_17849);
nand U18054 (N_18054,N_17950,N_17888);
nor U18055 (N_18055,N_17907,N_17800);
or U18056 (N_18056,N_17964,N_17918);
and U18057 (N_18057,N_17936,N_17989);
nand U18058 (N_18058,N_17925,N_17953);
or U18059 (N_18059,N_17971,N_17856);
nand U18060 (N_18060,N_17807,N_17983);
and U18061 (N_18061,N_17841,N_17996);
nor U18062 (N_18062,N_17816,N_17894);
and U18063 (N_18063,N_17981,N_17994);
nand U18064 (N_18064,N_17858,N_17811);
and U18065 (N_18065,N_17909,N_17948);
and U18066 (N_18066,N_17979,N_17897);
or U18067 (N_18067,N_17928,N_17966);
xor U18068 (N_18068,N_17804,N_17881);
nand U18069 (N_18069,N_17838,N_17999);
and U18070 (N_18070,N_17914,N_17893);
nor U18071 (N_18071,N_17969,N_17859);
nor U18072 (N_18072,N_17885,N_17870);
or U18073 (N_18073,N_17934,N_17877);
xnor U18074 (N_18074,N_17831,N_17904);
nor U18075 (N_18075,N_17997,N_17932);
and U18076 (N_18076,N_17910,N_17956);
nand U18077 (N_18077,N_17988,N_17839);
nand U18078 (N_18078,N_17933,N_17854);
or U18079 (N_18079,N_17967,N_17803);
nor U18080 (N_18080,N_17801,N_17843);
nand U18081 (N_18081,N_17903,N_17978);
nand U18082 (N_18082,N_17986,N_17846);
and U18083 (N_18083,N_17970,N_17882);
and U18084 (N_18084,N_17862,N_17912);
nand U18085 (N_18085,N_17876,N_17984);
nand U18086 (N_18086,N_17991,N_17957);
and U18087 (N_18087,N_17830,N_17819);
nor U18088 (N_18088,N_17901,N_17990);
or U18089 (N_18089,N_17832,N_17824);
nor U18090 (N_18090,N_17853,N_17940);
nand U18091 (N_18091,N_17972,N_17974);
nand U18092 (N_18092,N_17915,N_17946);
and U18093 (N_18093,N_17826,N_17814);
nor U18094 (N_18094,N_17868,N_17822);
nand U18095 (N_18095,N_17891,N_17884);
nand U18096 (N_18096,N_17892,N_17879);
or U18097 (N_18097,N_17987,N_17951);
or U18098 (N_18098,N_17851,N_17883);
nand U18099 (N_18099,N_17857,N_17812);
nand U18100 (N_18100,N_17958,N_17956);
or U18101 (N_18101,N_17975,N_17931);
or U18102 (N_18102,N_17860,N_17921);
nand U18103 (N_18103,N_17867,N_17952);
nand U18104 (N_18104,N_17918,N_17826);
nand U18105 (N_18105,N_17990,N_17927);
nor U18106 (N_18106,N_17919,N_17851);
and U18107 (N_18107,N_17963,N_17929);
and U18108 (N_18108,N_17959,N_17809);
nor U18109 (N_18109,N_17828,N_17833);
nand U18110 (N_18110,N_17884,N_17943);
and U18111 (N_18111,N_17940,N_17887);
or U18112 (N_18112,N_17830,N_17892);
nand U18113 (N_18113,N_17939,N_17867);
nand U18114 (N_18114,N_17959,N_17865);
nand U18115 (N_18115,N_17934,N_17836);
or U18116 (N_18116,N_17955,N_17807);
nand U18117 (N_18117,N_17993,N_17951);
and U18118 (N_18118,N_17920,N_17891);
nor U18119 (N_18119,N_17953,N_17985);
and U18120 (N_18120,N_17812,N_17956);
nor U18121 (N_18121,N_17824,N_17926);
or U18122 (N_18122,N_17979,N_17806);
and U18123 (N_18123,N_17907,N_17837);
and U18124 (N_18124,N_17846,N_17817);
and U18125 (N_18125,N_17848,N_17835);
or U18126 (N_18126,N_17931,N_17977);
nor U18127 (N_18127,N_17930,N_17925);
and U18128 (N_18128,N_17881,N_17970);
nor U18129 (N_18129,N_17850,N_17996);
and U18130 (N_18130,N_17936,N_17948);
or U18131 (N_18131,N_17862,N_17886);
nor U18132 (N_18132,N_17869,N_17827);
nand U18133 (N_18133,N_17804,N_17946);
and U18134 (N_18134,N_17844,N_17986);
nor U18135 (N_18135,N_17864,N_17988);
and U18136 (N_18136,N_17924,N_17984);
and U18137 (N_18137,N_17914,N_17994);
nand U18138 (N_18138,N_17816,N_17945);
nor U18139 (N_18139,N_17808,N_17986);
or U18140 (N_18140,N_17901,N_17865);
and U18141 (N_18141,N_17862,N_17973);
or U18142 (N_18142,N_17965,N_17929);
nand U18143 (N_18143,N_17930,N_17918);
and U18144 (N_18144,N_17898,N_17826);
nand U18145 (N_18145,N_17802,N_17836);
nor U18146 (N_18146,N_17804,N_17800);
nor U18147 (N_18147,N_17870,N_17812);
nand U18148 (N_18148,N_17972,N_17808);
nor U18149 (N_18149,N_17868,N_17892);
nand U18150 (N_18150,N_17973,N_17970);
and U18151 (N_18151,N_17861,N_17872);
or U18152 (N_18152,N_17850,N_17814);
nand U18153 (N_18153,N_17920,N_17979);
nor U18154 (N_18154,N_17976,N_17852);
nand U18155 (N_18155,N_17925,N_17923);
xor U18156 (N_18156,N_17986,N_17823);
or U18157 (N_18157,N_17803,N_17858);
nand U18158 (N_18158,N_17841,N_17810);
or U18159 (N_18159,N_17976,N_17858);
nand U18160 (N_18160,N_17972,N_17949);
nand U18161 (N_18161,N_17954,N_17923);
nor U18162 (N_18162,N_17860,N_17849);
nor U18163 (N_18163,N_17847,N_17882);
nor U18164 (N_18164,N_17894,N_17956);
nor U18165 (N_18165,N_17827,N_17969);
and U18166 (N_18166,N_17957,N_17810);
or U18167 (N_18167,N_17840,N_17926);
or U18168 (N_18168,N_17915,N_17876);
xnor U18169 (N_18169,N_17861,N_17964);
nor U18170 (N_18170,N_17832,N_17841);
nor U18171 (N_18171,N_17858,N_17817);
nor U18172 (N_18172,N_17973,N_17817);
xnor U18173 (N_18173,N_17869,N_17855);
nand U18174 (N_18174,N_17906,N_17892);
nand U18175 (N_18175,N_17833,N_17930);
xor U18176 (N_18176,N_17952,N_17928);
and U18177 (N_18177,N_17803,N_17832);
nand U18178 (N_18178,N_17902,N_17833);
nor U18179 (N_18179,N_17951,N_17969);
and U18180 (N_18180,N_17810,N_17899);
or U18181 (N_18181,N_17982,N_17844);
and U18182 (N_18182,N_17950,N_17808);
nor U18183 (N_18183,N_17875,N_17899);
nor U18184 (N_18184,N_17914,N_17925);
and U18185 (N_18185,N_17961,N_17804);
nor U18186 (N_18186,N_17979,N_17987);
or U18187 (N_18187,N_17837,N_17966);
nor U18188 (N_18188,N_17849,N_17983);
nand U18189 (N_18189,N_17868,N_17909);
or U18190 (N_18190,N_17861,N_17961);
nand U18191 (N_18191,N_17912,N_17964);
and U18192 (N_18192,N_17959,N_17893);
and U18193 (N_18193,N_17814,N_17959);
xor U18194 (N_18194,N_17918,N_17913);
or U18195 (N_18195,N_17867,N_17918);
and U18196 (N_18196,N_17921,N_17842);
or U18197 (N_18197,N_17878,N_17967);
nor U18198 (N_18198,N_17809,N_17995);
nor U18199 (N_18199,N_17969,N_17975);
nor U18200 (N_18200,N_18185,N_18112);
nand U18201 (N_18201,N_18107,N_18079);
nand U18202 (N_18202,N_18182,N_18068);
and U18203 (N_18203,N_18156,N_18008);
or U18204 (N_18204,N_18152,N_18189);
or U18205 (N_18205,N_18020,N_18052);
nor U18206 (N_18206,N_18061,N_18064);
nand U18207 (N_18207,N_18014,N_18188);
or U18208 (N_18208,N_18084,N_18148);
and U18209 (N_18209,N_18040,N_18081);
or U18210 (N_18210,N_18065,N_18038);
nor U18211 (N_18211,N_18173,N_18177);
nor U18212 (N_18212,N_18135,N_18066);
nor U18213 (N_18213,N_18159,N_18187);
and U18214 (N_18214,N_18138,N_18046);
and U18215 (N_18215,N_18006,N_18171);
and U18216 (N_18216,N_18158,N_18116);
and U18217 (N_18217,N_18113,N_18151);
and U18218 (N_18218,N_18060,N_18123);
nor U18219 (N_18219,N_18175,N_18047);
or U18220 (N_18220,N_18016,N_18163);
nor U18221 (N_18221,N_18125,N_18147);
or U18222 (N_18222,N_18074,N_18082);
or U18223 (N_18223,N_18161,N_18174);
nand U18224 (N_18224,N_18089,N_18190);
and U18225 (N_18225,N_18119,N_18143);
nand U18226 (N_18226,N_18098,N_18029);
nor U18227 (N_18227,N_18121,N_18166);
or U18228 (N_18228,N_18109,N_18165);
nand U18229 (N_18229,N_18067,N_18118);
nand U18230 (N_18230,N_18141,N_18128);
or U18231 (N_18231,N_18195,N_18018);
and U18232 (N_18232,N_18196,N_18051);
nor U18233 (N_18233,N_18027,N_18162);
and U18234 (N_18234,N_18150,N_18155);
or U18235 (N_18235,N_18055,N_18053);
nor U18236 (N_18236,N_18153,N_18117);
nand U18237 (N_18237,N_18180,N_18073);
and U18238 (N_18238,N_18045,N_18056);
or U18239 (N_18239,N_18160,N_18002);
and U18240 (N_18240,N_18087,N_18139);
and U18241 (N_18241,N_18086,N_18004);
or U18242 (N_18242,N_18134,N_18104);
nand U18243 (N_18243,N_18071,N_18048);
and U18244 (N_18244,N_18033,N_18194);
nand U18245 (N_18245,N_18193,N_18080);
nor U18246 (N_18246,N_18062,N_18168);
nand U18247 (N_18247,N_18090,N_18145);
and U18248 (N_18248,N_18043,N_18122);
nor U18249 (N_18249,N_18015,N_18093);
nand U18250 (N_18250,N_18179,N_18199);
and U18251 (N_18251,N_18085,N_18078);
and U18252 (N_18252,N_18176,N_18183);
or U18253 (N_18253,N_18019,N_18144);
or U18254 (N_18254,N_18026,N_18032);
and U18255 (N_18255,N_18181,N_18111);
and U18256 (N_18256,N_18088,N_18039);
and U18257 (N_18257,N_18131,N_18164);
or U18258 (N_18258,N_18096,N_18025);
nand U18259 (N_18259,N_18091,N_18154);
or U18260 (N_18260,N_18169,N_18110);
xnor U18261 (N_18261,N_18167,N_18184);
nor U18262 (N_18262,N_18009,N_18021);
nand U18263 (N_18263,N_18044,N_18013);
or U18264 (N_18264,N_18120,N_18108);
and U18265 (N_18265,N_18100,N_18102);
nor U18266 (N_18266,N_18172,N_18010);
and U18267 (N_18267,N_18037,N_18129);
or U18268 (N_18268,N_18124,N_18005);
and U18269 (N_18269,N_18149,N_18069);
nor U18270 (N_18270,N_18022,N_18140);
or U18271 (N_18271,N_18028,N_18198);
nand U18272 (N_18272,N_18103,N_18178);
and U18273 (N_18273,N_18105,N_18035);
and U18274 (N_18274,N_18097,N_18063);
nor U18275 (N_18275,N_18000,N_18083);
nor U18276 (N_18276,N_18126,N_18092);
nand U18277 (N_18277,N_18142,N_18030);
nor U18278 (N_18278,N_18114,N_18049);
nand U18279 (N_18279,N_18192,N_18099);
nor U18280 (N_18280,N_18031,N_18072);
nor U18281 (N_18281,N_18170,N_18001);
nand U18282 (N_18282,N_18095,N_18137);
nor U18283 (N_18283,N_18017,N_18057);
nor U18284 (N_18284,N_18136,N_18050);
and U18285 (N_18285,N_18003,N_18197);
nand U18286 (N_18286,N_18075,N_18146);
nor U18287 (N_18287,N_18186,N_18036);
or U18288 (N_18288,N_18094,N_18133);
nand U18289 (N_18289,N_18101,N_18023);
nor U18290 (N_18290,N_18191,N_18058);
nor U18291 (N_18291,N_18034,N_18070);
or U18292 (N_18292,N_18130,N_18012);
or U18293 (N_18293,N_18077,N_18041);
nand U18294 (N_18294,N_18115,N_18011);
xor U18295 (N_18295,N_18076,N_18007);
or U18296 (N_18296,N_18024,N_18042);
nand U18297 (N_18297,N_18059,N_18157);
nand U18298 (N_18298,N_18106,N_18132);
and U18299 (N_18299,N_18127,N_18054);
or U18300 (N_18300,N_18083,N_18064);
and U18301 (N_18301,N_18189,N_18079);
and U18302 (N_18302,N_18179,N_18088);
and U18303 (N_18303,N_18072,N_18055);
nand U18304 (N_18304,N_18086,N_18084);
nand U18305 (N_18305,N_18013,N_18061);
and U18306 (N_18306,N_18104,N_18052);
or U18307 (N_18307,N_18183,N_18135);
nand U18308 (N_18308,N_18120,N_18149);
and U18309 (N_18309,N_18113,N_18115);
and U18310 (N_18310,N_18155,N_18078);
nor U18311 (N_18311,N_18065,N_18125);
and U18312 (N_18312,N_18027,N_18097);
and U18313 (N_18313,N_18137,N_18021);
and U18314 (N_18314,N_18169,N_18138);
or U18315 (N_18315,N_18193,N_18161);
and U18316 (N_18316,N_18048,N_18028);
nand U18317 (N_18317,N_18026,N_18119);
and U18318 (N_18318,N_18191,N_18082);
and U18319 (N_18319,N_18093,N_18148);
nor U18320 (N_18320,N_18115,N_18057);
nand U18321 (N_18321,N_18127,N_18020);
and U18322 (N_18322,N_18094,N_18074);
nand U18323 (N_18323,N_18141,N_18138);
nand U18324 (N_18324,N_18084,N_18166);
or U18325 (N_18325,N_18148,N_18023);
and U18326 (N_18326,N_18095,N_18143);
nand U18327 (N_18327,N_18166,N_18111);
nand U18328 (N_18328,N_18066,N_18170);
and U18329 (N_18329,N_18186,N_18168);
nand U18330 (N_18330,N_18153,N_18144);
and U18331 (N_18331,N_18157,N_18118);
or U18332 (N_18332,N_18094,N_18160);
nor U18333 (N_18333,N_18138,N_18068);
and U18334 (N_18334,N_18128,N_18003);
xnor U18335 (N_18335,N_18027,N_18095);
nor U18336 (N_18336,N_18132,N_18033);
nand U18337 (N_18337,N_18061,N_18124);
or U18338 (N_18338,N_18144,N_18086);
or U18339 (N_18339,N_18097,N_18021);
nor U18340 (N_18340,N_18038,N_18112);
nor U18341 (N_18341,N_18141,N_18186);
nor U18342 (N_18342,N_18004,N_18194);
or U18343 (N_18343,N_18025,N_18149);
or U18344 (N_18344,N_18088,N_18122);
nand U18345 (N_18345,N_18194,N_18083);
nor U18346 (N_18346,N_18016,N_18034);
nor U18347 (N_18347,N_18138,N_18121);
or U18348 (N_18348,N_18164,N_18184);
nor U18349 (N_18349,N_18109,N_18121);
nand U18350 (N_18350,N_18122,N_18080);
nand U18351 (N_18351,N_18088,N_18124);
nor U18352 (N_18352,N_18003,N_18145);
nand U18353 (N_18353,N_18009,N_18046);
nand U18354 (N_18354,N_18144,N_18035);
and U18355 (N_18355,N_18167,N_18008);
and U18356 (N_18356,N_18011,N_18090);
nor U18357 (N_18357,N_18048,N_18184);
or U18358 (N_18358,N_18182,N_18032);
nor U18359 (N_18359,N_18044,N_18167);
and U18360 (N_18360,N_18197,N_18010);
nand U18361 (N_18361,N_18119,N_18187);
or U18362 (N_18362,N_18039,N_18114);
and U18363 (N_18363,N_18031,N_18035);
nand U18364 (N_18364,N_18030,N_18123);
nor U18365 (N_18365,N_18053,N_18132);
nand U18366 (N_18366,N_18132,N_18028);
nand U18367 (N_18367,N_18105,N_18054);
xor U18368 (N_18368,N_18080,N_18139);
or U18369 (N_18369,N_18142,N_18157);
or U18370 (N_18370,N_18154,N_18122);
nor U18371 (N_18371,N_18040,N_18048);
nand U18372 (N_18372,N_18034,N_18033);
nor U18373 (N_18373,N_18092,N_18134);
nor U18374 (N_18374,N_18180,N_18003);
nand U18375 (N_18375,N_18018,N_18178);
nand U18376 (N_18376,N_18022,N_18163);
and U18377 (N_18377,N_18136,N_18078);
nor U18378 (N_18378,N_18007,N_18056);
nor U18379 (N_18379,N_18085,N_18133);
or U18380 (N_18380,N_18142,N_18041);
or U18381 (N_18381,N_18067,N_18130);
nand U18382 (N_18382,N_18175,N_18016);
and U18383 (N_18383,N_18145,N_18155);
or U18384 (N_18384,N_18035,N_18117);
nand U18385 (N_18385,N_18133,N_18028);
nand U18386 (N_18386,N_18088,N_18028);
and U18387 (N_18387,N_18029,N_18146);
and U18388 (N_18388,N_18191,N_18124);
nand U18389 (N_18389,N_18017,N_18174);
xor U18390 (N_18390,N_18015,N_18120);
or U18391 (N_18391,N_18180,N_18123);
or U18392 (N_18392,N_18065,N_18046);
or U18393 (N_18393,N_18122,N_18066);
nor U18394 (N_18394,N_18138,N_18090);
xor U18395 (N_18395,N_18086,N_18172);
or U18396 (N_18396,N_18061,N_18087);
nor U18397 (N_18397,N_18023,N_18010);
nand U18398 (N_18398,N_18086,N_18089);
nor U18399 (N_18399,N_18110,N_18038);
nand U18400 (N_18400,N_18328,N_18350);
and U18401 (N_18401,N_18234,N_18275);
and U18402 (N_18402,N_18296,N_18207);
nand U18403 (N_18403,N_18363,N_18397);
and U18404 (N_18404,N_18264,N_18360);
nor U18405 (N_18405,N_18390,N_18210);
nor U18406 (N_18406,N_18224,N_18321);
nand U18407 (N_18407,N_18288,N_18374);
and U18408 (N_18408,N_18212,N_18385);
or U18409 (N_18409,N_18308,N_18380);
nor U18410 (N_18410,N_18272,N_18266);
nand U18411 (N_18411,N_18364,N_18230);
and U18412 (N_18412,N_18261,N_18376);
and U18413 (N_18413,N_18244,N_18311);
nor U18414 (N_18414,N_18344,N_18333);
nand U18415 (N_18415,N_18388,N_18375);
xor U18416 (N_18416,N_18250,N_18370);
and U18417 (N_18417,N_18218,N_18367);
and U18418 (N_18418,N_18322,N_18359);
nor U18419 (N_18419,N_18372,N_18211);
or U18420 (N_18420,N_18271,N_18317);
and U18421 (N_18421,N_18365,N_18209);
nor U18422 (N_18422,N_18253,N_18294);
nand U18423 (N_18423,N_18251,N_18238);
nand U18424 (N_18424,N_18320,N_18340);
and U18425 (N_18425,N_18221,N_18245);
nor U18426 (N_18426,N_18203,N_18304);
or U18427 (N_18427,N_18289,N_18237);
nor U18428 (N_18428,N_18332,N_18213);
nor U18429 (N_18429,N_18273,N_18260);
nor U18430 (N_18430,N_18287,N_18232);
or U18431 (N_18431,N_18334,N_18291);
and U18432 (N_18432,N_18371,N_18307);
or U18433 (N_18433,N_18248,N_18348);
nand U18434 (N_18434,N_18368,N_18356);
nor U18435 (N_18435,N_18231,N_18341);
or U18436 (N_18436,N_18262,N_18293);
or U18437 (N_18437,N_18292,N_18353);
nand U18438 (N_18438,N_18373,N_18338);
and U18439 (N_18439,N_18267,N_18270);
xnor U18440 (N_18440,N_18269,N_18255);
or U18441 (N_18441,N_18278,N_18243);
and U18442 (N_18442,N_18240,N_18205);
nand U18443 (N_18443,N_18215,N_18279);
and U18444 (N_18444,N_18301,N_18241);
or U18445 (N_18445,N_18233,N_18393);
nor U18446 (N_18446,N_18314,N_18217);
and U18447 (N_18447,N_18227,N_18327);
nand U18448 (N_18448,N_18225,N_18343);
and U18449 (N_18449,N_18208,N_18305);
nor U18450 (N_18450,N_18220,N_18357);
and U18451 (N_18451,N_18362,N_18342);
or U18452 (N_18452,N_18265,N_18242);
and U18453 (N_18453,N_18335,N_18202);
nand U18454 (N_18454,N_18358,N_18249);
and U18455 (N_18455,N_18354,N_18223);
nand U18456 (N_18456,N_18313,N_18377);
and U18457 (N_18457,N_18214,N_18396);
or U18458 (N_18458,N_18299,N_18226);
nand U18459 (N_18459,N_18298,N_18206);
nor U18460 (N_18460,N_18325,N_18352);
or U18461 (N_18461,N_18331,N_18235);
and U18462 (N_18462,N_18349,N_18310);
nor U18463 (N_18463,N_18336,N_18236);
or U18464 (N_18464,N_18200,N_18306);
nand U18465 (N_18465,N_18222,N_18398);
and U18466 (N_18466,N_18201,N_18295);
nor U18467 (N_18467,N_18346,N_18395);
and U18468 (N_18468,N_18285,N_18254);
and U18469 (N_18469,N_18282,N_18394);
and U18470 (N_18470,N_18284,N_18229);
and U18471 (N_18471,N_18309,N_18326);
and U18472 (N_18472,N_18280,N_18392);
nand U18473 (N_18473,N_18361,N_18247);
and U18474 (N_18474,N_18323,N_18258);
and U18475 (N_18475,N_18399,N_18312);
nor U18476 (N_18476,N_18339,N_18378);
nor U18477 (N_18477,N_18274,N_18281);
nor U18478 (N_18478,N_18246,N_18386);
nand U18479 (N_18479,N_18382,N_18263);
and U18480 (N_18480,N_18257,N_18276);
xnor U18481 (N_18481,N_18297,N_18239);
nor U18482 (N_18482,N_18391,N_18381);
nand U18483 (N_18483,N_18351,N_18366);
and U18484 (N_18484,N_18345,N_18318);
nand U18485 (N_18485,N_18355,N_18319);
or U18486 (N_18486,N_18369,N_18384);
nand U18487 (N_18487,N_18383,N_18316);
nor U18488 (N_18488,N_18303,N_18389);
nor U18489 (N_18489,N_18290,N_18315);
nand U18490 (N_18490,N_18329,N_18216);
and U18491 (N_18491,N_18286,N_18268);
xor U18492 (N_18492,N_18324,N_18330);
or U18493 (N_18493,N_18277,N_18259);
nand U18494 (N_18494,N_18300,N_18379);
or U18495 (N_18495,N_18387,N_18228);
and U18496 (N_18496,N_18219,N_18204);
nand U18497 (N_18497,N_18337,N_18252);
nand U18498 (N_18498,N_18302,N_18256);
nor U18499 (N_18499,N_18347,N_18283);
nor U18500 (N_18500,N_18307,N_18381);
or U18501 (N_18501,N_18209,N_18381);
or U18502 (N_18502,N_18396,N_18378);
nor U18503 (N_18503,N_18340,N_18262);
or U18504 (N_18504,N_18213,N_18269);
and U18505 (N_18505,N_18314,N_18283);
or U18506 (N_18506,N_18364,N_18302);
xnor U18507 (N_18507,N_18255,N_18303);
and U18508 (N_18508,N_18302,N_18376);
nand U18509 (N_18509,N_18306,N_18371);
and U18510 (N_18510,N_18223,N_18316);
nand U18511 (N_18511,N_18236,N_18275);
or U18512 (N_18512,N_18209,N_18235);
nand U18513 (N_18513,N_18219,N_18344);
and U18514 (N_18514,N_18326,N_18339);
nand U18515 (N_18515,N_18226,N_18385);
and U18516 (N_18516,N_18285,N_18362);
nand U18517 (N_18517,N_18372,N_18379);
and U18518 (N_18518,N_18292,N_18253);
nor U18519 (N_18519,N_18397,N_18239);
nor U18520 (N_18520,N_18287,N_18360);
nand U18521 (N_18521,N_18387,N_18333);
or U18522 (N_18522,N_18334,N_18374);
nor U18523 (N_18523,N_18361,N_18323);
nand U18524 (N_18524,N_18213,N_18271);
and U18525 (N_18525,N_18316,N_18399);
nand U18526 (N_18526,N_18226,N_18313);
or U18527 (N_18527,N_18390,N_18264);
and U18528 (N_18528,N_18331,N_18204);
nand U18529 (N_18529,N_18301,N_18203);
and U18530 (N_18530,N_18393,N_18350);
xnor U18531 (N_18531,N_18215,N_18345);
nand U18532 (N_18532,N_18266,N_18383);
nor U18533 (N_18533,N_18226,N_18324);
or U18534 (N_18534,N_18372,N_18316);
nand U18535 (N_18535,N_18351,N_18365);
and U18536 (N_18536,N_18368,N_18351);
nor U18537 (N_18537,N_18221,N_18302);
or U18538 (N_18538,N_18275,N_18360);
and U18539 (N_18539,N_18252,N_18359);
or U18540 (N_18540,N_18257,N_18336);
nand U18541 (N_18541,N_18238,N_18212);
nor U18542 (N_18542,N_18388,N_18234);
xnor U18543 (N_18543,N_18372,N_18356);
and U18544 (N_18544,N_18229,N_18244);
nor U18545 (N_18545,N_18381,N_18212);
and U18546 (N_18546,N_18226,N_18200);
nand U18547 (N_18547,N_18375,N_18315);
nor U18548 (N_18548,N_18292,N_18319);
nand U18549 (N_18549,N_18201,N_18365);
or U18550 (N_18550,N_18299,N_18237);
and U18551 (N_18551,N_18257,N_18271);
and U18552 (N_18552,N_18270,N_18289);
nand U18553 (N_18553,N_18308,N_18392);
or U18554 (N_18554,N_18263,N_18316);
nor U18555 (N_18555,N_18386,N_18345);
and U18556 (N_18556,N_18366,N_18236);
and U18557 (N_18557,N_18346,N_18384);
and U18558 (N_18558,N_18250,N_18200);
nor U18559 (N_18559,N_18394,N_18374);
or U18560 (N_18560,N_18203,N_18332);
or U18561 (N_18561,N_18203,N_18335);
nor U18562 (N_18562,N_18361,N_18243);
nand U18563 (N_18563,N_18299,N_18322);
or U18564 (N_18564,N_18329,N_18305);
nand U18565 (N_18565,N_18357,N_18299);
nand U18566 (N_18566,N_18202,N_18214);
nor U18567 (N_18567,N_18345,N_18374);
or U18568 (N_18568,N_18365,N_18312);
xor U18569 (N_18569,N_18212,N_18339);
nor U18570 (N_18570,N_18398,N_18297);
nor U18571 (N_18571,N_18239,N_18376);
nand U18572 (N_18572,N_18295,N_18220);
nor U18573 (N_18573,N_18338,N_18361);
or U18574 (N_18574,N_18314,N_18293);
and U18575 (N_18575,N_18228,N_18264);
or U18576 (N_18576,N_18380,N_18317);
and U18577 (N_18577,N_18339,N_18334);
or U18578 (N_18578,N_18204,N_18207);
nand U18579 (N_18579,N_18324,N_18395);
nor U18580 (N_18580,N_18202,N_18394);
and U18581 (N_18581,N_18249,N_18387);
nand U18582 (N_18582,N_18259,N_18289);
and U18583 (N_18583,N_18337,N_18310);
nand U18584 (N_18584,N_18396,N_18275);
and U18585 (N_18585,N_18354,N_18362);
nor U18586 (N_18586,N_18356,N_18337);
and U18587 (N_18587,N_18301,N_18345);
and U18588 (N_18588,N_18312,N_18227);
or U18589 (N_18589,N_18261,N_18217);
nor U18590 (N_18590,N_18307,N_18266);
and U18591 (N_18591,N_18248,N_18216);
nor U18592 (N_18592,N_18349,N_18309);
or U18593 (N_18593,N_18205,N_18322);
nand U18594 (N_18594,N_18356,N_18304);
and U18595 (N_18595,N_18266,N_18372);
and U18596 (N_18596,N_18279,N_18288);
or U18597 (N_18597,N_18365,N_18214);
nand U18598 (N_18598,N_18239,N_18374);
nand U18599 (N_18599,N_18339,N_18255);
or U18600 (N_18600,N_18451,N_18415);
or U18601 (N_18601,N_18544,N_18527);
and U18602 (N_18602,N_18556,N_18455);
or U18603 (N_18603,N_18557,N_18576);
nand U18604 (N_18604,N_18432,N_18426);
nand U18605 (N_18605,N_18550,N_18508);
or U18606 (N_18606,N_18506,N_18524);
and U18607 (N_18607,N_18536,N_18486);
nor U18608 (N_18608,N_18420,N_18489);
or U18609 (N_18609,N_18554,N_18428);
nand U18610 (N_18610,N_18439,N_18463);
nand U18611 (N_18611,N_18456,N_18573);
and U18612 (N_18612,N_18440,N_18492);
and U18613 (N_18613,N_18413,N_18582);
nand U18614 (N_18614,N_18497,N_18484);
or U18615 (N_18615,N_18520,N_18410);
or U18616 (N_18616,N_18470,N_18476);
nor U18617 (N_18617,N_18584,N_18490);
nor U18618 (N_18618,N_18472,N_18560);
nor U18619 (N_18619,N_18553,N_18412);
and U18620 (N_18620,N_18504,N_18485);
or U18621 (N_18621,N_18521,N_18431);
nand U18622 (N_18622,N_18534,N_18568);
nor U18623 (N_18623,N_18462,N_18468);
nor U18624 (N_18624,N_18575,N_18477);
and U18625 (N_18625,N_18459,N_18475);
nand U18626 (N_18626,N_18599,N_18539);
nand U18627 (N_18627,N_18518,N_18454);
or U18628 (N_18628,N_18586,N_18501);
or U18629 (N_18629,N_18530,N_18532);
or U18630 (N_18630,N_18466,N_18558);
nor U18631 (N_18631,N_18437,N_18494);
and U18632 (N_18632,N_18595,N_18538);
nand U18633 (N_18633,N_18419,N_18562);
xor U18634 (N_18634,N_18414,N_18563);
nand U18635 (N_18635,N_18528,N_18421);
or U18636 (N_18636,N_18591,N_18555);
nand U18637 (N_18637,N_18552,N_18479);
nor U18638 (N_18638,N_18445,N_18404);
nor U18639 (N_18639,N_18469,N_18511);
nor U18640 (N_18640,N_18549,N_18408);
nor U18641 (N_18641,N_18467,N_18525);
or U18642 (N_18642,N_18537,N_18516);
or U18643 (N_18643,N_18429,N_18403);
or U18644 (N_18644,N_18400,N_18566);
nand U18645 (N_18645,N_18487,N_18409);
or U18646 (N_18646,N_18502,N_18424);
and U18647 (N_18647,N_18513,N_18590);
nor U18648 (N_18648,N_18517,N_18448);
nor U18649 (N_18649,N_18540,N_18416);
or U18650 (N_18650,N_18567,N_18510);
or U18651 (N_18651,N_18594,N_18541);
nand U18652 (N_18652,N_18509,N_18435);
nor U18653 (N_18653,N_18401,N_18441);
nor U18654 (N_18654,N_18418,N_18458);
and U18655 (N_18655,N_18457,N_18425);
nand U18656 (N_18656,N_18491,N_18433);
or U18657 (N_18657,N_18499,N_18593);
xor U18658 (N_18658,N_18587,N_18507);
nor U18659 (N_18659,N_18407,N_18514);
nand U18660 (N_18660,N_18453,N_18564);
or U18661 (N_18661,N_18482,N_18411);
nor U18662 (N_18662,N_18548,N_18446);
or U18663 (N_18663,N_18559,N_18512);
and U18664 (N_18664,N_18434,N_18522);
or U18665 (N_18665,N_18542,N_18585);
nor U18666 (N_18666,N_18583,N_18447);
and U18667 (N_18667,N_18464,N_18452);
and U18668 (N_18668,N_18450,N_18526);
and U18669 (N_18669,N_18589,N_18442);
or U18670 (N_18670,N_18438,N_18543);
or U18671 (N_18671,N_18523,N_18444);
or U18672 (N_18672,N_18460,N_18496);
nor U18673 (N_18673,N_18579,N_18465);
and U18674 (N_18674,N_18443,N_18529);
and U18675 (N_18675,N_18474,N_18580);
nor U18676 (N_18676,N_18581,N_18545);
or U18677 (N_18677,N_18597,N_18570);
and U18678 (N_18678,N_18461,N_18473);
nand U18679 (N_18679,N_18533,N_18596);
nand U18680 (N_18680,N_18498,N_18436);
nor U18681 (N_18681,N_18519,N_18449);
or U18682 (N_18682,N_18423,N_18480);
nand U18683 (N_18683,N_18572,N_18500);
or U18684 (N_18684,N_18481,N_18471);
nor U18685 (N_18685,N_18571,N_18577);
nand U18686 (N_18686,N_18483,N_18495);
and U18687 (N_18687,N_18578,N_18488);
and U18688 (N_18688,N_18505,N_18592);
or U18689 (N_18689,N_18598,N_18574);
nor U18690 (N_18690,N_18547,N_18503);
or U18691 (N_18691,N_18551,N_18561);
nand U18692 (N_18692,N_18478,N_18588);
nor U18693 (N_18693,N_18405,N_18493);
and U18694 (N_18694,N_18406,N_18422);
or U18695 (N_18695,N_18569,N_18535);
xnor U18696 (N_18696,N_18430,N_18546);
and U18697 (N_18697,N_18531,N_18565);
nor U18698 (N_18698,N_18427,N_18402);
and U18699 (N_18699,N_18515,N_18417);
or U18700 (N_18700,N_18533,N_18495);
or U18701 (N_18701,N_18583,N_18530);
or U18702 (N_18702,N_18456,N_18526);
nor U18703 (N_18703,N_18546,N_18490);
or U18704 (N_18704,N_18544,N_18486);
nand U18705 (N_18705,N_18487,N_18539);
nor U18706 (N_18706,N_18452,N_18511);
and U18707 (N_18707,N_18473,N_18411);
nor U18708 (N_18708,N_18471,N_18446);
and U18709 (N_18709,N_18545,N_18424);
nand U18710 (N_18710,N_18572,N_18527);
nor U18711 (N_18711,N_18562,N_18507);
nand U18712 (N_18712,N_18464,N_18514);
or U18713 (N_18713,N_18511,N_18433);
and U18714 (N_18714,N_18593,N_18536);
and U18715 (N_18715,N_18553,N_18597);
or U18716 (N_18716,N_18422,N_18497);
and U18717 (N_18717,N_18412,N_18537);
nand U18718 (N_18718,N_18574,N_18522);
or U18719 (N_18719,N_18560,N_18480);
or U18720 (N_18720,N_18470,N_18536);
or U18721 (N_18721,N_18401,N_18488);
nor U18722 (N_18722,N_18551,N_18423);
nor U18723 (N_18723,N_18455,N_18487);
nor U18724 (N_18724,N_18499,N_18458);
nand U18725 (N_18725,N_18578,N_18400);
nor U18726 (N_18726,N_18464,N_18560);
nand U18727 (N_18727,N_18436,N_18562);
and U18728 (N_18728,N_18405,N_18534);
or U18729 (N_18729,N_18572,N_18592);
xnor U18730 (N_18730,N_18493,N_18575);
nand U18731 (N_18731,N_18588,N_18524);
or U18732 (N_18732,N_18582,N_18536);
nor U18733 (N_18733,N_18553,N_18492);
nor U18734 (N_18734,N_18412,N_18509);
or U18735 (N_18735,N_18520,N_18593);
nand U18736 (N_18736,N_18457,N_18501);
nor U18737 (N_18737,N_18555,N_18546);
and U18738 (N_18738,N_18411,N_18517);
and U18739 (N_18739,N_18494,N_18477);
nor U18740 (N_18740,N_18401,N_18554);
nor U18741 (N_18741,N_18593,N_18464);
and U18742 (N_18742,N_18451,N_18589);
xor U18743 (N_18743,N_18528,N_18512);
xnor U18744 (N_18744,N_18530,N_18450);
and U18745 (N_18745,N_18561,N_18447);
and U18746 (N_18746,N_18425,N_18552);
nand U18747 (N_18747,N_18586,N_18538);
or U18748 (N_18748,N_18508,N_18582);
nor U18749 (N_18749,N_18505,N_18456);
nand U18750 (N_18750,N_18469,N_18466);
nor U18751 (N_18751,N_18440,N_18507);
or U18752 (N_18752,N_18548,N_18448);
nand U18753 (N_18753,N_18404,N_18475);
nor U18754 (N_18754,N_18407,N_18420);
nand U18755 (N_18755,N_18523,N_18572);
or U18756 (N_18756,N_18422,N_18525);
xnor U18757 (N_18757,N_18599,N_18468);
or U18758 (N_18758,N_18534,N_18502);
or U18759 (N_18759,N_18422,N_18524);
nor U18760 (N_18760,N_18492,N_18434);
and U18761 (N_18761,N_18407,N_18425);
nor U18762 (N_18762,N_18533,N_18434);
nor U18763 (N_18763,N_18420,N_18495);
and U18764 (N_18764,N_18538,N_18511);
xnor U18765 (N_18765,N_18555,N_18500);
nor U18766 (N_18766,N_18506,N_18573);
and U18767 (N_18767,N_18546,N_18441);
nand U18768 (N_18768,N_18595,N_18481);
and U18769 (N_18769,N_18535,N_18471);
nor U18770 (N_18770,N_18445,N_18479);
nand U18771 (N_18771,N_18565,N_18533);
nor U18772 (N_18772,N_18541,N_18490);
and U18773 (N_18773,N_18423,N_18553);
or U18774 (N_18774,N_18447,N_18574);
and U18775 (N_18775,N_18480,N_18559);
and U18776 (N_18776,N_18465,N_18591);
nor U18777 (N_18777,N_18441,N_18544);
or U18778 (N_18778,N_18440,N_18546);
nor U18779 (N_18779,N_18457,N_18539);
or U18780 (N_18780,N_18564,N_18436);
or U18781 (N_18781,N_18416,N_18454);
or U18782 (N_18782,N_18450,N_18562);
nor U18783 (N_18783,N_18561,N_18583);
nor U18784 (N_18784,N_18535,N_18582);
and U18785 (N_18785,N_18561,N_18545);
nand U18786 (N_18786,N_18430,N_18465);
nand U18787 (N_18787,N_18446,N_18468);
nand U18788 (N_18788,N_18472,N_18580);
nor U18789 (N_18789,N_18575,N_18447);
or U18790 (N_18790,N_18462,N_18572);
nand U18791 (N_18791,N_18484,N_18534);
nand U18792 (N_18792,N_18518,N_18544);
and U18793 (N_18793,N_18595,N_18495);
and U18794 (N_18794,N_18579,N_18410);
or U18795 (N_18795,N_18415,N_18574);
nand U18796 (N_18796,N_18457,N_18573);
nor U18797 (N_18797,N_18559,N_18506);
or U18798 (N_18798,N_18432,N_18404);
nor U18799 (N_18799,N_18485,N_18437);
and U18800 (N_18800,N_18671,N_18603);
and U18801 (N_18801,N_18758,N_18685);
or U18802 (N_18802,N_18750,N_18627);
nor U18803 (N_18803,N_18609,N_18667);
nor U18804 (N_18804,N_18751,N_18770);
and U18805 (N_18805,N_18753,N_18641);
nor U18806 (N_18806,N_18654,N_18749);
or U18807 (N_18807,N_18767,N_18720);
nor U18808 (N_18808,N_18612,N_18786);
nand U18809 (N_18809,N_18707,N_18785);
nand U18810 (N_18810,N_18775,N_18634);
nand U18811 (N_18811,N_18605,N_18730);
and U18812 (N_18812,N_18613,N_18788);
and U18813 (N_18813,N_18742,N_18660);
nor U18814 (N_18814,N_18732,N_18664);
nor U18815 (N_18815,N_18624,N_18793);
and U18816 (N_18816,N_18661,N_18608);
or U18817 (N_18817,N_18737,N_18681);
and U18818 (N_18818,N_18666,N_18690);
nor U18819 (N_18819,N_18616,N_18650);
nor U18820 (N_18820,N_18714,N_18683);
or U18821 (N_18821,N_18710,N_18630);
nand U18822 (N_18822,N_18643,N_18761);
or U18823 (N_18823,N_18665,N_18736);
nand U18824 (N_18824,N_18629,N_18735);
or U18825 (N_18825,N_18653,N_18697);
nand U18826 (N_18826,N_18620,N_18618);
nand U18827 (N_18827,N_18734,N_18676);
or U18828 (N_18828,N_18696,N_18722);
nand U18829 (N_18829,N_18670,N_18717);
and U18830 (N_18830,N_18792,N_18600);
nor U18831 (N_18831,N_18674,N_18790);
nand U18832 (N_18832,N_18798,N_18655);
and U18833 (N_18833,N_18648,N_18748);
nand U18834 (N_18834,N_18754,N_18617);
and U18835 (N_18835,N_18614,N_18672);
nor U18836 (N_18836,N_18619,N_18724);
or U18837 (N_18837,N_18773,N_18601);
nand U18838 (N_18838,N_18662,N_18708);
and U18839 (N_18839,N_18631,N_18623);
nand U18840 (N_18840,N_18606,N_18760);
or U18841 (N_18841,N_18728,N_18621);
nand U18842 (N_18842,N_18778,N_18731);
nand U18843 (N_18843,N_18702,N_18698);
nor U18844 (N_18844,N_18649,N_18628);
or U18845 (N_18845,N_18658,N_18763);
and U18846 (N_18846,N_18700,N_18782);
nand U18847 (N_18847,N_18765,N_18604);
nor U18848 (N_18848,N_18689,N_18783);
nor U18849 (N_18849,N_18715,N_18680);
or U18850 (N_18850,N_18729,N_18651);
xor U18851 (N_18851,N_18602,N_18686);
nand U18852 (N_18852,N_18727,N_18644);
nor U18853 (N_18853,N_18647,N_18639);
nor U18854 (N_18854,N_18759,N_18733);
or U18855 (N_18855,N_18757,N_18615);
or U18856 (N_18856,N_18646,N_18688);
xor U18857 (N_18857,N_18622,N_18743);
nand U18858 (N_18858,N_18699,N_18755);
and U18859 (N_18859,N_18723,N_18725);
nor U18860 (N_18860,N_18679,N_18797);
nand U18861 (N_18861,N_18745,N_18721);
or U18862 (N_18862,N_18633,N_18640);
nor U18863 (N_18863,N_18626,N_18693);
nor U18864 (N_18864,N_18675,N_18668);
nor U18865 (N_18865,N_18692,N_18771);
or U18866 (N_18866,N_18796,N_18764);
and U18867 (N_18867,N_18645,N_18718);
and U18868 (N_18868,N_18752,N_18784);
or U18869 (N_18869,N_18787,N_18789);
nand U18870 (N_18870,N_18611,N_18704);
or U18871 (N_18871,N_18780,N_18659);
or U18872 (N_18872,N_18768,N_18632);
and U18873 (N_18873,N_18781,N_18772);
and U18874 (N_18874,N_18687,N_18779);
nand U18875 (N_18875,N_18794,N_18791);
nor U18876 (N_18876,N_18695,N_18774);
or U18877 (N_18877,N_18756,N_18610);
and U18878 (N_18878,N_18673,N_18677);
or U18879 (N_18879,N_18682,N_18625);
nand U18880 (N_18880,N_18739,N_18636);
nand U18881 (N_18881,N_18706,N_18777);
and U18882 (N_18882,N_18711,N_18642);
and U18883 (N_18883,N_18656,N_18607);
nand U18884 (N_18884,N_18726,N_18691);
nor U18885 (N_18885,N_18746,N_18766);
or U18886 (N_18886,N_18694,N_18678);
nor U18887 (N_18887,N_18740,N_18709);
or U18888 (N_18888,N_18712,N_18652);
nand U18889 (N_18889,N_18663,N_18747);
nand U18890 (N_18890,N_18762,N_18738);
nor U18891 (N_18891,N_18635,N_18799);
nor U18892 (N_18892,N_18719,N_18684);
and U18893 (N_18893,N_18741,N_18657);
nor U18894 (N_18894,N_18769,N_18637);
and U18895 (N_18895,N_18701,N_18669);
nand U18896 (N_18896,N_18638,N_18744);
and U18897 (N_18897,N_18716,N_18795);
or U18898 (N_18898,N_18703,N_18776);
nand U18899 (N_18899,N_18713,N_18705);
and U18900 (N_18900,N_18797,N_18669);
nor U18901 (N_18901,N_18757,N_18702);
nor U18902 (N_18902,N_18638,N_18795);
nor U18903 (N_18903,N_18703,N_18790);
and U18904 (N_18904,N_18741,N_18652);
or U18905 (N_18905,N_18748,N_18795);
nor U18906 (N_18906,N_18700,N_18697);
and U18907 (N_18907,N_18616,N_18767);
or U18908 (N_18908,N_18741,N_18650);
and U18909 (N_18909,N_18708,N_18725);
nand U18910 (N_18910,N_18667,N_18695);
nand U18911 (N_18911,N_18746,N_18743);
nor U18912 (N_18912,N_18760,N_18662);
nor U18913 (N_18913,N_18657,N_18723);
nor U18914 (N_18914,N_18779,N_18676);
and U18915 (N_18915,N_18698,N_18658);
nor U18916 (N_18916,N_18617,N_18651);
and U18917 (N_18917,N_18753,N_18610);
and U18918 (N_18918,N_18776,N_18779);
nor U18919 (N_18919,N_18796,N_18684);
or U18920 (N_18920,N_18677,N_18707);
and U18921 (N_18921,N_18725,N_18721);
or U18922 (N_18922,N_18766,N_18794);
nor U18923 (N_18923,N_18701,N_18799);
and U18924 (N_18924,N_18653,N_18724);
or U18925 (N_18925,N_18746,N_18662);
nand U18926 (N_18926,N_18672,N_18611);
nand U18927 (N_18927,N_18677,N_18689);
and U18928 (N_18928,N_18634,N_18668);
and U18929 (N_18929,N_18782,N_18702);
nand U18930 (N_18930,N_18679,N_18744);
nor U18931 (N_18931,N_18729,N_18737);
or U18932 (N_18932,N_18647,N_18728);
nor U18933 (N_18933,N_18650,N_18782);
or U18934 (N_18934,N_18648,N_18694);
or U18935 (N_18935,N_18677,N_18741);
or U18936 (N_18936,N_18745,N_18731);
or U18937 (N_18937,N_18740,N_18721);
and U18938 (N_18938,N_18748,N_18632);
nand U18939 (N_18939,N_18772,N_18783);
or U18940 (N_18940,N_18746,N_18654);
nand U18941 (N_18941,N_18739,N_18664);
nand U18942 (N_18942,N_18657,N_18790);
and U18943 (N_18943,N_18751,N_18641);
or U18944 (N_18944,N_18703,N_18728);
and U18945 (N_18945,N_18726,N_18605);
and U18946 (N_18946,N_18616,N_18701);
nor U18947 (N_18947,N_18778,N_18686);
nand U18948 (N_18948,N_18769,N_18638);
or U18949 (N_18949,N_18663,N_18666);
xnor U18950 (N_18950,N_18670,N_18737);
and U18951 (N_18951,N_18773,N_18706);
and U18952 (N_18952,N_18696,N_18618);
and U18953 (N_18953,N_18781,N_18767);
nand U18954 (N_18954,N_18615,N_18612);
or U18955 (N_18955,N_18796,N_18603);
nand U18956 (N_18956,N_18790,N_18682);
and U18957 (N_18957,N_18713,N_18727);
or U18958 (N_18958,N_18647,N_18786);
or U18959 (N_18959,N_18685,N_18610);
nand U18960 (N_18960,N_18647,N_18603);
nor U18961 (N_18961,N_18654,N_18766);
and U18962 (N_18962,N_18677,N_18732);
xnor U18963 (N_18963,N_18706,N_18682);
nor U18964 (N_18964,N_18792,N_18742);
nor U18965 (N_18965,N_18680,N_18621);
nand U18966 (N_18966,N_18640,N_18785);
nand U18967 (N_18967,N_18673,N_18707);
nor U18968 (N_18968,N_18664,N_18751);
nand U18969 (N_18969,N_18664,N_18611);
nor U18970 (N_18970,N_18681,N_18760);
or U18971 (N_18971,N_18756,N_18729);
nor U18972 (N_18972,N_18710,N_18758);
nand U18973 (N_18973,N_18606,N_18621);
or U18974 (N_18974,N_18732,N_18617);
nand U18975 (N_18975,N_18629,N_18775);
xor U18976 (N_18976,N_18720,N_18749);
or U18977 (N_18977,N_18619,N_18737);
nor U18978 (N_18978,N_18669,N_18716);
and U18979 (N_18979,N_18776,N_18605);
or U18980 (N_18980,N_18704,N_18793);
nor U18981 (N_18981,N_18607,N_18781);
nor U18982 (N_18982,N_18693,N_18623);
nor U18983 (N_18983,N_18670,N_18786);
or U18984 (N_18984,N_18791,N_18674);
nor U18985 (N_18985,N_18618,N_18772);
nand U18986 (N_18986,N_18670,N_18690);
xnor U18987 (N_18987,N_18605,N_18686);
or U18988 (N_18988,N_18764,N_18712);
and U18989 (N_18989,N_18736,N_18771);
nor U18990 (N_18990,N_18655,N_18613);
nor U18991 (N_18991,N_18607,N_18728);
or U18992 (N_18992,N_18705,N_18795);
xor U18993 (N_18993,N_18743,N_18792);
or U18994 (N_18994,N_18607,N_18628);
nor U18995 (N_18995,N_18680,N_18665);
and U18996 (N_18996,N_18652,N_18695);
and U18997 (N_18997,N_18715,N_18729);
nand U18998 (N_18998,N_18734,N_18763);
and U18999 (N_18999,N_18645,N_18613);
or U19000 (N_19000,N_18958,N_18924);
nand U19001 (N_19001,N_18995,N_18861);
nor U19002 (N_19002,N_18889,N_18965);
nand U19003 (N_19003,N_18884,N_18896);
xnor U19004 (N_19004,N_18880,N_18973);
nor U19005 (N_19005,N_18823,N_18916);
xor U19006 (N_19006,N_18801,N_18853);
and U19007 (N_19007,N_18942,N_18909);
nand U19008 (N_19008,N_18804,N_18867);
or U19009 (N_19009,N_18919,N_18922);
nor U19010 (N_19010,N_18888,N_18943);
and U19011 (N_19011,N_18964,N_18935);
nor U19012 (N_19012,N_18806,N_18951);
nor U19013 (N_19013,N_18895,N_18862);
nor U19014 (N_19014,N_18982,N_18821);
and U19015 (N_19015,N_18925,N_18944);
and U19016 (N_19016,N_18993,N_18932);
nor U19017 (N_19017,N_18915,N_18815);
xnor U19018 (N_19018,N_18968,N_18956);
nand U19019 (N_19019,N_18812,N_18937);
nand U19020 (N_19020,N_18908,N_18959);
and U19021 (N_19021,N_18855,N_18810);
nor U19022 (N_19022,N_18999,N_18988);
nand U19023 (N_19023,N_18962,N_18926);
or U19024 (N_19024,N_18848,N_18992);
and U19025 (N_19025,N_18912,N_18824);
and U19026 (N_19026,N_18840,N_18986);
and U19027 (N_19027,N_18831,N_18976);
nand U19028 (N_19028,N_18989,N_18891);
nor U19029 (N_19029,N_18886,N_18887);
nor U19030 (N_19030,N_18854,N_18826);
and U19031 (N_19031,N_18990,N_18903);
and U19032 (N_19032,N_18894,N_18825);
and U19033 (N_19033,N_18827,N_18914);
and U19034 (N_19034,N_18816,N_18910);
nand U19035 (N_19035,N_18822,N_18991);
or U19036 (N_19036,N_18869,N_18837);
or U19037 (N_19037,N_18979,N_18835);
or U19038 (N_19038,N_18817,N_18872);
nor U19039 (N_19039,N_18945,N_18953);
or U19040 (N_19040,N_18996,N_18949);
nand U19041 (N_19041,N_18875,N_18874);
xnor U19042 (N_19042,N_18923,N_18984);
nand U19043 (N_19043,N_18808,N_18948);
nand U19044 (N_19044,N_18900,N_18902);
nor U19045 (N_19045,N_18921,N_18936);
nor U19046 (N_19046,N_18966,N_18834);
nand U19047 (N_19047,N_18980,N_18829);
and U19048 (N_19048,N_18917,N_18941);
or U19049 (N_19049,N_18934,N_18885);
nand U19050 (N_19050,N_18849,N_18859);
nand U19051 (N_19051,N_18863,N_18851);
nand U19052 (N_19052,N_18929,N_18871);
nor U19053 (N_19053,N_18946,N_18905);
or U19054 (N_19054,N_18847,N_18836);
and U19055 (N_19055,N_18985,N_18950);
nand U19056 (N_19056,N_18960,N_18814);
nand U19057 (N_19057,N_18860,N_18899);
and U19058 (N_19058,N_18893,N_18839);
or U19059 (N_19059,N_18957,N_18911);
nor U19060 (N_19060,N_18832,N_18845);
or U19061 (N_19061,N_18805,N_18811);
and U19062 (N_19062,N_18846,N_18969);
nor U19063 (N_19063,N_18907,N_18938);
and U19064 (N_19064,N_18852,N_18975);
or U19065 (N_19065,N_18940,N_18920);
nand U19066 (N_19066,N_18819,N_18866);
nand U19067 (N_19067,N_18882,N_18898);
nor U19068 (N_19068,N_18865,N_18971);
nor U19069 (N_19069,N_18850,N_18987);
nor U19070 (N_19070,N_18952,N_18876);
nand U19071 (N_19071,N_18998,N_18809);
and U19072 (N_19072,N_18931,N_18833);
or U19073 (N_19073,N_18961,N_18955);
nor U19074 (N_19074,N_18890,N_18803);
and U19075 (N_19075,N_18967,N_18879);
nand U19076 (N_19076,N_18954,N_18830);
nor U19077 (N_19077,N_18906,N_18928);
and U19078 (N_19078,N_18930,N_18918);
nand U19079 (N_19079,N_18820,N_18807);
nand U19080 (N_19080,N_18870,N_18800);
nor U19081 (N_19081,N_18813,N_18970);
xor U19082 (N_19082,N_18972,N_18881);
or U19083 (N_19083,N_18818,N_18802);
nor U19084 (N_19084,N_18994,N_18939);
nand U19085 (N_19085,N_18978,N_18897);
nor U19086 (N_19086,N_18883,N_18864);
and U19087 (N_19087,N_18878,N_18873);
or U19088 (N_19088,N_18856,N_18828);
and U19089 (N_19089,N_18877,N_18858);
and U19090 (N_19090,N_18892,N_18843);
nand U19091 (N_19091,N_18868,N_18981);
nand U19092 (N_19092,N_18901,N_18841);
nand U19093 (N_19093,N_18844,N_18977);
and U19094 (N_19094,N_18838,N_18913);
and U19095 (N_19095,N_18947,N_18933);
nand U19096 (N_19096,N_18983,N_18842);
nor U19097 (N_19097,N_18857,N_18974);
nand U19098 (N_19098,N_18963,N_18904);
or U19099 (N_19099,N_18927,N_18997);
or U19100 (N_19100,N_18959,N_18950);
nand U19101 (N_19101,N_18989,N_18811);
nor U19102 (N_19102,N_18957,N_18880);
and U19103 (N_19103,N_18849,N_18993);
and U19104 (N_19104,N_18999,N_18890);
and U19105 (N_19105,N_18867,N_18824);
and U19106 (N_19106,N_18838,N_18979);
nor U19107 (N_19107,N_18973,N_18863);
and U19108 (N_19108,N_18889,N_18863);
nor U19109 (N_19109,N_18885,N_18978);
or U19110 (N_19110,N_18868,N_18856);
and U19111 (N_19111,N_18828,N_18854);
or U19112 (N_19112,N_18976,N_18933);
nand U19113 (N_19113,N_18874,N_18962);
or U19114 (N_19114,N_18944,N_18977);
nor U19115 (N_19115,N_18927,N_18800);
or U19116 (N_19116,N_18896,N_18809);
nor U19117 (N_19117,N_18840,N_18976);
and U19118 (N_19118,N_18824,N_18852);
or U19119 (N_19119,N_18855,N_18889);
nand U19120 (N_19120,N_18894,N_18925);
and U19121 (N_19121,N_18871,N_18857);
nor U19122 (N_19122,N_18864,N_18862);
and U19123 (N_19123,N_18854,N_18840);
nand U19124 (N_19124,N_18936,N_18999);
and U19125 (N_19125,N_18968,N_18929);
and U19126 (N_19126,N_18808,N_18935);
or U19127 (N_19127,N_18838,N_18934);
nand U19128 (N_19128,N_18876,N_18821);
xnor U19129 (N_19129,N_18965,N_18909);
nand U19130 (N_19130,N_18932,N_18960);
nor U19131 (N_19131,N_18972,N_18854);
and U19132 (N_19132,N_18908,N_18907);
nand U19133 (N_19133,N_18800,N_18807);
and U19134 (N_19134,N_18935,N_18834);
nor U19135 (N_19135,N_18831,N_18810);
nor U19136 (N_19136,N_18826,N_18803);
xor U19137 (N_19137,N_18867,N_18906);
nor U19138 (N_19138,N_18954,N_18851);
nor U19139 (N_19139,N_18996,N_18960);
and U19140 (N_19140,N_18817,N_18854);
or U19141 (N_19141,N_18817,N_18918);
or U19142 (N_19142,N_18998,N_18817);
nor U19143 (N_19143,N_18887,N_18843);
or U19144 (N_19144,N_18897,N_18981);
or U19145 (N_19145,N_18958,N_18994);
or U19146 (N_19146,N_18926,N_18978);
nor U19147 (N_19147,N_18860,N_18911);
nand U19148 (N_19148,N_18939,N_18847);
or U19149 (N_19149,N_18821,N_18864);
or U19150 (N_19150,N_18973,N_18821);
and U19151 (N_19151,N_18835,N_18919);
nand U19152 (N_19152,N_18950,N_18933);
and U19153 (N_19153,N_18894,N_18961);
nand U19154 (N_19154,N_18886,N_18868);
and U19155 (N_19155,N_18871,N_18829);
nand U19156 (N_19156,N_18886,N_18999);
or U19157 (N_19157,N_18913,N_18973);
or U19158 (N_19158,N_18903,N_18833);
and U19159 (N_19159,N_18923,N_18896);
nor U19160 (N_19160,N_18885,N_18810);
and U19161 (N_19161,N_18950,N_18805);
nand U19162 (N_19162,N_18824,N_18930);
nand U19163 (N_19163,N_18994,N_18977);
nor U19164 (N_19164,N_18971,N_18959);
or U19165 (N_19165,N_18860,N_18957);
or U19166 (N_19166,N_18886,N_18830);
nand U19167 (N_19167,N_18883,N_18911);
and U19168 (N_19168,N_18982,N_18957);
or U19169 (N_19169,N_18938,N_18902);
and U19170 (N_19170,N_18888,N_18815);
and U19171 (N_19171,N_18953,N_18853);
nor U19172 (N_19172,N_18814,N_18957);
nand U19173 (N_19173,N_18895,N_18850);
or U19174 (N_19174,N_18852,N_18826);
nor U19175 (N_19175,N_18943,N_18877);
nand U19176 (N_19176,N_18924,N_18957);
and U19177 (N_19177,N_18820,N_18946);
nand U19178 (N_19178,N_18875,N_18970);
nand U19179 (N_19179,N_18905,N_18920);
and U19180 (N_19180,N_18971,N_18938);
nor U19181 (N_19181,N_18896,N_18848);
nand U19182 (N_19182,N_18933,N_18841);
and U19183 (N_19183,N_18914,N_18886);
and U19184 (N_19184,N_18977,N_18878);
nor U19185 (N_19185,N_18932,N_18826);
nor U19186 (N_19186,N_18930,N_18979);
and U19187 (N_19187,N_18985,N_18885);
nor U19188 (N_19188,N_18893,N_18933);
or U19189 (N_19189,N_18951,N_18937);
and U19190 (N_19190,N_18865,N_18880);
nor U19191 (N_19191,N_18819,N_18878);
nor U19192 (N_19192,N_18863,N_18945);
and U19193 (N_19193,N_18987,N_18870);
nand U19194 (N_19194,N_18977,N_18806);
nor U19195 (N_19195,N_18845,N_18953);
nand U19196 (N_19196,N_18818,N_18853);
nor U19197 (N_19197,N_18991,N_18855);
or U19198 (N_19198,N_18852,N_18902);
and U19199 (N_19199,N_18943,N_18972);
or U19200 (N_19200,N_19083,N_19073);
or U19201 (N_19201,N_19037,N_19142);
or U19202 (N_19202,N_19040,N_19090);
or U19203 (N_19203,N_19026,N_19035);
nor U19204 (N_19204,N_19181,N_19050);
nand U19205 (N_19205,N_19059,N_19184);
nor U19206 (N_19206,N_19012,N_19192);
and U19207 (N_19207,N_19029,N_19109);
nand U19208 (N_19208,N_19137,N_19114);
nor U19209 (N_19209,N_19189,N_19097);
nor U19210 (N_19210,N_19062,N_19100);
nand U19211 (N_19211,N_19136,N_19128);
xnor U19212 (N_19212,N_19106,N_19158);
nand U19213 (N_19213,N_19197,N_19168);
and U19214 (N_19214,N_19198,N_19143);
nor U19215 (N_19215,N_19155,N_19081);
and U19216 (N_19216,N_19056,N_19044);
nand U19217 (N_19217,N_19048,N_19130);
nand U19218 (N_19218,N_19157,N_19084);
or U19219 (N_19219,N_19031,N_19135);
nor U19220 (N_19220,N_19166,N_19093);
xor U19221 (N_19221,N_19134,N_19153);
and U19222 (N_19222,N_19110,N_19161);
nand U19223 (N_19223,N_19057,N_19045);
nand U19224 (N_19224,N_19159,N_19116);
nor U19225 (N_19225,N_19022,N_19112);
xor U19226 (N_19226,N_19131,N_19160);
nor U19227 (N_19227,N_19186,N_19156);
or U19228 (N_19228,N_19065,N_19039);
or U19229 (N_19229,N_19077,N_19104);
xnor U19230 (N_19230,N_19041,N_19173);
nor U19231 (N_19231,N_19180,N_19177);
or U19232 (N_19232,N_19052,N_19194);
and U19233 (N_19233,N_19092,N_19047);
nor U19234 (N_19234,N_19170,N_19024);
nor U19235 (N_19235,N_19103,N_19095);
nor U19236 (N_19236,N_19054,N_19190);
nand U19237 (N_19237,N_19129,N_19108);
or U19238 (N_19238,N_19105,N_19094);
nor U19239 (N_19239,N_19008,N_19185);
nand U19240 (N_19240,N_19096,N_19145);
and U19241 (N_19241,N_19139,N_19033);
nand U19242 (N_19242,N_19066,N_19016);
and U19243 (N_19243,N_19119,N_19003);
nand U19244 (N_19244,N_19121,N_19150);
and U19245 (N_19245,N_19030,N_19085);
and U19246 (N_19246,N_19051,N_19027);
nor U19247 (N_19247,N_19006,N_19115);
or U19248 (N_19248,N_19034,N_19071);
nor U19249 (N_19249,N_19021,N_19068);
and U19250 (N_19250,N_19053,N_19148);
and U19251 (N_19251,N_19020,N_19078);
or U19252 (N_19252,N_19176,N_19009);
xnor U19253 (N_19253,N_19038,N_19175);
or U19254 (N_19254,N_19165,N_19069);
nor U19255 (N_19255,N_19018,N_19091);
nor U19256 (N_19256,N_19058,N_19144);
nand U19257 (N_19257,N_19087,N_19011);
nand U19258 (N_19258,N_19002,N_19042);
or U19259 (N_19259,N_19149,N_19064);
nand U19260 (N_19260,N_19147,N_19004);
nor U19261 (N_19261,N_19132,N_19079);
nor U19262 (N_19262,N_19179,N_19196);
nor U19263 (N_19263,N_19123,N_19111);
nor U19264 (N_19264,N_19086,N_19151);
nor U19265 (N_19265,N_19167,N_19099);
xor U19266 (N_19266,N_19082,N_19061);
nor U19267 (N_19267,N_19015,N_19074);
nor U19268 (N_19268,N_19023,N_19125);
and U19269 (N_19269,N_19017,N_19174);
or U19270 (N_19270,N_19001,N_19193);
nor U19271 (N_19271,N_19076,N_19140);
and U19272 (N_19272,N_19183,N_19113);
nand U19273 (N_19273,N_19182,N_19075);
or U19274 (N_19274,N_19010,N_19191);
nor U19275 (N_19275,N_19118,N_19098);
nand U19276 (N_19276,N_19032,N_19102);
xor U19277 (N_19277,N_19107,N_19163);
nor U19278 (N_19278,N_19172,N_19007);
and U19279 (N_19279,N_19138,N_19060);
nand U19280 (N_19280,N_19063,N_19000);
and U19281 (N_19281,N_19028,N_19127);
nand U19282 (N_19282,N_19164,N_19120);
nor U19283 (N_19283,N_19154,N_19014);
and U19284 (N_19284,N_19146,N_19055);
and U19285 (N_19285,N_19088,N_19133);
nand U19286 (N_19286,N_19178,N_19072);
nand U19287 (N_19287,N_19195,N_19043);
nor U19288 (N_19288,N_19122,N_19036);
or U19289 (N_19289,N_19199,N_19070);
or U19290 (N_19290,N_19117,N_19019);
and U19291 (N_19291,N_19162,N_19187);
and U19292 (N_19292,N_19171,N_19169);
nand U19293 (N_19293,N_19152,N_19188);
or U19294 (N_19294,N_19046,N_19013);
nand U19295 (N_19295,N_19005,N_19141);
and U19296 (N_19296,N_19126,N_19089);
nand U19297 (N_19297,N_19101,N_19049);
nor U19298 (N_19298,N_19067,N_19025);
or U19299 (N_19299,N_19080,N_19124);
or U19300 (N_19300,N_19009,N_19044);
nor U19301 (N_19301,N_19024,N_19184);
nor U19302 (N_19302,N_19170,N_19181);
nand U19303 (N_19303,N_19065,N_19080);
or U19304 (N_19304,N_19139,N_19188);
or U19305 (N_19305,N_19050,N_19105);
or U19306 (N_19306,N_19146,N_19141);
and U19307 (N_19307,N_19031,N_19123);
or U19308 (N_19308,N_19013,N_19020);
and U19309 (N_19309,N_19054,N_19195);
nand U19310 (N_19310,N_19175,N_19122);
and U19311 (N_19311,N_19131,N_19195);
nor U19312 (N_19312,N_19126,N_19197);
nand U19313 (N_19313,N_19074,N_19180);
and U19314 (N_19314,N_19129,N_19173);
or U19315 (N_19315,N_19070,N_19195);
nor U19316 (N_19316,N_19132,N_19023);
and U19317 (N_19317,N_19118,N_19129);
and U19318 (N_19318,N_19083,N_19026);
and U19319 (N_19319,N_19076,N_19104);
or U19320 (N_19320,N_19066,N_19099);
nor U19321 (N_19321,N_19125,N_19150);
and U19322 (N_19322,N_19183,N_19072);
nand U19323 (N_19323,N_19189,N_19039);
xnor U19324 (N_19324,N_19075,N_19149);
and U19325 (N_19325,N_19140,N_19115);
or U19326 (N_19326,N_19127,N_19077);
nor U19327 (N_19327,N_19116,N_19077);
or U19328 (N_19328,N_19053,N_19161);
nor U19329 (N_19329,N_19082,N_19098);
xnor U19330 (N_19330,N_19155,N_19089);
nor U19331 (N_19331,N_19016,N_19108);
nand U19332 (N_19332,N_19145,N_19052);
nor U19333 (N_19333,N_19145,N_19017);
nand U19334 (N_19334,N_19020,N_19025);
and U19335 (N_19335,N_19082,N_19010);
nand U19336 (N_19336,N_19146,N_19184);
and U19337 (N_19337,N_19066,N_19164);
or U19338 (N_19338,N_19041,N_19031);
or U19339 (N_19339,N_19063,N_19043);
nand U19340 (N_19340,N_19167,N_19184);
or U19341 (N_19341,N_19105,N_19003);
nand U19342 (N_19342,N_19055,N_19047);
and U19343 (N_19343,N_19037,N_19047);
nor U19344 (N_19344,N_19152,N_19079);
and U19345 (N_19345,N_19016,N_19124);
nand U19346 (N_19346,N_19092,N_19115);
nor U19347 (N_19347,N_19094,N_19039);
and U19348 (N_19348,N_19060,N_19132);
nand U19349 (N_19349,N_19040,N_19146);
or U19350 (N_19350,N_19132,N_19116);
nand U19351 (N_19351,N_19093,N_19175);
and U19352 (N_19352,N_19065,N_19082);
nor U19353 (N_19353,N_19193,N_19135);
nor U19354 (N_19354,N_19066,N_19071);
nor U19355 (N_19355,N_19007,N_19078);
or U19356 (N_19356,N_19125,N_19147);
nand U19357 (N_19357,N_19098,N_19085);
and U19358 (N_19358,N_19130,N_19163);
nor U19359 (N_19359,N_19185,N_19172);
nand U19360 (N_19360,N_19149,N_19044);
nand U19361 (N_19361,N_19185,N_19058);
or U19362 (N_19362,N_19147,N_19063);
nand U19363 (N_19363,N_19024,N_19199);
nand U19364 (N_19364,N_19113,N_19119);
nand U19365 (N_19365,N_19083,N_19031);
or U19366 (N_19366,N_19086,N_19132);
nor U19367 (N_19367,N_19176,N_19190);
nand U19368 (N_19368,N_19112,N_19090);
and U19369 (N_19369,N_19065,N_19093);
or U19370 (N_19370,N_19150,N_19113);
nor U19371 (N_19371,N_19149,N_19035);
or U19372 (N_19372,N_19168,N_19081);
nor U19373 (N_19373,N_19192,N_19153);
or U19374 (N_19374,N_19176,N_19037);
nor U19375 (N_19375,N_19026,N_19153);
or U19376 (N_19376,N_19136,N_19020);
nand U19377 (N_19377,N_19064,N_19183);
nor U19378 (N_19378,N_19085,N_19151);
and U19379 (N_19379,N_19046,N_19023);
nor U19380 (N_19380,N_19135,N_19018);
and U19381 (N_19381,N_19166,N_19196);
and U19382 (N_19382,N_19085,N_19027);
xnor U19383 (N_19383,N_19184,N_19078);
or U19384 (N_19384,N_19011,N_19175);
nor U19385 (N_19385,N_19062,N_19151);
nand U19386 (N_19386,N_19171,N_19095);
or U19387 (N_19387,N_19075,N_19143);
and U19388 (N_19388,N_19170,N_19107);
nor U19389 (N_19389,N_19141,N_19084);
or U19390 (N_19390,N_19183,N_19008);
or U19391 (N_19391,N_19094,N_19188);
and U19392 (N_19392,N_19171,N_19143);
and U19393 (N_19393,N_19114,N_19095);
and U19394 (N_19394,N_19026,N_19098);
or U19395 (N_19395,N_19130,N_19143);
and U19396 (N_19396,N_19085,N_19135);
and U19397 (N_19397,N_19150,N_19174);
nand U19398 (N_19398,N_19054,N_19035);
nand U19399 (N_19399,N_19043,N_19110);
nor U19400 (N_19400,N_19385,N_19367);
and U19401 (N_19401,N_19280,N_19334);
and U19402 (N_19402,N_19287,N_19341);
nand U19403 (N_19403,N_19298,N_19371);
and U19404 (N_19404,N_19309,N_19247);
nor U19405 (N_19405,N_19305,N_19318);
nand U19406 (N_19406,N_19275,N_19213);
and U19407 (N_19407,N_19366,N_19357);
nand U19408 (N_19408,N_19286,N_19231);
or U19409 (N_19409,N_19209,N_19325);
and U19410 (N_19410,N_19228,N_19375);
nor U19411 (N_19411,N_19246,N_19389);
or U19412 (N_19412,N_19251,N_19396);
and U19413 (N_19413,N_19290,N_19203);
nor U19414 (N_19414,N_19356,N_19360);
nand U19415 (N_19415,N_19259,N_19352);
or U19416 (N_19416,N_19380,N_19317);
nand U19417 (N_19417,N_19224,N_19250);
or U19418 (N_19418,N_19208,N_19379);
and U19419 (N_19419,N_19323,N_19358);
nand U19420 (N_19420,N_19265,N_19221);
nand U19421 (N_19421,N_19235,N_19321);
nand U19422 (N_19422,N_19350,N_19255);
nand U19423 (N_19423,N_19391,N_19292);
nand U19424 (N_19424,N_19272,N_19283);
or U19425 (N_19425,N_19273,N_19285);
and U19426 (N_19426,N_19328,N_19207);
nor U19427 (N_19427,N_19232,N_19218);
and U19428 (N_19428,N_19311,N_19374);
or U19429 (N_19429,N_19327,N_19266);
and U19430 (N_19430,N_19338,N_19288);
nand U19431 (N_19431,N_19210,N_19223);
nand U19432 (N_19432,N_19322,N_19234);
and U19433 (N_19433,N_19390,N_19348);
and U19434 (N_19434,N_19383,N_19336);
nor U19435 (N_19435,N_19227,N_19243);
or U19436 (N_19436,N_19204,N_19342);
or U19437 (N_19437,N_19282,N_19241);
nand U19438 (N_19438,N_19368,N_19351);
and U19439 (N_19439,N_19382,N_19245);
nand U19440 (N_19440,N_19284,N_19274);
or U19441 (N_19441,N_19212,N_19254);
nor U19442 (N_19442,N_19353,N_19363);
or U19443 (N_19443,N_19200,N_19315);
or U19444 (N_19444,N_19399,N_19258);
nor U19445 (N_19445,N_19222,N_19332);
nand U19446 (N_19446,N_19369,N_19316);
and U19447 (N_19447,N_19215,N_19278);
xnor U19448 (N_19448,N_19364,N_19248);
or U19449 (N_19449,N_19268,N_19202);
or U19450 (N_19450,N_19313,N_19238);
nand U19451 (N_19451,N_19307,N_19249);
nand U19452 (N_19452,N_19205,N_19392);
nand U19453 (N_19453,N_19393,N_19361);
nor U19454 (N_19454,N_19330,N_19310);
nor U19455 (N_19455,N_19340,N_19267);
or U19456 (N_19456,N_19263,N_19217);
and U19457 (N_19457,N_19201,N_19355);
nand U19458 (N_19458,N_19230,N_19312);
or U19459 (N_19459,N_19384,N_19314);
and U19460 (N_19460,N_19297,N_19291);
nand U19461 (N_19461,N_19395,N_19240);
and U19462 (N_19462,N_19387,N_19397);
and U19463 (N_19463,N_19377,N_19320);
nand U19464 (N_19464,N_19264,N_19252);
or U19465 (N_19465,N_19279,N_19372);
or U19466 (N_19466,N_19262,N_19378);
nor U19467 (N_19467,N_19304,N_19337);
and U19468 (N_19468,N_19226,N_19302);
and U19469 (N_19469,N_19236,N_19359);
nand U19470 (N_19470,N_19308,N_19333);
nand U19471 (N_19471,N_19244,N_19376);
and U19472 (N_19472,N_19370,N_19339);
or U19473 (N_19473,N_19270,N_19386);
and U19474 (N_19474,N_19261,N_19211);
nand U19475 (N_19475,N_19398,N_19242);
nand U19476 (N_19476,N_19281,N_19326);
nor U19477 (N_19477,N_19345,N_19219);
and U19478 (N_19478,N_19296,N_19239);
and U19479 (N_19479,N_19253,N_19394);
nand U19480 (N_19480,N_19344,N_19346);
nor U19481 (N_19481,N_19324,N_19329);
and U19482 (N_19482,N_19300,N_19225);
nor U19483 (N_19483,N_19256,N_19388);
and U19484 (N_19484,N_19293,N_19347);
or U19485 (N_19485,N_19303,N_19295);
nor U19486 (N_19486,N_19257,N_19260);
nor U19487 (N_19487,N_19276,N_19335);
and U19488 (N_19488,N_19354,N_19299);
nand U19489 (N_19489,N_19269,N_19216);
nor U19490 (N_19490,N_19349,N_19381);
or U19491 (N_19491,N_19331,N_19237);
nand U19492 (N_19492,N_19294,N_19319);
nand U19493 (N_19493,N_19373,N_19365);
nand U19494 (N_19494,N_19206,N_19306);
nor U19495 (N_19495,N_19362,N_19220);
or U19496 (N_19496,N_19214,N_19343);
or U19497 (N_19497,N_19289,N_19301);
nand U19498 (N_19498,N_19229,N_19277);
and U19499 (N_19499,N_19271,N_19233);
nor U19500 (N_19500,N_19396,N_19235);
or U19501 (N_19501,N_19381,N_19270);
and U19502 (N_19502,N_19378,N_19343);
nand U19503 (N_19503,N_19341,N_19226);
nor U19504 (N_19504,N_19256,N_19234);
nor U19505 (N_19505,N_19214,N_19363);
nand U19506 (N_19506,N_19305,N_19336);
and U19507 (N_19507,N_19395,N_19323);
nand U19508 (N_19508,N_19289,N_19240);
nor U19509 (N_19509,N_19284,N_19254);
nand U19510 (N_19510,N_19268,N_19208);
nand U19511 (N_19511,N_19246,N_19383);
or U19512 (N_19512,N_19222,N_19228);
or U19513 (N_19513,N_19242,N_19350);
and U19514 (N_19514,N_19386,N_19201);
and U19515 (N_19515,N_19265,N_19319);
and U19516 (N_19516,N_19378,N_19306);
nand U19517 (N_19517,N_19280,N_19295);
nand U19518 (N_19518,N_19318,N_19321);
or U19519 (N_19519,N_19349,N_19310);
nor U19520 (N_19520,N_19213,N_19361);
and U19521 (N_19521,N_19203,N_19258);
and U19522 (N_19522,N_19284,N_19309);
xnor U19523 (N_19523,N_19218,N_19319);
nand U19524 (N_19524,N_19337,N_19269);
xor U19525 (N_19525,N_19376,N_19367);
nand U19526 (N_19526,N_19268,N_19377);
nor U19527 (N_19527,N_19226,N_19219);
nor U19528 (N_19528,N_19273,N_19396);
nor U19529 (N_19529,N_19237,N_19349);
nand U19530 (N_19530,N_19220,N_19201);
or U19531 (N_19531,N_19240,N_19372);
nor U19532 (N_19532,N_19395,N_19350);
or U19533 (N_19533,N_19285,N_19238);
nand U19534 (N_19534,N_19284,N_19368);
nor U19535 (N_19535,N_19241,N_19332);
or U19536 (N_19536,N_19268,N_19393);
nand U19537 (N_19537,N_19335,N_19316);
and U19538 (N_19538,N_19264,N_19219);
nor U19539 (N_19539,N_19202,N_19321);
or U19540 (N_19540,N_19340,N_19258);
and U19541 (N_19541,N_19365,N_19285);
xor U19542 (N_19542,N_19312,N_19211);
nand U19543 (N_19543,N_19331,N_19246);
or U19544 (N_19544,N_19221,N_19272);
nor U19545 (N_19545,N_19327,N_19240);
and U19546 (N_19546,N_19229,N_19340);
nor U19547 (N_19547,N_19324,N_19220);
nand U19548 (N_19548,N_19295,N_19282);
and U19549 (N_19549,N_19294,N_19291);
and U19550 (N_19550,N_19367,N_19278);
or U19551 (N_19551,N_19223,N_19309);
nor U19552 (N_19552,N_19364,N_19318);
or U19553 (N_19553,N_19227,N_19383);
or U19554 (N_19554,N_19398,N_19369);
nor U19555 (N_19555,N_19217,N_19270);
nand U19556 (N_19556,N_19247,N_19320);
nand U19557 (N_19557,N_19316,N_19307);
nand U19558 (N_19558,N_19350,N_19292);
and U19559 (N_19559,N_19302,N_19201);
and U19560 (N_19560,N_19341,N_19360);
nand U19561 (N_19561,N_19299,N_19338);
nor U19562 (N_19562,N_19366,N_19340);
nor U19563 (N_19563,N_19361,N_19380);
nand U19564 (N_19564,N_19284,N_19395);
nand U19565 (N_19565,N_19354,N_19346);
or U19566 (N_19566,N_19385,N_19229);
or U19567 (N_19567,N_19295,N_19252);
and U19568 (N_19568,N_19296,N_19318);
or U19569 (N_19569,N_19348,N_19297);
or U19570 (N_19570,N_19381,N_19291);
nor U19571 (N_19571,N_19211,N_19351);
nand U19572 (N_19572,N_19225,N_19233);
nor U19573 (N_19573,N_19317,N_19352);
and U19574 (N_19574,N_19264,N_19335);
and U19575 (N_19575,N_19284,N_19223);
or U19576 (N_19576,N_19224,N_19302);
nand U19577 (N_19577,N_19352,N_19222);
nor U19578 (N_19578,N_19294,N_19256);
and U19579 (N_19579,N_19303,N_19209);
nor U19580 (N_19580,N_19346,N_19264);
and U19581 (N_19581,N_19235,N_19310);
nand U19582 (N_19582,N_19240,N_19225);
and U19583 (N_19583,N_19327,N_19219);
xor U19584 (N_19584,N_19265,N_19226);
nand U19585 (N_19585,N_19348,N_19304);
or U19586 (N_19586,N_19228,N_19260);
and U19587 (N_19587,N_19379,N_19255);
xnor U19588 (N_19588,N_19331,N_19299);
or U19589 (N_19589,N_19314,N_19233);
nand U19590 (N_19590,N_19314,N_19369);
and U19591 (N_19591,N_19256,N_19266);
or U19592 (N_19592,N_19342,N_19217);
nand U19593 (N_19593,N_19367,N_19201);
nand U19594 (N_19594,N_19371,N_19350);
nand U19595 (N_19595,N_19267,N_19314);
nand U19596 (N_19596,N_19285,N_19204);
nand U19597 (N_19597,N_19307,N_19383);
and U19598 (N_19598,N_19215,N_19343);
nand U19599 (N_19599,N_19224,N_19391);
and U19600 (N_19600,N_19593,N_19424);
nand U19601 (N_19601,N_19444,N_19463);
nand U19602 (N_19602,N_19540,N_19520);
nor U19603 (N_19603,N_19564,N_19488);
or U19604 (N_19604,N_19479,N_19402);
nor U19605 (N_19605,N_19582,N_19422);
nor U19606 (N_19606,N_19416,N_19465);
nand U19607 (N_19607,N_19468,N_19408);
and U19608 (N_19608,N_19525,N_19599);
and U19609 (N_19609,N_19576,N_19415);
nand U19610 (N_19610,N_19522,N_19443);
and U19611 (N_19611,N_19505,N_19403);
and U19612 (N_19612,N_19553,N_19453);
nand U19613 (N_19613,N_19501,N_19592);
or U19614 (N_19614,N_19458,N_19430);
nor U19615 (N_19615,N_19409,N_19476);
and U19616 (N_19616,N_19554,N_19542);
or U19617 (N_19617,N_19558,N_19496);
or U19618 (N_19618,N_19492,N_19438);
nor U19619 (N_19619,N_19419,N_19449);
nor U19620 (N_19620,N_19432,N_19507);
or U19621 (N_19621,N_19434,N_19551);
nand U19622 (N_19622,N_19474,N_19559);
xor U19623 (N_19623,N_19495,N_19568);
nand U19624 (N_19624,N_19555,N_19404);
xor U19625 (N_19625,N_19481,N_19497);
or U19626 (N_19626,N_19586,N_19509);
nor U19627 (N_19627,N_19452,N_19566);
or U19628 (N_19628,N_19562,N_19417);
or U19629 (N_19629,N_19462,N_19412);
and U19630 (N_19630,N_19508,N_19485);
nor U19631 (N_19631,N_19405,N_19470);
or U19632 (N_19632,N_19502,N_19513);
or U19633 (N_19633,N_19546,N_19538);
or U19634 (N_19634,N_19460,N_19528);
nor U19635 (N_19635,N_19441,N_19450);
and U19636 (N_19636,N_19596,N_19451);
nand U19637 (N_19637,N_19567,N_19503);
nand U19638 (N_19638,N_19590,N_19560);
and U19639 (N_19639,N_19445,N_19484);
or U19640 (N_19640,N_19550,N_19584);
or U19641 (N_19641,N_19521,N_19448);
and U19642 (N_19642,N_19523,N_19482);
or U19643 (N_19643,N_19585,N_19580);
or U19644 (N_19644,N_19545,N_19429);
or U19645 (N_19645,N_19464,N_19439);
xor U19646 (N_19646,N_19477,N_19428);
xor U19647 (N_19647,N_19537,N_19498);
nand U19648 (N_19648,N_19486,N_19530);
nand U19649 (N_19649,N_19515,N_19541);
and U19650 (N_19650,N_19573,N_19454);
nand U19651 (N_19651,N_19569,N_19570);
nor U19652 (N_19652,N_19561,N_19499);
nand U19653 (N_19653,N_19511,N_19597);
nor U19654 (N_19654,N_19427,N_19531);
or U19655 (N_19655,N_19556,N_19579);
or U19656 (N_19656,N_19544,N_19490);
and U19657 (N_19657,N_19472,N_19549);
nor U19658 (N_19658,N_19446,N_19480);
nor U19659 (N_19659,N_19598,N_19557);
nand U19660 (N_19660,N_19418,N_19413);
nor U19661 (N_19661,N_19519,N_19475);
nor U19662 (N_19662,N_19518,N_19407);
nand U19663 (N_19663,N_19431,N_19534);
nor U19664 (N_19664,N_19406,N_19469);
nand U19665 (N_19665,N_19466,N_19595);
and U19666 (N_19666,N_19423,N_19447);
and U19667 (N_19667,N_19527,N_19491);
or U19668 (N_19668,N_19440,N_19410);
nand U19669 (N_19669,N_19533,N_19442);
nand U19670 (N_19670,N_19548,N_19455);
or U19671 (N_19671,N_19425,N_19483);
nor U19672 (N_19672,N_19471,N_19524);
and U19673 (N_19673,N_19506,N_19411);
nand U19674 (N_19674,N_19433,N_19572);
or U19675 (N_19675,N_19588,N_19487);
or U19676 (N_19676,N_19489,N_19436);
nand U19677 (N_19677,N_19552,N_19478);
and U19678 (N_19678,N_19575,N_19421);
nor U19679 (N_19679,N_19581,N_19532);
nand U19680 (N_19680,N_19504,N_19563);
and U19681 (N_19681,N_19426,N_19543);
nand U19682 (N_19682,N_19461,N_19587);
nor U19683 (N_19683,N_19591,N_19459);
nand U19684 (N_19684,N_19583,N_19535);
and U19685 (N_19685,N_19577,N_19539);
and U19686 (N_19686,N_19414,N_19493);
nand U19687 (N_19687,N_19467,N_19516);
xnor U19688 (N_19688,N_19437,N_19574);
nand U19689 (N_19689,N_19401,N_19565);
and U19690 (N_19690,N_19589,N_19473);
and U19691 (N_19691,N_19517,N_19536);
xor U19692 (N_19692,N_19571,N_19494);
and U19693 (N_19693,N_19594,N_19510);
or U19694 (N_19694,N_19512,N_19435);
nand U19695 (N_19695,N_19514,N_19500);
and U19696 (N_19696,N_19456,N_19457);
and U19697 (N_19697,N_19547,N_19420);
and U19698 (N_19698,N_19578,N_19526);
and U19699 (N_19699,N_19529,N_19400);
nand U19700 (N_19700,N_19529,N_19444);
nor U19701 (N_19701,N_19468,N_19533);
and U19702 (N_19702,N_19543,N_19402);
or U19703 (N_19703,N_19506,N_19428);
and U19704 (N_19704,N_19576,N_19513);
nor U19705 (N_19705,N_19528,N_19438);
nand U19706 (N_19706,N_19545,N_19584);
nor U19707 (N_19707,N_19509,N_19576);
or U19708 (N_19708,N_19568,N_19497);
nor U19709 (N_19709,N_19491,N_19466);
or U19710 (N_19710,N_19514,N_19537);
nor U19711 (N_19711,N_19469,N_19461);
nor U19712 (N_19712,N_19578,N_19583);
or U19713 (N_19713,N_19566,N_19589);
nand U19714 (N_19714,N_19449,N_19525);
or U19715 (N_19715,N_19535,N_19504);
nor U19716 (N_19716,N_19530,N_19429);
nor U19717 (N_19717,N_19488,N_19465);
or U19718 (N_19718,N_19458,N_19539);
nor U19719 (N_19719,N_19427,N_19479);
nor U19720 (N_19720,N_19448,N_19404);
and U19721 (N_19721,N_19598,N_19458);
or U19722 (N_19722,N_19493,N_19543);
nor U19723 (N_19723,N_19407,N_19577);
and U19724 (N_19724,N_19484,N_19574);
and U19725 (N_19725,N_19438,N_19486);
xnor U19726 (N_19726,N_19442,N_19478);
or U19727 (N_19727,N_19481,N_19533);
or U19728 (N_19728,N_19529,N_19465);
or U19729 (N_19729,N_19543,N_19512);
or U19730 (N_19730,N_19566,N_19427);
nor U19731 (N_19731,N_19503,N_19590);
nand U19732 (N_19732,N_19592,N_19454);
nand U19733 (N_19733,N_19557,N_19447);
or U19734 (N_19734,N_19438,N_19515);
and U19735 (N_19735,N_19427,N_19543);
and U19736 (N_19736,N_19542,N_19541);
nor U19737 (N_19737,N_19410,N_19482);
and U19738 (N_19738,N_19421,N_19490);
and U19739 (N_19739,N_19596,N_19506);
nor U19740 (N_19740,N_19417,N_19415);
nand U19741 (N_19741,N_19511,N_19562);
and U19742 (N_19742,N_19565,N_19438);
and U19743 (N_19743,N_19511,N_19580);
and U19744 (N_19744,N_19597,N_19425);
nor U19745 (N_19745,N_19511,N_19411);
and U19746 (N_19746,N_19457,N_19563);
nor U19747 (N_19747,N_19511,N_19548);
nand U19748 (N_19748,N_19535,N_19534);
or U19749 (N_19749,N_19577,N_19519);
nor U19750 (N_19750,N_19495,N_19572);
and U19751 (N_19751,N_19431,N_19517);
nand U19752 (N_19752,N_19530,N_19450);
and U19753 (N_19753,N_19556,N_19451);
nor U19754 (N_19754,N_19452,N_19521);
nand U19755 (N_19755,N_19510,N_19595);
and U19756 (N_19756,N_19427,N_19474);
nor U19757 (N_19757,N_19569,N_19517);
or U19758 (N_19758,N_19422,N_19581);
nor U19759 (N_19759,N_19500,N_19405);
or U19760 (N_19760,N_19449,N_19427);
and U19761 (N_19761,N_19449,N_19413);
nand U19762 (N_19762,N_19544,N_19570);
xor U19763 (N_19763,N_19457,N_19573);
xnor U19764 (N_19764,N_19517,N_19560);
nand U19765 (N_19765,N_19552,N_19550);
or U19766 (N_19766,N_19487,N_19477);
and U19767 (N_19767,N_19578,N_19528);
nor U19768 (N_19768,N_19489,N_19447);
nor U19769 (N_19769,N_19538,N_19494);
nor U19770 (N_19770,N_19543,N_19595);
and U19771 (N_19771,N_19587,N_19422);
or U19772 (N_19772,N_19515,N_19549);
nand U19773 (N_19773,N_19485,N_19592);
nand U19774 (N_19774,N_19588,N_19547);
or U19775 (N_19775,N_19557,N_19527);
or U19776 (N_19776,N_19483,N_19486);
nor U19777 (N_19777,N_19564,N_19587);
or U19778 (N_19778,N_19519,N_19565);
nand U19779 (N_19779,N_19566,N_19525);
and U19780 (N_19780,N_19478,N_19594);
nand U19781 (N_19781,N_19442,N_19418);
nor U19782 (N_19782,N_19536,N_19430);
nor U19783 (N_19783,N_19440,N_19420);
and U19784 (N_19784,N_19423,N_19471);
nand U19785 (N_19785,N_19420,N_19452);
nor U19786 (N_19786,N_19493,N_19575);
nand U19787 (N_19787,N_19587,N_19598);
nor U19788 (N_19788,N_19453,N_19455);
or U19789 (N_19789,N_19409,N_19401);
and U19790 (N_19790,N_19590,N_19491);
xnor U19791 (N_19791,N_19485,N_19568);
nand U19792 (N_19792,N_19500,N_19560);
and U19793 (N_19793,N_19533,N_19464);
nor U19794 (N_19794,N_19434,N_19489);
nand U19795 (N_19795,N_19511,N_19528);
and U19796 (N_19796,N_19524,N_19545);
and U19797 (N_19797,N_19489,N_19598);
and U19798 (N_19798,N_19507,N_19504);
nand U19799 (N_19799,N_19400,N_19569);
or U19800 (N_19800,N_19676,N_19619);
nor U19801 (N_19801,N_19639,N_19702);
or U19802 (N_19802,N_19799,N_19612);
or U19803 (N_19803,N_19762,N_19746);
and U19804 (N_19804,N_19673,N_19649);
nor U19805 (N_19805,N_19665,N_19616);
nor U19806 (N_19806,N_19765,N_19758);
and U19807 (N_19807,N_19720,N_19716);
nand U19808 (N_19808,N_19696,N_19737);
or U19809 (N_19809,N_19733,N_19662);
or U19810 (N_19810,N_19734,N_19729);
nand U19811 (N_19811,N_19728,N_19667);
xnor U19812 (N_19812,N_19796,N_19689);
nand U19813 (N_19813,N_19644,N_19645);
nand U19814 (N_19814,N_19648,N_19745);
or U19815 (N_19815,N_19694,N_19610);
nor U19816 (N_19816,N_19744,N_19757);
nor U19817 (N_19817,N_19790,N_19766);
or U19818 (N_19818,N_19678,N_19764);
or U19819 (N_19819,N_19719,N_19769);
nor U19820 (N_19820,N_19726,N_19710);
nand U19821 (N_19821,N_19727,N_19660);
nor U19822 (N_19822,N_19767,N_19779);
nor U19823 (N_19823,N_19731,N_19672);
or U19824 (N_19824,N_19629,N_19627);
and U19825 (N_19825,N_19623,N_19699);
and U19826 (N_19826,N_19709,N_19756);
nand U19827 (N_19827,N_19742,N_19603);
nand U19828 (N_19828,N_19680,N_19791);
or U19829 (N_19829,N_19780,N_19788);
nand U19830 (N_19830,N_19703,N_19671);
nand U19831 (N_19831,N_19620,N_19732);
or U19832 (N_19832,N_19670,N_19604);
or U19833 (N_19833,N_19622,N_19773);
or U19834 (N_19834,N_19631,N_19721);
or U19835 (N_19835,N_19606,N_19641);
nor U19836 (N_19836,N_19736,N_19609);
nor U19837 (N_19837,N_19615,N_19657);
or U19838 (N_19838,N_19661,N_19752);
or U19839 (N_19839,N_19724,N_19748);
or U19840 (N_19840,N_19717,N_19647);
and U19841 (N_19841,N_19776,N_19789);
xnor U19842 (N_19842,N_19640,N_19698);
and U19843 (N_19843,N_19636,N_19621);
or U19844 (N_19844,N_19792,N_19674);
and U19845 (N_19845,N_19772,N_19785);
and U19846 (N_19846,N_19634,N_19675);
nor U19847 (N_19847,N_19658,N_19784);
or U19848 (N_19848,N_19701,N_19797);
nand U19849 (N_19849,N_19700,N_19656);
nor U19850 (N_19850,N_19695,N_19653);
nor U19851 (N_19851,N_19786,N_19730);
nand U19852 (N_19852,N_19740,N_19778);
or U19853 (N_19853,N_19685,N_19668);
or U19854 (N_19854,N_19614,N_19704);
nor U19855 (N_19855,N_19654,N_19669);
and U19856 (N_19856,N_19691,N_19611);
nand U19857 (N_19857,N_19659,N_19795);
and U19858 (N_19858,N_19687,N_19782);
nand U19859 (N_19859,N_19715,N_19625);
nor U19860 (N_19860,N_19725,N_19750);
and U19861 (N_19861,N_19753,N_19664);
or U19862 (N_19862,N_19690,N_19793);
nand U19863 (N_19863,N_19718,N_19618);
xnor U19864 (N_19864,N_19650,N_19638);
nor U19865 (N_19865,N_19711,N_19768);
nand U19866 (N_19866,N_19770,N_19602);
nor U19867 (N_19867,N_19713,N_19743);
nand U19868 (N_19868,N_19688,N_19794);
and U19869 (N_19869,N_19747,N_19738);
and U19870 (N_19870,N_19759,N_19751);
or U19871 (N_19871,N_19628,N_19775);
nor U19872 (N_19872,N_19643,N_19705);
nor U19873 (N_19873,N_19749,N_19755);
and U19874 (N_19874,N_19706,N_19771);
nor U19875 (N_19875,N_19708,N_19760);
or U19876 (N_19876,N_19783,N_19684);
xor U19877 (N_19877,N_19651,N_19714);
nor U19878 (N_19878,N_19787,N_19723);
nand U19879 (N_19879,N_19652,N_19735);
nor U19880 (N_19880,N_19693,N_19712);
or U19881 (N_19881,N_19781,N_19777);
nor U19882 (N_19882,N_19798,N_19697);
and U19883 (N_19883,N_19679,N_19707);
nand U19884 (N_19884,N_19605,N_19635);
and U19885 (N_19885,N_19663,N_19774);
nand U19886 (N_19886,N_19607,N_19601);
nand U19887 (N_19887,N_19763,N_19692);
nand U19888 (N_19888,N_19633,N_19686);
or U19889 (N_19889,N_19613,N_19642);
or U19890 (N_19890,N_19677,N_19754);
xnor U19891 (N_19891,N_19761,N_19646);
xor U19892 (N_19892,N_19630,N_19600);
nor U19893 (N_19893,N_19666,N_19741);
nor U19894 (N_19894,N_19681,N_19722);
nor U19895 (N_19895,N_19617,N_19608);
or U19896 (N_19896,N_19655,N_19626);
nand U19897 (N_19897,N_19637,N_19682);
nand U19898 (N_19898,N_19632,N_19624);
nand U19899 (N_19899,N_19683,N_19739);
nand U19900 (N_19900,N_19720,N_19706);
nand U19901 (N_19901,N_19643,N_19771);
nor U19902 (N_19902,N_19633,N_19780);
and U19903 (N_19903,N_19608,N_19634);
nand U19904 (N_19904,N_19680,N_19723);
nand U19905 (N_19905,N_19789,N_19763);
nand U19906 (N_19906,N_19612,N_19634);
or U19907 (N_19907,N_19777,N_19651);
nor U19908 (N_19908,N_19666,N_19783);
or U19909 (N_19909,N_19638,N_19770);
nor U19910 (N_19910,N_19736,N_19744);
or U19911 (N_19911,N_19703,N_19794);
and U19912 (N_19912,N_19652,N_19794);
nor U19913 (N_19913,N_19653,N_19678);
nand U19914 (N_19914,N_19705,N_19640);
and U19915 (N_19915,N_19613,N_19640);
and U19916 (N_19916,N_19629,N_19742);
nor U19917 (N_19917,N_19717,N_19678);
nand U19918 (N_19918,N_19681,N_19612);
nand U19919 (N_19919,N_19607,N_19783);
nand U19920 (N_19920,N_19693,N_19675);
nor U19921 (N_19921,N_19641,N_19722);
nor U19922 (N_19922,N_19715,N_19729);
or U19923 (N_19923,N_19708,N_19716);
or U19924 (N_19924,N_19705,N_19619);
and U19925 (N_19925,N_19788,N_19643);
and U19926 (N_19926,N_19658,N_19630);
nand U19927 (N_19927,N_19620,N_19654);
nand U19928 (N_19928,N_19797,N_19656);
and U19929 (N_19929,N_19636,N_19777);
nand U19930 (N_19930,N_19761,N_19740);
nand U19931 (N_19931,N_19624,N_19605);
nand U19932 (N_19932,N_19600,N_19627);
or U19933 (N_19933,N_19768,N_19787);
and U19934 (N_19934,N_19717,N_19736);
xnor U19935 (N_19935,N_19723,N_19746);
or U19936 (N_19936,N_19732,N_19632);
nand U19937 (N_19937,N_19750,N_19792);
nor U19938 (N_19938,N_19619,N_19711);
nand U19939 (N_19939,N_19606,N_19662);
and U19940 (N_19940,N_19667,N_19638);
or U19941 (N_19941,N_19631,N_19786);
nand U19942 (N_19942,N_19645,N_19786);
nand U19943 (N_19943,N_19705,N_19750);
and U19944 (N_19944,N_19689,N_19758);
nor U19945 (N_19945,N_19630,N_19700);
or U19946 (N_19946,N_19610,N_19671);
nand U19947 (N_19947,N_19737,N_19739);
nor U19948 (N_19948,N_19750,N_19648);
and U19949 (N_19949,N_19771,N_19723);
and U19950 (N_19950,N_19643,N_19627);
and U19951 (N_19951,N_19775,N_19785);
and U19952 (N_19952,N_19629,N_19652);
nand U19953 (N_19953,N_19651,N_19784);
or U19954 (N_19954,N_19716,N_19673);
and U19955 (N_19955,N_19665,N_19662);
nand U19956 (N_19956,N_19644,N_19737);
nor U19957 (N_19957,N_19764,N_19656);
and U19958 (N_19958,N_19729,N_19702);
and U19959 (N_19959,N_19724,N_19703);
nand U19960 (N_19960,N_19696,N_19699);
nand U19961 (N_19961,N_19665,N_19768);
nor U19962 (N_19962,N_19789,N_19703);
nand U19963 (N_19963,N_19788,N_19735);
or U19964 (N_19964,N_19791,N_19721);
nor U19965 (N_19965,N_19605,N_19653);
nor U19966 (N_19966,N_19738,N_19705);
and U19967 (N_19967,N_19676,N_19613);
or U19968 (N_19968,N_19620,N_19677);
nand U19969 (N_19969,N_19656,N_19698);
and U19970 (N_19970,N_19623,N_19604);
and U19971 (N_19971,N_19631,N_19683);
nand U19972 (N_19972,N_19638,N_19654);
and U19973 (N_19973,N_19794,N_19668);
and U19974 (N_19974,N_19728,N_19691);
and U19975 (N_19975,N_19792,N_19627);
and U19976 (N_19976,N_19791,N_19765);
nand U19977 (N_19977,N_19710,N_19758);
or U19978 (N_19978,N_19711,N_19616);
nand U19979 (N_19979,N_19779,N_19626);
and U19980 (N_19980,N_19658,N_19715);
and U19981 (N_19981,N_19709,N_19703);
nor U19982 (N_19982,N_19755,N_19657);
and U19983 (N_19983,N_19672,N_19761);
nor U19984 (N_19984,N_19665,N_19779);
nand U19985 (N_19985,N_19678,N_19706);
nand U19986 (N_19986,N_19756,N_19761);
or U19987 (N_19987,N_19662,N_19684);
and U19988 (N_19988,N_19772,N_19768);
and U19989 (N_19989,N_19657,N_19782);
or U19990 (N_19990,N_19641,N_19651);
nor U19991 (N_19991,N_19798,N_19745);
nor U19992 (N_19992,N_19680,N_19761);
nor U19993 (N_19993,N_19719,N_19695);
or U19994 (N_19994,N_19616,N_19765);
or U19995 (N_19995,N_19667,N_19602);
nand U19996 (N_19996,N_19626,N_19747);
nor U19997 (N_19997,N_19784,N_19665);
and U19998 (N_19998,N_19711,N_19794);
and U19999 (N_19999,N_19619,N_19791);
or UO_0 (O_0,N_19839,N_19890);
nor UO_1 (O_1,N_19879,N_19860);
nor UO_2 (O_2,N_19816,N_19831);
and UO_3 (O_3,N_19921,N_19974);
nand UO_4 (O_4,N_19836,N_19950);
and UO_5 (O_5,N_19861,N_19869);
and UO_6 (O_6,N_19865,N_19851);
nand UO_7 (O_7,N_19981,N_19937);
nor UO_8 (O_8,N_19903,N_19990);
and UO_9 (O_9,N_19947,N_19847);
nand UO_10 (O_10,N_19813,N_19966);
and UO_11 (O_11,N_19892,N_19992);
and UO_12 (O_12,N_19832,N_19987);
nor UO_13 (O_13,N_19993,N_19877);
nand UO_14 (O_14,N_19945,N_19959);
or UO_15 (O_15,N_19965,N_19932);
or UO_16 (O_16,N_19940,N_19918);
or UO_17 (O_17,N_19963,N_19872);
nor UO_18 (O_18,N_19837,N_19975);
and UO_19 (O_19,N_19922,N_19803);
nand UO_20 (O_20,N_19835,N_19896);
or UO_21 (O_21,N_19870,N_19926);
and UO_22 (O_22,N_19878,N_19935);
nor UO_23 (O_23,N_19994,N_19884);
nand UO_24 (O_24,N_19905,N_19828);
nor UO_25 (O_25,N_19876,N_19806);
and UO_26 (O_26,N_19881,N_19868);
and UO_27 (O_27,N_19980,N_19908);
nand UO_28 (O_28,N_19951,N_19907);
or UO_29 (O_29,N_19938,N_19886);
nor UO_30 (O_30,N_19991,N_19999);
and UO_31 (O_31,N_19997,N_19834);
nor UO_32 (O_32,N_19953,N_19961);
and UO_33 (O_33,N_19995,N_19809);
and UO_34 (O_34,N_19943,N_19856);
nand UO_35 (O_35,N_19821,N_19852);
nand UO_36 (O_36,N_19955,N_19913);
nor UO_37 (O_37,N_19925,N_19920);
nand UO_38 (O_38,N_19917,N_19928);
or UO_39 (O_39,N_19996,N_19958);
nor UO_40 (O_40,N_19988,N_19888);
or UO_41 (O_41,N_19874,N_19824);
nor UO_42 (O_42,N_19814,N_19811);
and UO_43 (O_43,N_19973,N_19957);
nand UO_44 (O_44,N_19822,N_19897);
nand UO_45 (O_45,N_19989,N_19929);
or UO_46 (O_46,N_19887,N_19889);
nand UO_47 (O_47,N_19915,N_19818);
and UO_48 (O_48,N_19894,N_19810);
and UO_49 (O_49,N_19805,N_19864);
or UO_50 (O_50,N_19904,N_19812);
and UO_51 (O_51,N_19895,N_19983);
and UO_52 (O_52,N_19825,N_19801);
nand UO_53 (O_53,N_19956,N_19998);
or UO_54 (O_54,N_19934,N_19944);
nor UO_55 (O_55,N_19848,N_19978);
or UO_56 (O_56,N_19863,N_19970);
nor UO_57 (O_57,N_19853,N_19979);
and UO_58 (O_58,N_19906,N_19817);
xnor UO_59 (O_59,N_19902,N_19880);
xor UO_60 (O_60,N_19962,N_19873);
or UO_61 (O_61,N_19866,N_19960);
nand UO_62 (O_62,N_19910,N_19844);
nand UO_63 (O_63,N_19909,N_19986);
and UO_64 (O_64,N_19854,N_19883);
nand UO_65 (O_65,N_19846,N_19941);
or UO_66 (O_66,N_19964,N_19972);
nor UO_67 (O_67,N_19899,N_19912);
and UO_68 (O_68,N_19841,N_19867);
or UO_69 (O_69,N_19850,N_19984);
and UO_70 (O_70,N_19919,N_19804);
or UO_71 (O_71,N_19842,N_19942);
nor UO_72 (O_72,N_19858,N_19936);
and UO_73 (O_73,N_19862,N_19807);
or UO_74 (O_74,N_19923,N_19914);
or UO_75 (O_75,N_19948,N_19815);
and UO_76 (O_76,N_19969,N_19833);
and UO_77 (O_77,N_19949,N_19827);
nand UO_78 (O_78,N_19802,N_19819);
nand UO_79 (O_79,N_19893,N_19800);
nand UO_80 (O_80,N_19857,N_19985);
and UO_81 (O_81,N_19900,N_19911);
xnor UO_82 (O_82,N_19820,N_19967);
nor UO_83 (O_83,N_19954,N_19885);
or UO_84 (O_84,N_19931,N_19891);
or UO_85 (O_85,N_19977,N_19939);
nand UO_86 (O_86,N_19849,N_19840);
or UO_87 (O_87,N_19830,N_19930);
nand UO_88 (O_88,N_19823,N_19875);
nand UO_89 (O_89,N_19946,N_19882);
and UO_90 (O_90,N_19808,N_19924);
nand UO_91 (O_91,N_19843,N_19901);
nand UO_92 (O_92,N_19898,N_19982);
or UO_93 (O_93,N_19855,N_19838);
or UO_94 (O_94,N_19871,N_19927);
and UO_95 (O_95,N_19916,N_19826);
and UO_96 (O_96,N_19968,N_19845);
and UO_97 (O_97,N_19933,N_19859);
nor UO_98 (O_98,N_19971,N_19976);
and UO_99 (O_99,N_19952,N_19829);
xnor UO_100 (O_100,N_19970,N_19813);
or UO_101 (O_101,N_19912,N_19827);
and UO_102 (O_102,N_19827,N_19972);
and UO_103 (O_103,N_19896,N_19861);
nand UO_104 (O_104,N_19821,N_19882);
and UO_105 (O_105,N_19905,N_19807);
or UO_106 (O_106,N_19844,N_19958);
nand UO_107 (O_107,N_19882,N_19909);
or UO_108 (O_108,N_19876,N_19891);
nand UO_109 (O_109,N_19829,N_19938);
nor UO_110 (O_110,N_19914,N_19958);
and UO_111 (O_111,N_19857,N_19962);
nand UO_112 (O_112,N_19803,N_19992);
nor UO_113 (O_113,N_19811,N_19881);
and UO_114 (O_114,N_19858,N_19829);
nand UO_115 (O_115,N_19808,N_19801);
nor UO_116 (O_116,N_19839,N_19938);
nor UO_117 (O_117,N_19846,N_19988);
nand UO_118 (O_118,N_19930,N_19980);
and UO_119 (O_119,N_19834,N_19866);
and UO_120 (O_120,N_19972,N_19968);
nand UO_121 (O_121,N_19979,N_19973);
nor UO_122 (O_122,N_19814,N_19806);
nor UO_123 (O_123,N_19925,N_19913);
or UO_124 (O_124,N_19950,N_19984);
nor UO_125 (O_125,N_19857,N_19945);
or UO_126 (O_126,N_19861,N_19882);
nand UO_127 (O_127,N_19911,N_19876);
or UO_128 (O_128,N_19969,N_19846);
nor UO_129 (O_129,N_19855,N_19861);
nand UO_130 (O_130,N_19948,N_19869);
and UO_131 (O_131,N_19919,N_19918);
nor UO_132 (O_132,N_19912,N_19888);
nor UO_133 (O_133,N_19873,N_19844);
nand UO_134 (O_134,N_19873,N_19924);
and UO_135 (O_135,N_19899,N_19840);
nor UO_136 (O_136,N_19993,N_19805);
nor UO_137 (O_137,N_19804,N_19879);
or UO_138 (O_138,N_19950,N_19919);
nand UO_139 (O_139,N_19895,N_19981);
and UO_140 (O_140,N_19926,N_19910);
nand UO_141 (O_141,N_19892,N_19958);
and UO_142 (O_142,N_19948,N_19831);
nor UO_143 (O_143,N_19828,N_19884);
or UO_144 (O_144,N_19857,N_19923);
nor UO_145 (O_145,N_19895,N_19867);
nand UO_146 (O_146,N_19912,N_19853);
and UO_147 (O_147,N_19960,N_19968);
and UO_148 (O_148,N_19945,N_19845);
and UO_149 (O_149,N_19892,N_19840);
or UO_150 (O_150,N_19934,N_19812);
nor UO_151 (O_151,N_19957,N_19910);
nor UO_152 (O_152,N_19890,N_19947);
or UO_153 (O_153,N_19811,N_19946);
nor UO_154 (O_154,N_19926,N_19981);
nand UO_155 (O_155,N_19822,N_19862);
and UO_156 (O_156,N_19814,N_19920);
nand UO_157 (O_157,N_19923,N_19882);
nand UO_158 (O_158,N_19924,N_19989);
nor UO_159 (O_159,N_19860,N_19894);
nand UO_160 (O_160,N_19807,N_19933);
or UO_161 (O_161,N_19888,N_19881);
or UO_162 (O_162,N_19839,N_19907);
or UO_163 (O_163,N_19980,N_19801);
nand UO_164 (O_164,N_19998,N_19892);
and UO_165 (O_165,N_19976,N_19915);
or UO_166 (O_166,N_19905,N_19943);
or UO_167 (O_167,N_19913,N_19830);
nand UO_168 (O_168,N_19924,N_19812);
nor UO_169 (O_169,N_19850,N_19950);
nand UO_170 (O_170,N_19857,N_19963);
or UO_171 (O_171,N_19953,N_19823);
and UO_172 (O_172,N_19954,N_19941);
or UO_173 (O_173,N_19932,N_19859);
nand UO_174 (O_174,N_19972,N_19990);
nand UO_175 (O_175,N_19944,N_19922);
or UO_176 (O_176,N_19805,N_19833);
and UO_177 (O_177,N_19927,N_19937);
nor UO_178 (O_178,N_19983,N_19980);
or UO_179 (O_179,N_19835,N_19984);
nand UO_180 (O_180,N_19807,N_19989);
and UO_181 (O_181,N_19958,N_19926);
xnor UO_182 (O_182,N_19937,N_19819);
nor UO_183 (O_183,N_19861,N_19827);
nand UO_184 (O_184,N_19913,N_19868);
or UO_185 (O_185,N_19861,N_19858);
or UO_186 (O_186,N_19861,N_19965);
xnor UO_187 (O_187,N_19841,N_19832);
xor UO_188 (O_188,N_19942,N_19887);
nor UO_189 (O_189,N_19941,N_19944);
and UO_190 (O_190,N_19910,N_19958);
and UO_191 (O_191,N_19834,N_19972);
nor UO_192 (O_192,N_19972,N_19881);
nor UO_193 (O_193,N_19920,N_19973);
or UO_194 (O_194,N_19881,N_19822);
or UO_195 (O_195,N_19890,N_19855);
nand UO_196 (O_196,N_19841,N_19910);
nor UO_197 (O_197,N_19848,N_19961);
or UO_198 (O_198,N_19860,N_19842);
or UO_199 (O_199,N_19818,N_19882);
and UO_200 (O_200,N_19904,N_19898);
nor UO_201 (O_201,N_19989,N_19803);
nand UO_202 (O_202,N_19881,N_19876);
and UO_203 (O_203,N_19868,N_19822);
or UO_204 (O_204,N_19801,N_19892);
nor UO_205 (O_205,N_19826,N_19895);
nor UO_206 (O_206,N_19842,N_19932);
and UO_207 (O_207,N_19953,N_19997);
nand UO_208 (O_208,N_19824,N_19834);
or UO_209 (O_209,N_19912,N_19907);
and UO_210 (O_210,N_19820,N_19803);
or UO_211 (O_211,N_19971,N_19818);
or UO_212 (O_212,N_19898,N_19842);
nor UO_213 (O_213,N_19828,N_19988);
or UO_214 (O_214,N_19893,N_19975);
nor UO_215 (O_215,N_19827,N_19900);
nand UO_216 (O_216,N_19900,N_19940);
and UO_217 (O_217,N_19837,N_19938);
nor UO_218 (O_218,N_19800,N_19905);
and UO_219 (O_219,N_19869,N_19898);
nand UO_220 (O_220,N_19843,N_19923);
or UO_221 (O_221,N_19967,N_19868);
or UO_222 (O_222,N_19932,N_19924);
nand UO_223 (O_223,N_19983,N_19869);
or UO_224 (O_224,N_19949,N_19817);
and UO_225 (O_225,N_19891,N_19947);
nor UO_226 (O_226,N_19926,N_19851);
and UO_227 (O_227,N_19940,N_19800);
nor UO_228 (O_228,N_19886,N_19952);
nor UO_229 (O_229,N_19989,N_19854);
nand UO_230 (O_230,N_19886,N_19936);
xor UO_231 (O_231,N_19880,N_19921);
nor UO_232 (O_232,N_19932,N_19951);
nor UO_233 (O_233,N_19807,N_19838);
nand UO_234 (O_234,N_19892,N_19857);
nor UO_235 (O_235,N_19943,N_19901);
and UO_236 (O_236,N_19826,N_19877);
nand UO_237 (O_237,N_19832,N_19961);
and UO_238 (O_238,N_19862,N_19813);
or UO_239 (O_239,N_19972,N_19988);
nor UO_240 (O_240,N_19860,N_19944);
nand UO_241 (O_241,N_19850,N_19925);
nand UO_242 (O_242,N_19992,N_19801);
nor UO_243 (O_243,N_19922,N_19924);
or UO_244 (O_244,N_19906,N_19992);
nor UO_245 (O_245,N_19910,N_19882);
nor UO_246 (O_246,N_19939,N_19971);
or UO_247 (O_247,N_19835,N_19824);
or UO_248 (O_248,N_19888,N_19832);
and UO_249 (O_249,N_19835,N_19924);
and UO_250 (O_250,N_19928,N_19849);
and UO_251 (O_251,N_19978,N_19865);
or UO_252 (O_252,N_19895,N_19929);
and UO_253 (O_253,N_19885,N_19828);
nor UO_254 (O_254,N_19908,N_19911);
or UO_255 (O_255,N_19922,N_19853);
and UO_256 (O_256,N_19813,N_19836);
or UO_257 (O_257,N_19949,N_19979);
and UO_258 (O_258,N_19991,N_19825);
or UO_259 (O_259,N_19880,N_19812);
nand UO_260 (O_260,N_19830,N_19890);
or UO_261 (O_261,N_19834,N_19996);
or UO_262 (O_262,N_19897,N_19908);
nor UO_263 (O_263,N_19857,N_19910);
or UO_264 (O_264,N_19995,N_19940);
nand UO_265 (O_265,N_19913,N_19943);
or UO_266 (O_266,N_19826,N_19814);
nor UO_267 (O_267,N_19929,N_19834);
and UO_268 (O_268,N_19811,N_19822);
and UO_269 (O_269,N_19973,N_19845);
nor UO_270 (O_270,N_19994,N_19807);
or UO_271 (O_271,N_19846,N_19946);
nor UO_272 (O_272,N_19953,N_19981);
and UO_273 (O_273,N_19931,N_19986);
or UO_274 (O_274,N_19943,N_19823);
and UO_275 (O_275,N_19854,N_19937);
or UO_276 (O_276,N_19882,N_19969);
and UO_277 (O_277,N_19942,N_19980);
and UO_278 (O_278,N_19965,N_19927);
or UO_279 (O_279,N_19889,N_19933);
and UO_280 (O_280,N_19898,N_19935);
nor UO_281 (O_281,N_19820,N_19914);
and UO_282 (O_282,N_19851,N_19928);
and UO_283 (O_283,N_19986,N_19838);
and UO_284 (O_284,N_19811,N_19830);
or UO_285 (O_285,N_19897,N_19937);
nand UO_286 (O_286,N_19800,N_19944);
nor UO_287 (O_287,N_19890,N_19926);
nor UO_288 (O_288,N_19866,N_19835);
and UO_289 (O_289,N_19904,N_19808);
nor UO_290 (O_290,N_19951,N_19917);
nand UO_291 (O_291,N_19956,N_19948);
nand UO_292 (O_292,N_19930,N_19801);
nand UO_293 (O_293,N_19901,N_19929);
nand UO_294 (O_294,N_19884,N_19890);
and UO_295 (O_295,N_19908,N_19984);
nand UO_296 (O_296,N_19961,N_19997);
and UO_297 (O_297,N_19970,N_19839);
and UO_298 (O_298,N_19905,N_19863);
or UO_299 (O_299,N_19961,N_19965);
or UO_300 (O_300,N_19844,N_19961);
or UO_301 (O_301,N_19949,N_19807);
and UO_302 (O_302,N_19972,N_19874);
and UO_303 (O_303,N_19970,N_19915);
nor UO_304 (O_304,N_19854,N_19982);
nor UO_305 (O_305,N_19948,N_19811);
or UO_306 (O_306,N_19931,N_19935);
or UO_307 (O_307,N_19965,N_19841);
and UO_308 (O_308,N_19882,N_19952);
or UO_309 (O_309,N_19811,N_19951);
and UO_310 (O_310,N_19868,N_19836);
nor UO_311 (O_311,N_19823,N_19843);
and UO_312 (O_312,N_19948,N_19918);
nor UO_313 (O_313,N_19880,N_19865);
nand UO_314 (O_314,N_19982,N_19865);
xor UO_315 (O_315,N_19904,N_19845);
nor UO_316 (O_316,N_19957,N_19995);
nor UO_317 (O_317,N_19847,N_19842);
nor UO_318 (O_318,N_19947,N_19910);
or UO_319 (O_319,N_19937,N_19866);
and UO_320 (O_320,N_19824,N_19986);
nor UO_321 (O_321,N_19950,N_19947);
nor UO_322 (O_322,N_19930,N_19958);
or UO_323 (O_323,N_19852,N_19941);
and UO_324 (O_324,N_19872,N_19940);
and UO_325 (O_325,N_19866,N_19901);
or UO_326 (O_326,N_19984,N_19828);
nand UO_327 (O_327,N_19929,N_19988);
and UO_328 (O_328,N_19916,N_19935);
nor UO_329 (O_329,N_19905,N_19802);
or UO_330 (O_330,N_19870,N_19911);
nor UO_331 (O_331,N_19848,N_19861);
nor UO_332 (O_332,N_19872,N_19830);
or UO_333 (O_333,N_19810,N_19934);
nor UO_334 (O_334,N_19943,N_19909);
and UO_335 (O_335,N_19867,N_19941);
nand UO_336 (O_336,N_19932,N_19837);
and UO_337 (O_337,N_19913,N_19926);
and UO_338 (O_338,N_19863,N_19910);
nor UO_339 (O_339,N_19813,N_19997);
nand UO_340 (O_340,N_19810,N_19951);
or UO_341 (O_341,N_19910,N_19824);
and UO_342 (O_342,N_19856,N_19951);
and UO_343 (O_343,N_19859,N_19922);
nor UO_344 (O_344,N_19952,N_19915);
and UO_345 (O_345,N_19825,N_19855);
nand UO_346 (O_346,N_19954,N_19857);
or UO_347 (O_347,N_19876,N_19963);
nand UO_348 (O_348,N_19903,N_19820);
or UO_349 (O_349,N_19800,N_19840);
nand UO_350 (O_350,N_19982,N_19843);
or UO_351 (O_351,N_19912,N_19974);
or UO_352 (O_352,N_19966,N_19904);
nand UO_353 (O_353,N_19992,N_19995);
and UO_354 (O_354,N_19959,N_19860);
nor UO_355 (O_355,N_19910,N_19832);
and UO_356 (O_356,N_19921,N_19981);
or UO_357 (O_357,N_19856,N_19955);
and UO_358 (O_358,N_19870,N_19914);
xor UO_359 (O_359,N_19830,N_19947);
nor UO_360 (O_360,N_19844,N_19894);
and UO_361 (O_361,N_19923,N_19859);
nor UO_362 (O_362,N_19853,N_19844);
or UO_363 (O_363,N_19956,N_19888);
or UO_364 (O_364,N_19881,N_19893);
nor UO_365 (O_365,N_19825,N_19955);
nand UO_366 (O_366,N_19932,N_19937);
or UO_367 (O_367,N_19897,N_19964);
nand UO_368 (O_368,N_19823,N_19882);
nor UO_369 (O_369,N_19866,N_19972);
nand UO_370 (O_370,N_19993,N_19835);
nor UO_371 (O_371,N_19941,N_19991);
or UO_372 (O_372,N_19874,N_19810);
nand UO_373 (O_373,N_19913,N_19917);
or UO_374 (O_374,N_19892,N_19809);
nor UO_375 (O_375,N_19978,N_19957);
nor UO_376 (O_376,N_19809,N_19931);
nor UO_377 (O_377,N_19880,N_19874);
nand UO_378 (O_378,N_19900,N_19966);
and UO_379 (O_379,N_19991,N_19826);
nand UO_380 (O_380,N_19992,N_19835);
and UO_381 (O_381,N_19989,N_19870);
and UO_382 (O_382,N_19986,N_19835);
nand UO_383 (O_383,N_19925,N_19961);
nand UO_384 (O_384,N_19998,N_19931);
or UO_385 (O_385,N_19859,N_19992);
nor UO_386 (O_386,N_19882,N_19963);
nor UO_387 (O_387,N_19947,N_19870);
xnor UO_388 (O_388,N_19934,N_19806);
nor UO_389 (O_389,N_19970,N_19950);
and UO_390 (O_390,N_19850,N_19941);
and UO_391 (O_391,N_19850,N_19815);
nor UO_392 (O_392,N_19804,N_19877);
or UO_393 (O_393,N_19931,N_19930);
and UO_394 (O_394,N_19828,N_19818);
nor UO_395 (O_395,N_19879,N_19967);
nor UO_396 (O_396,N_19976,N_19810);
nand UO_397 (O_397,N_19978,N_19974);
nand UO_398 (O_398,N_19873,N_19834);
nor UO_399 (O_399,N_19879,N_19973);
or UO_400 (O_400,N_19995,N_19843);
and UO_401 (O_401,N_19839,N_19830);
nor UO_402 (O_402,N_19979,N_19855);
nand UO_403 (O_403,N_19917,N_19990);
or UO_404 (O_404,N_19962,N_19938);
or UO_405 (O_405,N_19840,N_19936);
nor UO_406 (O_406,N_19961,N_19892);
and UO_407 (O_407,N_19924,N_19855);
nand UO_408 (O_408,N_19862,N_19828);
or UO_409 (O_409,N_19905,N_19926);
nand UO_410 (O_410,N_19837,N_19928);
or UO_411 (O_411,N_19852,N_19952);
or UO_412 (O_412,N_19924,N_19898);
nand UO_413 (O_413,N_19879,N_19824);
xnor UO_414 (O_414,N_19851,N_19868);
and UO_415 (O_415,N_19965,N_19916);
and UO_416 (O_416,N_19882,N_19892);
nand UO_417 (O_417,N_19822,N_19864);
nor UO_418 (O_418,N_19976,N_19806);
nor UO_419 (O_419,N_19907,N_19990);
or UO_420 (O_420,N_19886,N_19815);
and UO_421 (O_421,N_19978,N_19809);
nor UO_422 (O_422,N_19996,N_19928);
or UO_423 (O_423,N_19980,N_19854);
nand UO_424 (O_424,N_19924,N_19896);
nand UO_425 (O_425,N_19853,N_19870);
nor UO_426 (O_426,N_19895,N_19817);
or UO_427 (O_427,N_19889,N_19935);
nand UO_428 (O_428,N_19800,N_19826);
xor UO_429 (O_429,N_19941,N_19832);
nor UO_430 (O_430,N_19945,N_19877);
nor UO_431 (O_431,N_19842,N_19919);
or UO_432 (O_432,N_19972,N_19806);
and UO_433 (O_433,N_19911,N_19968);
or UO_434 (O_434,N_19860,N_19914);
or UO_435 (O_435,N_19987,N_19906);
and UO_436 (O_436,N_19978,N_19928);
and UO_437 (O_437,N_19936,N_19903);
or UO_438 (O_438,N_19965,N_19819);
nor UO_439 (O_439,N_19905,N_19859);
or UO_440 (O_440,N_19898,N_19862);
nor UO_441 (O_441,N_19965,N_19818);
nor UO_442 (O_442,N_19935,N_19865);
or UO_443 (O_443,N_19941,N_19895);
nand UO_444 (O_444,N_19887,N_19940);
nand UO_445 (O_445,N_19939,N_19877);
nor UO_446 (O_446,N_19958,N_19920);
nor UO_447 (O_447,N_19936,N_19993);
nor UO_448 (O_448,N_19857,N_19875);
nand UO_449 (O_449,N_19933,N_19816);
xor UO_450 (O_450,N_19960,N_19984);
and UO_451 (O_451,N_19881,N_19922);
nand UO_452 (O_452,N_19990,N_19927);
and UO_453 (O_453,N_19823,N_19892);
xor UO_454 (O_454,N_19995,N_19902);
and UO_455 (O_455,N_19807,N_19918);
nand UO_456 (O_456,N_19975,N_19826);
nand UO_457 (O_457,N_19902,N_19931);
nand UO_458 (O_458,N_19837,N_19870);
nand UO_459 (O_459,N_19839,N_19828);
and UO_460 (O_460,N_19829,N_19909);
and UO_461 (O_461,N_19908,N_19833);
and UO_462 (O_462,N_19810,N_19813);
nor UO_463 (O_463,N_19928,N_19895);
nor UO_464 (O_464,N_19944,N_19898);
nor UO_465 (O_465,N_19809,N_19837);
xor UO_466 (O_466,N_19987,N_19986);
nand UO_467 (O_467,N_19984,N_19991);
and UO_468 (O_468,N_19957,N_19901);
or UO_469 (O_469,N_19801,N_19823);
nor UO_470 (O_470,N_19917,N_19888);
or UO_471 (O_471,N_19988,N_19810);
xnor UO_472 (O_472,N_19959,N_19962);
nor UO_473 (O_473,N_19968,N_19826);
and UO_474 (O_474,N_19897,N_19878);
xor UO_475 (O_475,N_19815,N_19944);
nand UO_476 (O_476,N_19901,N_19925);
nor UO_477 (O_477,N_19846,N_19901);
nor UO_478 (O_478,N_19864,N_19937);
and UO_479 (O_479,N_19902,N_19956);
nand UO_480 (O_480,N_19860,N_19974);
nor UO_481 (O_481,N_19853,N_19822);
nand UO_482 (O_482,N_19946,N_19874);
nor UO_483 (O_483,N_19969,N_19918);
or UO_484 (O_484,N_19850,N_19928);
and UO_485 (O_485,N_19910,N_19801);
nand UO_486 (O_486,N_19888,N_19954);
nand UO_487 (O_487,N_19898,N_19936);
nand UO_488 (O_488,N_19836,N_19988);
and UO_489 (O_489,N_19900,N_19953);
and UO_490 (O_490,N_19853,N_19836);
nor UO_491 (O_491,N_19919,N_19887);
nand UO_492 (O_492,N_19916,N_19869);
and UO_493 (O_493,N_19870,N_19993);
nor UO_494 (O_494,N_19969,N_19901);
nand UO_495 (O_495,N_19993,N_19885);
nand UO_496 (O_496,N_19991,N_19813);
and UO_497 (O_497,N_19962,N_19840);
or UO_498 (O_498,N_19857,N_19862);
or UO_499 (O_499,N_19971,N_19973);
nor UO_500 (O_500,N_19907,N_19926);
nand UO_501 (O_501,N_19853,N_19896);
nand UO_502 (O_502,N_19966,N_19888);
nand UO_503 (O_503,N_19836,N_19968);
xor UO_504 (O_504,N_19957,N_19842);
or UO_505 (O_505,N_19883,N_19811);
or UO_506 (O_506,N_19976,N_19927);
nand UO_507 (O_507,N_19920,N_19850);
or UO_508 (O_508,N_19996,N_19964);
and UO_509 (O_509,N_19850,N_19977);
and UO_510 (O_510,N_19864,N_19806);
and UO_511 (O_511,N_19948,N_19823);
nand UO_512 (O_512,N_19845,N_19849);
and UO_513 (O_513,N_19838,N_19882);
and UO_514 (O_514,N_19941,N_19988);
nand UO_515 (O_515,N_19869,N_19939);
nor UO_516 (O_516,N_19975,N_19961);
nor UO_517 (O_517,N_19994,N_19849);
or UO_518 (O_518,N_19926,N_19902);
nor UO_519 (O_519,N_19980,N_19998);
and UO_520 (O_520,N_19836,N_19863);
nand UO_521 (O_521,N_19970,N_19819);
nor UO_522 (O_522,N_19956,N_19849);
or UO_523 (O_523,N_19802,N_19995);
and UO_524 (O_524,N_19967,N_19818);
and UO_525 (O_525,N_19804,N_19807);
or UO_526 (O_526,N_19829,N_19903);
nor UO_527 (O_527,N_19824,N_19814);
nor UO_528 (O_528,N_19924,N_19993);
and UO_529 (O_529,N_19829,N_19959);
or UO_530 (O_530,N_19849,N_19992);
nor UO_531 (O_531,N_19933,N_19890);
nor UO_532 (O_532,N_19808,N_19895);
and UO_533 (O_533,N_19823,N_19887);
or UO_534 (O_534,N_19943,N_19894);
nand UO_535 (O_535,N_19949,N_19992);
and UO_536 (O_536,N_19950,N_19861);
or UO_537 (O_537,N_19815,N_19902);
nand UO_538 (O_538,N_19839,N_19879);
or UO_539 (O_539,N_19857,N_19889);
nor UO_540 (O_540,N_19918,N_19861);
nand UO_541 (O_541,N_19940,N_19949);
and UO_542 (O_542,N_19822,N_19985);
nor UO_543 (O_543,N_19836,N_19983);
and UO_544 (O_544,N_19997,N_19815);
xnor UO_545 (O_545,N_19808,N_19835);
and UO_546 (O_546,N_19878,N_19954);
or UO_547 (O_547,N_19896,N_19995);
or UO_548 (O_548,N_19819,N_19901);
nand UO_549 (O_549,N_19811,N_19851);
nand UO_550 (O_550,N_19888,N_19990);
and UO_551 (O_551,N_19816,N_19996);
and UO_552 (O_552,N_19856,N_19879);
nand UO_553 (O_553,N_19962,N_19879);
or UO_554 (O_554,N_19879,N_19987);
and UO_555 (O_555,N_19815,N_19913);
and UO_556 (O_556,N_19868,N_19846);
or UO_557 (O_557,N_19804,N_19814);
nand UO_558 (O_558,N_19879,N_19845);
nor UO_559 (O_559,N_19871,N_19842);
or UO_560 (O_560,N_19889,N_19867);
or UO_561 (O_561,N_19926,N_19978);
and UO_562 (O_562,N_19904,N_19844);
nor UO_563 (O_563,N_19870,N_19842);
xnor UO_564 (O_564,N_19936,N_19951);
nor UO_565 (O_565,N_19991,N_19934);
and UO_566 (O_566,N_19957,N_19937);
nand UO_567 (O_567,N_19808,N_19979);
and UO_568 (O_568,N_19939,N_19853);
and UO_569 (O_569,N_19860,N_19934);
xor UO_570 (O_570,N_19950,N_19843);
nor UO_571 (O_571,N_19807,N_19942);
or UO_572 (O_572,N_19963,N_19877);
or UO_573 (O_573,N_19837,N_19862);
nor UO_574 (O_574,N_19893,N_19826);
or UO_575 (O_575,N_19988,N_19814);
or UO_576 (O_576,N_19882,N_19840);
nor UO_577 (O_577,N_19839,N_19993);
nand UO_578 (O_578,N_19909,N_19932);
and UO_579 (O_579,N_19896,N_19867);
xor UO_580 (O_580,N_19919,N_19876);
and UO_581 (O_581,N_19967,N_19954);
nor UO_582 (O_582,N_19954,N_19976);
or UO_583 (O_583,N_19924,N_19823);
nand UO_584 (O_584,N_19984,N_19827);
nand UO_585 (O_585,N_19931,N_19949);
or UO_586 (O_586,N_19853,N_19995);
nand UO_587 (O_587,N_19891,N_19873);
nand UO_588 (O_588,N_19925,N_19911);
nand UO_589 (O_589,N_19936,N_19838);
and UO_590 (O_590,N_19824,N_19870);
nor UO_591 (O_591,N_19987,N_19967);
nor UO_592 (O_592,N_19811,N_19810);
and UO_593 (O_593,N_19981,N_19885);
and UO_594 (O_594,N_19949,N_19975);
or UO_595 (O_595,N_19879,N_19976);
nor UO_596 (O_596,N_19996,N_19911);
nor UO_597 (O_597,N_19904,N_19922);
or UO_598 (O_598,N_19910,N_19870);
nor UO_599 (O_599,N_19960,N_19957);
and UO_600 (O_600,N_19984,N_19965);
nor UO_601 (O_601,N_19973,N_19870);
or UO_602 (O_602,N_19910,N_19825);
nand UO_603 (O_603,N_19903,N_19954);
nor UO_604 (O_604,N_19915,N_19926);
nand UO_605 (O_605,N_19923,N_19830);
and UO_606 (O_606,N_19869,N_19824);
or UO_607 (O_607,N_19912,N_19875);
nor UO_608 (O_608,N_19924,N_19848);
nor UO_609 (O_609,N_19878,N_19800);
and UO_610 (O_610,N_19900,N_19894);
or UO_611 (O_611,N_19807,N_19922);
and UO_612 (O_612,N_19990,N_19883);
nor UO_613 (O_613,N_19896,N_19888);
nand UO_614 (O_614,N_19962,N_19911);
nand UO_615 (O_615,N_19941,N_19808);
or UO_616 (O_616,N_19967,N_19848);
or UO_617 (O_617,N_19930,N_19887);
and UO_618 (O_618,N_19883,N_19961);
or UO_619 (O_619,N_19995,N_19987);
and UO_620 (O_620,N_19981,N_19802);
nor UO_621 (O_621,N_19990,N_19923);
nor UO_622 (O_622,N_19845,N_19941);
nor UO_623 (O_623,N_19874,N_19871);
and UO_624 (O_624,N_19837,N_19971);
nor UO_625 (O_625,N_19853,N_19925);
nand UO_626 (O_626,N_19821,N_19915);
nand UO_627 (O_627,N_19976,N_19889);
nand UO_628 (O_628,N_19840,N_19901);
nand UO_629 (O_629,N_19862,N_19843);
or UO_630 (O_630,N_19821,N_19823);
nand UO_631 (O_631,N_19931,N_19861);
nor UO_632 (O_632,N_19871,N_19937);
xnor UO_633 (O_633,N_19802,N_19894);
or UO_634 (O_634,N_19965,N_19809);
nand UO_635 (O_635,N_19809,N_19834);
nand UO_636 (O_636,N_19932,N_19969);
xor UO_637 (O_637,N_19858,N_19986);
nor UO_638 (O_638,N_19846,N_19942);
or UO_639 (O_639,N_19881,N_19801);
or UO_640 (O_640,N_19902,N_19971);
nand UO_641 (O_641,N_19812,N_19830);
and UO_642 (O_642,N_19989,N_19828);
nand UO_643 (O_643,N_19824,N_19978);
xor UO_644 (O_644,N_19802,N_19977);
nor UO_645 (O_645,N_19989,N_19927);
and UO_646 (O_646,N_19827,N_19936);
and UO_647 (O_647,N_19848,N_19903);
or UO_648 (O_648,N_19827,N_19903);
and UO_649 (O_649,N_19903,N_19919);
nor UO_650 (O_650,N_19889,N_19843);
and UO_651 (O_651,N_19849,N_19944);
nor UO_652 (O_652,N_19971,N_19923);
nand UO_653 (O_653,N_19864,N_19878);
nand UO_654 (O_654,N_19955,N_19828);
or UO_655 (O_655,N_19875,N_19852);
xor UO_656 (O_656,N_19830,N_19896);
nor UO_657 (O_657,N_19828,N_19913);
or UO_658 (O_658,N_19861,N_19887);
nor UO_659 (O_659,N_19830,N_19870);
nor UO_660 (O_660,N_19853,N_19996);
nor UO_661 (O_661,N_19978,N_19918);
nor UO_662 (O_662,N_19834,N_19915);
nand UO_663 (O_663,N_19888,N_19878);
and UO_664 (O_664,N_19941,N_19818);
and UO_665 (O_665,N_19823,N_19899);
nor UO_666 (O_666,N_19990,N_19909);
nand UO_667 (O_667,N_19985,N_19895);
or UO_668 (O_668,N_19852,N_19986);
nand UO_669 (O_669,N_19952,N_19950);
and UO_670 (O_670,N_19865,N_19929);
and UO_671 (O_671,N_19857,N_19950);
and UO_672 (O_672,N_19820,N_19862);
or UO_673 (O_673,N_19822,N_19914);
or UO_674 (O_674,N_19880,N_19841);
or UO_675 (O_675,N_19861,N_19901);
nor UO_676 (O_676,N_19869,N_19977);
nor UO_677 (O_677,N_19936,N_19891);
nand UO_678 (O_678,N_19894,N_19879);
nand UO_679 (O_679,N_19931,N_19954);
nand UO_680 (O_680,N_19853,N_19928);
nand UO_681 (O_681,N_19952,N_19917);
or UO_682 (O_682,N_19861,N_19819);
and UO_683 (O_683,N_19878,N_19930);
or UO_684 (O_684,N_19923,N_19955);
xnor UO_685 (O_685,N_19927,N_19946);
and UO_686 (O_686,N_19972,N_19861);
and UO_687 (O_687,N_19809,N_19884);
nor UO_688 (O_688,N_19829,N_19848);
nor UO_689 (O_689,N_19939,N_19880);
or UO_690 (O_690,N_19821,N_19956);
and UO_691 (O_691,N_19974,N_19807);
xnor UO_692 (O_692,N_19921,N_19976);
and UO_693 (O_693,N_19965,N_19866);
nor UO_694 (O_694,N_19933,N_19812);
or UO_695 (O_695,N_19920,N_19965);
nand UO_696 (O_696,N_19957,N_19909);
or UO_697 (O_697,N_19867,N_19863);
and UO_698 (O_698,N_19884,N_19874);
or UO_699 (O_699,N_19819,N_19984);
and UO_700 (O_700,N_19876,N_19813);
or UO_701 (O_701,N_19924,N_19857);
or UO_702 (O_702,N_19845,N_19897);
and UO_703 (O_703,N_19803,N_19822);
or UO_704 (O_704,N_19938,N_19864);
or UO_705 (O_705,N_19885,N_19847);
nand UO_706 (O_706,N_19923,N_19926);
or UO_707 (O_707,N_19987,N_19934);
and UO_708 (O_708,N_19863,N_19872);
and UO_709 (O_709,N_19854,N_19920);
xnor UO_710 (O_710,N_19971,N_19967);
nand UO_711 (O_711,N_19809,N_19805);
and UO_712 (O_712,N_19998,N_19895);
nand UO_713 (O_713,N_19969,N_19980);
or UO_714 (O_714,N_19988,N_19908);
xor UO_715 (O_715,N_19873,N_19893);
and UO_716 (O_716,N_19858,N_19873);
and UO_717 (O_717,N_19902,N_19894);
and UO_718 (O_718,N_19981,N_19955);
xor UO_719 (O_719,N_19954,N_19986);
and UO_720 (O_720,N_19975,N_19943);
nand UO_721 (O_721,N_19810,N_19843);
nand UO_722 (O_722,N_19984,N_19971);
nor UO_723 (O_723,N_19904,N_19970);
nand UO_724 (O_724,N_19820,N_19878);
and UO_725 (O_725,N_19813,N_19869);
or UO_726 (O_726,N_19821,N_19910);
and UO_727 (O_727,N_19965,N_19999);
and UO_728 (O_728,N_19838,N_19918);
and UO_729 (O_729,N_19834,N_19805);
nand UO_730 (O_730,N_19853,N_19812);
and UO_731 (O_731,N_19808,N_19850);
or UO_732 (O_732,N_19989,N_19886);
nand UO_733 (O_733,N_19872,N_19820);
nand UO_734 (O_734,N_19895,N_19825);
and UO_735 (O_735,N_19889,N_19813);
nand UO_736 (O_736,N_19934,N_19948);
nand UO_737 (O_737,N_19902,N_19801);
or UO_738 (O_738,N_19802,N_19896);
or UO_739 (O_739,N_19875,N_19911);
or UO_740 (O_740,N_19990,N_19851);
or UO_741 (O_741,N_19979,N_19869);
xnor UO_742 (O_742,N_19961,N_19852);
nor UO_743 (O_743,N_19870,N_19872);
nand UO_744 (O_744,N_19886,N_19934);
or UO_745 (O_745,N_19974,N_19929);
or UO_746 (O_746,N_19826,N_19886);
and UO_747 (O_747,N_19995,N_19994);
and UO_748 (O_748,N_19852,N_19990);
nand UO_749 (O_749,N_19900,N_19826);
nand UO_750 (O_750,N_19853,N_19831);
or UO_751 (O_751,N_19817,N_19950);
nand UO_752 (O_752,N_19972,N_19887);
nor UO_753 (O_753,N_19889,N_19957);
nand UO_754 (O_754,N_19858,N_19854);
nor UO_755 (O_755,N_19901,N_19873);
nor UO_756 (O_756,N_19875,N_19917);
or UO_757 (O_757,N_19919,N_19805);
and UO_758 (O_758,N_19918,N_19874);
nand UO_759 (O_759,N_19859,N_19828);
nor UO_760 (O_760,N_19861,N_19944);
or UO_761 (O_761,N_19820,N_19909);
and UO_762 (O_762,N_19942,N_19847);
nor UO_763 (O_763,N_19875,N_19998);
or UO_764 (O_764,N_19872,N_19813);
or UO_765 (O_765,N_19931,N_19990);
nand UO_766 (O_766,N_19924,N_19919);
or UO_767 (O_767,N_19973,N_19803);
nor UO_768 (O_768,N_19904,N_19917);
nor UO_769 (O_769,N_19960,N_19849);
and UO_770 (O_770,N_19939,N_19914);
xor UO_771 (O_771,N_19879,N_19970);
and UO_772 (O_772,N_19977,N_19884);
and UO_773 (O_773,N_19991,N_19930);
and UO_774 (O_774,N_19859,N_19812);
nor UO_775 (O_775,N_19992,N_19961);
nor UO_776 (O_776,N_19840,N_19811);
or UO_777 (O_777,N_19869,N_19833);
nand UO_778 (O_778,N_19827,N_19894);
or UO_779 (O_779,N_19833,N_19821);
nand UO_780 (O_780,N_19970,N_19984);
nor UO_781 (O_781,N_19812,N_19910);
and UO_782 (O_782,N_19883,N_19930);
or UO_783 (O_783,N_19823,N_19941);
nand UO_784 (O_784,N_19991,N_19928);
nand UO_785 (O_785,N_19860,N_19805);
or UO_786 (O_786,N_19920,N_19946);
nand UO_787 (O_787,N_19849,N_19817);
nand UO_788 (O_788,N_19859,N_19891);
xnor UO_789 (O_789,N_19929,N_19804);
or UO_790 (O_790,N_19823,N_19915);
nand UO_791 (O_791,N_19965,N_19937);
and UO_792 (O_792,N_19846,N_19813);
nor UO_793 (O_793,N_19897,N_19837);
nor UO_794 (O_794,N_19815,N_19973);
and UO_795 (O_795,N_19828,N_19947);
or UO_796 (O_796,N_19876,N_19851);
nor UO_797 (O_797,N_19985,N_19863);
nand UO_798 (O_798,N_19825,N_19970);
and UO_799 (O_799,N_19929,N_19803);
nand UO_800 (O_800,N_19904,N_19880);
and UO_801 (O_801,N_19946,N_19840);
and UO_802 (O_802,N_19896,N_19893);
or UO_803 (O_803,N_19873,N_19954);
nand UO_804 (O_804,N_19869,N_19863);
nor UO_805 (O_805,N_19885,N_19908);
or UO_806 (O_806,N_19835,N_19907);
or UO_807 (O_807,N_19960,N_19824);
or UO_808 (O_808,N_19913,N_19924);
nand UO_809 (O_809,N_19991,N_19822);
nor UO_810 (O_810,N_19819,N_19934);
or UO_811 (O_811,N_19981,N_19814);
and UO_812 (O_812,N_19931,N_19835);
nor UO_813 (O_813,N_19896,N_19862);
nor UO_814 (O_814,N_19884,N_19879);
or UO_815 (O_815,N_19984,N_19852);
or UO_816 (O_816,N_19906,N_19811);
nor UO_817 (O_817,N_19907,N_19979);
nor UO_818 (O_818,N_19825,N_19877);
and UO_819 (O_819,N_19928,N_19906);
or UO_820 (O_820,N_19961,N_19942);
nor UO_821 (O_821,N_19803,N_19909);
nor UO_822 (O_822,N_19816,N_19801);
nand UO_823 (O_823,N_19958,N_19850);
nor UO_824 (O_824,N_19958,N_19815);
xor UO_825 (O_825,N_19974,N_19853);
or UO_826 (O_826,N_19915,N_19890);
and UO_827 (O_827,N_19953,N_19861);
nand UO_828 (O_828,N_19993,N_19950);
nand UO_829 (O_829,N_19824,N_19857);
nand UO_830 (O_830,N_19909,N_19901);
nor UO_831 (O_831,N_19962,N_19980);
nor UO_832 (O_832,N_19998,N_19977);
nor UO_833 (O_833,N_19958,N_19873);
or UO_834 (O_834,N_19885,N_19888);
and UO_835 (O_835,N_19987,N_19999);
nor UO_836 (O_836,N_19889,N_19835);
xnor UO_837 (O_837,N_19887,N_19923);
or UO_838 (O_838,N_19818,N_19999);
nand UO_839 (O_839,N_19939,N_19829);
nand UO_840 (O_840,N_19953,N_19933);
nor UO_841 (O_841,N_19943,N_19991);
nor UO_842 (O_842,N_19987,N_19880);
nor UO_843 (O_843,N_19861,N_19974);
nor UO_844 (O_844,N_19932,N_19846);
nor UO_845 (O_845,N_19829,N_19988);
nand UO_846 (O_846,N_19800,N_19839);
or UO_847 (O_847,N_19832,N_19909);
and UO_848 (O_848,N_19936,N_19864);
or UO_849 (O_849,N_19984,N_19981);
and UO_850 (O_850,N_19941,N_19806);
or UO_851 (O_851,N_19972,N_19999);
nor UO_852 (O_852,N_19887,N_19929);
nand UO_853 (O_853,N_19932,N_19873);
and UO_854 (O_854,N_19946,N_19862);
nor UO_855 (O_855,N_19960,N_19905);
nor UO_856 (O_856,N_19845,N_19958);
nor UO_857 (O_857,N_19814,N_19986);
nor UO_858 (O_858,N_19898,N_19953);
xnor UO_859 (O_859,N_19814,N_19932);
or UO_860 (O_860,N_19991,N_19886);
or UO_861 (O_861,N_19987,N_19921);
nand UO_862 (O_862,N_19926,N_19839);
nor UO_863 (O_863,N_19877,N_19848);
and UO_864 (O_864,N_19872,N_19952);
and UO_865 (O_865,N_19821,N_19940);
and UO_866 (O_866,N_19803,N_19952);
or UO_867 (O_867,N_19829,N_19854);
nand UO_868 (O_868,N_19893,N_19917);
nor UO_869 (O_869,N_19897,N_19883);
and UO_870 (O_870,N_19998,N_19973);
nand UO_871 (O_871,N_19917,N_19831);
and UO_872 (O_872,N_19846,N_19979);
nand UO_873 (O_873,N_19909,N_19870);
nand UO_874 (O_874,N_19884,N_19841);
xor UO_875 (O_875,N_19895,N_19980);
nand UO_876 (O_876,N_19967,N_19931);
or UO_877 (O_877,N_19912,N_19932);
or UO_878 (O_878,N_19955,N_19937);
xor UO_879 (O_879,N_19856,N_19819);
or UO_880 (O_880,N_19985,N_19837);
or UO_881 (O_881,N_19850,N_19938);
nor UO_882 (O_882,N_19907,N_19906);
nand UO_883 (O_883,N_19962,N_19925);
nor UO_884 (O_884,N_19858,N_19845);
nand UO_885 (O_885,N_19864,N_19951);
or UO_886 (O_886,N_19867,N_19972);
and UO_887 (O_887,N_19968,N_19917);
nand UO_888 (O_888,N_19917,N_19998);
nor UO_889 (O_889,N_19813,N_19843);
or UO_890 (O_890,N_19962,N_19989);
nor UO_891 (O_891,N_19920,N_19975);
or UO_892 (O_892,N_19972,N_19890);
or UO_893 (O_893,N_19902,N_19979);
xor UO_894 (O_894,N_19970,N_19803);
nor UO_895 (O_895,N_19817,N_19887);
or UO_896 (O_896,N_19894,N_19909);
nand UO_897 (O_897,N_19964,N_19943);
and UO_898 (O_898,N_19891,N_19899);
nor UO_899 (O_899,N_19811,N_19953);
nor UO_900 (O_900,N_19849,N_19927);
nor UO_901 (O_901,N_19853,N_19887);
and UO_902 (O_902,N_19954,N_19909);
nand UO_903 (O_903,N_19922,N_19939);
or UO_904 (O_904,N_19874,N_19923);
nand UO_905 (O_905,N_19834,N_19939);
xor UO_906 (O_906,N_19995,N_19824);
or UO_907 (O_907,N_19822,N_19946);
nor UO_908 (O_908,N_19931,N_19955);
or UO_909 (O_909,N_19854,N_19861);
or UO_910 (O_910,N_19951,N_19914);
nor UO_911 (O_911,N_19852,N_19969);
nand UO_912 (O_912,N_19821,N_19974);
and UO_913 (O_913,N_19895,N_19898);
nand UO_914 (O_914,N_19870,N_19981);
nor UO_915 (O_915,N_19997,N_19922);
nand UO_916 (O_916,N_19803,N_19826);
and UO_917 (O_917,N_19870,N_19976);
or UO_918 (O_918,N_19809,N_19926);
or UO_919 (O_919,N_19914,N_19832);
nand UO_920 (O_920,N_19980,N_19924);
or UO_921 (O_921,N_19867,N_19885);
or UO_922 (O_922,N_19970,N_19809);
nor UO_923 (O_923,N_19883,N_19828);
and UO_924 (O_924,N_19873,N_19812);
and UO_925 (O_925,N_19891,N_19816);
nand UO_926 (O_926,N_19897,N_19873);
and UO_927 (O_927,N_19939,N_19948);
or UO_928 (O_928,N_19883,N_19853);
and UO_929 (O_929,N_19994,N_19970);
and UO_930 (O_930,N_19925,N_19941);
or UO_931 (O_931,N_19910,N_19872);
or UO_932 (O_932,N_19865,N_19850);
or UO_933 (O_933,N_19817,N_19824);
or UO_934 (O_934,N_19825,N_19886);
nor UO_935 (O_935,N_19985,N_19848);
or UO_936 (O_936,N_19815,N_19894);
and UO_937 (O_937,N_19988,N_19907);
or UO_938 (O_938,N_19991,N_19924);
or UO_939 (O_939,N_19820,N_19947);
or UO_940 (O_940,N_19999,N_19816);
nand UO_941 (O_941,N_19950,N_19972);
and UO_942 (O_942,N_19949,N_19862);
or UO_943 (O_943,N_19829,N_19819);
nand UO_944 (O_944,N_19864,N_19930);
or UO_945 (O_945,N_19832,N_19942);
and UO_946 (O_946,N_19892,N_19922);
and UO_947 (O_947,N_19861,N_19899);
or UO_948 (O_948,N_19919,N_19959);
or UO_949 (O_949,N_19810,N_19823);
nand UO_950 (O_950,N_19826,N_19980);
or UO_951 (O_951,N_19885,N_19942);
or UO_952 (O_952,N_19898,N_19850);
nor UO_953 (O_953,N_19827,N_19929);
nor UO_954 (O_954,N_19979,N_19961);
and UO_955 (O_955,N_19849,N_19940);
nor UO_956 (O_956,N_19817,N_19884);
or UO_957 (O_957,N_19960,N_19979);
nand UO_958 (O_958,N_19902,N_19835);
nand UO_959 (O_959,N_19972,N_19889);
nand UO_960 (O_960,N_19849,N_19912);
and UO_961 (O_961,N_19805,N_19966);
nor UO_962 (O_962,N_19959,N_19995);
and UO_963 (O_963,N_19941,N_19943);
nor UO_964 (O_964,N_19968,N_19822);
nor UO_965 (O_965,N_19980,N_19816);
and UO_966 (O_966,N_19827,N_19823);
nand UO_967 (O_967,N_19920,N_19985);
and UO_968 (O_968,N_19894,N_19865);
nand UO_969 (O_969,N_19837,N_19878);
or UO_970 (O_970,N_19963,N_19894);
or UO_971 (O_971,N_19963,N_19870);
nor UO_972 (O_972,N_19924,N_19935);
or UO_973 (O_973,N_19896,N_19824);
nor UO_974 (O_974,N_19878,N_19964);
or UO_975 (O_975,N_19911,N_19956);
and UO_976 (O_976,N_19886,N_19996);
nor UO_977 (O_977,N_19830,N_19949);
and UO_978 (O_978,N_19900,N_19915);
nor UO_979 (O_979,N_19863,N_19887);
nor UO_980 (O_980,N_19855,N_19956);
and UO_981 (O_981,N_19855,N_19918);
and UO_982 (O_982,N_19845,N_19818);
nor UO_983 (O_983,N_19999,N_19857);
and UO_984 (O_984,N_19917,N_19819);
or UO_985 (O_985,N_19903,N_19850);
or UO_986 (O_986,N_19885,N_19850);
and UO_987 (O_987,N_19809,N_19856);
nor UO_988 (O_988,N_19973,N_19819);
nor UO_989 (O_989,N_19876,N_19814);
nand UO_990 (O_990,N_19849,N_19888);
and UO_991 (O_991,N_19984,N_19933);
or UO_992 (O_992,N_19978,N_19826);
nor UO_993 (O_993,N_19943,N_19987);
or UO_994 (O_994,N_19916,N_19858);
or UO_995 (O_995,N_19997,N_19858);
or UO_996 (O_996,N_19848,N_19887);
and UO_997 (O_997,N_19909,N_19885);
and UO_998 (O_998,N_19920,N_19963);
and UO_999 (O_999,N_19859,N_19984);
nand UO_1000 (O_1000,N_19806,N_19951);
or UO_1001 (O_1001,N_19900,N_19877);
or UO_1002 (O_1002,N_19851,N_19892);
nor UO_1003 (O_1003,N_19858,N_19941);
or UO_1004 (O_1004,N_19875,N_19886);
or UO_1005 (O_1005,N_19884,N_19909);
and UO_1006 (O_1006,N_19954,N_19934);
and UO_1007 (O_1007,N_19893,N_19861);
nand UO_1008 (O_1008,N_19942,N_19806);
nand UO_1009 (O_1009,N_19894,N_19823);
or UO_1010 (O_1010,N_19952,N_19867);
and UO_1011 (O_1011,N_19890,N_19900);
nand UO_1012 (O_1012,N_19822,N_19999);
nor UO_1013 (O_1013,N_19897,N_19856);
nor UO_1014 (O_1014,N_19898,N_19876);
nor UO_1015 (O_1015,N_19823,N_19872);
nor UO_1016 (O_1016,N_19958,N_19915);
nor UO_1017 (O_1017,N_19885,N_19884);
and UO_1018 (O_1018,N_19875,N_19854);
nor UO_1019 (O_1019,N_19960,N_19835);
and UO_1020 (O_1020,N_19946,N_19969);
and UO_1021 (O_1021,N_19906,N_19914);
nor UO_1022 (O_1022,N_19971,N_19893);
and UO_1023 (O_1023,N_19813,N_19805);
and UO_1024 (O_1024,N_19913,N_19845);
or UO_1025 (O_1025,N_19990,N_19864);
nor UO_1026 (O_1026,N_19976,N_19890);
nor UO_1027 (O_1027,N_19869,N_19840);
or UO_1028 (O_1028,N_19944,N_19918);
nor UO_1029 (O_1029,N_19948,N_19868);
or UO_1030 (O_1030,N_19805,N_19932);
nand UO_1031 (O_1031,N_19836,N_19838);
or UO_1032 (O_1032,N_19889,N_19900);
nor UO_1033 (O_1033,N_19865,N_19889);
and UO_1034 (O_1034,N_19857,N_19871);
nor UO_1035 (O_1035,N_19861,N_19936);
nor UO_1036 (O_1036,N_19884,N_19924);
nor UO_1037 (O_1037,N_19952,N_19894);
or UO_1038 (O_1038,N_19912,N_19878);
nand UO_1039 (O_1039,N_19878,N_19942);
nor UO_1040 (O_1040,N_19941,N_19978);
nor UO_1041 (O_1041,N_19821,N_19981);
nand UO_1042 (O_1042,N_19815,N_19874);
nand UO_1043 (O_1043,N_19909,N_19903);
nor UO_1044 (O_1044,N_19986,N_19900);
nand UO_1045 (O_1045,N_19885,N_19921);
or UO_1046 (O_1046,N_19917,N_19812);
nor UO_1047 (O_1047,N_19962,N_19936);
or UO_1048 (O_1048,N_19850,N_19902);
nand UO_1049 (O_1049,N_19960,N_19876);
and UO_1050 (O_1050,N_19835,N_19858);
nor UO_1051 (O_1051,N_19984,N_19858);
xnor UO_1052 (O_1052,N_19998,N_19983);
nor UO_1053 (O_1053,N_19982,N_19943);
nand UO_1054 (O_1054,N_19974,N_19972);
nor UO_1055 (O_1055,N_19911,N_19810);
nand UO_1056 (O_1056,N_19890,N_19847);
and UO_1057 (O_1057,N_19880,N_19948);
and UO_1058 (O_1058,N_19959,N_19835);
or UO_1059 (O_1059,N_19907,N_19824);
nand UO_1060 (O_1060,N_19885,N_19965);
and UO_1061 (O_1061,N_19896,N_19922);
and UO_1062 (O_1062,N_19822,N_19810);
and UO_1063 (O_1063,N_19936,N_19940);
and UO_1064 (O_1064,N_19903,N_19856);
and UO_1065 (O_1065,N_19805,N_19998);
nor UO_1066 (O_1066,N_19939,N_19919);
nor UO_1067 (O_1067,N_19963,N_19922);
nor UO_1068 (O_1068,N_19873,N_19803);
nor UO_1069 (O_1069,N_19897,N_19853);
nand UO_1070 (O_1070,N_19942,N_19865);
nand UO_1071 (O_1071,N_19908,N_19930);
nor UO_1072 (O_1072,N_19831,N_19902);
and UO_1073 (O_1073,N_19804,N_19869);
or UO_1074 (O_1074,N_19997,N_19974);
and UO_1075 (O_1075,N_19962,N_19966);
and UO_1076 (O_1076,N_19993,N_19954);
or UO_1077 (O_1077,N_19982,N_19812);
or UO_1078 (O_1078,N_19919,N_19984);
nand UO_1079 (O_1079,N_19924,N_19907);
nand UO_1080 (O_1080,N_19800,N_19876);
nand UO_1081 (O_1081,N_19965,N_19947);
and UO_1082 (O_1082,N_19885,N_19975);
nand UO_1083 (O_1083,N_19922,N_19813);
or UO_1084 (O_1084,N_19955,N_19843);
nand UO_1085 (O_1085,N_19939,N_19938);
or UO_1086 (O_1086,N_19959,N_19839);
and UO_1087 (O_1087,N_19902,N_19978);
or UO_1088 (O_1088,N_19996,N_19936);
or UO_1089 (O_1089,N_19942,N_19935);
nand UO_1090 (O_1090,N_19947,N_19807);
nand UO_1091 (O_1091,N_19948,N_19884);
nand UO_1092 (O_1092,N_19939,N_19979);
nor UO_1093 (O_1093,N_19928,N_19847);
and UO_1094 (O_1094,N_19993,N_19939);
or UO_1095 (O_1095,N_19844,N_19817);
nor UO_1096 (O_1096,N_19857,N_19848);
nor UO_1097 (O_1097,N_19810,N_19965);
nor UO_1098 (O_1098,N_19891,N_19915);
or UO_1099 (O_1099,N_19991,N_19862);
nor UO_1100 (O_1100,N_19921,N_19992);
nor UO_1101 (O_1101,N_19961,N_19838);
and UO_1102 (O_1102,N_19960,N_19843);
nor UO_1103 (O_1103,N_19838,N_19867);
nor UO_1104 (O_1104,N_19970,N_19838);
nand UO_1105 (O_1105,N_19840,N_19837);
nand UO_1106 (O_1106,N_19848,N_19979);
or UO_1107 (O_1107,N_19812,N_19952);
and UO_1108 (O_1108,N_19903,N_19988);
or UO_1109 (O_1109,N_19875,N_19907);
or UO_1110 (O_1110,N_19889,N_19837);
and UO_1111 (O_1111,N_19808,N_19967);
nand UO_1112 (O_1112,N_19836,N_19960);
or UO_1113 (O_1113,N_19882,N_19929);
nor UO_1114 (O_1114,N_19871,N_19941);
and UO_1115 (O_1115,N_19953,N_19885);
nor UO_1116 (O_1116,N_19887,N_19825);
nor UO_1117 (O_1117,N_19871,N_19974);
nor UO_1118 (O_1118,N_19959,N_19924);
and UO_1119 (O_1119,N_19818,N_19844);
nor UO_1120 (O_1120,N_19869,N_19860);
nand UO_1121 (O_1121,N_19973,N_19829);
and UO_1122 (O_1122,N_19971,N_19867);
nand UO_1123 (O_1123,N_19883,N_19964);
or UO_1124 (O_1124,N_19945,N_19852);
or UO_1125 (O_1125,N_19939,N_19847);
nor UO_1126 (O_1126,N_19967,N_19957);
nand UO_1127 (O_1127,N_19859,N_19838);
nor UO_1128 (O_1128,N_19833,N_19827);
nor UO_1129 (O_1129,N_19854,N_19977);
and UO_1130 (O_1130,N_19855,N_19823);
and UO_1131 (O_1131,N_19964,N_19966);
nor UO_1132 (O_1132,N_19819,N_19823);
and UO_1133 (O_1133,N_19841,N_19950);
nand UO_1134 (O_1134,N_19966,N_19998);
and UO_1135 (O_1135,N_19860,N_19875);
nand UO_1136 (O_1136,N_19982,N_19995);
and UO_1137 (O_1137,N_19909,N_19808);
or UO_1138 (O_1138,N_19953,N_19800);
or UO_1139 (O_1139,N_19990,N_19943);
and UO_1140 (O_1140,N_19810,N_19829);
nand UO_1141 (O_1141,N_19914,N_19842);
nor UO_1142 (O_1142,N_19868,N_19806);
and UO_1143 (O_1143,N_19825,N_19812);
nor UO_1144 (O_1144,N_19936,N_19872);
and UO_1145 (O_1145,N_19906,N_19894);
nand UO_1146 (O_1146,N_19923,N_19913);
or UO_1147 (O_1147,N_19882,N_19935);
nand UO_1148 (O_1148,N_19911,N_19838);
nand UO_1149 (O_1149,N_19928,N_19893);
nand UO_1150 (O_1150,N_19809,N_19940);
and UO_1151 (O_1151,N_19872,N_19878);
nand UO_1152 (O_1152,N_19845,N_19948);
and UO_1153 (O_1153,N_19813,N_19918);
nor UO_1154 (O_1154,N_19856,N_19971);
xor UO_1155 (O_1155,N_19882,N_19869);
nand UO_1156 (O_1156,N_19999,N_19804);
or UO_1157 (O_1157,N_19973,N_19942);
xnor UO_1158 (O_1158,N_19846,N_19812);
nor UO_1159 (O_1159,N_19912,N_19877);
nor UO_1160 (O_1160,N_19996,N_19866);
nand UO_1161 (O_1161,N_19835,N_19983);
nor UO_1162 (O_1162,N_19945,N_19944);
nor UO_1163 (O_1163,N_19960,N_19912);
nor UO_1164 (O_1164,N_19934,N_19811);
nand UO_1165 (O_1165,N_19839,N_19917);
nor UO_1166 (O_1166,N_19898,N_19804);
and UO_1167 (O_1167,N_19927,N_19820);
nor UO_1168 (O_1168,N_19871,N_19938);
and UO_1169 (O_1169,N_19887,N_19846);
nand UO_1170 (O_1170,N_19969,N_19907);
or UO_1171 (O_1171,N_19927,N_19921);
and UO_1172 (O_1172,N_19918,N_19866);
nand UO_1173 (O_1173,N_19953,N_19846);
nand UO_1174 (O_1174,N_19949,N_19839);
nand UO_1175 (O_1175,N_19890,N_19838);
nand UO_1176 (O_1176,N_19963,N_19889);
and UO_1177 (O_1177,N_19876,N_19887);
and UO_1178 (O_1178,N_19989,N_19822);
nand UO_1179 (O_1179,N_19879,N_19993);
nor UO_1180 (O_1180,N_19969,N_19811);
nand UO_1181 (O_1181,N_19898,N_19921);
or UO_1182 (O_1182,N_19983,N_19876);
or UO_1183 (O_1183,N_19830,N_19823);
nor UO_1184 (O_1184,N_19962,N_19917);
nand UO_1185 (O_1185,N_19834,N_19813);
nor UO_1186 (O_1186,N_19869,N_19801);
nor UO_1187 (O_1187,N_19807,N_19957);
or UO_1188 (O_1188,N_19954,N_19854);
or UO_1189 (O_1189,N_19863,N_19901);
or UO_1190 (O_1190,N_19812,N_19879);
and UO_1191 (O_1191,N_19905,N_19958);
or UO_1192 (O_1192,N_19822,N_19804);
nor UO_1193 (O_1193,N_19935,N_19825);
nor UO_1194 (O_1194,N_19849,N_19984);
nand UO_1195 (O_1195,N_19809,N_19934);
or UO_1196 (O_1196,N_19801,N_19920);
nand UO_1197 (O_1197,N_19883,N_19953);
nand UO_1198 (O_1198,N_19933,N_19966);
or UO_1199 (O_1199,N_19991,N_19836);
nand UO_1200 (O_1200,N_19800,N_19895);
nand UO_1201 (O_1201,N_19812,N_19989);
and UO_1202 (O_1202,N_19977,N_19913);
nand UO_1203 (O_1203,N_19960,N_19851);
nand UO_1204 (O_1204,N_19996,N_19954);
nor UO_1205 (O_1205,N_19885,N_19955);
xnor UO_1206 (O_1206,N_19838,N_19947);
or UO_1207 (O_1207,N_19842,N_19967);
and UO_1208 (O_1208,N_19887,N_19833);
and UO_1209 (O_1209,N_19866,N_19968);
or UO_1210 (O_1210,N_19947,N_19987);
nor UO_1211 (O_1211,N_19944,N_19986);
nand UO_1212 (O_1212,N_19851,N_19920);
nand UO_1213 (O_1213,N_19821,N_19972);
xor UO_1214 (O_1214,N_19970,N_19933);
nor UO_1215 (O_1215,N_19862,N_19859);
nand UO_1216 (O_1216,N_19836,N_19804);
xor UO_1217 (O_1217,N_19904,N_19874);
and UO_1218 (O_1218,N_19827,N_19879);
nor UO_1219 (O_1219,N_19827,N_19869);
or UO_1220 (O_1220,N_19848,N_19971);
nand UO_1221 (O_1221,N_19817,N_19996);
nor UO_1222 (O_1222,N_19816,N_19879);
nor UO_1223 (O_1223,N_19984,N_19876);
nor UO_1224 (O_1224,N_19865,N_19841);
nor UO_1225 (O_1225,N_19927,N_19811);
and UO_1226 (O_1226,N_19903,N_19866);
nor UO_1227 (O_1227,N_19945,N_19900);
and UO_1228 (O_1228,N_19975,N_19813);
nor UO_1229 (O_1229,N_19976,N_19917);
nand UO_1230 (O_1230,N_19870,N_19996);
or UO_1231 (O_1231,N_19925,N_19816);
nand UO_1232 (O_1232,N_19906,N_19805);
nor UO_1233 (O_1233,N_19980,N_19934);
or UO_1234 (O_1234,N_19860,N_19961);
xnor UO_1235 (O_1235,N_19976,N_19824);
nor UO_1236 (O_1236,N_19972,N_19814);
nand UO_1237 (O_1237,N_19937,N_19883);
nor UO_1238 (O_1238,N_19880,N_19923);
or UO_1239 (O_1239,N_19997,N_19853);
xnor UO_1240 (O_1240,N_19853,N_19842);
nor UO_1241 (O_1241,N_19809,N_19929);
nand UO_1242 (O_1242,N_19845,N_19875);
and UO_1243 (O_1243,N_19941,N_19888);
nor UO_1244 (O_1244,N_19887,N_19958);
nand UO_1245 (O_1245,N_19899,N_19892);
or UO_1246 (O_1246,N_19819,N_19922);
and UO_1247 (O_1247,N_19875,N_19805);
nor UO_1248 (O_1248,N_19905,N_19949);
xor UO_1249 (O_1249,N_19954,N_19919);
or UO_1250 (O_1250,N_19853,N_19813);
and UO_1251 (O_1251,N_19874,N_19986);
nor UO_1252 (O_1252,N_19987,N_19863);
and UO_1253 (O_1253,N_19854,N_19818);
or UO_1254 (O_1254,N_19923,N_19941);
or UO_1255 (O_1255,N_19845,N_19955);
and UO_1256 (O_1256,N_19861,N_19979);
or UO_1257 (O_1257,N_19852,N_19981);
nand UO_1258 (O_1258,N_19988,N_19826);
and UO_1259 (O_1259,N_19988,N_19820);
nand UO_1260 (O_1260,N_19973,N_19850);
nand UO_1261 (O_1261,N_19835,N_19836);
and UO_1262 (O_1262,N_19890,N_19925);
and UO_1263 (O_1263,N_19929,N_19869);
or UO_1264 (O_1264,N_19934,N_19868);
nor UO_1265 (O_1265,N_19946,N_19841);
and UO_1266 (O_1266,N_19870,N_19892);
nand UO_1267 (O_1267,N_19934,N_19925);
xnor UO_1268 (O_1268,N_19845,N_19892);
nand UO_1269 (O_1269,N_19946,N_19805);
nand UO_1270 (O_1270,N_19961,N_19888);
nand UO_1271 (O_1271,N_19823,N_19998);
and UO_1272 (O_1272,N_19876,N_19927);
or UO_1273 (O_1273,N_19818,N_19830);
and UO_1274 (O_1274,N_19802,N_19961);
xor UO_1275 (O_1275,N_19855,N_19994);
or UO_1276 (O_1276,N_19915,N_19853);
or UO_1277 (O_1277,N_19877,N_19983);
or UO_1278 (O_1278,N_19985,N_19818);
and UO_1279 (O_1279,N_19832,N_19893);
and UO_1280 (O_1280,N_19820,N_19930);
nand UO_1281 (O_1281,N_19999,N_19955);
nand UO_1282 (O_1282,N_19908,N_19852);
or UO_1283 (O_1283,N_19871,N_19849);
nand UO_1284 (O_1284,N_19911,N_19939);
nand UO_1285 (O_1285,N_19876,N_19802);
nand UO_1286 (O_1286,N_19889,N_19978);
nand UO_1287 (O_1287,N_19863,N_19816);
nand UO_1288 (O_1288,N_19914,N_19952);
nor UO_1289 (O_1289,N_19808,N_19902);
nand UO_1290 (O_1290,N_19808,N_19969);
nand UO_1291 (O_1291,N_19808,N_19958);
nor UO_1292 (O_1292,N_19997,N_19936);
nand UO_1293 (O_1293,N_19939,N_19861);
nor UO_1294 (O_1294,N_19834,N_19961);
or UO_1295 (O_1295,N_19822,N_19885);
xor UO_1296 (O_1296,N_19838,N_19904);
nor UO_1297 (O_1297,N_19829,N_19976);
and UO_1298 (O_1298,N_19871,N_19940);
nor UO_1299 (O_1299,N_19869,N_19902);
or UO_1300 (O_1300,N_19940,N_19839);
and UO_1301 (O_1301,N_19847,N_19802);
nand UO_1302 (O_1302,N_19846,N_19967);
nand UO_1303 (O_1303,N_19906,N_19886);
nand UO_1304 (O_1304,N_19963,N_19851);
nand UO_1305 (O_1305,N_19851,N_19959);
nor UO_1306 (O_1306,N_19900,N_19897);
or UO_1307 (O_1307,N_19895,N_19812);
or UO_1308 (O_1308,N_19928,N_19817);
and UO_1309 (O_1309,N_19877,N_19978);
xor UO_1310 (O_1310,N_19839,N_19946);
nand UO_1311 (O_1311,N_19931,N_19884);
or UO_1312 (O_1312,N_19850,N_19910);
and UO_1313 (O_1313,N_19985,N_19808);
nand UO_1314 (O_1314,N_19954,N_19876);
or UO_1315 (O_1315,N_19998,N_19883);
or UO_1316 (O_1316,N_19840,N_19874);
or UO_1317 (O_1317,N_19805,N_19899);
nand UO_1318 (O_1318,N_19826,N_19974);
and UO_1319 (O_1319,N_19825,N_19872);
xnor UO_1320 (O_1320,N_19957,N_19876);
nand UO_1321 (O_1321,N_19972,N_19810);
and UO_1322 (O_1322,N_19926,N_19807);
xnor UO_1323 (O_1323,N_19851,N_19919);
xor UO_1324 (O_1324,N_19944,N_19821);
nor UO_1325 (O_1325,N_19975,N_19968);
or UO_1326 (O_1326,N_19820,N_19816);
nor UO_1327 (O_1327,N_19940,N_19895);
or UO_1328 (O_1328,N_19818,N_19803);
nor UO_1329 (O_1329,N_19890,N_19857);
or UO_1330 (O_1330,N_19802,N_19815);
nor UO_1331 (O_1331,N_19865,N_19991);
and UO_1332 (O_1332,N_19979,N_19862);
nor UO_1333 (O_1333,N_19855,N_19822);
or UO_1334 (O_1334,N_19910,N_19859);
and UO_1335 (O_1335,N_19949,N_19853);
and UO_1336 (O_1336,N_19837,N_19852);
or UO_1337 (O_1337,N_19987,N_19881);
or UO_1338 (O_1338,N_19883,N_19851);
nor UO_1339 (O_1339,N_19896,N_19866);
and UO_1340 (O_1340,N_19912,N_19979);
and UO_1341 (O_1341,N_19938,N_19900);
nand UO_1342 (O_1342,N_19933,N_19839);
or UO_1343 (O_1343,N_19876,N_19862);
nor UO_1344 (O_1344,N_19903,N_19849);
nor UO_1345 (O_1345,N_19856,N_19872);
nand UO_1346 (O_1346,N_19811,N_19938);
and UO_1347 (O_1347,N_19826,N_19914);
or UO_1348 (O_1348,N_19811,N_19897);
and UO_1349 (O_1349,N_19996,N_19804);
nor UO_1350 (O_1350,N_19848,N_19810);
xor UO_1351 (O_1351,N_19815,N_19962);
nand UO_1352 (O_1352,N_19890,N_19853);
nand UO_1353 (O_1353,N_19927,N_19933);
or UO_1354 (O_1354,N_19911,N_19890);
nand UO_1355 (O_1355,N_19940,N_19818);
and UO_1356 (O_1356,N_19902,N_19852);
and UO_1357 (O_1357,N_19811,N_19915);
nand UO_1358 (O_1358,N_19894,N_19821);
and UO_1359 (O_1359,N_19914,N_19932);
or UO_1360 (O_1360,N_19948,N_19892);
nand UO_1361 (O_1361,N_19843,N_19834);
and UO_1362 (O_1362,N_19991,N_19868);
nand UO_1363 (O_1363,N_19871,N_19823);
and UO_1364 (O_1364,N_19906,N_19808);
and UO_1365 (O_1365,N_19996,N_19881);
nor UO_1366 (O_1366,N_19965,N_19895);
nor UO_1367 (O_1367,N_19879,N_19996);
nor UO_1368 (O_1368,N_19848,N_19820);
xnor UO_1369 (O_1369,N_19803,N_19984);
or UO_1370 (O_1370,N_19906,N_19812);
nor UO_1371 (O_1371,N_19983,N_19912);
and UO_1372 (O_1372,N_19823,N_19861);
nand UO_1373 (O_1373,N_19901,N_19804);
nor UO_1374 (O_1374,N_19860,N_19815);
or UO_1375 (O_1375,N_19946,N_19909);
and UO_1376 (O_1376,N_19886,N_19889);
nor UO_1377 (O_1377,N_19979,N_19906);
and UO_1378 (O_1378,N_19823,N_19912);
and UO_1379 (O_1379,N_19980,N_19915);
and UO_1380 (O_1380,N_19958,N_19911);
nor UO_1381 (O_1381,N_19868,N_19983);
nand UO_1382 (O_1382,N_19987,N_19807);
or UO_1383 (O_1383,N_19984,N_19818);
nand UO_1384 (O_1384,N_19955,N_19870);
or UO_1385 (O_1385,N_19852,N_19894);
xnor UO_1386 (O_1386,N_19897,N_19889);
nand UO_1387 (O_1387,N_19968,N_19965);
nor UO_1388 (O_1388,N_19813,N_19952);
or UO_1389 (O_1389,N_19861,N_19802);
nand UO_1390 (O_1390,N_19816,N_19939);
and UO_1391 (O_1391,N_19867,N_19960);
xnor UO_1392 (O_1392,N_19878,N_19844);
nand UO_1393 (O_1393,N_19883,N_19852);
nand UO_1394 (O_1394,N_19885,N_19945);
or UO_1395 (O_1395,N_19815,N_19856);
and UO_1396 (O_1396,N_19878,N_19949);
nand UO_1397 (O_1397,N_19954,N_19824);
and UO_1398 (O_1398,N_19896,N_19955);
nor UO_1399 (O_1399,N_19860,N_19933);
nor UO_1400 (O_1400,N_19852,N_19898);
or UO_1401 (O_1401,N_19836,N_19986);
or UO_1402 (O_1402,N_19820,N_19875);
and UO_1403 (O_1403,N_19993,N_19994);
or UO_1404 (O_1404,N_19904,N_19889);
and UO_1405 (O_1405,N_19803,N_19886);
or UO_1406 (O_1406,N_19809,N_19955);
nand UO_1407 (O_1407,N_19977,N_19867);
nor UO_1408 (O_1408,N_19831,N_19931);
nand UO_1409 (O_1409,N_19824,N_19892);
nor UO_1410 (O_1410,N_19816,N_19865);
nor UO_1411 (O_1411,N_19875,N_19950);
nand UO_1412 (O_1412,N_19851,N_19970);
nand UO_1413 (O_1413,N_19955,N_19997);
nor UO_1414 (O_1414,N_19965,N_19862);
xnor UO_1415 (O_1415,N_19888,N_19841);
and UO_1416 (O_1416,N_19989,N_19956);
nor UO_1417 (O_1417,N_19814,N_19965);
nor UO_1418 (O_1418,N_19944,N_19873);
nor UO_1419 (O_1419,N_19830,N_19968);
and UO_1420 (O_1420,N_19878,N_19866);
nor UO_1421 (O_1421,N_19924,N_19946);
or UO_1422 (O_1422,N_19926,N_19968);
xnor UO_1423 (O_1423,N_19965,N_19850);
nor UO_1424 (O_1424,N_19949,N_19938);
and UO_1425 (O_1425,N_19804,N_19868);
nor UO_1426 (O_1426,N_19990,N_19960);
and UO_1427 (O_1427,N_19907,N_19955);
nand UO_1428 (O_1428,N_19916,N_19978);
nand UO_1429 (O_1429,N_19945,N_19948);
or UO_1430 (O_1430,N_19820,N_19983);
or UO_1431 (O_1431,N_19982,N_19860);
nand UO_1432 (O_1432,N_19931,N_19940);
or UO_1433 (O_1433,N_19877,N_19889);
or UO_1434 (O_1434,N_19953,N_19847);
or UO_1435 (O_1435,N_19890,N_19950);
nand UO_1436 (O_1436,N_19883,N_19881);
nor UO_1437 (O_1437,N_19922,N_19976);
xor UO_1438 (O_1438,N_19868,N_19979);
or UO_1439 (O_1439,N_19841,N_19842);
nand UO_1440 (O_1440,N_19814,N_19812);
or UO_1441 (O_1441,N_19823,N_19951);
nor UO_1442 (O_1442,N_19946,N_19960);
nand UO_1443 (O_1443,N_19898,N_19836);
nor UO_1444 (O_1444,N_19858,N_19847);
nand UO_1445 (O_1445,N_19863,N_19918);
nand UO_1446 (O_1446,N_19940,N_19898);
and UO_1447 (O_1447,N_19840,N_19818);
or UO_1448 (O_1448,N_19924,N_19905);
nor UO_1449 (O_1449,N_19896,N_19869);
nor UO_1450 (O_1450,N_19957,N_19880);
nand UO_1451 (O_1451,N_19807,N_19916);
or UO_1452 (O_1452,N_19804,N_19889);
nor UO_1453 (O_1453,N_19950,N_19918);
nand UO_1454 (O_1454,N_19854,N_19844);
nand UO_1455 (O_1455,N_19846,N_19943);
and UO_1456 (O_1456,N_19959,N_19917);
or UO_1457 (O_1457,N_19960,N_19880);
and UO_1458 (O_1458,N_19832,N_19974);
nand UO_1459 (O_1459,N_19840,N_19856);
or UO_1460 (O_1460,N_19976,N_19947);
nor UO_1461 (O_1461,N_19812,N_19993);
nor UO_1462 (O_1462,N_19821,N_19859);
and UO_1463 (O_1463,N_19804,N_19920);
and UO_1464 (O_1464,N_19902,N_19805);
and UO_1465 (O_1465,N_19996,N_19856);
and UO_1466 (O_1466,N_19943,N_19929);
nor UO_1467 (O_1467,N_19948,N_19959);
and UO_1468 (O_1468,N_19932,N_19854);
nor UO_1469 (O_1469,N_19961,N_19854);
nand UO_1470 (O_1470,N_19946,N_19935);
nor UO_1471 (O_1471,N_19845,N_19824);
and UO_1472 (O_1472,N_19884,N_19894);
nand UO_1473 (O_1473,N_19855,N_19876);
xor UO_1474 (O_1474,N_19893,N_19977);
and UO_1475 (O_1475,N_19997,N_19844);
and UO_1476 (O_1476,N_19899,N_19991);
xnor UO_1477 (O_1477,N_19839,N_19853);
nand UO_1478 (O_1478,N_19866,N_19952);
nand UO_1479 (O_1479,N_19882,N_19899);
and UO_1480 (O_1480,N_19934,N_19936);
nand UO_1481 (O_1481,N_19963,N_19865);
nand UO_1482 (O_1482,N_19904,N_19993);
nand UO_1483 (O_1483,N_19844,N_19924);
or UO_1484 (O_1484,N_19921,N_19956);
nor UO_1485 (O_1485,N_19852,N_19853);
or UO_1486 (O_1486,N_19800,N_19985);
or UO_1487 (O_1487,N_19859,N_19826);
or UO_1488 (O_1488,N_19849,N_19914);
nand UO_1489 (O_1489,N_19855,N_19803);
nand UO_1490 (O_1490,N_19901,N_19999);
and UO_1491 (O_1491,N_19882,N_19988);
nor UO_1492 (O_1492,N_19975,N_19946);
nor UO_1493 (O_1493,N_19803,N_19918);
nand UO_1494 (O_1494,N_19859,N_19938);
nor UO_1495 (O_1495,N_19921,N_19911);
nor UO_1496 (O_1496,N_19932,N_19985);
and UO_1497 (O_1497,N_19927,N_19968);
and UO_1498 (O_1498,N_19919,N_19920);
nor UO_1499 (O_1499,N_19804,N_19971);
nand UO_1500 (O_1500,N_19911,N_19946);
and UO_1501 (O_1501,N_19985,N_19803);
xnor UO_1502 (O_1502,N_19842,N_19887);
nand UO_1503 (O_1503,N_19938,N_19964);
or UO_1504 (O_1504,N_19915,N_19909);
or UO_1505 (O_1505,N_19973,N_19849);
nand UO_1506 (O_1506,N_19882,N_19851);
nand UO_1507 (O_1507,N_19826,N_19899);
and UO_1508 (O_1508,N_19885,N_19808);
nand UO_1509 (O_1509,N_19836,N_19959);
or UO_1510 (O_1510,N_19916,N_19941);
nor UO_1511 (O_1511,N_19833,N_19964);
and UO_1512 (O_1512,N_19907,N_19855);
and UO_1513 (O_1513,N_19916,N_19824);
or UO_1514 (O_1514,N_19994,N_19905);
or UO_1515 (O_1515,N_19939,N_19967);
or UO_1516 (O_1516,N_19884,N_19932);
and UO_1517 (O_1517,N_19817,N_19981);
xor UO_1518 (O_1518,N_19873,N_19930);
nor UO_1519 (O_1519,N_19809,N_19914);
and UO_1520 (O_1520,N_19847,N_19877);
or UO_1521 (O_1521,N_19910,N_19912);
nor UO_1522 (O_1522,N_19837,N_19990);
or UO_1523 (O_1523,N_19903,N_19973);
or UO_1524 (O_1524,N_19970,N_19945);
and UO_1525 (O_1525,N_19914,N_19824);
nand UO_1526 (O_1526,N_19914,N_19805);
nand UO_1527 (O_1527,N_19922,N_19979);
or UO_1528 (O_1528,N_19961,N_19812);
and UO_1529 (O_1529,N_19844,N_19935);
nand UO_1530 (O_1530,N_19960,N_19975);
or UO_1531 (O_1531,N_19949,N_19893);
or UO_1532 (O_1532,N_19917,N_19903);
or UO_1533 (O_1533,N_19838,N_19801);
or UO_1534 (O_1534,N_19996,N_19890);
and UO_1535 (O_1535,N_19837,N_19838);
or UO_1536 (O_1536,N_19887,N_19947);
nor UO_1537 (O_1537,N_19823,N_19816);
nor UO_1538 (O_1538,N_19938,N_19986);
nand UO_1539 (O_1539,N_19825,N_19996);
or UO_1540 (O_1540,N_19808,N_19931);
or UO_1541 (O_1541,N_19992,N_19896);
nand UO_1542 (O_1542,N_19983,N_19939);
nand UO_1543 (O_1543,N_19874,N_19978);
nor UO_1544 (O_1544,N_19857,N_19951);
nand UO_1545 (O_1545,N_19856,N_19817);
nand UO_1546 (O_1546,N_19892,N_19965);
nand UO_1547 (O_1547,N_19882,N_19922);
or UO_1548 (O_1548,N_19838,N_19818);
nand UO_1549 (O_1549,N_19909,N_19862);
or UO_1550 (O_1550,N_19822,N_19879);
nor UO_1551 (O_1551,N_19987,N_19990);
nand UO_1552 (O_1552,N_19995,N_19978);
xnor UO_1553 (O_1553,N_19989,N_19967);
nand UO_1554 (O_1554,N_19814,N_19947);
nor UO_1555 (O_1555,N_19889,N_19985);
and UO_1556 (O_1556,N_19878,N_19849);
or UO_1557 (O_1557,N_19807,N_19801);
and UO_1558 (O_1558,N_19849,N_19893);
nor UO_1559 (O_1559,N_19991,N_19932);
nor UO_1560 (O_1560,N_19903,N_19996);
and UO_1561 (O_1561,N_19804,N_19863);
xnor UO_1562 (O_1562,N_19877,N_19941);
nand UO_1563 (O_1563,N_19868,N_19887);
nand UO_1564 (O_1564,N_19853,N_19832);
nor UO_1565 (O_1565,N_19838,N_19833);
and UO_1566 (O_1566,N_19939,N_19845);
or UO_1567 (O_1567,N_19802,N_19865);
nand UO_1568 (O_1568,N_19918,N_19930);
nand UO_1569 (O_1569,N_19832,N_19819);
nand UO_1570 (O_1570,N_19987,N_19922);
and UO_1571 (O_1571,N_19928,N_19857);
nand UO_1572 (O_1572,N_19862,N_19955);
and UO_1573 (O_1573,N_19919,N_19882);
nand UO_1574 (O_1574,N_19825,N_19843);
and UO_1575 (O_1575,N_19934,N_19879);
nor UO_1576 (O_1576,N_19808,N_19804);
nand UO_1577 (O_1577,N_19901,N_19872);
and UO_1578 (O_1578,N_19850,N_19951);
and UO_1579 (O_1579,N_19883,N_19842);
and UO_1580 (O_1580,N_19970,N_19952);
nand UO_1581 (O_1581,N_19821,N_19848);
or UO_1582 (O_1582,N_19930,N_19926);
and UO_1583 (O_1583,N_19867,N_19907);
or UO_1584 (O_1584,N_19954,N_19860);
or UO_1585 (O_1585,N_19845,N_19853);
and UO_1586 (O_1586,N_19812,N_19999);
and UO_1587 (O_1587,N_19810,N_19947);
nor UO_1588 (O_1588,N_19902,N_19867);
nand UO_1589 (O_1589,N_19899,N_19928);
or UO_1590 (O_1590,N_19955,N_19967);
nand UO_1591 (O_1591,N_19808,N_19892);
and UO_1592 (O_1592,N_19933,N_19881);
or UO_1593 (O_1593,N_19984,N_19985);
and UO_1594 (O_1594,N_19965,N_19988);
or UO_1595 (O_1595,N_19801,N_19928);
or UO_1596 (O_1596,N_19803,N_19807);
nor UO_1597 (O_1597,N_19919,N_19880);
and UO_1598 (O_1598,N_19840,N_19916);
nand UO_1599 (O_1599,N_19888,N_19860);
or UO_1600 (O_1600,N_19896,N_19984);
and UO_1601 (O_1601,N_19851,N_19836);
nor UO_1602 (O_1602,N_19972,N_19813);
nor UO_1603 (O_1603,N_19976,N_19996);
and UO_1604 (O_1604,N_19970,N_19864);
nand UO_1605 (O_1605,N_19900,N_19958);
nand UO_1606 (O_1606,N_19907,N_19914);
nor UO_1607 (O_1607,N_19945,N_19911);
and UO_1608 (O_1608,N_19846,N_19914);
nor UO_1609 (O_1609,N_19810,N_19860);
and UO_1610 (O_1610,N_19800,N_19950);
and UO_1611 (O_1611,N_19840,N_19898);
and UO_1612 (O_1612,N_19833,N_19904);
or UO_1613 (O_1613,N_19989,N_19879);
and UO_1614 (O_1614,N_19937,N_19982);
or UO_1615 (O_1615,N_19884,N_19899);
or UO_1616 (O_1616,N_19883,N_19955);
nand UO_1617 (O_1617,N_19961,N_19811);
nand UO_1618 (O_1618,N_19806,N_19952);
nand UO_1619 (O_1619,N_19872,N_19846);
and UO_1620 (O_1620,N_19974,N_19881);
nand UO_1621 (O_1621,N_19832,N_19960);
and UO_1622 (O_1622,N_19994,N_19937);
nor UO_1623 (O_1623,N_19903,N_19901);
nor UO_1624 (O_1624,N_19914,N_19808);
or UO_1625 (O_1625,N_19910,N_19922);
or UO_1626 (O_1626,N_19986,N_19935);
nor UO_1627 (O_1627,N_19985,N_19901);
or UO_1628 (O_1628,N_19848,N_19856);
nor UO_1629 (O_1629,N_19911,N_19994);
nand UO_1630 (O_1630,N_19871,N_19909);
xnor UO_1631 (O_1631,N_19853,N_19926);
nand UO_1632 (O_1632,N_19882,N_19901);
and UO_1633 (O_1633,N_19867,N_19805);
and UO_1634 (O_1634,N_19992,N_19970);
or UO_1635 (O_1635,N_19923,N_19937);
nand UO_1636 (O_1636,N_19839,N_19852);
nor UO_1637 (O_1637,N_19838,N_19869);
or UO_1638 (O_1638,N_19981,N_19948);
and UO_1639 (O_1639,N_19823,N_19826);
or UO_1640 (O_1640,N_19910,N_19864);
nor UO_1641 (O_1641,N_19844,N_19939);
nand UO_1642 (O_1642,N_19991,N_19828);
nor UO_1643 (O_1643,N_19906,N_19831);
nor UO_1644 (O_1644,N_19900,N_19923);
nand UO_1645 (O_1645,N_19884,N_19859);
nor UO_1646 (O_1646,N_19835,N_19834);
nor UO_1647 (O_1647,N_19922,N_19946);
nand UO_1648 (O_1648,N_19810,N_19892);
or UO_1649 (O_1649,N_19805,N_19823);
or UO_1650 (O_1650,N_19982,N_19979);
and UO_1651 (O_1651,N_19917,N_19874);
nor UO_1652 (O_1652,N_19886,N_19963);
or UO_1653 (O_1653,N_19868,N_19816);
and UO_1654 (O_1654,N_19864,N_19956);
nand UO_1655 (O_1655,N_19803,N_19890);
or UO_1656 (O_1656,N_19942,N_19820);
xnor UO_1657 (O_1657,N_19875,N_19881);
nor UO_1658 (O_1658,N_19966,N_19907);
or UO_1659 (O_1659,N_19977,N_19933);
or UO_1660 (O_1660,N_19925,N_19960);
or UO_1661 (O_1661,N_19956,N_19832);
nand UO_1662 (O_1662,N_19903,N_19933);
nor UO_1663 (O_1663,N_19890,N_19931);
nor UO_1664 (O_1664,N_19882,N_19826);
nand UO_1665 (O_1665,N_19841,N_19957);
and UO_1666 (O_1666,N_19900,N_19971);
or UO_1667 (O_1667,N_19908,N_19883);
nor UO_1668 (O_1668,N_19856,N_19924);
nor UO_1669 (O_1669,N_19892,N_19910);
or UO_1670 (O_1670,N_19809,N_19967);
and UO_1671 (O_1671,N_19807,N_19906);
nand UO_1672 (O_1672,N_19874,N_19805);
nand UO_1673 (O_1673,N_19802,N_19898);
nor UO_1674 (O_1674,N_19878,N_19874);
nor UO_1675 (O_1675,N_19991,N_19942);
nor UO_1676 (O_1676,N_19911,N_19846);
or UO_1677 (O_1677,N_19850,N_19890);
and UO_1678 (O_1678,N_19861,N_19815);
or UO_1679 (O_1679,N_19841,N_19997);
nand UO_1680 (O_1680,N_19957,N_19839);
or UO_1681 (O_1681,N_19906,N_19842);
and UO_1682 (O_1682,N_19893,N_19872);
nor UO_1683 (O_1683,N_19842,N_19856);
or UO_1684 (O_1684,N_19866,N_19875);
and UO_1685 (O_1685,N_19967,N_19928);
nor UO_1686 (O_1686,N_19981,N_19806);
and UO_1687 (O_1687,N_19950,N_19924);
nand UO_1688 (O_1688,N_19892,N_19928);
and UO_1689 (O_1689,N_19887,N_19990);
nand UO_1690 (O_1690,N_19872,N_19814);
nand UO_1691 (O_1691,N_19816,N_19856);
nand UO_1692 (O_1692,N_19824,N_19902);
and UO_1693 (O_1693,N_19929,N_19948);
and UO_1694 (O_1694,N_19955,N_19861);
and UO_1695 (O_1695,N_19800,N_19984);
nor UO_1696 (O_1696,N_19929,N_19916);
nand UO_1697 (O_1697,N_19892,N_19955);
nor UO_1698 (O_1698,N_19851,N_19911);
xor UO_1699 (O_1699,N_19907,N_19834);
nor UO_1700 (O_1700,N_19987,N_19954);
or UO_1701 (O_1701,N_19904,N_19823);
nor UO_1702 (O_1702,N_19826,N_19865);
xnor UO_1703 (O_1703,N_19891,N_19829);
and UO_1704 (O_1704,N_19897,N_19962);
nor UO_1705 (O_1705,N_19872,N_19852);
and UO_1706 (O_1706,N_19825,N_19830);
or UO_1707 (O_1707,N_19910,N_19931);
nand UO_1708 (O_1708,N_19915,N_19882);
or UO_1709 (O_1709,N_19816,N_19825);
and UO_1710 (O_1710,N_19954,N_19892);
nor UO_1711 (O_1711,N_19869,N_19936);
nor UO_1712 (O_1712,N_19861,N_19824);
nor UO_1713 (O_1713,N_19984,N_19899);
and UO_1714 (O_1714,N_19866,N_19970);
nor UO_1715 (O_1715,N_19926,N_19880);
nor UO_1716 (O_1716,N_19934,N_19862);
and UO_1717 (O_1717,N_19868,N_19937);
or UO_1718 (O_1718,N_19914,N_19848);
nor UO_1719 (O_1719,N_19841,N_19902);
nor UO_1720 (O_1720,N_19849,N_19859);
and UO_1721 (O_1721,N_19948,N_19803);
and UO_1722 (O_1722,N_19896,N_19929);
nor UO_1723 (O_1723,N_19886,N_19914);
nand UO_1724 (O_1724,N_19844,N_19883);
nor UO_1725 (O_1725,N_19844,N_19889);
nand UO_1726 (O_1726,N_19833,N_19956);
nor UO_1727 (O_1727,N_19937,N_19934);
or UO_1728 (O_1728,N_19853,N_19877);
or UO_1729 (O_1729,N_19940,N_19984);
nor UO_1730 (O_1730,N_19835,N_19950);
xor UO_1731 (O_1731,N_19805,N_19950);
xnor UO_1732 (O_1732,N_19944,N_19840);
or UO_1733 (O_1733,N_19865,N_19955);
or UO_1734 (O_1734,N_19928,N_19994);
nor UO_1735 (O_1735,N_19873,N_19884);
or UO_1736 (O_1736,N_19976,N_19840);
nor UO_1737 (O_1737,N_19831,N_19857);
or UO_1738 (O_1738,N_19963,N_19981);
nor UO_1739 (O_1739,N_19937,N_19884);
and UO_1740 (O_1740,N_19839,N_19954);
nor UO_1741 (O_1741,N_19968,N_19954);
and UO_1742 (O_1742,N_19821,N_19890);
and UO_1743 (O_1743,N_19822,N_19887);
or UO_1744 (O_1744,N_19869,N_19811);
and UO_1745 (O_1745,N_19842,N_19933);
or UO_1746 (O_1746,N_19993,N_19894);
nand UO_1747 (O_1747,N_19945,N_19960);
nand UO_1748 (O_1748,N_19816,N_19885);
or UO_1749 (O_1749,N_19843,N_19835);
and UO_1750 (O_1750,N_19987,N_19923);
nand UO_1751 (O_1751,N_19916,N_19846);
nor UO_1752 (O_1752,N_19838,N_19815);
nand UO_1753 (O_1753,N_19863,N_19822);
or UO_1754 (O_1754,N_19996,N_19847);
nor UO_1755 (O_1755,N_19845,N_19829);
and UO_1756 (O_1756,N_19811,N_19874);
xor UO_1757 (O_1757,N_19810,N_19948);
nand UO_1758 (O_1758,N_19815,N_19979);
or UO_1759 (O_1759,N_19806,N_19911);
xor UO_1760 (O_1760,N_19865,N_19846);
nand UO_1761 (O_1761,N_19821,N_19997);
nand UO_1762 (O_1762,N_19957,N_19991);
and UO_1763 (O_1763,N_19985,N_19851);
nor UO_1764 (O_1764,N_19896,N_19945);
or UO_1765 (O_1765,N_19899,N_19850);
nor UO_1766 (O_1766,N_19816,N_19975);
or UO_1767 (O_1767,N_19947,N_19864);
xor UO_1768 (O_1768,N_19874,N_19832);
nor UO_1769 (O_1769,N_19900,N_19924);
or UO_1770 (O_1770,N_19842,N_19956);
and UO_1771 (O_1771,N_19850,N_19878);
nor UO_1772 (O_1772,N_19843,N_19856);
nor UO_1773 (O_1773,N_19888,N_19873);
nor UO_1774 (O_1774,N_19878,N_19934);
xor UO_1775 (O_1775,N_19921,N_19993);
and UO_1776 (O_1776,N_19998,N_19841);
or UO_1777 (O_1777,N_19886,N_19856);
nor UO_1778 (O_1778,N_19845,N_19867);
or UO_1779 (O_1779,N_19875,N_19888);
or UO_1780 (O_1780,N_19862,N_19882);
and UO_1781 (O_1781,N_19918,N_19912);
or UO_1782 (O_1782,N_19829,N_19817);
or UO_1783 (O_1783,N_19930,N_19955);
and UO_1784 (O_1784,N_19988,N_19839);
and UO_1785 (O_1785,N_19944,N_19917);
and UO_1786 (O_1786,N_19997,N_19814);
or UO_1787 (O_1787,N_19813,N_19861);
nand UO_1788 (O_1788,N_19855,N_19963);
or UO_1789 (O_1789,N_19926,N_19995);
or UO_1790 (O_1790,N_19970,N_19828);
nand UO_1791 (O_1791,N_19885,N_19914);
nor UO_1792 (O_1792,N_19979,N_19983);
nand UO_1793 (O_1793,N_19873,N_19815);
nor UO_1794 (O_1794,N_19848,N_19880);
and UO_1795 (O_1795,N_19840,N_19950);
and UO_1796 (O_1796,N_19804,N_19818);
or UO_1797 (O_1797,N_19966,N_19976);
and UO_1798 (O_1798,N_19867,N_19839);
or UO_1799 (O_1799,N_19895,N_19902);
and UO_1800 (O_1800,N_19940,N_19920);
or UO_1801 (O_1801,N_19938,N_19961);
and UO_1802 (O_1802,N_19980,N_19946);
xor UO_1803 (O_1803,N_19934,N_19889);
nor UO_1804 (O_1804,N_19938,N_19895);
nand UO_1805 (O_1805,N_19866,N_19876);
nand UO_1806 (O_1806,N_19835,N_19915);
or UO_1807 (O_1807,N_19944,N_19933);
nor UO_1808 (O_1808,N_19977,N_19819);
and UO_1809 (O_1809,N_19969,N_19816);
nor UO_1810 (O_1810,N_19978,N_19844);
nand UO_1811 (O_1811,N_19876,N_19861);
nand UO_1812 (O_1812,N_19930,N_19853);
or UO_1813 (O_1813,N_19999,N_19836);
and UO_1814 (O_1814,N_19946,N_19884);
and UO_1815 (O_1815,N_19821,N_19906);
or UO_1816 (O_1816,N_19950,N_19951);
or UO_1817 (O_1817,N_19846,N_19937);
xor UO_1818 (O_1818,N_19997,N_19999);
and UO_1819 (O_1819,N_19854,N_19963);
or UO_1820 (O_1820,N_19913,N_19852);
or UO_1821 (O_1821,N_19892,N_19988);
nor UO_1822 (O_1822,N_19972,N_19983);
or UO_1823 (O_1823,N_19830,N_19820);
xnor UO_1824 (O_1824,N_19947,N_19898);
and UO_1825 (O_1825,N_19807,N_19901);
nand UO_1826 (O_1826,N_19832,N_19814);
and UO_1827 (O_1827,N_19898,N_19970);
and UO_1828 (O_1828,N_19812,N_19874);
and UO_1829 (O_1829,N_19888,N_19871);
nand UO_1830 (O_1830,N_19952,N_19815);
xnor UO_1831 (O_1831,N_19856,N_19926);
nor UO_1832 (O_1832,N_19832,N_19843);
nor UO_1833 (O_1833,N_19978,N_19867);
or UO_1834 (O_1834,N_19848,N_19940);
and UO_1835 (O_1835,N_19936,N_19815);
or UO_1836 (O_1836,N_19809,N_19994);
and UO_1837 (O_1837,N_19819,N_19801);
or UO_1838 (O_1838,N_19835,N_19926);
or UO_1839 (O_1839,N_19991,N_19925);
nor UO_1840 (O_1840,N_19997,N_19892);
xnor UO_1841 (O_1841,N_19985,N_19875);
nand UO_1842 (O_1842,N_19864,N_19812);
or UO_1843 (O_1843,N_19816,N_19924);
nor UO_1844 (O_1844,N_19948,N_19995);
nand UO_1845 (O_1845,N_19939,N_19959);
and UO_1846 (O_1846,N_19987,N_19899);
nand UO_1847 (O_1847,N_19824,N_19838);
or UO_1848 (O_1848,N_19906,N_19990);
or UO_1849 (O_1849,N_19874,N_19902);
nand UO_1850 (O_1850,N_19892,N_19962);
nor UO_1851 (O_1851,N_19964,N_19936);
and UO_1852 (O_1852,N_19860,N_19905);
nand UO_1853 (O_1853,N_19855,N_19824);
or UO_1854 (O_1854,N_19849,N_19855);
or UO_1855 (O_1855,N_19837,N_19853);
nand UO_1856 (O_1856,N_19978,N_19997);
and UO_1857 (O_1857,N_19831,N_19939);
nand UO_1858 (O_1858,N_19956,N_19962);
nor UO_1859 (O_1859,N_19861,N_19946);
nor UO_1860 (O_1860,N_19857,N_19946);
nand UO_1861 (O_1861,N_19988,N_19835);
nor UO_1862 (O_1862,N_19866,N_19998);
and UO_1863 (O_1863,N_19933,N_19862);
nor UO_1864 (O_1864,N_19803,N_19997);
nor UO_1865 (O_1865,N_19800,N_19830);
or UO_1866 (O_1866,N_19879,N_19850);
and UO_1867 (O_1867,N_19897,N_19946);
nor UO_1868 (O_1868,N_19924,N_19972);
or UO_1869 (O_1869,N_19805,N_19955);
and UO_1870 (O_1870,N_19972,N_19858);
nand UO_1871 (O_1871,N_19986,N_19875);
or UO_1872 (O_1872,N_19954,N_19974);
and UO_1873 (O_1873,N_19895,N_19882);
nand UO_1874 (O_1874,N_19961,N_19855);
nand UO_1875 (O_1875,N_19993,N_19915);
and UO_1876 (O_1876,N_19865,N_19905);
nor UO_1877 (O_1877,N_19991,N_19893);
or UO_1878 (O_1878,N_19866,N_19884);
nand UO_1879 (O_1879,N_19967,N_19893);
nand UO_1880 (O_1880,N_19833,N_19860);
and UO_1881 (O_1881,N_19932,N_19966);
or UO_1882 (O_1882,N_19917,N_19849);
or UO_1883 (O_1883,N_19823,N_19897);
and UO_1884 (O_1884,N_19800,N_19991);
and UO_1885 (O_1885,N_19899,N_19920);
or UO_1886 (O_1886,N_19969,N_19802);
nor UO_1887 (O_1887,N_19858,N_19857);
nor UO_1888 (O_1888,N_19936,N_19885);
or UO_1889 (O_1889,N_19981,N_19892);
or UO_1890 (O_1890,N_19812,N_19826);
nand UO_1891 (O_1891,N_19875,N_19996);
or UO_1892 (O_1892,N_19845,N_19863);
nand UO_1893 (O_1893,N_19956,N_19976);
or UO_1894 (O_1894,N_19944,N_19811);
or UO_1895 (O_1895,N_19923,N_19960);
nand UO_1896 (O_1896,N_19820,N_19920);
nor UO_1897 (O_1897,N_19931,N_19977);
nand UO_1898 (O_1898,N_19814,N_19898);
nand UO_1899 (O_1899,N_19896,N_19870);
or UO_1900 (O_1900,N_19848,N_19828);
xnor UO_1901 (O_1901,N_19876,N_19988);
nand UO_1902 (O_1902,N_19930,N_19837);
nor UO_1903 (O_1903,N_19859,N_19811);
or UO_1904 (O_1904,N_19953,N_19911);
nor UO_1905 (O_1905,N_19812,N_19840);
nor UO_1906 (O_1906,N_19930,N_19859);
or UO_1907 (O_1907,N_19868,N_19856);
or UO_1908 (O_1908,N_19910,N_19856);
and UO_1909 (O_1909,N_19942,N_19953);
xor UO_1910 (O_1910,N_19995,N_19914);
and UO_1911 (O_1911,N_19857,N_19960);
nand UO_1912 (O_1912,N_19883,N_19985);
nor UO_1913 (O_1913,N_19928,N_19838);
and UO_1914 (O_1914,N_19916,N_19884);
and UO_1915 (O_1915,N_19838,N_19879);
nand UO_1916 (O_1916,N_19911,N_19826);
nand UO_1917 (O_1917,N_19812,N_19942);
nand UO_1918 (O_1918,N_19900,N_19990);
nand UO_1919 (O_1919,N_19903,N_19991);
nor UO_1920 (O_1920,N_19880,N_19940);
or UO_1921 (O_1921,N_19885,N_19933);
or UO_1922 (O_1922,N_19958,N_19819);
nand UO_1923 (O_1923,N_19921,N_19859);
nor UO_1924 (O_1924,N_19821,N_19916);
nor UO_1925 (O_1925,N_19847,N_19990);
or UO_1926 (O_1926,N_19854,N_19923);
and UO_1927 (O_1927,N_19975,N_19982);
and UO_1928 (O_1928,N_19862,N_19967);
nand UO_1929 (O_1929,N_19893,N_19810);
and UO_1930 (O_1930,N_19894,N_19885);
and UO_1931 (O_1931,N_19997,N_19826);
nand UO_1932 (O_1932,N_19988,N_19918);
and UO_1933 (O_1933,N_19878,N_19804);
and UO_1934 (O_1934,N_19971,N_19972);
nor UO_1935 (O_1935,N_19883,N_19872);
and UO_1936 (O_1936,N_19801,N_19942);
and UO_1937 (O_1937,N_19979,N_19977);
and UO_1938 (O_1938,N_19948,N_19839);
or UO_1939 (O_1939,N_19931,N_19860);
and UO_1940 (O_1940,N_19810,N_19975);
nand UO_1941 (O_1941,N_19966,N_19969);
nor UO_1942 (O_1942,N_19910,N_19818);
nand UO_1943 (O_1943,N_19821,N_19991);
or UO_1944 (O_1944,N_19984,N_19951);
and UO_1945 (O_1945,N_19886,N_19970);
xor UO_1946 (O_1946,N_19836,N_19962);
or UO_1947 (O_1947,N_19912,N_19839);
or UO_1948 (O_1948,N_19962,N_19842);
nor UO_1949 (O_1949,N_19866,N_19826);
nand UO_1950 (O_1950,N_19936,N_19995);
and UO_1951 (O_1951,N_19869,N_19943);
and UO_1952 (O_1952,N_19899,N_19827);
nor UO_1953 (O_1953,N_19946,N_19999);
nand UO_1954 (O_1954,N_19997,N_19944);
nand UO_1955 (O_1955,N_19819,N_19966);
nor UO_1956 (O_1956,N_19904,N_19912);
and UO_1957 (O_1957,N_19822,N_19995);
nor UO_1958 (O_1958,N_19830,N_19868);
nand UO_1959 (O_1959,N_19831,N_19973);
nor UO_1960 (O_1960,N_19951,N_19952);
or UO_1961 (O_1961,N_19928,N_19887);
nor UO_1962 (O_1962,N_19946,N_19993);
or UO_1963 (O_1963,N_19840,N_19853);
nand UO_1964 (O_1964,N_19895,N_19877);
nand UO_1965 (O_1965,N_19939,N_19926);
nor UO_1966 (O_1966,N_19923,N_19800);
or UO_1967 (O_1967,N_19947,N_19966);
and UO_1968 (O_1968,N_19822,N_19828);
nor UO_1969 (O_1969,N_19980,N_19994);
nor UO_1970 (O_1970,N_19978,N_19984);
nor UO_1971 (O_1971,N_19968,N_19967);
nor UO_1972 (O_1972,N_19999,N_19897);
or UO_1973 (O_1973,N_19990,N_19948);
nand UO_1974 (O_1974,N_19830,N_19998);
and UO_1975 (O_1975,N_19844,N_19974);
or UO_1976 (O_1976,N_19829,N_19813);
nand UO_1977 (O_1977,N_19957,N_19816);
and UO_1978 (O_1978,N_19867,N_19919);
nand UO_1979 (O_1979,N_19971,N_19954);
or UO_1980 (O_1980,N_19847,N_19915);
or UO_1981 (O_1981,N_19985,N_19876);
or UO_1982 (O_1982,N_19992,N_19922);
nor UO_1983 (O_1983,N_19921,N_19810);
and UO_1984 (O_1984,N_19899,N_19821);
and UO_1985 (O_1985,N_19889,N_19870);
and UO_1986 (O_1986,N_19943,N_19830);
nand UO_1987 (O_1987,N_19914,N_19857);
nand UO_1988 (O_1988,N_19831,N_19947);
nand UO_1989 (O_1989,N_19882,N_19822);
and UO_1990 (O_1990,N_19950,N_19944);
and UO_1991 (O_1991,N_19994,N_19803);
nor UO_1992 (O_1992,N_19920,N_19937);
nand UO_1993 (O_1993,N_19930,N_19993);
and UO_1994 (O_1994,N_19922,N_19840);
or UO_1995 (O_1995,N_19937,N_19805);
nor UO_1996 (O_1996,N_19979,N_19888);
or UO_1997 (O_1997,N_19985,N_19946);
nand UO_1998 (O_1998,N_19846,N_19996);
or UO_1999 (O_1999,N_19842,N_19968);
and UO_2000 (O_2000,N_19926,N_19800);
and UO_2001 (O_2001,N_19984,N_19996);
nor UO_2002 (O_2002,N_19887,N_19856);
nor UO_2003 (O_2003,N_19840,N_19994);
and UO_2004 (O_2004,N_19947,N_19859);
or UO_2005 (O_2005,N_19923,N_19852);
nand UO_2006 (O_2006,N_19975,N_19868);
and UO_2007 (O_2007,N_19986,N_19979);
nor UO_2008 (O_2008,N_19899,N_19852);
and UO_2009 (O_2009,N_19825,N_19960);
xnor UO_2010 (O_2010,N_19848,N_19911);
or UO_2011 (O_2011,N_19916,N_19827);
nor UO_2012 (O_2012,N_19987,N_19868);
nand UO_2013 (O_2013,N_19888,N_19863);
nand UO_2014 (O_2014,N_19859,N_19998);
or UO_2015 (O_2015,N_19877,N_19938);
or UO_2016 (O_2016,N_19856,N_19863);
and UO_2017 (O_2017,N_19919,N_19946);
or UO_2018 (O_2018,N_19935,N_19952);
or UO_2019 (O_2019,N_19940,N_19905);
and UO_2020 (O_2020,N_19942,N_19912);
or UO_2021 (O_2021,N_19987,N_19835);
and UO_2022 (O_2022,N_19947,N_19809);
or UO_2023 (O_2023,N_19981,N_19965);
or UO_2024 (O_2024,N_19831,N_19847);
nor UO_2025 (O_2025,N_19963,N_19818);
xnor UO_2026 (O_2026,N_19803,N_19840);
or UO_2027 (O_2027,N_19959,N_19998);
and UO_2028 (O_2028,N_19932,N_19907);
nand UO_2029 (O_2029,N_19807,N_19979);
nand UO_2030 (O_2030,N_19973,N_19914);
nor UO_2031 (O_2031,N_19933,N_19997);
nor UO_2032 (O_2032,N_19977,N_19822);
nor UO_2033 (O_2033,N_19992,N_19812);
or UO_2034 (O_2034,N_19859,N_19927);
and UO_2035 (O_2035,N_19988,N_19928);
or UO_2036 (O_2036,N_19873,N_19810);
and UO_2037 (O_2037,N_19972,N_19917);
nand UO_2038 (O_2038,N_19832,N_19959);
and UO_2039 (O_2039,N_19992,N_19912);
and UO_2040 (O_2040,N_19850,N_19991);
and UO_2041 (O_2041,N_19805,N_19818);
nor UO_2042 (O_2042,N_19964,N_19880);
nand UO_2043 (O_2043,N_19853,N_19867);
nand UO_2044 (O_2044,N_19889,N_19930);
nand UO_2045 (O_2045,N_19836,N_19859);
or UO_2046 (O_2046,N_19882,N_19905);
nor UO_2047 (O_2047,N_19885,N_19944);
or UO_2048 (O_2048,N_19989,N_19957);
or UO_2049 (O_2049,N_19944,N_19901);
or UO_2050 (O_2050,N_19927,N_19807);
or UO_2051 (O_2051,N_19904,N_19847);
and UO_2052 (O_2052,N_19984,N_19964);
and UO_2053 (O_2053,N_19808,N_19883);
nand UO_2054 (O_2054,N_19904,N_19909);
and UO_2055 (O_2055,N_19990,N_19804);
or UO_2056 (O_2056,N_19876,N_19842);
or UO_2057 (O_2057,N_19937,N_19861);
nor UO_2058 (O_2058,N_19929,N_19853);
or UO_2059 (O_2059,N_19900,N_19870);
nand UO_2060 (O_2060,N_19871,N_19863);
nor UO_2061 (O_2061,N_19814,N_19800);
and UO_2062 (O_2062,N_19800,N_19812);
and UO_2063 (O_2063,N_19877,N_19927);
nand UO_2064 (O_2064,N_19907,N_19976);
nand UO_2065 (O_2065,N_19815,N_19920);
nand UO_2066 (O_2066,N_19859,N_19876);
nor UO_2067 (O_2067,N_19982,N_19927);
or UO_2068 (O_2068,N_19911,N_19899);
nor UO_2069 (O_2069,N_19932,N_19812);
and UO_2070 (O_2070,N_19933,N_19943);
and UO_2071 (O_2071,N_19881,N_19880);
nand UO_2072 (O_2072,N_19906,N_19888);
nor UO_2073 (O_2073,N_19869,N_19812);
nand UO_2074 (O_2074,N_19990,N_19879);
and UO_2075 (O_2075,N_19894,N_19888);
nand UO_2076 (O_2076,N_19895,N_19907);
or UO_2077 (O_2077,N_19841,N_19858);
nand UO_2078 (O_2078,N_19883,N_19878);
nand UO_2079 (O_2079,N_19822,N_19998);
or UO_2080 (O_2080,N_19927,N_19874);
and UO_2081 (O_2081,N_19831,N_19913);
and UO_2082 (O_2082,N_19864,N_19988);
nand UO_2083 (O_2083,N_19842,N_19937);
and UO_2084 (O_2084,N_19822,N_19932);
nand UO_2085 (O_2085,N_19991,N_19904);
nand UO_2086 (O_2086,N_19973,N_19951);
nand UO_2087 (O_2087,N_19876,N_19832);
nor UO_2088 (O_2088,N_19860,N_19977);
or UO_2089 (O_2089,N_19983,N_19959);
or UO_2090 (O_2090,N_19930,N_19983);
nand UO_2091 (O_2091,N_19959,N_19871);
and UO_2092 (O_2092,N_19944,N_19908);
and UO_2093 (O_2093,N_19943,N_19842);
or UO_2094 (O_2094,N_19856,N_19803);
and UO_2095 (O_2095,N_19963,N_19841);
or UO_2096 (O_2096,N_19828,N_19957);
nor UO_2097 (O_2097,N_19936,N_19959);
nand UO_2098 (O_2098,N_19975,N_19839);
and UO_2099 (O_2099,N_19929,N_19977);
xor UO_2100 (O_2100,N_19913,N_19876);
and UO_2101 (O_2101,N_19989,N_19999);
and UO_2102 (O_2102,N_19943,N_19821);
or UO_2103 (O_2103,N_19890,N_19856);
and UO_2104 (O_2104,N_19969,N_19815);
or UO_2105 (O_2105,N_19884,N_19887);
nand UO_2106 (O_2106,N_19929,N_19846);
or UO_2107 (O_2107,N_19838,N_19934);
nand UO_2108 (O_2108,N_19936,N_19966);
nand UO_2109 (O_2109,N_19906,N_19802);
nor UO_2110 (O_2110,N_19985,N_19809);
or UO_2111 (O_2111,N_19835,N_19833);
or UO_2112 (O_2112,N_19995,N_19952);
nand UO_2113 (O_2113,N_19926,N_19834);
nand UO_2114 (O_2114,N_19977,N_19922);
or UO_2115 (O_2115,N_19974,N_19975);
or UO_2116 (O_2116,N_19837,N_19907);
and UO_2117 (O_2117,N_19999,N_19820);
nand UO_2118 (O_2118,N_19971,N_19996);
nor UO_2119 (O_2119,N_19832,N_19879);
nor UO_2120 (O_2120,N_19930,N_19973);
or UO_2121 (O_2121,N_19984,N_19839);
nor UO_2122 (O_2122,N_19850,N_19884);
and UO_2123 (O_2123,N_19804,N_19881);
or UO_2124 (O_2124,N_19967,N_19824);
or UO_2125 (O_2125,N_19929,N_19979);
and UO_2126 (O_2126,N_19866,N_19930);
nand UO_2127 (O_2127,N_19940,N_19847);
nor UO_2128 (O_2128,N_19940,N_19841);
nand UO_2129 (O_2129,N_19887,N_19922);
nor UO_2130 (O_2130,N_19878,N_19943);
or UO_2131 (O_2131,N_19876,N_19907);
nor UO_2132 (O_2132,N_19802,N_19862);
nor UO_2133 (O_2133,N_19872,N_19954);
and UO_2134 (O_2134,N_19867,N_19961);
and UO_2135 (O_2135,N_19898,N_19927);
nand UO_2136 (O_2136,N_19870,N_19922);
nand UO_2137 (O_2137,N_19917,N_19800);
and UO_2138 (O_2138,N_19854,N_19912);
nor UO_2139 (O_2139,N_19900,N_19964);
nor UO_2140 (O_2140,N_19919,N_19976);
nand UO_2141 (O_2141,N_19821,N_19965);
nor UO_2142 (O_2142,N_19999,N_19876);
xor UO_2143 (O_2143,N_19834,N_19841);
and UO_2144 (O_2144,N_19964,N_19858);
or UO_2145 (O_2145,N_19905,N_19987);
nor UO_2146 (O_2146,N_19920,N_19932);
nor UO_2147 (O_2147,N_19840,N_19969);
or UO_2148 (O_2148,N_19809,N_19957);
and UO_2149 (O_2149,N_19988,N_19800);
or UO_2150 (O_2150,N_19933,N_19950);
and UO_2151 (O_2151,N_19924,N_19822);
or UO_2152 (O_2152,N_19881,N_19839);
nand UO_2153 (O_2153,N_19843,N_19828);
or UO_2154 (O_2154,N_19935,N_19808);
or UO_2155 (O_2155,N_19826,N_19972);
or UO_2156 (O_2156,N_19873,N_19881);
or UO_2157 (O_2157,N_19892,N_19933);
and UO_2158 (O_2158,N_19894,N_19987);
nor UO_2159 (O_2159,N_19941,N_19934);
nand UO_2160 (O_2160,N_19916,N_19857);
or UO_2161 (O_2161,N_19827,N_19805);
or UO_2162 (O_2162,N_19958,N_19990);
nand UO_2163 (O_2163,N_19912,N_19998);
nor UO_2164 (O_2164,N_19911,N_19988);
and UO_2165 (O_2165,N_19839,N_19950);
nor UO_2166 (O_2166,N_19833,N_19895);
or UO_2167 (O_2167,N_19805,N_19841);
or UO_2168 (O_2168,N_19952,N_19844);
and UO_2169 (O_2169,N_19962,N_19893);
or UO_2170 (O_2170,N_19965,N_19855);
nand UO_2171 (O_2171,N_19852,N_19838);
or UO_2172 (O_2172,N_19953,N_19986);
and UO_2173 (O_2173,N_19992,N_19815);
nand UO_2174 (O_2174,N_19916,N_19812);
nor UO_2175 (O_2175,N_19904,N_19945);
or UO_2176 (O_2176,N_19988,N_19949);
nor UO_2177 (O_2177,N_19883,N_19905);
and UO_2178 (O_2178,N_19905,N_19999);
nand UO_2179 (O_2179,N_19978,N_19942);
and UO_2180 (O_2180,N_19842,N_19913);
nor UO_2181 (O_2181,N_19895,N_19823);
and UO_2182 (O_2182,N_19974,N_19988);
nor UO_2183 (O_2183,N_19919,N_19850);
nand UO_2184 (O_2184,N_19973,N_19896);
nor UO_2185 (O_2185,N_19891,N_19989);
or UO_2186 (O_2186,N_19933,N_19856);
nand UO_2187 (O_2187,N_19963,N_19977);
and UO_2188 (O_2188,N_19851,N_19806);
nand UO_2189 (O_2189,N_19836,N_19810);
nor UO_2190 (O_2190,N_19912,N_19821);
nand UO_2191 (O_2191,N_19809,N_19869);
nand UO_2192 (O_2192,N_19809,N_19865);
nand UO_2193 (O_2193,N_19904,N_19910);
and UO_2194 (O_2194,N_19937,N_19850);
or UO_2195 (O_2195,N_19804,N_19994);
nand UO_2196 (O_2196,N_19909,N_19965);
and UO_2197 (O_2197,N_19861,N_19996);
nand UO_2198 (O_2198,N_19815,N_19935);
nand UO_2199 (O_2199,N_19814,N_19959);
nor UO_2200 (O_2200,N_19890,N_19983);
nor UO_2201 (O_2201,N_19865,N_19918);
or UO_2202 (O_2202,N_19970,N_19811);
or UO_2203 (O_2203,N_19917,N_19889);
and UO_2204 (O_2204,N_19801,N_19812);
nor UO_2205 (O_2205,N_19861,N_19935);
nand UO_2206 (O_2206,N_19889,N_19995);
nand UO_2207 (O_2207,N_19894,N_19870);
or UO_2208 (O_2208,N_19849,N_19898);
or UO_2209 (O_2209,N_19944,N_19851);
nor UO_2210 (O_2210,N_19995,N_19909);
nor UO_2211 (O_2211,N_19894,N_19824);
nand UO_2212 (O_2212,N_19822,N_19872);
and UO_2213 (O_2213,N_19964,N_19967);
or UO_2214 (O_2214,N_19904,N_19857);
or UO_2215 (O_2215,N_19804,N_19980);
nor UO_2216 (O_2216,N_19889,N_19946);
and UO_2217 (O_2217,N_19906,N_19973);
and UO_2218 (O_2218,N_19900,N_19949);
nor UO_2219 (O_2219,N_19823,N_19865);
nand UO_2220 (O_2220,N_19919,N_19837);
or UO_2221 (O_2221,N_19979,N_19998);
or UO_2222 (O_2222,N_19838,N_19908);
nor UO_2223 (O_2223,N_19843,N_19854);
nand UO_2224 (O_2224,N_19931,N_19947);
nor UO_2225 (O_2225,N_19826,N_19903);
nand UO_2226 (O_2226,N_19825,N_19907);
and UO_2227 (O_2227,N_19941,N_19951);
nor UO_2228 (O_2228,N_19838,N_19949);
nand UO_2229 (O_2229,N_19984,N_19817);
nand UO_2230 (O_2230,N_19866,N_19945);
nand UO_2231 (O_2231,N_19965,N_19946);
or UO_2232 (O_2232,N_19865,N_19917);
nand UO_2233 (O_2233,N_19897,N_19952);
or UO_2234 (O_2234,N_19923,N_19949);
nand UO_2235 (O_2235,N_19915,N_19825);
nor UO_2236 (O_2236,N_19959,N_19941);
and UO_2237 (O_2237,N_19829,N_19835);
nor UO_2238 (O_2238,N_19842,N_19907);
and UO_2239 (O_2239,N_19801,N_19839);
nor UO_2240 (O_2240,N_19985,N_19894);
nor UO_2241 (O_2241,N_19846,N_19957);
nor UO_2242 (O_2242,N_19939,N_19901);
and UO_2243 (O_2243,N_19918,N_19841);
or UO_2244 (O_2244,N_19814,N_19853);
or UO_2245 (O_2245,N_19916,N_19977);
nor UO_2246 (O_2246,N_19858,N_19943);
and UO_2247 (O_2247,N_19879,N_19977);
and UO_2248 (O_2248,N_19831,N_19920);
nand UO_2249 (O_2249,N_19940,N_19980);
nor UO_2250 (O_2250,N_19880,N_19928);
nand UO_2251 (O_2251,N_19940,N_19960);
nand UO_2252 (O_2252,N_19928,N_19852);
or UO_2253 (O_2253,N_19912,N_19915);
nand UO_2254 (O_2254,N_19829,N_19996);
nand UO_2255 (O_2255,N_19809,N_19831);
nand UO_2256 (O_2256,N_19981,N_19865);
or UO_2257 (O_2257,N_19952,N_19969);
nand UO_2258 (O_2258,N_19928,N_19995);
and UO_2259 (O_2259,N_19871,N_19817);
nor UO_2260 (O_2260,N_19811,N_19893);
or UO_2261 (O_2261,N_19854,N_19880);
nand UO_2262 (O_2262,N_19929,N_19870);
nand UO_2263 (O_2263,N_19959,N_19843);
and UO_2264 (O_2264,N_19924,N_19929);
nand UO_2265 (O_2265,N_19800,N_19961);
and UO_2266 (O_2266,N_19975,N_19897);
and UO_2267 (O_2267,N_19958,N_19901);
xor UO_2268 (O_2268,N_19821,N_19913);
nand UO_2269 (O_2269,N_19945,N_19899);
nand UO_2270 (O_2270,N_19888,N_19877);
and UO_2271 (O_2271,N_19883,N_19922);
nor UO_2272 (O_2272,N_19900,N_19943);
nor UO_2273 (O_2273,N_19857,N_19883);
nor UO_2274 (O_2274,N_19990,N_19840);
nand UO_2275 (O_2275,N_19879,N_19974);
nand UO_2276 (O_2276,N_19881,N_19955);
or UO_2277 (O_2277,N_19815,N_19901);
or UO_2278 (O_2278,N_19893,N_19996);
or UO_2279 (O_2279,N_19874,N_19861);
or UO_2280 (O_2280,N_19925,N_19858);
and UO_2281 (O_2281,N_19846,N_19870);
nor UO_2282 (O_2282,N_19925,N_19918);
or UO_2283 (O_2283,N_19880,N_19925);
nor UO_2284 (O_2284,N_19961,N_19985);
nand UO_2285 (O_2285,N_19803,N_19975);
nor UO_2286 (O_2286,N_19885,N_19892);
or UO_2287 (O_2287,N_19952,N_19999);
nor UO_2288 (O_2288,N_19843,N_19820);
nor UO_2289 (O_2289,N_19858,N_19918);
nand UO_2290 (O_2290,N_19832,N_19818);
nand UO_2291 (O_2291,N_19850,N_19895);
or UO_2292 (O_2292,N_19949,N_19889);
or UO_2293 (O_2293,N_19958,N_19893);
or UO_2294 (O_2294,N_19822,N_19952);
nand UO_2295 (O_2295,N_19936,N_19877);
nand UO_2296 (O_2296,N_19867,N_19962);
nor UO_2297 (O_2297,N_19867,N_19959);
and UO_2298 (O_2298,N_19970,N_19964);
and UO_2299 (O_2299,N_19967,N_19974);
and UO_2300 (O_2300,N_19900,N_19973);
nand UO_2301 (O_2301,N_19972,N_19987);
and UO_2302 (O_2302,N_19906,N_19946);
or UO_2303 (O_2303,N_19911,N_19823);
nand UO_2304 (O_2304,N_19855,N_19937);
or UO_2305 (O_2305,N_19874,N_19935);
or UO_2306 (O_2306,N_19806,N_19913);
nand UO_2307 (O_2307,N_19883,N_19935);
nand UO_2308 (O_2308,N_19891,N_19897);
nand UO_2309 (O_2309,N_19997,N_19912);
and UO_2310 (O_2310,N_19927,N_19887);
nand UO_2311 (O_2311,N_19858,N_19842);
nor UO_2312 (O_2312,N_19979,N_19930);
nand UO_2313 (O_2313,N_19877,N_19800);
or UO_2314 (O_2314,N_19864,N_19856);
or UO_2315 (O_2315,N_19965,N_19958);
or UO_2316 (O_2316,N_19900,N_19967);
nand UO_2317 (O_2317,N_19836,N_19841);
and UO_2318 (O_2318,N_19942,N_19867);
nor UO_2319 (O_2319,N_19937,N_19847);
xnor UO_2320 (O_2320,N_19876,N_19946);
nor UO_2321 (O_2321,N_19852,N_19826);
or UO_2322 (O_2322,N_19927,N_19909);
nor UO_2323 (O_2323,N_19843,N_19864);
and UO_2324 (O_2324,N_19977,N_19974);
and UO_2325 (O_2325,N_19949,N_19908);
and UO_2326 (O_2326,N_19854,N_19895);
or UO_2327 (O_2327,N_19952,N_19929);
nand UO_2328 (O_2328,N_19933,N_19850);
nor UO_2329 (O_2329,N_19922,N_19802);
nor UO_2330 (O_2330,N_19813,N_19990);
nor UO_2331 (O_2331,N_19892,N_19807);
and UO_2332 (O_2332,N_19848,N_19929);
and UO_2333 (O_2333,N_19888,N_19968);
nor UO_2334 (O_2334,N_19944,N_19899);
and UO_2335 (O_2335,N_19988,N_19926);
nand UO_2336 (O_2336,N_19806,N_19938);
or UO_2337 (O_2337,N_19848,N_19851);
and UO_2338 (O_2338,N_19960,N_19944);
nand UO_2339 (O_2339,N_19869,N_19956);
nand UO_2340 (O_2340,N_19855,N_19881);
or UO_2341 (O_2341,N_19928,N_19860);
and UO_2342 (O_2342,N_19891,N_19843);
nand UO_2343 (O_2343,N_19832,N_19922);
or UO_2344 (O_2344,N_19859,N_19874);
or UO_2345 (O_2345,N_19849,N_19951);
nand UO_2346 (O_2346,N_19902,N_19940);
xnor UO_2347 (O_2347,N_19839,N_19883);
nand UO_2348 (O_2348,N_19938,N_19845);
or UO_2349 (O_2349,N_19919,N_19855);
nand UO_2350 (O_2350,N_19961,N_19857);
and UO_2351 (O_2351,N_19971,N_19964);
xnor UO_2352 (O_2352,N_19952,N_19927);
or UO_2353 (O_2353,N_19864,N_19865);
or UO_2354 (O_2354,N_19915,N_19857);
xor UO_2355 (O_2355,N_19948,N_19844);
and UO_2356 (O_2356,N_19832,N_19821);
xor UO_2357 (O_2357,N_19952,N_19883);
nor UO_2358 (O_2358,N_19877,N_19836);
or UO_2359 (O_2359,N_19849,N_19921);
and UO_2360 (O_2360,N_19866,N_19815);
nor UO_2361 (O_2361,N_19998,N_19970);
xnor UO_2362 (O_2362,N_19872,N_19875);
or UO_2363 (O_2363,N_19940,N_19854);
and UO_2364 (O_2364,N_19829,N_19941);
nand UO_2365 (O_2365,N_19892,N_19822);
and UO_2366 (O_2366,N_19928,N_19948);
and UO_2367 (O_2367,N_19884,N_19804);
nand UO_2368 (O_2368,N_19952,N_19855);
nor UO_2369 (O_2369,N_19829,N_19886);
nor UO_2370 (O_2370,N_19952,N_19899);
nand UO_2371 (O_2371,N_19889,N_19939);
or UO_2372 (O_2372,N_19864,N_19899);
xnor UO_2373 (O_2373,N_19912,N_19879);
and UO_2374 (O_2374,N_19935,N_19827);
nor UO_2375 (O_2375,N_19992,N_19884);
nand UO_2376 (O_2376,N_19863,N_19838);
nor UO_2377 (O_2377,N_19902,N_19842);
and UO_2378 (O_2378,N_19887,N_19917);
nor UO_2379 (O_2379,N_19924,N_19930);
nor UO_2380 (O_2380,N_19906,N_19847);
nor UO_2381 (O_2381,N_19896,N_19898);
or UO_2382 (O_2382,N_19834,N_19931);
nand UO_2383 (O_2383,N_19911,N_19835);
or UO_2384 (O_2384,N_19989,N_19926);
xnor UO_2385 (O_2385,N_19919,N_19807);
and UO_2386 (O_2386,N_19964,N_19864);
nand UO_2387 (O_2387,N_19952,N_19847);
nand UO_2388 (O_2388,N_19902,N_19946);
and UO_2389 (O_2389,N_19949,N_19912);
nor UO_2390 (O_2390,N_19817,N_19841);
nor UO_2391 (O_2391,N_19888,N_19857);
nor UO_2392 (O_2392,N_19950,N_19991);
nor UO_2393 (O_2393,N_19874,N_19846);
nand UO_2394 (O_2394,N_19859,N_19972);
nand UO_2395 (O_2395,N_19958,N_19890);
or UO_2396 (O_2396,N_19955,N_19908);
or UO_2397 (O_2397,N_19924,N_19977);
nand UO_2398 (O_2398,N_19850,N_19926);
and UO_2399 (O_2399,N_19839,N_19844);
or UO_2400 (O_2400,N_19842,N_19939);
and UO_2401 (O_2401,N_19866,N_19885);
and UO_2402 (O_2402,N_19943,N_19974);
and UO_2403 (O_2403,N_19851,N_19969);
nor UO_2404 (O_2404,N_19935,N_19833);
nand UO_2405 (O_2405,N_19813,N_19819);
nand UO_2406 (O_2406,N_19986,N_19915);
nor UO_2407 (O_2407,N_19929,N_19990);
and UO_2408 (O_2408,N_19914,N_19924);
or UO_2409 (O_2409,N_19943,N_19945);
nor UO_2410 (O_2410,N_19938,N_19825);
or UO_2411 (O_2411,N_19985,N_19828);
nand UO_2412 (O_2412,N_19860,N_19854);
or UO_2413 (O_2413,N_19990,N_19959);
nor UO_2414 (O_2414,N_19825,N_19992);
nand UO_2415 (O_2415,N_19857,N_19827);
nand UO_2416 (O_2416,N_19876,N_19924);
nand UO_2417 (O_2417,N_19935,N_19811);
and UO_2418 (O_2418,N_19962,N_19958);
nand UO_2419 (O_2419,N_19902,N_19802);
or UO_2420 (O_2420,N_19879,N_19914);
nor UO_2421 (O_2421,N_19901,N_19884);
or UO_2422 (O_2422,N_19915,N_19979);
or UO_2423 (O_2423,N_19949,N_19901);
or UO_2424 (O_2424,N_19811,N_19887);
and UO_2425 (O_2425,N_19916,N_19861);
nand UO_2426 (O_2426,N_19928,N_19986);
or UO_2427 (O_2427,N_19952,N_19986);
or UO_2428 (O_2428,N_19902,N_19888);
and UO_2429 (O_2429,N_19972,N_19960);
nand UO_2430 (O_2430,N_19956,N_19870);
nand UO_2431 (O_2431,N_19976,N_19903);
nor UO_2432 (O_2432,N_19912,N_19885);
or UO_2433 (O_2433,N_19864,N_19854);
nand UO_2434 (O_2434,N_19837,N_19964);
nor UO_2435 (O_2435,N_19999,N_19846);
and UO_2436 (O_2436,N_19833,N_19866);
and UO_2437 (O_2437,N_19938,N_19904);
or UO_2438 (O_2438,N_19985,N_19801);
nor UO_2439 (O_2439,N_19835,N_19891);
or UO_2440 (O_2440,N_19891,N_19937);
or UO_2441 (O_2441,N_19815,N_19859);
nand UO_2442 (O_2442,N_19910,N_19961);
and UO_2443 (O_2443,N_19867,N_19938);
xor UO_2444 (O_2444,N_19857,N_19990);
nor UO_2445 (O_2445,N_19866,N_19816);
nor UO_2446 (O_2446,N_19893,N_19863);
nor UO_2447 (O_2447,N_19829,N_19934);
and UO_2448 (O_2448,N_19891,N_19929);
nor UO_2449 (O_2449,N_19857,N_19811);
and UO_2450 (O_2450,N_19951,N_19851);
nand UO_2451 (O_2451,N_19957,N_19849);
or UO_2452 (O_2452,N_19933,N_19857);
nand UO_2453 (O_2453,N_19976,N_19874);
nand UO_2454 (O_2454,N_19925,N_19992);
xor UO_2455 (O_2455,N_19866,N_19867);
and UO_2456 (O_2456,N_19963,N_19996);
nor UO_2457 (O_2457,N_19901,N_19858);
or UO_2458 (O_2458,N_19909,N_19891);
nor UO_2459 (O_2459,N_19875,N_19949);
nor UO_2460 (O_2460,N_19893,N_19817);
and UO_2461 (O_2461,N_19985,N_19833);
and UO_2462 (O_2462,N_19838,N_19944);
nand UO_2463 (O_2463,N_19902,N_19862);
nand UO_2464 (O_2464,N_19898,N_19907);
nand UO_2465 (O_2465,N_19811,N_19802);
and UO_2466 (O_2466,N_19827,N_19850);
or UO_2467 (O_2467,N_19960,N_19895);
or UO_2468 (O_2468,N_19972,N_19820);
nor UO_2469 (O_2469,N_19813,N_19981);
or UO_2470 (O_2470,N_19999,N_19854);
nand UO_2471 (O_2471,N_19955,N_19943);
or UO_2472 (O_2472,N_19842,N_19988);
and UO_2473 (O_2473,N_19862,N_19892);
or UO_2474 (O_2474,N_19987,N_19920);
and UO_2475 (O_2475,N_19985,N_19983);
and UO_2476 (O_2476,N_19931,N_19859);
and UO_2477 (O_2477,N_19857,N_19836);
nand UO_2478 (O_2478,N_19810,N_19816);
or UO_2479 (O_2479,N_19810,N_19837);
or UO_2480 (O_2480,N_19816,N_19935);
nand UO_2481 (O_2481,N_19891,N_19926);
or UO_2482 (O_2482,N_19906,N_19877);
xor UO_2483 (O_2483,N_19919,N_19966);
and UO_2484 (O_2484,N_19990,N_19902);
nand UO_2485 (O_2485,N_19856,N_19935);
nand UO_2486 (O_2486,N_19811,N_19980);
nand UO_2487 (O_2487,N_19851,N_19917);
or UO_2488 (O_2488,N_19910,N_19899);
and UO_2489 (O_2489,N_19882,N_19945);
nand UO_2490 (O_2490,N_19988,N_19901);
xnor UO_2491 (O_2491,N_19825,N_19883);
nand UO_2492 (O_2492,N_19990,N_19881);
and UO_2493 (O_2493,N_19855,N_19816);
xor UO_2494 (O_2494,N_19951,N_19976);
and UO_2495 (O_2495,N_19868,N_19831);
and UO_2496 (O_2496,N_19801,N_19842);
and UO_2497 (O_2497,N_19884,N_19895);
or UO_2498 (O_2498,N_19902,N_19917);
nand UO_2499 (O_2499,N_19887,N_19847);
endmodule