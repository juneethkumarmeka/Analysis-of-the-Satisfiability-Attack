module basic_2500_25000_3000_8_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nand U0 (N_0,In_408,In_242);
nor U1 (N_1,In_1765,In_2439);
and U2 (N_2,In_914,In_1824);
nor U3 (N_3,In_351,In_2417);
or U4 (N_4,In_1530,In_2496);
nor U5 (N_5,In_540,In_1093);
and U6 (N_6,In_1827,In_101);
and U7 (N_7,In_500,In_485);
nand U8 (N_8,In_1621,In_2307);
xor U9 (N_9,In_694,In_173);
or U10 (N_10,In_894,In_2244);
or U11 (N_11,In_289,In_1032);
nor U12 (N_12,In_1430,In_72);
and U13 (N_13,In_737,In_1089);
or U14 (N_14,In_1578,In_565);
or U15 (N_15,In_138,In_2116);
and U16 (N_16,In_768,In_1076);
xor U17 (N_17,In_2453,In_1100);
and U18 (N_18,In_2077,In_1444);
xnor U19 (N_19,In_469,In_1091);
and U20 (N_20,In_1067,In_559);
and U21 (N_21,In_499,In_1731);
nor U22 (N_22,In_1106,In_786);
nand U23 (N_23,In_1348,In_1748);
or U24 (N_24,In_2029,In_1445);
or U25 (N_25,In_573,In_2100);
or U26 (N_26,In_2205,In_470);
or U27 (N_27,In_477,In_1454);
nand U28 (N_28,In_846,In_794);
or U29 (N_29,In_1528,In_1634);
nand U30 (N_30,In_2112,In_531);
and U31 (N_31,In_2451,In_1836);
or U32 (N_32,In_613,In_1154);
nand U33 (N_33,In_797,In_1262);
and U34 (N_34,In_576,In_2023);
and U35 (N_35,In_1047,In_161);
and U36 (N_36,In_2384,In_1215);
nor U37 (N_37,In_2234,In_2061);
and U38 (N_38,In_1995,In_1819);
and U39 (N_39,In_1838,In_1708);
nand U40 (N_40,In_281,In_1096);
nand U41 (N_41,In_2273,In_1338);
or U42 (N_42,In_986,In_980);
or U43 (N_43,In_287,In_2144);
or U44 (N_44,In_644,In_639);
or U45 (N_45,In_856,In_1685);
nand U46 (N_46,In_2041,In_1479);
or U47 (N_47,In_396,In_537);
nor U48 (N_48,In_1974,In_2348);
nand U49 (N_49,In_54,In_444);
nand U50 (N_50,In_896,In_89);
or U51 (N_51,In_1048,In_409);
and U52 (N_52,In_2175,In_325);
or U53 (N_53,In_2305,In_736);
and U54 (N_54,In_988,In_2036);
or U55 (N_55,In_2193,In_1144);
nand U56 (N_56,In_2267,In_216);
nor U57 (N_57,In_144,In_1107);
or U58 (N_58,In_1160,In_1341);
or U59 (N_59,In_215,In_458);
xnor U60 (N_60,In_1113,In_1894);
and U61 (N_61,In_1226,In_827);
nand U62 (N_62,In_557,In_2182);
and U63 (N_63,In_2055,In_1441);
and U64 (N_64,In_2458,In_526);
and U65 (N_65,In_1651,In_81);
nor U66 (N_66,In_1388,In_2468);
xor U67 (N_67,In_640,In_1551);
and U68 (N_68,In_804,In_1169);
nor U69 (N_69,In_624,In_1428);
nand U70 (N_70,In_1461,In_1527);
nand U71 (N_71,In_1500,In_1079);
nand U72 (N_72,In_2378,In_508);
nand U73 (N_73,In_232,In_2216);
nand U74 (N_74,In_1652,In_525);
nor U75 (N_75,In_619,In_735);
nor U76 (N_76,In_1072,In_1679);
or U77 (N_77,In_478,In_2038);
and U78 (N_78,In_230,In_1702);
nand U79 (N_79,In_2225,In_2042);
and U80 (N_80,In_2350,In_599);
and U81 (N_81,In_2314,In_1227);
or U82 (N_82,In_2212,In_954);
nor U83 (N_83,In_1565,In_501);
nand U84 (N_84,In_331,In_109);
and U85 (N_85,In_1312,In_1177);
nor U86 (N_86,In_166,In_1778);
nor U87 (N_87,In_1153,In_2110);
nor U88 (N_88,In_1673,In_407);
or U89 (N_89,In_916,In_200);
and U90 (N_90,In_1889,In_1409);
and U91 (N_91,In_104,In_1097);
or U92 (N_92,In_974,In_102);
or U93 (N_93,In_1739,In_2452);
and U94 (N_94,In_1236,In_2475);
or U95 (N_95,In_861,In_299);
and U96 (N_96,In_1640,In_953);
nor U97 (N_97,In_2121,In_669);
nand U98 (N_98,In_872,In_2166);
or U99 (N_99,In_967,In_753);
nor U100 (N_100,In_1482,In_897);
nor U101 (N_101,In_427,In_2429);
and U102 (N_102,In_670,In_1534);
or U103 (N_103,In_1490,In_197);
nand U104 (N_104,In_1537,In_298);
or U105 (N_105,In_1367,In_1768);
and U106 (N_106,In_2007,In_467);
xnor U107 (N_107,In_1234,In_1495);
nor U108 (N_108,In_965,In_15);
xnor U109 (N_109,In_419,In_686);
nand U110 (N_110,In_2471,In_1420);
nor U111 (N_111,In_1466,In_1346);
xnor U112 (N_112,In_1850,In_680);
or U113 (N_113,In_92,In_1059);
nor U114 (N_114,In_491,In_566);
and U115 (N_115,In_609,In_823);
nor U116 (N_116,In_453,In_530);
xor U117 (N_117,In_574,In_1735);
nand U118 (N_118,In_9,In_463);
and U119 (N_119,In_664,In_715);
nor U120 (N_120,In_223,In_103);
and U121 (N_121,In_1951,In_468);
or U122 (N_122,In_1233,In_402);
and U123 (N_123,In_796,In_749);
nand U124 (N_124,In_1460,In_586);
nor U125 (N_125,In_69,In_1309);
and U126 (N_126,In_1925,In_1696);
and U127 (N_127,In_1485,In_940);
and U128 (N_128,In_1992,In_1725);
nor U129 (N_129,In_2329,In_249);
and U130 (N_130,In_1835,In_443);
nor U131 (N_131,In_2047,In_973);
nand U132 (N_132,In_1985,In_51);
and U133 (N_133,In_601,In_1321);
nand U134 (N_134,In_1011,In_1390);
xnor U135 (N_135,In_1684,In_1826);
nand U136 (N_136,In_2472,In_1357);
nand U137 (N_137,In_1639,In_288);
or U138 (N_138,In_21,In_2437);
and U139 (N_139,In_1423,In_2242);
xnor U140 (N_140,In_868,In_1763);
or U141 (N_141,In_1614,In_1128);
nor U142 (N_142,In_693,In_365);
and U143 (N_143,In_1038,In_115);
nand U144 (N_144,In_291,In_1373);
nor U145 (N_145,In_113,In_2300);
or U146 (N_146,In_1549,In_1542);
nand U147 (N_147,In_615,In_1724);
nor U148 (N_148,In_48,In_265);
and U149 (N_149,In_511,In_663);
nor U150 (N_150,In_218,In_1954);
nand U151 (N_151,In_1884,In_927);
or U152 (N_152,In_1174,In_2297);
nand U153 (N_153,In_548,In_1328);
and U154 (N_154,In_1303,In_1413);
or U155 (N_155,In_1241,In_303);
and U156 (N_156,In_2365,In_1976);
xor U157 (N_157,In_2330,In_1396);
nor U158 (N_158,In_522,In_2396);
or U159 (N_159,In_160,In_1298);
or U160 (N_160,In_2174,In_744);
and U161 (N_161,In_2089,In_2251);
nand U162 (N_162,In_44,In_1637);
or U163 (N_163,In_302,In_626);
nor U164 (N_164,In_702,In_1502);
nor U165 (N_165,In_439,In_2333);
and U166 (N_166,In_492,In_2399);
or U167 (N_167,In_1264,In_36);
nand U168 (N_168,In_824,In_898);
xnor U169 (N_169,In_406,In_428);
xnor U170 (N_170,In_2258,In_106);
nor U171 (N_171,In_517,In_139);
xor U172 (N_172,In_1631,In_556);
or U173 (N_173,In_2433,In_2084);
and U174 (N_174,In_1465,In_1507);
xor U175 (N_175,In_1035,In_875);
nand U176 (N_176,In_455,In_1031);
nand U177 (N_177,In_1515,In_1489);
nor U178 (N_178,In_1410,In_1987);
and U179 (N_179,In_2277,In_1650);
and U180 (N_180,In_1676,In_985);
xor U181 (N_181,In_1204,In_539);
nor U182 (N_182,In_1541,In_1592);
and U183 (N_183,In_438,In_1707);
nand U184 (N_184,In_2190,In_78);
or U185 (N_185,In_1111,In_2264);
or U186 (N_186,In_755,In_1936);
nand U187 (N_187,In_2315,In_486);
or U188 (N_188,In_2480,In_1082);
nand U189 (N_189,In_641,In_2156);
and U190 (N_190,In_1643,In_1845);
xor U191 (N_191,In_905,In_546);
or U192 (N_192,In_2178,In_1400);
nor U193 (N_193,In_231,In_1314);
nand U194 (N_194,In_1133,In_2195);
or U195 (N_195,In_2400,In_1855);
and U196 (N_196,In_589,In_1921);
or U197 (N_197,In_497,In_143);
nand U198 (N_198,In_2105,In_2133);
and U199 (N_199,In_1155,In_1857);
nor U200 (N_200,In_826,In_1480);
nor U201 (N_201,In_1586,In_535);
nor U202 (N_202,In_1315,In_2176);
or U203 (N_203,In_1284,In_2370);
nand U204 (N_204,In_675,In_398);
nand U205 (N_205,In_1045,In_1810);
xnor U206 (N_206,In_659,In_5);
xor U207 (N_207,In_1131,In_1316);
nor U208 (N_208,In_229,In_1398);
nand U209 (N_209,In_2372,In_2293);
xor U210 (N_210,In_123,In_2421);
nor U211 (N_211,In_1546,In_1605);
nor U212 (N_212,In_1268,In_1102);
xnor U213 (N_213,In_1783,In_812);
and U214 (N_214,In_1170,In_1232);
nor U215 (N_215,In_2463,In_1548);
or U216 (N_216,In_2076,In_2034);
nor U217 (N_217,In_1034,In_2292);
nand U218 (N_218,In_1692,In_2303);
and U219 (N_219,In_1190,In_2422);
and U220 (N_220,In_668,In_93);
or U221 (N_221,In_2002,In_2210);
nand U222 (N_222,In_2013,In_1447);
or U223 (N_223,In_1254,In_2331);
nor U224 (N_224,In_1820,In_364);
nor U225 (N_225,In_1167,In_1501);
and U226 (N_226,In_1422,In_235);
nor U227 (N_227,In_2196,In_1833);
or U228 (N_228,In_2252,In_1435);
or U229 (N_229,In_1335,In_278);
nor U230 (N_230,In_2153,In_2294);
nor U231 (N_231,In_476,In_1095);
nand U232 (N_232,In_1116,In_2169);
and U233 (N_233,In_2493,In_1667);
or U234 (N_234,In_814,In_1825);
xor U235 (N_235,In_667,In_527);
xnor U236 (N_236,In_1112,In_528);
nand U237 (N_237,In_867,In_1164);
nor U238 (N_238,In_2498,In_1520);
or U239 (N_239,In_612,In_938);
xor U240 (N_240,In_1701,In_2265);
nand U241 (N_241,In_295,In_1218);
and U242 (N_242,In_1257,In_579);
or U243 (N_243,In_400,In_1516);
nor U244 (N_244,In_1814,In_2270);
or U245 (N_245,In_401,In_1004);
or U246 (N_246,In_750,In_130);
nand U247 (N_247,In_1970,In_1275);
and U248 (N_248,In_1881,In_2164);
or U249 (N_249,In_2402,In_1389);
nor U250 (N_250,In_809,In_859);
nand U251 (N_251,In_1939,In_100);
or U252 (N_252,In_1104,In_1785);
and U253 (N_253,In_328,In_1442);
and U254 (N_254,In_136,In_2483);
xnor U255 (N_255,In_1929,In_1121);
and U256 (N_256,In_2332,In_801);
xnor U257 (N_257,In_97,In_789);
nor U258 (N_258,In_2407,In_1406);
or U259 (N_259,In_730,In_2389);
or U260 (N_260,In_1455,In_213);
nand U261 (N_261,In_2342,In_881);
xor U262 (N_262,In_684,In_181);
and U263 (N_263,In_820,In_704);
and U264 (N_264,In_1469,In_892);
nor U265 (N_265,In_2403,In_1755);
and U266 (N_266,In_2319,In_1784);
or U267 (N_267,In_1386,In_627);
and U268 (N_268,In_1296,In_55);
nor U269 (N_269,In_588,In_284);
or U270 (N_270,In_1536,In_2306);
or U271 (N_271,In_395,In_979);
xnor U272 (N_272,In_251,In_1687);
nor U273 (N_273,In_2425,In_2096);
nand U274 (N_274,In_1581,In_2302);
or U275 (N_275,In_2397,In_1867);
nor U276 (N_276,In_2441,In_2470);
or U277 (N_277,In_884,In_1364);
and U278 (N_278,In_777,In_1737);
and U279 (N_279,In_696,In_441);
or U280 (N_280,In_214,In_332);
nor U281 (N_281,In_310,In_2494);
or U282 (N_282,In_1677,In_1437);
nor U283 (N_283,In_902,In_2159);
nor U284 (N_284,In_203,In_1187);
or U285 (N_285,In_2367,In_2461);
nand U286 (N_286,In_2206,In_177);
or U287 (N_287,In_555,In_785);
nand U288 (N_288,In_1329,In_729);
nand U289 (N_289,In_16,In_1418);
or U290 (N_290,In_1175,In_637);
nand U291 (N_291,In_1165,In_2401);
xor U292 (N_292,In_918,In_1387);
nand U293 (N_293,In_636,In_87);
or U294 (N_294,In_150,In_1286);
nor U295 (N_295,In_1874,In_1620);
nor U296 (N_296,In_1083,In_417);
nand U297 (N_297,In_2291,In_751);
xnor U298 (N_298,In_2489,In_2394);
and U299 (N_299,In_519,In_320);
and U300 (N_300,In_2262,In_1832);
nand U301 (N_301,In_1271,In_521);
or U302 (N_302,In_1365,In_734);
nor U303 (N_303,In_169,In_152);
nor U304 (N_304,In_264,In_1522);
nand U305 (N_305,In_323,In_1796);
and U306 (N_306,In_268,In_440);
or U307 (N_307,In_1745,In_1007);
xnor U308 (N_308,In_2428,In_1023);
or U309 (N_309,In_1394,In_1941);
or U310 (N_310,In_1998,In_710);
and U311 (N_311,In_2308,In_196);
nand U312 (N_312,In_1024,In_1180);
and U313 (N_313,In_2122,In_1595);
nor U314 (N_314,In_1660,In_1686);
nor U315 (N_315,In_1267,In_356);
nand U316 (N_316,In_2215,In_1744);
or U317 (N_317,In_1790,In_758);
and U318 (N_318,In_1540,In_2448);
and U319 (N_319,In_915,In_941);
xnor U320 (N_320,In_1887,In_1648);
nand U321 (N_321,In_357,In_1355);
xnor U322 (N_322,In_1068,In_1054);
xor U323 (N_323,In_424,In_2028);
nor U324 (N_324,In_314,In_935);
nand U325 (N_325,In_1844,In_776);
nor U326 (N_326,In_1729,In_1963);
nor U327 (N_327,In_962,In_1572);
nand U328 (N_328,In_1179,In_761);
and U329 (N_329,In_1519,In_118);
xnor U330 (N_330,In_77,In_480);
or U331 (N_331,In_1403,In_2261);
xor U332 (N_332,In_813,In_665);
or U333 (N_333,In_1919,In_784);
nor U334 (N_334,In_2341,In_296);
nand U335 (N_335,In_2373,In_2414);
nor U336 (N_336,In_378,In_1957);
or U337 (N_337,In_1608,In_745);
and U338 (N_338,In_841,In_2266);
nand U339 (N_339,In_2135,In_919);
and U340 (N_340,In_975,In_504);
nor U341 (N_341,In_1216,In_273);
and U342 (N_342,In_1671,In_372);
nor U343 (N_343,In_958,In_2086);
nor U344 (N_344,In_413,In_2181);
nor U345 (N_345,In_1788,In_1483);
and U346 (N_346,In_607,In_802);
xnor U347 (N_347,In_198,In_2194);
and U348 (N_348,In_1185,In_193);
or U349 (N_349,In_647,In_2465);
and U350 (N_350,In_1277,In_274);
nor U351 (N_351,In_2046,In_2091);
and U352 (N_352,In_95,In_1659);
xor U353 (N_353,In_1869,In_1554);
nand U354 (N_354,In_790,In_2025);
or U355 (N_355,In_1431,In_1834);
or U356 (N_356,In_1099,In_1901);
nor U357 (N_357,In_1623,In_1973);
xnor U358 (N_358,In_550,In_2413);
or U359 (N_359,In_1775,In_853);
and U360 (N_360,In_2213,In_1205);
nor U361 (N_361,In_1597,In_1883);
and U362 (N_362,In_1734,In_948);
and U363 (N_363,In_538,In_399);
and U364 (N_364,In_805,In_890);
nor U365 (N_365,In_957,In_1663);
and U366 (N_366,In_1473,In_587);
xor U367 (N_367,In_27,In_2039);
nor U368 (N_368,In_250,In_1580);
nand U369 (N_369,In_1764,In_1282);
or U370 (N_370,In_2085,In_1186);
and U371 (N_371,In_2187,In_1641);
or U372 (N_372,In_2426,In_1361);
nor U373 (N_373,In_739,In_909);
nor U374 (N_374,In_1063,In_2104);
nor U375 (N_375,In_1379,In_842);
and U376 (N_376,In_623,In_1847);
nand U377 (N_377,In_561,In_1767);
xnor U378 (N_378,In_1301,In_1203);
nor U379 (N_379,In_2005,In_1959);
nor U380 (N_380,In_932,In_1488);
xnor U381 (N_381,In_552,In_452);
and U382 (N_382,In_2000,In_532);
or U383 (N_383,In_47,In_376);
nand U384 (N_384,In_1664,In_125);
and U385 (N_385,In_2312,In_1900);
and U386 (N_386,In_2481,In_1451);
xnor U387 (N_387,In_2345,In_1449);
xor U388 (N_388,In_2382,In_1782);
nand U389 (N_389,In_1715,In_2211);
or U390 (N_390,In_1560,In_2462);
or U391 (N_391,In_879,In_2068);
nand U392 (N_392,In_863,In_1557);
nand U393 (N_393,In_13,In_280);
and U394 (N_394,In_1757,In_1397);
or U395 (N_395,In_2058,In_1108);
and U396 (N_396,In_1021,In_1349);
and U397 (N_397,In_1304,In_516);
xnor U398 (N_398,In_931,In_2171);
nor U399 (N_399,In_2035,In_2014);
and U400 (N_400,In_543,In_1088);
xor U401 (N_401,In_933,In_1066);
or U402 (N_402,In_1201,In_949);
xor U403 (N_403,In_2201,In_893);
xnor U404 (N_404,In_2044,In_2198);
and U405 (N_405,In_717,In_509);
nand U406 (N_406,In_2405,In_1074);
nor U407 (N_407,In_1084,In_42);
and U408 (N_408,In_20,In_645);
xor U409 (N_409,In_317,In_2486);
nand U410 (N_410,In_269,In_1305);
nor U411 (N_411,In_283,In_1197);
and U412 (N_412,In_819,In_560);
xnor U413 (N_413,In_1851,In_1162);
nand U414 (N_414,In_738,In_2129);
and U415 (N_415,In_506,In_2209);
nor U416 (N_416,In_2119,In_38);
nor U417 (N_417,In_830,In_1665);
or U418 (N_418,In_1436,In_159);
or U419 (N_419,In_2454,In_1274);
and U420 (N_420,In_2098,In_2324);
and U421 (N_421,In_85,In_2063);
xnor U422 (N_422,In_316,In_674);
and U423 (N_423,In_1042,In_1075);
nand U424 (N_424,In_959,In_2376);
and U425 (N_425,In_1086,In_2395);
or U426 (N_426,In_676,In_2418);
xnor U427 (N_427,In_858,In_361);
or U428 (N_428,In_330,In_1142);
nor U429 (N_429,In_1746,In_1117);
or U430 (N_430,In_917,In_989);
or U431 (N_431,In_1794,In_991);
xor U432 (N_432,In_1991,In_436);
nor U433 (N_433,In_83,In_1716);
and U434 (N_434,In_493,In_995);
or U435 (N_435,In_2059,In_34);
or U436 (N_436,In_889,In_825);
and U437 (N_437,In_621,In_1340);
nand U438 (N_438,In_2346,In_425);
or U439 (N_439,In_1459,In_2409);
or U440 (N_440,In_2219,In_1908);
nand U441 (N_441,In_1994,In_544);
xnor U442 (N_442,In_860,In_633);
or U443 (N_443,In_114,In_1616);
nand U444 (N_444,In_192,In_847);
nor U445 (N_445,In_1758,In_35);
xnor U446 (N_446,In_2257,In_791);
or U447 (N_447,In_30,In_1375);
or U448 (N_448,In_1852,In_1585);
or U449 (N_449,In_209,In_558);
xor U450 (N_450,In_10,In_2456);
and U451 (N_451,In_2167,In_585);
or U452 (N_452,In_2377,In_437);
or U453 (N_453,In_134,In_1989);
and U454 (N_454,In_2322,In_2466);
nor U455 (N_455,In_926,In_1292);
nor U456 (N_456,In_2043,In_1661);
nor U457 (N_457,In_1849,In_808);
or U458 (N_458,In_799,In_241);
or U459 (N_459,In_628,In_1094);
nor U460 (N_460,In_2124,In_279);
xor U461 (N_461,In_970,In_141);
and U462 (N_462,In_195,In_1535);
and U463 (N_463,In_2339,In_913);
or U464 (N_464,In_1342,In_1016);
and U465 (N_465,In_1747,In_1324);
or U466 (N_466,In_912,In_1934);
nand U467 (N_467,In_459,In_1051);
nor U468 (N_468,In_1143,In_90);
nor U469 (N_469,In_910,In_224);
and U470 (N_470,In_787,In_1158);
nand U471 (N_471,In_185,In_1478);
and U472 (N_472,In_2298,In_1440);
nor U473 (N_473,In_712,In_1371);
nor U474 (N_474,In_523,In_336);
nor U475 (N_475,In_1087,In_2152);
nor U476 (N_476,In_743,In_1923);
or U477 (N_477,In_2048,In_2391);
nor U478 (N_478,In_1902,In_699);
nand U479 (N_479,In_1750,In_792);
and U480 (N_480,In_1730,In_839);
nor U481 (N_481,In_687,In_1517);
nand U482 (N_482,In_31,In_2488);
nor U483 (N_483,In_1193,In_1049);
nand U484 (N_484,In_259,In_6);
or U485 (N_485,In_2473,In_201);
nand U486 (N_486,In_2021,In_335);
nand U487 (N_487,In_53,In_4);
xor U488 (N_488,In_1967,In_1843);
nor U489 (N_489,In_2081,In_507);
nor U490 (N_490,In_1635,In_1374);
nor U491 (N_491,In_1879,In_2150);
and U492 (N_492,In_2185,In_1253);
nand U493 (N_493,In_204,In_2260);
and U494 (N_494,In_267,In_0);
and U495 (N_495,In_1882,In_1841);
or U496 (N_496,In_1070,In_1446);
and U497 (N_497,In_757,In_2214);
or U498 (N_498,In_1071,In_154);
nand U499 (N_499,In_649,In_1988);
nand U500 (N_500,In_434,In_2485);
or U501 (N_501,In_1911,In_1720);
and U502 (N_502,In_2310,In_1053);
xnor U503 (N_503,In_1242,In_1182);
nand U504 (N_504,In_582,In_2253);
nor U505 (N_505,In_2286,In_2151);
nor U506 (N_506,In_416,In_2388);
nand U507 (N_507,In_260,In_366);
and U508 (N_508,In_404,In_1713);
nand U509 (N_509,In_82,In_176);
nor U510 (N_510,In_968,In_1372);
nor U511 (N_511,In_1424,In_1774);
or U512 (N_512,In_2321,In_2027);
or U513 (N_513,In_1828,In_1858);
xnor U514 (N_514,In_1839,In_170);
nand U515 (N_515,In_1965,In_494);
and U516 (N_516,In_2246,In_1496);
xnor U517 (N_517,In_924,In_904);
nand U518 (N_518,In_844,In_1933);
and U519 (N_519,In_1848,In_671);
or U520 (N_520,In_1276,In_1571);
and U521 (N_521,In_1136,In_2435);
and U522 (N_522,In_245,In_1065);
nand U523 (N_523,In_2097,In_391);
nand U524 (N_524,In_1829,In_319);
nand U525 (N_525,In_1598,In_1915);
nor U526 (N_526,In_312,In_387);
nor U527 (N_527,In_2326,In_545);
nor U528 (N_528,In_293,In_1780);
and U529 (N_529,In_1191,In_1503);
and U530 (N_530,In_1950,In_370);
xor U531 (N_531,In_1013,In_891);
xnor U532 (N_532,In_107,In_1945);
nor U533 (N_533,In_1633,In_551);
or U534 (N_534,In_2087,In_1497);
nor U535 (N_535,In_724,In_1680);
nand U536 (N_536,In_233,In_2066);
and U537 (N_537,In_2499,In_1166);
or U538 (N_538,In_770,In_1256);
or U539 (N_539,In_14,In_2102);
and U540 (N_540,In_75,In_1124);
nand U541 (N_541,In_1903,In_1351);
nand U542 (N_542,In_1948,In_833);
nand U543 (N_543,In_711,In_1999);
or U544 (N_544,In_594,In_1217);
and U545 (N_545,In_1977,In_307);
or U546 (N_546,In_944,In_1809);
xor U547 (N_547,In_1359,In_1464);
or U548 (N_548,In_581,In_1358);
nand U549 (N_549,In_2233,In_1064);
and U550 (N_550,In_1896,In_362);
nand U551 (N_551,In_1395,In_206);
nand U552 (N_552,In_1531,In_37);
nor U553 (N_553,In_488,In_1886);
or U554 (N_554,In_1584,In_1208);
and U555 (N_555,In_1802,In_1225);
and U556 (N_556,In_653,In_1682);
or U557 (N_557,In_2450,In_815);
or U558 (N_558,In_2343,In_708);
nand U559 (N_559,In_1090,In_642);
or U560 (N_560,In_720,In_2410);
or U561 (N_561,In_513,In_187);
nand U562 (N_562,In_1429,In_1694);
xnor U563 (N_563,In_2362,In_747);
or U564 (N_564,In_2238,In_1699);
nand U565 (N_565,In_179,In_1363);
xnor U566 (N_566,In_194,In_661);
nand U567 (N_567,In_2139,In_2170);
nor U568 (N_568,In_2158,In_1690);
and U569 (N_569,In_2271,In_1533);
or U570 (N_570,In_907,In_29);
and U571 (N_571,In_420,In_1964);
or U572 (N_572,In_2224,In_2430);
and U573 (N_573,In_1808,In_1545);
nor U574 (N_574,In_1115,In_1392);
nor U575 (N_575,In_2016,In_2383);
nor U576 (N_576,In_595,In_190);
and U577 (N_577,In_1791,In_133);
nor U578 (N_578,In_276,In_2204);
or U579 (N_579,In_1354,In_1003);
and U580 (N_580,In_650,In_1823);
or U581 (N_581,In_217,In_2255);
or U582 (N_582,In_1317,In_1022);
nand U583 (N_583,In_1779,In_2334);
or U584 (N_584,In_2445,In_562);
or U585 (N_585,In_1041,In_956);
nand U586 (N_586,In_460,In_2064);
xnor U587 (N_587,In_2235,In_1279);
xnor U588 (N_588,In_726,In_65);
nand U589 (N_589,In_1868,In_2432);
nand U590 (N_590,In_885,In_1615);
nand U591 (N_591,In_244,In_1583);
and U592 (N_592,In_1110,In_226);
xor U593 (N_593,In_1514,In_2427);
nand U594 (N_594,In_184,In_124);
nor U595 (N_595,In_1830,In_253);
nand U596 (N_596,In_503,In_1453);
nor U597 (N_597,In_2247,In_1669);
and U598 (N_598,In_1140,In_275);
and U599 (N_599,In_2126,In_660);
nor U600 (N_600,In_1700,In_2008);
or U601 (N_601,In_709,In_2154);
nand U602 (N_602,In_110,In_308);
nor U603 (N_603,In_1493,In_2325);
nand U604 (N_604,In_512,In_1956);
or U605 (N_605,In_17,In_1981);
nand U606 (N_606,In_1156,In_779);
nor U607 (N_607,In_285,In_1119);
xor U608 (N_608,In_2120,In_411);
and U609 (N_609,In_658,In_473);
or U610 (N_610,In_2017,In_418);
xnor U611 (N_611,In_2184,In_1697);
or U612 (N_612,In_2050,In_1009);
and U613 (N_613,In_1741,In_874);
and U614 (N_614,In_2335,In_381);
nand U615 (N_615,In_1714,In_1930);
xnor U616 (N_616,In_129,In_1594);
or U617 (N_617,In_2033,In_168);
nor U618 (N_618,In_2065,In_1521);
xor U619 (N_619,In_225,In_373);
nand U620 (N_620,In_359,In_688);
nor U621 (N_621,In_390,In_1240);
nor U622 (N_622,In_2420,In_1378);
or U623 (N_623,In_2269,In_1622);
and U624 (N_624,In_2368,In_1897);
nand U625 (N_625,In_128,In_1753);
nand U626 (N_626,In_1269,In_383);
xor U627 (N_627,In_2375,In_1955);
and U628 (N_628,In_1006,In_1202);
and U629 (N_629,In_2360,In_2369);
nand U630 (N_630,In_282,In_746);
and U631 (N_631,In_149,In_8);
nand U632 (N_632,In_983,In_1411);
nand U633 (N_633,In_1481,In_1738);
nand U634 (N_634,In_1138,In_84);
or U635 (N_635,In_341,In_1538);
nor U636 (N_636,In_333,In_2024);
nand U637 (N_637,In_2220,In_2103);
and U638 (N_638,In_322,In_1600);
and U639 (N_639,In_943,In_1052);
nor U640 (N_640,In_2082,In_1854);
xor U641 (N_641,In_1647,In_851);
or U642 (N_642,In_79,In_1058);
and U643 (N_643,In_929,In_865);
nor U644 (N_644,In_564,In_446);
or U645 (N_645,In_1675,In_292);
or U646 (N_646,In_1433,In_1081);
nand U647 (N_647,In_277,In_237);
nand U648 (N_648,In_1603,In_240);
or U649 (N_649,In_382,In_1926);
and U650 (N_650,In_1151,In_2344);
nor U651 (N_651,In_1475,In_146);
and U652 (N_652,In_119,In_596);
or U653 (N_653,In_1996,In_1712);
or U654 (N_654,In_732,In_678);
and U655 (N_655,In_767,In_180);
nand U656 (N_656,In_2132,In_1026);
or U657 (N_657,In_648,In_741);
and U658 (N_658,In_2309,In_111);
and U659 (N_659,In_64,In_1570);
nor U660 (N_660,In_1683,In_2349);
and U661 (N_661,In_643,In_1508);
nor U662 (N_662,In_1875,In_622);
nor U663 (N_663,In_1895,In_1544);
nand U664 (N_664,In_1448,In_1080);
and U665 (N_665,In_603,In_155);
xor U666 (N_666,In_553,In_1025);
nand U667 (N_667,In_1295,In_1990);
xnor U668 (N_668,In_346,In_186);
nand U669 (N_669,In_1822,In_719);
or U670 (N_670,In_2037,In_1972);
xor U671 (N_671,In_442,In_831);
or U672 (N_672,In_1842,In_1366);
or U673 (N_673,In_1412,In_1368);
nand U674 (N_674,In_969,In_294);
and U675 (N_675,In_1470,In_1347);
or U676 (N_676,In_1468,In_1740);
nand U677 (N_677,In_911,In_618);
and U678 (N_678,In_2015,In_725);
nand U679 (N_679,In_7,In_2392);
nand U680 (N_680,In_2186,In_1904);
nor U681 (N_681,In_1125,In_2364);
and U682 (N_682,In_1721,In_1118);
xnor U683 (N_683,In_1247,In_1602);
or U684 (N_684,In_1229,In_992);
and U685 (N_685,In_151,In_2282);
nand U686 (N_686,In_1245,In_1123);
xor U687 (N_687,In_175,In_2416);
nor U688 (N_688,In_1327,In_1610);
or U689 (N_689,In_403,In_1344);
or U690 (N_690,In_429,In_763);
and U691 (N_691,In_228,In_1002);
and U692 (N_692,In_1550,In_1927);
and U693 (N_693,In_864,In_487);
nand U694 (N_694,In_654,In_1653);
or U695 (N_695,In_1417,In_11);
nand U696 (N_696,In_1861,In_1333);
nor U697 (N_697,In_338,In_1265);
and U698 (N_698,In_703,In_243);
and U699 (N_699,In_59,In_1198);
and U700 (N_700,In_91,In_1624);
or U701 (N_701,In_1280,In_1222);
and U702 (N_702,In_2474,In_1582);
and U703 (N_703,In_1710,In_2295);
or U704 (N_704,In_1762,In_2492);
nor U705 (N_705,In_1801,In_1512);
and U706 (N_706,In_2228,In_994);
or U707 (N_707,In_629,In_300);
xor U708 (N_708,In_379,In_96);
xnor U709 (N_709,In_1878,In_368);
nor U710 (N_710,In_73,In_1678);
and U711 (N_711,In_2078,In_1916);
and U712 (N_712,In_2320,In_2108);
or U713 (N_713,In_2200,In_2268);
nand U714 (N_714,In_2250,In_2199);
and U715 (N_715,In_2022,In_1322);
nor U716 (N_716,In_52,In_2241);
and U717 (N_717,In_677,In_1028);
nand U718 (N_718,In_1139,In_937);
or U719 (N_719,In_1273,In_1103);
or U720 (N_720,In_2387,In_423);
nor U721 (N_721,In_1971,In_1261);
nand U722 (N_722,In_1294,In_449);
nand U723 (N_723,In_12,In_2189);
nor U724 (N_724,In_1674,In_2197);
and U725 (N_725,In_1206,In_656);
and U726 (N_726,In_2128,In_1281);
or U727 (N_727,In_900,In_583);
and U728 (N_728,In_2351,In_472);
nand U729 (N_729,In_635,In_1288);
and U730 (N_730,In_705,In_1689);
nand U731 (N_731,In_1427,In_1593);
nor U732 (N_732,In_454,In_610);
nand U733 (N_733,In_1636,In_1212);
and U734 (N_734,In_1463,In_32);
and U735 (N_735,In_580,In_707);
nor U736 (N_736,In_1968,In_2245);
and U737 (N_737,In_1326,In_657);
or U738 (N_738,In_577,In_1248);
nand U739 (N_739,In_1766,In_255);
xnor U740 (N_740,In_662,In_369);
nand U741 (N_741,In_2354,In_2117);
or U742 (N_742,In_222,In_672);
nand U743 (N_743,In_1210,In_731);
and U744 (N_744,In_2328,In_142);
nor U745 (N_745,In_2083,In_2455);
xnor U746 (N_746,In_246,In_355);
nand U747 (N_747,In_2374,In_315);
and U748 (N_748,In_339,In_981);
nor U749 (N_749,In_385,In_1050);
nor U750 (N_750,In_1330,In_50);
and U751 (N_751,In_1383,In_1287);
and U752 (N_752,In_2003,In_837);
or U753 (N_753,In_482,In_1982);
and U754 (N_754,In_1628,In_164);
or U755 (N_755,In_1642,In_1944);
xor U756 (N_756,In_2056,In_2398);
or U757 (N_757,In_1574,In_261);
or U758 (N_758,In_752,In_1698);
or U759 (N_759,In_2054,In_1733);
nand U760 (N_760,In_262,In_1362);
or U761 (N_761,In_930,In_1399);
and U762 (N_762,In_489,In_886);
and U763 (N_763,In_848,In_939);
or U764 (N_764,In_714,In_286);
xor U765 (N_765,In_24,In_1718);
and U766 (N_766,In_2001,In_575);
xnor U767 (N_767,In_2467,In_49);
nor U768 (N_768,In_254,In_547);
nand U769 (N_769,In_2440,In_2101);
nor U770 (N_770,In_1943,In_2436);
and U771 (N_771,In_388,In_1318);
nand U772 (N_772,In_1983,In_1609);
and U773 (N_773,In_1693,In_1246);
nor U774 (N_774,In_1037,In_1529);
and U775 (N_775,In_869,In_74);
or U776 (N_776,In_1310,In_1239);
nor U777 (N_777,In_450,In_882);
nand U778 (N_778,In_572,In_389);
xor U779 (N_779,In_247,In_600);
and U780 (N_780,In_1719,In_1543);
and U781 (N_781,In_1062,In_972);
nand U782 (N_782,In_1356,In_2071);
nand U783 (N_783,In_2012,In_604);
and U784 (N_784,In_1591,In_2142);
nand U785 (N_785,In_397,In_2272);
nor U786 (N_786,In_1953,In_923);
nor U787 (N_787,In_1419,In_1800);
nand U788 (N_788,In_344,In_1877);
and U789 (N_789,In_1817,In_2073);
or U790 (N_790,In_1283,In_2287);
nor U791 (N_791,In_1770,In_1408);
and U792 (N_792,In_2353,In_466);
and U793 (N_793,In_1816,In_2130);
and U794 (N_794,In_350,In_318);
or U795 (N_795,In_1711,In_908);
nand U796 (N_796,In_1061,In_1014);
nand U797 (N_797,In_132,In_1029);
or U798 (N_798,In_337,In_793);
xor U799 (N_799,In_977,In_534);
nand U800 (N_800,In_1126,In_1918);
xor U801 (N_801,In_1325,In_1122);
or U802 (N_802,In_2236,In_474);
and U803 (N_803,In_19,In_1704);
or U804 (N_804,In_1942,In_67);
and U805 (N_805,In_1057,In_2227);
or U806 (N_806,In_682,In_1590);
and U807 (N_807,In_1188,In_505);
and U808 (N_808,In_1589,In_490);
and U809 (N_809,In_591,In_2385);
nand U810 (N_810,In_2229,In_3);
and U811 (N_811,In_1781,In_1147);
nor U812 (N_812,In_1567,In_1458);
nor U813 (N_813,In_987,In_148);
and U814 (N_814,In_1909,In_2340);
nand U815 (N_815,In_584,In_611);
nand U816 (N_816,In_520,In_2138);
xnor U817 (N_817,In_1360,In_880);
and U818 (N_818,In_1913,In_188);
xor U819 (N_819,In_1777,In_140);
and U820 (N_820,In_1382,In_1853);
nor U821 (N_821,In_1821,In_1214);
and U822 (N_822,In_2188,In_723);
and U823 (N_823,In_608,In_2231);
nand U824 (N_824,In_2131,In_1772);
nand U825 (N_825,In_1805,In_1732);
or U826 (N_826,In_1150,In_88);
and U827 (N_827,In_510,In_895);
nand U828 (N_828,In_1339,In_901);
nor U829 (N_829,In_782,In_1644);
or U830 (N_830,In_422,In_2143);
or U831 (N_831,In_1069,In_1960);
nor U832 (N_832,In_1935,In_1691);
or U833 (N_833,In_171,In_367);
nand U834 (N_834,In_1209,In_1561);
or U835 (N_835,In_256,In_1914);
or U836 (N_836,In_405,In_1056);
nor U837 (N_837,In_1290,In_2338);
nand U838 (N_838,In_2051,In_920);
xnor U839 (N_839,In_99,In_2090);
and U840 (N_840,In_1627,In_2478);
nor U841 (N_841,In_928,In_105);
or U842 (N_842,In_1806,In_1085);
nor U843 (N_843,In_1152,In_1752);
nor U844 (N_844,In_1506,In_788);
and U845 (N_845,In_1907,In_471);
or U846 (N_846,In_321,In_2031);
or U847 (N_847,In_1060,In_2226);
and U848 (N_848,In_1771,In_208);
and U849 (N_849,In_843,In_2248);
or U850 (N_850,In_773,In_1812);
nor U851 (N_851,In_2040,In_829);
and U852 (N_852,In_1015,In_514);
xor U853 (N_853,In_2304,In_2230);
or U854 (N_854,In_1759,In_1958);
nand U855 (N_855,In_2316,In_1172);
and U856 (N_856,In_598,In_1525);
nor U857 (N_857,In_1471,In_1937);
nor U858 (N_858,In_2032,In_542);
and U859 (N_859,In_765,In_2457);
and U860 (N_860,In_1947,In_888);
or U861 (N_861,In_836,In_1494);
nor U862 (N_862,In_2495,In_1798);
nand U863 (N_863,In_655,In_1859);
nand U864 (N_864,In_1604,In_1414);
xnor U865 (N_865,In_1688,In_1352);
nor U866 (N_866,In_1405,In_1949);
or U867 (N_867,In_936,In_327);
and U868 (N_868,In_945,In_1952);
nand U869 (N_869,In_2217,In_1426);
nand U870 (N_870,In_108,In_2114);
or U871 (N_871,In_1039,In_1192);
and U872 (N_872,In_754,In_380);
or U873 (N_873,In_2289,In_1932);
or U874 (N_874,In_1457,In_202);
and U875 (N_875,In_2327,In_2207);
nand U876 (N_876,In_1504,In_993);
nor U877 (N_877,In_1505,In_2160);
and U878 (N_878,In_1486,In_2415);
nand U879 (N_879,In_1818,In_2296);
nor U880 (N_880,In_28,In_1840);
and U881 (N_881,In_2380,In_1866);
or U882 (N_882,In_2411,In_1289);
or U883 (N_883,In_1980,In_2162);
and U884 (N_884,In_1211,In_112);
nand U885 (N_885,In_2444,In_481);
nand U886 (N_886,In_1984,In_183);
or U887 (N_887,In_156,In_950);
xnor U888 (N_888,In_2191,In_248);
nor U889 (N_889,In_1658,In_2168);
nand U890 (N_890,In_2075,In_1979);
and U891 (N_891,In_2203,In_1563);
nor U892 (N_892,In_1803,In_2095);
nor U893 (N_893,In_592,In_616);
and U894 (N_894,In_2127,In_2145);
nor U895 (N_895,In_1044,In_721);
or U896 (N_896,In_212,In_821);
and U897 (N_897,In_1587,In_1010);
or U898 (N_898,In_877,In_1425);
and U899 (N_899,In_2301,In_1146);
and U900 (N_900,In_1860,In_2113);
or U901 (N_901,In_1467,In_878);
or U902 (N_902,In_1231,In_2053);
xor U903 (N_903,In_220,In_798);
nor U904 (N_904,In_701,In_828);
nand U905 (N_905,In_147,In_1195);
nand U906 (N_906,In_227,In_990);
nand U907 (N_907,In_567,In_984);
nand U908 (N_908,In_1862,In_1649);
nand U909 (N_909,In_1452,In_614);
nor U910 (N_910,In_1632,In_2459);
nor U911 (N_911,In_1114,In_1601);
or U912 (N_912,In_2469,In_1319);
nor U913 (N_913,In_834,In_727);
and U914 (N_914,In_1157,In_2254);
and U915 (N_915,In_2256,In_2431);
nor U916 (N_916,In_1332,In_1539);
xnor U917 (N_917,In_1311,In_1846);
or U918 (N_918,In_713,In_2239);
and U919 (N_919,In_1336,In_2140);
xnor U920 (N_920,In_1588,In_1176);
nand U921 (N_921,In_691,In_1353);
nand U922 (N_922,In_2284,In_996);
nor U923 (N_923,In_165,In_2192);
xor U924 (N_924,In_1132,In_1259);
or U925 (N_925,In_1619,In_1524);
nand U926 (N_926,In_313,In_1751);
nor U927 (N_927,In_2490,In_963);
or U928 (N_928,In_2180,In_1235);
or U929 (N_929,In_2442,In_475);
or U930 (N_930,In_817,In_1098);
and U931 (N_931,In_876,In_1300);
or U932 (N_932,In_305,In_1078);
or U933 (N_933,In_2311,In_690);
and U934 (N_934,In_1556,In_326);
nand U935 (N_935,In_1892,In_290);
and U936 (N_936,In_733,In_1434);
and U937 (N_937,In_1200,In_41);
nand U938 (N_938,In_2177,In_1173);
or U939 (N_939,In_2218,In_1159);
nor U940 (N_940,In_301,In_810);
nor U941 (N_941,In_22,In_1001);
nor U942 (N_942,In_157,In_541);
nor U943 (N_943,In_392,In_818);
nor U944 (N_944,In_1402,In_1163);
nand U945 (N_945,In_174,In_120);
nor U946 (N_946,In_976,In_1092);
nor U947 (N_947,In_1562,In_563);
nand U948 (N_948,In_1439,In_2434);
and U949 (N_949,In_903,In_352);
xor U950 (N_950,In_692,In_1807);
nor U951 (N_951,In_2020,In_153);
nand U952 (N_952,In_1509,In_807);
and U953 (N_953,In_2476,In_759);
xor U954 (N_954,In_706,In_1263);
nand U955 (N_955,In_652,In_178);
or U956 (N_956,In_2412,In_1105);
or U957 (N_957,In_1393,In_2408);
or U958 (N_958,In_2381,In_1272);
and U959 (N_959,In_2363,In_219);
nand U960 (N_960,In_772,In_971);
xor U961 (N_961,In_966,In_1761);
xor U962 (N_962,In_1345,In_960);
xor U963 (N_963,In_1421,In_1137);
nand U964 (N_964,In_1607,In_61);
nand U965 (N_965,In_66,In_386);
nor U966 (N_966,In_234,In_722);
nand U967 (N_967,In_698,In_2336);
and U968 (N_968,In_1706,In_2123);
xnor U969 (N_969,In_1230,In_1555);
nor U970 (N_970,In_484,In_56);
nand U971 (N_971,In_1975,In_116);
nor U972 (N_972,In_1966,In_272);
or U973 (N_973,In_2479,In_571);
and U974 (N_974,In_554,In_1199);
nand U975 (N_975,In_1532,In_1726);
nor U976 (N_976,In_271,In_775);
nand U977 (N_977,In_1993,In_257);
nor U978 (N_978,In_2165,In_1129);
and U979 (N_979,In_2072,In_1456);
nor U980 (N_980,In_855,In_68);
nand U981 (N_981,In_1670,In_2323);
or U982 (N_982,In_2406,In_870);
and U983 (N_983,In_1888,In_1579);
or U984 (N_984,In_1787,In_358);
and U985 (N_985,In_740,In_756);
and U986 (N_986,In_1221,In_2099);
xor U987 (N_987,In_1027,In_1873);
or U988 (N_988,In_2359,In_297);
xor U989 (N_989,In_816,In_2137);
nor U990 (N_990,In_163,In_1773);
nand U991 (N_991,In_1599,In_1183);
nand U992 (N_992,In_363,In_1404);
and U993 (N_993,In_18,In_2497);
and U994 (N_994,In_2221,In_1969);
nor U995 (N_995,In_1334,In_311);
nor U996 (N_996,In_2278,In_342);
xnor U997 (N_997,In_1297,In_838);
and U998 (N_998,In_632,In_1130);
nor U999 (N_999,In_651,In_252);
or U1000 (N_1000,In_2018,In_1266);
nand U1001 (N_1001,In_1376,In_524);
or U1002 (N_1002,In_1922,In_1224);
and U1003 (N_1003,In_1552,In_309);
or U1004 (N_1004,In_2276,In_430);
and U1005 (N_1005,In_57,In_631);
nor U1006 (N_1006,In_634,In_1906);
nor U1007 (N_1007,In_2049,In_39);
or U1008 (N_1008,In_375,In_354);
nor U1009 (N_1009,In_172,In_1474);
xnor U1010 (N_1010,In_432,In_1695);
and U1011 (N_1011,In_1559,In_1019);
nand U1012 (N_1012,In_2134,In_1238);
nand U1013 (N_1013,In_1033,In_1898);
and U1014 (N_1014,In_1722,In_2109);
nand U1015 (N_1015,In_1168,In_205);
nor U1016 (N_1016,In_947,In_2240);
and U1017 (N_1017,In_2347,In_1055);
xnor U1018 (N_1018,In_1564,In_862);
nor U1019 (N_1019,In_1331,In_1244);
nand U1020 (N_1020,In_845,In_964);
xnor U1021 (N_1021,In_742,In_1223);
or U1022 (N_1022,In_1668,In_1101);
nor U1023 (N_1023,In_94,In_1510);
or U1024 (N_1024,In_978,In_2317);
nand U1025 (N_1025,In_1709,In_666);
and U1026 (N_1026,In_86,In_630);
or U1027 (N_1027,In_207,In_2067);
nand U1028 (N_1028,In_2118,In_465);
xnor U1029 (N_1029,In_1036,In_871);
nor U1030 (N_1030,In_2274,In_2464);
nand U1031 (N_1031,In_1769,In_2115);
nor U1032 (N_1032,In_1912,In_456);
nand U1033 (N_1033,In_121,In_1728);
or U1034 (N_1034,In_1171,In_1705);
or U1035 (N_1035,In_1487,In_518);
nor U1036 (N_1036,In_98,In_1498);
and U1037 (N_1037,In_25,In_1385);
and U1038 (N_1038,In_2356,In_2357);
nor U1039 (N_1039,In_1492,In_1484);
xor U1040 (N_1040,In_63,In_1756);
or U1041 (N_1041,In_1135,In_748);
or U1042 (N_1042,In_2149,In_1885);
nand U1043 (N_1043,In_1120,In_1613);
nor U1044 (N_1044,In_1012,In_2106);
nand U1045 (N_1045,In_906,In_1703);
nor U1046 (N_1046,In_1020,In_1596);
nor U1047 (N_1047,In_1381,In_2477);
nor U1048 (N_1048,In_2141,In_1630);
nor U1049 (N_1049,In_1308,In_131);
nor U1050 (N_1050,In_840,In_2275);
nor U1051 (N_1051,In_1178,In_1391);
and U1052 (N_1052,In_1337,In_270);
nand U1053 (N_1053,In_2318,In_2237);
nor U1054 (N_1054,In_191,In_1871);
nor U1055 (N_1055,In_1837,In_857);
nor U1056 (N_1056,In_2045,In_210);
and U1057 (N_1057,In_1511,In_182);
nor U1058 (N_1058,In_1890,In_1742);
or U1059 (N_1059,In_568,In_1000);
nand U1060 (N_1060,In_410,In_1285);
nand U1061 (N_1061,In_1401,In_1797);
nand U1062 (N_1062,In_1573,In_2011);
and U1063 (N_1063,In_1864,In_1865);
xor U1064 (N_1064,In_1776,In_1196);
or U1065 (N_1065,In_2390,In_2379);
xor U1066 (N_1066,In_2371,In_2352);
or U1067 (N_1067,In_1618,In_955);
or U1068 (N_1068,In_1547,In_414);
or U1069 (N_1069,In_1617,In_2088);
nand U1070 (N_1070,In_1320,In_1343);
xor U1071 (N_1071,In_605,In_1611);
nor U1072 (N_1072,In_1723,In_1491);
nor U1073 (N_1073,In_2393,In_679);
or U1074 (N_1074,In_1250,In_431);
nor U1075 (N_1075,In_2074,In_1194);
or U1076 (N_1076,In_394,In_1499);
nor U1077 (N_1077,In_1576,In_2069);
nand U1078 (N_1078,In_2222,In_2172);
nand U1079 (N_1079,In_1804,In_1577);
nor U1080 (N_1080,In_1477,In_2438);
or U1081 (N_1081,In_1207,In_1384);
or U1082 (N_1082,In_1638,In_2243);
nand U1083 (N_1083,In_393,In_762);
or U1084 (N_1084,In_445,In_1030);
nand U1085 (N_1085,In_2337,In_1717);
or U1086 (N_1086,In_1946,In_1018);
nand U1087 (N_1087,In_26,In_127);
or U1088 (N_1088,In_1299,In_1228);
nand U1089 (N_1089,In_822,In_1380);
and U1090 (N_1090,In_2030,In_1831);
and U1091 (N_1091,In_1962,In_457);
or U1092 (N_1092,In_1568,In_2161);
nor U1093 (N_1093,In_462,In_697);
and U1094 (N_1094,In_76,In_2249);
or U1095 (N_1095,In_1252,In_2386);
nand U1096 (N_1096,In_1815,In_360);
xor U1097 (N_1097,In_999,In_1237);
and U1098 (N_1098,In_1872,In_2281);
and U1099 (N_1099,In_502,In_263);
or U1100 (N_1100,In_951,In_700);
nor U1101 (N_1101,In_2404,In_415);
nor U1102 (N_1102,In_1811,In_942);
nand U1103 (N_1103,In_2060,In_1938);
and U1104 (N_1104,In_1672,In_2484);
or U1105 (N_1105,In_800,In_1040);
nor U1106 (N_1106,In_1795,In_1880);
and U1107 (N_1107,In_1876,In_1754);
or U1108 (N_1108,In_716,In_1432);
or U1109 (N_1109,In_617,In_447);
xnor U1110 (N_1110,In_852,In_1077);
nor U1111 (N_1111,In_451,In_412);
nor U1112 (N_1112,In_728,In_536);
and U1113 (N_1113,In_1220,In_2157);
xor U1114 (N_1114,In_1017,In_998);
nor U1115 (N_1115,In_495,In_1476);
or U1116 (N_1116,In_835,In_40);
nand U1117 (N_1117,In_1073,In_1450);
and U1118 (N_1118,In_1145,In_1986);
xnor U1119 (N_1119,In_1251,In_345);
or U1120 (N_1120,In_1863,In_1043);
or U1121 (N_1121,In_1369,In_695);
or U1122 (N_1122,In_2285,In_45);
and U1123 (N_1123,In_199,In_2183);
nand U1124 (N_1124,In_883,In_1189);
nand U1125 (N_1125,In_33,In_2419);
or U1126 (N_1126,In_1219,In_1526);
or U1127 (N_1127,In_2057,In_258);
and U1128 (N_1128,In_1891,In_2019);
nand U1129 (N_1129,In_221,In_1307);
and U1130 (N_1130,In_2259,In_1258);
and U1131 (N_1131,In_2080,In_2290);
nand U1132 (N_1132,In_2263,In_1443);
nor U1133 (N_1133,In_1243,In_334);
or U1134 (N_1134,In_1793,In_2093);
nor U1135 (N_1135,In_348,In_866);
or U1136 (N_1136,In_2449,In_783);
or U1137 (N_1137,In_1666,In_1656);
or U1138 (N_1138,In_934,In_681);
and U1139 (N_1139,In_1148,In_1905);
and U1140 (N_1140,In_340,In_1293);
xnor U1141 (N_1141,In_2446,In_1213);
xnor U1142 (N_1142,In_1255,In_1657);
nor U1143 (N_1143,In_2208,In_43);
and U1144 (N_1144,In_464,In_1645);
or U1145 (N_1145,In_925,In_1569);
nand U1146 (N_1146,In_1997,In_570);
nand U1147 (N_1147,In_1181,In_1518);
or U1148 (N_1148,In_211,In_1920);
nand U1149 (N_1149,In_2361,In_2491);
nor U1150 (N_1150,In_854,In_2111);
nor U1151 (N_1151,In_2006,In_2009);
or U1152 (N_1152,In_689,In_1270);
or U1153 (N_1153,In_625,In_1302);
nand U1154 (N_1154,In_832,In_2163);
or U1155 (N_1155,In_126,In_1961);
or U1156 (N_1156,In_117,In_1462);
nand U1157 (N_1157,In_1513,In_1566);
nand U1158 (N_1158,In_766,In_774);
and U1159 (N_1159,In_122,In_62);
or U1160 (N_1160,In_1260,In_46);
and U1161 (N_1161,In_1407,In_329);
nand U1162 (N_1162,In_1743,In_1416);
nor U1163 (N_1163,In_921,In_2232);
nand U1164 (N_1164,In_1978,In_529);
or U1165 (N_1165,In_2424,In_2299);
or U1166 (N_1166,In_1893,In_685);
or U1167 (N_1167,In_1149,In_2070);
nand U1168 (N_1168,In_1625,In_533);
nor U1169 (N_1169,In_371,In_374);
nor U1170 (N_1170,In_377,In_1899);
nor U1171 (N_1171,In_1749,In_1005);
and U1172 (N_1172,In_1323,In_496);
and U1173 (N_1173,In_1575,In_2136);
or U1174 (N_1174,In_2443,In_1629);
and U1175 (N_1175,In_2094,In_1553);
or U1176 (N_1176,In_2173,In_135);
nor U1177 (N_1177,In_2223,In_1856);
and U1178 (N_1178,In_435,In_1626);
nand U1179 (N_1179,In_498,In_236);
nor U1180 (N_1180,In_479,In_646);
and U1181 (N_1181,In_1928,In_602);
or U1182 (N_1182,In_1606,In_2447);
xnor U1183 (N_1183,In_718,In_1792);
or U1184 (N_1184,In_811,In_961);
and U1185 (N_1185,In_162,In_549);
nand U1186 (N_1186,In_1109,In_2026);
nand U1187 (N_1187,In_2147,In_2313);
and U1188 (N_1188,In_887,In_2355);
and U1189 (N_1189,In_683,In_1931);
and U1190 (N_1190,In_2052,In_324);
xnor U1191 (N_1191,In_1046,In_2179);
xor U1192 (N_1192,In_2423,In_946);
or U1193 (N_1193,In_2202,In_593);
or U1194 (N_1194,In_2010,In_997);
nand U1195 (N_1195,In_1370,In_1662);
nor U1196 (N_1196,In_2107,In_2004);
nand U1197 (N_1197,In_1127,In_71);
nand U1198 (N_1198,In_304,In_2);
nor U1199 (N_1199,In_2487,In_806);
nand U1200 (N_1200,In_2358,In_1646);
nand U1201 (N_1201,In_1161,In_1278);
or U1202 (N_1202,In_781,In_384);
nand U1203 (N_1203,In_769,In_347);
nand U1204 (N_1204,In_1813,In_1313);
nand U1205 (N_1205,In_1727,In_760);
and U1206 (N_1206,In_2092,In_764);
nor U1207 (N_1207,In_80,In_58);
or U1208 (N_1208,In_982,In_1141);
or U1209 (N_1209,In_448,In_145);
and U1210 (N_1210,In_1736,In_578);
and U1211 (N_1211,In_606,In_1523);
and U1212 (N_1212,In_238,In_353);
nor U1213 (N_1213,In_771,In_1558);
or U1214 (N_1214,In_1870,In_1917);
nor U1215 (N_1215,In_2155,In_2279);
or U1216 (N_1216,In_2146,In_1306);
nand U1217 (N_1217,In_849,In_673);
nor U1218 (N_1218,In_1612,In_2125);
nor U1219 (N_1219,In_343,In_1924);
or U1220 (N_1220,In_1472,In_1799);
nand U1221 (N_1221,In_515,In_2482);
or U1222 (N_1222,In_1415,In_189);
or U1223 (N_1223,In_850,In_433);
nor U1224 (N_1224,In_2062,In_620);
and U1225 (N_1225,In_349,In_2366);
nand U1226 (N_1226,In_1681,In_1291);
nand U1227 (N_1227,In_1377,In_1760);
nand U1228 (N_1228,In_922,In_2280);
nor U1229 (N_1229,In_483,In_1008);
or U1230 (N_1230,In_1789,In_1);
and U1231 (N_1231,In_803,In_778);
nand U1232 (N_1232,In_597,In_1786);
nor U1233 (N_1233,In_873,In_1655);
nand U1234 (N_1234,In_239,In_306);
and U1235 (N_1235,In_1134,In_2148);
or U1236 (N_1236,In_795,In_1438);
nand U1237 (N_1237,In_2460,In_2283);
or U1238 (N_1238,In_590,In_2079);
and U1239 (N_1239,In_780,In_1940);
nor U1240 (N_1240,In_158,In_137);
or U1241 (N_1241,In_1350,In_899);
or U1242 (N_1242,In_569,In_1654);
xnor U1243 (N_1243,In_60,In_23);
or U1244 (N_1244,In_638,In_70);
and U1245 (N_1245,In_2288,In_1249);
nor U1246 (N_1246,In_426,In_461);
nand U1247 (N_1247,In_952,In_1910);
and U1248 (N_1248,In_266,In_1184);
or U1249 (N_1249,In_167,In_421);
nand U1250 (N_1250,In_464,In_1023);
nor U1251 (N_1251,In_2270,In_1668);
nor U1252 (N_1252,In_1823,In_410);
or U1253 (N_1253,In_2291,In_1555);
and U1254 (N_1254,In_1163,In_1622);
and U1255 (N_1255,In_340,In_239);
or U1256 (N_1256,In_1206,In_159);
nor U1257 (N_1257,In_780,In_1659);
nor U1258 (N_1258,In_1565,In_2451);
nor U1259 (N_1259,In_437,In_137);
or U1260 (N_1260,In_1038,In_1303);
or U1261 (N_1261,In_4,In_1116);
xor U1262 (N_1262,In_2306,In_336);
and U1263 (N_1263,In_1970,In_2349);
nand U1264 (N_1264,In_1107,In_1003);
nand U1265 (N_1265,In_916,In_1971);
or U1266 (N_1266,In_2402,In_33);
or U1267 (N_1267,In_2384,In_1031);
nand U1268 (N_1268,In_1726,In_1037);
or U1269 (N_1269,In_1528,In_1033);
and U1270 (N_1270,In_2108,In_1328);
and U1271 (N_1271,In_820,In_1285);
or U1272 (N_1272,In_29,In_1664);
nor U1273 (N_1273,In_1615,In_898);
and U1274 (N_1274,In_739,In_282);
or U1275 (N_1275,In_1178,In_998);
nor U1276 (N_1276,In_548,In_863);
nand U1277 (N_1277,In_1690,In_851);
or U1278 (N_1278,In_1353,In_680);
nand U1279 (N_1279,In_813,In_429);
and U1280 (N_1280,In_1643,In_697);
xnor U1281 (N_1281,In_1420,In_2097);
xor U1282 (N_1282,In_267,In_255);
or U1283 (N_1283,In_2029,In_1354);
and U1284 (N_1284,In_222,In_961);
nand U1285 (N_1285,In_373,In_468);
or U1286 (N_1286,In_2285,In_510);
and U1287 (N_1287,In_176,In_2232);
nor U1288 (N_1288,In_1104,In_426);
xnor U1289 (N_1289,In_2441,In_1725);
nand U1290 (N_1290,In_1475,In_2006);
xnor U1291 (N_1291,In_898,In_1520);
and U1292 (N_1292,In_982,In_388);
nor U1293 (N_1293,In_885,In_1725);
and U1294 (N_1294,In_2292,In_1938);
and U1295 (N_1295,In_856,In_207);
or U1296 (N_1296,In_540,In_1981);
nand U1297 (N_1297,In_1532,In_838);
or U1298 (N_1298,In_388,In_1208);
xnor U1299 (N_1299,In_1225,In_215);
nor U1300 (N_1300,In_219,In_1003);
or U1301 (N_1301,In_1517,In_313);
nand U1302 (N_1302,In_862,In_1846);
and U1303 (N_1303,In_1112,In_301);
nand U1304 (N_1304,In_2282,In_1758);
and U1305 (N_1305,In_2279,In_2248);
nor U1306 (N_1306,In_2227,In_1478);
nand U1307 (N_1307,In_444,In_1756);
nor U1308 (N_1308,In_2322,In_2253);
or U1309 (N_1309,In_1612,In_1923);
nor U1310 (N_1310,In_1668,In_1298);
nand U1311 (N_1311,In_663,In_2117);
nand U1312 (N_1312,In_177,In_2275);
and U1313 (N_1313,In_1865,In_2216);
or U1314 (N_1314,In_605,In_1325);
nor U1315 (N_1315,In_1409,In_839);
and U1316 (N_1316,In_987,In_246);
or U1317 (N_1317,In_671,In_1650);
xor U1318 (N_1318,In_2476,In_352);
and U1319 (N_1319,In_2449,In_1499);
nand U1320 (N_1320,In_454,In_770);
nand U1321 (N_1321,In_221,In_2096);
nand U1322 (N_1322,In_750,In_1624);
or U1323 (N_1323,In_2181,In_1363);
nor U1324 (N_1324,In_139,In_636);
nor U1325 (N_1325,In_1097,In_517);
and U1326 (N_1326,In_1627,In_357);
or U1327 (N_1327,In_778,In_118);
or U1328 (N_1328,In_252,In_1521);
or U1329 (N_1329,In_523,In_2473);
xor U1330 (N_1330,In_349,In_1095);
xor U1331 (N_1331,In_447,In_174);
xor U1332 (N_1332,In_2198,In_1168);
xor U1333 (N_1333,In_543,In_372);
or U1334 (N_1334,In_1839,In_827);
and U1335 (N_1335,In_434,In_650);
or U1336 (N_1336,In_666,In_1142);
and U1337 (N_1337,In_627,In_945);
nand U1338 (N_1338,In_1540,In_2020);
nor U1339 (N_1339,In_188,In_637);
or U1340 (N_1340,In_777,In_1880);
or U1341 (N_1341,In_984,In_1229);
and U1342 (N_1342,In_1106,In_2244);
nand U1343 (N_1343,In_25,In_1568);
nand U1344 (N_1344,In_972,In_2484);
or U1345 (N_1345,In_808,In_2371);
xor U1346 (N_1346,In_103,In_1130);
or U1347 (N_1347,In_35,In_1750);
nand U1348 (N_1348,In_746,In_2427);
and U1349 (N_1349,In_2366,In_245);
nor U1350 (N_1350,In_78,In_687);
nor U1351 (N_1351,In_1527,In_320);
xor U1352 (N_1352,In_2136,In_1109);
or U1353 (N_1353,In_770,In_2074);
and U1354 (N_1354,In_439,In_857);
or U1355 (N_1355,In_90,In_1202);
and U1356 (N_1356,In_905,In_406);
or U1357 (N_1357,In_1088,In_737);
and U1358 (N_1358,In_943,In_809);
nor U1359 (N_1359,In_807,In_816);
and U1360 (N_1360,In_1204,In_841);
nand U1361 (N_1361,In_502,In_939);
or U1362 (N_1362,In_919,In_492);
or U1363 (N_1363,In_2368,In_1161);
nor U1364 (N_1364,In_1721,In_980);
xor U1365 (N_1365,In_485,In_789);
and U1366 (N_1366,In_2131,In_2159);
and U1367 (N_1367,In_947,In_1365);
or U1368 (N_1368,In_1813,In_2409);
and U1369 (N_1369,In_378,In_2357);
or U1370 (N_1370,In_2439,In_1037);
nor U1371 (N_1371,In_834,In_359);
xnor U1372 (N_1372,In_1790,In_482);
nor U1373 (N_1373,In_828,In_2255);
or U1374 (N_1374,In_876,In_386);
or U1375 (N_1375,In_2228,In_2066);
nor U1376 (N_1376,In_818,In_537);
nand U1377 (N_1377,In_209,In_992);
and U1378 (N_1378,In_1235,In_1346);
or U1379 (N_1379,In_1527,In_1780);
nor U1380 (N_1380,In_542,In_2265);
or U1381 (N_1381,In_2400,In_1104);
and U1382 (N_1382,In_2320,In_1647);
and U1383 (N_1383,In_770,In_2047);
and U1384 (N_1384,In_572,In_489);
and U1385 (N_1385,In_1913,In_84);
or U1386 (N_1386,In_916,In_2420);
nor U1387 (N_1387,In_272,In_706);
nand U1388 (N_1388,In_1900,In_1649);
nand U1389 (N_1389,In_1386,In_1734);
and U1390 (N_1390,In_249,In_1575);
nand U1391 (N_1391,In_2056,In_2269);
nor U1392 (N_1392,In_28,In_25);
or U1393 (N_1393,In_700,In_1334);
nor U1394 (N_1394,In_541,In_1102);
nor U1395 (N_1395,In_1078,In_2381);
and U1396 (N_1396,In_1474,In_1564);
and U1397 (N_1397,In_13,In_967);
nor U1398 (N_1398,In_2421,In_2339);
xnor U1399 (N_1399,In_608,In_1740);
nor U1400 (N_1400,In_1050,In_777);
nor U1401 (N_1401,In_1178,In_570);
or U1402 (N_1402,In_1611,In_58);
nand U1403 (N_1403,In_1697,In_1411);
nand U1404 (N_1404,In_2308,In_2226);
or U1405 (N_1405,In_264,In_889);
nand U1406 (N_1406,In_1660,In_1929);
nand U1407 (N_1407,In_1077,In_2428);
and U1408 (N_1408,In_1749,In_1106);
xor U1409 (N_1409,In_1997,In_1350);
and U1410 (N_1410,In_368,In_503);
or U1411 (N_1411,In_1664,In_567);
and U1412 (N_1412,In_653,In_2107);
or U1413 (N_1413,In_211,In_1120);
nor U1414 (N_1414,In_1678,In_2293);
or U1415 (N_1415,In_766,In_15);
xnor U1416 (N_1416,In_851,In_699);
nor U1417 (N_1417,In_663,In_2380);
xnor U1418 (N_1418,In_1879,In_248);
or U1419 (N_1419,In_569,In_676);
nor U1420 (N_1420,In_2403,In_1463);
xnor U1421 (N_1421,In_263,In_348);
xnor U1422 (N_1422,In_748,In_2399);
or U1423 (N_1423,In_490,In_1942);
nand U1424 (N_1424,In_2273,In_1912);
xnor U1425 (N_1425,In_2495,In_564);
nor U1426 (N_1426,In_72,In_968);
or U1427 (N_1427,In_2048,In_1733);
nand U1428 (N_1428,In_2444,In_2397);
nor U1429 (N_1429,In_1549,In_2023);
nand U1430 (N_1430,In_397,In_1989);
or U1431 (N_1431,In_1368,In_1684);
and U1432 (N_1432,In_962,In_1650);
nor U1433 (N_1433,In_1720,In_425);
and U1434 (N_1434,In_1599,In_1009);
or U1435 (N_1435,In_366,In_2451);
nand U1436 (N_1436,In_324,In_2482);
and U1437 (N_1437,In_20,In_2013);
or U1438 (N_1438,In_1920,In_2241);
or U1439 (N_1439,In_1763,In_1720);
nor U1440 (N_1440,In_2397,In_1663);
and U1441 (N_1441,In_415,In_2095);
nor U1442 (N_1442,In_2341,In_1774);
and U1443 (N_1443,In_876,In_942);
or U1444 (N_1444,In_1365,In_2167);
and U1445 (N_1445,In_1887,In_1195);
nor U1446 (N_1446,In_1135,In_681);
or U1447 (N_1447,In_1228,In_1726);
and U1448 (N_1448,In_464,In_685);
nand U1449 (N_1449,In_1780,In_1831);
nor U1450 (N_1450,In_151,In_2101);
nand U1451 (N_1451,In_2069,In_1320);
nor U1452 (N_1452,In_1018,In_894);
nor U1453 (N_1453,In_442,In_1566);
and U1454 (N_1454,In_1056,In_1701);
nor U1455 (N_1455,In_1884,In_761);
or U1456 (N_1456,In_2423,In_34);
or U1457 (N_1457,In_1364,In_2457);
and U1458 (N_1458,In_1147,In_495);
or U1459 (N_1459,In_2403,In_378);
or U1460 (N_1460,In_1520,In_491);
xor U1461 (N_1461,In_1655,In_1076);
nor U1462 (N_1462,In_2345,In_1325);
nand U1463 (N_1463,In_403,In_2277);
nand U1464 (N_1464,In_1234,In_919);
and U1465 (N_1465,In_1430,In_1821);
xor U1466 (N_1466,In_1190,In_1738);
and U1467 (N_1467,In_2094,In_445);
nand U1468 (N_1468,In_1568,In_1160);
nor U1469 (N_1469,In_2051,In_1173);
nor U1470 (N_1470,In_1767,In_1194);
or U1471 (N_1471,In_1022,In_2469);
nor U1472 (N_1472,In_989,In_1572);
xor U1473 (N_1473,In_627,In_922);
and U1474 (N_1474,In_369,In_1165);
and U1475 (N_1475,In_984,In_929);
and U1476 (N_1476,In_1851,In_724);
nor U1477 (N_1477,In_2380,In_1014);
nor U1478 (N_1478,In_1742,In_597);
or U1479 (N_1479,In_732,In_1889);
or U1480 (N_1480,In_334,In_567);
or U1481 (N_1481,In_1517,In_849);
nor U1482 (N_1482,In_1354,In_1259);
or U1483 (N_1483,In_608,In_1546);
nand U1484 (N_1484,In_1500,In_499);
nand U1485 (N_1485,In_1496,In_1410);
or U1486 (N_1486,In_1636,In_133);
nor U1487 (N_1487,In_715,In_782);
and U1488 (N_1488,In_633,In_555);
xnor U1489 (N_1489,In_676,In_1003);
nand U1490 (N_1490,In_1822,In_440);
and U1491 (N_1491,In_1459,In_304);
and U1492 (N_1492,In_2236,In_440);
or U1493 (N_1493,In_2069,In_1478);
nand U1494 (N_1494,In_760,In_176);
nor U1495 (N_1495,In_1887,In_1872);
and U1496 (N_1496,In_2488,In_1278);
nand U1497 (N_1497,In_1175,In_2428);
nor U1498 (N_1498,In_439,In_493);
nor U1499 (N_1499,In_1753,In_1789);
or U1500 (N_1500,In_1902,In_975);
and U1501 (N_1501,In_1939,In_1636);
nand U1502 (N_1502,In_2229,In_5);
nand U1503 (N_1503,In_1048,In_1688);
or U1504 (N_1504,In_865,In_709);
or U1505 (N_1505,In_765,In_1229);
nor U1506 (N_1506,In_1562,In_1538);
xnor U1507 (N_1507,In_1101,In_1076);
nor U1508 (N_1508,In_2022,In_791);
or U1509 (N_1509,In_776,In_1374);
and U1510 (N_1510,In_343,In_1949);
or U1511 (N_1511,In_562,In_787);
and U1512 (N_1512,In_574,In_2215);
and U1513 (N_1513,In_454,In_100);
or U1514 (N_1514,In_886,In_1686);
and U1515 (N_1515,In_1124,In_1261);
or U1516 (N_1516,In_1672,In_736);
xor U1517 (N_1517,In_791,In_733);
and U1518 (N_1518,In_2199,In_909);
or U1519 (N_1519,In_1447,In_1781);
or U1520 (N_1520,In_2475,In_753);
or U1521 (N_1521,In_293,In_120);
nor U1522 (N_1522,In_1039,In_889);
and U1523 (N_1523,In_945,In_1562);
or U1524 (N_1524,In_1903,In_1313);
and U1525 (N_1525,In_1248,In_1992);
xor U1526 (N_1526,In_1670,In_373);
nor U1527 (N_1527,In_1106,In_99);
and U1528 (N_1528,In_521,In_715);
and U1529 (N_1529,In_126,In_1515);
nand U1530 (N_1530,In_1102,In_2055);
or U1531 (N_1531,In_1313,In_2038);
or U1532 (N_1532,In_2075,In_820);
or U1533 (N_1533,In_1117,In_539);
or U1534 (N_1534,In_1388,In_2333);
nor U1535 (N_1535,In_283,In_388);
nand U1536 (N_1536,In_891,In_1074);
and U1537 (N_1537,In_646,In_1060);
and U1538 (N_1538,In_1065,In_551);
and U1539 (N_1539,In_1968,In_1730);
nand U1540 (N_1540,In_159,In_2339);
nor U1541 (N_1541,In_454,In_308);
nor U1542 (N_1542,In_1482,In_2350);
or U1543 (N_1543,In_648,In_967);
nand U1544 (N_1544,In_372,In_1748);
nor U1545 (N_1545,In_630,In_2412);
and U1546 (N_1546,In_2149,In_27);
and U1547 (N_1547,In_1594,In_458);
nor U1548 (N_1548,In_2271,In_798);
nand U1549 (N_1549,In_510,In_224);
nor U1550 (N_1550,In_750,In_1719);
nand U1551 (N_1551,In_1186,In_841);
nand U1552 (N_1552,In_410,In_2318);
and U1553 (N_1553,In_1040,In_2186);
nand U1554 (N_1554,In_421,In_1991);
or U1555 (N_1555,In_1572,In_1641);
or U1556 (N_1556,In_781,In_332);
or U1557 (N_1557,In_673,In_546);
and U1558 (N_1558,In_2162,In_162);
or U1559 (N_1559,In_2101,In_373);
and U1560 (N_1560,In_1820,In_2168);
xor U1561 (N_1561,In_1299,In_624);
or U1562 (N_1562,In_1102,In_1820);
and U1563 (N_1563,In_707,In_200);
or U1564 (N_1564,In_302,In_1619);
or U1565 (N_1565,In_1904,In_259);
and U1566 (N_1566,In_526,In_988);
nor U1567 (N_1567,In_2143,In_2272);
and U1568 (N_1568,In_1621,In_139);
nand U1569 (N_1569,In_1415,In_154);
xor U1570 (N_1570,In_2392,In_874);
and U1571 (N_1571,In_409,In_422);
nand U1572 (N_1572,In_216,In_2037);
nor U1573 (N_1573,In_1561,In_841);
nor U1574 (N_1574,In_462,In_1362);
and U1575 (N_1575,In_339,In_2282);
or U1576 (N_1576,In_869,In_1914);
or U1577 (N_1577,In_1320,In_2420);
nand U1578 (N_1578,In_326,In_637);
nor U1579 (N_1579,In_1338,In_1485);
nor U1580 (N_1580,In_82,In_2242);
xor U1581 (N_1581,In_1634,In_2090);
nor U1582 (N_1582,In_2240,In_667);
nor U1583 (N_1583,In_880,In_2220);
nand U1584 (N_1584,In_1368,In_1608);
nor U1585 (N_1585,In_2161,In_908);
xor U1586 (N_1586,In_530,In_1391);
nor U1587 (N_1587,In_164,In_342);
or U1588 (N_1588,In_1771,In_50);
nor U1589 (N_1589,In_1450,In_2283);
nor U1590 (N_1590,In_920,In_1275);
and U1591 (N_1591,In_1865,In_1463);
or U1592 (N_1592,In_2235,In_1567);
or U1593 (N_1593,In_1824,In_740);
xnor U1594 (N_1594,In_2134,In_2141);
or U1595 (N_1595,In_1620,In_1012);
nor U1596 (N_1596,In_363,In_1127);
or U1597 (N_1597,In_1013,In_102);
nor U1598 (N_1598,In_1683,In_1979);
nor U1599 (N_1599,In_426,In_253);
and U1600 (N_1600,In_1452,In_883);
and U1601 (N_1601,In_306,In_1924);
and U1602 (N_1602,In_498,In_2226);
and U1603 (N_1603,In_1372,In_1431);
or U1604 (N_1604,In_1440,In_2454);
or U1605 (N_1605,In_211,In_1784);
nand U1606 (N_1606,In_2214,In_278);
nor U1607 (N_1607,In_2492,In_861);
nand U1608 (N_1608,In_2032,In_275);
nor U1609 (N_1609,In_779,In_1387);
xor U1610 (N_1610,In_1432,In_2173);
xnor U1611 (N_1611,In_2130,In_1474);
nor U1612 (N_1612,In_452,In_1724);
xnor U1613 (N_1613,In_252,In_1237);
nor U1614 (N_1614,In_583,In_1646);
or U1615 (N_1615,In_1460,In_2040);
nor U1616 (N_1616,In_1543,In_470);
xnor U1617 (N_1617,In_525,In_92);
xor U1618 (N_1618,In_1599,In_1654);
nand U1619 (N_1619,In_898,In_1104);
and U1620 (N_1620,In_167,In_409);
nand U1621 (N_1621,In_1332,In_601);
and U1622 (N_1622,In_2383,In_1656);
nor U1623 (N_1623,In_1758,In_1467);
or U1624 (N_1624,In_2491,In_1991);
nand U1625 (N_1625,In_1654,In_1449);
nand U1626 (N_1626,In_2112,In_690);
and U1627 (N_1627,In_2060,In_1601);
nor U1628 (N_1628,In_818,In_1550);
and U1629 (N_1629,In_77,In_2157);
and U1630 (N_1630,In_2442,In_2098);
and U1631 (N_1631,In_203,In_1071);
nand U1632 (N_1632,In_1580,In_2192);
nand U1633 (N_1633,In_1382,In_1968);
nor U1634 (N_1634,In_1266,In_846);
nor U1635 (N_1635,In_889,In_1849);
or U1636 (N_1636,In_1981,In_846);
and U1637 (N_1637,In_2110,In_1595);
or U1638 (N_1638,In_1673,In_1965);
and U1639 (N_1639,In_1630,In_2041);
nand U1640 (N_1640,In_2453,In_108);
and U1641 (N_1641,In_1173,In_35);
nand U1642 (N_1642,In_1708,In_2493);
or U1643 (N_1643,In_1555,In_2479);
and U1644 (N_1644,In_1714,In_167);
and U1645 (N_1645,In_2357,In_90);
and U1646 (N_1646,In_596,In_7);
or U1647 (N_1647,In_2112,In_300);
or U1648 (N_1648,In_2137,In_2082);
nor U1649 (N_1649,In_2038,In_576);
and U1650 (N_1650,In_1554,In_751);
xor U1651 (N_1651,In_601,In_2080);
and U1652 (N_1652,In_1512,In_2245);
or U1653 (N_1653,In_641,In_118);
xor U1654 (N_1654,In_875,In_2451);
and U1655 (N_1655,In_683,In_102);
or U1656 (N_1656,In_1938,In_1896);
and U1657 (N_1657,In_598,In_198);
nor U1658 (N_1658,In_2061,In_1031);
xor U1659 (N_1659,In_680,In_386);
nor U1660 (N_1660,In_207,In_211);
nand U1661 (N_1661,In_678,In_2156);
or U1662 (N_1662,In_1888,In_1205);
and U1663 (N_1663,In_1966,In_2177);
or U1664 (N_1664,In_630,In_1063);
or U1665 (N_1665,In_2062,In_2441);
or U1666 (N_1666,In_192,In_2051);
or U1667 (N_1667,In_2096,In_737);
and U1668 (N_1668,In_1068,In_1955);
nand U1669 (N_1669,In_2430,In_702);
and U1670 (N_1670,In_2306,In_155);
nand U1671 (N_1671,In_1409,In_803);
and U1672 (N_1672,In_2312,In_1222);
nand U1673 (N_1673,In_968,In_1077);
or U1674 (N_1674,In_1303,In_1476);
or U1675 (N_1675,In_1326,In_1408);
nand U1676 (N_1676,In_1815,In_1996);
nor U1677 (N_1677,In_1241,In_1417);
and U1678 (N_1678,In_81,In_2169);
nor U1679 (N_1679,In_735,In_1886);
nand U1680 (N_1680,In_1760,In_231);
and U1681 (N_1681,In_1921,In_1522);
nor U1682 (N_1682,In_1061,In_798);
and U1683 (N_1683,In_1789,In_1575);
or U1684 (N_1684,In_1831,In_1577);
nor U1685 (N_1685,In_2103,In_725);
nor U1686 (N_1686,In_587,In_1467);
nand U1687 (N_1687,In_2095,In_909);
nand U1688 (N_1688,In_1934,In_830);
and U1689 (N_1689,In_170,In_1046);
nand U1690 (N_1690,In_1708,In_789);
nor U1691 (N_1691,In_1355,In_2399);
nor U1692 (N_1692,In_628,In_1506);
and U1693 (N_1693,In_796,In_2464);
nand U1694 (N_1694,In_2169,In_2367);
nand U1695 (N_1695,In_1788,In_11);
nand U1696 (N_1696,In_607,In_240);
and U1697 (N_1697,In_459,In_377);
xor U1698 (N_1698,In_108,In_1981);
and U1699 (N_1699,In_959,In_1197);
nor U1700 (N_1700,In_1532,In_698);
nor U1701 (N_1701,In_1952,In_1297);
or U1702 (N_1702,In_2431,In_129);
or U1703 (N_1703,In_1041,In_1097);
nand U1704 (N_1704,In_1126,In_1269);
nand U1705 (N_1705,In_2250,In_2494);
and U1706 (N_1706,In_1189,In_1287);
xor U1707 (N_1707,In_2487,In_1473);
nand U1708 (N_1708,In_458,In_1879);
nand U1709 (N_1709,In_2361,In_730);
or U1710 (N_1710,In_1992,In_1890);
and U1711 (N_1711,In_1382,In_2395);
or U1712 (N_1712,In_2024,In_1225);
or U1713 (N_1713,In_1634,In_36);
nand U1714 (N_1714,In_1028,In_1898);
xnor U1715 (N_1715,In_1904,In_2057);
xnor U1716 (N_1716,In_156,In_726);
nor U1717 (N_1717,In_712,In_1158);
nand U1718 (N_1718,In_1989,In_1250);
nand U1719 (N_1719,In_175,In_1096);
nor U1720 (N_1720,In_337,In_694);
xor U1721 (N_1721,In_103,In_1435);
nand U1722 (N_1722,In_2106,In_1827);
and U1723 (N_1723,In_687,In_777);
nor U1724 (N_1724,In_1100,In_476);
or U1725 (N_1725,In_2128,In_899);
nor U1726 (N_1726,In_586,In_1012);
and U1727 (N_1727,In_1825,In_817);
xnor U1728 (N_1728,In_53,In_2358);
or U1729 (N_1729,In_522,In_2170);
and U1730 (N_1730,In_2355,In_467);
nand U1731 (N_1731,In_616,In_2007);
and U1732 (N_1732,In_304,In_601);
nand U1733 (N_1733,In_1405,In_1352);
xor U1734 (N_1734,In_1171,In_1861);
and U1735 (N_1735,In_600,In_251);
and U1736 (N_1736,In_219,In_1394);
nand U1737 (N_1737,In_720,In_607);
nor U1738 (N_1738,In_384,In_2089);
nand U1739 (N_1739,In_2368,In_2460);
nand U1740 (N_1740,In_2253,In_2345);
and U1741 (N_1741,In_1383,In_1198);
nand U1742 (N_1742,In_706,In_134);
or U1743 (N_1743,In_704,In_716);
or U1744 (N_1744,In_821,In_1473);
nor U1745 (N_1745,In_221,In_1702);
nor U1746 (N_1746,In_1858,In_96);
nand U1747 (N_1747,In_1772,In_1806);
and U1748 (N_1748,In_1954,In_1285);
or U1749 (N_1749,In_2422,In_812);
nand U1750 (N_1750,In_1232,In_287);
nor U1751 (N_1751,In_352,In_1519);
nor U1752 (N_1752,In_928,In_1594);
or U1753 (N_1753,In_2248,In_498);
and U1754 (N_1754,In_246,In_636);
nand U1755 (N_1755,In_1231,In_1299);
and U1756 (N_1756,In_612,In_1048);
nand U1757 (N_1757,In_72,In_1160);
or U1758 (N_1758,In_584,In_458);
and U1759 (N_1759,In_2047,In_492);
nand U1760 (N_1760,In_2309,In_2214);
or U1761 (N_1761,In_497,In_2207);
nor U1762 (N_1762,In_1599,In_1269);
nand U1763 (N_1763,In_685,In_1425);
xor U1764 (N_1764,In_990,In_284);
xor U1765 (N_1765,In_434,In_1190);
and U1766 (N_1766,In_613,In_1711);
or U1767 (N_1767,In_1224,In_2360);
and U1768 (N_1768,In_176,In_943);
nand U1769 (N_1769,In_1232,In_72);
nand U1770 (N_1770,In_2046,In_2143);
nor U1771 (N_1771,In_1910,In_1812);
nand U1772 (N_1772,In_1509,In_266);
and U1773 (N_1773,In_201,In_328);
and U1774 (N_1774,In_1743,In_425);
nor U1775 (N_1775,In_257,In_275);
and U1776 (N_1776,In_1250,In_1831);
nor U1777 (N_1777,In_1036,In_1181);
and U1778 (N_1778,In_1659,In_1317);
nand U1779 (N_1779,In_446,In_2069);
and U1780 (N_1780,In_1385,In_2402);
and U1781 (N_1781,In_1468,In_1571);
xnor U1782 (N_1782,In_361,In_2418);
or U1783 (N_1783,In_747,In_1853);
nor U1784 (N_1784,In_986,In_2062);
xnor U1785 (N_1785,In_1979,In_586);
and U1786 (N_1786,In_1643,In_2488);
or U1787 (N_1787,In_982,In_1947);
and U1788 (N_1788,In_2077,In_192);
and U1789 (N_1789,In_960,In_1075);
nand U1790 (N_1790,In_425,In_2022);
nand U1791 (N_1791,In_1649,In_1079);
nand U1792 (N_1792,In_202,In_328);
or U1793 (N_1793,In_1963,In_252);
or U1794 (N_1794,In_704,In_2434);
nor U1795 (N_1795,In_678,In_2003);
and U1796 (N_1796,In_188,In_1811);
and U1797 (N_1797,In_1120,In_1145);
nand U1798 (N_1798,In_431,In_1557);
nand U1799 (N_1799,In_21,In_44);
and U1800 (N_1800,In_1818,In_1535);
or U1801 (N_1801,In_819,In_660);
nand U1802 (N_1802,In_2318,In_1869);
nand U1803 (N_1803,In_1642,In_1963);
nand U1804 (N_1804,In_490,In_1160);
and U1805 (N_1805,In_2033,In_839);
xor U1806 (N_1806,In_801,In_426);
and U1807 (N_1807,In_2009,In_1957);
or U1808 (N_1808,In_180,In_2226);
nand U1809 (N_1809,In_469,In_2076);
nand U1810 (N_1810,In_1164,In_1179);
xnor U1811 (N_1811,In_2462,In_2043);
or U1812 (N_1812,In_161,In_1932);
and U1813 (N_1813,In_910,In_428);
nor U1814 (N_1814,In_2319,In_1881);
or U1815 (N_1815,In_833,In_344);
xnor U1816 (N_1816,In_1650,In_1057);
nand U1817 (N_1817,In_2101,In_563);
and U1818 (N_1818,In_1449,In_144);
xnor U1819 (N_1819,In_359,In_2009);
nand U1820 (N_1820,In_2239,In_726);
or U1821 (N_1821,In_300,In_1861);
and U1822 (N_1822,In_1915,In_1000);
and U1823 (N_1823,In_2446,In_392);
nand U1824 (N_1824,In_1986,In_1048);
or U1825 (N_1825,In_264,In_689);
xnor U1826 (N_1826,In_1491,In_394);
or U1827 (N_1827,In_314,In_404);
and U1828 (N_1828,In_2173,In_1041);
and U1829 (N_1829,In_1286,In_667);
or U1830 (N_1830,In_86,In_204);
and U1831 (N_1831,In_2072,In_1025);
and U1832 (N_1832,In_10,In_1025);
nand U1833 (N_1833,In_1080,In_1797);
nor U1834 (N_1834,In_2174,In_743);
or U1835 (N_1835,In_1475,In_334);
or U1836 (N_1836,In_1351,In_858);
or U1837 (N_1837,In_36,In_1823);
nor U1838 (N_1838,In_2412,In_2488);
xnor U1839 (N_1839,In_51,In_2470);
and U1840 (N_1840,In_955,In_865);
nor U1841 (N_1841,In_981,In_1739);
nor U1842 (N_1842,In_1244,In_2285);
and U1843 (N_1843,In_1090,In_1719);
nor U1844 (N_1844,In_1757,In_202);
and U1845 (N_1845,In_1548,In_1763);
xnor U1846 (N_1846,In_242,In_742);
nand U1847 (N_1847,In_1686,In_1015);
nor U1848 (N_1848,In_972,In_1350);
or U1849 (N_1849,In_1959,In_1585);
nor U1850 (N_1850,In_1696,In_1926);
nand U1851 (N_1851,In_1297,In_9);
or U1852 (N_1852,In_2488,In_1503);
nor U1853 (N_1853,In_2370,In_1356);
nor U1854 (N_1854,In_228,In_2073);
nand U1855 (N_1855,In_2168,In_1544);
nor U1856 (N_1856,In_1830,In_2174);
and U1857 (N_1857,In_1948,In_342);
xor U1858 (N_1858,In_458,In_1747);
nor U1859 (N_1859,In_539,In_764);
xnor U1860 (N_1860,In_1849,In_2241);
nand U1861 (N_1861,In_409,In_1638);
and U1862 (N_1862,In_323,In_1290);
nor U1863 (N_1863,In_1286,In_1126);
or U1864 (N_1864,In_748,In_2005);
nand U1865 (N_1865,In_2462,In_1627);
or U1866 (N_1866,In_153,In_1962);
and U1867 (N_1867,In_1021,In_926);
and U1868 (N_1868,In_1985,In_1414);
xor U1869 (N_1869,In_1281,In_1937);
nor U1870 (N_1870,In_1965,In_2431);
and U1871 (N_1871,In_388,In_2351);
nand U1872 (N_1872,In_1150,In_1875);
or U1873 (N_1873,In_1336,In_292);
and U1874 (N_1874,In_2108,In_1434);
xor U1875 (N_1875,In_46,In_2312);
nand U1876 (N_1876,In_777,In_1933);
nor U1877 (N_1877,In_1529,In_1639);
nand U1878 (N_1878,In_2067,In_892);
nor U1879 (N_1879,In_1233,In_936);
and U1880 (N_1880,In_885,In_630);
nor U1881 (N_1881,In_1894,In_1103);
and U1882 (N_1882,In_1163,In_2483);
and U1883 (N_1883,In_188,In_1052);
or U1884 (N_1884,In_1000,In_1458);
nand U1885 (N_1885,In_1601,In_23);
and U1886 (N_1886,In_6,In_2154);
or U1887 (N_1887,In_2183,In_2269);
or U1888 (N_1888,In_256,In_1508);
nand U1889 (N_1889,In_2466,In_1827);
or U1890 (N_1890,In_605,In_193);
and U1891 (N_1891,In_103,In_1419);
nand U1892 (N_1892,In_577,In_2197);
and U1893 (N_1893,In_731,In_1702);
and U1894 (N_1894,In_1615,In_1856);
or U1895 (N_1895,In_1966,In_461);
and U1896 (N_1896,In_1130,In_167);
nand U1897 (N_1897,In_1743,In_1386);
or U1898 (N_1898,In_951,In_441);
and U1899 (N_1899,In_1574,In_51);
xor U1900 (N_1900,In_2380,In_995);
nand U1901 (N_1901,In_789,In_1338);
nor U1902 (N_1902,In_1952,In_2065);
or U1903 (N_1903,In_829,In_556);
and U1904 (N_1904,In_442,In_861);
or U1905 (N_1905,In_2330,In_2228);
and U1906 (N_1906,In_2241,In_327);
nand U1907 (N_1907,In_497,In_315);
or U1908 (N_1908,In_2418,In_643);
nor U1909 (N_1909,In_568,In_401);
nand U1910 (N_1910,In_301,In_1597);
nand U1911 (N_1911,In_631,In_964);
nor U1912 (N_1912,In_1810,In_257);
nand U1913 (N_1913,In_1584,In_1405);
nand U1914 (N_1914,In_1062,In_169);
nor U1915 (N_1915,In_295,In_2294);
nor U1916 (N_1916,In_1914,In_535);
nor U1917 (N_1917,In_2,In_38);
or U1918 (N_1918,In_514,In_1029);
nand U1919 (N_1919,In_622,In_10);
and U1920 (N_1920,In_539,In_1291);
nor U1921 (N_1921,In_2375,In_137);
and U1922 (N_1922,In_1526,In_1649);
nand U1923 (N_1923,In_1619,In_1443);
and U1924 (N_1924,In_691,In_2164);
and U1925 (N_1925,In_2289,In_1482);
nand U1926 (N_1926,In_1124,In_268);
and U1927 (N_1927,In_55,In_655);
nor U1928 (N_1928,In_2284,In_385);
or U1929 (N_1929,In_2376,In_2414);
and U1930 (N_1930,In_1092,In_197);
nor U1931 (N_1931,In_1786,In_1102);
or U1932 (N_1932,In_2130,In_1824);
or U1933 (N_1933,In_1097,In_696);
nor U1934 (N_1934,In_548,In_428);
nand U1935 (N_1935,In_1134,In_1357);
and U1936 (N_1936,In_379,In_1536);
or U1937 (N_1937,In_1894,In_1816);
or U1938 (N_1938,In_1298,In_1428);
nand U1939 (N_1939,In_1339,In_752);
nand U1940 (N_1940,In_253,In_2345);
or U1941 (N_1941,In_1762,In_405);
nand U1942 (N_1942,In_1821,In_416);
or U1943 (N_1943,In_579,In_1621);
and U1944 (N_1944,In_1961,In_1484);
nor U1945 (N_1945,In_14,In_908);
nor U1946 (N_1946,In_2110,In_685);
nor U1947 (N_1947,In_1915,In_408);
or U1948 (N_1948,In_186,In_1759);
and U1949 (N_1949,In_1400,In_1126);
nor U1950 (N_1950,In_240,In_1641);
or U1951 (N_1951,In_62,In_1582);
or U1952 (N_1952,In_1330,In_2124);
nor U1953 (N_1953,In_2017,In_1406);
and U1954 (N_1954,In_2469,In_373);
nand U1955 (N_1955,In_174,In_1295);
and U1956 (N_1956,In_166,In_891);
nand U1957 (N_1957,In_2351,In_1502);
nand U1958 (N_1958,In_561,In_177);
nor U1959 (N_1959,In_949,In_2198);
nand U1960 (N_1960,In_1135,In_212);
or U1961 (N_1961,In_1901,In_2348);
and U1962 (N_1962,In_191,In_785);
or U1963 (N_1963,In_1,In_1031);
nor U1964 (N_1964,In_152,In_2015);
or U1965 (N_1965,In_2186,In_2488);
nand U1966 (N_1966,In_1370,In_1015);
or U1967 (N_1967,In_661,In_454);
and U1968 (N_1968,In_751,In_846);
nand U1969 (N_1969,In_1149,In_1503);
nor U1970 (N_1970,In_2164,In_396);
and U1971 (N_1971,In_2163,In_1767);
or U1972 (N_1972,In_763,In_821);
or U1973 (N_1973,In_916,In_1248);
and U1974 (N_1974,In_1357,In_1775);
nand U1975 (N_1975,In_1572,In_786);
or U1976 (N_1976,In_1403,In_433);
nor U1977 (N_1977,In_2160,In_846);
xnor U1978 (N_1978,In_1302,In_1887);
and U1979 (N_1979,In_524,In_91);
nor U1980 (N_1980,In_1220,In_564);
or U1981 (N_1981,In_1830,In_320);
or U1982 (N_1982,In_335,In_924);
and U1983 (N_1983,In_200,In_1239);
nor U1984 (N_1984,In_1636,In_530);
xnor U1985 (N_1985,In_279,In_1441);
and U1986 (N_1986,In_854,In_1800);
and U1987 (N_1987,In_2127,In_985);
and U1988 (N_1988,In_1734,In_712);
nand U1989 (N_1989,In_1328,In_2301);
nand U1990 (N_1990,In_577,In_295);
or U1991 (N_1991,In_1885,In_2213);
nand U1992 (N_1992,In_1069,In_1972);
xor U1993 (N_1993,In_1048,In_350);
nand U1994 (N_1994,In_1802,In_563);
nor U1995 (N_1995,In_1146,In_30);
nand U1996 (N_1996,In_1327,In_879);
or U1997 (N_1997,In_52,In_1585);
nor U1998 (N_1998,In_1745,In_394);
or U1999 (N_1999,In_2112,In_1427);
and U2000 (N_2000,In_1291,In_1906);
nor U2001 (N_2001,In_1790,In_2142);
or U2002 (N_2002,In_234,In_2149);
xor U2003 (N_2003,In_1713,In_1443);
nor U2004 (N_2004,In_2140,In_1129);
nand U2005 (N_2005,In_1591,In_2242);
and U2006 (N_2006,In_940,In_1132);
or U2007 (N_2007,In_2400,In_286);
or U2008 (N_2008,In_410,In_626);
and U2009 (N_2009,In_478,In_2180);
nand U2010 (N_2010,In_1686,In_346);
or U2011 (N_2011,In_1848,In_2415);
nor U2012 (N_2012,In_1318,In_2495);
nand U2013 (N_2013,In_811,In_2385);
nand U2014 (N_2014,In_1061,In_2096);
or U2015 (N_2015,In_263,In_1969);
or U2016 (N_2016,In_2110,In_14);
nand U2017 (N_2017,In_1546,In_1444);
or U2018 (N_2018,In_1100,In_841);
nor U2019 (N_2019,In_1943,In_454);
nor U2020 (N_2020,In_283,In_805);
and U2021 (N_2021,In_2473,In_1455);
and U2022 (N_2022,In_293,In_1391);
or U2023 (N_2023,In_907,In_2403);
nand U2024 (N_2024,In_2417,In_472);
nor U2025 (N_2025,In_1984,In_683);
and U2026 (N_2026,In_1338,In_165);
or U2027 (N_2027,In_1290,In_422);
nand U2028 (N_2028,In_1957,In_1860);
xor U2029 (N_2029,In_993,In_754);
or U2030 (N_2030,In_1861,In_1945);
xnor U2031 (N_2031,In_678,In_1263);
and U2032 (N_2032,In_1832,In_2123);
nand U2033 (N_2033,In_1410,In_180);
or U2034 (N_2034,In_1286,In_1213);
xor U2035 (N_2035,In_689,In_105);
nor U2036 (N_2036,In_1306,In_1264);
and U2037 (N_2037,In_1749,In_606);
nand U2038 (N_2038,In_1744,In_2054);
nand U2039 (N_2039,In_690,In_1840);
nand U2040 (N_2040,In_74,In_106);
or U2041 (N_2041,In_427,In_1640);
nor U2042 (N_2042,In_950,In_2118);
and U2043 (N_2043,In_1874,In_1904);
and U2044 (N_2044,In_2093,In_1379);
nand U2045 (N_2045,In_2022,In_937);
nor U2046 (N_2046,In_1698,In_1816);
nor U2047 (N_2047,In_1317,In_1051);
nor U2048 (N_2048,In_2293,In_2445);
nand U2049 (N_2049,In_878,In_1002);
nand U2050 (N_2050,In_1635,In_1893);
or U2051 (N_2051,In_545,In_1132);
nand U2052 (N_2052,In_901,In_1933);
and U2053 (N_2053,In_732,In_1247);
nor U2054 (N_2054,In_2237,In_198);
nand U2055 (N_2055,In_1253,In_2422);
and U2056 (N_2056,In_1212,In_1295);
xnor U2057 (N_2057,In_1169,In_1516);
or U2058 (N_2058,In_2373,In_431);
nor U2059 (N_2059,In_842,In_494);
nand U2060 (N_2060,In_1015,In_587);
and U2061 (N_2061,In_1840,In_1945);
or U2062 (N_2062,In_113,In_994);
nor U2063 (N_2063,In_1009,In_552);
or U2064 (N_2064,In_1624,In_1958);
and U2065 (N_2065,In_941,In_467);
and U2066 (N_2066,In_1844,In_1149);
nand U2067 (N_2067,In_2136,In_715);
and U2068 (N_2068,In_1375,In_309);
nand U2069 (N_2069,In_896,In_1533);
nor U2070 (N_2070,In_976,In_1980);
xor U2071 (N_2071,In_1034,In_420);
nand U2072 (N_2072,In_269,In_2055);
xor U2073 (N_2073,In_864,In_1635);
nor U2074 (N_2074,In_1212,In_125);
nand U2075 (N_2075,In_1326,In_2360);
and U2076 (N_2076,In_217,In_816);
or U2077 (N_2077,In_433,In_1217);
nor U2078 (N_2078,In_235,In_2454);
nand U2079 (N_2079,In_2456,In_1655);
nand U2080 (N_2080,In_1179,In_1119);
nor U2081 (N_2081,In_2337,In_1013);
nor U2082 (N_2082,In_794,In_39);
or U2083 (N_2083,In_1085,In_487);
nor U2084 (N_2084,In_1191,In_1598);
nand U2085 (N_2085,In_1760,In_259);
nand U2086 (N_2086,In_2267,In_1729);
nor U2087 (N_2087,In_836,In_2422);
nor U2088 (N_2088,In_1334,In_1728);
or U2089 (N_2089,In_564,In_189);
nor U2090 (N_2090,In_1340,In_390);
nand U2091 (N_2091,In_1125,In_189);
nor U2092 (N_2092,In_2060,In_1249);
and U2093 (N_2093,In_2414,In_869);
xnor U2094 (N_2094,In_1323,In_372);
and U2095 (N_2095,In_736,In_193);
or U2096 (N_2096,In_17,In_739);
nor U2097 (N_2097,In_2153,In_1873);
nand U2098 (N_2098,In_1381,In_1587);
nand U2099 (N_2099,In_1832,In_455);
nor U2100 (N_2100,In_479,In_1442);
nor U2101 (N_2101,In_1217,In_2220);
nand U2102 (N_2102,In_614,In_2484);
nand U2103 (N_2103,In_118,In_2239);
and U2104 (N_2104,In_584,In_1158);
and U2105 (N_2105,In_2312,In_1036);
and U2106 (N_2106,In_1139,In_421);
nand U2107 (N_2107,In_2162,In_2369);
nor U2108 (N_2108,In_1772,In_2075);
or U2109 (N_2109,In_2403,In_2005);
and U2110 (N_2110,In_829,In_504);
nor U2111 (N_2111,In_1464,In_2138);
or U2112 (N_2112,In_186,In_1177);
nor U2113 (N_2113,In_2287,In_189);
nand U2114 (N_2114,In_1846,In_2059);
nand U2115 (N_2115,In_326,In_918);
xnor U2116 (N_2116,In_1184,In_1674);
or U2117 (N_2117,In_233,In_1653);
nand U2118 (N_2118,In_1678,In_1030);
and U2119 (N_2119,In_1550,In_1464);
and U2120 (N_2120,In_39,In_2025);
or U2121 (N_2121,In_2415,In_1081);
nor U2122 (N_2122,In_1032,In_247);
nand U2123 (N_2123,In_1869,In_188);
nand U2124 (N_2124,In_2204,In_1766);
nor U2125 (N_2125,In_201,In_115);
or U2126 (N_2126,In_1626,In_1328);
or U2127 (N_2127,In_158,In_948);
and U2128 (N_2128,In_1492,In_1183);
xnor U2129 (N_2129,In_236,In_1839);
nor U2130 (N_2130,In_726,In_1735);
nor U2131 (N_2131,In_900,In_1922);
or U2132 (N_2132,In_232,In_66);
or U2133 (N_2133,In_1722,In_528);
or U2134 (N_2134,In_1520,In_1308);
and U2135 (N_2135,In_1156,In_1198);
nor U2136 (N_2136,In_2223,In_1577);
nor U2137 (N_2137,In_1128,In_132);
and U2138 (N_2138,In_300,In_1200);
or U2139 (N_2139,In_74,In_115);
or U2140 (N_2140,In_2074,In_1155);
xnor U2141 (N_2141,In_809,In_986);
xnor U2142 (N_2142,In_2074,In_1665);
nand U2143 (N_2143,In_2216,In_1944);
nand U2144 (N_2144,In_451,In_1663);
xnor U2145 (N_2145,In_475,In_1525);
xor U2146 (N_2146,In_1195,In_2199);
and U2147 (N_2147,In_963,In_627);
nand U2148 (N_2148,In_767,In_787);
nand U2149 (N_2149,In_80,In_1377);
or U2150 (N_2150,In_1602,In_328);
xor U2151 (N_2151,In_2442,In_1252);
and U2152 (N_2152,In_1081,In_703);
nand U2153 (N_2153,In_2409,In_1070);
or U2154 (N_2154,In_822,In_1522);
and U2155 (N_2155,In_924,In_312);
nand U2156 (N_2156,In_905,In_1739);
or U2157 (N_2157,In_1241,In_1243);
nand U2158 (N_2158,In_2355,In_231);
and U2159 (N_2159,In_48,In_64);
nor U2160 (N_2160,In_1924,In_1321);
or U2161 (N_2161,In_1981,In_2110);
nor U2162 (N_2162,In_1342,In_257);
or U2163 (N_2163,In_634,In_1368);
nor U2164 (N_2164,In_2036,In_451);
and U2165 (N_2165,In_898,In_2339);
and U2166 (N_2166,In_1591,In_2193);
nor U2167 (N_2167,In_2400,In_2362);
nand U2168 (N_2168,In_370,In_2496);
and U2169 (N_2169,In_1450,In_913);
nor U2170 (N_2170,In_921,In_294);
nand U2171 (N_2171,In_2488,In_324);
nor U2172 (N_2172,In_1506,In_1538);
nor U2173 (N_2173,In_1764,In_1199);
and U2174 (N_2174,In_2093,In_1603);
nand U2175 (N_2175,In_265,In_1421);
or U2176 (N_2176,In_2341,In_2436);
or U2177 (N_2177,In_883,In_2096);
nor U2178 (N_2178,In_1235,In_1567);
and U2179 (N_2179,In_1217,In_371);
nand U2180 (N_2180,In_2349,In_2384);
xnor U2181 (N_2181,In_239,In_188);
nor U2182 (N_2182,In_1742,In_51);
nand U2183 (N_2183,In_413,In_2254);
xor U2184 (N_2184,In_1889,In_1956);
nand U2185 (N_2185,In_2015,In_1931);
and U2186 (N_2186,In_214,In_772);
nand U2187 (N_2187,In_125,In_1418);
nor U2188 (N_2188,In_1486,In_30);
nand U2189 (N_2189,In_1102,In_153);
nor U2190 (N_2190,In_1264,In_1058);
nor U2191 (N_2191,In_1162,In_963);
nand U2192 (N_2192,In_1585,In_2269);
or U2193 (N_2193,In_695,In_901);
nor U2194 (N_2194,In_1777,In_1392);
or U2195 (N_2195,In_2023,In_657);
or U2196 (N_2196,In_1682,In_839);
nor U2197 (N_2197,In_1231,In_504);
and U2198 (N_2198,In_466,In_1624);
or U2199 (N_2199,In_1776,In_374);
nand U2200 (N_2200,In_694,In_1867);
and U2201 (N_2201,In_1245,In_928);
or U2202 (N_2202,In_755,In_601);
nor U2203 (N_2203,In_1925,In_2294);
nand U2204 (N_2204,In_124,In_650);
nor U2205 (N_2205,In_1773,In_657);
nand U2206 (N_2206,In_2216,In_312);
nor U2207 (N_2207,In_130,In_1433);
and U2208 (N_2208,In_2057,In_1720);
or U2209 (N_2209,In_286,In_2014);
nor U2210 (N_2210,In_59,In_1977);
nand U2211 (N_2211,In_2117,In_1138);
and U2212 (N_2212,In_518,In_1792);
xnor U2213 (N_2213,In_2352,In_1239);
nor U2214 (N_2214,In_1198,In_2048);
xor U2215 (N_2215,In_1972,In_984);
and U2216 (N_2216,In_2283,In_230);
nand U2217 (N_2217,In_2264,In_54);
and U2218 (N_2218,In_1282,In_1005);
nor U2219 (N_2219,In_1957,In_2176);
or U2220 (N_2220,In_1118,In_1959);
or U2221 (N_2221,In_857,In_834);
xor U2222 (N_2222,In_1735,In_1319);
and U2223 (N_2223,In_2206,In_1479);
or U2224 (N_2224,In_1870,In_1092);
nor U2225 (N_2225,In_1318,In_2122);
and U2226 (N_2226,In_1580,In_527);
and U2227 (N_2227,In_1142,In_2005);
nor U2228 (N_2228,In_1710,In_821);
nand U2229 (N_2229,In_1684,In_308);
nor U2230 (N_2230,In_33,In_2217);
or U2231 (N_2231,In_256,In_1956);
and U2232 (N_2232,In_1554,In_863);
nand U2233 (N_2233,In_882,In_372);
nor U2234 (N_2234,In_823,In_1012);
nand U2235 (N_2235,In_1539,In_197);
nand U2236 (N_2236,In_1518,In_785);
nand U2237 (N_2237,In_2285,In_2350);
or U2238 (N_2238,In_965,In_2);
or U2239 (N_2239,In_998,In_2218);
and U2240 (N_2240,In_2300,In_293);
and U2241 (N_2241,In_412,In_1958);
xor U2242 (N_2242,In_1764,In_2392);
nor U2243 (N_2243,In_2130,In_293);
and U2244 (N_2244,In_2319,In_999);
and U2245 (N_2245,In_227,In_1840);
nand U2246 (N_2246,In_394,In_896);
or U2247 (N_2247,In_2298,In_656);
nand U2248 (N_2248,In_660,In_2163);
and U2249 (N_2249,In_1843,In_1900);
nand U2250 (N_2250,In_1469,In_1866);
nor U2251 (N_2251,In_1154,In_1063);
nor U2252 (N_2252,In_1685,In_81);
nor U2253 (N_2253,In_1474,In_279);
or U2254 (N_2254,In_340,In_1397);
nand U2255 (N_2255,In_1369,In_1023);
or U2256 (N_2256,In_215,In_2246);
nand U2257 (N_2257,In_979,In_291);
xnor U2258 (N_2258,In_803,In_1849);
nor U2259 (N_2259,In_1194,In_1979);
nand U2260 (N_2260,In_1270,In_373);
or U2261 (N_2261,In_2241,In_1695);
xnor U2262 (N_2262,In_1652,In_1629);
nor U2263 (N_2263,In_11,In_2334);
or U2264 (N_2264,In_1322,In_1158);
and U2265 (N_2265,In_1370,In_448);
xor U2266 (N_2266,In_17,In_20);
nand U2267 (N_2267,In_2165,In_731);
nand U2268 (N_2268,In_192,In_394);
nand U2269 (N_2269,In_1190,In_51);
nor U2270 (N_2270,In_265,In_1300);
or U2271 (N_2271,In_293,In_1362);
nand U2272 (N_2272,In_936,In_622);
nor U2273 (N_2273,In_932,In_1654);
nor U2274 (N_2274,In_50,In_973);
and U2275 (N_2275,In_1095,In_1866);
nand U2276 (N_2276,In_2241,In_1143);
nand U2277 (N_2277,In_2295,In_1526);
nor U2278 (N_2278,In_1963,In_732);
or U2279 (N_2279,In_332,In_1964);
or U2280 (N_2280,In_1864,In_320);
or U2281 (N_2281,In_141,In_1564);
and U2282 (N_2282,In_1755,In_915);
and U2283 (N_2283,In_2483,In_1202);
nand U2284 (N_2284,In_856,In_2222);
nor U2285 (N_2285,In_326,In_867);
nor U2286 (N_2286,In_2020,In_1456);
and U2287 (N_2287,In_1114,In_344);
and U2288 (N_2288,In_1689,In_2173);
or U2289 (N_2289,In_1916,In_173);
or U2290 (N_2290,In_1879,In_1912);
and U2291 (N_2291,In_2232,In_376);
xnor U2292 (N_2292,In_2099,In_1458);
or U2293 (N_2293,In_2085,In_1126);
nor U2294 (N_2294,In_1432,In_449);
xor U2295 (N_2295,In_1481,In_870);
nor U2296 (N_2296,In_1463,In_1573);
nand U2297 (N_2297,In_1031,In_1301);
and U2298 (N_2298,In_191,In_1359);
xnor U2299 (N_2299,In_816,In_2358);
and U2300 (N_2300,In_1106,In_242);
nand U2301 (N_2301,In_1244,In_1037);
nand U2302 (N_2302,In_2489,In_2232);
or U2303 (N_2303,In_1951,In_509);
and U2304 (N_2304,In_866,In_1994);
and U2305 (N_2305,In_1506,In_2369);
and U2306 (N_2306,In_229,In_2088);
or U2307 (N_2307,In_604,In_2245);
or U2308 (N_2308,In_2417,In_359);
xnor U2309 (N_2309,In_2007,In_1061);
or U2310 (N_2310,In_1820,In_1768);
or U2311 (N_2311,In_1120,In_2140);
or U2312 (N_2312,In_487,In_1735);
nor U2313 (N_2313,In_1526,In_651);
or U2314 (N_2314,In_1230,In_2282);
nand U2315 (N_2315,In_842,In_433);
nor U2316 (N_2316,In_1163,In_886);
nor U2317 (N_2317,In_1167,In_1356);
xnor U2318 (N_2318,In_2060,In_1494);
or U2319 (N_2319,In_1567,In_815);
or U2320 (N_2320,In_1522,In_2067);
nand U2321 (N_2321,In_822,In_660);
nand U2322 (N_2322,In_1597,In_2370);
xor U2323 (N_2323,In_1502,In_1657);
nand U2324 (N_2324,In_2087,In_2199);
xor U2325 (N_2325,In_439,In_1188);
nor U2326 (N_2326,In_393,In_860);
xor U2327 (N_2327,In_424,In_1076);
or U2328 (N_2328,In_2169,In_1308);
nor U2329 (N_2329,In_1623,In_214);
nor U2330 (N_2330,In_2486,In_1862);
or U2331 (N_2331,In_772,In_779);
nor U2332 (N_2332,In_1533,In_535);
and U2333 (N_2333,In_2412,In_1010);
nor U2334 (N_2334,In_2321,In_858);
nand U2335 (N_2335,In_13,In_1492);
xnor U2336 (N_2336,In_2374,In_271);
or U2337 (N_2337,In_1817,In_2165);
or U2338 (N_2338,In_2376,In_1529);
and U2339 (N_2339,In_2254,In_1404);
or U2340 (N_2340,In_2231,In_2076);
nand U2341 (N_2341,In_2474,In_655);
or U2342 (N_2342,In_277,In_701);
and U2343 (N_2343,In_1571,In_1356);
xor U2344 (N_2344,In_552,In_2410);
nor U2345 (N_2345,In_927,In_2440);
or U2346 (N_2346,In_2262,In_1758);
nor U2347 (N_2347,In_836,In_748);
xnor U2348 (N_2348,In_1703,In_661);
nor U2349 (N_2349,In_2327,In_1452);
or U2350 (N_2350,In_1116,In_2232);
or U2351 (N_2351,In_2098,In_377);
and U2352 (N_2352,In_779,In_287);
xnor U2353 (N_2353,In_1467,In_1031);
and U2354 (N_2354,In_2349,In_2146);
nor U2355 (N_2355,In_2108,In_763);
nand U2356 (N_2356,In_2177,In_1963);
and U2357 (N_2357,In_711,In_2214);
and U2358 (N_2358,In_513,In_341);
xnor U2359 (N_2359,In_849,In_735);
nand U2360 (N_2360,In_1557,In_1717);
or U2361 (N_2361,In_2184,In_2230);
or U2362 (N_2362,In_1069,In_839);
or U2363 (N_2363,In_1960,In_1945);
and U2364 (N_2364,In_1855,In_2030);
nand U2365 (N_2365,In_19,In_962);
nand U2366 (N_2366,In_2009,In_770);
or U2367 (N_2367,In_167,In_1008);
nor U2368 (N_2368,In_1907,In_285);
nand U2369 (N_2369,In_242,In_797);
nand U2370 (N_2370,In_2264,In_2209);
and U2371 (N_2371,In_1413,In_953);
nand U2372 (N_2372,In_2038,In_2403);
nand U2373 (N_2373,In_508,In_850);
and U2374 (N_2374,In_903,In_2406);
or U2375 (N_2375,In_217,In_2157);
xnor U2376 (N_2376,In_64,In_1735);
or U2377 (N_2377,In_1838,In_443);
xnor U2378 (N_2378,In_567,In_978);
nand U2379 (N_2379,In_1946,In_1761);
xnor U2380 (N_2380,In_472,In_1981);
nor U2381 (N_2381,In_1137,In_1301);
and U2382 (N_2382,In_1500,In_2342);
nor U2383 (N_2383,In_1029,In_2374);
nand U2384 (N_2384,In_1175,In_68);
nand U2385 (N_2385,In_1119,In_1879);
or U2386 (N_2386,In_255,In_1129);
and U2387 (N_2387,In_844,In_1596);
or U2388 (N_2388,In_1348,In_1909);
nor U2389 (N_2389,In_2097,In_1525);
nor U2390 (N_2390,In_661,In_664);
nor U2391 (N_2391,In_1197,In_828);
or U2392 (N_2392,In_1251,In_465);
or U2393 (N_2393,In_1154,In_1172);
nor U2394 (N_2394,In_1629,In_1923);
nand U2395 (N_2395,In_1193,In_166);
or U2396 (N_2396,In_2452,In_507);
and U2397 (N_2397,In_1159,In_448);
nand U2398 (N_2398,In_2303,In_268);
nor U2399 (N_2399,In_576,In_1065);
and U2400 (N_2400,In_158,In_1369);
or U2401 (N_2401,In_145,In_327);
nor U2402 (N_2402,In_1091,In_83);
or U2403 (N_2403,In_1467,In_415);
and U2404 (N_2404,In_1794,In_162);
xor U2405 (N_2405,In_401,In_793);
nand U2406 (N_2406,In_1901,In_1567);
and U2407 (N_2407,In_1192,In_343);
or U2408 (N_2408,In_634,In_1700);
and U2409 (N_2409,In_1742,In_1941);
and U2410 (N_2410,In_815,In_1653);
nor U2411 (N_2411,In_2068,In_477);
nor U2412 (N_2412,In_2372,In_1250);
and U2413 (N_2413,In_2065,In_866);
and U2414 (N_2414,In_1307,In_878);
or U2415 (N_2415,In_87,In_2064);
or U2416 (N_2416,In_774,In_1604);
nor U2417 (N_2417,In_938,In_2324);
nor U2418 (N_2418,In_1857,In_1464);
or U2419 (N_2419,In_749,In_349);
and U2420 (N_2420,In_1519,In_215);
nor U2421 (N_2421,In_608,In_2079);
nor U2422 (N_2422,In_1299,In_1143);
xnor U2423 (N_2423,In_1736,In_1902);
or U2424 (N_2424,In_1512,In_1568);
or U2425 (N_2425,In_663,In_2303);
nand U2426 (N_2426,In_1588,In_1982);
xnor U2427 (N_2427,In_896,In_2092);
xor U2428 (N_2428,In_939,In_1800);
nand U2429 (N_2429,In_16,In_405);
nand U2430 (N_2430,In_2073,In_1293);
nand U2431 (N_2431,In_1676,In_1311);
or U2432 (N_2432,In_686,In_1881);
and U2433 (N_2433,In_2414,In_184);
and U2434 (N_2434,In_155,In_1265);
nor U2435 (N_2435,In_369,In_264);
nor U2436 (N_2436,In_1033,In_790);
nand U2437 (N_2437,In_2093,In_1811);
and U2438 (N_2438,In_789,In_2396);
nor U2439 (N_2439,In_290,In_1981);
nor U2440 (N_2440,In_204,In_2208);
xor U2441 (N_2441,In_1094,In_1703);
nand U2442 (N_2442,In_1662,In_447);
nor U2443 (N_2443,In_2114,In_2040);
or U2444 (N_2444,In_176,In_2335);
nand U2445 (N_2445,In_2325,In_1120);
or U2446 (N_2446,In_242,In_1928);
or U2447 (N_2447,In_2057,In_2390);
nand U2448 (N_2448,In_1912,In_533);
nand U2449 (N_2449,In_238,In_1920);
xnor U2450 (N_2450,In_2143,In_1611);
or U2451 (N_2451,In_1172,In_2041);
and U2452 (N_2452,In_31,In_1413);
nor U2453 (N_2453,In_523,In_1911);
and U2454 (N_2454,In_39,In_1313);
nor U2455 (N_2455,In_192,In_1890);
xnor U2456 (N_2456,In_1767,In_307);
nand U2457 (N_2457,In_1678,In_422);
or U2458 (N_2458,In_1034,In_1871);
or U2459 (N_2459,In_419,In_2236);
nand U2460 (N_2460,In_490,In_84);
and U2461 (N_2461,In_579,In_1093);
and U2462 (N_2462,In_94,In_1698);
xnor U2463 (N_2463,In_164,In_77);
nor U2464 (N_2464,In_807,In_206);
and U2465 (N_2465,In_1889,In_573);
or U2466 (N_2466,In_2367,In_2192);
or U2467 (N_2467,In_808,In_2127);
or U2468 (N_2468,In_1286,In_1117);
or U2469 (N_2469,In_1982,In_42);
xnor U2470 (N_2470,In_667,In_2175);
or U2471 (N_2471,In_2479,In_2130);
nor U2472 (N_2472,In_342,In_889);
nand U2473 (N_2473,In_990,In_583);
nor U2474 (N_2474,In_423,In_2295);
nand U2475 (N_2475,In_919,In_383);
or U2476 (N_2476,In_268,In_855);
or U2477 (N_2477,In_2089,In_2288);
and U2478 (N_2478,In_2079,In_248);
and U2479 (N_2479,In_256,In_735);
or U2480 (N_2480,In_477,In_1952);
xnor U2481 (N_2481,In_1031,In_1011);
nor U2482 (N_2482,In_1028,In_120);
nor U2483 (N_2483,In_2054,In_1336);
and U2484 (N_2484,In_1930,In_1400);
and U2485 (N_2485,In_1056,In_1373);
nor U2486 (N_2486,In_1331,In_548);
nand U2487 (N_2487,In_2417,In_888);
or U2488 (N_2488,In_721,In_960);
or U2489 (N_2489,In_744,In_1185);
nand U2490 (N_2490,In_856,In_1037);
and U2491 (N_2491,In_1086,In_2479);
and U2492 (N_2492,In_771,In_1600);
xnor U2493 (N_2493,In_1938,In_1802);
or U2494 (N_2494,In_813,In_754);
or U2495 (N_2495,In_180,In_1698);
nand U2496 (N_2496,In_44,In_2362);
nor U2497 (N_2497,In_1378,In_283);
nand U2498 (N_2498,In_1351,In_5);
or U2499 (N_2499,In_1504,In_105);
and U2500 (N_2500,In_1809,In_1964);
or U2501 (N_2501,In_1548,In_2068);
or U2502 (N_2502,In_1854,In_837);
nand U2503 (N_2503,In_1214,In_1117);
nor U2504 (N_2504,In_39,In_847);
or U2505 (N_2505,In_1988,In_380);
nand U2506 (N_2506,In_1671,In_2223);
nand U2507 (N_2507,In_975,In_1362);
or U2508 (N_2508,In_1924,In_136);
or U2509 (N_2509,In_234,In_1093);
nor U2510 (N_2510,In_1409,In_590);
or U2511 (N_2511,In_269,In_1223);
xor U2512 (N_2512,In_2397,In_2086);
nor U2513 (N_2513,In_568,In_1906);
xor U2514 (N_2514,In_2343,In_506);
nor U2515 (N_2515,In_669,In_1824);
or U2516 (N_2516,In_481,In_337);
nand U2517 (N_2517,In_2435,In_21);
and U2518 (N_2518,In_1077,In_1268);
or U2519 (N_2519,In_2164,In_1191);
xnor U2520 (N_2520,In_2440,In_528);
or U2521 (N_2521,In_1178,In_834);
xor U2522 (N_2522,In_2133,In_681);
nor U2523 (N_2523,In_1188,In_2371);
nand U2524 (N_2524,In_667,In_101);
nor U2525 (N_2525,In_1886,In_640);
nor U2526 (N_2526,In_2404,In_1099);
and U2527 (N_2527,In_766,In_104);
and U2528 (N_2528,In_2032,In_2002);
nand U2529 (N_2529,In_1494,In_466);
nor U2530 (N_2530,In_624,In_613);
xnor U2531 (N_2531,In_585,In_297);
and U2532 (N_2532,In_2167,In_687);
nor U2533 (N_2533,In_1667,In_1258);
or U2534 (N_2534,In_437,In_978);
or U2535 (N_2535,In_2421,In_1280);
xor U2536 (N_2536,In_812,In_23);
nand U2537 (N_2537,In_239,In_2005);
nor U2538 (N_2538,In_1776,In_384);
and U2539 (N_2539,In_2369,In_1846);
or U2540 (N_2540,In_1087,In_842);
nand U2541 (N_2541,In_1853,In_2494);
or U2542 (N_2542,In_923,In_2071);
and U2543 (N_2543,In_2194,In_946);
nor U2544 (N_2544,In_2319,In_1913);
nand U2545 (N_2545,In_514,In_311);
and U2546 (N_2546,In_1153,In_2405);
nand U2547 (N_2547,In_1151,In_540);
nor U2548 (N_2548,In_407,In_2301);
or U2549 (N_2549,In_262,In_735);
or U2550 (N_2550,In_206,In_527);
nand U2551 (N_2551,In_572,In_1879);
nor U2552 (N_2552,In_155,In_527);
or U2553 (N_2553,In_524,In_1628);
or U2554 (N_2554,In_1921,In_1718);
or U2555 (N_2555,In_40,In_1811);
nor U2556 (N_2556,In_2244,In_1282);
nand U2557 (N_2557,In_1509,In_951);
xnor U2558 (N_2558,In_300,In_2120);
nor U2559 (N_2559,In_1277,In_1294);
xor U2560 (N_2560,In_1815,In_743);
nor U2561 (N_2561,In_2455,In_2421);
and U2562 (N_2562,In_1195,In_712);
or U2563 (N_2563,In_1337,In_1986);
xor U2564 (N_2564,In_2372,In_1095);
nand U2565 (N_2565,In_628,In_273);
nor U2566 (N_2566,In_851,In_1778);
and U2567 (N_2567,In_1633,In_1767);
nand U2568 (N_2568,In_1393,In_1941);
or U2569 (N_2569,In_837,In_991);
nand U2570 (N_2570,In_2449,In_1605);
nand U2571 (N_2571,In_2152,In_835);
nor U2572 (N_2572,In_2332,In_741);
or U2573 (N_2573,In_2304,In_2361);
nor U2574 (N_2574,In_1906,In_281);
and U2575 (N_2575,In_639,In_574);
and U2576 (N_2576,In_931,In_361);
or U2577 (N_2577,In_1421,In_1288);
nand U2578 (N_2578,In_86,In_1584);
or U2579 (N_2579,In_1721,In_1175);
or U2580 (N_2580,In_137,In_433);
nand U2581 (N_2581,In_1226,In_597);
nor U2582 (N_2582,In_442,In_1133);
nand U2583 (N_2583,In_657,In_1289);
nand U2584 (N_2584,In_752,In_2112);
and U2585 (N_2585,In_2217,In_1310);
xnor U2586 (N_2586,In_1465,In_957);
nor U2587 (N_2587,In_1726,In_555);
and U2588 (N_2588,In_727,In_341);
and U2589 (N_2589,In_1494,In_2318);
nor U2590 (N_2590,In_889,In_1863);
nor U2591 (N_2591,In_2327,In_2167);
nand U2592 (N_2592,In_2203,In_778);
or U2593 (N_2593,In_1600,In_1377);
or U2594 (N_2594,In_1914,In_724);
and U2595 (N_2595,In_2253,In_184);
nor U2596 (N_2596,In_604,In_1381);
xor U2597 (N_2597,In_189,In_2437);
or U2598 (N_2598,In_167,In_948);
or U2599 (N_2599,In_5,In_1040);
nor U2600 (N_2600,In_32,In_2481);
or U2601 (N_2601,In_1943,In_996);
nor U2602 (N_2602,In_40,In_430);
and U2603 (N_2603,In_132,In_177);
nor U2604 (N_2604,In_2371,In_489);
xnor U2605 (N_2605,In_2027,In_750);
nand U2606 (N_2606,In_1685,In_1341);
nand U2607 (N_2607,In_622,In_1625);
or U2608 (N_2608,In_241,In_460);
xor U2609 (N_2609,In_2398,In_2061);
or U2610 (N_2610,In_1895,In_596);
or U2611 (N_2611,In_1298,In_1672);
or U2612 (N_2612,In_1815,In_766);
and U2613 (N_2613,In_1166,In_1273);
nor U2614 (N_2614,In_1446,In_2306);
and U2615 (N_2615,In_804,In_392);
nand U2616 (N_2616,In_2032,In_1861);
nand U2617 (N_2617,In_131,In_1464);
or U2618 (N_2618,In_622,In_1051);
nor U2619 (N_2619,In_550,In_2410);
xnor U2620 (N_2620,In_390,In_2078);
nand U2621 (N_2621,In_1341,In_1505);
nor U2622 (N_2622,In_1557,In_628);
nor U2623 (N_2623,In_1817,In_1380);
nand U2624 (N_2624,In_1063,In_6);
or U2625 (N_2625,In_145,In_906);
nor U2626 (N_2626,In_940,In_362);
nor U2627 (N_2627,In_1075,In_1926);
nor U2628 (N_2628,In_298,In_1349);
or U2629 (N_2629,In_1013,In_2390);
nand U2630 (N_2630,In_702,In_1888);
xor U2631 (N_2631,In_471,In_2498);
and U2632 (N_2632,In_458,In_1686);
and U2633 (N_2633,In_2420,In_1075);
and U2634 (N_2634,In_2196,In_261);
and U2635 (N_2635,In_1314,In_1811);
and U2636 (N_2636,In_483,In_553);
nand U2637 (N_2637,In_42,In_1118);
xor U2638 (N_2638,In_868,In_29);
or U2639 (N_2639,In_2155,In_2228);
xor U2640 (N_2640,In_1388,In_2120);
and U2641 (N_2641,In_309,In_307);
and U2642 (N_2642,In_1917,In_2450);
nor U2643 (N_2643,In_1065,In_2439);
and U2644 (N_2644,In_1324,In_722);
or U2645 (N_2645,In_2176,In_1112);
and U2646 (N_2646,In_926,In_1115);
and U2647 (N_2647,In_1698,In_1267);
and U2648 (N_2648,In_407,In_2256);
or U2649 (N_2649,In_1022,In_1104);
nand U2650 (N_2650,In_1764,In_1132);
or U2651 (N_2651,In_149,In_1929);
nand U2652 (N_2652,In_1730,In_1021);
nand U2653 (N_2653,In_1467,In_1837);
or U2654 (N_2654,In_1451,In_714);
and U2655 (N_2655,In_1801,In_665);
xor U2656 (N_2656,In_1133,In_147);
nand U2657 (N_2657,In_1469,In_1462);
and U2658 (N_2658,In_2395,In_1824);
and U2659 (N_2659,In_1596,In_95);
xor U2660 (N_2660,In_41,In_423);
or U2661 (N_2661,In_1937,In_1234);
xnor U2662 (N_2662,In_855,In_200);
nor U2663 (N_2663,In_1534,In_1067);
or U2664 (N_2664,In_43,In_2011);
nor U2665 (N_2665,In_521,In_1561);
and U2666 (N_2666,In_919,In_1528);
nand U2667 (N_2667,In_2160,In_1150);
or U2668 (N_2668,In_1010,In_830);
and U2669 (N_2669,In_181,In_2347);
xor U2670 (N_2670,In_2115,In_27);
xor U2671 (N_2671,In_798,In_2469);
nand U2672 (N_2672,In_894,In_822);
and U2673 (N_2673,In_2266,In_1231);
and U2674 (N_2674,In_1598,In_1977);
nor U2675 (N_2675,In_448,In_428);
xor U2676 (N_2676,In_636,In_1800);
and U2677 (N_2677,In_185,In_1540);
nor U2678 (N_2678,In_488,In_951);
and U2679 (N_2679,In_877,In_1802);
or U2680 (N_2680,In_806,In_777);
xor U2681 (N_2681,In_1812,In_860);
or U2682 (N_2682,In_2390,In_63);
xor U2683 (N_2683,In_483,In_314);
nand U2684 (N_2684,In_1371,In_794);
and U2685 (N_2685,In_836,In_2458);
and U2686 (N_2686,In_338,In_443);
nand U2687 (N_2687,In_1670,In_2490);
nor U2688 (N_2688,In_1828,In_1673);
nor U2689 (N_2689,In_1004,In_1636);
and U2690 (N_2690,In_1719,In_1820);
xor U2691 (N_2691,In_2259,In_2003);
and U2692 (N_2692,In_1260,In_405);
xor U2693 (N_2693,In_374,In_1408);
nor U2694 (N_2694,In_1820,In_1109);
or U2695 (N_2695,In_1666,In_2343);
nor U2696 (N_2696,In_2100,In_468);
nor U2697 (N_2697,In_541,In_2490);
and U2698 (N_2698,In_2077,In_855);
or U2699 (N_2699,In_1681,In_232);
and U2700 (N_2700,In_177,In_1190);
xor U2701 (N_2701,In_725,In_2044);
and U2702 (N_2702,In_1740,In_2238);
nand U2703 (N_2703,In_1932,In_1779);
nor U2704 (N_2704,In_367,In_215);
nand U2705 (N_2705,In_700,In_1118);
nand U2706 (N_2706,In_1087,In_2491);
and U2707 (N_2707,In_1762,In_11);
and U2708 (N_2708,In_2161,In_2232);
nor U2709 (N_2709,In_2374,In_2101);
or U2710 (N_2710,In_2313,In_1096);
xnor U2711 (N_2711,In_2309,In_1306);
and U2712 (N_2712,In_206,In_1331);
or U2713 (N_2713,In_2228,In_1312);
nand U2714 (N_2714,In_2130,In_933);
nor U2715 (N_2715,In_1052,In_2117);
nor U2716 (N_2716,In_1101,In_642);
nor U2717 (N_2717,In_14,In_2323);
nand U2718 (N_2718,In_1747,In_522);
and U2719 (N_2719,In_6,In_732);
or U2720 (N_2720,In_1907,In_1500);
nand U2721 (N_2721,In_1821,In_1142);
and U2722 (N_2722,In_1786,In_528);
or U2723 (N_2723,In_71,In_2222);
or U2724 (N_2724,In_2385,In_48);
nor U2725 (N_2725,In_2286,In_2354);
and U2726 (N_2726,In_823,In_855);
nand U2727 (N_2727,In_2319,In_1312);
nor U2728 (N_2728,In_2324,In_445);
nand U2729 (N_2729,In_1136,In_530);
or U2730 (N_2730,In_1113,In_769);
or U2731 (N_2731,In_1926,In_1897);
nor U2732 (N_2732,In_1755,In_796);
or U2733 (N_2733,In_1121,In_599);
nor U2734 (N_2734,In_2395,In_375);
xor U2735 (N_2735,In_994,In_762);
nand U2736 (N_2736,In_2286,In_18);
and U2737 (N_2737,In_637,In_750);
or U2738 (N_2738,In_54,In_1622);
nand U2739 (N_2739,In_1669,In_647);
nor U2740 (N_2740,In_1570,In_1868);
nor U2741 (N_2741,In_2268,In_785);
nand U2742 (N_2742,In_2022,In_1080);
and U2743 (N_2743,In_1987,In_74);
and U2744 (N_2744,In_1214,In_367);
nor U2745 (N_2745,In_518,In_725);
nand U2746 (N_2746,In_1970,In_145);
xnor U2747 (N_2747,In_1540,In_1395);
nor U2748 (N_2748,In_2053,In_231);
xnor U2749 (N_2749,In_2196,In_2087);
and U2750 (N_2750,In_602,In_1526);
nor U2751 (N_2751,In_165,In_108);
nand U2752 (N_2752,In_1191,In_1791);
xor U2753 (N_2753,In_1698,In_1588);
nor U2754 (N_2754,In_1196,In_2075);
nor U2755 (N_2755,In_1478,In_1838);
and U2756 (N_2756,In_1123,In_1028);
xnor U2757 (N_2757,In_348,In_351);
or U2758 (N_2758,In_610,In_484);
and U2759 (N_2759,In_807,In_578);
or U2760 (N_2760,In_1455,In_1720);
nor U2761 (N_2761,In_400,In_863);
nand U2762 (N_2762,In_1147,In_1632);
and U2763 (N_2763,In_2296,In_959);
and U2764 (N_2764,In_2401,In_1439);
and U2765 (N_2765,In_318,In_2245);
or U2766 (N_2766,In_692,In_1064);
nand U2767 (N_2767,In_629,In_1809);
or U2768 (N_2768,In_1262,In_129);
nand U2769 (N_2769,In_863,In_1058);
and U2770 (N_2770,In_1736,In_2430);
nand U2771 (N_2771,In_2119,In_1009);
nor U2772 (N_2772,In_511,In_2226);
xnor U2773 (N_2773,In_1246,In_2135);
nor U2774 (N_2774,In_274,In_202);
and U2775 (N_2775,In_1276,In_501);
nand U2776 (N_2776,In_766,In_504);
or U2777 (N_2777,In_337,In_1547);
or U2778 (N_2778,In_1626,In_993);
xor U2779 (N_2779,In_650,In_183);
nand U2780 (N_2780,In_1294,In_1565);
nand U2781 (N_2781,In_1544,In_899);
or U2782 (N_2782,In_1963,In_945);
xnor U2783 (N_2783,In_675,In_1729);
nor U2784 (N_2784,In_1590,In_1067);
and U2785 (N_2785,In_1521,In_47);
nor U2786 (N_2786,In_2208,In_703);
nand U2787 (N_2787,In_121,In_1451);
and U2788 (N_2788,In_447,In_889);
and U2789 (N_2789,In_1140,In_392);
or U2790 (N_2790,In_1451,In_2425);
nand U2791 (N_2791,In_383,In_492);
nand U2792 (N_2792,In_1436,In_2436);
nand U2793 (N_2793,In_666,In_2131);
or U2794 (N_2794,In_1202,In_1641);
or U2795 (N_2795,In_770,In_1899);
nand U2796 (N_2796,In_627,In_334);
and U2797 (N_2797,In_2144,In_1315);
nand U2798 (N_2798,In_1939,In_967);
nor U2799 (N_2799,In_2058,In_1896);
nor U2800 (N_2800,In_436,In_1919);
and U2801 (N_2801,In_570,In_1831);
nor U2802 (N_2802,In_260,In_1179);
or U2803 (N_2803,In_2347,In_2408);
nor U2804 (N_2804,In_2016,In_1224);
or U2805 (N_2805,In_2376,In_1578);
xor U2806 (N_2806,In_1369,In_724);
or U2807 (N_2807,In_1372,In_2001);
nand U2808 (N_2808,In_1820,In_487);
or U2809 (N_2809,In_2461,In_504);
nor U2810 (N_2810,In_2446,In_2375);
nor U2811 (N_2811,In_162,In_124);
and U2812 (N_2812,In_452,In_1285);
nand U2813 (N_2813,In_299,In_1191);
or U2814 (N_2814,In_1669,In_707);
or U2815 (N_2815,In_2350,In_1321);
and U2816 (N_2816,In_607,In_1288);
nand U2817 (N_2817,In_1388,In_578);
nand U2818 (N_2818,In_279,In_686);
nand U2819 (N_2819,In_860,In_71);
or U2820 (N_2820,In_760,In_1633);
nor U2821 (N_2821,In_545,In_489);
and U2822 (N_2822,In_1353,In_2439);
nor U2823 (N_2823,In_1681,In_1197);
and U2824 (N_2824,In_1190,In_2259);
and U2825 (N_2825,In_733,In_1329);
or U2826 (N_2826,In_1531,In_1484);
or U2827 (N_2827,In_178,In_871);
or U2828 (N_2828,In_1784,In_165);
and U2829 (N_2829,In_404,In_2430);
nand U2830 (N_2830,In_996,In_129);
or U2831 (N_2831,In_249,In_1899);
nand U2832 (N_2832,In_377,In_1468);
or U2833 (N_2833,In_204,In_1218);
nor U2834 (N_2834,In_994,In_100);
nor U2835 (N_2835,In_361,In_1264);
xnor U2836 (N_2836,In_1074,In_968);
and U2837 (N_2837,In_722,In_1707);
or U2838 (N_2838,In_1883,In_359);
or U2839 (N_2839,In_2085,In_2276);
nor U2840 (N_2840,In_2007,In_1231);
and U2841 (N_2841,In_126,In_1294);
or U2842 (N_2842,In_1267,In_1077);
xor U2843 (N_2843,In_262,In_257);
or U2844 (N_2844,In_1784,In_2421);
and U2845 (N_2845,In_2196,In_821);
nand U2846 (N_2846,In_1499,In_1482);
nor U2847 (N_2847,In_2063,In_84);
nor U2848 (N_2848,In_1016,In_908);
and U2849 (N_2849,In_1097,In_1717);
nand U2850 (N_2850,In_545,In_385);
and U2851 (N_2851,In_1225,In_482);
nor U2852 (N_2852,In_29,In_982);
and U2853 (N_2853,In_1492,In_708);
nor U2854 (N_2854,In_1044,In_1014);
or U2855 (N_2855,In_324,In_892);
or U2856 (N_2856,In_2203,In_569);
and U2857 (N_2857,In_2496,In_1287);
nor U2858 (N_2858,In_618,In_1990);
nor U2859 (N_2859,In_241,In_590);
nor U2860 (N_2860,In_1192,In_2089);
and U2861 (N_2861,In_277,In_569);
xor U2862 (N_2862,In_1642,In_317);
and U2863 (N_2863,In_1666,In_2036);
nor U2864 (N_2864,In_361,In_1637);
or U2865 (N_2865,In_73,In_1825);
and U2866 (N_2866,In_735,In_2458);
nor U2867 (N_2867,In_1407,In_2193);
nand U2868 (N_2868,In_1378,In_298);
nand U2869 (N_2869,In_2018,In_230);
nand U2870 (N_2870,In_1189,In_368);
nor U2871 (N_2871,In_1048,In_1042);
or U2872 (N_2872,In_49,In_744);
and U2873 (N_2873,In_2015,In_1116);
or U2874 (N_2874,In_0,In_2269);
or U2875 (N_2875,In_807,In_1211);
or U2876 (N_2876,In_483,In_2074);
and U2877 (N_2877,In_2306,In_2426);
or U2878 (N_2878,In_1803,In_1363);
nor U2879 (N_2879,In_1922,In_2347);
and U2880 (N_2880,In_2232,In_841);
or U2881 (N_2881,In_919,In_2140);
nor U2882 (N_2882,In_1376,In_1907);
and U2883 (N_2883,In_2,In_217);
nor U2884 (N_2884,In_495,In_2311);
and U2885 (N_2885,In_1256,In_1905);
or U2886 (N_2886,In_680,In_2086);
nand U2887 (N_2887,In_221,In_1299);
or U2888 (N_2888,In_899,In_837);
nand U2889 (N_2889,In_2276,In_2119);
and U2890 (N_2890,In_1593,In_709);
nand U2891 (N_2891,In_1277,In_648);
or U2892 (N_2892,In_1891,In_380);
or U2893 (N_2893,In_1687,In_1758);
nand U2894 (N_2894,In_1115,In_1820);
or U2895 (N_2895,In_1713,In_1357);
nand U2896 (N_2896,In_2307,In_941);
nor U2897 (N_2897,In_2270,In_1123);
or U2898 (N_2898,In_945,In_444);
nand U2899 (N_2899,In_700,In_29);
and U2900 (N_2900,In_125,In_1766);
and U2901 (N_2901,In_1526,In_2237);
and U2902 (N_2902,In_80,In_2028);
nor U2903 (N_2903,In_1956,In_2267);
and U2904 (N_2904,In_2324,In_433);
nand U2905 (N_2905,In_354,In_1421);
nand U2906 (N_2906,In_188,In_156);
and U2907 (N_2907,In_2389,In_620);
nor U2908 (N_2908,In_1046,In_559);
nand U2909 (N_2909,In_1089,In_1422);
or U2910 (N_2910,In_455,In_221);
nand U2911 (N_2911,In_2297,In_217);
nand U2912 (N_2912,In_317,In_614);
or U2913 (N_2913,In_263,In_1142);
and U2914 (N_2914,In_1221,In_2408);
nand U2915 (N_2915,In_15,In_1786);
nor U2916 (N_2916,In_428,In_345);
nand U2917 (N_2917,In_2187,In_1202);
nor U2918 (N_2918,In_951,In_670);
and U2919 (N_2919,In_1931,In_928);
or U2920 (N_2920,In_2074,In_586);
or U2921 (N_2921,In_372,In_2327);
or U2922 (N_2922,In_945,In_570);
nand U2923 (N_2923,In_1936,In_750);
and U2924 (N_2924,In_742,In_1196);
nor U2925 (N_2925,In_2233,In_291);
nor U2926 (N_2926,In_1454,In_2409);
nor U2927 (N_2927,In_2146,In_1180);
nand U2928 (N_2928,In_900,In_1706);
nand U2929 (N_2929,In_1734,In_91);
nand U2930 (N_2930,In_664,In_1286);
nor U2931 (N_2931,In_2221,In_764);
or U2932 (N_2932,In_1142,In_1412);
nor U2933 (N_2933,In_431,In_112);
or U2934 (N_2934,In_887,In_434);
nor U2935 (N_2935,In_684,In_1943);
nand U2936 (N_2936,In_554,In_65);
xnor U2937 (N_2937,In_2112,In_783);
nor U2938 (N_2938,In_148,In_274);
or U2939 (N_2939,In_723,In_1593);
and U2940 (N_2940,In_131,In_1583);
xnor U2941 (N_2941,In_712,In_1197);
or U2942 (N_2942,In_2221,In_1506);
nor U2943 (N_2943,In_1339,In_1126);
or U2944 (N_2944,In_31,In_1044);
xnor U2945 (N_2945,In_1243,In_2141);
xnor U2946 (N_2946,In_986,In_40);
or U2947 (N_2947,In_926,In_2167);
nand U2948 (N_2948,In_2451,In_849);
or U2949 (N_2949,In_259,In_1898);
nand U2950 (N_2950,In_246,In_244);
and U2951 (N_2951,In_749,In_98);
and U2952 (N_2952,In_983,In_988);
nor U2953 (N_2953,In_1052,In_1330);
and U2954 (N_2954,In_1819,In_336);
nor U2955 (N_2955,In_132,In_2249);
or U2956 (N_2956,In_946,In_2351);
and U2957 (N_2957,In_287,In_2460);
nor U2958 (N_2958,In_1389,In_811);
nor U2959 (N_2959,In_1916,In_1227);
or U2960 (N_2960,In_92,In_1502);
xor U2961 (N_2961,In_1234,In_1);
and U2962 (N_2962,In_1151,In_2395);
nor U2963 (N_2963,In_1689,In_2166);
nand U2964 (N_2964,In_2130,In_1275);
or U2965 (N_2965,In_1077,In_1382);
nor U2966 (N_2966,In_199,In_1892);
nand U2967 (N_2967,In_2042,In_1513);
or U2968 (N_2968,In_132,In_1015);
nand U2969 (N_2969,In_878,In_2474);
or U2970 (N_2970,In_1082,In_82);
or U2971 (N_2971,In_1259,In_1382);
nor U2972 (N_2972,In_852,In_2226);
and U2973 (N_2973,In_1293,In_459);
and U2974 (N_2974,In_253,In_299);
or U2975 (N_2975,In_88,In_2470);
nor U2976 (N_2976,In_1463,In_915);
nand U2977 (N_2977,In_617,In_61);
or U2978 (N_2978,In_10,In_1279);
or U2979 (N_2979,In_2031,In_29);
or U2980 (N_2980,In_198,In_654);
or U2981 (N_2981,In_698,In_1186);
nand U2982 (N_2982,In_1934,In_1159);
or U2983 (N_2983,In_2169,In_1);
or U2984 (N_2984,In_98,In_2489);
and U2985 (N_2985,In_570,In_511);
xor U2986 (N_2986,In_1287,In_1386);
or U2987 (N_2987,In_441,In_549);
nor U2988 (N_2988,In_304,In_2451);
nor U2989 (N_2989,In_1830,In_725);
nand U2990 (N_2990,In_1759,In_531);
or U2991 (N_2991,In_1428,In_1462);
nor U2992 (N_2992,In_126,In_1502);
nand U2993 (N_2993,In_941,In_2173);
nor U2994 (N_2994,In_1591,In_1224);
nand U2995 (N_2995,In_2490,In_1972);
nor U2996 (N_2996,In_2323,In_506);
and U2997 (N_2997,In_2294,In_1677);
nand U2998 (N_2998,In_1899,In_812);
nand U2999 (N_2999,In_2326,In_540);
or U3000 (N_3000,In_1722,In_1130);
xnor U3001 (N_3001,In_865,In_1180);
nand U3002 (N_3002,In_2267,In_70);
and U3003 (N_3003,In_357,In_1830);
and U3004 (N_3004,In_1996,In_1363);
or U3005 (N_3005,In_1591,In_1344);
or U3006 (N_3006,In_1783,In_1875);
or U3007 (N_3007,In_1762,In_2037);
and U3008 (N_3008,In_870,In_897);
and U3009 (N_3009,In_1412,In_82);
and U3010 (N_3010,In_2096,In_473);
nand U3011 (N_3011,In_753,In_2448);
nor U3012 (N_3012,In_1700,In_307);
xnor U3013 (N_3013,In_2258,In_2298);
nand U3014 (N_3014,In_709,In_1787);
or U3015 (N_3015,In_1340,In_1159);
or U3016 (N_3016,In_365,In_1413);
or U3017 (N_3017,In_2433,In_1011);
or U3018 (N_3018,In_2143,In_399);
or U3019 (N_3019,In_983,In_196);
nand U3020 (N_3020,In_897,In_1608);
nand U3021 (N_3021,In_2186,In_1519);
nor U3022 (N_3022,In_5,In_2305);
nand U3023 (N_3023,In_1862,In_2325);
and U3024 (N_3024,In_344,In_162);
and U3025 (N_3025,In_1457,In_212);
nand U3026 (N_3026,In_244,In_1265);
or U3027 (N_3027,In_870,In_2148);
xor U3028 (N_3028,In_1280,In_2305);
and U3029 (N_3029,In_983,In_948);
or U3030 (N_3030,In_458,In_1318);
and U3031 (N_3031,In_411,In_302);
nand U3032 (N_3032,In_1838,In_1620);
or U3033 (N_3033,In_84,In_524);
and U3034 (N_3034,In_710,In_1613);
xnor U3035 (N_3035,In_1563,In_757);
nand U3036 (N_3036,In_371,In_396);
or U3037 (N_3037,In_1280,In_12);
and U3038 (N_3038,In_1439,In_2389);
and U3039 (N_3039,In_2270,In_2223);
or U3040 (N_3040,In_392,In_2275);
xor U3041 (N_3041,In_1566,In_25);
or U3042 (N_3042,In_1589,In_86);
xor U3043 (N_3043,In_1701,In_2429);
nand U3044 (N_3044,In_770,In_1598);
and U3045 (N_3045,In_921,In_1121);
nor U3046 (N_3046,In_1368,In_1537);
nor U3047 (N_3047,In_908,In_267);
or U3048 (N_3048,In_1717,In_292);
nor U3049 (N_3049,In_807,In_1952);
xnor U3050 (N_3050,In_956,In_97);
and U3051 (N_3051,In_1459,In_2480);
nor U3052 (N_3052,In_2396,In_1055);
and U3053 (N_3053,In_733,In_2271);
nor U3054 (N_3054,In_1639,In_2472);
nand U3055 (N_3055,In_519,In_1550);
and U3056 (N_3056,In_91,In_1504);
and U3057 (N_3057,In_347,In_1524);
and U3058 (N_3058,In_248,In_1585);
or U3059 (N_3059,In_1783,In_2401);
xnor U3060 (N_3060,In_115,In_1437);
nor U3061 (N_3061,In_727,In_1296);
and U3062 (N_3062,In_337,In_927);
or U3063 (N_3063,In_627,In_1846);
nor U3064 (N_3064,In_2457,In_1805);
nor U3065 (N_3065,In_1896,In_453);
and U3066 (N_3066,In_2065,In_42);
or U3067 (N_3067,In_2026,In_128);
nand U3068 (N_3068,In_1393,In_644);
and U3069 (N_3069,In_104,In_509);
or U3070 (N_3070,In_721,In_1511);
and U3071 (N_3071,In_733,In_1780);
or U3072 (N_3072,In_1067,In_2461);
and U3073 (N_3073,In_395,In_1316);
and U3074 (N_3074,In_1643,In_698);
nand U3075 (N_3075,In_1254,In_1173);
or U3076 (N_3076,In_2166,In_1244);
or U3077 (N_3077,In_1878,In_2384);
nand U3078 (N_3078,In_1413,In_863);
or U3079 (N_3079,In_22,In_763);
and U3080 (N_3080,In_904,In_778);
nor U3081 (N_3081,In_223,In_2212);
or U3082 (N_3082,In_1248,In_185);
or U3083 (N_3083,In_2220,In_794);
nand U3084 (N_3084,In_1564,In_2288);
nand U3085 (N_3085,In_2054,In_486);
nand U3086 (N_3086,In_2337,In_1292);
nor U3087 (N_3087,In_443,In_2479);
and U3088 (N_3088,In_1937,In_1438);
nor U3089 (N_3089,In_1214,In_356);
or U3090 (N_3090,In_1128,In_291);
nor U3091 (N_3091,In_664,In_683);
nor U3092 (N_3092,In_2031,In_2316);
and U3093 (N_3093,In_1907,In_1378);
nor U3094 (N_3094,In_216,In_1097);
and U3095 (N_3095,In_1845,In_289);
nand U3096 (N_3096,In_600,In_57);
and U3097 (N_3097,In_1469,In_1181);
nor U3098 (N_3098,In_1314,In_844);
nand U3099 (N_3099,In_1906,In_1594);
nand U3100 (N_3100,In_844,In_2495);
and U3101 (N_3101,In_741,In_1930);
nor U3102 (N_3102,In_386,In_99);
and U3103 (N_3103,In_2075,In_781);
nor U3104 (N_3104,In_1753,In_1719);
or U3105 (N_3105,In_2165,In_1686);
nor U3106 (N_3106,In_2002,In_304);
or U3107 (N_3107,In_399,In_1802);
or U3108 (N_3108,In_2196,In_1638);
or U3109 (N_3109,In_1075,In_394);
xnor U3110 (N_3110,In_340,In_516);
nand U3111 (N_3111,In_1940,In_1263);
nor U3112 (N_3112,In_1865,In_1573);
nor U3113 (N_3113,In_1957,In_13);
nor U3114 (N_3114,In_1623,In_1042);
nand U3115 (N_3115,In_713,In_1975);
and U3116 (N_3116,In_2158,In_962);
nand U3117 (N_3117,In_1541,In_1258);
or U3118 (N_3118,In_759,In_1741);
nor U3119 (N_3119,In_1104,In_1371);
nand U3120 (N_3120,In_870,In_1720);
or U3121 (N_3121,In_108,In_1234);
nand U3122 (N_3122,In_842,In_852);
or U3123 (N_3123,In_1414,In_211);
nand U3124 (N_3124,In_2284,In_2235);
xnor U3125 (N_3125,N_872,N_1484);
xor U3126 (N_3126,N_2220,N_1785);
and U3127 (N_3127,N_2057,N_797);
and U3128 (N_3128,N_1026,N_2957);
xor U3129 (N_3129,N_2367,N_1167);
nand U3130 (N_3130,N_899,N_2167);
and U3131 (N_3131,N_2649,N_2169);
or U3132 (N_3132,N_1033,N_2961);
or U3133 (N_3133,N_2773,N_2480);
nand U3134 (N_3134,N_485,N_2245);
and U3135 (N_3135,N_2016,N_599);
nand U3136 (N_3136,N_1809,N_247);
and U3137 (N_3137,N_2607,N_1731);
or U3138 (N_3138,N_1481,N_817);
or U3139 (N_3139,N_1926,N_821);
nor U3140 (N_3140,N_1909,N_1937);
and U3141 (N_3141,N_2261,N_2684);
nor U3142 (N_3142,N_1504,N_2902);
and U3143 (N_3143,N_2890,N_1202);
and U3144 (N_3144,N_1983,N_1276);
nor U3145 (N_3145,N_2692,N_97);
nor U3146 (N_3146,N_904,N_1257);
nor U3147 (N_3147,N_1805,N_74);
and U3148 (N_3148,N_1599,N_761);
and U3149 (N_3149,N_2519,N_1806);
nand U3150 (N_3150,N_1549,N_2206);
nor U3151 (N_3151,N_2217,N_547);
or U3152 (N_3152,N_951,N_2403);
nand U3153 (N_3153,N_2048,N_1993);
and U3154 (N_3154,N_2710,N_2462);
and U3155 (N_3155,N_331,N_2296);
nor U3156 (N_3156,N_1839,N_1954);
or U3157 (N_3157,N_1596,N_2826);
nor U3158 (N_3158,N_1380,N_2198);
or U3159 (N_3159,N_2465,N_2588);
nor U3160 (N_3160,N_1323,N_668);
nand U3161 (N_3161,N_1096,N_2639);
or U3162 (N_3162,N_812,N_1821);
xor U3163 (N_3163,N_524,N_2471);
nand U3164 (N_3164,N_2407,N_528);
nor U3165 (N_3165,N_553,N_1247);
nand U3166 (N_3166,N_1992,N_2022);
and U3167 (N_3167,N_2627,N_2557);
nor U3168 (N_3168,N_799,N_1774);
and U3169 (N_3169,N_2676,N_2771);
xor U3170 (N_3170,N_1958,N_2674);
nand U3171 (N_3171,N_2443,N_173);
or U3172 (N_3172,N_1246,N_1070);
or U3173 (N_3173,N_447,N_911);
and U3174 (N_3174,N_52,N_2078);
and U3175 (N_3175,N_138,N_1157);
or U3176 (N_3176,N_2663,N_2528);
nor U3177 (N_3177,N_357,N_339);
nand U3178 (N_3178,N_2130,N_360);
nand U3179 (N_3179,N_1294,N_98);
and U3180 (N_3180,N_1870,N_16);
or U3181 (N_3181,N_2833,N_3089);
nor U3182 (N_3182,N_1517,N_2321);
and U3183 (N_3183,N_809,N_2909);
nor U3184 (N_3184,N_733,N_1892);
nor U3185 (N_3185,N_3092,N_111);
or U3186 (N_3186,N_1694,N_1828);
and U3187 (N_3187,N_328,N_216);
nand U3188 (N_3188,N_1123,N_1317);
nand U3189 (N_3189,N_2014,N_1637);
or U3190 (N_3190,N_236,N_1492);
nor U3191 (N_3191,N_3038,N_2160);
and U3192 (N_3192,N_944,N_2106);
nand U3193 (N_3193,N_1829,N_155);
xnor U3194 (N_3194,N_2521,N_2186);
and U3195 (N_3195,N_660,N_801);
nor U3196 (N_3196,N_1568,N_1501);
xor U3197 (N_3197,N_418,N_1746);
nor U3198 (N_3198,N_2230,N_859);
xnor U3199 (N_3199,N_248,N_197);
nor U3200 (N_3200,N_2887,N_463);
xor U3201 (N_3201,N_2794,N_2857);
or U3202 (N_3202,N_609,N_1188);
nor U3203 (N_3203,N_12,N_2327);
or U3204 (N_3204,N_2747,N_1547);
nor U3205 (N_3205,N_1154,N_1527);
or U3206 (N_3206,N_2455,N_321);
and U3207 (N_3207,N_1652,N_424);
or U3208 (N_3208,N_1303,N_263);
or U3209 (N_3209,N_2615,N_223);
nor U3210 (N_3210,N_2181,N_2533);
nor U3211 (N_3211,N_564,N_2702);
nor U3212 (N_3212,N_1150,N_2091);
nor U3213 (N_3213,N_1091,N_1251);
nand U3214 (N_3214,N_2193,N_2038);
and U3215 (N_3215,N_1689,N_87);
and U3216 (N_3216,N_2872,N_276);
nand U3217 (N_3217,N_1665,N_1301);
and U3218 (N_3218,N_390,N_1949);
xor U3219 (N_3219,N_370,N_243);
nor U3220 (N_3220,N_2073,N_1716);
and U3221 (N_3221,N_1739,N_1505);
nor U3222 (N_3222,N_180,N_2527);
and U3223 (N_3223,N_487,N_2147);
and U3224 (N_3224,N_2373,N_664);
nor U3225 (N_3225,N_2779,N_3035);
and U3226 (N_3226,N_2659,N_1600);
nand U3227 (N_3227,N_129,N_536);
and U3228 (N_3228,N_1006,N_1106);
nor U3229 (N_3229,N_2232,N_1864);
or U3230 (N_3230,N_1094,N_771);
or U3231 (N_3231,N_1268,N_324);
and U3232 (N_3232,N_2817,N_1795);
and U3233 (N_3233,N_2041,N_2545);
nor U3234 (N_3234,N_1927,N_1262);
or U3235 (N_3235,N_569,N_565);
nor U3236 (N_3236,N_946,N_3009);
and U3237 (N_3237,N_127,N_1868);
nor U3238 (N_3238,N_685,N_2955);
or U3239 (N_3239,N_240,N_158);
or U3240 (N_3240,N_2845,N_1728);
xor U3241 (N_3241,N_375,N_2379);
nor U3242 (N_3242,N_1978,N_1046);
or U3243 (N_3243,N_2675,N_3050);
nor U3244 (N_3244,N_2020,N_2582);
nor U3245 (N_3245,N_2156,N_193);
nor U3246 (N_3246,N_915,N_1312);
or U3247 (N_3247,N_304,N_1942);
or U3248 (N_3248,N_786,N_394);
or U3249 (N_3249,N_3001,N_742);
or U3250 (N_3250,N_64,N_1922);
nor U3251 (N_3251,N_2489,N_199);
or U3252 (N_3252,N_787,N_459);
or U3253 (N_3253,N_2138,N_2405);
and U3254 (N_3254,N_1789,N_120);
and U3255 (N_3255,N_1292,N_577);
or U3256 (N_3256,N_2170,N_1277);
nand U3257 (N_3257,N_1855,N_1567);
or U3258 (N_3258,N_1972,N_943);
and U3259 (N_3259,N_2903,N_1351);
nand U3260 (N_3260,N_2974,N_54);
and U3261 (N_3261,N_839,N_23);
or U3262 (N_3262,N_1379,N_2302);
nor U3263 (N_3263,N_1895,N_3046);
or U3264 (N_3264,N_2458,N_3004);
nand U3265 (N_3265,N_453,N_3000);
nor U3266 (N_3266,N_2700,N_2286);
and U3267 (N_3267,N_169,N_2430);
nor U3268 (N_3268,N_456,N_1743);
nor U3269 (N_3269,N_3062,N_1069);
and U3270 (N_3270,N_665,N_470);
or U3271 (N_3271,N_250,N_813);
nor U3272 (N_3272,N_2592,N_208);
nor U3273 (N_3273,N_527,N_1664);
xnor U3274 (N_3274,N_932,N_2237);
and U3275 (N_3275,N_2882,N_306);
nor U3276 (N_3276,N_1705,N_1462);
or U3277 (N_3277,N_1437,N_1245);
or U3278 (N_3278,N_2113,N_1095);
nor U3279 (N_3279,N_2337,N_1348);
and U3280 (N_3280,N_1945,N_1563);
nor U3281 (N_3281,N_1745,N_992);
or U3282 (N_3282,N_873,N_2531);
or U3283 (N_3283,N_995,N_1410);
nor U3284 (N_3284,N_2419,N_1963);
nand U3285 (N_3285,N_3066,N_2459);
nor U3286 (N_3286,N_1024,N_343);
nand U3287 (N_3287,N_631,N_1853);
nor U3288 (N_3288,N_1889,N_403);
nand U3289 (N_3289,N_1990,N_39);
nand U3290 (N_3290,N_1555,N_604);
or U3291 (N_3291,N_763,N_847);
or U3292 (N_3292,N_607,N_1820);
xnor U3293 (N_3293,N_2028,N_1620);
nand U3294 (N_3294,N_2435,N_2049);
nor U3295 (N_3295,N_2103,N_218);
and U3296 (N_3296,N_989,N_2287);
and U3297 (N_3297,N_2668,N_918);
nand U3298 (N_3298,N_1622,N_1908);
nor U3299 (N_3299,N_2197,N_618);
and U3300 (N_3300,N_66,N_719);
and U3301 (N_3301,N_1695,N_1152);
nor U3302 (N_3302,N_2412,N_363);
or U3303 (N_3303,N_1766,N_427);
and U3304 (N_3304,N_175,N_766);
xnor U3305 (N_3305,N_2324,N_1229);
nor U3306 (N_3306,N_1956,N_691);
and U3307 (N_3307,N_796,N_2381);
and U3308 (N_3308,N_1242,N_349);
nand U3309 (N_3309,N_1976,N_1191);
or U3310 (N_3310,N_1604,N_2716);
nor U3311 (N_3311,N_3095,N_49);
nor U3312 (N_3312,N_1102,N_2852);
nand U3313 (N_3313,N_886,N_746);
nand U3314 (N_3314,N_2602,N_2297);
or U3315 (N_3315,N_2553,N_793);
nand U3316 (N_3316,N_1987,N_682);
nor U3317 (N_3317,N_2919,N_1944);
or U3318 (N_3318,N_2670,N_389);
xnor U3319 (N_3319,N_1635,N_106);
or U3320 (N_3320,N_597,N_29);
nand U3321 (N_3321,N_1019,N_2240);
nand U3322 (N_3322,N_119,N_3090);
nand U3323 (N_3323,N_85,N_2671);
xnor U3324 (N_3324,N_1285,N_1421);
or U3325 (N_3325,N_1856,N_2939);
nand U3326 (N_3326,N_117,N_1640);
nand U3327 (N_3327,N_294,N_2927);
and U3328 (N_3328,N_1712,N_2848);
xor U3329 (N_3329,N_2040,N_2142);
nand U3330 (N_3330,N_1479,N_1030);
and U3331 (N_3331,N_2564,N_2139);
and U3332 (N_3332,N_426,N_2714);
nand U3333 (N_3333,N_983,N_2841);
nor U3334 (N_3334,N_1482,N_1588);
nor U3335 (N_3335,N_1316,N_2488);
and U3336 (N_3336,N_268,N_709);
or U3337 (N_3337,N_406,N_2479);
nor U3338 (N_3338,N_1736,N_1684);
and U3339 (N_3339,N_2356,N_2154);
nand U3340 (N_3340,N_883,N_1538);
or U3341 (N_3341,N_2086,N_2425);
nor U3342 (N_3342,N_1930,N_2177);
or U3343 (N_3343,N_641,N_1283);
nor U3344 (N_3344,N_945,N_889);
xor U3345 (N_3345,N_1562,N_2941);
nand U3346 (N_3346,N_2234,N_77);
or U3347 (N_3347,N_2829,N_458);
nand U3348 (N_3348,N_2474,N_1758);
nor U3349 (N_3349,N_341,N_1180);
and U3350 (N_3350,N_2188,N_388);
and U3351 (N_3351,N_2983,N_2605);
or U3352 (N_3352,N_474,N_1417);
or U3353 (N_3353,N_404,N_2594);
or U3354 (N_3354,N_2910,N_2062);
or U3355 (N_3355,N_2775,N_19);
or U3356 (N_3356,N_1430,N_2331);
nand U3357 (N_3357,N_1841,N_1066);
nor U3358 (N_3358,N_712,N_2242);
nand U3359 (N_3359,N_1867,N_1280);
or U3360 (N_3360,N_1392,N_3024);
or U3361 (N_3361,N_2359,N_2896);
or U3362 (N_3362,N_2473,N_2394);
nor U3363 (N_3363,N_566,N_2768);
or U3364 (N_3364,N_1548,N_2399);
and U3365 (N_3365,N_1063,N_2212);
nor U3366 (N_3366,N_2210,N_1438);
xnor U3367 (N_3367,N_1452,N_1584);
and U3368 (N_3368,N_2850,N_2013);
nand U3369 (N_3369,N_1439,N_104);
nor U3370 (N_3370,N_1387,N_184);
and U3371 (N_3371,N_806,N_420);
nand U3372 (N_3372,N_36,N_78);
and U3373 (N_3373,N_1896,N_598);
or U3374 (N_3374,N_1151,N_2618);
xnor U3375 (N_3375,N_2752,N_822);
and U3376 (N_3376,N_1556,N_2087);
or U3377 (N_3377,N_578,N_1675);
and U3378 (N_3378,N_3117,N_1884);
or U3379 (N_3379,N_1784,N_189);
xor U3380 (N_3380,N_2691,N_810);
nand U3381 (N_3381,N_2025,N_1209);
or U3382 (N_3382,N_225,N_1815);
xnor U3383 (N_3383,N_2076,N_1244);
nand U3384 (N_3384,N_1237,N_625);
nor U3385 (N_3385,N_2883,N_953);
or U3386 (N_3386,N_2348,N_200);
nor U3387 (N_3387,N_2556,N_1068);
or U3388 (N_3388,N_2309,N_2270);
nor U3389 (N_3389,N_1376,N_2165);
nor U3390 (N_3390,N_1529,N_1087);
or U3391 (N_3391,N_1441,N_1748);
nand U3392 (N_3392,N_2226,N_214);
nor U3393 (N_3393,N_2836,N_2370);
nor U3394 (N_3394,N_2898,N_1476);
and U3395 (N_3395,N_1878,N_764);
xnor U3396 (N_3396,N_1149,N_2783);
nor U3397 (N_3397,N_563,N_2427);
nand U3398 (N_3398,N_818,N_2942);
nand U3399 (N_3399,N_3064,N_2968);
or U3400 (N_3400,N_931,N_1733);
nor U3401 (N_3401,N_1638,N_715);
nor U3402 (N_3402,N_2662,N_1770);
nand U3403 (N_3403,N_884,N_716);
or U3404 (N_3404,N_209,N_227);
nand U3405 (N_3405,N_1647,N_1022);
xnor U3406 (N_3406,N_108,N_414);
or U3407 (N_3407,N_2544,N_1579);
or U3408 (N_3408,N_549,N_1175);
and U3409 (N_3409,N_1816,N_2257);
xor U3410 (N_3410,N_533,N_1118);
or U3411 (N_3411,N_3078,N_2301);
or U3412 (N_3412,N_653,N_2892);
nor U3413 (N_3413,N_2808,N_1539);
nand U3414 (N_3414,N_1718,N_1212);
and U3415 (N_3415,N_3053,N_457);
or U3416 (N_3416,N_1726,N_280);
or U3417 (N_3417,N_2908,N_3091);
nor U3418 (N_3418,N_115,N_2965);
or U3419 (N_3419,N_415,N_1402);
nand U3420 (N_3420,N_3122,N_881);
and U3421 (N_3421,N_2837,N_136);
nand U3422 (N_3422,N_1724,N_267);
and U3423 (N_3423,N_188,N_68);
and U3424 (N_3424,N_878,N_95);
and U3425 (N_3425,N_2858,N_823);
xor U3426 (N_3426,N_190,N_1776);
nor U3427 (N_3427,N_1080,N_2574);
and U3428 (N_3428,N_1398,N_534);
nand U3429 (N_3429,N_1271,N_2661);
nand U3430 (N_3430,N_1365,N_2935);
nand U3431 (N_3431,N_2061,N_2828);
nor U3432 (N_3432,N_2352,N_2901);
or U3433 (N_3433,N_425,N_1759);
xnor U3434 (N_3434,N_2772,N_3094);
nand U3435 (N_3435,N_2863,N_2164);
or U3436 (N_3436,N_868,N_1749);
xor U3437 (N_3437,N_649,N_555);
nand U3438 (N_3438,N_1198,N_141);
nor U3439 (N_3439,N_438,N_2767);
or U3440 (N_3440,N_2037,N_2314);
nand U3441 (N_3441,N_409,N_1170);
and U3442 (N_3442,N_638,N_269);
and U3443 (N_3443,N_701,N_45);
or U3444 (N_3444,N_2499,N_3068);
nand U3445 (N_3445,N_2264,N_2753);
nor U3446 (N_3446,N_819,N_2224);
nor U3447 (N_3447,N_2102,N_2922);
nand U3448 (N_3448,N_844,N_1626);
nand U3449 (N_3449,N_1557,N_2416);
nand U3450 (N_3450,N_956,N_571);
or U3451 (N_3451,N_2687,N_1617);
or U3452 (N_3452,N_504,N_1953);
or U3453 (N_3453,N_131,N_135);
nand U3454 (N_3454,N_61,N_271);
or U3455 (N_3455,N_3036,N_1830);
nor U3456 (N_3456,N_2135,N_288);
xor U3457 (N_3457,N_2024,N_1060);
nand U3458 (N_3458,N_1844,N_5);
and U3459 (N_3459,N_273,N_67);
nand U3460 (N_3460,N_2704,N_356);
and U3461 (N_3461,N_2283,N_2899);
and U3462 (N_3462,N_1148,N_14);
nor U3463 (N_3463,N_882,N_2105);
nor U3464 (N_3464,N_639,N_1863);
nand U3465 (N_3465,N_2548,N_2140);
nand U3466 (N_3466,N_205,N_655);
nand U3467 (N_3467,N_1140,N_336);
and U3468 (N_3468,N_378,N_411);
or U3469 (N_3469,N_1645,N_1898);
or U3470 (N_3470,N_382,N_2623);
or U3471 (N_3471,N_949,N_2354);
and U3472 (N_3472,N_2127,N_678);
nor U3473 (N_3473,N_1491,N_1221);
or U3474 (N_3474,N_1660,N_230);
nand U3475 (N_3475,N_1193,N_303);
nand U3476 (N_3476,N_1797,N_957);
nand U3477 (N_3477,N_2295,N_2547);
and U3478 (N_3478,N_2422,N_50);
or U3479 (N_3479,N_1509,N_1925);
nor U3480 (N_3480,N_798,N_515);
nor U3481 (N_3481,N_1593,N_1359);
nand U3482 (N_3482,N_1015,N_1888);
nor U3483 (N_3483,N_2822,N_3077);
nor U3484 (N_3484,N_22,N_1667);
nor U3485 (N_3485,N_2967,N_292);
nand U3486 (N_3486,N_258,N_2884);
or U3487 (N_3487,N_1999,N_2006);
and U3488 (N_3488,N_465,N_1056);
nor U3489 (N_3489,N_2997,N_1488);
or U3490 (N_3490,N_803,N_2298);
nor U3491 (N_3491,N_3069,N_1083);
nor U3492 (N_3492,N_2940,N_708);
or U3493 (N_3493,N_2930,N_2386);
nor U3494 (N_3494,N_21,N_550);
or U3495 (N_3495,N_322,N_2218);
or U3496 (N_3496,N_102,N_2677);
and U3497 (N_3497,N_2820,N_916);
nand U3498 (N_3498,N_2308,N_2995);
nand U3499 (N_3499,N_183,N_907);
or U3500 (N_3500,N_3016,N_126);
xnor U3501 (N_3501,N_320,N_2570);
or U3502 (N_3502,N_1835,N_3055);
nand U3503 (N_3503,N_2727,N_2401);
or U3504 (N_3504,N_608,N_170);
nand U3505 (N_3505,N_1606,N_1383);
nand U3506 (N_3506,N_830,N_1269);
or U3507 (N_3507,N_2256,N_1425);
nor U3508 (N_3508,N_1516,N_2015);
or U3509 (N_3509,N_2325,N_2318);
nor U3510 (N_3510,N_1525,N_1852);
nand U3511 (N_3511,N_1764,N_1882);
and U3512 (N_3512,N_610,N_2228);
nor U3513 (N_3513,N_690,N_1176);
and U3514 (N_3514,N_1319,N_1796);
nor U3515 (N_3515,N_662,N_1814);
or U3516 (N_3516,N_2996,N_2083);
or U3517 (N_3517,N_2757,N_699);
nand U3518 (N_3518,N_1499,N_3124);
or U3519 (N_3519,N_1636,N_1754);
and U3520 (N_3520,N_1536,N_1623);
nor U3521 (N_3521,N_2561,N_1763);
or U3522 (N_3522,N_1840,N_1744);
nor U3523 (N_3523,N_2111,N_1381);
nand U3524 (N_3524,N_3003,N_1740);
or U3525 (N_3525,N_773,N_2760);
and U3526 (N_3526,N_172,N_1296);
or U3527 (N_3527,N_758,N_2338);
nand U3528 (N_3528,N_192,N_2);
xnor U3529 (N_3529,N_905,N_3102);
nor U3530 (N_3530,N_1912,N_2635);
and U3531 (N_3531,N_311,N_431);
or U3532 (N_3532,N_2213,N_71);
and U3533 (N_3533,N_2158,N_1813);
or U3534 (N_3534,N_970,N_1669);
nand U3535 (N_3535,N_140,N_1966);
and U3536 (N_3536,N_1164,N_2924);
nand U3537 (N_3537,N_1769,N_467);
and U3538 (N_3538,N_2926,N_1649);
and U3539 (N_3539,N_930,N_2109);
or U3540 (N_3540,N_552,N_1985);
xor U3541 (N_3541,N_1132,N_2736);
or U3542 (N_3542,N_1451,N_2002);
and U3543 (N_3543,N_2614,N_1683);
nor U3544 (N_3544,N_31,N_1655);
nand U3545 (N_3545,N_3019,N_2789);
nand U3546 (N_3546,N_42,N_2653);
xnor U3547 (N_3547,N_1061,N_413);
nand U3548 (N_3548,N_482,N_2770);
or U3549 (N_3549,N_1799,N_2993);
xor U3550 (N_3550,N_3111,N_2391);
nor U3551 (N_3551,N_2569,N_1017);
or U3552 (N_3552,N_961,N_1103);
and U3553 (N_3553,N_1613,N_2268);
and U3554 (N_3554,N_857,N_2179);
or U3555 (N_3555,N_1394,N_232);
nand U3556 (N_3556,N_1270,N_2529);
nand U3557 (N_3557,N_740,N_264);
nor U3558 (N_3558,N_2263,N_755);
nand U3559 (N_3559,N_157,N_1363);
nor U3560 (N_3560,N_2056,N_1977);
and U3561 (N_3561,N_2696,N_1115);
and U3562 (N_3562,N_3098,N_2320);
xor U3563 (N_3563,N_2629,N_2498);
nor U3564 (N_3564,N_2917,N_2577);
xnor U3565 (N_3565,N_925,N_2648);
and U3566 (N_3566,N_1998,N_2063);
nand U3567 (N_3567,N_481,N_2291);
and U3568 (N_3568,N_2492,N_3052);
or U3569 (N_3569,N_1223,N_2428);
nor U3570 (N_3570,N_2617,N_697);
nand U3571 (N_3571,N_450,N_3123);
nand U3572 (N_3572,N_1207,N_1752);
nand U3573 (N_3573,N_567,N_151);
or U3574 (N_3574,N_1634,N_2542);
and U3575 (N_3575,N_2460,N_1357);
xor U3576 (N_3576,N_2766,N_1012);
and U3577 (N_3577,N_444,N_750);
xnor U3578 (N_3578,N_2970,N_1495);
nor U3579 (N_3579,N_2843,N_1933);
and U3580 (N_3580,N_2233,N_2801);
nor U3581 (N_3581,N_2952,N_659);
nand U3582 (N_3582,N_2503,N_2375);
nand U3583 (N_3583,N_15,N_681);
or U3584 (N_3584,N_1881,N_1952);
nand U3585 (N_3585,N_2010,N_2200);
and U3586 (N_3586,N_2364,N_1447);
xor U3587 (N_3587,N_2027,N_2721);
nor U3588 (N_3588,N_392,N_2440);
and U3589 (N_3589,N_2634,N_1506);
or U3590 (N_3590,N_1920,N_1058);
and U3591 (N_3591,N_1619,N_1013);
and U3592 (N_3592,N_2537,N_1122);
and U3593 (N_3593,N_2163,N_460);
nand U3594 (N_3594,N_1234,N_2420);
nor U3595 (N_3595,N_2021,N_2340);
or U3596 (N_3596,N_2797,N_2005);
nor U3597 (N_3597,N_285,N_1399);
or U3598 (N_3598,N_1045,N_926);
or U3599 (N_3599,N_496,N_785);
or U3600 (N_3600,N_1824,N_2842);
nor U3601 (N_3601,N_1996,N_3041);
or U3602 (N_3602,N_579,N_82);
nor U3603 (N_3603,N_1875,N_2094);
nor U3604 (N_3604,N_1897,N_1334);
and U3605 (N_3605,N_408,N_2238);
nor U3606 (N_3606,N_1048,N_1420);
and U3607 (N_3607,N_616,N_1227);
and U3608 (N_3608,N_1943,N_1656);
xor U3609 (N_3609,N_291,N_2377);
nand U3610 (N_3610,N_233,N_760);
and U3611 (N_3611,N_2121,N_829);
and U3612 (N_3612,N_391,N_2129);
nand U3613 (N_3613,N_2708,N_2991);
and U3614 (N_3614,N_72,N_2853);
nand U3615 (N_3615,N_947,N_1885);
and U3616 (N_3616,N_977,N_1971);
nand U3617 (N_3617,N_212,N_972);
or U3618 (N_3618,N_436,N_2125);
and U3619 (N_3619,N_257,N_1435);
nand U3620 (N_3620,N_1366,N_2496);
or U3621 (N_3621,N_942,N_1515);
or U3622 (N_3622,N_1325,N_1948);
nand U3623 (N_3623,N_1757,N_261);
nor U3624 (N_3624,N_2493,N_2579);
nor U3625 (N_3625,N_2312,N_789);
nor U3626 (N_3626,N_1166,N_228);
nor U3627 (N_3627,N_1373,N_1085);
nand U3628 (N_3628,N_540,N_150);
nand U3629 (N_3629,N_1589,N_1710);
nand U3630 (N_3630,N_1051,N_132);
and U3631 (N_3631,N_2000,N_3088);
or U3632 (N_3632,N_2840,N_3065);
or U3633 (N_3633,N_1217,N_1475);
nor U3634 (N_3634,N_832,N_84);
nand U3635 (N_3635,N_6,N_1213);
and U3636 (N_3636,N_2609,N_1137);
nand U3637 (N_3637,N_3120,N_603);
and U3638 (N_3638,N_134,N_2580);
and U3639 (N_3639,N_484,N_1463);
nand U3640 (N_3640,N_2089,N_2393);
and U3641 (N_3641,N_2748,N_2478);
nor U3642 (N_3642,N_130,N_2053);
and U3643 (N_3643,N_123,N_635);
nor U3644 (N_3644,N_1682,N_1706);
nand U3645 (N_3645,N_2520,N_3096);
or U3646 (N_3646,N_310,N_2642);
nand U3647 (N_3647,N_2423,N_3081);
nand U3648 (N_3648,N_2806,N_1003);
nor U3649 (N_3649,N_1225,N_2728);
nand U3650 (N_3650,N_367,N_999);
nor U3651 (N_3651,N_2215,N_833);
nand U3652 (N_3652,N_377,N_1862);
nand U3653 (N_3653,N_3043,N_2055);
nor U3654 (N_3654,N_1541,N_2637);
or U3655 (N_3655,N_477,N_2491);
nand U3656 (N_3656,N_2711,N_1018);
nand U3657 (N_3657,N_2984,N_711);
xnor U3658 (N_3658,N_3101,N_96);
nor U3659 (N_3659,N_231,N_2856);
xnor U3660 (N_3660,N_221,N_1629);
and U3661 (N_3661,N_556,N_1838);
and U3662 (N_3662,N_842,N_206);
or U3663 (N_3663,N_3045,N_2762);
nand U3664 (N_3664,N_585,N_3017);
nor U3665 (N_3665,N_741,N_2402);
or U3666 (N_3666,N_2538,N_1891);
and U3667 (N_3667,N_2698,N_2690);
nor U3668 (N_3668,N_1480,N_2467);
or U3669 (N_3669,N_198,N_3047);
and U3670 (N_3670,N_689,N_2011);
nand U3671 (N_3671,N_1576,N_1627);
nor U3672 (N_3672,N_1672,N_1356);
nor U3673 (N_3673,N_1940,N_1616);
or U3674 (N_3674,N_396,N_202);
or U3675 (N_3675,N_2067,N_1500);
and U3676 (N_3676,N_47,N_3109);
nand U3677 (N_3677,N_702,N_2575);
nand U3678 (N_3678,N_397,N_2072);
and U3679 (N_3679,N_449,N_677);
nor U3680 (N_3680,N_2506,N_455);
or U3681 (N_3681,N_1704,N_2382);
or U3682 (N_3682,N_2384,N_1585);
nand U3683 (N_3683,N_2593,N_2632);
nor U3684 (N_3684,N_51,N_734);
and U3685 (N_3685,N_3026,N_69);
or U3686 (N_3686,N_2631,N_634);
nor U3687 (N_3687,N_2715,N_272);
nand U3688 (N_3688,N_1162,N_1642);
nor U3689 (N_3689,N_299,N_2070);
nor U3690 (N_3690,N_871,N_2765);
or U3691 (N_3691,N_952,N_530);
xnor U3692 (N_3692,N_76,N_2483);
nand U3693 (N_3693,N_28,N_2791);
nor U3694 (N_3694,N_1295,N_1044);
and U3695 (N_3695,N_237,N_2616);
nand U3696 (N_3696,N_2601,N_860);
nand U3697 (N_3697,N_672,N_2551);
and U3698 (N_3698,N_1362,N_18);
or U3699 (N_3699,N_1719,N_371);
nor U3700 (N_3700,N_2369,N_680);
and U3701 (N_3701,N_2380,N_1471);
and U3702 (N_3702,N_159,N_516);
and U3703 (N_3703,N_717,N_1092);
or U3704 (N_3704,N_387,N_854);
and U3705 (N_3705,N_2448,N_2811);
nand U3706 (N_3706,N_142,N_1641);
xor U3707 (N_3707,N_2487,N_1062);
xnor U3708 (N_3708,N_936,N_698);
or U3709 (N_3709,N_622,N_1413);
xnor U3710 (N_3710,N_2960,N_3100);
nor U3711 (N_3711,N_544,N_1540);
nor U3712 (N_3712,N_1980,N_1729);
nor U3713 (N_3713,N_433,N_1508);
or U3714 (N_3714,N_2358,N_1964);
xnor U3715 (N_3715,N_242,N_1615);
xnor U3716 (N_3716,N_2559,N_2221);
and U3717 (N_3717,N_1747,N_2274);
nor U3718 (N_3718,N_1768,N_1582);
or U3719 (N_3719,N_671,N_2724);
nor U3720 (N_3720,N_2151,N_1537);
or U3721 (N_3721,N_1232,N_3039);
nor U3722 (N_3722,N_2918,N_1361);
nand U3723 (N_3723,N_2680,N_41);
and U3724 (N_3724,N_1146,N_1023);
xor U3725 (N_3725,N_650,N_2349);
or U3726 (N_3726,N_2873,N_554);
nor U3727 (N_3727,N_348,N_2964);
or U3728 (N_3728,N_1238,N_890);
or U3729 (N_3729,N_1084,N_2973);
nor U3730 (N_3730,N_2718,N_2054);
and U3731 (N_3731,N_2457,N_2205);
xnor U3732 (N_3732,N_1968,N_774);
and U3733 (N_3733,N_91,N_848);
nor U3734 (N_3734,N_1419,N_1281);
or U3735 (N_3735,N_1981,N_2330);
or U3736 (N_3736,N_2793,N_2253);
and U3737 (N_3737,N_2958,N_1906);
nor U3738 (N_3738,N_628,N_466);
or U3739 (N_3739,N_968,N_2695);
or U3740 (N_3740,N_93,N_2172);
nor U3741 (N_3741,N_1822,N_1142);
nor U3742 (N_3742,N_2007,N_1859);
and U3743 (N_3743,N_2516,N_2651);
nand U3744 (N_3744,N_2351,N_2641);
nand U3745 (N_3745,N_1924,N_1668);
or U3746 (N_3746,N_2039,N_1291);
nand U3747 (N_3747,N_1676,N_1876);
nor U3748 (N_3748,N_2733,N_783);
or U3749 (N_3749,N_606,N_784);
xor U3750 (N_3750,N_2667,N_2413);
or U3751 (N_3751,N_1591,N_2916);
or U3752 (N_3752,N_1101,N_617);
nand U3753 (N_3753,N_56,N_2814);
nand U3754 (N_3754,N_2239,N_1034);
nor U3755 (N_3755,N_1513,N_1324);
nand U3756 (N_3756,N_2148,N_2758);
or U3757 (N_3757,N_2796,N_3058);
nor U3758 (N_3758,N_1075,N_1534);
nand U3759 (N_3759,N_1583,N_2476);
or U3760 (N_3760,N_841,N_2243);
and U3761 (N_3761,N_1477,N_2441);
nor U3762 (N_3762,N_963,N_2595);
or U3763 (N_3763,N_667,N_2081);
and U3764 (N_3764,N_2907,N_3119);
nor U3765 (N_3765,N_744,N_423);
and U3766 (N_3766,N_877,N_3028);
and U3767 (N_3767,N_94,N_1382);
nor U3768 (N_3768,N_480,N_676);
nand U3769 (N_3769,N_888,N_1767);
and U3770 (N_3770,N_2068,N_1468);
nor U3771 (N_3771,N_601,N_1512);
nor U3772 (N_3772,N_301,N_731);
xnor U3773 (N_3773,N_575,N_2332);
or U3774 (N_3774,N_1233,N_2562);
and U3775 (N_3775,N_313,N_279);
xor U3776 (N_3776,N_929,N_2293);
or U3777 (N_3777,N_790,N_1732);
nor U3778 (N_3778,N_1520,N_705);
or U3779 (N_3779,N_2682,N_2679);
nor U3780 (N_3780,N_2485,N_2241);
or U3781 (N_3781,N_3073,N_2119);
and U3782 (N_3782,N_749,N_1318);
or U3783 (N_3783,N_514,N_2626);
nor U3784 (N_3784,N_2943,N_981);
nor U3785 (N_3785,N_1711,N_1812);
or U3786 (N_3786,N_3103,N_2622);
or U3787 (N_3787,N_3030,N_174);
or U3788 (N_3788,N_33,N_1341);
nand U3789 (N_3789,N_1400,N_109);
and U3790 (N_3790,N_1511,N_3002);
and U3791 (N_3791,N_2865,N_153);
nor U3792 (N_3792,N_2871,N_57);
nor U3793 (N_3793,N_1760,N_2880);
or U3794 (N_3794,N_1893,N_3108);
or U3795 (N_3795,N_919,N_1258);
and U3796 (N_3796,N_118,N_988);
nor U3797 (N_3797,N_1833,N_2482);
and U3798 (N_3798,N_1384,N_2180);
nor U3799 (N_3799,N_1478,N_2316);
and U3800 (N_3800,N_2824,N_2799);
and U3801 (N_3801,N_826,N_2994);
nand U3802 (N_3802,N_1586,N_2012);
or U3803 (N_3803,N_1792,N_1391);
and U3804 (N_3804,N_562,N_781);
nor U3805 (N_3805,N_2050,N_627);
nor U3806 (N_3806,N_405,N_2173);
nand U3807 (N_3807,N_2987,N_494);
xor U3808 (N_3808,N_2502,N_2155);
nor U3809 (N_3809,N_2150,N_2395);
nand U3810 (N_3810,N_2347,N_1039);
nor U3811 (N_3811,N_401,N_2437);
nor U3812 (N_3812,N_644,N_1901);
nand U3813 (N_3813,N_2439,N_692);
nand U3814 (N_3814,N_1773,N_3014);
and U3815 (N_3815,N_998,N_2500);
nor U3816 (N_3816,N_2329,N_570);
nand U3817 (N_3817,N_262,N_2803);
or U3818 (N_3818,N_430,N_2665);
or U3819 (N_3819,N_2161,N_2928);
nor U3820 (N_3820,N_1762,N_3113);
and U3821 (N_3821,N_724,N_2894);
nand U3822 (N_3822,N_253,N_1021);
xnor U3823 (N_3823,N_1308,N_732);
nor U3824 (N_3824,N_2844,N_90);
xor U3825 (N_3825,N_2681,N_2854);
and U3826 (N_3826,N_201,N_355);
and U3827 (N_3827,N_1214,N_1161);
nor U3828 (N_3828,N_2578,N_955);
or U3829 (N_3829,N_1098,N_1130);
nor U3830 (N_3830,N_1375,N_921);
or U3831 (N_3831,N_2279,N_2168);
and U3832 (N_3832,N_2819,N_1305);
nand U3833 (N_3833,N_238,N_314);
or U3834 (N_3834,N_1699,N_114);
or U3835 (N_3835,N_1036,N_2108);
and U3836 (N_3836,N_548,N_923);
xor U3837 (N_3837,N_195,N_2305);
and U3838 (N_3838,N_1401,N_2713);
or U3839 (N_3839,N_1037,N_27);
or U3840 (N_3840,N_10,N_1750);
and U3841 (N_3841,N_1218,N_2672);
nor U3842 (N_3842,N_2472,N_1367);
xnor U3843 (N_3843,N_2655,N_1445);
and U3844 (N_3844,N_1526,N_2137);
and U3845 (N_3845,N_20,N_1340);
and U3846 (N_3846,N_2742,N_546);
and U3847 (N_3847,N_1679,N_2043);
or U3848 (N_3848,N_1650,N_2761);
nor U3849 (N_3849,N_167,N_1786);
nor U3850 (N_3850,N_1861,N_2859);
nor U3851 (N_3851,N_2058,N_317);
and U3852 (N_3852,N_2036,N_281);
nand U3853 (N_3853,N_695,N_1089);
and U3854 (N_3854,N_1950,N_2246);
or U3855 (N_3855,N_1531,N_1761);
nor U3856 (N_3856,N_794,N_1135);
nand U3857 (N_3857,N_1848,N_2079);
and U3858 (N_3858,N_1932,N_2265);
nor U3859 (N_3859,N_2343,N_663);
xnor U3860 (N_3860,N_2805,N_2510);
xnor U3861 (N_3861,N_332,N_1239);
nor U3862 (N_3862,N_1995,N_1020);
nor U3863 (N_3863,N_1602,N_855);
or U3864 (N_3864,N_2357,N_1697);
nor U3865 (N_3865,N_726,N_1755);
nand U3866 (N_3866,N_1936,N_0);
nor U3867 (N_3867,N_1934,N_359);
nor U3868 (N_3868,N_2250,N_3106);
nand U3869 (N_3869,N_2451,N_2378);
or U3870 (N_3870,N_1782,N_2581);
nand U3871 (N_3871,N_675,N_88);
and U3872 (N_3872,N_296,N_1266);
nand U3873 (N_3873,N_376,N_1337);
nand U3874 (N_3874,N_3072,N_55);
and U3875 (N_3875,N_1955,N_2589);
nor U3876 (N_3876,N_1474,N_1565);
xor U3877 (N_3877,N_521,N_2678);
and U3878 (N_3878,N_217,N_928);
and U3879 (N_3879,N_2273,N_1723);
nor U3880 (N_3880,N_1184,N_2535);
and U3881 (N_3881,N_2795,N_182);
nor U3882 (N_3882,N_1643,N_1575);
and U3883 (N_3883,N_531,N_2088);
nor U3884 (N_3884,N_1494,N_756);
nand U3885 (N_3885,N_2342,N_1331);
or U3886 (N_3886,N_1975,N_1960);
and U3887 (N_3887,N_1335,N_876);
nand U3888 (N_3888,N_2744,N_1594);
or U3889 (N_3889,N_2344,N_791);
or U3890 (N_3890,N_2524,N_468);
or U3891 (N_3891,N_3011,N_2755);
nor U3892 (N_3892,N_2585,N_154);
and U3893 (N_3893,N_2084,N_2328);
nand U3894 (N_3894,N_611,N_2208);
nor U3895 (N_3895,N_139,N_2445);
nor U3896 (N_3896,N_558,N_17);
nor U3897 (N_3897,N_335,N_2390);
or U3898 (N_3898,N_727,N_1573);
or U3899 (N_3899,N_2019,N_3110);
or U3900 (N_3900,N_35,N_780);
xnor U3901 (N_3901,N_2784,N_2563);
xor U3902 (N_3902,N_1078,N_643);
nand U3903 (N_3903,N_1553,N_2720);
nand U3904 (N_3904,N_1670,N_60);
or U3905 (N_3905,N_1552,N_2541);
nor U3906 (N_3906,N_1309,N_13);
nand U3907 (N_3907,N_1440,N_1328);
nor U3908 (N_3908,N_984,N_1355);
nor U3909 (N_3909,N_1545,N_502);
nand U3910 (N_3910,N_1923,N_2566);
or U3911 (N_3911,N_1116,N_1624);
nor U3912 (N_3912,N_2953,N_879);
xor U3913 (N_3913,N_975,N_1454);
nand U3914 (N_3914,N_1104,N_1709);
and U3915 (N_3915,N_2552,N_1442);
nand U3916 (N_3916,N_2227,N_1658);
xnor U3917 (N_3917,N_2397,N_510);
nand U3918 (N_3918,N_1053,N_776);
nand U3919 (N_3919,N_145,N_2948);
nand U3920 (N_3920,N_2514,N_461);
and U3921 (N_3921,N_561,N_2195);
nor U3922 (N_3922,N_2666,N_2278);
and U3923 (N_3923,N_584,N_80);
and U3924 (N_3924,N_2624,N_1354);
nor U3925 (N_3925,N_1172,N_619);
nand U3926 (N_3926,N_2992,N_1406);
and U3927 (N_3927,N_3008,N_985);
and U3928 (N_3928,N_1299,N_2870);
or U3929 (N_3929,N_808,N_1979);
nand U3930 (N_3930,N_493,N_1255);
nor U3931 (N_3931,N_2949,N_2114);
and U3932 (N_3932,N_1374,N_497);
xnor U3933 (N_3933,N_1486,N_1107);
nand U3934 (N_3934,N_347,N_2294);
nor U3935 (N_3935,N_2255,N_312);
nand U3936 (N_3936,N_1657,N_2630);
and U3937 (N_3937,N_330,N_858);
xor U3938 (N_3938,N_1231,N_315);
nor U3939 (N_3939,N_2534,N_1077);
nor U3940 (N_3940,N_2565,N_2932);
or U3941 (N_3941,N_379,N_2956);
nor U3942 (N_3942,N_1825,N_2866);
nand U3943 (N_3943,N_2951,N_2625);
and U3944 (N_3944,N_2885,N_954);
xnor U3945 (N_3945,N_1052,N_2477);
and U3946 (N_3946,N_827,N_100);
or U3947 (N_3947,N_1289,N_1422);
or U3948 (N_3948,N_752,N_2414);
or U3949 (N_3949,N_535,N_2353);
nor U3950 (N_3950,N_490,N_2669);
or U3951 (N_3951,N_2606,N_730);
xnor U3952 (N_3952,N_287,N_1857);
or U3953 (N_3953,N_1533,N_448);
xnor U3954 (N_3954,N_1141,N_836);
nor U3955 (N_3955,N_2804,N_940);
nand U3956 (N_3956,N_2456,N_2619);
xor U3957 (N_3957,N_2846,N_165);
and U3958 (N_3958,N_2185,N_2051);
nand U3959 (N_3959,N_2745,N_1195);
nand U3960 (N_3960,N_738,N_2558);
nand U3961 (N_3961,N_2816,N_333);
and U3962 (N_3962,N_2284,N_2400);
nor U3963 (N_3963,N_2855,N_640);
nand U3964 (N_3964,N_624,N_996);
nand U3965 (N_3965,N_334,N_327);
nand U3966 (N_3966,N_1917,N_1612);
or U3967 (N_3967,N_559,N_1201);
and U3968 (N_3968,N_1073,N_1842);
xnor U3969 (N_3969,N_11,N_220);
xnor U3970 (N_3970,N_2576,N_2954);
or U3971 (N_3971,N_1514,N_79);
xnor U3972 (N_3972,N_2247,N_2825);
nor U3973 (N_3973,N_48,N_2149);
or U3974 (N_3974,N_1609,N_1253);
nand U3975 (N_3975,N_1991,N_3044);
and U3976 (N_3976,N_1997,N_9);
nand U3977 (N_3977,N_1001,N_2620);
or U3978 (N_3978,N_2363,N_3059);
or U3979 (N_3979,N_816,N_1286);
and U3980 (N_3980,N_1055,N_1871);
nor U3981 (N_3981,N_1065,N_1378);
nor U3982 (N_3982,N_2034,N_1630);
or U3983 (N_3983,N_1064,N_820);
or U3984 (N_3984,N_1427,N_2199);
or U3985 (N_3985,N_1158,N_1038);
nor U3986 (N_3986,N_3060,N_286);
nand U3987 (N_3987,N_412,N_1364);
nand U3988 (N_3988,N_1005,N_2734);
nand U3989 (N_3989,N_2097,N_2699);
nor U3990 (N_3990,N_3034,N_1578);
nor U3991 (N_3991,N_2026,N_2654);
nand U3992 (N_3992,N_44,N_2269);
nor U3993 (N_3993,N_1467,N_1566);
and U3994 (N_3994,N_2436,N_2790);
and U3995 (N_3995,N_2821,N_1330);
nand U3996 (N_3996,N_1811,N_1189);
nor U3997 (N_3997,N_1646,N_2976);
nand U3998 (N_3998,N_179,N_2044);
nand U3999 (N_3999,N_2408,N_693);
nand U4000 (N_4000,N_1858,N_1715);
xor U4001 (N_4001,N_2299,N_2518);
and U4002 (N_4002,N_293,N_1686);
or U4003 (N_4003,N_1423,N_2809);
and U4004 (N_4004,N_3071,N_3033);
nor U4005 (N_4005,N_1220,N_2033);
and U4006 (N_4006,N_2732,N_2759);
or U4007 (N_4007,N_2990,N_144);
nor U4008 (N_4008,N_1874,N_1941);
or U4009 (N_4009,N_1072,N_1249);
nand U4010 (N_4010,N_2640,N_2937);
or U4011 (N_4011,N_2860,N_2392);
nand U4012 (N_4012,N_1698,N_419);
nand U4013 (N_4013,N_1320,N_498);
nand U4014 (N_4014,N_1088,N_595);
or U4015 (N_4015,N_1720,N_658);
nand U4016 (N_4016,N_700,N_2339);
xor U4017 (N_4017,N_3079,N_46);
or U4018 (N_4018,N_2599,N_1854);
or U4019 (N_4019,N_2417,N_3029);
xnor U4020 (N_4020,N_1311,N_2530);
and U4021 (N_4021,N_73,N_1333);
nor U4022 (N_4022,N_1178,N_2509);
or U4023 (N_4023,N_1674,N_473);
xor U4024 (N_4024,N_2554,N_864);
nor U4025 (N_4025,N_2756,N_1000);
nor U4026 (N_4026,N_1775,N_440);
or U4027 (N_4027,N_1028,N_3085);
nand U4028 (N_4028,N_1031,N_3084);
and U4029 (N_4029,N_421,N_2481);
nor U4030 (N_4030,N_853,N_384);
or U4031 (N_4031,N_1887,N_979);
nor U4032 (N_4032,N_2920,N_464);
nor U4033 (N_4033,N_1765,N_229);
nand U4034 (N_4034,N_2603,N_2429);
and U4035 (N_4035,N_3018,N_1302);
nand U4036 (N_4036,N_2107,N_1702);
nor U4037 (N_4037,N_958,N_124);
nand U4038 (N_4038,N_2319,N_679);
nand U4039 (N_4039,N_501,N_316);
xnor U4040 (N_4040,N_260,N_880);
nand U4041 (N_4041,N_2881,N_210);
and U4042 (N_4042,N_1263,N_2132);
nor U4043 (N_4043,N_492,N_59);
or U4044 (N_4044,N_2741,N_2746);
xnor U4045 (N_4045,N_2830,N_400);
or U4046 (N_4046,N_2042,N_239);
nand U4047 (N_4047,N_1487,N_2262);
or U4048 (N_4048,N_912,N_1519);
nand U4049 (N_4049,N_26,N_1273);
or U4050 (N_4050,N_1389,N_1168);
or U4051 (N_4051,N_1110,N_2176);
and U4052 (N_4052,N_1143,N_3076);
or U4053 (N_4053,N_2468,N_863);
nor U4054 (N_4054,N_1701,N_1332);
nor U4055 (N_4055,N_1127,N_778);
nand U4056 (N_4056,N_2074,N_2432);
and U4057 (N_4057,N_2504,N_488);
nor U4058 (N_4058,N_207,N_1313);
nor U4059 (N_4059,N_633,N_959);
nor U4060 (N_4060,N_1136,N_2202);
nand U4061 (N_4061,N_275,N_835);
nand U4062 (N_4062,N_612,N_2366);
nand U4063 (N_4063,N_1282,N_1173);
or U4064 (N_4064,N_1967,N_2060);
nand U4065 (N_4065,N_491,N_1185);
or U4066 (N_4066,N_443,N_1497);
or U4067 (N_4067,N_2643,N_1986);
nor U4068 (N_4068,N_2505,N_1230);
nor U4069 (N_4069,N_2219,N_2145);
nand U4070 (N_4070,N_2571,N_2586);
nor U4071 (N_4071,N_2800,N_894);
or U4072 (N_4072,N_373,N_1714);
and U4073 (N_4073,N_1570,N_2192);
nand U4074 (N_4074,N_2120,N_1787);
or U4075 (N_4075,N_656,N_976);
or U4076 (N_4076,N_3022,N_2071);
xor U4077 (N_4077,N_1315,N_1946);
or U4078 (N_4078,N_1577,N_2688);
nor U4079 (N_4079,N_32,N_234);
or U4080 (N_4080,N_2355,N_1466);
and U4081 (N_4081,N_1560,N_2864);
nor U4082 (N_4082,N_1456,N_2223);
xor U4083 (N_4083,N_2095,N_148);
nor U4084 (N_4084,N_121,N_1360);
or U4085 (N_4085,N_1338,N_1507);
and U4086 (N_4086,N_2879,N_1428);
xnor U4087 (N_4087,N_2567,N_342);
nand U4088 (N_4088,N_245,N_518);
or U4089 (N_4089,N_714,N_2689);
nor U4090 (N_4090,N_2410,N_1707);
nor U4091 (N_4091,N_1260,N_290);
xor U4092 (N_4092,N_1082,N_1008);
nand U4093 (N_4093,N_1708,N_1605);
and U4094 (N_4094,N_246,N_1872);
nand U4095 (N_4095,N_3010,N_688);
nand U4096 (N_4096,N_300,N_350);
xor U4097 (N_4097,N_2144,N_163);
and U4098 (N_4098,N_1197,N_2590);
and U4099 (N_4099,N_1226,N_647);
xnor U4100 (N_4100,N_1011,N_364);
xnor U4101 (N_4101,N_137,N_2009);
and U4102 (N_4102,N_1126,N_2921);
or U4103 (N_4103,N_1090,N_3067);
nand U4104 (N_4104,N_1911,N_1204);
nor U4105 (N_4105,N_1431,N_834);
and U4106 (N_4106,N_2818,N_249);
nor U4107 (N_4107,N_2849,N_737);
nor U4108 (N_4108,N_993,N_3027);
xnor U4109 (N_4109,N_542,N_539);
nor U4110 (N_4110,N_2646,N_933);
or U4111 (N_4111,N_2196,N_4);
nand U4112 (N_4112,N_1673,N_1903);
or U4113 (N_4113,N_768,N_2187);
xnor U4114 (N_4114,N_1121,N_775);
nand U4115 (N_4115,N_2418,N_2082);
nor U4116 (N_4116,N_1685,N_1259);
nand U4117 (N_4117,N_428,N_107);
or U4118 (N_4118,N_1409,N_2989);
xor U4119 (N_4119,N_2867,N_621);
nand U4120 (N_4120,N_112,N_875);
and U4121 (N_4121,N_1493,N_2449);
or U4122 (N_4122,N_2707,N_2031);
nor U4123 (N_4123,N_895,N_1558);
xnor U4124 (N_4124,N_1035,N_185);
and U4125 (N_4125,N_1436,N_2115);
nand U4126 (N_4126,N_2368,N_792);
xnor U4127 (N_4127,N_3116,N_3040);
or U4128 (N_4128,N_1256,N_462);
and U4129 (N_4129,N_2549,N_2782);
and U4130 (N_4130,N_1032,N_511);
or U4131 (N_4131,N_2875,N_583);
and U4132 (N_4132,N_2446,N_2513);
nand U4133 (N_4133,N_92,N_2543);
or U4134 (N_4134,N_1951,N_1692);
or U4135 (N_4135,N_1002,N_2862);
and U4136 (N_4136,N_1688,N_1722);
and U4137 (N_4137,N_2116,N_352);
nand U4138 (N_4138,N_194,N_747);
xnor U4139 (N_4139,N_1004,N_256);
and U4140 (N_4140,N_802,N_3013);
xor U4141 (N_4141,N_1831,N_3086);
nor U4142 (N_4142,N_125,N_2915);
or U4143 (N_4143,N_2934,N_980);
or U4144 (N_4144,N_1788,N_1783);
xor U4145 (N_4145,N_2911,N_576);
nand U4146 (N_4146,N_3057,N_2281);
or U4147 (N_4147,N_1329,N_2999);
xnor U4148 (N_4148,N_769,N_935);
and U4149 (N_4149,N_2434,N_2608);
xor U4150 (N_4150,N_86,N_2750);
xnor U4151 (N_4151,N_522,N_308);
xnor U4152 (N_4152,N_2568,N_2868);
nor U4153 (N_4153,N_2431,N_893);
or U4154 (N_4154,N_2555,N_1272);
or U4155 (N_4155,N_2786,N_439);
or U4156 (N_4156,N_1794,N_2933);
nand U4157 (N_4157,N_2406,N_1434);
or U4158 (N_4158,N_1114,N_2387);
or U4159 (N_4159,N_101,N_652);
or U4160 (N_4160,N_1472,N_416);
and U4161 (N_4161,N_489,N_203);
xor U4162 (N_4162,N_143,N_1801);
and U4163 (N_4163,N_1734,N_295);
xor U4164 (N_4164,N_3006,N_3104);
and U4165 (N_4165,N_441,N_630);
nor U4166 (N_4166,N_666,N_187);
xnor U4167 (N_4167,N_398,N_1342);
or U4168 (N_4168,N_1628,N_1931);
nand U4169 (N_4169,N_251,N_1503);
and U4170 (N_4170,N_1298,N_2511);
nand U4171 (N_4171,N_3087,N_2171);
nand U4172 (N_4172,N_2191,N_3042);
or U4173 (N_4173,N_399,N_1860);
nand U4174 (N_4174,N_620,N_843);
nor U4175 (N_4175,N_1192,N_486);
nand U4176 (N_4176,N_1388,N_2454);
xor U4177 (N_4177,N_2981,N_2209);
nand U4178 (N_4178,N_2763,N_582);
nor U4179 (N_4179,N_2174,N_765);
nand U4180 (N_4180,N_446,N_1349);
nor U4181 (N_4181,N_156,N_2812);
or U4182 (N_4182,N_2673,N_1393);
or U4183 (N_4183,N_503,N_1969);
and U4184 (N_4184,N_2584,N_2597);
xnor U4185 (N_4185,N_1554,N_3093);
and U4186 (N_4186,N_934,N_344);
nor U4187 (N_4187,N_222,N_651);
xor U4188 (N_4188,N_898,N_1306);
nand U4189 (N_4189,N_2802,N_2717);
nor U4190 (N_4190,N_2017,N_2396);
and U4191 (N_4191,N_1790,N_2123);
and U4192 (N_4192,N_901,N_2104);
nor U4193 (N_4193,N_2982,N_2633);
xor U4194 (N_4194,N_1321,N_1808);
nor U4195 (N_4195,N_2315,N_2272);
or U4196 (N_4196,N_684,N_2737);
nor U4197 (N_4197,N_805,N_1100);
nor U4198 (N_4198,N_706,N_2183);
or U4199 (N_4199,N_2433,N_1254);
and U4200 (N_4200,N_75,N_2494);
and U4201 (N_4201,N_429,N_1677);
and U4202 (N_4202,N_900,N_1490);
or U4203 (N_4203,N_1464,N_1800);
nand U4204 (N_4204,N_2484,N_1700);
and U4205 (N_4205,N_2936,N_2810);
or U4206 (N_4206,N_2938,N_2190);
nor U4207 (N_4207,N_1390,N_1662);
and U4208 (N_4208,N_728,N_687);
nor U4209 (N_4209,N_1648,N_297);
nand U4210 (N_4210,N_1343,N_1631);
and U4211 (N_4211,N_654,N_319);
nand U4212 (N_4212,N_2304,N_3107);
or U4213 (N_4213,N_866,N_366);
nor U4214 (N_4214,N_1278,N_1819);
or U4215 (N_4215,N_1433,N_1461);
nor U4216 (N_4216,N_2101,N_1965);
nand U4217 (N_4217,N_2236,N_2235);
xnor U4218 (N_4218,N_3037,N_2876);
or U4219 (N_4219,N_753,N_2497);
nand U4220 (N_4220,N_2469,N_602);
nand U4221 (N_4221,N_70,N_694);
nand U4222 (N_4222,N_309,N_149);
xnor U4223 (N_4223,N_1982,N_289);
or U4224 (N_4224,N_596,N_1370);
nor U4225 (N_4225,N_417,N_478);
and U4226 (N_4226,N_1580,N_1448);
or U4227 (N_4227,N_938,N_2656);
and U4228 (N_4228,N_1252,N_2975);
or U4229 (N_4229,N_1186,N_432);
nor U4230 (N_4230,N_1372,N_2143);
nor U4231 (N_4231,N_541,N_1866);
nand U4232 (N_4232,N_1200,N_1581);
or U4233 (N_4233,N_1502,N_2372);
nand U4234 (N_4234,N_2442,N_2341);
nor U4235 (N_4235,N_2166,N_1543);
and U4236 (N_4236,N_1780,N_1465);
nand U4237 (N_4237,N_2029,N_445);
or U4238 (N_4238,N_1415,N_1826);
xor U4239 (N_4239,N_2946,N_807);
and U4240 (N_4240,N_2869,N_1518);
nand U4241 (N_4241,N_506,N_903);
xor U4242 (N_4242,N_1153,N_283);
and U4243 (N_4243,N_1603,N_2229);
nor U4244 (N_4244,N_3048,N_1165);
and U4245 (N_4245,N_500,N_2075);
xnor U4246 (N_4246,N_1610,N_1879);
or U4247 (N_4247,N_613,N_1429);
or U4248 (N_4248,N_2251,N_593);
and U4249 (N_4249,N_2785,N_1611);
or U4250 (N_4250,N_2495,N_1962);
and U4251 (N_4251,N_1524,N_282);
or U4252 (N_4252,N_2895,N_777);
nor U4253 (N_4253,N_211,N_2931);
nor U4254 (N_4254,N_2466,N_255);
nand U4255 (N_4255,N_2136,N_657);
nand U4256 (N_4256,N_1994,N_1873);
xor U4257 (N_4257,N_2539,N_2045);
nand U4258 (N_4258,N_2788,N_2360);
nand U4259 (N_4259,N_1713,N_2839);
and U4260 (N_4260,N_704,N_495);
nor U4261 (N_4261,N_278,N_846);
nand U4262 (N_4262,N_648,N_2798);
and U4263 (N_4263,N_1029,N_589);
or U4264 (N_4264,N_1798,N_939);
or U4265 (N_4265,N_1105,N_1919);
and U4266 (N_4266,N_2925,N_1725);
xor U4267 (N_4267,N_937,N_146);
xnor U4268 (N_4268,N_1900,N_2512);
nand U4269 (N_4269,N_2686,N_2573);
and U4270 (N_4270,N_922,N_1124);
nor U4271 (N_4271,N_1368,N_1693);
or U4272 (N_4272,N_1300,N_815);
and U4273 (N_4273,N_2326,N_1928);
nor U4274 (N_4274,N_1279,N_337);
or U4275 (N_4275,N_2612,N_2636);
nor U4276 (N_4276,N_2046,N_1804);
nor U4277 (N_4277,N_508,N_669);
nand U4278 (N_4278,N_3054,N_2317);
and U4279 (N_4279,N_2764,N_1322);
nor U4280 (N_4280,N_1043,N_588);
nor U4281 (N_4281,N_1275,N_2658);
or U4282 (N_4282,N_2311,N_2303);
or U4283 (N_4283,N_177,N_1009);
nor U4284 (N_4284,N_850,N_965);
or U4285 (N_4285,N_2781,N_1458);
nor U4286 (N_4286,N_1532,N_2739);
nor U4287 (N_4287,N_852,N_1210);
nor U4288 (N_4288,N_512,N_1139);
xnor U4289 (N_4289,N_2703,N_3114);
or U4290 (N_4290,N_1510,N_1426);
nand U4291 (N_4291,N_1250,N_2252);
nor U4292 (N_4292,N_1957,N_759);
and U4293 (N_4293,N_326,N_2133);
or U4294 (N_4294,N_2141,N_636);
nand U4295 (N_4295,N_374,N_3021);
nor U4296 (N_4296,N_252,N_2735);
xor U4297 (N_4297,N_1097,N_1791);
nor U4298 (N_4298,N_1666,N_1040);
and U4299 (N_4299,N_1935,N_2838);
and U4300 (N_4300,N_1449,N_2313);
nand U4301 (N_4301,N_385,N_892);
and U4302 (N_4302,N_3097,N_1929);
and U4303 (N_4303,N_586,N_703);
nor U4304 (N_4304,N_1219,N_340);
nor U4305 (N_4305,N_909,N_2152);
nand U4306 (N_4306,N_3051,N_1915);
nor U4307 (N_4307,N_748,N_1651);
nor U4308 (N_4308,N_3070,N_605);
xnor U4309 (N_4309,N_1194,N_2065);
or U4310 (N_4310,N_1886,N_2421);
and U4311 (N_4311,N_615,N_1432);
nor U4312 (N_4312,N_395,N_2371);
and U4313 (N_4313,N_2726,N_1042);
nor U4314 (N_4314,N_851,N_2706);
nor U4315 (N_4315,N_1460,N_191);
nor U4316 (N_4316,N_2277,N_2159);
and U4317 (N_4317,N_557,N_1850);
and U4318 (N_4318,N_3032,N_1469);
or U4319 (N_4319,N_380,N_2540);
and U4320 (N_4320,N_1753,N_2888);
nand U4321 (N_4321,N_302,N_824);
or U4322 (N_4322,N_1086,N_3118);
and U4323 (N_4323,N_2923,N_1159);
and U4324 (N_4324,N_353,N_767);
or U4325 (N_4325,N_422,N_772);
xor U4326 (N_4326,N_637,N_2383);
or U4327 (N_4327,N_2628,N_2664);
or U4328 (N_4328,N_178,N_2335);
or U4329 (N_4329,N_3082,N_1846);
xor U4330 (N_4330,N_1235,N_2962);
nand U4331 (N_4331,N_1131,N_241);
or U4332 (N_4332,N_1559,N_2945);
nor U4333 (N_4333,N_580,N_686);
and U4334 (N_4334,N_2310,N_2098);
nor U4335 (N_4335,N_116,N_997);
or U4336 (N_4336,N_434,N_2093);
nor U4337 (N_4337,N_574,N_1125);
nand U4338 (N_4338,N_3005,N_1444);
xnor U4339 (N_4339,N_2572,N_870);
nand U4340 (N_4340,N_2231,N_2526);
nand U4341 (N_4341,N_2712,N_1883);
nor U4342 (N_4342,N_1569,N_2685);
and U4343 (N_4343,N_1345,N_1974);
nand U4344 (N_4344,N_1894,N_1395);
or U4345 (N_4345,N_1117,N_1010);
nand U4346 (N_4346,N_2134,N_532);
nor U4347 (N_4347,N_673,N_323);
or U4348 (N_4348,N_831,N_2182);
and U4349 (N_4349,N_529,N_2389);
nor U4350 (N_4350,N_1307,N_1211);
and U4351 (N_4351,N_43,N_3020);
or U4352 (N_4352,N_2453,N_2905);
and U4353 (N_4353,N_1408,N_1455);
nand U4354 (N_4354,N_2470,N_2404);
nand U4355 (N_4355,N_2201,N_2085);
and U4356 (N_4356,N_38,N_1099);
nand U4357 (N_4357,N_2776,N_849);
nor U4358 (N_4358,N_1174,N_1703);
nor U4359 (N_4359,N_885,N_811);
or U4360 (N_4360,N_2189,N_1339);
and U4361 (N_4361,N_1550,N_891);
nor U4362 (N_4362,N_25,N_2532);
or U4363 (N_4363,N_2211,N_1443);
and U4364 (N_4364,N_1346,N_986);
nor U4365 (N_4365,N_2769,N_1498);
nor U4366 (N_4366,N_1424,N_3105);
xnor U4367 (N_4367,N_2267,N_2385);
nand U4368 (N_4368,N_476,N_1314);
nand U4369 (N_4369,N_720,N_1741);
or U4370 (N_4370,N_53,N_381);
nand U4371 (N_4371,N_1396,N_2099);
or U4372 (N_4372,N_573,N_1595);
nor U4373 (N_4373,N_2904,N_729);
and U4374 (N_4374,N_368,N_3031);
nand U4375 (N_4375,N_83,N_2978);
nand U4376 (N_4376,N_2100,N_1522);
or U4377 (N_4377,N_2254,N_2077);
nand U4378 (N_4378,N_2069,N_2376);
and U4379 (N_4379,N_1632,N_2248);
nor U4380 (N_4380,N_509,N_1205);
or U4381 (N_4381,N_626,N_1717);
nand U4382 (N_4382,N_1076,N_974);
and U4383 (N_4383,N_1284,N_1847);
nor U4384 (N_4384,N_1050,N_1119);
and U4385 (N_4385,N_1411,N_2730);
xor U4386 (N_4386,N_2743,N_1057);
nor U4387 (N_4387,N_1206,N_2447);
nand U4388 (N_4388,N_1156,N_1243);
and U4389 (N_4389,N_1597,N_614);
nor U4390 (N_4390,N_2096,N_722);
nand U4391 (N_4391,N_161,N_2906);
xor U4392 (N_4392,N_2729,N_372);
nand U4393 (N_4393,N_483,N_2266);
nand U4394 (N_4394,N_828,N_2207);
or U4395 (N_4395,N_1049,N_927);
xnor U4396 (N_4396,N_2346,N_537);
and U4397 (N_4397,N_2288,N_969);
and U4398 (N_4398,N_754,N_869);
and U4399 (N_4399,N_1678,N_1293);
or U4400 (N_4400,N_1353,N_2792);
and U4401 (N_4401,N_2475,N_1910);
nor U4402 (N_4402,N_2184,N_710);
nand U4403 (N_4403,N_592,N_164);
nor U4404 (N_4404,N_1989,N_1199);
or U4405 (N_4405,N_2259,N_1222);
nor U4406 (N_4406,N_475,N_2508);
nand U4407 (N_4407,N_1145,N_361);
nor U4408 (N_4408,N_259,N_2831);
and U4409 (N_4409,N_2290,N_1241);
nor U4410 (N_4410,N_2153,N_3075);
nor U4411 (N_4411,N_2030,N_1310);
or U4412 (N_4412,N_1129,N_1248);
nor U4413 (N_4413,N_2900,N_1027);
nand U4414 (N_4414,N_2258,N_2709);
or U4415 (N_4415,N_795,N_948);
and U4416 (N_4416,N_266,N_991);
nor U4417 (N_4417,N_1544,N_2322);
and U4418 (N_4418,N_2731,N_1644);
nand U4419 (N_4419,N_519,N_2550);
or U4420 (N_4420,N_2587,N_743);
xnor U4421 (N_4421,N_590,N_745);
nor U4422 (N_4422,N_982,N_274);
or U4423 (N_4423,N_307,N_994);
nor U4424 (N_4424,N_1071,N_2886);
and U4425 (N_4425,N_325,N_1687);
and U4426 (N_4426,N_435,N_2004);
nand U4427 (N_4427,N_2157,N_1485);
and U4428 (N_4428,N_587,N_707);
xnor U4429 (N_4429,N_1183,N_1690);
or U4430 (N_4430,N_757,N_1877);
nor U4431 (N_4431,N_964,N_1772);
or U4432 (N_4432,N_2117,N_1109);
or U4433 (N_4433,N_967,N_1681);
or U4434 (N_4434,N_2985,N_804);
and U4435 (N_4435,N_2280,N_1914);
xor U4436 (N_4436,N_1618,N_1240);
nor U4437 (N_4437,N_551,N_2289);
or U4438 (N_4438,N_1727,N_1890);
and U4439 (N_4439,N_2610,N_837);
or U4440 (N_4440,N_897,N_1224);
or U4441 (N_4441,N_1216,N_1654);
or U4442 (N_4442,N_1405,N_345);
or U4443 (N_4443,N_2591,N_1781);
nand U4444 (N_4444,N_365,N_1453);
or U4445 (N_4445,N_2878,N_1112);
or U4446 (N_4446,N_1181,N_181);
or U4447 (N_4447,N_674,N_523);
or U4448 (N_4448,N_751,N_1182);
and U4449 (N_4449,N_914,N_2362);
nor U4450 (N_4450,N_736,N_1169);
and U4451 (N_4451,N_538,N_1134);
and U4452 (N_4452,N_1081,N_1921);
or U4453 (N_4453,N_1592,N_2988);
nor U4454 (N_4454,N_393,N_196);
xor U4455 (N_4455,N_2697,N_1196);
nand U4456 (N_4456,N_162,N_788);
and U4457 (N_4457,N_2203,N_2507);
or U4458 (N_4458,N_147,N_1574);
nand U4459 (N_4459,N_1528,N_3115);
and U4460 (N_4460,N_2126,N_2950);
nand U4461 (N_4461,N_1938,N_133);
or U4462 (N_4462,N_1793,N_34);
xor U4463 (N_4463,N_1913,N_1404);
xor U4464 (N_4464,N_2971,N_2861);
nor U4465 (N_4465,N_2282,N_1208);
nand U4466 (N_4466,N_1344,N_244);
and U4467 (N_4467,N_2972,N_1771);
nand U4468 (N_4468,N_3063,N_3061);
xnor U4469 (N_4469,N_3012,N_1827);
xor U4470 (N_4470,N_2560,N_3049);
nor U4471 (N_4471,N_1267,N_924);
and U4472 (N_4472,N_941,N_762);
or U4473 (N_4473,N_629,N_2947);
nor U4474 (N_4474,N_318,N_896);
nand U4475 (N_4475,N_867,N_623);
nor U4476 (N_4476,N_2644,N_2683);
xnor U4477 (N_4477,N_213,N_1621);
or U4478 (N_4478,N_2411,N_1457);
nor U4479 (N_4479,N_1899,N_277);
nor U4480 (N_4480,N_442,N_2336);
nor U4481 (N_4481,N_2124,N_1601);
or U4482 (N_4482,N_2003,N_451);
nand U4483 (N_4483,N_2701,N_2415);
nand U4484 (N_4484,N_37,N_452);
xor U4485 (N_4485,N_1802,N_1691);
nand U4486 (N_4486,N_2052,N_2118);
or U4487 (N_4487,N_113,N_62);
nor U4488 (N_4488,N_3099,N_2780);
and U4489 (N_4489,N_2080,N_1625);
or U4490 (N_4490,N_1661,N_1633);
and U4491 (N_4491,N_2583,N_2464);
xor U4492 (N_4492,N_3025,N_8);
or U4493 (N_4493,N_2122,N_874);
nor U4494 (N_4494,N_1093,N_2693);
and U4495 (N_4495,N_1014,N_560);
or U4496 (N_4496,N_1155,N_105);
xnor U4497 (N_4497,N_1521,N_2426);
nor U4498 (N_4498,N_1163,N_1653);
nand U4499 (N_4499,N_971,N_2807);
nor U4500 (N_4500,N_978,N_2660);
or U4501 (N_4501,N_2835,N_358);
nor U4502 (N_4502,N_3080,N_1939);
nand U4503 (N_4503,N_2444,N_642);
nand U4504 (N_4504,N_645,N_1542);
xor U4505 (N_4505,N_2832,N_1120);
nand U4506 (N_4506,N_1865,N_1845);
and U4507 (N_4507,N_632,N_1551);
nand U4508 (N_4508,N_479,N_1386);
nor U4509 (N_4509,N_2023,N_1297);
xnor U4510 (N_4510,N_1007,N_3);
nor U4511 (N_4511,N_2977,N_2777);
and U4512 (N_4512,N_1147,N_383);
and U4513 (N_4513,N_2522,N_1489);
or U4514 (N_4514,N_65,N_2128);
or U4515 (N_4515,N_735,N_58);
nor U4516 (N_4516,N_1918,N_1738);
and U4517 (N_4517,N_2914,N_2090);
nand U4518 (N_4518,N_2194,N_1236);
nand U4519 (N_4519,N_2450,N_3007);
and U4520 (N_4520,N_1352,N_1614);
nand U4521 (N_4521,N_865,N_572);
xnor U4522 (N_4522,N_2323,N_2959);
xor U4523 (N_4523,N_2891,N_2047);
nand U4524 (N_4524,N_2092,N_1041);
nand U4525 (N_4525,N_2647,N_505);
nor U4526 (N_4526,N_2112,N_1138);
nand U4527 (N_4527,N_721,N_1659);
and U4528 (N_4528,N_545,N_2979);
nor U4529 (N_4529,N_507,N_63);
or U4530 (N_4530,N_1179,N_2066);
nor U4531 (N_4531,N_1025,N_472);
and U4532 (N_4532,N_1397,N_543);
xnor U4533 (N_4533,N_591,N_910);
xor U4534 (N_4534,N_1663,N_1988);
nand U4535 (N_4535,N_1358,N_2611);
nand U4536 (N_4536,N_840,N_235);
and U4537 (N_4537,N_2216,N_887);
or U4538 (N_4538,N_739,N_2650);
or U4539 (N_4539,N_1779,N_1496);
and U4540 (N_4540,N_1778,N_2361);
nor U4541 (N_4541,N_354,N_2271);
and U4542 (N_4542,N_2969,N_1113);
nor U4543 (N_4543,N_2598,N_861);
or U4544 (N_4544,N_2300,N_2032);
and U4545 (N_4545,N_1228,N_2008);
and U4546 (N_4546,N_1823,N_2596);
nand U4547 (N_4547,N_1108,N_2749);
or U4548 (N_4548,N_1851,N_103);
nand U4549 (N_4549,N_2225,N_2657);
and U4550 (N_4550,N_1916,N_215);
nand U4551 (N_4551,N_2214,N_718);
nor U4552 (N_4552,N_226,N_1907);
and U4553 (N_4553,N_1843,N_2064);
nand U4554 (N_4554,N_2517,N_1837);
nor U4555 (N_4555,N_369,N_1564);
and U4556 (N_4556,N_2244,N_329);
and U4557 (N_4557,N_1696,N_1047);
and U4558 (N_4558,N_2621,N_1818);
or U4559 (N_4559,N_2645,N_1133);
and U4560 (N_4560,N_2851,N_1530);
and U4561 (N_4561,N_1403,N_1265);
nand U4562 (N_4562,N_2815,N_2723);
nor U4563 (N_4563,N_1190,N_2452);
or U4564 (N_4564,N_2162,N_1144);
nor U4565 (N_4565,N_2350,N_1177);
nand U4566 (N_4566,N_2249,N_499);
and U4567 (N_4567,N_1561,N_581);
nor U4568 (N_4568,N_1111,N_987);
nand U4569 (N_4569,N_2897,N_1016);
nor U4570 (N_4570,N_1160,N_2307);
nand U4571 (N_4571,N_1304,N_3121);
and U4572 (N_4572,N_1737,N_782);
nor U4573 (N_4573,N_284,N_2929);
or U4574 (N_4574,N_661,N_990);
and U4575 (N_4575,N_3083,N_3015);
or U4576 (N_4576,N_1832,N_1803);
nand U4577 (N_4577,N_2694,N_713);
or U4578 (N_4578,N_3112,N_1834);
and U4579 (N_4579,N_471,N_2980);
or U4580 (N_4580,N_204,N_2285);
nor U4581 (N_4581,N_1680,N_2652);
and U4582 (N_4582,N_168,N_2638);
nor U4583 (N_4583,N_800,N_1350);
nor U4584 (N_4584,N_1947,N_7);
nand U4585 (N_4585,N_2613,N_2604);
nor U4586 (N_4586,N_2398,N_2525);
xnor U4587 (N_4587,N_973,N_2834);
and U4588 (N_4588,N_1751,N_2889);
and U4589 (N_4589,N_1587,N_1473);
nor U4590 (N_4590,N_1671,N_2966);
and U4591 (N_4591,N_906,N_1459);
nor U4592 (N_4592,N_517,N_3023);
xor U4593 (N_4593,N_298,N_2754);
or U4594 (N_4594,N_908,N_1535);
or U4595 (N_4595,N_814,N_2740);
nor U4596 (N_4596,N_2823,N_2738);
or U4597 (N_4597,N_407,N_1079);
nand U4598 (N_4598,N_2847,N_1446);
or U4599 (N_4599,N_683,N_670);
and U4600 (N_4600,N_3056,N_2501);
nor U4601 (N_4601,N_696,N_1067);
or U4602 (N_4602,N_346,N_437);
nor U4603 (N_4603,N_1735,N_1385);
and U4604 (N_4604,N_2334,N_2438);
nor U4605 (N_4605,N_1959,N_219);
or U4606 (N_4606,N_725,N_1326);
or U4607 (N_4607,N_2787,N_2001);
nor U4608 (N_4608,N_1054,N_2523);
and U4609 (N_4609,N_1290,N_2913);
nor U4610 (N_4610,N_2751,N_1416);
nand U4611 (N_4611,N_2345,N_568);
and U4612 (N_4612,N_1721,N_24);
nor U4613 (N_4613,N_1880,N_2963);
and U4614 (N_4614,N_469,N_779);
nor U4615 (N_4615,N_2292,N_305);
nand U4616 (N_4616,N_2725,N_1171);
nor U4617 (N_4617,N_99,N_1414);
nor U4618 (N_4618,N_2388,N_513);
nor U4619 (N_4619,N_1369,N_2178);
and U4620 (N_4620,N_186,N_1639);
or U4621 (N_4621,N_1904,N_2813);
nand U4622 (N_4622,N_2463,N_1807);
nor U4623 (N_4623,N_2515,N_2018);
nand U4624 (N_4624,N_410,N_2874);
nor U4625 (N_4625,N_2893,N_1327);
and U4626 (N_4626,N_1523,N_845);
xnor U4627 (N_4627,N_1905,N_2365);
nand U4628 (N_4628,N_1973,N_1590);
nor U4629 (N_4629,N_856,N_1869);
or U4630 (N_4630,N_2222,N_1607);
nand U4631 (N_4631,N_166,N_723);
nor U4632 (N_4632,N_1470,N_1970);
and U4633 (N_4633,N_770,N_2827);
or U4634 (N_4634,N_950,N_386);
or U4635 (N_4635,N_2035,N_2719);
nor U4636 (N_4636,N_2131,N_270);
or U4637 (N_4637,N_362,N_2912);
and U4638 (N_4638,N_1377,N_89);
or U4639 (N_4639,N_1059,N_594);
nand U4640 (N_4640,N_1961,N_1817);
nor U4641 (N_4641,N_2333,N_966);
and U4642 (N_4642,N_2986,N_160);
and U4643 (N_4643,N_1371,N_1742);
nor U4644 (N_4644,N_1274,N_960);
or U4645 (N_4645,N_1128,N_2260);
nand U4646 (N_4646,N_2409,N_526);
or U4647 (N_4647,N_1730,N_1984);
xnor U4648 (N_4648,N_1598,N_1571);
or U4649 (N_4649,N_1347,N_1849);
or U4650 (N_4650,N_1483,N_2600);
nand U4651 (N_4651,N_1074,N_838);
nor U4652 (N_4652,N_1412,N_1902);
nand U4653 (N_4653,N_1336,N_2490);
nor U4654 (N_4654,N_1756,N_525);
and U4655 (N_4655,N_920,N_1777);
xnor U4656 (N_4656,N_128,N_338);
or U4657 (N_4657,N_2722,N_962);
nand U4658 (N_4658,N_2424,N_2486);
nor U4659 (N_4659,N_2275,N_917);
or U4660 (N_4660,N_3074,N_2374);
or U4661 (N_4661,N_351,N_1572);
nand U4662 (N_4662,N_110,N_2778);
and U4663 (N_4663,N_2705,N_1836);
xnor U4664 (N_4664,N_402,N_122);
nor U4665 (N_4665,N_454,N_825);
nor U4666 (N_4666,N_1450,N_30);
xnor U4667 (N_4667,N_2204,N_2276);
or U4668 (N_4668,N_1546,N_1418);
nand U4669 (N_4669,N_1187,N_254);
nand U4670 (N_4670,N_1608,N_2536);
nand U4671 (N_4671,N_2546,N_2146);
and U4672 (N_4672,N_902,N_600);
and U4673 (N_4673,N_862,N_81);
or U4674 (N_4674,N_1215,N_913);
and U4675 (N_4675,N_1407,N_1288);
and U4676 (N_4676,N_646,N_2059);
xnor U4677 (N_4677,N_2175,N_2306);
nor U4678 (N_4678,N_1203,N_1287);
and U4679 (N_4679,N_520,N_2774);
or U4680 (N_4680,N_2944,N_2110);
or U4681 (N_4681,N_2461,N_171);
nand U4682 (N_4682,N_265,N_152);
and U4683 (N_4683,N_1261,N_40);
nor U4684 (N_4684,N_1,N_2998);
or U4685 (N_4685,N_176,N_1264);
or U4686 (N_4686,N_224,N_1810);
nor U4687 (N_4687,N_2877,N_1242);
and U4688 (N_4688,N_2378,N_1636);
or U4689 (N_4689,N_2491,N_224);
nor U4690 (N_4690,N_2910,N_2196);
or U4691 (N_4691,N_1082,N_1579);
or U4692 (N_4692,N_1929,N_2472);
and U4693 (N_4693,N_715,N_1870);
or U4694 (N_4694,N_12,N_1233);
nand U4695 (N_4695,N_211,N_474);
nor U4696 (N_4696,N_3044,N_2243);
or U4697 (N_4697,N_2245,N_828);
nor U4698 (N_4698,N_2620,N_888);
nand U4699 (N_4699,N_1666,N_1102);
xnor U4700 (N_4700,N_1682,N_2156);
nor U4701 (N_4701,N_1938,N_1727);
xor U4702 (N_4702,N_1043,N_460);
and U4703 (N_4703,N_309,N_1038);
or U4704 (N_4704,N_3035,N_1148);
nand U4705 (N_4705,N_547,N_2325);
nand U4706 (N_4706,N_1881,N_2224);
or U4707 (N_4707,N_686,N_2520);
nand U4708 (N_4708,N_1797,N_801);
and U4709 (N_4709,N_2774,N_162);
nor U4710 (N_4710,N_676,N_1730);
and U4711 (N_4711,N_2968,N_291);
xnor U4712 (N_4712,N_1161,N_3118);
or U4713 (N_4713,N_2819,N_825);
or U4714 (N_4714,N_2355,N_2198);
nor U4715 (N_4715,N_2798,N_598);
and U4716 (N_4716,N_1351,N_2573);
or U4717 (N_4717,N_2436,N_629);
and U4718 (N_4718,N_2178,N_1062);
nand U4719 (N_4719,N_1517,N_2654);
and U4720 (N_4720,N_2242,N_1148);
nor U4721 (N_4721,N_422,N_2504);
nand U4722 (N_4722,N_379,N_1390);
nand U4723 (N_4723,N_1282,N_537);
and U4724 (N_4724,N_1011,N_278);
and U4725 (N_4725,N_1141,N_857);
nand U4726 (N_4726,N_207,N_1931);
xor U4727 (N_4727,N_1064,N_2144);
or U4728 (N_4728,N_2923,N_1826);
nand U4729 (N_4729,N_2760,N_1831);
xor U4730 (N_4730,N_887,N_1132);
xor U4731 (N_4731,N_1089,N_2536);
nand U4732 (N_4732,N_555,N_2661);
nor U4733 (N_4733,N_2350,N_1223);
or U4734 (N_4734,N_2041,N_810);
nand U4735 (N_4735,N_2538,N_2490);
or U4736 (N_4736,N_2025,N_2488);
and U4737 (N_4737,N_2327,N_973);
nor U4738 (N_4738,N_2028,N_1024);
nor U4739 (N_4739,N_1980,N_248);
or U4740 (N_4740,N_1113,N_3018);
and U4741 (N_4741,N_37,N_2583);
xnor U4742 (N_4742,N_937,N_1669);
nand U4743 (N_4743,N_1434,N_2417);
nor U4744 (N_4744,N_1967,N_788);
nor U4745 (N_4745,N_3081,N_1875);
or U4746 (N_4746,N_2130,N_3065);
or U4747 (N_4747,N_1466,N_53);
and U4748 (N_4748,N_1963,N_2947);
nor U4749 (N_4749,N_2047,N_2607);
and U4750 (N_4750,N_2509,N_2525);
or U4751 (N_4751,N_1144,N_501);
or U4752 (N_4752,N_2790,N_2077);
nand U4753 (N_4753,N_1636,N_1558);
nor U4754 (N_4754,N_329,N_1893);
or U4755 (N_4755,N_92,N_1095);
or U4756 (N_4756,N_2334,N_73);
xnor U4757 (N_4757,N_1650,N_890);
or U4758 (N_4758,N_2765,N_998);
nor U4759 (N_4759,N_1010,N_2469);
nor U4760 (N_4760,N_2031,N_446);
or U4761 (N_4761,N_118,N_204);
nand U4762 (N_4762,N_573,N_701);
nand U4763 (N_4763,N_635,N_1942);
nor U4764 (N_4764,N_2533,N_2401);
nand U4765 (N_4765,N_2812,N_545);
or U4766 (N_4766,N_604,N_1203);
nand U4767 (N_4767,N_3104,N_405);
xnor U4768 (N_4768,N_2415,N_838);
or U4769 (N_4769,N_1138,N_1733);
nand U4770 (N_4770,N_1290,N_207);
nor U4771 (N_4771,N_2226,N_1177);
nor U4772 (N_4772,N_2480,N_1817);
and U4773 (N_4773,N_240,N_1660);
and U4774 (N_4774,N_25,N_231);
nand U4775 (N_4775,N_715,N_1483);
or U4776 (N_4776,N_1452,N_3108);
xor U4777 (N_4777,N_469,N_107);
nor U4778 (N_4778,N_602,N_2612);
or U4779 (N_4779,N_1732,N_1993);
nor U4780 (N_4780,N_499,N_2768);
nand U4781 (N_4781,N_1427,N_2015);
and U4782 (N_4782,N_111,N_1172);
nor U4783 (N_4783,N_1204,N_132);
or U4784 (N_4784,N_1574,N_1111);
nand U4785 (N_4785,N_2279,N_2593);
or U4786 (N_4786,N_215,N_1311);
nand U4787 (N_4787,N_1074,N_1593);
and U4788 (N_4788,N_1102,N_2372);
xor U4789 (N_4789,N_519,N_743);
or U4790 (N_4790,N_2489,N_1341);
nand U4791 (N_4791,N_2387,N_1622);
and U4792 (N_4792,N_2646,N_905);
xor U4793 (N_4793,N_58,N_630);
or U4794 (N_4794,N_179,N_355);
nand U4795 (N_4795,N_1310,N_568);
and U4796 (N_4796,N_2248,N_956);
nand U4797 (N_4797,N_538,N_1384);
and U4798 (N_4798,N_3092,N_1349);
nor U4799 (N_4799,N_716,N_1890);
or U4800 (N_4800,N_1171,N_248);
and U4801 (N_4801,N_872,N_1472);
nor U4802 (N_4802,N_1745,N_591);
or U4803 (N_4803,N_2161,N_2812);
nand U4804 (N_4804,N_2052,N_884);
nand U4805 (N_4805,N_379,N_1949);
nor U4806 (N_4806,N_2306,N_1873);
nor U4807 (N_4807,N_1983,N_2020);
nand U4808 (N_4808,N_1425,N_2548);
or U4809 (N_4809,N_2471,N_2644);
xnor U4810 (N_4810,N_510,N_1564);
nand U4811 (N_4811,N_142,N_1189);
nor U4812 (N_4812,N_2479,N_2011);
and U4813 (N_4813,N_2301,N_1866);
nor U4814 (N_4814,N_2323,N_2316);
and U4815 (N_4815,N_556,N_1295);
or U4816 (N_4816,N_1261,N_1138);
nor U4817 (N_4817,N_1565,N_2011);
nand U4818 (N_4818,N_3059,N_503);
and U4819 (N_4819,N_2650,N_2363);
and U4820 (N_4820,N_2126,N_2970);
or U4821 (N_4821,N_2741,N_626);
or U4822 (N_4822,N_2727,N_2566);
xor U4823 (N_4823,N_2666,N_621);
or U4824 (N_4824,N_2495,N_1327);
nor U4825 (N_4825,N_1934,N_786);
nand U4826 (N_4826,N_536,N_1961);
nor U4827 (N_4827,N_3079,N_925);
nor U4828 (N_4828,N_417,N_373);
nand U4829 (N_4829,N_3029,N_283);
xnor U4830 (N_4830,N_2096,N_1807);
nand U4831 (N_4831,N_637,N_1464);
nor U4832 (N_4832,N_2996,N_2360);
and U4833 (N_4833,N_1673,N_2409);
or U4834 (N_4834,N_783,N_1387);
and U4835 (N_4835,N_1623,N_421);
nor U4836 (N_4836,N_1805,N_1107);
nor U4837 (N_4837,N_1666,N_1534);
xnor U4838 (N_4838,N_1715,N_920);
and U4839 (N_4839,N_553,N_809);
nand U4840 (N_4840,N_1380,N_2646);
nand U4841 (N_4841,N_712,N_1515);
or U4842 (N_4842,N_1169,N_1028);
nor U4843 (N_4843,N_1004,N_2916);
and U4844 (N_4844,N_1225,N_1449);
and U4845 (N_4845,N_3084,N_2351);
nand U4846 (N_4846,N_2885,N_1875);
nor U4847 (N_4847,N_417,N_3120);
or U4848 (N_4848,N_2531,N_1836);
nor U4849 (N_4849,N_1707,N_1506);
and U4850 (N_4850,N_3117,N_33);
or U4851 (N_4851,N_2897,N_1396);
or U4852 (N_4852,N_2857,N_1787);
xor U4853 (N_4853,N_859,N_1376);
or U4854 (N_4854,N_967,N_1512);
or U4855 (N_4855,N_2759,N_646);
nand U4856 (N_4856,N_820,N_898);
and U4857 (N_4857,N_11,N_1088);
or U4858 (N_4858,N_2261,N_2270);
or U4859 (N_4859,N_2495,N_2433);
nand U4860 (N_4860,N_1086,N_2173);
nor U4861 (N_4861,N_1483,N_895);
nor U4862 (N_4862,N_1221,N_138);
or U4863 (N_4863,N_516,N_874);
nor U4864 (N_4864,N_1766,N_2086);
or U4865 (N_4865,N_2849,N_1598);
xnor U4866 (N_4866,N_146,N_1619);
nor U4867 (N_4867,N_1281,N_2428);
nor U4868 (N_4868,N_1512,N_2728);
nand U4869 (N_4869,N_2626,N_178);
or U4870 (N_4870,N_1765,N_1044);
and U4871 (N_4871,N_1845,N_1512);
nand U4872 (N_4872,N_2519,N_965);
nor U4873 (N_4873,N_1788,N_286);
or U4874 (N_4874,N_2384,N_1658);
nor U4875 (N_4875,N_2042,N_1435);
xor U4876 (N_4876,N_2022,N_3068);
or U4877 (N_4877,N_1224,N_1442);
and U4878 (N_4878,N_29,N_437);
and U4879 (N_4879,N_816,N_1058);
and U4880 (N_4880,N_842,N_1937);
or U4881 (N_4881,N_474,N_2490);
xor U4882 (N_4882,N_1118,N_3039);
or U4883 (N_4883,N_546,N_1848);
nor U4884 (N_4884,N_2419,N_3080);
nor U4885 (N_4885,N_2426,N_1081);
or U4886 (N_4886,N_2378,N_624);
nor U4887 (N_4887,N_3024,N_2161);
nand U4888 (N_4888,N_2154,N_723);
nor U4889 (N_4889,N_1880,N_2148);
nor U4890 (N_4890,N_2293,N_393);
nand U4891 (N_4891,N_2488,N_2841);
or U4892 (N_4892,N_315,N_1446);
nand U4893 (N_4893,N_1701,N_643);
or U4894 (N_4894,N_387,N_902);
nor U4895 (N_4895,N_981,N_610);
nand U4896 (N_4896,N_458,N_2560);
nand U4897 (N_4897,N_2619,N_2470);
nor U4898 (N_4898,N_3033,N_3097);
or U4899 (N_4899,N_790,N_994);
nand U4900 (N_4900,N_2736,N_1368);
nor U4901 (N_4901,N_1425,N_2389);
and U4902 (N_4902,N_1379,N_1638);
nor U4903 (N_4903,N_2666,N_2035);
nor U4904 (N_4904,N_424,N_2129);
or U4905 (N_4905,N_801,N_1477);
nor U4906 (N_4906,N_2108,N_2815);
or U4907 (N_4907,N_2028,N_2726);
and U4908 (N_4908,N_2400,N_2264);
and U4909 (N_4909,N_2905,N_2201);
xor U4910 (N_4910,N_2767,N_926);
or U4911 (N_4911,N_3082,N_2957);
nand U4912 (N_4912,N_2803,N_1090);
nand U4913 (N_4913,N_2033,N_1074);
nand U4914 (N_4914,N_3101,N_2845);
or U4915 (N_4915,N_947,N_1345);
xnor U4916 (N_4916,N_1565,N_66);
nand U4917 (N_4917,N_1635,N_2703);
nor U4918 (N_4918,N_1295,N_1183);
nand U4919 (N_4919,N_1731,N_151);
nor U4920 (N_4920,N_2287,N_2447);
and U4921 (N_4921,N_2553,N_1181);
or U4922 (N_4922,N_105,N_549);
or U4923 (N_4923,N_1968,N_43);
or U4924 (N_4924,N_1261,N_1190);
nor U4925 (N_4925,N_1741,N_2956);
nand U4926 (N_4926,N_707,N_1552);
nor U4927 (N_4927,N_1973,N_971);
or U4928 (N_4928,N_1054,N_1198);
nand U4929 (N_4929,N_1077,N_2240);
nor U4930 (N_4930,N_1925,N_412);
and U4931 (N_4931,N_240,N_1034);
and U4932 (N_4932,N_366,N_1093);
nor U4933 (N_4933,N_902,N_532);
and U4934 (N_4934,N_3056,N_2343);
and U4935 (N_4935,N_147,N_2658);
or U4936 (N_4936,N_2113,N_1031);
nand U4937 (N_4937,N_2257,N_2281);
or U4938 (N_4938,N_2061,N_602);
or U4939 (N_4939,N_285,N_287);
nor U4940 (N_4940,N_623,N_1032);
nand U4941 (N_4941,N_2655,N_2554);
and U4942 (N_4942,N_2162,N_830);
or U4943 (N_4943,N_2221,N_1015);
xnor U4944 (N_4944,N_1475,N_1301);
nor U4945 (N_4945,N_1833,N_731);
and U4946 (N_4946,N_452,N_2170);
and U4947 (N_4947,N_734,N_1688);
xor U4948 (N_4948,N_1604,N_2060);
xor U4949 (N_4949,N_1113,N_1676);
nor U4950 (N_4950,N_2201,N_203);
nor U4951 (N_4951,N_505,N_1222);
or U4952 (N_4952,N_2102,N_2939);
nand U4953 (N_4953,N_1970,N_1919);
nor U4954 (N_4954,N_2125,N_2977);
xnor U4955 (N_4955,N_1063,N_1832);
and U4956 (N_4956,N_2244,N_231);
and U4957 (N_4957,N_1900,N_2833);
nand U4958 (N_4958,N_1544,N_3012);
and U4959 (N_4959,N_2413,N_1163);
nor U4960 (N_4960,N_1533,N_2361);
xnor U4961 (N_4961,N_2490,N_518);
nand U4962 (N_4962,N_2965,N_1049);
nand U4963 (N_4963,N_2381,N_2819);
and U4964 (N_4964,N_663,N_973);
nand U4965 (N_4965,N_495,N_1213);
nand U4966 (N_4966,N_864,N_2139);
nand U4967 (N_4967,N_236,N_1245);
nor U4968 (N_4968,N_230,N_2855);
nand U4969 (N_4969,N_3001,N_504);
nor U4970 (N_4970,N_363,N_2457);
or U4971 (N_4971,N_756,N_1534);
and U4972 (N_4972,N_1087,N_1933);
nand U4973 (N_4973,N_1087,N_1103);
xnor U4974 (N_4974,N_2038,N_968);
and U4975 (N_4975,N_61,N_1752);
nand U4976 (N_4976,N_1938,N_2504);
nand U4977 (N_4977,N_2335,N_2038);
nand U4978 (N_4978,N_2462,N_897);
xnor U4979 (N_4979,N_1347,N_937);
nor U4980 (N_4980,N_2789,N_783);
or U4981 (N_4981,N_342,N_2309);
and U4982 (N_4982,N_1134,N_301);
or U4983 (N_4983,N_1339,N_792);
nand U4984 (N_4984,N_1414,N_104);
nor U4985 (N_4985,N_1447,N_2586);
nor U4986 (N_4986,N_1870,N_3061);
xor U4987 (N_4987,N_1922,N_1587);
and U4988 (N_4988,N_2725,N_1705);
nand U4989 (N_4989,N_2778,N_278);
nand U4990 (N_4990,N_564,N_1616);
xor U4991 (N_4991,N_1744,N_2594);
nand U4992 (N_4992,N_142,N_13);
nor U4993 (N_4993,N_2314,N_2232);
nor U4994 (N_4994,N_1513,N_825);
xnor U4995 (N_4995,N_2566,N_1455);
nor U4996 (N_4996,N_52,N_2848);
and U4997 (N_4997,N_2445,N_2740);
and U4998 (N_4998,N_491,N_2161);
or U4999 (N_4999,N_851,N_419);
or U5000 (N_5000,N_583,N_766);
and U5001 (N_5001,N_2831,N_425);
or U5002 (N_5002,N_1649,N_1572);
nand U5003 (N_5003,N_1293,N_2902);
or U5004 (N_5004,N_1963,N_1041);
or U5005 (N_5005,N_1518,N_782);
and U5006 (N_5006,N_849,N_1665);
nand U5007 (N_5007,N_2414,N_1906);
nor U5008 (N_5008,N_1725,N_911);
and U5009 (N_5009,N_2695,N_2642);
and U5010 (N_5010,N_1168,N_1103);
nand U5011 (N_5011,N_2208,N_400);
nand U5012 (N_5012,N_1017,N_2273);
xnor U5013 (N_5013,N_283,N_1645);
nand U5014 (N_5014,N_2715,N_1743);
xnor U5015 (N_5015,N_1584,N_2115);
nand U5016 (N_5016,N_419,N_2211);
nand U5017 (N_5017,N_735,N_1305);
nand U5018 (N_5018,N_1972,N_2441);
or U5019 (N_5019,N_293,N_384);
or U5020 (N_5020,N_951,N_1214);
nand U5021 (N_5021,N_2986,N_1290);
or U5022 (N_5022,N_1490,N_1445);
nand U5023 (N_5023,N_822,N_782);
nor U5024 (N_5024,N_2312,N_73);
xnor U5025 (N_5025,N_2173,N_1522);
or U5026 (N_5026,N_2650,N_1877);
or U5027 (N_5027,N_1610,N_843);
or U5028 (N_5028,N_3004,N_2315);
or U5029 (N_5029,N_1865,N_1663);
xnor U5030 (N_5030,N_514,N_2024);
xor U5031 (N_5031,N_1681,N_2663);
and U5032 (N_5032,N_487,N_237);
or U5033 (N_5033,N_2086,N_59);
nand U5034 (N_5034,N_1181,N_2030);
nor U5035 (N_5035,N_538,N_2747);
nand U5036 (N_5036,N_1962,N_1443);
nand U5037 (N_5037,N_2081,N_3018);
nand U5038 (N_5038,N_1832,N_1632);
nand U5039 (N_5039,N_1531,N_1550);
and U5040 (N_5040,N_2876,N_620);
nor U5041 (N_5041,N_2131,N_1714);
xor U5042 (N_5042,N_2343,N_1493);
nand U5043 (N_5043,N_3008,N_548);
and U5044 (N_5044,N_867,N_2313);
xor U5045 (N_5045,N_928,N_456);
xor U5046 (N_5046,N_1076,N_2524);
or U5047 (N_5047,N_2239,N_2043);
and U5048 (N_5048,N_213,N_2882);
and U5049 (N_5049,N_903,N_743);
nor U5050 (N_5050,N_220,N_3105);
nor U5051 (N_5051,N_2782,N_3026);
or U5052 (N_5052,N_519,N_165);
or U5053 (N_5053,N_2868,N_1924);
nor U5054 (N_5054,N_1864,N_2292);
nand U5055 (N_5055,N_1572,N_2407);
nand U5056 (N_5056,N_624,N_1920);
and U5057 (N_5057,N_1424,N_392);
nor U5058 (N_5058,N_3028,N_1437);
or U5059 (N_5059,N_531,N_1874);
xor U5060 (N_5060,N_1368,N_2350);
nand U5061 (N_5061,N_2340,N_2397);
nand U5062 (N_5062,N_1988,N_2730);
and U5063 (N_5063,N_543,N_1322);
or U5064 (N_5064,N_382,N_1227);
and U5065 (N_5065,N_72,N_1647);
xor U5066 (N_5066,N_2556,N_1985);
nand U5067 (N_5067,N_714,N_1003);
nand U5068 (N_5068,N_1764,N_2903);
nor U5069 (N_5069,N_2834,N_1893);
nor U5070 (N_5070,N_2337,N_775);
or U5071 (N_5071,N_2100,N_2516);
nor U5072 (N_5072,N_2670,N_2210);
nor U5073 (N_5073,N_2052,N_2175);
nand U5074 (N_5074,N_1868,N_1543);
or U5075 (N_5075,N_1934,N_993);
nor U5076 (N_5076,N_1377,N_2765);
and U5077 (N_5077,N_974,N_1250);
nand U5078 (N_5078,N_1005,N_643);
or U5079 (N_5079,N_875,N_688);
or U5080 (N_5080,N_213,N_678);
or U5081 (N_5081,N_2898,N_3004);
or U5082 (N_5082,N_2337,N_1978);
or U5083 (N_5083,N_2041,N_3078);
nand U5084 (N_5084,N_304,N_1435);
xor U5085 (N_5085,N_1543,N_3049);
nor U5086 (N_5086,N_2113,N_494);
nand U5087 (N_5087,N_900,N_1171);
nand U5088 (N_5088,N_2018,N_776);
nand U5089 (N_5089,N_1449,N_1722);
or U5090 (N_5090,N_1707,N_431);
nor U5091 (N_5091,N_1121,N_1509);
or U5092 (N_5092,N_1181,N_393);
and U5093 (N_5093,N_1596,N_2035);
nor U5094 (N_5094,N_42,N_457);
nand U5095 (N_5095,N_2097,N_660);
nor U5096 (N_5096,N_1367,N_2623);
nand U5097 (N_5097,N_2321,N_2853);
and U5098 (N_5098,N_1521,N_1718);
or U5099 (N_5099,N_564,N_1689);
or U5100 (N_5100,N_1285,N_1143);
nor U5101 (N_5101,N_1922,N_628);
and U5102 (N_5102,N_2641,N_2646);
or U5103 (N_5103,N_2769,N_1720);
and U5104 (N_5104,N_477,N_133);
or U5105 (N_5105,N_170,N_724);
and U5106 (N_5106,N_1346,N_2313);
nor U5107 (N_5107,N_1304,N_946);
or U5108 (N_5108,N_462,N_1804);
nand U5109 (N_5109,N_151,N_2414);
nor U5110 (N_5110,N_45,N_2431);
or U5111 (N_5111,N_2713,N_1079);
nand U5112 (N_5112,N_426,N_2818);
and U5113 (N_5113,N_1687,N_525);
and U5114 (N_5114,N_1579,N_609);
xnor U5115 (N_5115,N_1832,N_2875);
or U5116 (N_5116,N_923,N_1940);
nor U5117 (N_5117,N_2724,N_677);
xor U5118 (N_5118,N_82,N_1239);
or U5119 (N_5119,N_898,N_671);
or U5120 (N_5120,N_2492,N_925);
or U5121 (N_5121,N_1120,N_1886);
nor U5122 (N_5122,N_3104,N_1663);
nor U5123 (N_5123,N_2151,N_1104);
or U5124 (N_5124,N_2090,N_1110);
nor U5125 (N_5125,N_1783,N_1170);
nand U5126 (N_5126,N_3111,N_614);
nor U5127 (N_5127,N_1769,N_1975);
xnor U5128 (N_5128,N_236,N_1297);
nand U5129 (N_5129,N_1813,N_1673);
xor U5130 (N_5130,N_998,N_1626);
and U5131 (N_5131,N_1639,N_2684);
nand U5132 (N_5132,N_1250,N_2731);
xnor U5133 (N_5133,N_1878,N_124);
nand U5134 (N_5134,N_43,N_920);
xnor U5135 (N_5135,N_344,N_1960);
nand U5136 (N_5136,N_2599,N_875);
nand U5137 (N_5137,N_2467,N_1075);
nand U5138 (N_5138,N_899,N_685);
nand U5139 (N_5139,N_485,N_768);
nor U5140 (N_5140,N_356,N_714);
nand U5141 (N_5141,N_2460,N_97);
nand U5142 (N_5142,N_1143,N_576);
and U5143 (N_5143,N_1842,N_2816);
nor U5144 (N_5144,N_2529,N_2895);
nor U5145 (N_5145,N_3047,N_2517);
nor U5146 (N_5146,N_2085,N_2668);
and U5147 (N_5147,N_3093,N_1565);
and U5148 (N_5148,N_257,N_1598);
or U5149 (N_5149,N_1762,N_2726);
xnor U5150 (N_5150,N_1078,N_1033);
nor U5151 (N_5151,N_1817,N_634);
or U5152 (N_5152,N_715,N_1046);
and U5153 (N_5153,N_3086,N_2219);
xnor U5154 (N_5154,N_1577,N_115);
nand U5155 (N_5155,N_2091,N_1456);
or U5156 (N_5156,N_2347,N_844);
nor U5157 (N_5157,N_823,N_2088);
or U5158 (N_5158,N_939,N_2049);
or U5159 (N_5159,N_1933,N_2613);
nand U5160 (N_5160,N_2769,N_2020);
and U5161 (N_5161,N_566,N_1286);
nand U5162 (N_5162,N_2613,N_1861);
or U5163 (N_5163,N_132,N_2046);
nor U5164 (N_5164,N_675,N_3028);
xnor U5165 (N_5165,N_198,N_1974);
nor U5166 (N_5166,N_206,N_349);
or U5167 (N_5167,N_1597,N_1135);
or U5168 (N_5168,N_2438,N_2868);
nor U5169 (N_5169,N_2213,N_2211);
and U5170 (N_5170,N_1711,N_1463);
nor U5171 (N_5171,N_877,N_663);
and U5172 (N_5172,N_837,N_2661);
xnor U5173 (N_5173,N_1379,N_2766);
and U5174 (N_5174,N_2774,N_1563);
and U5175 (N_5175,N_2498,N_1652);
xnor U5176 (N_5176,N_2098,N_1148);
and U5177 (N_5177,N_113,N_1160);
nor U5178 (N_5178,N_1133,N_3023);
nand U5179 (N_5179,N_1011,N_852);
xnor U5180 (N_5180,N_1399,N_2087);
and U5181 (N_5181,N_1840,N_2806);
and U5182 (N_5182,N_1060,N_307);
and U5183 (N_5183,N_731,N_525);
or U5184 (N_5184,N_949,N_1247);
or U5185 (N_5185,N_2013,N_2750);
nand U5186 (N_5186,N_2439,N_2456);
nor U5187 (N_5187,N_1974,N_1683);
and U5188 (N_5188,N_2428,N_330);
and U5189 (N_5189,N_1634,N_2216);
nand U5190 (N_5190,N_172,N_2311);
nand U5191 (N_5191,N_1108,N_1861);
nand U5192 (N_5192,N_81,N_957);
and U5193 (N_5193,N_2095,N_2898);
nand U5194 (N_5194,N_1912,N_1380);
and U5195 (N_5195,N_1948,N_2510);
and U5196 (N_5196,N_2258,N_813);
and U5197 (N_5197,N_2860,N_1219);
nor U5198 (N_5198,N_1089,N_2451);
xnor U5199 (N_5199,N_498,N_407);
xnor U5200 (N_5200,N_1852,N_1249);
nand U5201 (N_5201,N_1198,N_843);
and U5202 (N_5202,N_318,N_1300);
nand U5203 (N_5203,N_849,N_1876);
nand U5204 (N_5204,N_819,N_679);
or U5205 (N_5205,N_319,N_2846);
nand U5206 (N_5206,N_1520,N_445);
nor U5207 (N_5207,N_275,N_875);
nor U5208 (N_5208,N_425,N_791);
nor U5209 (N_5209,N_2884,N_801);
and U5210 (N_5210,N_1328,N_788);
nand U5211 (N_5211,N_380,N_196);
nand U5212 (N_5212,N_468,N_2081);
nand U5213 (N_5213,N_34,N_211);
and U5214 (N_5214,N_1527,N_1853);
nand U5215 (N_5215,N_3080,N_1777);
and U5216 (N_5216,N_2211,N_2586);
nand U5217 (N_5217,N_630,N_671);
or U5218 (N_5218,N_2715,N_105);
and U5219 (N_5219,N_1529,N_1984);
xnor U5220 (N_5220,N_1130,N_3022);
and U5221 (N_5221,N_585,N_1788);
nand U5222 (N_5222,N_2637,N_2470);
nand U5223 (N_5223,N_1409,N_195);
and U5224 (N_5224,N_3042,N_630);
nand U5225 (N_5225,N_2421,N_1132);
nor U5226 (N_5226,N_1602,N_2465);
or U5227 (N_5227,N_1490,N_1025);
nor U5228 (N_5228,N_1606,N_1510);
nand U5229 (N_5229,N_844,N_1612);
or U5230 (N_5230,N_2104,N_1772);
and U5231 (N_5231,N_2492,N_416);
and U5232 (N_5232,N_2887,N_2202);
xnor U5233 (N_5233,N_3102,N_1592);
and U5234 (N_5234,N_905,N_789);
or U5235 (N_5235,N_305,N_304);
or U5236 (N_5236,N_1887,N_2569);
nand U5237 (N_5237,N_2630,N_2618);
or U5238 (N_5238,N_1343,N_2845);
or U5239 (N_5239,N_126,N_77);
or U5240 (N_5240,N_526,N_1584);
nand U5241 (N_5241,N_915,N_2476);
and U5242 (N_5242,N_511,N_1157);
nand U5243 (N_5243,N_3073,N_486);
or U5244 (N_5244,N_719,N_1198);
nand U5245 (N_5245,N_1859,N_790);
nand U5246 (N_5246,N_2758,N_2614);
nor U5247 (N_5247,N_2040,N_2850);
nor U5248 (N_5248,N_2540,N_1199);
nand U5249 (N_5249,N_2848,N_2690);
nand U5250 (N_5250,N_2321,N_1366);
nor U5251 (N_5251,N_1794,N_1993);
or U5252 (N_5252,N_414,N_238);
nand U5253 (N_5253,N_603,N_2028);
nor U5254 (N_5254,N_2347,N_2943);
nor U5255 (N_5255,N_3050,N_1936);
and U5256 (N_5256,N_844,N_1247);
nor U5257 (N_5257,N_1329,N_2155);
or U5258 (N_5258,N_882,N_2827);
or U5259 (N_5259,N_660,N_507);
nor U5260 (N_5260,N_1379,N_941);
nor U5261 (N_5261,N_731,N_1035);
nor U5262 (N_5262,N_2442,N_2781);
nand U5263 (N_5263,N_123,N_2461);
and U5264 (N_5264,N_2024,N_2959);
xnor U5265 (N_5265,N_1191,N_2571);
nor U5266 (N_5266,N_3074,N_699);
nand U5267 (N_5267,N_767,N_1155);
nand U5268 (N_5268,N_2504,N_841);
or U5269 (N_5269,N_286,N_117);
nand U5270 (N_5270,N_2668,N_1000);
nor U5271 (N_5271,N_1989,N_1821);
nand U5272 (N_5272,N_2402,N_2012);
nor U5273 (N_5273,N_326,N_3027);
nand U5274 (N_5274,N_118,N_771);
or U5275 (N_5275,N_2921,N_507);
nor U5276 (N_5276,N_633,N_1092);
and U5277 (N_5277,N_1002,N_1079);
nand U5278 (N_5278,N_2856,N_2142);
and U5279 (N_5279,N_1085,N_2961);
nand U5280 (N_5280,N_3122,N_2119);
nor U5281 (N_5281,N_733,N_2666);
and U5282 (N_5282,N_112,N_2915);
nand U5283 (N_5283,N_2835,N_1521);
nor U5284 (N_5284,N_2440,N_1084);
or U5285 (N_5285,N_2825,N_1217);
and U5286 (N_5286,N_1609,N_1978);
nor U5287 (N_5287,N_1786,N_662);
nand U5288 (N_5288,N_143,N_735);
nand U5289 (N_5289,N_1484,N_1518);
xnor U5290 (N_5290,N_206,N_2146);
nand U5291 (N_5291,N_2788,N_1922);
nor U5292 (N_5292,N_686,N_2087);
and U5293 (N_5293,N_2629,N_1511);
and U5294 (N_5294,N_2716,N_2793);
or U5295 (N_5295,N_898,N_40);
nor U5296 (N_5296,N_607,N_1482);
nor U5297 (N_5297,N_122,N_1386);
nor U5298 (N_5298,N_1911,N_1583);
nor U5299 (N_5299,N_2347,N_326);
nand U5300 (N_5300,N_1245,N_3044);
nor U5301 (N_5301,N_2064,N_846);
nor U5302 (N_5302,N_442,N_2901);
or U5303 (N_5303,N_1668,N_2389);
and U5304 (N_5304,N_2422,N_2813);
nand U5305 (N_5305,N_2748,N_1577);
nand U5306 (N_5306,N_2509,N_2048);
nor U5307 (N_5307,N_106,N_868);
xnor U5308 (N_5308,N_509,N_499);
and U5309 (N_5309,N_3009,N_2338);
nand U5310 (N_5310,N_1304,N_2172);
and U5311 (N_5311,N_2850,N_2660);
or U5312 (N_5312,N_1879,N_1973);
xnor U5313 (N_5313,N_6,N_2457);
and U5314 (N_5314,N_281,N_2108);
nor U5315 (N_5315,N_2036,N_2039);
nor U5316 (N_5316,N_1542,N_1437);
nor U5317 (N_5317,N_3105,N_556);
nor U5318 (N_5318,N_2863,N_1856);
or U5319 (N_5319,N_744,N_2544);
nand U5320 (N_5320,N_1677,N_1345);
nor U5321 (N_5321,N_1196,N_2133);
nand U5322 (N_5322,N_1386,N_2778);
nor U5323 (N_5323,N_294,N_821);
nor U5324 (N_5324,N_169,N_218);
or U5325 (N_5325,N_2722,N_1880);
nor U5326 (N_5326,N_761,N_569);
or U5327 (N_5327,N_1194,N_3040);
and U5328 (N_5328,N_2292,N_2136);
nand U5329 (N_5329,N_1491,N_2030);
or U5330 (N_5330,N_130,N_865);
nand U5331 (N_5331,N_980,N_398);
and U5332 (N_5332,N_2603,N_553);
and U5333 (N_5333,N_2874,N_284);
nand U5334 (N_5334,N_539,N_1098);
nand U5335 (N_5335,N_3110,N_2407);
nor U5336 (N_5336,N_1008,N_117);
or U5337 (N_5337,N_1404,N_2952);
nor U5338 (N_5338,N_1439,N_1913);
and U5339 (N_5339,N_1064,N_1112);
xnor U5340 (N_5340,N_1020,N_1159);
and U5341 (N_5341,N_1634,N_46);
xnor U5342 (N_5342,N_3097,N_1527);
nor U5343 (N_5343,N_2798,N_354);
nand U5344 (N_5344,N_649,N_222);
xor U5345 (N_5345,N_2656,N_1429);
nand U5346 (N_5346,N_197,N_2986);
nor U5347 (N_5347,N_2806,N_2403);
nor U5348 (N_5348,N_92,N_2840);
or U5349 (N_5349,N_1209,N_399);
nor U5350 (N_5350,N_3013,N_656);
nor U5351 (N_5351,N_1657,N_1584);
or U5352 (N_5352,N_1077,N_2855);
or U5353 (N_5353,N_1543,N_2835);
nand U5354 (N_5354,N_95,N_2098);
or U5355 (N_5355,N_557,N_2409);
xnor U5356 (N_5356,N_729,N_424);
and U5357 (N_5357,N_1201,N_1536);
nor U5358 (N_5358,N_2272,N_362);
nor U5359 (N_5359,N_556,N_241);
xor U5360 (N_5360,N_2938,N_241);
nor U5361 (N_5361,N_1519,N_405);
and U5362 (N_5362,N_2528,N_2733);
nor U5363 (N_5363,N_1812,N_779);
nor U5364 (N_5364,N_2287,N_1780);
nor U5365 (N_5365,N_1853,N_2490);
nor U5366 (N_5366,N_539,N_424);
xor U5367 (N_5367,N_1905,N_1852);
and U5368 (N_5368,N_1574,N_824);
xor U5369 (N_5369,N_2618,N_1233);
or U5370 (N_5370,N_1770,N_180);
nand U5371 (N_5371,N_42,N_2177);
xor U5372 (N_5372,N_2763,N_1819);
or U5373 (N_5373,N_1967,N_328);
xor U5374 (N_5374,N_1811,N_1058);
nor U5375 (N_5375,N_949,N_2078);
nor U5376 (N_5376,N_1694,N_2005);
and U5377 (N_5377,N_2704,N_2175);
nand U5378 (N_5378,N_2683,N_96);
and U5379 (N_5379,N_2079,N_2435);
nor U5380 (N_5380,N_460,N_712);
nor U5381 (N_5381,N_2162,N_672);
nand U5382 (N_5382,N_1510,N_1626);
and U5383 (N_5383,N_1751,N_2420);
and U5384 (N_5384,N_2985,N_1802);
and U5385 (N_5385,N_250,N_1806);
or U5386 (N_5386,N_2233,N_1360);
and U5387 (N_5387,N_2545,N_424);
or U5388 (N_5388,N_2876,N_2701);
and U5389 (N_5389,N_2860,N_1643);
or U5390 (N_5390,N_1770,N_864);
nor U5391 (N_5391,N_2537,N_2756);
and U5392 (N_5392,N_1057,N_1655);
nand U5393 (N_5393,N_1659,N_2584);
and U5394 (N_5394,N_2714,N_3055);
or U5395 (N_5395,N_1399,N_2633);
or U5396 (N_5396,N_2984,N_2373);
and U5397 (N_5397,N_835,N_242);
nor U5398 (N_5398,N_3072,N_720);
or U5399 (N_5399,N_971,N_179);
or U5400 (N_5400,N_2236,N_800);
nand U5401 (N_5401,N_534,N_2711);
nor U5402 (N_5402,N_1627,N_2807);
or U5403 (N_5403,N_1893,N_1567);
and U5404 (N_5404,N_2928,N_2932);
nor U5405 (N_5405,N_506,N_3102);
xor U5406 (N_5406,N_2428,N_1017);
or U5407 (N_5407,N_1740,N_810);
or U5408 (N_5408,N_2069,N_1022);
and U5409 (N_5409,N_2392,N_1681);
xnor U5410 (N_5410,N_554,N_434);
nand U5411 (N_5411,N_2739,N_2090);
and U5412 (N_5412,N_772,N_13);
and U5413 (N_5413,N_2380,N_622);
nand U5414 (N_5414,N_1662,N_2648);
and U5415 (N_5415,N_1268,N_109);
and U5416 (N_5416,N_1965,N_1106);
nor U5417 (N_5417,N_1171,N_42);
or U5418 (N_5418,N_2371,N_2499);
nand U5419 (N_5419,N_136,N_426);
nand U5420 (N_5420,N_667,N_158);
and U5421 (N_5421,N_1417,N_682);
xnor U5422 (N_5422,N_1489,N_2338);
nor U5423 (N_5423,N_3015,N_532);
or U5424 (N_5424,N_985,N_944);
and U5425 (N_5425,N_3012,N_367);
nor U5426 (N_5426,N_1344,N_231);
or U5427 (N_5427,N_2852,N_566);
or U5428 (N_5428,N_1210,N_1025);
or U5429 (N_5429,N_2314,N_1793);
nor U5430 (N_5430,N_1057,N_3065);
nand U5431 (N_5431,N_857,N_395);
nand U5432 (N_5432,N_1135,N_2716);
nor U5433 (N_5433,N_680,N_2728);
nor U5434 (N_5434,N_3071,N_2524);
nand U5435 (N_5435,N_876,N_2194);
nand U5436 (N_5436,N_1506,N_1002);
and U5437 (N_5437,N_2403,N_1129);
nand U5438 (N_5438,N_706,N_2982);
xnor U5439 (N_5439,N_494,N_940);
nand U5440 (N_5440,N_15,N_1118);
xor U5441 (N_5441,N_1025,N_2132);
and U5442 (N_5442,N_3073,N_1148);
nor U5443 (N_5443,N_1753,N_19);
and U5444 (N_5444,N_721,N_1366);
or U5445 (N_5445,N_980,N_2160);
nand U5446 (N_5446,N_2706,N_879);
or U5447 (N_5447,N_1240,N_573);
nand U5448 (N_5448,N_2351,N_1406);
nand U5449 (N_5449,N_274,N_562);
nand U5450 (N_5450,N_758,N_2759);
or U5451 (N_5451,N_2942,N_1059);
or U5452 (N_5452,N_2544,N_1402);
and U5453 (N_5453,N_660,N_894);
and U5454 (N_5454,N_2010,N_2728);
nor U5455 (N_5455,N_266,N_426);
or U5456 (N_5456,N_2421,N_2273);
and U5457 (N_5457,N_948,N_2203);
or U5458 (N_5458,N_2284,N_3095);
or U5459 (N_5459,N_719,N_2664);
or U5460 (N_5460,N_2951,N_2816);
and U5461 (N_5461,N_82,N_377);
xnor U5462 (N_5462,N_1175,N_2378);
and U5463 (N_5463,N_2396,N_1982);
nand U5464 (N_5464,N_850,N_203);
or U5465 (N_5465,N_2974,N_1981);
or U5466 (N_5466,N_2210,N_2348);
or U5467 (N_5467,N_2675,N_2882);
nand U5468 (N_5468,N_455,N_1938);
nand U5469 (N_5469,N_2132,N_2333);
or U5470 (N_5470,N_3102,N_1108);
or U5471 (N_5471,N_1726,N_593);
nand U5472 (N_5472,N_2321,N_764);
nor U5473 (N_5473,N_2789,N_2824);
or U5474 (N_5474,N_1302,N_2099);
nand U5475 (N_5475,N_2624,N_509);
and U5476 (N_5476,N_1843,N_2953);
nand U5477 (N_5477,N_2022,N_1023);
nor U5478 (N_5478,N_2406,N_2772);
nand U5479 (N_5479,N_2814,N_632);
nand U5480 (N_5480,N_899,N_2759);
and U5481 (N_5481,N_2418,N_1923);
and U5482 (N_5482,N_945,N_2167);
nor U5483 (N_5483,N_239,N_1216);
nor U5484 (N_5484,N_644,N_2536);
nor U5485 (N_5485,N_2036,N_1720);
nor U5486 (N_5486,N_619,N_395);
nand U5487 (N_5487,N_63,N_1436);
and U5488 (N_5488,N_2235,N_2302);
or U5489 (N_5489,N_1284,N_123);
nand U5490 (N_5490,N_719,N_416);
nand U5491 (N_5491,N_2467,N_1380);
or U5492 (N_5492,N_1305,N_1917);
nor U5493 (N_5493,N_806,N_2549);
and U5494 (N_5494,N_2466,N_1292);
and U5495 (N_5495,N_655,N_800);
nor U5496 (N_5496,N_361,N_1086);
nor U5497 (N_5497,N_2236,N_2506);
and U5498 (N_5498,N_156,N_1576);
nand U5499 (N_5499,N_327,N_3006);
or U5500 (N_5500,N_2457,N_906);
nor U5501 (N_5501,N_2923,N_508);
nand U5502 (N_5502,N_927,N_1814);
or U5503 (N_5503,N_1121,N_491);
nor U5504 (N_5504,N_1230,N_2964);
nand U5505 (N_5505,N_579,N_1783);
and U5506 (N_5506,N_1792,N_2194);
and U5507 (N_5507,N_1987,N_649);
and U5508 (N_5508,N_893,N_1265);
nor U5509 (N_5509,N_2103,N_3022);
nor U5510 (N_5510,N_254,N_386);
and U5511 (N_5511,N_610,N_1021);
nor U5512 (N_5512,N_1298,N_566);
and U5513 (N_5513,N_2102,N_669);
or U5514 (N_5514,N_1418,N_3020);
and U5515 (N_5515,N_2825,N_1769);
or U5516 (N_5516,N_2893,N_1871);
nor U5517 (N_5517,N_1937,N_1350);
nand U5518 (N_5518,N_2409,N_2621);
or U5519 (N_5519,N_1624,N_1672);
xor U5520 (N_5520,N_2160,N_921);
and U5521 (N_5521,N_1889,N_3122);
nand U5522 (N_5522,N_1544,N_2433);
nor U5523 (N_5523,N_2247,N_1649);
nand U5524 (N_5524,N_2127,N_3062);
nor U5525 (N_5525,N_1127,N_624);
nor U5526 (N_5526,N_3093,N_635);
and U5527 (N_5527,N_73,N_1744);
nand U5528 (N_5528,N_1188,N_2232);
nor U5529 (N_5529,N_2961,N_1868);
nor U5530 (N_5530,N_609,N_2028);
nand U5531 (N_5531,N_930,N_3103);
or U5532 (N_5532,N_341,N_1121);
and U5533 (N_5533,N_2629,N_2758);
and U5534 (N_5534,N_2743,N_1361);
nor U5535 (N_5535,N_1136,N_2868);
and U5536 (N_5536,N_654,N_2037);
and U5537 (N_5537,N_2837,N_1200);
nand U5538 (N_5538,N_363,N_788);
and U5539 (N_5539,N_939,N_1494);
and U5540 (N_5540,N_1904,N_943);
and U5541 (N_5541,N_794,N_839);
or U5542 (N_5542,N_2310,N_1478);
and U5543 (N_5543,N_2934,N_2958);
or U5544 (N_5544,N_1566,N_2261);
nand U5545 (N_5545,N_2420,N_2099);
or U5546 (N_5546,N_2594,N_54);
nand U5547 (N_5547,N_1989,N_1598);
nor U5548 (N_5548,N_385,N_1549);
xor U5549 (N_5549,N_688,N_625);
nand U5550 (N_5550,N_1269,N_1522);
nor U5551 (N_5551,N_2413,N_2858);
nand U5552 (N_5552,N_2882,N_1471);
or U5553 (N_5553,N_1935,N_1614);
and U5554 (N_5554,N_2452,N_1674);
nor U5555 (N_5555,N_2182,N_11);
and U5556 (N_5556,N_2231,N_2547);
nor U5557 (N_5557,N_2046,N_55);
and U5558 (N_5558,N_540,N_1552);
and U5559 (N_5559,N_2702,N_1543);
and U5560 (N_5560,N_791,N_1169);
and U5561 (N_5561,N_43,N_816);
or U5562 (N_5562,N_785,N_1533);
or U5563 (N_5563,N_243,N_1611);
nor U5564 (N_5564,N_2679,N_2054);
and U5565 (N_5565,N_261,N_767);
nand U5566 (N_5566,N_896,N_193);
or U5567 (N_5567,N_809,N_2426);
or U5568 (N_5568,N_2133,N_846);
and U5569 (N_5569,N_1684,N_829);
nor U5570 (N_5570,N_493,N_822);
nand U5571 (N_5571,N_2947,N_1051);
xnor U5572 (N_5572,N_3078,N_2852);
or U5573 (N_5573,N_2867,N_793);
nor U5574 (N_5574,N_3016,N_1096);
nand U5575 (N_5575,N_412,N_577);
and U5576 (N_5576,N_2792,N_1792);
and U5577 (N_5577,N_1234,N_3020);
nand U5578 (N_5578,N_2794,N_2777);
xor U5579 (N_5579,N_1196,N_1800);
and U5580 (N_5580,N_1963,N_2024);
and U5581 (N_5581,N_2623,N_722);
nor U5582 (N_5582,N_2948,N_2666);
and U5583 (N_5583,N_2820,N_1394);
xor U5584 (N_5584,N_1775,N_1956);
and U5585 (N_5585,N_1983,N_2664);
and U5586 (N_5586,N_2883,N_3071);
and U5587 (N_5587,N_2315,N_2750);
and U5588 (N_5588,N_1310,N_1614);
nand U5589 (N_5589,N_59,N_1935);
nor U5590 (N_5590,N_1523,N_1609);
nand U5591 (N_5591,N_3056,N_19);
or U5592 (N_5592,N_1851,N_2551);
nor U5593 (N_5593,N_1793,N_1535);
nand U5594 (N_5594,N_845,N_1828);
nor U5595 (N_5595,N_1378,N_1477);
or U5596 (N_5596,N_3077,N_933);
and U5597 (N_5597,N_935,N_568);
or U5598 (N_5598,N_3033,N_2355);
nand U5599 (N_5599,N_1373,N_1803);
nor U5600 (N_5600,N_1431,N_2888);
and U5601 (N_5601,N_23,N_2062);
or U5602 (N_5602,N_1496,N_1602);
or U5603 (N_5603,N_1454,N_1780);
and U5604 (N_5604,N_2709,N_708);
or U5605 (N_5605,N_1273,N_3094);
nor U5606 (N_5606,N_263,N_380);
or U5607 (N_5607,N_616,N_2004);
or U5608 (N_5608,N_728,N_2094);
and U5609 (N_5609,N_1270,N_66);
or U5610 (N_5610,N_43,N_1035);
or U5611 (N_5611,N_126,N_2667);
and U5612 (N_5612,N_1874,N_1706);
nand U5613 (N_5613,N_24,N_2670);
and U5614 (N_5614,N_2757,N_187);
xnor U5615 (N_5615,N_2612,N_818);
or U5616 (N_5616,N_1486,N_905);
xnor U5617 (N_5617,N_1004,N_597);
and U5618 (N_5618,N_3068,N_2485);
xnor U5619 (N_5619,N_734,N_1185);
nor U5620 (N_5620,N_1736,N_2205);
and U5621 (N_5621,N_1510,N_98);
and U5622 (N_5622,N_38,N_495);
or U5623 (N_5623,N_1515,N_828);
and U5624 (N_5624,N_2886,N_1038);
xor U5625 (N_5625,N_2889,N_1244);
and U5626 (N_5626,N_926,N_1660);
nor U5627 (N_5627,N_553,N_2905);
and U5628 (N_5628,N_396,N_1811);
xnor U5629 (N_5629,N_110,N_2191);
and U5630 (N_5630,N_2626,N_2809);
xor U5631 (N_5631,N_198,N_1700);
nand U5632 (N_5632,N_1084,N_1676);
xor U5633 (N_5633,N_1115,N_182);
or U5634 (N_5634,N_1790,N_768);
and U5635 (N_5635,N_1399,N_2071);
nand U5636 (N_5636,N_2091,N_1636);
nor U5637 (N_5637,N_685,N_710);
nand U5638 (N_5638,N_2982,N_1441);
xnor U5639 (N_5639,N_1097,N_2223);
nand U5640 (N_5640,N_974,N_1468);
and U5641 (N_5641,N_693,N_3101);
nor U5642 (N_5642,N_2572,N_2192);
and U5643 (N_5643,N_3122,N_2637);
nand U5644 (N_5644,N_784,N_197);
and U5645 (N_5645,N_1207,N_2272);
or U5646 (N_5646,N_1365,N_2616);
nor U5647 (N_5647,N_1830,N_3086);
and U5648 (N_5648,N_2561,N_2510);
nand U5649 (N_5649,N_230,N_476);
and U5650 (N_5650,N_2704,N_2013);
nand U5651 (N_5651,N_3065,N_2478);
or U5652 (N_5652,N_1403,N_2187);
and U5653 (N_5653,N_1938,N_202);
nor U5654 (N_5654,N_2080,N_436);
nor U5655 (N_5655,N_1297,N_1328);
nor U5656 (N_5656,N_2444,N_658);
nand U5657 (N_5657,N_2395,N_2931);
xnor U5658 (N_5658,N_2444,N_1607);
xnor U5659 (N_5659,N_2491,N_1134);
or U5660 (N_5660,N_1987,N_2621);
or U5661 (N_5661,N_3042,N_1095);
nor U5662 (N_5662,N_532,N_2583);
nand U5663 (N_5663,N_2531,N_351);
or U5664 (N_5664,N_656,N_1757);
nand U5665 (N_5665,N_964,N_1715);
and U5666 (N_5666,N_1010,N_2401);
or U5667 (N_5667,N_1368,N_3051);
nand U5668 (N_5668,N_1646,N_2229);
nand U5669 (N_5669,N_573,N_1701);
and U5670 (N_5670,N_2038,N_2490);
nand U5671 (N_5671,N_1444,N_1745);
and U5672 (N_5672,N_1762,N_1169);
and U5673 (N_5673,N_2777,N_1783);
or U5674 (N_5674,N_1691,N_128);
or U5675 (N_5675,N_3042,N_2759);
and U5676 (N_5676,N_925,N_2523);
xnor U5677 (N_5677,N_2191,N_2999);
xnor U5678 (N_5678,N_3,N_2744);
and U5679 (N_5679,N_566,N_1956);
nor U5680 (N_5680,N_1518,N_2175);
and U5681 (N_5681,N_677,N_1221);
nand U5682 (N_5682,N_3071,N_106);
and U5683 (N_5683,N_1616,N_2266);
nor U5684 (N_5684,N_2758,N_173);
and U5685 (N_5685,N_2578,N_1272);
nand U5686 (N_5686,N_2192,N_1731);
and U5687 (N_5687,N_1769,N_1758);
nand U5688 (N_5688,N_1889,N_2044);
nand U5689 (N_5689,N_2745,N_973);
or U5690 (N_5690,N_2829,N_2212);
nand U5691 (N_5691,N_619,N_2514);
or U5692 (N_5692,N_2338,N_2070);
or U5693 (N_5693,N_3104,N_1831);
and U5694 (N_5694,N_1347,N_1579);
or U5695 (N_5695,N_1341,N_1105);
and U5696 (N_5696,N_2362,N_2822);
or U5697 (N_5697,N_900,N_986);
nand U5698 (N_5698,N_1747,N_1062);
nor U5699 (N_5699,N_1977,N_549);
nor U5700 (N_5700,N_588,N_1272);
nand U5701 (N_5701,N_701,N_387);
nand U5702 (N_5702,N_2418,N_517);
or U5703 (N_5703,N_2752,N_2397);
and U5704 (N_5704,N_1524,N_757);
or U5705 (N_5705,N_27,N_2541);
or U5706 (N_5706,N_1818,N_1648);
and U5707 (N_5707,N_1009,N_1975);
nand U5708 (N_5708,N_2916,N_1663);
xnor U5709 (N_5709,N_2504,N_3061);
and U5710 (N_5710,N_566,N_2184);
nor U5711 (N_5711,N_423,N_1903);
nand U5712 (N_5712,N_1437,N_2794);
or U5713 (N_5713,N_2265,N_319);
nand U5714 (N_5714,N_2349,N_2088);
and U5715 (N_5715,N_2682,N_275);
nor U5716 (N_5716,N_2637,N_1238);
and U5717 (N_5717,N_2683,N_1328);
xnor U5718 (N_5718,N_1795,N_1165);
and U5719 (N_5719,N_171,N_155);
nand U5720 (N_5720,N_2813,N_2853);
and U5721 (N_5721,N_3100,N_3038);
and U5722 (N_5722,N_1103,N_139);
nor U5723 (N_5723,N_2556,N_1710);
and U5724 (N_5724,N_2416,N_188);
xnor U5725 (N_5725,N_2153,N_838);
nor U5726 (N_5726,N_534,N_1324);
and U5727 (N_5727,N_2837,N_1408);
nor U5728 (N_5728,N_2179,N_1620);
or U5729 (N_5729,N_1990,N_1949);
xor U5730 (N_5730,N_1950,N_633);
and U5731 (N_5731,N_1646,N_957);
nand U5732 (N_5732,N_255,N_1708);
or U5733 (N_5733,N_2701,N_2539);
nand U5734 (N_5734,N_619,N_1045);
and U5735 (N_5735,N_1874,N_1144);
or U5736 (N_5736,N_3111,N_805);
nand U5737 (N_5737,N_2956,N_687);
nand U5738 (N_5738,N_1250,N_2861);
nand U5739 (N_5739,N_795,N_372);
nor U5740 (N_5740,N_1721,N_375);
xnor U5741 (N_5741,N_17,N_1186);
and U5742 (N_5742,N_122,N_445);
xor U5743 (N_5743,N_814,N_2736);
nor U5744 (N_5744,N_471,N_1600);
nand U5745 (N_5745,N_2400,N_1438);
and U5746 (N_5746,N_234,N_1616);
and U5747 (N_5747,N_787,N_2591);
nand U5748 (N_5748,N_867,N_786);
or U5749 (N_5749,N_1786,N_1371);
or U5750 (N_5750,N_2793,N_2355);
nand U5751 (N_5751,N_2817,N_1201);
xnor U5752 (N_5752,N_2152,N_2509);
nor U5753 (N_5753,N_332,N_2390);
nor U5754 (N_5754,N_1330,N_640);
nor U5755 (N_5755,N_1820,N_1484);
nor U5756 (N_5756,N_2557,N_2250);
or U5757 (N_5757,N_3124,N_41);
nand U5758 (N_5758,N_2754,N_1208);
nor U5759 (N_5759,N_1852,N_2560);
nor U5760 (N_5760,N_542,N_943);
or U5761 (N_5761,N_1626,N_910);
nand U5762 (N_5762,N_1527,N_1982);
nor U5763 (N_5763,N_621,N_530);
and U5764 (N_5764,N_2803,N_698);
and U5765 (N_5765,N_419,N_383);
and U5766 (N_5766,N_2603,N_2463);
nor U5767 (N_5767,N_3029,N_2251);
xor U5768 (N_5768,N_2523,N_583);
or U5769 (N_5769,N_1112,N_354);
or U5770 (N_5770,N_2521,N_2279);
nor U5771 (N_5771,N_1590,N_1789);
nor U5772 (N_5772,N_1397,N_1248);
nor U5773 (N_5773,N_2989,N_1269);
or U5774 (N_5774,N_1111,N_1191);
nor U5775 (N_5775,N_2044,N_1445);
nand U5776 (N_5776,N_3010,N_1597);
nor U5777 (N_5777,N_1766,N_1220);
and U5778 (N_5778,N_3091,N_344);
and U5779 (N_5779,N_1065,N_1401);
nor U5780 (N_5780,N_1551,N_2926);
and U5781 (N_5781,N_1418,N_1214);
or U5782 (N_5782,N_2712,N_2331);
and U5783 (N_5783,N_634,N_1337);
nor U5784 (N_5784,N_3120,N_546);
nor U5785 (N_5785,N_2113,N_1885);
or U5786 (N_5786,N_3091,N_1368);
nor U5787 (N_5787,N_2437,N_907);
nand U5788 (N_5788,N_1403,N_2883);
and U5789 (N_5789,N_2963,N_2124);
or U5790 (N_5790,N_2615,N_1338);
nor U5791 (N_5791,N_3001,N_1726);
or U5792 (N_5792,N_889,N_1859);
nand U5793 (N_5793,N_1095,N_152);
or U5794 (N_5794,N_2677,N_1597);
nand U5795 (N_5795,N_2178,N_1895);
xnor U5796 (N_5796,N_1585,N_1881);
and U5797 (N_5797,N_1311,N_471);
nand U5798 (N_5798,N_1041,N_1033);
nand U5799 (N_5799,N_2650,N_2955);
xor U5800 (N_5800,N_1574,N_1870);
nor U5801 (N_5801,N_1466,N_1346);
and U5802 (N_5802,N_188,N_2725);
nor U5803 (N_5803,N_683,N_939);
nor U5804 (N_5804,N_1293,N_1209);
xnor U5805 (N_5805,N_2351,N_321);
or U5806 (N_5806,N_823,N_3025);
or U5807 (N_5807,N_2677,N_1967);
or U5808 (N_5808,N_774,N_118);
nor U5809 (N_5809,N_2428,N_233);
and U5810 (N_5810,N_1500,N_234);
nor U5811 (N_5811,N_992,N_377);
xor U5812 (N_5812,N_2897,N_20);
and U5813 (N_5813,N_1507,N_1891);
nand U5814 (N_5814,N_2311,N_2444);
nand U5815 (N_5815,N_2293,N_1412);
or U5816 (N_5816,N_297,N_910);
xnor U5817 (N_5817,N_386,N_111);
and U5818 (N_5818,N_2459,N_2215);
nor U5819 (N_5819,N_2171,N_117);
nor U5820 (N_5820,N_986,N_539);
or U5821 (N_5821,N_1951,N_452);
nand U5822 (N_5822,N_537,N_2781);
nand U5823 (N_5823,N_1458,N_2362);
nand U5824 (N_5824,N_2195,N_2986);
or U5825 (N_5825,N_37,N_125);
and U5826 (N_5826,N_203,N_1011);
nand U5827 (N_5827,N_2871,N_2121);
nand U5828 (N_5828,N_2827,N_711);
or U5829 (N_5829,N_969,N_2100);
xnor U5830 (N_5830,N_2162,N_2946);
nand U5831 (N_5831,N_527,N_284);
nand U5832 (N_5832,N_2891,N_3045);
or U5833 (N_5833,N_1076,N_2171);
or U5834 (N_5834,N_1643,N_676);
nand U5835 (N_5835,N_1494,N_1252);
and U5836 (N_5836,N_2881,N_232);
or U5837 (N_5837,N_37,N_47);
nor U5838 (N_5838,N_910,N_2654);
or U5839 (N_5839,N_2785,N_497);
xnor U5840 (N_5840,N_1086,N_3029);
and U5841 (N_5841,N_259,N_675);
nand U5842 (N_5842,N_2885,N_2527);
xnor U5843 (N_5843,N_1973,N_359);
and U5844 (N_5844,N_1600,N_1584);
and U5845 (N_5845,N_782,N_1712);
and U5846 (N_5846,N_2388,N_2662);
nor U5847 (N_5847,N_2784,N_455);
nor U5848 (N_5848,N_1684,N_1986);
or U5849 (N_5849,N_939,N_133);
nor U5850 (N_5850,N_458,N_2689);
or U5851 (N_5851,N_597,N_2879);
or U5852 (N_5852,N_2938,N_2291);
nor U5853 (N_5853,N_841,N_2892);
and U5854 (N_5854,N_2816,N_2521);
and U5855 (N_5855,N_2840,N_2971);
nand U5856 (N_5856,N_2055,N_2919);
nand U5857 (N_5857,N_909,N_2078);
and U5858 (N_5858,N_1259,N_810);
or U5859 (N_5859,N_2207,N_961);
or U5860 (N_5860,N_2443,N_254);
and U5861 (N_5861,N_48,N_1629);
and U5862 (N_5862,N_2426,N_900);
nand U5863 (N_5863,N_1655,N_3105);
and U5864 (N_5864,N_327,N_2746);
and U5865 (N_5865,N_2024,N_2277);
and U5866 (N_5866,N_2483,N_362);
xor U5867 (N_5867,N_1738,N_2330);
nand U5868 (N_5868,N_2022,N_260);
and U5869 (N_5869,N_2688,N_1107);
nand U5870 (N_5870,N_1065,N_137);
nor U5871 (N_5871,N_472,N_536);
nand U5872 (N_5872,N_2787,N_1083);
nor U5873 (N_5873,N_854,N_485);
nand U5874 (N_5874,N_240,N_2141);
and U5875 (N_5875,N_1111,N_876);
nand U5876 (N_5876,N_2384,N_42);
nand U5877 (N_5877,N_1032,N_2286);
and U5878 (N_5878,N_839,N_1112);
xnor U5879 (N_5879,N_1306,N_2883);
and U5880 (N_5880,N_2878,N_1894);
or U5881 (N_5881,N_2361,N_2503);
and U5882 (N_5882,N_322,N_132);
nor U5883 (N_5883,N_1547,N_1277);
nand U5884 (N_5884,N_1835,N_2866);
nor U5885 (N_5885,N_95,N_307);
nand U5886 (N_5886,N_2887,N_2284);
or U5887 (N_5887,N_1351,N_808);
or U5888 (N_5888,N_1964,N_1784);
nor U5889 (N_5889,N_1845,N_1768);
or U5890 (N_5890,N_1552,N_1166);
nor U5891 (N_5891,N_2440,N_1671);
or U5892 (N_5892,N_310,N_105);
nand U5893 (N_5893,N_3092,N_1956);
nand U5894 (N_5894,N_123,N_821);
nor U5895 (N_5895,N_1740,N_451);
xnor U5896 (N_5896,N_823,N_1306);
or U5897 (N_5897,N_1728,N_1110);
xnor U5898 (N_5898,N_3072,N_194);
nor U5899 (N_5899,N_823,N_1767);
and U5900 (N_5900,N_3091,N_2573);
and U5901 (N_5901,N_240,N_2672);
or U5902 (N_5902,N_2452,N_1988);
nand U5903 (N_5903,N_1592,N_2860);
nand U5904 (N_5904,N_1796,N_18);
nor U5905 (N_5905,N_2440,N_2150);
nand U5906 (N_5906,N_1807,N_1615);
xor U5907 (N_5907,N_1165,N_2503);
nor U5908 (N_5908,N_2540,N_578);
nor U5909 (N_5909,N_2628,N_1517);
nand U5910 (N_5910,N_1556,N_1774);
xnor U5911 (N_5911,N_2626,N_1145);
nor U5912 (N_5912,N_1448,N_136);
or U5913 (N_5913,N_1837,N_2213);
or U5914 (N_5914,N_2660,N_333);
and U5915 (N_5915,N_2293,N_1052);
nor U5916 (N_5916,N_729,N_835);
xnor U5917 (N_5917,N_2675,N_2732);
nor U5918 (N_5918,N_2683,N_1820);
nand U5919 (N_5919,N_2171,N_2221);
and U5920 (N_5920,N_2711,N_1104);
nor U5921 (N_5921,N_579,N_483);
nand U5922 (N_5922,N_336,N_542);
nor U5923 (N_5923,N_1360,N_2325);
or U5924 (N_5924,N_1082,N_2710);
and U5925 (N_5925,N_504,N_2362);
nand U5926 (N_5926,N_1380,N_1152);
and U5927 (N_5927,N_1886,N_2369);
or U5928 (N_5928,N_655,N_2467);
nand U5929 (N_5929,N_1977,N_909);
xor U5930 (N_5930,N_2881,N_2423);
xnor U5931 (N_5931,N_1201,N_1021);
or U5932 (N_5932,N_196,N_2716);
nand U5933 (N_5933,N_930,N_2224);
nand U5934 (N_5934,N_1888,N_818);
or U5935 (N_5935,N_2896,N_1638);
nand U5936 (N_5936,N_1123,N_419);
or U5937 (N_5937,N_714,N_1709);
and U5938 (N_5938,N_1927,N_2772);
nand U5939 (N_5939,N_786,N_2884);
or U5940 (N_5940,N_502,N_2245);
nor U5941 (N_5941,N_2231,N_2517);
and U5942 (N_5942,N_102,N_2198);
nor U5943 (N_5943,N_617,N_1329);
or U5944 (N_5944,N_1759,N_321);
or U5945 (N_5945,N_603,N_1287);
or U5946 (N_5946,N_2692,N_2760);
nor U5947 (N_5947,N_1207,N_2253);
and U5948 (N_5948,N_180,N_1279);
and U5949 (N_5949,N_2940,N_2633);
nand U5950 (N_5950,N_1531,N_718);
nand U5951 (N_5951,N_2158,N_1091);
nor U5952 (N_5952,N_994,N_2194);
and U5953 (N_5953,N_2407,N_1608);
or U5954 (N_5954,N_619,N_887);
nand U5955 (N_5955,N_2246,N_2874);
nand U5956 (N_5956,N_922,N_1249);
nand U5957 (N_5957,N_347,N_2078);
or U5958 (N_5958,N_1304,N_2803);
nor U5959 (N_5959,N_874,N_290);
nor U5960 (N_5960,N_2272,N_1216);
nor U5961 (N_5961,N_2086,N_2429);
and U5962 (N_5962,N_440,N_2985);
nor U5963 (N_5963,N_2784,N_1576);
nor U5964 (N_5964,N_3106,N_2663);
nand U5965 (N_5965,N_257,N_744);
xnor U5966 (N_5966,N_3029,N_1649);
nor U5967 (N_5967,N_1664,N_2572);
nor U5968 (N_5968,N_1314,N_2882);
nand U5969 (N_5969,N_523,N_2153);
and U5970 (N_5970,N_1533,N_250);
nand U5971 (N_5971,N_805,N_2690);
xor U5972 (N_5972,N_1484,N_3063);
and U5973 (N_5973,N_1004,N_2870);
xor U5974 (N_5974,N_1992,N_2276);
and U5975 (N_5975,N_1309,N_2730);
nor U5976 (N_5976,N_594,N_779);
and U5977 (N_5977,N_3064,N_802);
and U5978 (N_5978,N_1265,N_2205);
and U5979 (N_5979,N_697,N_2729);
nor U5980 (N_5980,N_2364,N_875);
xnor U5981 (N_5981,N_208,N_231);
or U5982 (N_5982,N_174,N_1293);
and U5983 (N_5983,N_278,N_1522);
or U5984 (N_5984,N_371,N_1593);
and U5985 (N_5985,N_2273,N_1563);
or U5986 (N_5986,N_1525,N_2805);
nand U5987 (N_5987,N_1170,N_947);
or U5988 (N_5988,N_2409,N_1612);
or U5989 (N_5989,N_225,N_2604);
nor U5990 (N_5990,N_79,N_2388);
and U5991 (N_5991,N_41,N_1026);
and U5992 (N_5992,N_821,N_2843);
and U5993 (N_5993,N_1148,N_2515);
and U5994 (N_5994,N_605,N_1616);
nor U5995 (N_5995,N_2291,N_755);
nor U5996 (N_5996,N_1282,N_52);
or U5997 (N_5997,N_1500,N_439);
or U5998 (N_5998,N_917,N_2228);
nand U5999 (N_5999,N_1890,N_35);
and U6000 (N_6000,N_950,N_2451);
or U6001 (N_6001,N_1820,N_2235);
and U6002 (N_6002,N_2926,N_1905);
nand U6003 (N_6003,N_1677,N_2210);
and U6004 (N_6004,N_617,N_1305);
nor U6005 (N_6005,N_2557,N_2072);
nand U6006 (N_6006,N_1785,N_1009);
nor U6007 (N_6007,N_628,N_135);
or U6008 (N_6008,N_1420,N_429);
nand U6009 (N_6009,N_1277,N_177);
or U6010 (N_6010,N_2675,N_971);
or U6011 (N_6011,N_2290,N_518);
xor U6012 (N_6012,N_334,N_2987);
or U6013 (N_6013,N_1802,N_3079);
nand U6014 (N_6014,N_1944,N_2488);
or U6015 (N_6015,N_209,N_1763);
or U6016 (N_6016,N_818,N_1788);
nor U6017 (N_6017,N_2414,N_1743);
nor U6018 (N_6018,N_1938,N_969);
or U6019 (N_6019,N_1250,N_1148);
or U6020 (N_6020,N_1078,N_1810);
or U6021 (N_6021,N_1918,N_3117);
nand U6022 (N_6022,N_365,N_770);
nor U6023 (N_6023,N_2771,N_749);
and U6024 (N_6024,N_3024,N_1169);
and U6025 (N_6025,N_2505,N_2757);
or U6026 (N_6026,N_2175,N_2248);
nand U6027 (N_6027,N_2279,N_2297);
nor U6028 (N_6028,N_1559,N_80);
or U6029 (N_6029,N_3035,N_2582);
or U6030 (N_6030,N_98,N_1413);
nand U6031 (N_6031,N_211,N_679);
and U6032 (N_6032,N_879,N_1168);
nor U6033 (N_6033,N_2543,N_2002);
and U6034 (N_6034,N_115,N_2287);
and U6035 (N_6035,N_2700,N_1763);
nand U6036 (N_6036,N_1990,N_1134);
or U6037 (N_6037,N_638,N_1642);
or U6038 (N_6038,N_2851,N_2995);
nor U6039 (N_6039,N_1936,N_2068);
and U6040 (N_6040,N_148,N_772);
nor U6041 (N_6041,N_279,N_819);
or U6042 (N_6042,N_1938,N_973);
xor U6043 (N_6043,N_231,N_1288);
or U6044 (N_6044,N_1952,N_113);
xor U6045 (N_6045,N_812,N_1966);
or U6046 (N_6046,N_368,N_913);
or U6047 (N_6047,N_1235,N_86);
nand U6048 (N_6048,N_676,N_2069);
nor U6049 (N_6049,N_2442,N_919);
or U6050 (N_6050,N_2384,N_2037);
or U6051 (N_6051,N_2500,N_1323);
or U6052 (N_6052,N_1407,N_1532);
and U6053 (N_6053,N_1569,N_2261);
nor U6054 (N_6054,N_2326,N_2395);
or U6055 (N_6055,N_413,N_1503);
or U6056 (N_6056,N_939,N_2047);
nor U6057 (N_6057,N_735,N_421);
nand U6058 (N_6058,N_2871,N_521);
and U6059 (N_6059,N_295,N_769);
and U6060 (N_6060,N_445,N_2576);
and U6061 (N_6061,N_825,N_2678);
or U6062 (N_6062,N_1948,N_2452);
xnor U6063 (N_6063,N_2363,N_1858);
nor U6064 (N_6064,N_1962,N_838);
and U6065 (N_6065,N_810,N_63);
nand U6066 (N_6066,N_2376,N_1274);
or U6067 (N_6067,N_514,N_361);
nor U6068 (N_6068,N_1953,N_127);
nand U6069 (N_6069,N_1445,N_470);
nand U6070 (N_6070,N_941,N_363);
or U6071 (N_6071,N_1608,N_1235);
nor U6072 (N_6072,N_1717,N_2463);
or U6073 (N_6073,N_1076,N_3077);
xnor U6074 (N_6074,N_1031,N_1566);
and U6075 (N_6075,N_2618,N_188);
or U6076 (N_6076,N_1644,N_2660);
nand U6077 (N_6077,N_115,N_2976);
nor U6078 (N_6078,N_296,N_2146);
xor U6079 (N_6079,N_2488,N_2803);
nor U6080 (N_6080,N_2669,N_2350);
nor U6081 (N_6081,N_1992,N_2340);
xnor U6082 (N_6082,N_2741,N_590);
nor U6083 (N_6083,N_1600,N_2862);
xor U6084 (N_6084,N_1238,N_690);
nand U6085 (N_6085,N_46,N_1644);
nor U6086 (N_6086,N_2511,N_2901);
nand U6087 (N_6087,N_2747,N_2425);
nor U6088 (N_6088,N_1994,N_123);
nor U6089 (N_6089,N_2223,N_1732);
and U6090 (N_6090,N_2993,N_2315);
nand U6091 (N_6091,N_1642,N_528);
nor U6092 (N_6092,N_459,N_2049);
nor U6093 (N_6093,N_1825,N_775);
or U6094 (N_6094,N_883,N_504);
and U6095 (N_6095,N_347,N_539);
nor U6096 (N_6096,N_1603,N_2061);
and U6097 (N_6097,N_906,N_2727);
nor U6098 (N_6098,N_1699,N_216);
nand U6099 (N_6099,N_2656,N_2608);
and U6100 (N_6100,N_2167,N_263);
nand U6101 (N_6101,N_1443,N_596);
and U6102 (N_6102,N_416,N_3044);
nor U6103 (N_6103,N_830,N_1933);
or U6104 (N_6104,N_2920,N_1839);
and U6105 (N_6105,N_1536,N_1231);
and U6106 (N_6106,N_2761,N_1782);
nor U6107 (N_6107,N_1147,N_2105);
xor U6108 (N_6108,N_3011,N_807);
nor U6109 (N_6109,N_639,N_591);
or U6110 (N_6110,N_2464,N_1232);
nor U6111 (N_6111,N_838,N_2106);
or U6112 (N_6112,N_789,N_421);
or U6113 (N_6113,N_3052,N_1364);
and U6114 (N_6114,N_1385,N_886);
nand U6115 (N_6115,N_2751,N_3063);
xnor U6116 (N_6116,N_314,N_50);
xnor U6117 (N_6117,N_2753,N_499);
nand U6118 (N_6118,N_127,N_2553);
or U6119 (N_6119,N_1022,N_2746);
xnor U6120 (N_6120,N_1354,N_980);
nor U6121 (N_6121,N_1735,N_2117);
and U6122 (N_6122,N_3110,N_923);
nor U6123 (N_6123,N_1408,N_2045);
nand U6124 (N_6124,N_1178,N_1300);
and U6125 (N_6125,N_2526,N_153);
nor U6126 (N_6126,N_1318,N_2865);
xnor U6127 (N_6127,N_2197,N_648);
and U6128 (N_6128,N_254,N_718);
or U6129 (N_6129,N_322,N_462);
and U6130 (N_6130,N_1594,N_1456);
or U6131 (N_6131,N_8,N_1707);
and U6132 (N_6132,N_2382,N_1333);
and U6133 (N_6133,N_2849,N_344);
nand U6134 (N_6134,N_2897,N_668);
nand U6135 (N_6135,N_669,N_147);
nand U6136 (N_6136,N_362,N_315);
nand U6137 (N_6137,N_2518,N_3013);
nand U6138 (N_6138,N_254,N_2714);
and U6139 (N_6139,N_2407,N_2538);
nand U6140 (N_6140,N_189,N_379);
xnor U6141 (N_6141,N_168,N_7);
xor U6142 (N_6142,N_945,N_412);
nor U6143 (N_6143,N_1482,N_806);
nand U6144 (N_6144,N_1164,N_2133);
and U6145 (N_6145,N_2317,N_1335);
xnor U6146 (N_6146,N_1905,N_1880);
nand U6147 (N_6147,N_2011,N_2092);
and U6148 (N_6148,N_1433,N_869);
nand U6149 (N_6149,N_856,N_299);
nand U6150 (N_6150,N_627,N_1766);
and U6151 (N_6151,N_214,N_527);
and U6152 (N_6152,N_2464,N_208);
nand U6153 (N_6153,N_3010,N_153);
xnor U6154 (N_6154,N_323,N_1591);
nand U6155 (N_6155,N_2623,N_3110);
and U6156 (N_6156,N_1427,N_2795);
or U6157 (N_6157,N_2238,N_2367);
nor U6158 (N_6158,N_2308,N_2076);
xor U6159 (N_6159,N_1973,N_704);
nor U6160 (N_6160,N_1038,N_1254);
or U6161 (N_6161,N_1295,N_2691);
nor U6162 (N_6162,N_177,N_485);
nand U6163 (N_6163,N_2626,N_328);
and U6164 (N_6164,N_1281,N_727);
or U6165 (N_6165,N_1614,N_1861);
nor U6166 (N_6166,N_1220,N_1363);
nor U6167 (N_6167,N_2483,N_1699);
or U6168 (N_6168,N_175,N_2285);
nor U6169 (N_6169,N_602,N_157);
and U6170 (N_6170,N_1062,N_1215);
nand U6171 (N_6171,N_1378,N_1747);
and U6172 (N_6172,N_2960,N_1505);
nand U6173 (N_6173,N_142,N_251);
nand U6174 (N_6174,N_2354,N_1685);
nor U6175 (N_6175,N_410,N_3064);
nor U6176 (N_6176,N_2565,N_270);
nand U6177 (N_6177,N_3112,N_3036);
nor U6178 (N_6178,N_409,N_1659);
xor U6179 (N_6179,N_1498,N_2322);
nand U6180 (N_6180,N_389,N_1760);
xnor U6181 (N_6181,N_1168,N_2756);
nand U6182 (N_6182,N_250,N_716);
and U6183 (N_6183,N_1063,N_1391);
nor U6184 (N_6184,N_1115,N_1091);
nor U6185 (N_6185,N_724,N_165);
nand U6186 (N_6186,N_2641,N_2166);
nand U6187 (N_6187,N_590,N_1566);
nand U6188 (N_6188,N_2190,N_28);
or U6189 (N_6189,N_1981,N_2139);
or U6190 (N_6190,N_1571,N_1343);
nand U6191 (N_6191,N_2520,N_1690);
and U6192 (N_6192,N_1487,N_2062);
or U6193 (N_6193,N_1997,N_631);
nand U6194 (N_6194,N_1684,N_1483);
nand U6195 (N_6195,N_1671,N_2725);
or U6196 (N_6196,N_2714,N_853);
or U6197 (N_6197,N_1414,N_1205);
and U6198 (N_6198,N_2285,N_438);
nor U6199 (N_6199,N_2849,N_1891);
or U6200 (N_6200,N_2606,N_439);
or U6201 (N_6201,N_1851,N_774);
nor U6202 (N_6202,N_119,N_2470);
and U6203 (N_6203,N_1217,N_2252);
or U6204 (N_6204,N_1692,N_1784);
or U6205 (N_6205,N_1903,N_1423);
or U6206 (N_6206,N_2050,N_2653);
nand U6207 (N_6207,N_2873,N_160);
and U6208 (N_6208,N_72,N_1482);
nor U6209 (N_6209,N_2717,N_503);
and U6210 (N_6210,N_668,N_525);
xnor U6211 (N_6211,N_2805,N_2771);
nor U6212 (N_6212,N_2873,N_1347);
nor U6213 (N_6213,N_2027,N_2070);
nor U6214 (N_6214,N_2761,N_608);
xor U6215 (N_6215,N_1623,N_2922);
and U6216 (N_6216,N_245,N_128);
nor U6217 (N_6217,N_720,N_2393);
nor U6218 (N_6218,N_2779,N_2802);
or U6219 (N_6219,N_898,N_1901);
nand U6220 (N_6220,N_791,N_323);
or U6221 (N_6221,N_1395,N_2746);
and U6222 (N_6222,N_1498,N_1659);
nor U6223 (N_6223,N_1017,N_2720);
and U6224 (N_6224,N_1292,N_424);
or U6225 (N_6225,N_2685,N_86);
or U6226 (N_6226,N_1927,N_415);
or U6227 (N_6227,N_587,N_364);
or U6228 (N_6228,N_2363,N_1370);
and U6229 (N_6229,N_1770,N_2818);
or U6230 (N_6230,N_671,N_1903);
nand U6231 (N_6231,N_1357,N_1158);
and U6232 (N_6232,N_2441,N_1084);
and U6233 (N_6233,N_2520,N_361);
nand U6234 (N_6234,N_1524,N_884);
nand U6235 (N_6235,N_1508,N_2328);
nor U6236 (N_6236,N_2104,N_2691);
or U6237 (N_6237,N_3115,N_247);
nor U6238 (N_6238,N_2432,N_707);
nand U6239 (N_6239,N_1910,N_1140);
or U6240 (N_6240,N_1410,N_1057);
and U6241 (N_6241,N_2483,N_324);
nand U6242 (N_6242,N_799,N_368);
and U6243 (N_6243,N_1718,N_196);
nor U6244 (N_6244,N_2951,N_702);
nor U6245 (N_6245,N_2636,N_2655);
nor U6246 (N_6246,N_874,N_435);
nand U6247 (N_6247,N_1824,N_1357);
nand U6248 (N_6248,N_227,N_973);
nor U6249 (N_6249,N_2694,N_564);
nand U6250 (N_6250,N_5381,N_3608);
or U6251 (N_6251,N_6234,N_3230);
and U6252 (N_6252,N_4462,N_5780);
or U6253 (N_6253,N_3178,N_3697);
nand U6254 (N_6254,N_3856,N_4684);
nand U6255 (N_6255,N_4700,N_5206);
or U6256 (N_6256,N_4236,N_5695);
or U6257 (N_6257,N_5337,N_6088);
and U6258 (N_6258,N_4591,N_4532);
xnor U6259 (N_6259,N_5533,N_3583);
and U6260 (N_6260,N_5476,N_3367);
xnor U6261 (N_6261,N_3813,N_3366);
nor U6262 (N_6262,N_5866,N_5768);
or U6263 (N_6263,N_5443,N_5700);
or U6264 (N_6264,N_3911,N_5336);
nand U6265 (N_6265,N_4194,N_4877);
and U6266 (N_6266,N_5123,N_4812);
and U6267 (N_6267,N_5873,N_5774);
xnor U6268 (N_6268,N_4606,N_5257);
and U6269 (N_6269,N_4637,N_4414);
and U6270 (N_6270,N_5924,N_3532);
xnor U6271 (N_6271,N_3896,N_4614);
or U6272 (N_6272,N_4324,N_5815);
or U6273 (N_6273,N_5893,N_4650);
nand U6274 (N_6274,N_3933,N_4670);
or U6275 (N_6275,N_4165,N_5937);
nand U6276 (N_6276,N_3199,N_4796);
and U6277 (N_6277,N_4379,N_5687);
nand U6278 (N_6278,N_5878,N_4091);
or U6279 (N_6279,N_4663,N_4367);
and U6280 (N_6280,N_5142,N_5931);
or U6281 (N_6281,N_6173,N_4973);
and U6282 (N_6282,N_4003,N_4264);
or U6283 (N_6283,N_3486,N_3257);
or U6284 (N_6284,N_3320,N_3333);
or U6285 (N_6285,N_6110,N_5560);
nand U6286 (N_6286,N_4951,N_6170);
or U6287 (N_6287,N_5602,N_4911);
nand U6288 (N_6288,N_6013,N_5761);
nor U6289 (N_6289,N_4660,N_3809);
xnor U6290 (N_6290,N_3397,N_5694);
nor U6291 (N_6291,N_4238,N_6019);
and U6292 (N_6292,N_4043,N_5391);
or U6293 (N_6293,N_3742,N_4335);
or U6294 (N_6294,N_5124,N_3679);
or U6295 (N_6295,N_3248,N_3326);
nand U6296 (N_6296,N_6080,N_6249);
and U6297 (N_6297,N_3187,N_3473);
nor U6298 (N_6298,N_4035,N_5184);
nor U6299 (N_6299,N_6078,N_3940);
or U6300 (N_6300,N_5788,N_3380);
and U6301 (N_6301,N_3400,N_3800);
nand U6302 (N_6302,N_3368,N_3492);
and U6303 (N_6303,N_3871,N_5906);
nand U6304 (N_6304,N_4653,N_3146);
nor U6305 (N_6305,N_3381,N_4084);
nand U6306 (N_6306,N_5351,N_3711);
or U6307 (N_6307,N_4546,N_3131);
or U6308 (N_6308,N_6193,N_5222);
and U6309 (N_6309,N_3924,N_4031);
or U6310 (N_6310,N_4867,N_3716);
nand U6311 (N_6311,N_5753,N_4064);
nor U6312 (N_6312,N_4348,N_4480);
nand U6313 (N_6313,N_3195,N_5935);
or U6314 (N_6314,N_5287,N_3653);
nor U6315 (N_6315,N_4928,N_5224);
nand U6316 (N_6316,N_5959,N_3233);
nor U6317 (N_6317,N_4328,N_6021);
or U6318 (N_6318,N_4799,N_6201);
xor U6319 (N_6319,N_4548,N_5590);
nor U6320 (N_6320,N_5892,N_5739);
nor U6321 (N_6321,N_5288,N_4069);
nor U6322 (N_6322,N_5290,N_3929);
or U6323 (N_6323,N_4890,N_5423);
xnor U6324 (N_6324,N_4547,N_4773);
and U6325 (N_6325,N_3701,N_4390);
and U6326 (N_6326,N_5395,N_3151);
nor U6327 (N_6327,N_4932,N_3126);
and U6328 (N_6328,N_3755,N_4057);
and U6329 (N_6329,N_3884,N_4125);
or U6330 (N_6330,N_4242,N_3877);
nor U6331 (N_6331,N_5131,N_3694);
nand U6332 (N_6332,N_4166,N_5660);
and U6333 (N_6333,N_5238,N_4254);
nor U6334 (N_6334,N_4876,N_4387);
or U6335 (N_6335,N_4730,N_5921);
or U6336 (N_6336,N_4446,N_4572);
xnor U6337 (N_6337,N_5281,N_3689);
nand U6338 (N_6338,N_5200,N_6075);
nand U6339 (N_6339,N_3406,N_5862);
or U6340 (N_6340,N_6211,N_4195);
nand U6341 (N_6341,N_6017,N_4474);
or U6342 (N_6342,N_3338,N_5932);
or U6343 (N_6343,N_4272,N_5625);
and U6344 (N_6344,N_3311,N_6095);
or U6345 (N_6345,N_4226,N_4163);
nand U6346 (N_6346,N_5562,N_4962);
or U6347 (N_6347,N_3942,N_4169);
nand U6348 (N_6348,N_6109,N_5059);
nor U6349 (N_6349,N_4409,N_4327);
or U6350 (N_6350,N_4838,N_3916);
nor U6351 (N_6351,N_5865,N_3547);
nand U6352 (N_6352,N_5332,N_3798);
and U6353 (N_6353,N_4120,N_3594);
nor U6354 (N_6354,N_3510,N_3231);
nand U6355 (N_6355,N_3518,N_4981);
nand U6356 (N_6356,N_6083,N_4837);
nor U6357 (N_6357,N_3585,N_5573);
and U6358 (N_6358,N_4600,N_3279);
xnor U6359 (N_6359,N_4373,N_4997);
nand U6360 (N_6360,N_5568,N_3981);
and U6361 (N_6361,N_5690,N_4174);
or U6362 (N_6362,N_5116,N_5601);
and U6363 (N_6363,N_4610,N_6217);
xnor U6364 (N_6364,N_4842,N_3729);
xnor U6365 (N_6365,N_4630,N_6244);
xor U6366 (N_6366,N_5555,N_3165);
xor U6367 (N_6367,N_5756,N_5699);
and U6368 (N_6368,N_5745,N_5772);
nand U6369 (N_6369,N_5249,N_3502);
and U6370 (N_6370,N_4384,N_3853);
xor U6371 (N_6371,N_3391,N_4449);
and U6372 (N_6372,N_3521,N_3150);
and U6373 (N_6373,N_4819,N_6206);
nand U6374 (N_6374,N_4252,N_5449);
or U6375 (N_6375,N_4419,N_5090);
nand U6376 (N_6376,N_4578,N_4185);
or U6377 (N_6377,N_5159,N_5017);
nand U6378 (N_6378,N_5913,N_5737);
nand U6379 (N_6379,N_3698,N_4398);
or U6380 (N_6380,N_5342,N_5556);
or U6381 (N_6381,N_5520,N_4427);
and U6382 (N_6382,N_5842,N_4391);
and U6383 (N_6383,N_5538,N_3321);
nor U6384 (N_6384,N_4726,N_4229);
nor U6385 (N_6385,N_4464,N_4960);
or U6386 (N_6386,N_3953,N_3720);
nor U6387 (N_6387,N_3724,N_5736);
nand U6388 (N_6388,N_4022,N_3703);
xor U6389 (N_6389,N_5604,N_4457);
nand U6390 (N_6390,N_5161,N_4692);
xor U6391 (N_6391,N_3444,N_5480);
or U6392 (N_6392,N_5528,N_3985);
xor U6393 (N_6393,N_6241,N_3948);
or U6394 (N_6394,N_4127,N_4790);
xor U6395 (N_6395,N_4130,N_5995);
and U6396 (N_6396,N_4400,N_4710);
xor U6397 (N_6397,N_3374,N_5697);
nand U6398 (N_6398,N_5759,N_5997);
or U6399 (N_6399,N_3616,N_4787);
or U6400 (N_6400,N_3978,N_3892);
or U6401 (N_6401,N_5554,N_3312);
and U6402 (N_6402,N_4941,N_3354);
nor U6403 (N_6403,N_3750,N_3261);
nand U6404 (N_6404,N_4622,N_3297);
or U6405 (N_6405,N_5484,N_3386);
or U6406 (N_6406,N_3474,N_5198);
and U6407 (N_6407,N_4098,N_3964);
nor U6408 (N_6408,N_4293,N_4370);
xnor U6409 (N_6409,N_4891,N_4786);
nand U6410 (N_6410,N_3991,N_5171);
or U6411 (N_6411,N_4306,N_3456);
and U6412 (N_6412,N_5872,N_5647);
nor U6413 (N_6413,N_5170,N_6068);
xnor U6414 (N_6414,N_6132,N_3427);
and U6415 (N_6415,N_4027,N_5269);
and U6416 (N_6416,N_5195,N_4055);
and U6417 (N_6417,N_4109,N_6098);
xor U6418 (N_6418,N_3967,N_4744);
nand U6419 (N_6419,N_5838,N_3707);
or U6420 (N_6420,N_3515,N_3477);
and U6421 (N_6421,N_4080,N_5707);
and U6422 (N_6422,N_4143,N_4586);
nand U6423 (N_6423,N_5466,N_5631);
nand U6424 (N_6424,N_5826,N_4683);
nor U6425 (N_6425,N_4643,N_5905);
or U6426 (N_6426,N_4340,N_5855);
nor U6427 (N_6427,N_3822,N_5596);
nor U6428 (N_6428,N_3905,N_3169);
nand U6429 (N_6429,N_6090,N_5714);
nor U6430 (N_6430,N_5851,N_3156);
nor U6431 (N_6431,N_4281,N_4524);
and U6432 (N_6432,N_4249,N_3251);
or U6433 (N_6433,N_3268,N_5672);
and U6434 (N_6434,N_3635,N_4447);
nand U6435 (N_6435,N_4346,N_6000);
or U6436 (N_6436,N_5722,N_5091);
or U6437 (N_6437,N_4804,N_4216);
nor U6438 (N_6438,N_4171,N_3392);
and U6439 (N_6439,N_3776,N_4571);
nor U6440 (N_6440,N_5086,N_3954);
nand U6441 (N_6441,N_4605,N_3564);
or U6442 (N_6442,N_3936,N_4705);
or U6443 (N_6443,N_3470,N_3791);
nand U6444 (N_6444,N_3795,N_4312);
nand U6445 (N_6445,N_5369,N_4843);
or U6446 (N_6446,N_5296,N_4634);
nand U6447 (N_6447,N_5825,N_5819);
and U6448 (N_6448,N_5233,N_3399);
xnor U6449 (N_6449,N_5444,N_5472);
xnor U6450 (N_6450,N_3715,N_4679);
nand U6451 (N_6451,N_3203,N_5664);
xor U6452 (N_6452,N_5817,N_3580);
xor U6453 (N_6453,N_5505,N_4501);
and U6454 (N_6454,N_3134,N_4523);
or U6455 (N_6455,N_4051,N_4018);
xor U6456 (N_6456,N_3555,N_4428);
nor U6457 (N_6457,N_4158,N_3304);
nor U6458 (N_6458,N_5183,N_4826);
nand U6459 (N_6459,N_4193,N_3331);
nand U6460 (N_6460,N_4302,N_3420);
and U6461 (N_6461,N_5529,N_6099);
nand U6462 (N_6462,N_5909,N_6200);
xnor U6463 (N_6463,N_5082,N_3272);
and U6464 (N_6464,N_6199,N_3970);
or U6465 (N_6465,N_5470,N_4349);
nor U6466 (N_6466,N_4511,N_4270);
and U6467 (N_6467,N_6052,N_3699);
nor U6468 (N_6468,N_5080,N_5823);
nor U6469 (N_6469,N_4994,N_4934);
nand U6470 (N_6470,N_4062,N_5122);
and U6471 (N_6471,N_5039,N_5532);
nor U6472 (N_6472,N_5515,N_3411);
or U6473 (N_6473,N_4023,N_4658);
nor U6474 (N_6474,N_5534,N_5099);
and U6475 (N_6475,N_3834,N_3211);
or U6476 (N_6476,N_4386,N_3686);
xnor U6477 (N_6477,N_5278,N_5521);
or U6478 (N_6478,N_4296,N_4138);
nor U6479 (N_6479,N_4694,N_4937);
or U6480 (N_6480,N_5936,N_4082);
nand U6481 (N_6481,N_3641,N_5957);
or U6482 (N_6482,N_3620,N_5225);
nand U6483 (N_6483,N_4543,N_4963);
xnor U6484 (N_6484,N_4151,N_5055);
and U6485 (N_6485,N_5552,N_3757);
nor U6486 (N_6486,N_6005,N_6081);
and U6487 (N_6487,N_5510,N_4186);
xnor U6488 (N_6488,N_5158,N_5971);
nor U6489 (N_6489,N_4172,N_3493);
and U6490 (N_6490,N_3622,N_5375);
and U6491 (N_6491,N_4331,N_4835);
or U6492 (N_6492,N_4682,N_4800);
and U6493 (N_6493,N_5926,N_4823);
and U6494 (N_6494,N_5495,N_3524);
or U6495 (N_6495,N_5329,N_4781);
nor U6496 (N_6496,N_5481,N_6062);
or U6497 (N_6497,N_5946,N_3219);
nor U6498 (N_6498,N_3952,N_6187);
nor U6499 (N_6499,N_4639,N_4797);
nor U6500 (N_6500,N_5689,N_3447);
and U6501 (N_6501,N_4515,N_5175);
nor U6502 (N_6502,N_4265,N_4661);
and U6503 (N_6503,N_5945,N_5150);
nor U6504 (N_6504,N_3475,N_4103);
nor U6505 (N_6505,N_4013,N_5379);
xnor U6506 (N_6506,N_5255,N_5034);
xnor U6507 (N_6507,N_4672,N_3300);
nand U6508 (N_6508,N_5377,N_5852);
or U6509 (N_6509,N_3323,N_3566);
nor U6510 (N_6510,N_6014,N_6054);
and U6511 (N_6511,N_6022,N_5447);
xnor U6512 (N_6512,N_6100,N_5477);
and U6513 (N_6513,N_5634,N_4279);
xnor U6514 (N_6514,N_4609,N_4319);
nor U6515 (N_6515,N_3874,N_4540);
nor U6516 (N_6516,N_5570,N_6148);
and U6517 (N_6517,N_3693,N_4521);
nor U6518 (N_6518,N_3543,N_4649);
or U6519 (N_6519,N_4137,N_3271);
or U6520 (N_6520,N_3783,N_3662);
nor U6521 (N_6521,N_3844,N_5733);
nand U6522 (N_6522,N_5147,N_4045);
nor U6523 (N_6523,N_3173,N_5637);
or U6524 (N_6524,N_6191,N_6026);
and U6525 (N_6525,N_5574,N_4341);
or U6526 (N_6526,N_5084,N_3328);
nand U6527 (N_6527,N_5681,N_4536);
or U6528 (N_6528,N_4121,N_6006);
and U6529 (N_6529,N_4374,N_5870);
xor U6530 (N_6530,N_6167,N_4453);
xor U6531 (N_6531,N_5209,N_6036);
and U6532 (N_6532,N_4085,N_5092);
nand U6533 (N_6533,N_3973,N_3557);
and U6534 (N_6534,N_4263,N_4714);
nor U6535 (N_6535,N_3604,N_4231);
or U6536 (N_6536,N_3295,N_3968);
nand U6537 (N_6537,N_4984,N_3546);
nor U6538 (N_6538,N_5954,N_4383);
nor U6539 (N_6539,N_3784,N_3476);
and U6540 (N_6540,N_3868,N_4982);
and U6541 (N_6541,N_4198,N_3728);
and U6542 (N_6542,N_3434,N_5758);
and U6543 (N_6543,N_3950,N_5857);
nor U6544 (N_6544,N_3215,N_4320);
and U6545 (N_6545,N_4880,N_3225);
or U6546 (N_6546,N_4844,N_4607);
or U6547 (N_6547,N_5322,N_4757);
nor U6548 (N_6548,N_3269,N_3188);
or U6549 (N_6549,N_5478,N_5833);
nor U6550 (N_6550,N_3445,N_5549);
xnor U6551 (N_6551,N_4778,N_5891);
nor U6552 (N_6552,N_4645,N_5008);
or U6553 (N_6553,N_3607,N_3569);
nor U6554 (N_6554,N_5112,N_4758);
and U6555 (N_6555,N_4197,N_4865);
and U6556 (N_6556,N_4030,N_5302);
nand U6557 (N_6557,N_3627,N_4215);
nor U6558 (N_6558,N_3424,N_4104);
xor U6559 (N_6559,N_3988,N_3930);
xor U6560 (N_6560,N_3530,N_4228);
nand U6561 (N_6561,N_6057,N_3598);
nand U6562 (N_6562,N_4925,N_3529);
nand U6563 (N_6563,N_4581,N_5939);
nor U6564 (N_6564,N_5769,N_5189);
and U6565 (N_6565,N_6015,N_3505);
and U6566 (N_6566,N_4316,N_4184);
xor U6567 (N_6567,N_4514,N_4957);
nand U6568 (N_6568,N_5650,N_4967);
xnor U6569 (N_6569,N_3992,N_3370);
or U6570 (N_6570,N_5474,N_3390);
and U6571 (N_6571,N_4820,N_4140);
or U6572 (N_6572,N_4841,N_4964);
nand U6573 (N_6573,N_5215,N_5718);
nor U6574 (N_6574,N_6212,N_4564);
nand U6575 (N_6575,N_3943,N_5176);
nor U6576 (N_6576,N_5600,N_5900);
xor U6577 (N_6577,N_3623,N_5847);
or U6578 (N_6578,N_4202,N_4741);
and U6579 (N_6579,N_4971,N_3612);
nor U6580 (N_6580,N_4083,N_3654);
or U6581 (N_6581,N_4274,N_3639);
or U6582 (N_6582,N_3717,N_5916);
and U6583 (N_6583,N_4931,N_5339);
nor U6584 (N_6584,N_5599,N_5563);
nand U6585 (N_6585,N_5607,N_3408);
nor U6586 (N_6586,N_3153,N_3266);
or U6587 (N_6587,N_5103,N_5557);
and U6588 (N_6588,N_3565,N_5543);
nand U6589 (N_6589,N_5948,N_6119);
or U6590 (N_6590,N_3241,N_4845);
nor U6591 (N_6591,N_5861,N_3306);
or U6592 (N_6592,N_4821,N_3168);
nand U6593 (N_6593,N_3252,N_3850);
nand U6594 (N_6594,N_4164,N_4351);
and U6595 (N_6595,N_3223,N_4979);
nand U6596 (N_6596,N_3920,N_3522);
and U6597 (N_6597,N_3377,N_4834);
and U6598 (N_6598,N_5965,N_5797);
nor U6599 (N_6599,N_4525,N_5187);
nand U6600 (N_6600,N_5335,N_6242);
or U6601 (N_6601,N_4577,N_4853);
and U6602 (N_6602,N_5307,N_4733);
or U6603 (N_6603,N_4950,N_3365);
nor U6604 (N_6604,N_4106,N_5778);
and U6605 (N_6605,N_3576,N_3862);
or U6606 (N_6606,N_6011,N_4095);
and U6607 (N_6607,N_4918,N_5007);
and U6608 (N_6608,N_4053,N_4422);
and U6609 (N_6609,N_6016,N_5723);
or U6610 (N_6610,N_4396,N_3253);
nor U6611 (N_6611,N_4305,N_5950);
and U6612 (N_6612,N_5360,N_4065);
nand U6613 (N_6613,N_3431,N_3334);
or U6614 (N_6614,N_3976,N_3708);
nor U6615 (N_6615,N_5386,N_5999);
and U6616 (N_6616,N_4233,N_3472);
nand U6617 (N_6617,N_5643,N_4776);
nor U6618 (N_6618,N_4795,N_4680);
nand U6619 (N_6619,N_5422,N_4872);
nand U6620 (N_6620,N_5834,N_5076);
and U6621 (N_6621,N_4015,N_3881);
and U6622 (N_6622,N_5621,N_5575);
and U6623 (N_6623,N_4417,N_5160);
and U6624 (N_6624,N_4459,N_5194);
nand U6625 (N_6625,N_5345,N_4775);
xnor U6626 (N_6626,N_3925,N_5738);
and U6627 (N_6627,N_5294,N_3574);
or U6628 (N_6628,N_5720,N_5874);
or U6629 (N_6629,N_5743,N_3221);
nand U6630 (N_6630,N_4128,N_4308);
nand U6631 (N_6631,N_3739,N_3305);
xnor U6632 (N_6632,N_4731,N_4557);
xnor U6633 (N_6633,N_4291,N_5791);
and U6634 (N_6634,N_4580,N_5393);
nor U6635 (N_6635,N_4256,N_5668);
and U6636 (N_6636,N_5514,N_4874);
or U6637 (N_6637,N_5982,N_5646);
nor U6638 (N_6638,N_4033,N_6227);
nand U6639 (N_6639,N_5418,N_4756);
xor U6640 (N_6640,N_3861,N_4531);
and U6641 (N_6641,N_3316,N_4538);
nand U6642 (N_6642,N_3412,N_4519);
or U6643 (N_6643,N_3175,N_3176);
nor U6644 (N_6644,N_4403,N_4839);
nor U6645 (N_6645,N_6152,N_3944);
nand U6646 (N_6646,N_4850,N_4401);
and U6647 (N_6647,N_4569,N_6065);
nand U6648 (N_6648,N_5093,N_5106);
or U6649 (N_6649,N_4440,N_5485);
and U6650 (N_6650,N_5962,N_4750);
nor U6651 (N_6651,N_5615,N_4155);
nand U6652 (N_6652,N_5102,N_5306);
nor U6653 (N_6653,N_3688,N_3875);
xor U6654 (N_6654,N_3563,N_5657);
and U6655 (N_6655,N_4977,N_6149);
xor U6656 (N_6656,N_3945,N_3603);
and U6657 (N_6657,N_4878,N_4259);
nor U6658 (N_6658,N_5289,N_3197);
nand U6659 (N_6659,N_5513,N_3632);
and U6660 (N_6660,N_4154,N_3586);
nand U6661 (N_6661,N_4014,N_5108);
nor U6662 (N_6662,N_4418,N_5998);
and U6663 (N_6663,N_5491,N_5760);
nand U6664 (N_6664,N_4101,N_5585);
or U6665 (N_6665,N_4528,N_5859);
nand U6666 (N_6666,N_5312,N_4000);
or U6667 (N_6667,N_4412,N_4631);
or U6668 (N_6668,N_3143,N_5250);
and U6669 (N_6669,N_4587,N_3613);
nand U6670 (N_6670,N_5830,N_3413);
nor U6671 (N_6671,N_4004,N_3651);
or U6672 (N_6672,N_5490,N_4475);
nand U6673 (N_6673,N_3805,N_5276);
nor U6674 (N_6674,N_3907,N_6060);
or U6675 (N_6675,N_4005,N_4170);
or U6676 (N_6676,N_6174,N_5373);
nand U6677 (N_6677,N_5070,N_3696);
or U6678 (N_6678,N_4503,N_3423);
nand U6679 (N_6679,N_5938,N_4300);
and U6680 (N_6680,N_4240,N_3573);
and U6681 (N_6681,N_5029,N_4992);
or U6682 (N_6682,N_5078,N_4722);
nand U6683 (N_6683,N_3508,N_3509);
or U6684 (N_6684,N_5144,N_3275);
nor U6685 (N_6685,N_5525,N_4806);
nand U6686 (N_6686,N_4460,N_5002);
and U6687 (N_6687,N_4477,N_5115);
nand U6688 (N_6688,N_4991,N_4691);
nor U6689 (N_6689,N_5344,N_3733);
and U6690 (N_6690,N_3799,N_6131);
nand U6691 (N_6691,N_6116,N_4421);
nor U6692 (N_6692,N_3990,N_4554);
xor U6693 (N_6693,N_4869,N_3719);
and U6694 (N_6694,N_5710,N_5219);
nand U6695 (N_6695,N_6144,N_3900);
nand U6696 (N_6696,N_5740,N_5911);
and U6697 (N_6697,N_5450,N_5097);
nand U6698 (N_6698,N_3727,N_5058);
or U6699 (N_6699,N_5064,N_6097);
and U6700 (N_6700,N_3910,N_3644);
nor U6701 (N_6701,N_5026,N_5612);
nor U6702 (N_6702,N_3352,N_4136);
nand U6703 (N_6703,N_3647,N_5915);
and U6704 (N_6704,N_6111,N_5461);
nor U6705 (N_6705,N_3845,N_5502);
xnor U6706 (N_6706,N_5149,N_4956);
or U6707 (N_6707,N_4555,N_5241);
nand U6708 (N_6708,N_3702,N_3244);
and U6709 (N_6709,N_3359,N_3155);
nand U6710 (N_6710,N_5109,N_3571);
nand U6711 (N_6711,N_4150,N_4006);
xnor U6712 (N_6712,N_3414,N_5440);
or U6713 (N_6713,N_5696,N_5676);
or U6714 (N_6714,N_4219,N_4513);
nor U6715 (N_6715,N_4613,N_6164);
nand U6716 (N_6716,N_6226,N_3303);
nand U6717 (N_6717,N_5500,N_4881);
xor U6718 (N_6718,N_3590,N_4445);
nor U6719 (N_6719,N_3764,N_5885);
or U6720 (N_6720,N_6045,N_6176);
nor U6721 (N_6721,N_4073,N_5782);
nand U6722 (N_6722,N_5776,N_5114);
or U6723 (N_6723,N_5677,N_5035);
and U6724 (N_6724,N_4489,N_3914);
or U6725 (N_6725,N_4725,N_5263);
or U6726 (N_6726,N_4141,N_5271);
or U6727 (N_6727,N_5519,N_4811);
nor U6728 (N_6728,N_5894,N_4719);
nor U6729 (N_6729,N_4019,N_3322);
and U6730 (N_6730,N_4598,N_3227);
or U6731 (N_6731,N_3148,N_5617);
nand U6732 (N_6732,N_5104,N_3676);
nand U6733 (N_6733,N_3852,N_5280);
nor U6734 (N_6734,N_3684,N_4632);
nand U6735 (N_6735,N_4404,N_4798);
nor U6736 (N_6736,N_5436,N_3706);
and U6737 (N_6737,N_5839,N_3759);
nor U6738 (N_6738,N_5488,N_5914);
nand U6739 (N_6739,N_4189,N_3483);
nor U6740 (N_6740,N_4153,N_3356);
nor U6741 (N_6741,N_3544,N_4640);
nor U6742 (N_6742,N_3927,N_4350);
or U6743 (N_6743,N_3130,N_5473);
or U6744 (N_6744,N_3226,N_3749);
or U6745 (N_6745,N_5498,N_3831);
and U6746 (N_6746,N_4667,N_4146);
nor U6747 (N_6747,N_5662,N_5348);
or U6748 (N_6748,N_5688,N_3440);
nor U6749 (N_6749,N_5037,N_4668);
or U6750 (N_6750,N_6033,N_3705);
and U6751 (N_6751,N_4251,N_6168);
or U6752 (N_6752,N_4774,N_4855);
and U6753 (N_6753,N_4468,N_4058);
and U6754 (N_6754,N_5813,N_4070);
or U6755 (N_6755,N_4659,N_6118);
nor U6756 (N_6756,N_5486,N_4802);
nand U6757 (N_6757,N_3873,N_4875);
nand U6758 (N_6758,N_4448,N_4135);
nand U6759 (N_6759,N_4735,N_4126);
nand U6760 (N_6760,N_5433,N_4192);
nor U6761 (N_6761,N_4830,N_3235);
nand U6762 (N_6762,N_5648,N_5889);
and U6763 (N_6763,N_4119,N_5057);
and U6764 (N_6764,N_5191,N_4945);
nand U6765 (N_6765,N_5493,N_3606);
nor U6766 (N_6766,N_4914,N_3194);
xor U6767 (N_6767,N_4688,N_5185);
nor U6768 (N_6768,N_3490,N_4225);
nor U6769 (N_6769,N_4717,N_5432);
and U6770 (N_6770,N_5275,N_6042);
nand U6771 (N_6771,N_6020,N_6221);
nand U6772 (N_6772,N_4323,N_4675);
nand U6773 (N_6773,N_3670,N_4870);
and U6774 (N_6774,N_4618,N_6114);
nor U6775 (N_6775,N_6072,N_3329);
or U6776 (N_6776,N_3682,N_3640);
and U6777 (N_6777,N_4970,N_5445);
or U6778 (N_6778,N_5483,N_3232);
nor U6779 (N_6779,N_3299,N_3164);
nor U6780 (N_6780,N_3288,N_4534);
and U6781 (N_6781,N_4708,N_4552);
and U6782 (N_6782,N_4212,N_4282);
or U6783 (N_6783,N_5096,N_4122);
nand U6784 (N_6784,N_5441,N_5412);
or U6785 (N_6785,N_3821,N_3779);
and U6786 (N_6786,N_5934,N_5073);
or U6787 (N_6787,N_5674,N_4326);
or U6788 (N_6788,N_5673,N_3658);
nand U6789 (N_6789,N_4885,N_6117);
nor U6790 (N_6790,N_5392,N_5989);
nor U6791 (N_6791,N_5616,N_3315);
nor U6792 (N_6792,N_3752,N_5282);
nor U6793 (N_6793,N_4368,N_5409);
xor U6794 (N_6794,N_4026,N_5179);
or U6795 (N_6795,N_3216,N_5460);
and U6796 (N_6796,N_3541,N_3828);
or U6797 (N_6797,N_4451,N_5884);
nand U6798 (N_6798,N_3403,N_3959);
or U6799 (N_6799,N_6240,N_5136);
or U6800 (N_6800,N_4042,N_5651);
nand U6801 (N_6801,N_4793,N_4338);
nand U6802 (N_6802,N_5917,N_4913);
xnor U6803 (N_6803,N_6163,N_5658);
and U6804 (N_6804,N_5414,N_6082);
nor U6805 (N_6805,N_5779,N_3963);
nand U6806 (N_6806,N_4673,N_6179);
or U6807 (N_6807,N_3888,N_5614);
or U6808 (N_6808,N_4676,N_4160);
nor U6809 (N_6809,N_5321,N_6048);
or U6810 (N_6810,N_4686,N_4079);
nand U6811 (N_6811,N_5065,N_5652);
and U6812 (N_6812,N_5050,N_5221);
nand U6813 (N_6813,N_3401,N_4309);
or U6814 (N_6814,N_4167,N_4333);
and U6815 (N_6815,N_3325,N_4039);
nand U6816 (N_6816,N_3382,N_4727);
and U6817 (N_6817,N_4582,N_5589);
nand U6818 (N_6818,N_4092,N_4180);
nand U6819 (N_6819,N_6077,N_4310);
nor U6820 (N_6820,N_5877,N_4585);
nand U6821 (N_6821,N_3840,N_5749);
nor U6822 (N_6822,N_4638,N_3767);
and U6823 (N_6823,N_5388,N_5069);
nor U6824 (N_6824,N_3860,N_5773);
or U6825 (N_6825,N_3723,N_6051);
and U6826 (N_6826,N_6120,N_4280);
nor U6827 (N_6827,N_6123,N_4801);
nor U6828 (N_6828,N_3673,N_4900);
and U6829 (N_6829,N_4247,N_4220);
nor U6830 (N_6830,N_3931,N_5644);
and U6831 (N_6831,N_5169,N_4243);
nor U6832 (N_6832,N_4199,N_3897);
or U6833 (N_6833,N_6053,N_4919);
or U6834 (N_6834,N_5357,N_6038);
nor U6835 (N_6835,N_5795,N_5794);
nor U6836 (N_6836,N_6030,N_6230);
nand U6837 (N_6837,N_3637,N_4807);
and U6838 (N_6838,N_4205,N_5875);
and U6839 (N_6839,N_4382,N_4846);
and U6840 (N_6840,N_4187,N_5374);
or U6841 (N_6841,N_3903,N_5014);
and U6842 (N_6842,N_3344,N_3738);
nand U6843 (N_6843,N_3672,N_3584);
nand U6844 (N_6844,N_6247,N_5633);
xor U6845 (N_6845,N_5202,N_5622);
and U6846 (N_6846,N_3245,N_4235);
or U6847 (N_6847,N_6073,N_4810);
or U6848 (N_6848,N_3204,N_3436);
or U6849 (N_6849,N_5820,N_4353);
or U6850 (N_6850,N_3770,N_3499);
or U6851 (N_6851,N_4856,N_5802);
and U6852 (N_6852,N_3763,N_5558);
nand U6853 (N_6853,N_5553,N_5805);
nor U6854 (N_6854,N_6223,N_3934);
nor U6855 (N_6855,N_3885,N_4413);
xor U6856 (N_6856,N_5990,N_5299);
xnor U6857 (N_6857,N_5033,N_3928);
and U6858 (N_6858,N_5027,N_4635);
nand U6859 (N_6859,N_4500,N_5804);
nand U6860 (N_6860,N_3298,N_5462);
nor U6861 (N_6861,N_3904,N_4123);
nand U6862 (N_6862,N_3213,N_5132);
nand U6863 (N_6863,N_3357,N_4953);
nand U6864 (N_6864,N_4737,N_4828);
and U6865 (N_6865,N_3459,N_4753);
and U6866 (N_6866,N_3319,N_3558);
xor U6867 (N_6867,N_3296,N_5579);
and U6868 (N_6868,N_4207,N_3506);
nand U6869 (N_6869,N_5085,N_5693);
and U6870 (N_6870,N_3249,N_5811);
nor U6871 (N_6871,N_5846,N_3207);
nor U6872 (N_6872,N_4752,N_4294);
nor U6873 (N_6873,N_5783,N_3777);
nand U6874 (N_6874,N_4224,N_3376);
or U6875 (N_6875,N_5487,N_4077);
or U6876 (N_6876,N_4822,N_5992);
and U6877 (N_6877,N_3250,N_5364);
and U6878 (N_6878,N_4740,N_5709);
xnor U6879 (N_6879,N_6074,N_4481);
nand U6880 (N_6880,N_4952,N_4048);
and U6881 (N_6881,N_3274,N_4943);
nand U6882 (N_6882,N_3210,N_4176);
or U6883 (N_6883,N_3388,N_5972);
nand U6884 (N_6884,N_5904,N_5564);
nor U6885 (N_6885,N_5214,N_5829);
or U6886 (N_6886,N_5654,N_5787);
xnor U6887 (N_6887,N_3866,N_5716);
nand U6888 (N_6888,N_3807,N_5793);
nand U6889 (N_6889,N_4388,N_4720);
nor U6890 (N_6890,N_6198,N_5223);
xnor U6891 (N_6891,N_5667,N_6222);
nand U6892 (N_6892,N_3602,N_3307);
and U6893 (N_6893,N_5535,N_3731);
and U6894 (N_6894,N_5721,N_4888);
xnor U6895 (N_6895,N_3535,N_5244);
nand U6896 (N_6896,N_5272,N_5352);
nand U6897 (N_6897,N_5400,N_3318);
nand U6898 (N_6898,N_6153,N_4483);
nand U6899 (N_6899,N_4407,N_6007);
nand U6900 (N_6900,N_4873,N_5456);
nor U6901 (N_6901,N_4627,N_4611);
nor U6902 (N_6902,N_3171,N_5624);
or U6903 (N_6903,N_5482,N_4336);
and U6904 (N_6904,N_3495,N_4012);
and U6905 (N_6905,N_4271,N_6209);
and U6906 (N_6906,N_4861,N_5207);
nand U6907 (N_6907,N_4268,N_4078);
and U6908 (N_6908,N_3137,N_6246);
nor U6909 (N_6909,N_5049,N_5863);
nand U6910 (N_6910,N_3200,N_5338);
nand U6911 (N_6911,N_5266,N_5446);
nand U6912 (N_6912,N_4895,N_5277);
or U6913 (N_6913,N_4434,N_5626);
or U6914 (N_6914,N_5671,N_3190);
or U6915 (N_6915,N_5188,N_3457);
xnor U6916 (N_6916,N_4375,N_5524);
and U6917 (N_6917,N_3561,N_4779);
nand U6918 (N_6918,N_3196,N_4258);
nor U6919 (N_6919,N_4458,N_4208);
nand U6920 (N_6920,N_3977,N_3246);
and U6921 (N_6921,N_5711,N_5105);
nand U6922 (N_6922,N_3814,N_5719);
xor U6923 (N_6923,N_3396,N_6093);
xnor U6924 (N_6924,N_5967,N_5358);
or U6925 (N_6925,N_5978,N_5330);
or U6926 (N_6926,N_6184,N_5051);
nand U6927 (N_6927,N_4655,N_3935);
and U6928 (N_6928,N_5569,N_4652);
and U6929 (N_6929,N_6183,N_5196);
nand U6930 (N_6930,N_5153,N_4759);
nand U6931 (N_6931,N_6229,N_6142);
nand U6932 (N_6932,N_3138,N_5956);
or U6933 (N_6933,N_4736,N_3174);
nand U6934 (N_6934,N_3410,N_3238);
and U6935 (N_6935,N_5403,N_4946);
xnor U6936 (N_6936,N_5592,N_3479);
or U6937 (N_6937,N_3732,N_3554);
and U6938 (N_6938,N_5193,N_5887);
or U6939 (N_6939,N_5315,N_3768);
xnor U6940 (N_6940,N_4009,N_4492);
xnor U6941 (N_6941,N_3466,N_5910);
nand U6942 (N_6942,N_4502,N_5094);
or U6943 (N_6943,N_5886,N_3346);
or U6944 (N_6944,N_5765,N_5501);
xor U6945 (N_6945,N_3833,N_5832);
and U6946 (N_6946,N_3540,N_5229);
nand U6947 (N_6947,N_3422,N_4152);
or U6948 (N_6948,N_5098,N_6225);
nor U6949 (N_6949,N_3747,N_4961);
nand U6950 (N_6950,N_5044,N_6044);
or U6951 (N_6951,N_4729,N_4342);
or U6952 (N_6952,N_6195,N_4966);
nor U6953 (N_6953,N_5240,N_6181);
nand U6954 (N_6954,N_6239,N_4295);
or U6955 (N_6955,N_5750,N_3618);
and U6956 (N_6956,N_5228,N_6087);
or U6957 (N_6957,N_3562,N_5670);
and U6958 (N_6958,N_4408,N_3157);
or U6959 (N_6959,N_5593,N_5426);
nor U6960 (N_6960,N_3497,N_4411);
or U6961 (N_6961,N_5212,N_3726);
nand U6962 (N_6962,N_3278,N_4938);
nor U6963 (N_6963,N_3857,N_3974);
or U6964 (N_6964,N_4097,N_6189);
nand U6965 (N_6965,N_5610,N_4993);
nor U6966 (N_6966,N_6001,N_3762);
or U6967 (N_6967,N_5100,N_3291);
or U6968 (N_6968,N_4406,N_5245);
nor U6969 (N_6969,N_4399,N_4505);
nor U6970 (N_6970,N_4974,N_5043);
or U6971 (N_6971,N_4562,N_5353);
and U6972 (N_6972,N_5468,N_4542);
nand U6973 (N_6973,N_5816,N_3517);
or U6974 (N_6974,N_6186,N_5517);
or U6975 (N_6975,N_4149,N_4292);
and U6976 (N_6976,N_3551,N_4780);
and U6977 (N_6977,N_3657,N_3995);
nor U6978 (N_6978,N_6165,N_3591);
nand U6979 (N_6979,N_4442,N_4763);
nor U6980 (N_6980,N_4760,N_3465);
or U6981 (N_6981,N_3837,N_4955);
nor U6982 (N_6982,N_4232,N_4988);
and U6983 (N_6983,N_4332,N_6190);
xor U6984 (N_6984,N_5713,N_3349);
and U6985 (N_6985,N_5119,N_4990);
nor U6986 (N_6986,N_5201,N_6237);
nor U6987 (N_6987,N_5264,N_5767);
nand U6988 (N_6988,N_3969,N_3906);
nor U6989 (N_6989,N_4689,N_5645);
or U6990 (N_6990,N_5199,N_3542);
nor U6991 (N_6991,N_3849,N_4203);
nor U6992 (N_6992,N_3525,N_4443);
nor U6993 (N_6993,N_5442,N_5083);
or U6994 (N_6994,N_5691,N_4372);
nand U6995 (N_6995,N_6041,N_3678);
or U6996 (N_6996,N_3625,N_6008);
and U6997 (N_6997,N_5611,N_5363);
nand U6998 (N_6998,N_5056,N_5130);
and U6999 (N_6999,N_3690,N_3787);
or U7000 (N_7000,N_6202,N_5389);
nand U7001 (N_7001,N_3957,N_6208);
xnor U7002 (N_7002,N_5424,N_4965);
nor U7003 (N_7003,N_3824,N_3166);
nand U7004 (N_7004,N_3870,N_4743);
nand U7005 (N_7005,N_5708,N_5174);
or U7006 (N_7006,N_3956,N_3217);
nand U7007 (N_7007,N_4738,N_3534);
nand U7008 (N_7008,N_3941,N_3514);
or U7009 (N_7009,N_5331,N_4817);
or U7010 (N_7010,N_6124,N_3922);
nand U7011 (N_7011,N_6066,N_5325);
nor U7012 (N_7012,N_4892,N_5496);
nand U7013 (N_7013,N_4864,N_5996);
nand U7014 (N_7014,N_5499,N_3984);
or U7015 (N_7015,N_3765,N_3154);
nor U7016 (N_7016,N_6185,N_4766);
nor U7017 (N_7017,N_4617,N_5942);
or U7018 (N_7018,N_4604,N_4420);
or U7019 (N_7019,N_3375,N_3416);
nor U7020 (N_7020,N_4040,N_4879);
nand U7021 (N_7021,N_5620,N_4433);
or U7022 (N_7022,N_4191,N_5453);
or U7023 (N_7023,N_4923,N_4196);
or U7024 (N_7024,N_3421,N_3441);
or U7025 (N_7025,N_3961,N_3867);
nand U7026 (N_7026,N_5744,N_5507);
and U7027 (N_7027,N_5807,N_5781);
and U7028 (N_7028,N_5941,N_3484);
or U7029 (N_7029,N_4011,N_3839);
xor U7030 (N_7030,N_5291,N_3189);
nor U7031 (N_7031,N_5966,N_3258);
and U7032 (N_7032,N_4530,N_3438);
nand U7033 (N_7033,N_5853,N_5416);
or U7034 (N_7034,N_3222,N_5385);
and U7035 (N_7035,N_4887,N_3993);
xor U7036 (N_7036,N_4473,N_5741);
nor U7037 (N_7037,N_3281,N_5974);
or U7038 (N_7038,N_3224,N_4910);
xor U7039 (N_7039,N_6126,N_3671);
and U7040 (N_7040,N_4921,N_5698);
or U7041 (N_7041,N_3149,N_3327);
nand U7042 (N_7042,N_3145,N_5582);
nand U7043 (N_7043,N_5157,N_5304);
and U7044 (N_7044,N_6177,N_5679);
nand U7045 (N_7045,N_3549,N_3343);
or U7046 (N_7046,N_3259,N_4666);
or U7047 (N_7047,N_3982,N_3780);
xnor U7048 (N_7048,N_5113,N_3577);
nand U7049 (N_7049,N_5042,N_5712);
nor U7050 (N_7050,N_5818,N_3668);
or U7051 (N_7051,N_4132,N_5506);
nand U7052 (N_7052,N_3615,N_4574);
nor U7053 (N_7053,N_5952,N_4250);
and U7054 (N_7054,N_5211,N_3369);
nor U7055 (N_7055,N_5927,N_5204);
and U7056 (N_7056,N_6236,N_5869);
nand U7057 (N_7057,N_3921,N_4597);
nand U7058 (N_7058,N_3949,N_4358);
nand U7059 (N_7059,N_4550,N_6219);
or U7060 (N_7060,N_4624,N_4142);
nand U7061 (N_7061,N_3206,N_3528);
nor U7062 (N_7062,N_5584,N_4431);
nor U7063 (N_7063,N_5134,N_3309);
xor U7064 (N_7064,N_5578,N_6182);
or U7065 (N_7065,N_4486,N_4724);
or U7066 (N_7066,N_4693,N_5933);
xnor U7067 (N_7067,N_3313,N_4922);
nor U7068 (N_7068,N_4579,N_5190);
and U7069 (N_7069,N_6169,N_3433);
and U7070 (N_7070,N_3285,N_4063);
or U7071 (N_7071,N_5354,N_4437);
and U7072 (N_7072,N_4110,N_4772);
xor U7073 (N_7073,N_6150,N_4339);
nand U7074 (N_7074,N_3289,N_4222);
xor U7075 (N_7075,N_3718,N_3437);
xnor U7076 (N_7076,N_4261,N_4721);
nand U7077 (N_7077,N_3342,N_4785);
nor U7078 (N_7078,N_3277,N_4698);
or U7079 (N_7079,N_5048,N_6238);
and U7080 (N_7080,N_5730,N_4898);
xnor U7081 (N_7081,N_4381,N_5117);
or U7082 (N_7082,N_5947,N_5020);
xnor U7083 (N_7083,N_4244,N_4678);
nor U7084 (N_7084,N_4699,N_3994);
nor U7085 (N_7085,N_5635,N_5394);
and U7086 (N_7086,N_5438,N_4697);
nor U7087 (N_7087,N_5798,N_4924);
nand U7088 (N_7088,N_5448,N_5071);
nor U7089 (N_7089,N_5896,N_4337);
nand U7090 (N_7090,N_5430,N_4038);
nor U7091 (N_7091,N_4848,N_5036);
nand U7092 (N_7092,N_4541,N_5248);
or U7093 (N_7093,N_4001,N_4036);
nand U7094 (N_7094,N_4284,N_6010);
and U7095 (N_7095,N_5308,N_5040);
nand U7096 (N_7096,N_6049,N_5148);
nor U7097 (N_7097,N_5283,N_5128);
nor U7098 (N_7098,N_4329,N_3663);
and U7099 (N_7099,N_5052,N_3142);
or U7100 (N_7100,N_4628,N_3882);
xor U7101 (N_7101,N_4423,N_3980);
and U7102 (N_7102,N_5786,N_4636);
nor U7103 (N_7103,N_4702,N_6086);
or U7104 (N_7104,N_4954,N_3185);
or U7105 (N_7105,N_3597,N_6210);
nor U7106 (N_7106,N_4852,N_5561);
nor U7107 (N_7107,N_3898,N_3132);
nand U7108 (N_7108,N_3979,N_6154);
nand U7109 (N_7109,N_5881,N_3649);
nand U7110 (N_7110,N_5796,N_5066);
nor U7111 (N_7111,N_3478,N_3996);
and U7112 (N_7112,N_5365,N_4131);
xor U7113 (N_7113,N_5138,N_4245);
nand U7114 (N_7114,N_6047,N_3803);
nand U7115 (N_7115,N_5883,N_6063);
nand U7116 (N_7116,N_4463,N_5692);
nand U7117 (N_7117,N_4754,N_3704);
nand U7118 (N_7118,N_5405,N_5587);
nor U7119 (N_7119,N_4527,N_5685);
nor U7120 (N_7120,N_4405,N_5362);
nand U7121 (N_7121,N_4017,N_3141);
nor U7122 (N_7122,N_5981,N_4516);
nand U7123 (N_7123,N_6151,N_4499);
xnor U7124 (N_7124,N_4936,N_5382);
nor U7125 (N_7125,N_4866,N_3452);
and U7126 (N_7126,N_4767,N_4430);
nand U7127 (N_7127,N_3796,N_5239);
and U7128 (N_7128,N_4498,N_5822);
nor U7129 (N_7129,N_6156,N_4595);
and U7130 (N_7130,N_5594,N_3158);
and U7131 (N_7131,N_6205,N_3254);
nand U7132 (N_7132,N_5751,N_4944);
nand U7133 (N_7133,N_5273,N_4755);
nor U7134 (N_7134,N_4748,N_4010);
or U7135 (N_7135,N_5680,N_4517);
nand U7136 (N_7136,N_3409,N_5735);
nand U7137 (N_7137,N_5435,N_4602);
and U7138 (N_7138,N_4558,N_3491);
nand U7139 (N_7139,N_4813,N_5523);
nor U7140 (N_7140,N_3820,N_4986);
and U7141 (N_7141,N_3687,N_6113);
or U7142 (N_7142,N_3778,N_3462);
nor U7143 (N_7143,N_4410,N_6012);
nor U7144 (N_7144,N_4476,N_3485);
and U7145 (N_7145,N_4360,N_4642);
nand U7146 (N_7146,N_5608,N_4393);
and U7147 (N_7147,N_4076,N_3958);
xor U7148 (N_7148,N_3843,N_3516);
or U7149 (N_7149,N_3364,N_4704);
or U7150 (N_7150,N_6055,N_6136);
nand U7151 (N_7151,N_5192,N_3746);
nand U7152 (N_7152,N_5095,N_5827);
nor U7153 (N_7153,N_3301,N_4816);
or U7154 (N_7154,N_3407,N_3592);
or U7155 (N_7155,N_3363,N_5429);
or U7156 (N_7156,N_5704,N_4504);
xnor U7157 (N_7157,N_4599,N_5016);
nor U7158 (N_7158,N_5023,N_5895);
or U7159 (N_7159,N_5638,N_3205);
nand U7160 (N_7160,N_3443,N_6248);
xnor U7161 (N_7161,N_4677,N_4794);
nand U7162 (N_7162,N_5327,N_4311);
nand U7163 (N_7163,N_6161,N_5799);
nand U7164 (N_7164,N_5636,N_4262);
and U7165 (N_7165,N_5930,N_5951);
or U7166 (N_7166,N_3287,N_6231);
and U7167 (N_7167,N_5572,N_3489);
nor U7168 (N_7168,N_5133,N_5976);
and U7169 (N_7169,N_5434,N_4929);
and U7170 (N_7170,N_4690,N_4972);
and U7171 (N_7171,N_3918,N_5143);
xor U7172 (N_7172,N_5655,N_5376);
nand U7173 (N_7173,N_4402,N_4713);
nor U7174 (N_7174,N_3793,N_3152);
xnor U7175 (N_7175,N_4479,N_5237);
nand U7176 (N_7176,N_4432,N_3202);
nand U7177 (N_7177,N_4248,N_4090);
or U7178 (N_7178,N_5785,N_6112);
xnor U7179 (N_7179,N_5988,N_5928);
nand U7180 (N_7180,N_3680,N_3220);
nand U7181 (N_7181,N_3552,N_5848);
nor U7182 (N_7182,N_5539,N_6037);
or U7183 (N_7183,N_5571,N_6216);
nor U7184 (N_7184,N_4533,N_5032);
or U7185 (N_7185,N_4363,N_3519);
nor U7186 (N_7186,N_5701,N_3236);
nand U7187 (N_7187,N_4777,N_3913);
xor U7188 (N_7188,N_4825,N_5107);
and U7189 (N_7189,N_4539,N_5943);
nor U7190 (N_7190,N_4567,N_4948);
nand U7191 (N_7191,N_5489,N_5763);
or U7192 (N_7192,N_6214,N_6220);
nor U7193 (N_7193,N_5022,N_5876);
nor U7194 (N_7194,N_5411,N_4314);
nand U7195 (N_7195,N_4742,N_3139);
nor U7196 (N_7196,N_4118,N_6122);
xor U7197 (N_7197,N_5868,N_4267);
and U7198 (N_7198,N_5326,N_5208);
and U7199 (N_7199,N_3751,N_4669);
or U7200 (N_7200,N_5203,N_5279);
or U7201 (N_7201,N_5653,N_5837);
or U7202 (N_7202,N_4029,N_3270);
nor U7203 (N_7203,N_3817,N_4072);
nor U7204 (N_7204,N_5087,N_4857);
nand U7205 (N_7205,N_3209,N_3894);
and U7206 (N_7206,N_5541,N_3167);
nor U7207 (N_7207,N_5843,N_5213);
or U7208 (N_7208,N_4111,N_3480);
xnor U7209 (N_7209,N_4510,N_4487);
or U7210 (N_7210,N_3599,N_3570);
or U7211 (N_7211,N_3610,N_3290);
nor U7212 (N_7212,N_3162,N_3912);
nand U7213 (N_7213,N_3387,N_5013);
nand U7214 (N_7214,N_5060,N_4425);
and U7215 (N_7215,N_5588,N_4860);
nor U7216 (N_7216,N_5828,N_6143);
nor U7217 (N_7217,N_3402,N_5028);
or U7218 (N_7218,N_5319,N_5746);
and U7219 (N_7219,N_4380,N_3454);
and U7220 (N_7220,N_6130,N_4603);
and U7221 (N_7221,N_3435,N_4218);
xnor U7222 (N_7222,N_4046,N_6138);
and U7223 (N_7223,N_4424,N_4148);
and U7224 (N_7224,N_5151,N_3503);
nand U7225 (N_7225,N_4253,N_4495);
nor U7226 (N_7226,N_3314,N_5258);
nor U7227 (N_7227,N_4553,N_4575);
nand U7228 (N_7228,N_5018,N_5770);
nor U7229 (N_7229,N_5497,N_5724);
nor U7230 (N_7230,N_4344,N_4998);
and U7231 (N_7231,N_5469,N_4330);
nand U7232 (N_7232,N_4260,N_4145);
nand U7233 (N_7233,N_4620,N_5841);
nand U7234 (N_7234,N_5366,N_3237);
and U7235 (N_7235,N_5669,N_4392);
nand U7236 (N_7236,N_3630,N_5546);
nand U7237 (N_7237,N_4210,N_3193);
and U7238 (N_7238,N_5726,N_5300);
and U7239 (N_7239,N_4723,N_4301);
nor U7240 (N_7240,N_4978,N_5313);
xnor U7241 (N_7241,N_5010,N_6079);
and U7242 (N_7242,N_5856,N_4436);
xor U7243 (N_7243,N_3214,N_4906);
or U7244 (N_7244,N_3371,N_4859);
nor U7245 (N_7245,N_3674,N_5821);
nor U7246 (N_7246,N_3553,N_5850);
nand U7247 (N_7247,N_4315,N_5619);
and U7248 (N_7248,N_6172,N_3548);
nand U7249 (N_7249,N_5542,N_5882);
and U7250 (N_7250,N_3802,N_3451);
and U7251 (N_7251,N_3172,N_5340);
or U7252 (N_7252,N_5072,N_3582);
nor U7253 (N_7253,N_5314,N_4478);
nand U7254 (N_7254,N_3661,N_4129);
nand U7255 (N_7255,N_4469,N_4321);
nor U7256 (N_7256,N_4854,N_3520);
or U7257 (N_7257,N_5437,N_3841);
or U7258 (N_7258,N_3572,N_5235);
xor U7259 (N_7259,N_4814,N_5125);
or U7260 (N_7260,N_3946,N_3669);
and U7261 (N_7261,N_3125,N_4246);
or U7262 (N_7262,N_5025,N_3966);
nor U7263 (N_7263,N_5504,N_5297);
and U7264 (N_7264,N_4352,N_5511);
nand U7265 (N_7265,N_5577,N_4619);
xor U7266 (N_7266,N_4903,N_4901);
nor U7267 (N_7267,N_5268,N_3769);
nor U7268 (N_7268,N_3617,N_6076);
nand U7269 (N_7269,N_3737,N_3685);
nor U7270 (N_7270,N_3494,N_4450);
nand U7271 (N_7271,N_6046,N_6039);
nor U7272 (N_7272,N_5068,N_4116);
nand U7273 (N_7273,N_5459,N_5024);
nor U7274 (N_7274,N_5227,N_5661);
xnor U7275 (N_7275,N_3761,N_5372);
nand U7276 (N_7276,N_4529,N_4535);
or U7277 (N_7277,N_5784,N_4912);
and U7278 (N_7278,N_4290,N_3709);
nand U7279 (N_7279,N_4902,N_4512);
or U7280 (N_7280,N_3847,N_5531);
or U7281 (N_7281,N_3488,N_5627);
and U7282 (N_7282,N_3192,N_6160);
or U7283 (N_7283,N_5567,N_4840);
nand U7284 (N_7284,N_5285,N_5041);
nor U7285 (N_7285,N_5075,N_5421);
and U7286 (N_7286,N_4930,N_6089);
or U7287 (N_7287,N_3634,N_5605);
and U7288 (N_7288,N_3450,N_4976);
or U7289 (N_7289,N_3267,N_3198);
or U7290 (N_7290,N_4361,N_5980);
nand U7291 (N_7291,N_4134,N_4059);
nand U7292 (N_7292,N_4920,N_4144);
or U7293 (N_7293,N_5955,N_4275);
xnor U7294 (N_7294,N_5246,N_5186);
nor U7295 (N_7295,N_5452,N_6141);
and U7296 (N_7296,N_3665,N_6031);
and U7297 (N_7297,N_4664,N_4701);
and U7298 (N_7298,N_5210,N_4762);
xnor U7299 (N_7299,N_5754,N_4508);
and U7300 (N_7300,N_5021,N_4507);
nor U7301 (N_7301,N_3960,N_4371);
nand U7302 (N_7302,N_6102,N_4933);
nor U7303 (N_7303,N_6207,N_5349);
xor U7304 (N_7304,N_3302,N_4985);
nand U7305 (N_7305,N_5110,N_4695);
nand U7306 (N_7306,N_4893,N_4020);
or U7307 (N_7307,N_4803,N_3614);
xnor U7308 (N_7308,N_4102,N_3816);
and U7309 (N_7309,N_4034,N_3394);
and U7310 (N_7310,N_5686,N_4188);
xnor U7311 (N_7311,N_3596,N_5439);
nor U7312 (N_7312,N_6203,N_3575);
and U7313 (N_7313,N_6056,N_5218);
nor U7314 (N_7314,N_5925,N_3815);
or U7315 (N_7315,N_3360,N_3848);
and U7316 (N_7316,N_4556,N_5551);
nand U7317 (N_7317,N_5341,N_5178);
and U7318 (N_7318,N_3419,N_5355);
nand U7319 (N_7319,N_3545,N_5597);
nor U7320 (N_7320,N_4100,N_6002);
or U7321 (N_7321,N_3712,N_6125);
and U7322 (N_7322,N_4050,N_3876);
xnor U7323 (N_7323,N_5305,N_4908);
nand U7324 (N_7324,N_4052,N_5053);
or U7325 (N_7325,N_3760,N_3878);
or U7326 (N_7326,N_6228,N_6106);
and U7327 (N_7327,N_5417,N_4768);
and U7328 (N_7328,N_4454,N_5755);
or U7329 (N_7329,N_4177,N_6104);
nand U7330 (N_7330,N_3425,N_3336);
and U7331 (N_7331,N_5408,N_6158);
and U7332 (N_7332,N_3901,N_6115);
and U7333 (N_7333,N_4438,N_5301);
and U7334 (N_7334,N_3987,N_3611);
xnor U7335 (N_7335,N_5231,N_3247);
xnor U7336 (N_7336,N_4159,N_4060);
and U7337 (N_7337,N_4592,N_6194);
nor U7338 (N_7338,N_3983,N_5232);
nand U7339 (N_7339,N_5135,N_6155);
nand U7340 (N_7340,N_3786,N_3487);
and U7341 (N_7341,N_4147,N_3255);
or U7342 (N_7342,N_5479,N_6196);
nand U7343 (N_7343,N_3939,N_5993);
and U7344 (N_7344,N_4376,N_3794);
and U7345 (N_7345,N_3330,N_3926);
and U7346 (N_7346,N_3593,N_3341);
or U7347 (N_7347,N_3832,N_4318);
and U7348 (N_7348,N_5079,N_5898);
or U7349 (N_7349,N_5011,N_3186);
or U7350 (N_7350,N_4644,N_6050);
nor U7351 (N_7351,N_4886,N_3823);
nor U7352 (N_7352,N_3471,N_5309);
nor U7353 (N_7353,N_4633,N_4718);
or U7354 (N_7354,N_5220,N_4506);
xor U7355 (N_7355,N_4537,N_4889);
and U7356 (N_7356,N_5969,N_4863);
and U7357 (N_7357,N_4862,N_3656);
or U7358 (N_7358,N_3645,N_4178);
or U7359 (N_7359,N_6024,N_5067);
or U7360 (N_7360,N_5270,N_3496);
xor U7361 (N_7361,N_3182,N_5518);
nor U7362 (N_7362,N_6128,N_4745);
or U7363 (N_7363,N_4182,N_6145);
nand U7364 (N_7364,N_4112,N_4565);
nand U7365 (N_7365,N_4883,N_5920);
nand U7366 (N_7366,N_4739,N_4217);
xor U7367 (N_7367,N_4286,N_3523);
nor U7368 (N_7368,N_3191,N_6235);
or U7369 (N_7369,N_5262,N_4028);
and U7370 (N_7370,N_3619,N_3513);
nor U7371 (N_7371,N_5899,N_4471);
nand U7372 (N_7372,N_4646,N_3650);
and U7373 (N_7373,N_3917,N_3937);
nand U7374 (N_7374,N_5045,N_5140);
nand U7375 (N_7375,N_3439,N_5127);
or U7376 (N_7376,N_4563,N_4435);
or U7377 (N_7377,N_4851,N_6243);
nand U7378 (N_7378,N_5154,N_4313);
xor U7379 (N_7379,N_3695,N_6107);
or U7380 (N_7380,N_4926,N_3890);
nand U7381 (N_7381,N_4827,N_3710);
or U7382 (N_7382,N_6035,N_3830);
nor U7383 (N_7383,N_5404,N_5146);
nor U7384 (N_7384,N_4179,N_3998);
nand U7385 (N_7385,N_5165,N_5985);
and U7386 (N_7386,N_4615,N_5629);
or U7387 (N_7387,N_3633,N_3389);
nor U7388 (N_7388,N_4255,N_4223);
and U7389 (N_7389,N_5961,N_5001);
nor U7390 (N_7390,N_3511,N_4734);
nand U7391 (N_7391,N_5234,N_4882);
and U7392 (N_7392,N_3883,N_4175);
nor U7393 (N_7393,N_3811,N_5897);
nand U7394 (N_7394,N_5800,N_3398);
xnor U7395 (N_7395,N_5019,N_4809);
xnor U7396 (N_7396,N_3538,N_6178);
nand U7397 (N_7397,N_6146,N_3468);
nand U7398 (N_7398,N_5649,N_6094);
and U7399 (N_7399,N_3642,N_3384);
or U7400 (N_7400,N_3405,N_5004);
or U7401 (N_7401,N_3355,N_3448);
or U7402 (N_7402,N_5298,N_5923);
or U7403 (N_7403,N_5254,N_4485);
nor U7404 (N_7404,N_5402,N_4369);
nor U7405 (N_7405,N_4162,N_4596);
nor U7406 (N_7406,N_4273,N_5632);
and U7407 (N_7407,N_5731,N_4899);
or U7408 (N_7408,N_3902,N_5912);
nor U7409 (N_7409,N_5790,N_4975);
or U7410 (N_7410,N_5455,N_5428);
and U7411 (N_7411,N_5463,N_4544);
nand U7412 (N_7412,N_3430,N_4989);
nor U7413 (N_7413,N_5139,N_3938);
and U7414 (N_7414,N_4808,N_4343);
xor U7415 (N_7415,N_4764,N_5979);
and U7416 (N_7416,N_4378,N_4493);
or U7417 (N_7417,N_5559,N_5922);
nand U7418 (N_7418,N_3887,N_3864);
xor U7419 (N_7419,N_4429,N_3722);
nand U7420 (N_7420,N_5591,N_4747);
nand U7421 (N_7421,N_3818,N_3426);
nand U7422 (N_7422,N_3537,N_4549);
nand U7423 (N_7423,N_3859,N_3629);
nand U7424 (N_7424,N_6040,N_3965);
and U7425 (N_7425,N_3631,N_5370);
nand U7426 (N_7426,N_5129,N_5173);
nor U7427 (N_7427,N_4884,N_3161);
xnor U7428 (N_7428,N_4016,N_5703);
or U7429 (N_7429,N_4576,N_5919);
or U7430 (N_7430,N_3501,N_4426);
or U7431 (N_7431,N_3785,N_3373);
nor U7432 (N_7432,N_4746,N_4227);
xor U7433 (N_7433,N_3886,N_4560);
nor U7434 (N_7434,N_6121,N_4354);
or U7435 (N_7435,N_5803,N_3147);
or U7436 (N_7436,N_5323,N_4707);
nor U7437 (N_7437,N_6061,N_4214);
xnor U7438 (N_7438,N_3404,N_4395);
nor U7439 (N_7439,N_3133,N_5831);
nor U7440 (N_7440,N_4490,N_4829);
nor U7441 (N_7441,N_5522,N_5427);
and U7442 (N_7442,N_3643,N_4959);
nand U7443 (N_7443,N_5728,N_6137);
and U7444 (N_7444,N_4894,N_5613);
nor U7445 (N_7445,N_3358,N_5267);
nand U7446 (N_7446,N_5512,N_6233);
xnor U7447 (N_7447,N_5964,N_5111);
nand U7448 (N_7448,N_5766,N_5261);
nor U7449 (N_7449,N_4322,N_4211);
nor U7450 (N_7450,N_5929,N_3560);
and U7451 (N_7451,N_5944,N_5406);
nand U7452 (N_7452,N_6029,N_3228);
nand U7453 (N_7453,N_5666,N_5180);
nor U7454 (N_7454,N_3744,N_5516);
nor U7455 (N_7455,N_6140,N_4824);
or U7456 (N_7456,N_3442,N_5141);
and U7457 (N_7457,N_3340,N_4007);
and U7458 (N_7458,N_5378,N_3997);
nand U7459 (N_7459,N_4008,N_5860);
or U7460 (N_7460,N_4066,N_4298);
and U7461 (N_7461,N_4241,N_5458);
nor U7462 (N_7462,N_4345,N_4213);
nand U7463 (N_7463,N_5545,N_5958);
nor U7464 (N_7464,N_3418,N_5457);
xnor U7465 (N_7465,N_6025,N_4094);
nand U7466 (N_7466,N_3308,N_3595);
and U7467 (N_7467,N_5530,N_4916);
nand U7468 (N_7468,N_5401,N_3812);
and U7469 (N_7469,N_5550,N_3748);
nor U7470 (N_7470,N_4488,N_4032);
or U7471 (N_7471,N_3567,N_3638);
or U7472 (N_7472,N_4087,N_4608);
and U7473 (N_7473,N_3184,N_3527);
or U7474 (N_7474,N_5015,N_4573);
nand U7475 (N_7475,N_5260,N_5236);
nand U7476 (N_7476,N_5618,N_3667);
or U7477 (N_7477,N_5350,N_4765);
nand U7478 (N_7478,N_3539,N_5840);
nand U7479 (N_7479,N_5274,N_3256);
or U7480 (N_7480,N_4496,N_4980);
nand U7481 (N_7481,N_5580,N_3129);
nand U7482 (N_7482,N_5940,N_3891);
or U7483 (N_7483,N_4656,N_4792);
nand U7484 (N_7484,N_5295,N_3838);
nand U7485 (N_7485,N_3144,N_5252);
and U7486 (N_7486,N_5888,N_3932);
and U7487 (N_7487,N_4783,N_3652);
nand U7488 (N_7488,N_4056,N_3282);
nand U7489 (N_7489,N_3332,N_4139);
or U7490 (N_7490,N_4221,N_3683);
nand U7491 (N_7491,N_3469,N_4049);
nor U7492 (N_7492,N_5247,N_4947);
and U7493 (N_7493,N_3660,N_4968);
and U7494 (N_7494,N_3754,N_5005);
xor U7495 (N_7495,N_5715,N_5464);
or U7496 (N_7496,N_5994,N_4716);
and U7497 (N_7497,N_3339,N_5983);
or U7498 (N_7498,N_5177,N_4071);
nor U7499 (N_7499,N_3646,N_5732);
nand U7500 (N_7500,N_3735,N_3362);
or U7501 (N_7501,N_3428,N_4647);
or U7502 (N_7502,N_5734,N_4441);
nand U7503 (N_7503,N_3774,N_4818);
or U7504 (N_7504,N_4209,N_3589);
nor U7505 (N_7505,N_3775,N_6009);
nor U7506 (N_7506,N_5121,N_3526);
nor U7507 (N_7507,N_4200,N_6108);
xnor U7508 (N_7508,N_5536,N_4230);
xnor U7509 (N_7509,N_4299,N_5752);
nand U7510 (N_7510,N_5665,N_4927);
nand U7511 (N_7511,N_5317,N_4415);
nand U7512 (N_7512,N_4239,N_4761);
nor U7513 (N_7513,N_5492,N_3578);
nor U7514 (N_7514,N_4362,N_6127);
nor U7515 (N_7515,N_5918,N_5871);
or U7516 (N_7516,N_3556,N_6135);
or U7517 (N_7517,N_5384,N_6085);
nand U7518 (N_7518,N_5705,N_6101);
and U7519 (N_7519,N_4377,N_5320);
or U7520 (N_7520,N_3714,N_5725);
nand U7521 (N_7521,N_3498,N_5361);
or U7522 (N_7522,N_4484,N_5396);
and U7523 (N_7523,N_3675,N_3743);
or U7524 (N_7524,N_3201,N_5397);
nand U7525 (N_7525,N_4317,N_6034);
or U7526 (N_7526,N_5030,N_3276);
and U7527 (N_7527,N_4303,N_4616);
nand U7528 (N_7528,N_5641,N_6070);
and U7529 (N_7529,N_4551,N_3609);
and U7530 (N_7530,N_5845,N_5836);
and U7531 (N_7531,N_3458,N_4365);
nor U7532 (N_7532,N_5031,N_5963);
nor U7533 (N_7533,N_5771,N_5509);
nand U7534 (N_7534,N_5880,N_5226);
and U7535 (N_7535,N_3395,N_3504);
or U7536 (N_7536,N_3788,N_3533);
nor U7537 (N_7537,N_4917,N_5903);
and U7538 (N_7538,N_6245,N_4099);
and U7539 (N_7539,N_5089,N_5012);
or U7540 (N_7540,N_6067,N_4709);
and U7541 (N_7541,N_3692,N_5253);
nand U7542 (N_7542,N_3835,N_5000);
or U7543 (N_7543,N_3531,N_4237);
and U7544 (N_7544,N_5808,N_4266);
or U7545 (N_7545,N_5717,N_3208);
nor U7546 (N_7546,N_4711,N_5764);
and U7547 (N_7547,N_3773,N_6069);
and U7548 (N_7548,N_3240,N_5908);
nand U7549 (N_7549,N_5467,N_5126);
nor U7550 (N_7550,N_4681,N_5970);
nand U7551 (N_7551,N_5775,N_6215);
or U7552 (N_7552,N_3681,N_3804);
nand U7553 (N_7553,N_3700,N_3842);
nor U7554 (N_7554,N_5729,N_5814);
nand U7555 (N_7555,N_6204,N_4096);
nand U7556 (N_7556,N_5286,N_3753);
or U7557 (N_7557,N_3481,N_3242);
and U7558 (N_7558,N_3734,N_5425);
or U7559 (N_7559,N_4589,N_5155);
and U7560 (N_7560,N_5328,N_4385);
nor U7561 (N_7561,N_4896,N_3262);
nand U7562 (N_7562,N_6166,N_5061);
nand U7563 (N_7563,N_3691,N_6043);
and U7564 (N_7564,N_5508,N_4124);
xnor U7565 (N_7565,N_3624,N_4805);
nor U7566 (N_7566,N_3600,N_4789);
xnor U7567 (N_7567,N_3863,N_4356);
nand U7568 (N_7568,N_4455,N_3858);
nor U7569 (N_7569,N_5901,N_5242);
nand U7570 (N_7570,N_3721,N_5062);
nand U7571 (N_7571,N_5540,N_4467);
nor U7572 (N_7572,N_5678,N_4394);
nand U7573 (N_7573,N_6197,N_3666);
and U7574 (N_7574,N_5801,N_4566);
nand U7575 (N_7575,N_4325,N_5399);
or U7576 (N_7576,N_4559,N_4105);
or U7577 (N_7577,N_5675,N_6159);
nor U7578 (N_7578,N_5684,N_3801);
or U7579 (N_7579,N_3999,N_3908);
nand U7580 (N_7580,N_5063,N_3163);
or U7581 (N_7581,N_4522,N_4289);
xnor U7582 (N_7582,N_5606,N_5683);
nor U7583 (N_7583,N_3507,N_3626);
nand U7584 (N_7584,N_3587,N_5367);
or U7585 (N_7585,N_3846,N_4108);
nor U7586 (N_7586,N_5088,N_5145);
and U7587 (N_7587,N_3292,N_5431);
or U7588 (N_7588,N_3636,N_4024);
nor U7589 (N_7589,N_5292,N_5475);
xor U7590 (N_7590,N_3810,N_5991);
or U7591 (N_7591,N_3449,N_4482);
nor U7592 (N_7592,N_5603,N_5359);
nor U7593 (N_7593,N_3889,N_4206);
and U7594 (N_7594,N_3872,N_5973);
nor U7595 (N_7595,N_4788,N_3170);
nor U7596 (N_7596,N_3855,N_3467);
and U7597 (N_7597,N_3736,N_3664);
or U7598 (N_7598,N_4958,N_4509);
nor U7599 (N_7599,N_4397,N_4939);
and U7600 (N_7600,N_5390,N_3865);
nand U7601 (N_7601,N_4161,N_4791);
nand U7602 (N_7602,N_5074,N_3895);
or U7603 (N_7603,N_4909,N_3337);
nor U7604 (N_7604,N_5565,N_3879);
nand U7605 (N_7605,N_5727,N_6213);
or U7606 (N_7606,N_5777,N_4897);
nor U7607 (N_7607,N_4297,N_5742);
nor U7608 (N_7608,N_5879,N_5120);
and U7609 (N_7609,N_5663,N_5642);
xor U7610 (N_7610,N_5256,N_5975);
nand U7611 (N_7611,N_3179,N_4641);
nor U7612 (N_7612,N_3345,N_4671);
and U7613 (N_7613,N_3393,N_6218);
and U7614 (N_7614,N_5659,N_4021);
and U7615 (N_7615,N_4568,N_3265);
or U7616 (N_7616,N_5806,N_4355);
or U7617 (N_7617,N_5216,N_3461);
nand U7618 (N_7618,N_3955,N_5586);
nand U7619 (N_7619,N_6103,N_3909);
nand U7620 (N_7620,N_5182,N_3361);
nand U7621 (N_7621,N_4002,N_4117);
or U7622 (N_7622,N_6023,N_6188);
or U7623 (N_7623,N_4366,N_3829);
nand U7624 (N_7624,N_4067,N_5639);
nor U7625 (N_7625,N_5038,N_3919);
and U7626 (N_7626,N_5630,N_5205);
nand U7627 (N_7627,N_4089,N_4987);
and U7628 (N_7628,N_5316,N_5454);
and U7629 (N_7629,N_4621,N_6139);
and U7630 (N_7630,N_4047,N_3280);
and U7631 (N_7631,N_5420,N_3127);
or U7632 (N_7632,N_5706,N_5046);
xnor U7633 (N_7633,N_4784,N_4465);
and U7634 (N_7634,N_5810,N_4044);
nor U7635 (N_7635,N_3159,N_4497);
and U7636 (N_7636,N_3851,N_4612);
nand U7637 (N_7637,N_4114,N_3460);
or U7638 (N_7638,N_4081,N_3819);
or U7639 (N_7639,N_3808,N_3601);
nor U7640 (N_7640,N_3745,N_4601);
and U7641 (N_7641,N_4285,N_4657);
nor U7642 (N_7642,N_3324,N_3293);
or U7643 (N_7643,N_5566,N_5324);
xnor U7644 (N_7644,N_4983,N_3869);
or U7645 (N_7645,N_3550,N_3771);
nand U7646 (N_7646,N_5544,N_5547);
nand U7647 (N_7647,N_4706,N_5371);
nor U7648 (N_7648,N_4687,N_4364);
xor U7649 (N_7649,N_4452,N_3464);
xor U7650 (N_7650,N_5581,N_4283);
nor U7651 (N_7651,N_5054,N_4915);
or U7652 (N_7652,N_4570,N_6091);
xnor U7653 (N_7653,N_5419,N_3229);
or U7654 (N_7654,N_3180,N_3772);
nand U7655 (N_7655,N_3383,N_4996);
or U7656 (N_7656,N_3353,N_6071);
xor U7657 (N_7657,N_4849,N_4935);
and U7658 (N_7658,N_5890,N_3263);
or U7659 (N_7659,N_4115,N_6084);
or U7660 (N_7660,N_4995,N_6157);
nand U7661 (N_7661,N_3135,N_4868);
or U7662 (N_7662,N_5006,N_4782);
nor U7663 (N_7663,N_5537,N_4183);
nor U7664 (N_7664,N_3183,N_4940);
nor U7665 (N_7665,N_4969,N_4086);
nand U7666 (N_7666,N_3781,N_3260);
or U7667 (N_7667,N_5682,N_5809);
and U7668 (N_7668,N_3659,N_4836);
nand U7669 (N_7669,N_4770,N_3972);
nand U7670 (N_7670,N_5792,N_5168);
or U7671 (N_7671,N_4771,N_4204);
xor U7672 (N_7672,N_3128,N_3782);
and U7673 (N_7673,N_5265,N_5849);
nor U7674 (N_7674,N_3455,N_5310);
xnor U7675 (N_7675,N_6147,N_5867);
nor U7676 (N_7676,N_5987,N_3559);
nor U7677 (N_7677,N_4584,N_3899);
or U7678 (N_7678,N_5410,N_3446);
or U7679 (N_7679,N_5101,N_4075);
nand U7680 (N_7680,N_3962,N_5368);
and U7681 (N_7681,N_3986,N_4461);
and U7682 (N_7682,N_5380,N_5318);
or U7683 (N_7683,N_4287,N_4625);
and U7684 (N_7684,N_5583,N_3512);
xor U7685 (N_7685,N_3947,N_3350);
and U7686 (N_7686,N_4696,N_4732);
nand U7687 (N_7687,N_5347,N_5844);
nand U7688 (N_7688,N_4665,N_4871);
and U7689 (N_7689,N_3284,N_6096);
and U7690 (N_7690,N_5812,N_6171);
nor U7691 (N_7691,N_3648,N_5854);
nand U7692 (N_7692,N_4257,N_5949);
nor U7693 (N_7693,N_4623,N_5789);
nor U7694 (N_7694,N_3378,N_3605);
or U7695 (N_7695,N_6018,N_5960);
or U7696 (N_7696,N_4201,N_3283);
and U7697 (N_7697,N_3417,N_5003);
and U7698 (N_7698,N_4068,N_4728);
nand U7699 (N_7699,N_3975,N_4168);
nor U7700 (N_7700,N_4269,N_5181);
nor U7701 (N_7701,N_3741,N_4054);
nand U7702 (N_7702,N_4999,N_4278);
nor U7703 (N_7703,N_4466,N_4907);
nand U7704 (N_7704,N_5387,N_3140);
and U7705 (N_7705,N_4173,N_3792);
or U7706 (N_7706,N_3351,N_4416);
or U7707 (N_7707,N_5640,N_5527);
nor U7708 (N_7708,N_4359,N_5243);
nor U7709 (N_7709,N_5628,N_6027);
nand U7710 (N_7710,N_5230,N_4751);
xnor U7711 (N_7711,N_5494,N_3536);
or U7712 (N_7712,N_4674,N_5623);
xnor U7713 (N_7713,N_6162,N_4334);
or U7714 (N_7714,N_5747,N_5548);
nand U7715 (N_7715,N_3806,N_5907);
nand U7716 (N_7716,N_5077,N_3628);
and U7717 (N_7717,N_6192,N_5259);
or U7718 (N_7718,N_3218,N_3713);
nor U7719 (N_7719,N_3239,N_5167);
and U7720 (N_7720,N_3655,N_4472);
xor U7721 (N_7721,N_4304,N_5118);
nand U7722 (N_7722,N_3500,N_3463);
or U7723 (N_7723,N_3725,N_6092);
and U7724 (N_7724,N_3880,N_3317);
nand U7725 (N_7725,N_4389,N_4648);
and U7726 (N_7726,N_4858,N_3579);
and U7727 (N_7727,N_6232,N_5311);
nor U7728 (N_7728,N_5503,N_3758);
nor U7729 (N_7729,N_5383,N_3827);
and U7730 (N_7730,N_4904,N_4444);
and U7731 (N_7731,N_4594,N_4157);
nor U7732 (N_7732,N_3893,N_3212);
xor U7733 (N_7733,N_4526,N_4088);
xor U7734 (N_7734,N_4277,N_4093);
nand U7735 (N_7735,N_5526,N_5953);
or U7736 (N_7736,N_6180,N_4847);
nor U7737 (N_7737,N_5166,N_4491);
or U7738 (N_7738,N_5609,N_6032);
xnor U7739 (N_7739,N_4156,N_6058);
nor U7740 (N_7740,N_6105,N_4181);
nand U7741 (N_7741,N_3379,N_4831);
and U7742 (N_7742,N_3766,N_5284);
or U7743 (N_7743,N_4276,N_5762);
and U7744 (N_7744,N_4037,N_4061);
xnor U7745 (N_7745,N_3797,N_4749);
or U7746 (N_7746,N_5081,N_3677);
and U7747 (N_7747,N_5858,N_5163);
nand U7748 (N_7748,N_6175,N_4593);
and U7749 (N_7749,N_5415,N_3294);
or U7750 (N_7750,N_4703,N_4654);
and U7751 (N_7751,N_5172,N_3482);
nand U7752 (N_7752,N_4942,N_6003);
and U7753 (N_7753,N_6129,N_4107);
xor U7754 (N_7754,N_5576,N_5356);
nand U7755 (N_7755,N_3825,N_6028);
xnor U7756 (N_7756,N_5343,N_3989);
nand U7757 (N_7757,N_5398,N_4025);
nor U7758 (N_7758,N_3789,N_5047);
nand U7759 (N_7759,N_6133,N_5217);
xor U7760 (N_7760,N_4905,N_3286);
nor U7761 (N_7761,N_3415,N_3273);
nand U7762 (N_7762,N_3581,N_3971);
or U7763 (N_7763,N_3568,N_3588);
xor U7764 (N_7764,N_5137,N_6059);
or U7765 (N_7765,N_4833,N_4588);
or U7766 (N_7766,N_5598,N_4074);
nand U7767 (N_7767,N_4133,N_5251);
nor U7768 (N_7768,N_4518,N_3756);
nand U7769 (N_7769,N_5595,N_3453);
and U7770 (N_7770,N_5864,N_3730);
nor U7771 (N_7771,N_5656,N_3385);
nand U7772 (N_7772,N_6004,N_5162);
and U7773 (N_7773,N_4769,N_4041);
and U7774 (N_7774,N_5293,N_3621);
or U7775 (N_7775,N_3923,N_6134);
and U7776 (N_7776,N_4651,N_3951);
xnor U7777 (N_7777,N_5835,N_4288);
and U7778 (N_7778,N_4662,N_5471);
and U7779 (N_7779,N_5156,N_5465);
nor U7780 (N_7780,N_3915,N_3836);
nand U7781 (N_7781,N_5977,N_4357);
nor U7782 (N_7782,N_4520,N_6064);
and U7783 (N_7783,N_5346,N_4439);
xnor U7784 (N_7784,N_5824,N_4590);
nand U7785 (N_7785,N_4561,N_5757);
nand U7786 (N_7786,N_5009,N_4715);
xnor U7787 (N_7787,N_3740,N_4626);
nand U7788 (N_7788,N_3429,N_3432);
and U7789 (N_7789,N_5968,N_5152);
nand U7790 (N_7790,N_3234,N_3335);
or U7791 (N_7791,N_3160,N_4583);
nand U7792 (N_7792,N_4190,N_5984);
nand U7793 (N_7793,N_4815,N_3136);
nor U7794 (N_7794,N_4545,N_4712);
or U7795 (N_7795,N_5333,N_3310);
and U7796 (N_7796,N_5986,N_5702);
nor U7797 (N_7797,N_5748,N_5902);
and U7798 (N_7798,N_4347,N_4949);
nand U7799 (N_7799,N_4113,N_3347);
or U7800 (N_7800,N_3854,N_4456);
and U7801 (N_7801,N_3177,N_3243);
nand U7802 (N_7802,N_5197,N_5407);
nor U7803 (N_7803,N_4832,N_4470);
nor U7804 (N_7804,N_4234,N_3348);
nand U7805 (N_7805,N_3264,N_5164);
nand U7806 (N_7806,N_6224,N_4494);
and U7807 (N_7807,N_3372,N_5413);
and U7808 (N_7808,N_3181,N_4629);
xnor U7809 (N_7809,N_5451,N_5303);
or U7810 (N_7810,N_3826,N_5334);
and U7811 (N_7811,N_4685,N_4307);
and U7812 (N_7812,N_3790,N_5936);
or U7813 (N_7813,N_4489,N_6009);
nand U7814 (N_7814,N_5601,N_3411);
or U7815 (N_7815,N_3476,N_5700);
or U7816 (N_7816,N_5162,N_3183);
nand U7817 (N_7817,N_6002,N_6070);
and U7818 (N_7818,N_5445,N_3188);
nand U7819 (N_7819,N_4599,N_5820);
nand U7820 (N_7820,N_3163,N_4482);
or U7821 (N_7821,N_4192,N_5118);
and U7822 (N_7822,N_5728,N_4816);
nor U7823 (N_7823,N_3871,N_5358);
nor U7824 (N_7824,N_5893,N_5568);
nor U7825 (N_7825,N_3766,N_5919);
nand U7826 (N_7826,N_4149,N_6011);
or U7827 (N_7827,N_5820,N_5586);
or U7828 (N_7828,N_5190,N_4112);
and U7829 (N_7829,N_4688,N_5610);
or U7830 (N_7830,N_4374,N_4684);
and U7831 (N_7831,N_3876,N_5732);
or U7832 (N_7832,N_6158,N_5131);
or U7833 (N_7833,N_4176,N_3429);
and U7834 (N_7834,N_5379,N_6058);
and U7835 (N_7835,N_3449,N_6009);
and U7836 (N_7836,N_5165,N_5318);
or U7837 (N_7837,N_5794,N_6132);
nand U7838 (N_7838,N_5504,N_5010);
or U7839 (N_7839,N_4124,N_5423);
nor U7840 (N_7840,N_3742,N_4932);
and U7841 (N_7841,N_4011,N_5108);
nor U7842 (N_7842,N_5338,N_5074);
and U7843 (N_7843,N_3338,N_5783);
nor U7844 (N_7844,N_3644,N_4836);
nand U7845 (N_7845,N_5435,N_6156);
nor U7846 (N_7846,N_4064,N_4750);
or U7847 (N_7847,N_5626,N_4720);
nor U7848 (N_7848,N_5621,N_4986);
and U7849 (N_7849,N_4648,N_3322);
or U7850 (N_7850,N_4426,N_5727);
or U7851 (N_7851,N_4759,N_5112);
or U7852 (N_7852,N_3907,N_5887);
and U7853 (N_7853,N_3449,N_5167);
or U7854 (N_7854,N_4718,N_3159);
or U7855 (N_7855,N_3932,N_4785);
and U7856 (N_7856,N_4999,N_4270);
nand U7857 (N_7857,N_5340,N_5339);
nand U7858 (N_7858,N_5741,N_5211);
or U7859 (N_7859,N_5922,N_5037);
nand U7860 (N_7860,N_4039,N_3665);
and U7861 (N_7861,N_5202,N_4239);
nand U7862 (N_7862,N_4058,N_3758);
nor U7863 (N_7863,N_3535,N_4280);
nand U7864 (N_7864,N_3407,N_4695);
nand U7865 (N_7865,N_5112,N_5178);
or U7866 (N_7866,N_4587,N_4805);
and U7867 (N_7867,N_3774,N_4785);
nand U7868 (N_7868,N_5117,N_3746);
nand U7869 (N_7869,N_3630,N_5512);
nand U7870 (N_7870,N_4681,N_6124);
xor U7871 (N_7871,N_5542,N_5491);
nand U7872 (N_7872,N_5615,N_4613);
and U7873 (N_7873,N_4622,N_5300);
and U7874 (N_7874,N_4437,N_3918);
and U7875 (N_7875,N_4967,N_5357);
or U7876 (N_7876,N_3192,N_3466);
or U7877 (N_7877,N_4932,N_5396);
or U7878 (N_7878,N_4616,N_4275);
nand U7879 (N_7879,N_3762,N_5906);
nor U7880 (N_7880,N_5712,N_5675);
nor U7881 (N_7881,N_3349,N_4159);
and U7882 (N_7882,N_5284,N_3785);
xor U7883 (N_7883,N_6013,N_3205);
nand U7884 (N_7884,N_5307,N_4607);
or U7885 (N_7885,N_5298,N_3336);
and U7886 (N_7886,N_4809,N_3180);
or U7887 (N_7887,N_4932,N_5243);
or U7888 (N_7888,N_5129,N_3883);
or U7889 (N_7889,N_4455,N_3364);
nor U7890 (N_7890,N_4174,N_4230);
nor U7891 (N_7891,N_5136,N_3454);
nand U7892 (N_7892,N_5173,N_5130);
nor U7893 (N_7893,N_4061,N_3901);
or U7894 (N_7894,N_3474,N_6094);
nor U7895 (N_7895,N_5102,N_3168);
or U7896 (N_7896,N_4472,N_4567);
xor U7897 (N_7897,N_4800,N_5199);
nor U7898 (N_7898,N_4481,N_4755);
or U7899 (N_7899,N_3238,N_4994);
or U7900 (N_7900,N_5443,N_5248);
nor U7901 (N_7901,N_5612,N_3143);
nor U7902 (N_7902,N_4340,N_3427);
and U7903 (N_7903,N_5027,N_4161);
nand U7904 (N_7904,N_5550,N_3908);
and U7905 (N_7905,N_3606,N_4116);
and U7906 (N_7906,N_5154,N_3297);
nand U7907 (N_7907,N_4930,N_4019);
or U7908 (N_7908,N_6130,N_5234);
nor U7909 (N_7909,N_3587,N_4698);
xor U7910 (N_7910,N_6090,N_4672);
xnor U7911 (N_7911,N_3356,N_5330);
or U7912 (N_7912,N_5063,N_4114);
nor U7913 (N_7913,N_5656,N_3351);
and U7914 (N_7914,N_5344,N_4384);
or U7915 (N_7915,N_5765,N_4277);
xnor U7916 (N_7916,N_4102,N_3178);
nor U7917 (N_7917,N_4378,N_4836);
or U7918 (N_7918,N_3793,N_3174);
or U7919 (N_7919,N_6100,N_4180);
or U7920 (N_7920,N_4159,N_5450);
and U7921 (N_7921,N_4083,N_5550);
xnor U7922 (N_7922,N_3282,N_5087);
and U7923 (N_7923,N_4146,N_3912);
and U7924 (N_7924,N_5731,N_4050);
or U7925 (N_7925,N_4815,N_3609);
nor U7926 (N_7926,N_4742,N_5769);
nand U7927 (N_7927,N_4392,N_4909);
and U7928 (N_7928,N_3994,N_5054);
and U7929 (N_7929,N_5509,N_4911);
or U7930 (N_7930,N_5553,N_5567);
nor U7931 (N_7931,N_4523,N_6126);
or U7932 (N_7932,N_5885,N_3247);
nand U7933 (N_7933,N_4624,N_5357);
or U7934 (N_7934,N_5409,N_3153);
nand U7935 (N_7935,N_4027,N_5334);
nor U7936 (N_7936,N_4932,N_4530);
or U7937 (N_7937,N_5077,N_3832);
nor U7938 (N_7938,N_5807,N_5662);
nand U7939 (N_7939,N_4349,N_5665);
nand U7940 (N_7940,N_6149,N_4738);
nor U7941 (N_7941,N_3382,N_3330);
or U7942 (N_7942,N_5140,N_5112);
nand U7943 (N_7943,N_5264,N_6158);
nand U7944 (N_7944,N_5937,N_3998);
or U7945 (N_7945,N_3241,N_4274);
and U7946 (N_7946,N_3904,N_5204);
and U7947 (N_7947,N_6232,N_6089);
nor U7948 (N_7948,N_5597,N_4675);
or U7949 (N_7949,N_3766,N_4715);
nor U7950 (N_7950,N_5757,N_5253);
nor U7951 (N_7951,N_4817,N_5949);
nor U7952 (N_7952,N_5337,N_4694);
and U7953 (N_7953,N_3690,N_3591);
or U7954 (N_7954,N_5138,N_4485);
and U7955 (N_7955,N_4674,N_4223);
or U7956 (N_7956,N_5884,N_5518);
and U7957 (N_7957,N_5924,N_5307);
or U7958 (N_7958,N_4710,N_5835);
or U7959 (N_7959,N_3625,N_3943);
or U7960 (N_7960,N_4634,N_3160);
nand U7961 (N_7961,N_3826,N_3801);
and U7962 (N_7962,N_4712,N_4783);
nor U7963 (N_7963,N_4736,N_3336);
or U7964 (N_7964,N_3948,N_3204);
or U7965 (N_7965,N_5131,N_5539);
nand U7966 (N_7966,N_6195,N_4151);
or U7967 (N_7967,N_5488,N_5062);
and U7968 (N_7968,N_3270,N_5994);
nand U7969 (N_7969,N_5812,N_3191);
and U7970 (N_7970,N_4985,N_5664);
or U7971 (N_7971,N_4766,N_5178);
xnor U7972 (N_7972,N_5908,N_5584);
xor U7973 (N_7973,N_4062,N_5546);
nor U7974 (N_7974,N_5049,N_4578);
nor U7975 (N_7975,N_5919,N_5054);
or U7976 (N_7976,N_4146,N_5302);
or U7977 (N_7977,N_4322,N_5581);
or U7978 (N_7978,N_5248,N_5930);
or U7979 (N_7979,N_3813,N_4356);
xnor U7980 (N_7980,N_4669,N_6016);
nand U7981 (N_7981,N_5861,N_6077);
xnor U7982 (N_7982,N_5233,N_5069);
and U7983 (N_7983,N_5771,N_5197);
nor U7984 (N_7984,N_4657,N_3908);
and U7985 (N_7985,N_6150,N_6003);
or U7986 (N_7986,N_5477,N_5391);
xor U7987 (N_7987,N_3630,N_3660);
and U7988 (N_7988,N_4630,N_5544);
xor U7989 (N_7989,N_6107,N_4959);
nand U7990 (N_7990,N_5760,N_3171);
nor U7991 (N_7991,N_4880,N_4581);
and U7992 (N_7992,N_4137,N_5964);
and U7993 (N_7993,N_4308,N_3728);
and U7994 (N_7994,N_3723,N_5516);
and U7995 (N_7995,N_3785,N_3812);
or U7996 (N_7996,N_3184,N_5783);
nand U7997 (N_7997,N_4911,N_3854);
nand U7998 (N_7998,N_6051,N_3991);
nor U7999 (N_7999,N_5988,N_6011);
or U8000 (N_8000,N_4727,N_3977);
xnor U8001 (N_8001,N_4488,N_4694);
nand U8002 (N_8002,N_4515,N_5201);
nand U8003 (N_8003,N_6162,N_4671);
xnor U8004 (N_8004,N_3814,N_4563);
or U8005 (N_8005,N_4349,N_4400);
or U8006 (N_8006,N_5967,N_3284);
nand U8007 (N_8007,N_6207,N_4344);
or U8008 (N_8008,N_4623,N_4699);
and U8009 (N_8009,N_3941,N_4455);
nand U8010 (N_8010,N_5108,N_4186);
and U8011 (N_8011,N_3684,N_3227);
or U8012 (N_8012,N_3449,N_5296);
and U8013 (N_8013,N_6222,N_5900);
nand U8014 (N_8014,N_5468,N_5640);
nand U8015 (N_8015,N_3885,N_6236);
nor U8016 (N_8016,N_3801,N_5041);
nor U8017 (N_8017,N_4219,N_4627);
nand U8018 (N_8018,N_4645,N_3220);
nand U8019 (N_8019,N_5736,N_4482);
or U8020 (N_8020,N_3604,N_4943);
nand U8021 (N_8021,N_5094,N_3376);
nand U8022 (N_8022,N_5086,N_4353);
or U8023 (N_8023,N_4400,N_5941);
nand U8024 (N_8024,N_5707,N_5964);
and U8025 (N_8025,N_3351,N_3910);
nand U8026 (N_8026,N_3781,N_6038);
or U8027 (N_8027,N_6127,N_5904);
nor U8028 (N_8028,N_3810,N_3633);
nand U8029 (N_8029,N_4413,N_3669);
nand U8030 (N_8030,N_4513,N_5631);
nand U8031 (N_8031,N_3250,N_4729);
and U8032 (N_8032,N_3220,N_3387);
and U8033 (N_8033,N_4114,N_4417);
nor U8034 (N_8034,N_5723,N_6157);
xor U8035 (N_8035,N_5562,N_3972);
and U8036 (N_8036,N_4099,N_4767);
or U8037 (N_8037,N_4358,N_4017);
and U8038 (N_8038,N_5414,N_5543);
nand U8039 (N_8039,N_5573,N_4155);
and U8040 (N_8040,N_3976,N_3885);
nand U8041 (N_8041,N_5578,N_3211);
and U8042 (N_8042,N_3308,N_5924);
or U8043 (N_8043,N_3883,N_3888);
nand U8044 (N_8044,N_3139,N_5228);
and U8045 (N_8045,N_4201,N_5873);
or U8046 (N_8046,N_4367,N_3555);
and U8047 (N_8047,N_5489,N_4675);
or U8048 (N_8048,N_4191,N_4994);
or U8049 (N_8049,N_3249,N_5991);
nand U8050 (N_8050,N_4473,N_4183);
nand U8051 (N_8051,N_4525,N_4716);
nand U8052 (N_8052,N_4828,N_5269);
nor U8053 (N_8053,N_5636,N_5838);
nand U8054 (N_8054,N_4095,N_5017);
xnor U8055 (N_8055,N_5607,N_3211);
and U8056 (N_8056,N_4768,N_5469);
nor U8057 (N_8057,N_5808,N_5409);
nand U8058 (N_8058,N_3455,N_5783);
or U8059 (N_8059,N_3470,N_3466);
and U8060 (N_8060,N_5225,N_5219);
nor U8061 (N_8061,N_3418,N_5100);
and U8062 (N_8062,N_4682,N_4730);
nand U8063 (N_8063,N_3662,N_4059);
and U8064 (N_8064,N_3184,N_4551);
nor U8065 (N_8065,N_4159,N_4275);
nor U8066 (N_8066,N_5650,N_4042);
nand U8067 (N_8067,N_5149,N_5343);
nand U8068 (N_8068,N_4376,N_4503);
nand U8069 (N_8069,N_5136,N_4936);
nor U8070 (N_8070,N_4335,N_5927);
and U8071 (N_8071,N_4933,N_4902);
or U8072 (N_8072,N_5412,N_4944);
or U8073 (N_8073,N_6117,N_5359);
nand U8074 (N_8074,N_5953,N_5015);
nand U8075 (N_8075,N_5679,N_3756);
nand U8076 (N_8076,N_5805,N_5956);
and U8077 (N_8077,N_5989,N_5861);
nand U8078 (N_8078,N_5475,N_5873);
nor U8079 (N_8079,N_3156,N_3841);
xor U8080 (N_8080,N_5839,N_3181);
and U8081 (N_8081,N_3265,N_5387);
nor U8082 (N_8082,N_4104,N_5445);
nor U8083 (N_8083,N_6127,N_3301);
or U8084 (N_8084,N_4504,N_3721);
and U8085 (N_8085,N_5484,N_4142);
nor U8086 (N_8086,N_3200,N_5409);
or U8087 (N_8087,N_6102,N_4303);
nand U8088 (N_8088,N_3604,N_3561);
and U8089 (N_8089,N_3287,N_3496);
nand U8090 (N_8090,N_4831,N_3805);
and U8091 (N_8091,N_5785,N_5413);
nor U8092 (N_8092,N_4058,N_4160);
or U8093 (N_8093,N_4862,N_3208);
or U8094 (N_8094,N_4537,N_3849);
nor U8095 (N_8095,N_5440,N_6109);
nand U8096 (N_8096,N_4986,N_5533);
nor U8097 (N_8097,N_3652,N_5122);
and U8098 (N_8098,N_5523,N_4426);
xnor U8099 (N_8099,N_5720,N_6041);
nand U8100 (N_8100,N_4486,N_4671);
and U8101 (N_8101,N_6152,N_5476);
or U8102 (N_8102,N_6104,N_5714);
nor U8103 (N_8103,N_4812,N_5828);
or U8104 (N_8104,N_4228,N_4978);
nand U8105 (N_8105,N_4986,N_6196);
or U8106 (N_8106,N_5624,N_5336);
and U8107 (N_8107,N_3872,N_5399);
xnor U8108 (N_8108,N_4304,N_3595);
or U8109 (N_8109,N_4706,N_4000);
nand U8110 (N_8110,N_4687,N_5472);
or U8111 (N_8111,N_5788,N_3563);
nand U8112 (N_8112,N_3712,N_4862);
or U8113 (N_8113,N_5130,N_4852);
or U8114 (N_8114,N_5026,N_4939);
xnor U8115 (N_8115,N_5259,N_5993);
nor U8116 (N_8116,N_5765,N_5319);
or U8117 (N_8117,N_5590,N_5899);
or U8118 (N_8118,N_5325,N_3430);
nand U8119 (N_8119,N_3567,N_3860);
and U8120 (N_8120,N_4600,N_4423);
nand U8121 (N_8121,N_5835,N_3364);
or U8122 (N_8122,N_4725,N_5043);
nand U8123 (N_8123,N_4264,N_5897);
and U8124 (N_8124,N_4388,N_3499);
nand U8125 (N_8125,N_4382,N_3917);
nand U8126 (N_8126,N_4550,N_3596);
xor U8127 (N_8127,N_3918,N_4830);
nor U8128 (N_8128,N_3885,N_5854);
nand U8129 (N_8129,N_4591,N_3548);
nor U8130 (N_8130,N_5608,N_4322);
and U8131 (N_8131,N_3173,N_5236);
or U8132 (N_8132,N_3359,N_3939);
and U8133 (N_8133,N_3214,N_4290);
nor U8134 (N_8134,N_4267,N_5927);
nor U8135 (N_8135,N_5598,N_4792);
nand U8136 (N_8136,N_3127,N_5076);
nand U8137 (N_8137,N_6153,N_5387);
xnor U8138 (N_8138,N_3672,N_3898);
and U8139 (N_8139,N_4288,N_5786);
or U8140 (N_8140,N_5187,N_3326);
or U8141 (N_8141,N_6061,N_5875);
and U8142 (N_8142,N_4444,N_5753);
nand U8143 (N_8143,N_3749,N_5217);
nor U8144 (N_8144,N_5050,N_4380);
nor U8145 (N_8145,N_6083,N_3655);
and U8146 (N_8146,N_5981,N_6110);
nand U8147 (N_8147,N_5596,N_4146);
xor U8148 (N_8148,N_5717,N_3354);
or U8149 (N_8149,N_3985,N_3558);
and U8150 (N_8150,N_4555,N_5567);
nand U8151 (N_8151,N_4413,N_4207);
nand U8152 (N_8152,N_4317,N_5171);
and U8153 (N_8153,N_4078,N_5299);
or U8154 (N_8154,N_4620,N_3300);
xnor U8155 (N_8155,N_5349,N_4792);
or U8156 (N_8156,N_4504,N_3363);
nor U8157 (N_8157,N_5267,N_6004);
and U8158 (N_8158,N_5363,N_4793);
xor U8159 (N_8159,N_3499,N_4238);
xnor U8160 (N_8160,N_4238,N_4063);
and U8161 (N_8161,N_4736,N_5417);
nor U8162 (N_8162,N_4646,N_3513);
and U8163 (N_8163,N_4813,N_5318);
xnor U8164 (N_8164,N_6154,N_3472);
nor U8165 (N_8165,N_5115,N_4571);
nand U8166 (N_8166,N_6085,N_5225);
xor U8167 (N_8167,N_6182,N_5150);
or U8168 (N_8168,N_5415,N_4919);
xnor U8169 (N_8169,N_3329,N_3820);
nand U8170 (N_8170,N_6141,N_3287);
nor U8171 (N_8171,N_5409,N_4119);
nand U8172 (N_8172,N_3802,N_5525);
nor U8173 (N_8173,N_5859,N_4595);
nor U8174 (N_8174,N_6080,N_4135);
or U8175 (N_8175,N_6062,N_5714);
or U8176 (N_8176,N_4382,N_5737);
xnor U8177 (N_8177,N_6218,N_5854);
nand U8178 (N_8178,N_5589,N_4038);
or U8179 (N_8179,N_3714,N_3729);
nor U8180 (N_8180,N_3193,N_4656);
and U8181 (N_8181,N_4432,N_5075);
nand U8182 (N_8182,N_5284,N_5152);
nand U8183 (N_8183,N_3725,N_4226);
or U8184 (N_8184,N_5916,N_5976);
and U8185 (N_8185,N_5724,N_3303);
or U8186 (N_8186,N_3754,N_3657);
nor U8187 (N_8187,N_5146,N_5680);
and U8188 (N_8188,N_3616,N_3283);
nand U8189 (N_8189,N_5845,N_3491);
nand U8190 (N_8190,N_5762,N_6131);
nor U8191 (N_8191,N_3806,N_4102);
and U8192 (N_8192,N_4382,N_4725);
nand U8193 (N_8193,N_3623,N_4888);
nor U8194 (N_8194,N_4858,N_5039);
or U8195 (N_8195,N_5417,N_5749);
or U8196 (N_8196,N_4863,N_4037);
or U8197 (N_8197,N_3453,N_3679);
or U8198 (N_8198,N_3968,N_4100);
nand U8199 (N_8199,N_4055,N_5995);
or U8200 (N_8200,N_3843,N_3664);
nand U8201 (N_8201,N_5182,N_6011);
or U8202 (N_8202,N_4724,N_5506);
nand U8203 (N_8203,N_5719,N_4032);
xnor U8204 (N_8204,N_5695,N_4984);
xor U8205 (N_8205,N_5478,N_3878);
and U8206 (N_8206,N_6057,N_4405);
nor U8207 (N_8207,N_4253,N_3582);
nand U8208 (N_8208,N_5720,N_5665);
nor U8209 (N_8209,N_3353,N_5846);
and U8210 (N_8210,N_5665,N_3501);
and U8211 (N_8211,N_5970,N_4880);
nand U8212 (N_8212,N_3582,N_3934);
nor U8213 (N_8213,N_6052,N_4112);
nor U8214 (N_8214,N_3358,N_5089);
and U8215 (N_8215,N_5399,N_4422);
or U8216 (N_8216,N_4352,N_5072);
or U8217 (N_8217,N_5352,N_3155);
nor U8218 (N_8218,N_4422,N_5439);
or U8219 (N_8219,N_4724,N_4218);
or U8220 (N_8220,N_5754,N_3627);
nand U8221 (N_8221,N_3748,N_5826);
or U8222 (N_8222,N_4151,N_4641);
nand U8223 (N_8223,N_3410,N_4332);
and U8224 (N_8224,N_4222,N_6004);
nor U8225 (N_8225,N_3427,N_6032);
and U8226 (N_8226,N_4349,N_3256);
nor U8227 (N_8227,N_4352,N_5677);
and U8228 (N_8228,N_3665,N_3798);
nand U8229 (N_8229,N_5310,N_4607);
nor U8230 (N_8230,N_3472,N_4054);
and U8231 (N_8231,N_4436,N_5125);
or U8232 (N_8232,N_5643,N_5386);
and U8233 (N_8233,N_6080,N_4948);
nand U8234 (N_8234,N_4967,N_3787);
and U8235 (N_8235,N_6221,N_3343);
and U8236 (N_8236,N_4517,N_3225);
nor U8237 (N_8237,N_3690,N_5077);
and U8238 (N_8238,N_5286,N_6204);
or U8239 (N_8239,N_4854,N_3412);
nor U8240 (N_8240,N_3356,N_6222);
xnor U8241 (N_8241,N_5061,N_4539);
xnor U8242 (N_8242,N_4285,N_4709);
or U8243 (N_8243,N_3719,N_4680);
and U8244 (N_8244,N_3938,N_3379);
nand U8245 (N_8245,N_5819,N_5563);
or U8246 (N_8246,N_4435,N_4236);
and U8247 (N_8247,N_4316,N_6049);
or U8248 (N_8248,N_4556,N_4117);
nand U8249 (N_8249,N_5201,N_3659);
nor U8250 (N_8250,N_6208,N_3217);
or U8251 (N_8251,N_4130,N_6087);
nor U8252 (N_8252,N_3537,N_5823);
nor U8253 (N_8253,N_3558,N_3337);
nor U8254 (N_8254,N_3484,N_5281);
nand U8255 (N_8255,N_6085,N_3439);
nor U8256 (N_8256,N_6249,N_5130);
nand U8257 (N_8257,N_3949,N_4970);
or U8258 (N_8258,N_3925,N_6031);
nor U8259 (N_8259,N_3741,N_5208);
nor U8260 (N_8260,N_5817,N_3891);
and U8261 (N_8261,N_5797,N_4788);
and U8262 (N_8262,N_4041,N_5913);
nor U8263 (N_8263,N_5260,N_3373);
nor U8264 (N_8264,N_4656,N_4562);
nor U8265 (N_8265,N_5868,N_5675);
nand U8266 (N_8266,N_5546,N_3255);
nand U8267 (N_8267,N_3568,N_6194);
or U8268 (N_8268,N_4564,N_5107);
nand U8269 (N_8269,N_3671,N_4421);
or U8270 (N_8270,N_4285,N_3633);
or U8271 (N_8271,N_3344,N_4311);
and U8272 (N_8272,N_3748,N_5698);
nand U8273 (N_8273,N_3538,N_3161);
nor U8274 (N_8274,N_4873,N_6009);
nor U8275 (N_8275,N_5746,N_3173);
or U8276 (N_8276,N_6151,N_5057);
nor U8277 (N_8277,N_5570,N_4965);
nor U8278 (N_8278,N_3294,N_5121);
and U8279 (N_8279,N_6230,N_4301);
nor U8280 (N_8280,N_5389,N_4996);
and U8281 (N_8281,N_5352,N_5896);
xnor U8282 (N_8282,N_5677,N_3853);
or U8283 (N_8283,N_3170,N_6172);
or U8284 (N_8284,N_5675,N_3147);
nor U8285 (N_8285,N_5883,N_4915);
nor U8286 (N_8286,N_4521,N_3255);
or U8287 (N_8287,N_3272,N_5432);
or U8288 (N_8288,N_5818,N_4768);
and U8289 (N_8289,N_5191,N_5506);
or U8290 (N_8290,N_3795,N_6063);
xor U8291 (N_8291,N_5503,N_4725);
nor U8292 (N_8292,N_5057,N_4743);
or U8293 (N_8293,N_4326,N_6243);
and U8294 (N_8294,N_5776,N_3825);
nor U8295 (N_8295,N_4146,N_4792);
nand U8296 (N_8296,N_4513,N_5425);
xnor U8297 (N_8297,N_6100,N_5868);
nand U8298 (N_8298,N_5292,N_5870);
or U8299 (N_8299,N_3525,N_5486);
or U8300 (N_8300,N_3385,N_3663);
xor U8301 (N_8301,N_4247,N_6245);
nor U8302 (N_8302,N_5280,N_5422);
nand U8303 (N_8303,N_3908,N_4098);
nand U8304 (N_8304,N_5849,N_3490);
or U8305 (N_8305,N_5941,N_5294);
and U8306 (N_8306,N_3386,N_3399);
nor U8307 (N_8307,N_4780,N_4673);
nor U8308 (N_8308,N_3953,N_3458);
and U8309 (N_8309,N_4288,N_4398);
nor U8310 (N_8310,N_3750,N_5936);
nor U8311 (N_8311,N_3629,N_4353);
or U8312 (N_8312,N_5469,N_5878);
or U8313 (N_8313,N_6178,N_4232);
or U8314 (N_8314,N_6224,N_3167);
nor U8315 (N_8315,N_5096,N_6025);
xor U8316 (N_8316,N_5028,N_6071);
nor U8317 (N_8317,N_4239,N_3644);
nor U8318 (N_8318,N_4964,N_4472);
and U8319 (N_8319,N_4700,N_4568);
or U8320 (N_8320,N_3859,N_4461);
or U8321 (N_8321,N_4353,N_3882);
nor U8322 (N_8322,N_3225,N_4394);
nand U8323 (N_8323,N_5550,N_6134);
or U8324 (N_8324,N_3815,N_5441);
nor U8325 (N_8325,N_4405,N_5144);
nand U8326 (N_8326,N_5487,N_4205);
or U8327 (N_8327,N_5972,N_4279);
nand U8328 (N_8328,N_5758,N_3720);
nor U8329 (N_8329,N_3507,N_3468);
nor U8330 (N_8330,N_5302,N_4251);
and U8331 (N_8331,N_3729,N_4006);
or U8332 (N_8332,N_3398,N_6033);
xnor U8333 (N_8333,N_6005,N_3826);
and U8334 (N_8334,N_3267,N_4624);
xnor U8335 (N_8335,N_4200,N_4949);
and U8336 (N_8336,N_5490,N_4773);
and U8337 (N_8337,N_4883,N_5490);
nand U8338 (N_8338,N_3467,N_5734);
xnor U8339 (N_8339,N_5349,N_5149);
nand U8340 (N_8340,N_4351,N_3272);
or U8341 (N_8341,N_4491,N_4451);
or U8342 (N_8342,N_4145,N_5905);
and U8343 (N_8343,N_5556,N_3710);
xor U8344 (N_8344,N_3773,N_5993);
or U8345 (N_8345,N_6207,N_5342);
nor U8346 (N_8346,N_3916,N_3914);
nor U8347 (N_8347,N_3750,N_3504);
and U8348 (N_8348,N_3690,N_4184);
and U8349 (N_8349,N_3405,N_4758);
and U8350 (N_8350,N_5278,N_5410);
nand U8351 (N_8351,N_4142,N_5738);
nand U8352 (N_8352,N_5591,N_5444);
nor U8353 (N_8353,N_3996,N_5403);
xor U8354 (N_8354,N_3643,N_3729);
nor U8355 (N_8355,N_4139,N_3198);
nand U8356 (N_8356,N_5274,N_4739);
nand U8357 (N_8357,N_5867,N_4730);
or U8358 (N_8358,N_5585,N_3291);
and U8359 (N_8359,N_5476,N_5402);
or U8360 (N_8360,N_5822,N_4246);
or U8361 (N_8361,N_3573,N_3586);
nor U8362 (N_8362,N_4029,N_6226);
and U8363 (N_8363,N_3179,N_5765);
nand U8364 (N_8364,N_4604,N_4199);
nand U8365 (N_8365,N_6006,N_3373);
or U8366 (N_8366,N_3409,N_6222);
xnor U8367 (N_8367,N_3999,N_3601);
xor U8368 (N_8368,N_5950,N_3508);
nand U8369 (N_8369,N_5811,N_4323);
xor U8370 (N_8370,N_4693,N_6226);
nor U8371 (N_8371,N_5425,N_4599);
and U8372 (N_8372,N_3263,N_4097);
nor U8373 (N_8373,N_5073,N_4493);
and U8374 (N_8374,N_3924,N_5385);
nand U8375 (N_8375,N_5979,N_4437);
and U8376 (N_8376,N_5774,N_5744);
nand U8377 (N_8377,N_3233,N_4212);
or U8378 (N_8378,N_5405,N_4254);
nand U8379 (N_8379,N_5229,N_5947);
and U8380 (N_8380,N_5198,N_4436);
nand U8381 (N_8381,N_5315,N_3978);
or U8382 (N_8382,N_4799,N_3190);
xnor U8383 (N_8383,N_5845,N_4340);
or U8384 (N_8384,N_4780,N_4120);
and U8385 (N_8385,N_5116,N_3282);
or U8386 (N_8386,N_4870,N_5177);
nor U8387 (N_8387,N_3659,N_5872);
nor U8388 (N_8388,N_6116,N_5118);
nor U8389 (N_8389,N_4420,N_5633);
xnor U8390 (N_8390,N_4731,N_4069);
xnor U8391 (N_8391,N_3803,N_5903);
nor U8392 (N_8392,N_5506,N_5260);
nor U8393 (N_8393,N_3207,N_5372);
or U8394 (N_8394,N_4318,N_5590);
nand U8395 (N_8395,N_4575,N_3327);
nand U8396 (N_8396,N_5515,N_4746);
or U8397 (N_8397,N_3892,N_5854);
and U8398 (N_8398,N_3564,N_5963);
xnor U8399 (N_8399,N_4638,N_3790);
and U8400 (N_8400,N_5955,N_5444);
and U8401 (N_8401,N_5361,N_5821);
nor U8402 (N_8402,N_3136,N_5407);
or U8403 (N_8403,N_4542,N_3880);
nand U8404 (N_8404,N_3582,N_5674);
and U8405 (N_8405,N_3958,N_5093);
nand U8406 (N_8406,N_6065,N_5751);
xnor U8407 (N_8407,N_3448,N_4562);
nand U8408 (N_8408,N_5819,N_4754);
nor U8409 (N_8409,N_3257,N_5114);
xnor U8410 (N_8410,N_5505,N_5895);
xor U8411 (N_8411,N_3244,N_4169);
xor U8412 (N_8412,N_4025,N_3303);
nor U8413 (N_8413,N_5317,N_5483);
nand U8414 (N_8414,N_3469,N_4996);
nor U8415 (N_8415,N_5374,N_3133);
nor U8416 (N_8416,N_3700,N_3856);
and U8417 (N_8417,N_3763,N_5900);
nand U8418 (N_8418,N_4399,N_3492);
or U8419 (N_8419,N_5607,N_4489);
and U8420 (N_8420,N_3868,N_4908);
or U8421 (N_8421,N_4759,N_4972);
and U8422 (N_8422,N_4751,N_3796);
or U8423 (N_8423,N_3556,N_5335);
and U8424 (N_8424,N_4839,N_5922);
nand U8425 (N_8425,N_4558,N_3341);
nand U8426 (N_8426,N_3322,N_3401);
or U8427 (N_8427,N_4789,N_3544);
and U8428 (N_8428,N_3423,N_4581);
and U8429 (N_8429,N_5685,N_5977);
xor U8430 (N_8430,N_3705,N_5837);
nor U8431 (N_8431,N_4597,N_4057);
nand U8432 (N_8432,N_5552,N_3265);
and U8433 (N_8433,N_5522,N_5794);
xnor U8434 (N_8434,N_4322,N_4306);
xnor U8435 (N_8435,N_5947,N_5181);
and U8436 (N_8436,N_4453,N_3550);
or U8437 (N_8437,N_4176,N_3174);
and U8438 (N_8438,N_3455,N_4996);
and U8439 (N_8439,N_3442,N_3598);
nor U8440 (N_8440,N_3361,N_5949);
nor U8441 (N_8441,N_5707,N_5915);
nand U8442 (N_8442,N_6007,N_5159);
xor U8443 (N_8443,N_3551,N_4870);
or U8444 (N_8444,N_3417,N_4596);
nand U8445 (N_8445,N_3540,N_6148);
and U8446 (N_8446,N_5109,N_4002);
or U8447 (N_8447,N_5884,N_6138);
and U8448 (N_8448,N_3436,N_3963);
and U8449 (N_8449,N_5164,N_3831);
or U8450 (N_8450,N_4380,N_4712);
and U8451 (N_8451,N_4093,N_3263);
and U8452 (N_8452,N_5310,N_4379);
nor U8453 (N_8453,N_6138,N_3774);
nor U8454 (N_8454,N_4185,N_5516);
or U8455 (N_8455,N_5376,N_5047);
nor U8456 (N_8456,N_3770,N_5032);
or U8457 (N_8457,N_3791,N_3166);
nor U8458 (N_8458,N_4699,N_6035);
or U8459 (N_8459,N_6031,N_3370);
nand U8460 (N_8460,N_4050,N_3238);
or U8461 (N_8461,N_4448,N_6205);
nor U8462 (N_8462,N_4093,N_3469);
or U8463 (N_8463,N_5322,N_4773);
or U8464 (N_8464,N_4028,N_4162);
or U8465 (N_8465,N_3457,N_5068);
and U8466 (N_8466,N_4569,N_4589);
and U8467 (N_8467,N_5115,N_4811);
nand U8468 (N_8468,N_3508,N_5122);
and U8469 (N_8469,N_4183,N_5683);
xnor U8470 (N_8470,N_4853,N_6080);
nand U8471 (N_8471,N_5016,N_3520);
nand U8472 (N_8472,N_4294,N_4570);
nand U8473 (N_8473,N_5875,N_3917);
nand U8474 (N_8474,N_3863,N_4031);
xnor U8475 (N_8475,N_4713,N_4964);
nor U8476 (N_8476,N_4551,N_4581);
nand U8477 (N_8477,N_4398,N_3821);
xor U8478 (N_8478,N_3446,N_4524);
nand U8479 (N_8479,N_3545,N_5753);
and U8480 (N_8480,N_5000,N_4230);
nor U8481 (N_8481,N_5105,N_3134);
and U8482 (N_8482,N_3929,N_5586);
or U8483 (N_8483,N_6236,N_5167);
nor U8484 (N_8484,N_3896,N_3324);
and U8485 (N_8485,N_5876,N_5466);
and U8486 (N_8486,N_6245,N_6109);
xor U8487 (N_8487,N_3147,N_5973);
and U8488 (N_8488,N_6205,N_3393);
nand U8489 (N_8489,N_3650,N_6002);
nor U8490 (N_8490,N_4896,N_3370);
nand U8491 (N_8491,N_3211,N_3961);
nand U8492 (N_8492,N_5876,N_3569);
and U8493 (N_8493,N_4836,N_4265);
or U8494 (N_8494,N_6218,N_3700);
or U8495 (N_8495,N_5864,N_4773);
and U8496 (N_8496,N_3169,N_5879);
or U8497 (N_8497,N_4702,N_4992);
nand U8498 (N_8498,N_3340,N_6221);
nor U8499 (N_8499,N_4159,N_4621);
or U8500 (N_8500,N_4046,N_5173);
or U8501 (N_8501,N_6119,N_4521);
or U8502 (N_8502,N_5559,N_3703);
or U8503 (N_8503,N_3325,N_4954);
nor U8504 (N_8504,N_3865,N_4415);
nor U8505 (N_8505,N_5619,N_4758);
nor U8506 (N_8506,N_3859,N_6236);
nor U8507 (N_8507,N_5248,N_4011);
nand U8508 (N_8508,N_5111,N_6019);
and U8509 (N_8509,N_4218,N_3814);
nand U8510 (N_8510,N_5641,N_4216);
and U8511 (N_8511,N_3475,N_4019);
xor U8512 (N_8512,N_3411,N_5082);
or U8513 (N_8513,N_5709,N_4526);
or U8514 (N_8514,N_4274,N_5719);
and U8515 (N_8515,N_3254,N_5340);
nand U8516 (N_8516,N_6247,N_3148);
or U8517 (N_8517,N_3701,N_5881);
or U8518 (N_8518,N_4179,N_4703);
nand U8519 (N_8519,N_3220,N_4407);
or U8520 (N_8520,N_4590,N_3991);
nand U8521 (N_8521,N_4729,N_4655);
xnor U8522 (N_8522,N_5613,N_5445);
and U8523 (N_8523,N_4949,N_3916);
nand U8524 (N_8524,N_6182,N_4854);
xnor U8525 (N_8525,N_3780,N_3785);
and U8526 (N_8526,N_4476,N_6104);
xnor U8527 (N_8527,N_5198,N_3167);
or U8528 (N_8528,N_3830,N_5466);
nand U8529 (N_8529,N_3833,N_3762);
nand U8530 (N_8530,N_5769,N_4806);
and U8531 (N_8531,N_5162,N_4211);
or U8532 (N_8532,N_5441,N_5298);
nor U8533 (N_8533,N_4386,N_4481);
and U8534 (N_8534,N_5841,N_4235);
and U8535 (N_8535,N_3395,N_6177);
nand U8536 (N_8536,N_3847,N_4282);
xnor U8537 (N_8537,N_5779,N_4409);
or U8538 (N_8538,N_5051,N_4244);
nand U8539 (N_8539,N_4526,N_4593);
and U8540 (N_8540,N_5253,N_5282);
nand U8541 (N_8541,N_3848,N_3632);
or U8542 (N_8542,N_4337,N_6012);
and U8543 (N_8543,N_6232,N_4419);
nor U8544 (N_8544,N_4893,N_5886);
and U8545 (N_8545,N_3981,N_4485);
or U8546 (N_8546,N_5257,N_3514);
nor U8547 (N_8547,N_5337,N_3189);
nand U8548 (N_8548,N_4958,N_4327);
nor U8549 (N_8549,N_3796,N_5458);
or U8550 (N_8550,N_4240,N_4344);
and U8551 (N_8551,N_3798,N_4044);
and U8552 (N_8552,N_3180,N_6192);
or U8553 (N_8553,N_4151,N_6219);
xnor U8554 (N_8554,N_5898,N_5455);
nand U8555 (N_8555,N_4753,N_3803);
nand U8556 (N_8556,N_5954,N_6204);
nand U8557 (N_8557,N_4558,N_5142);
and U8558 (N_8558,N_4517,N_5327);
xnor U8559 (N_8559,N_4809,N_5367);
nand U8560 (N_8560,N_6185,N_6081);
and U8561 (N_8561,N_5346,N_3919);
or U8562 (N_8562,N_4570,N_5059);
or U8563 (N_8563,N_5670,N_3299);
and U8564 (N_8564,N_4189,N_4966);
nand U8565 (N_8565,N_3445,N_5751);
or U8566 (N_8566,N_4289,N_3499);
nor U8567 (N_8567,N_4085,N_4912);
xor U8568 (N_8568,N_4793,N_4815);
and U8569 (N_8569,N_4700,N_4286);
or U8570 (N_8570,N_4907,N_6151);
xor U8571 (N_8571,N_4331,N_3576);
or U8572 (N_8572,N_4458,N_4169);
or U8573 (N_8573,N_5064,N_3401);
nor U8574 (N_8574,N_3979,N_3433);
and U8575 (N_8575,N_5842,N_4975);
nand U8576 (N_8576,N_4752,N_5106);
and U8577 (N_8577,N_3936,N_5934);
nor U8578 (N_8578,N_4806,N_5617);
nor U8579 (N_8579,N_3385,N_5319);
or U8580 (N_8580,N_3298,N_6022);
nor U8581 (N_8581,N_5336,N_4231);
or U8582 (N_8582,N_4248,N_5111);
or U8583 (N_8583,N_4965,N_5146);
nand U8584 (N_8584,N_3934,N_4680);
nand U8585 (N_8585,N_3225,N_4386);
nand U8586 (N_8586,N_5494,N_3339);
nand U8587 (N_8587,N_3486,N_6237);
nand U8588 (N_8588,N_4091,N_5394);
xnor U8589 (N_8589,N_6121,N_6143);
and U8590 (N_8590,N_4477,N_5184);
xor U8591 (N_8591,N_4803,N_3256);
nor U8592 (N_8592,N_5493,N_4131);
nor U8593 (N_8593,N_6123,N_3813);
nor U8594 (N_8594,N_4740,N_5006);
nor U8595 (N_8595,N_4413,N_3925);
nand U8596 (N_8596,N_3780,N_3140);
nand U8597 (N_8597,N_3415,N_3873);
nand U8598 (N_8598,N_5262,N_5213);
nand U8599 (N_8599,N_4903,N_4141);
nand U8600 (N_8600,N_4233,N_4235);
or U8601 (N_8601,N_3404,N_3502);
and U8602 (N_8602,N_4017,N_5632);
nand U8603 (N_8603,N_5576,N_5287);
nand U8604 (N_8604,N_3847,N_4611);
nand U8605 (N_8605,N_3244,N_5606);
nor U8606 (N_8606,N_4317,N_6111);
and U8607 (N_8607,N_5374,N_5880);
or U8608 (N_8608,N_5846,N_3916);
and U8609 (N_8609,N_5264,N_3479);
or U8610 (N_8610,N_5976,N_3420);
nand U8611 (N_8611,N_4699,N_3358);
nor U8612 (N_8612,N_3810,N_6126);
nor U8613 (N_8613,N_3962,N_4186);
and U8614 (N_8614,N_3403,N_4582);
nor U8615 (N_8615,N_3514,N_4386);
or U8616 (N_8616,N_3611,N_5848);
nand U8617 (N_8617,N_4748,N_3625);
nor U8618 (N_8618,N_3683,N_4443);
nor U8619 (N_8619,N_4867,N_5067);
and U8620 (N_8620,N_5162,N_4522);
or U8621 (N_8621,N_5003,N_3968);
xor U8622 (N_8622,N_5352,N_4960);
nor U8623 (N_8623,N_3205,N_5191);
or U8624 (N_8624,N_4727,N_5379);
nor U8625 (N_8625,N_3629,N_3510);
nor U8626 (N_8626,N_4941,N_5534);
xor U8627 (N_8627,N_5856,N_5173);
or U8628 (N_8628,N_5171,N_4138);
nand U8629 (N_8629,N_3391,N_5744);
nor U8630 (N_8630,N_3632,N_5373);
or U8631 (N_8631,N_4105,N_3449);
nand U8632 (N_8632,N_3894,N_5982);
or U8633 (N_8633,N_6161,N_5178);
nand U8634 (N_8634,N_4341,N_4635);
nand U8635 (N_8635,N_4248,N_5902);
nor U8636 (N_8636,N_5390,N_5024);
nor U8637 (N_8637,N_5937,N_3754);
and U8638 (N_8638,N_5837,N_4839);
nand U8639 (N_8639,N_5521,N_6180);
nand U8640 (N_8640,N_3381,N_4296);
nor U8641 (N_8641,N_4105,N_4758);
nand U8642 (N_8642,N_4616,N_4052);
or U8643 (N_8643,N_4034,N_4588);
nand U8644 (N_8644,N_4325,N_5858);
and U8645 (N_8645,N_5268,N_3453);
nor U8646 (N_8646,N_5186,N_4740);
and U8647 (N_8647,N_4324,N_3345);
nor U8648 (N_8648,N_4430,N_4643);
nand U8649 (N_8649,N_3303,N_5275);
and U8650 (N_8650,N_4163,N_5800);
nand U8651 (N_8651,N_3800,N_4996);
and U8652 (N_8652,N_4504,N_4228);
nand U8653 (N_8653,N_6114,N_3208);
nor U8654 (N_8654,N_4206,N_4452);
and U8655 (N_8655,N_4477,N_5466);
nor U8656 (N_8656,N_4509,N_5083);
or U8657 (N_8657,N_4083,N_5170);
and U8658 (N_8658,N_4527,N_5523);
nand U8659 (N_8659,N_5129,N_5241);
nand U8660 (N_8660,N_5872,N_5093);
nor U8661 (N_8661,N_4934,N_4203);
and U8662 (N_8662,N_4661,N_4821);
xor U8663 (N_8663,N_5707,N_5262);
nor U8664 (N_8664,N_4658,N_5960);
and U8665 (N_8665,N_4226,N_4238);
and U8666 (N_8666,N_5931,N_4245);
xnor U8667 (N_8667,N_4294,N_4694);
and U8668 (N_8668,N_4239,N_5467);
and U8669 (N_8669,N_3171,N_5454);
xor U8670 (N_8670,N_5833,N_4431);
and U8671 (N_8671,N_5387,N_4812);
nor U8672 (N_8672,N_4701,N_4533);
nand U8673 (N_8673,N_3769,N_4217);
or U8674 (N_8674,N_6180,N_4356);
nor U8675 (N_8675,N_4983,N_5561);
nor U8676 (N_8676,N_5178,N_3564);
nor U8677 (N_8677,N_5236,N_4148);
xor U8678 (N_8678,N_4030,N_3309);
nor U8679 (N_8679,N_5564,N_3365);
and U8680 (N_8680,N_5120,N_3746);
nand U8681 (N_8681,N_5975,N_5009);
nand U8682 (N_8682,N_5311,N_3419);
nand U8683 (N_8683,N_4619,N_6158);
nor U8684 (N_8684,N_3870,N_5739);
xor U8685 (N_8685,N_5462,N_5227);
or U8686 (N_8686,N_3680,N_4469);
nor U8687 (N_8687,N_3584,N_3560);
and U8688 (N_8688,N_5541,N_3429);
or U8689 (N_8689,N_5883,N_4103);
nor U8690 (N_8690,N_4512,N_3307);
nor U8691 (N_8691,N_4218,N_3819);
nand U8692 (N_8692,N_4773,N_4144);
or U8693 (N_8693,N_3536,N_4379);
or U8694 (N_8694,N_6155,N_4705);
nor U8695 (N_8695,N_4228,N_5471);
and U8696 (N_8696,N_3215,N_5414);
or U8697 (N_8697,N_5510,N_4460);
nand U8698 (N_8698,N_3913,N_3572);
and U8699 (N_8699,N_3729,N_3505);
xor U8700 (N_8700,N_3744,N_3916);
and U8701 (N_8701,N_3448,N_6004);
nor U8702 (N_8702,N_3889,N_4229);
or U8703 (N_8703,N_4689,N_3927);
and U8704 (N_8704,N_5954,N_6069);
nor U8705 (N_8705,N_3234,N_5930);
nand U8706 (N_8706,N_3850,N_5533);
or U8707 (N_8707,N_5332,N_4366);
nand U8708 (N_8708,N_3633,N_4290);
nand U8709 (N_8709,N_5902,N_5635);
or U8710 (N_8710,N_3839,N_3292);
xor U8711 (N_8711,N_3439,N_4137);
or U8712 (N_8712,N_6229,N_5195);
and U8713 (N_8713,N_5741,N_6018);
nand U8714 (N_8714,N_5304,N_4023);
xor U8715 (N_8715,N_4686,N_5637);
or U8716 (N_8716,N_3578,N_5816);
and U8717 (N_8717,N_3315,N_4656);
and U8718 (N_8718,N_4303,N_5064);
nor U8719 (N_8719,N_5714,N_5034);
and U8720 (N_8720,N_5996,N_3354);
and U8721 (N_8721,N_4162,N_4423);
or U8722 (N_8722,N_3649,N_4383);
nand U8723 (N_8723,N_3803,N_4901);
xor U8724 (N_8724,N_5642,N_4490);
or U8725 (N_8725,N_4361,N_5849);
and U8726 (N_8726,N_5503,N_4286);
nand U8727 (N_8727,N_4674,N_4559);
or U8728 (N_8728,N_4606,N_4350);
nor U8729 (N_8729,N_4355,N_5648);
xnor U8730 (N_8730,N_4235,N_6075);
nand U8731 (N_8731,N_4346,N_4886);
nor U8732 (N_8732,N_4489,N_5692);
nor U8733 (N_8733,N_4892,N_3445);
or U8734 (N_8734,N_5684,N_6120);
nand U8735 (N_8735,N_5488,N_3797);
or U8736 (N_8736,N_5355,N_3337);
or U8737 (N_8737,N_3936,N_5362);
nand U8738 (N_8738,N_4389,N_4808);
and U8739 (N_8739,N_5136,N_3265);
nor U8740 (N_8740,N_4914,N_4031);
or U8741 (N_8741,N_5226,N_5969);
nand U8742 (N_8742,N_3173,N_4668);
or U8743 (N_8743,N_3929,N_3263);
and U8744 (N_8744,N_5115,N_3423);
xnor U8745 (N_8745,N_6206,N_4443);
nor U8746 (N_8746,N_5316,N_4739);
and U8747 (N_8747,N_5715,N_6122);
or U8748 (N_8748,N_5537,N_5258);
or U8749 (N_8749,N_4421,N_6121);
or U8750 (N_8750,N_4956,N_3817);
nand U8751 (N_8751,N_6114,N_5824);
or U8752 (N_8752,N_4505,N_5705);
and U8753 (N_8753,N_4867,N_3862);
nor U8754 (N_8754,N_4816,N_6029);
or U8755 (N_8755,N_4807,N_3140);
or U8756 (N_8756,N_4352,N_5752);
and U8757 (N_8757,N_3183,N_3810);
or U8758 (N_8758,N_3656,N_5611);
and U8759 (N_8759,N_5750,N_5345);
xnor U8760 (N_8760,N_3254,N_6218);
or U8761 (N_8761,N_3580,N_4383);
or U8762 (N_8762,N_4048,N_3273);
or U8763 (N_8763,N_3619,N_4539);
nor U8764 (N_8764,N_4086,N_4117);
or U8765 (N_8765,N_4542,N_5306);
nor U8766 (N_8766,N_4657,N_4957);
nor U8767 (N_8767,N_3825,N_4768);
xnor U8768 (N_8768,N_3510,N_5304);
nor U8769 (N_8769,N_4412,N_3949);
nand U8770 (N_8770,N_3272,N_5450);
nand U8771 (N_8771,N_5953,N_5441);
and U8772 (N_8772,N_5607,N_3716);
nand U8773 (N_8773,N_3308,N_3893);
xnor U8774 (N_8774,N_3810,N_3913);
nand U8775 (N_8775,N_5675,N_3561);
nand U8776 (N_8776,N_3278,N_5271);
nand U8777 (N_8777,N_5821,N_3598);
nor U8778 (N_8778,N_4553,N_6186);
or U8779 (N_8779,N_3392,N_3461);
nor U8780 (N_8780,N_6224,N_5724);
nor U8781 (N_8781,N_3175,N_4587);
or U8782 (N_8782,N_3779,N_3962);
nor U8783 (N_8783,N_4958,N_5119);
nor U8784 (N_8784,N_3960,N_3860);
xnor U8785 (N_8785,N_5184,N_5394);
or U8786 (N_8786,N_3317,N_3293);
nor U8787 (N_8787,N_4027,N_5817);
or U8788 (N_8788,N_4310,N_5889);
nor U8789 (N_8789,N_4959,N_3199);
nand U8790 (N_8790,N_4171,N_4813);
nand U8791 (N_8791,N_3388,N_3667);
nor U8792 (N_8792,N_4294,N_6103);
or U8793 (N_8793,N_4075,N_5428);
nand U8794 (N_8794,N_4154,N_4484);
nor U8795 (N_8795,N_3741,N_5898);
and U8796 (N_8796,N_5196,N_5685);
nor U8797 (N_8797,N_4905,N_4553);
nand U8798 (N_8798,N_3270,N_6175);
or U8799 (N_8799,N_3304,N_4338);
nand U8800 (N_8800,N_3574,N_6146);
and U8801 (N_8801,N_3458,N_4891);
nor U8802 (N_8802,N_4230,N_4965);
or U8803 (N_8803,N_5408,N_4746);
and U8804 (N_8804,N_4715,N_3768);
nor U8805 (N_8805,N_5010,N_4398);
nor U8806 (N_8806,N_3908,N_5116);
xor U8807 (N_8807,N_3297,N_4305);
nor U8808 (N_8808,N_5164,N_4651);
or U8809 (N_8809,N_3472,N_4669);
or U8810 (N_8810,N_3603,N_5172);
nor U8811 (N_8811,N_4550,N_4051);
nand U8812 (N_8812,N_5329,N_5231);
and U8813 (N_8813,N_3182,N_3155);
and U8814 (N_8814,N_4317,N_5230);
and U8815 (N_8815,N_5060,N_4056);
or U8816 (N_8816,N_4691,N_4814);
nor U8817 (N_8817,N_4172,N_5623);
and U8818 (N_8818,N_5390,N_4074);
nor U8819 (N_8819,N_3748,N_3681);
or U8820 (N_8820,N_3873,N_3741);
and U8821 (N_8821,N_5946,N_3884);
or U8822 (N_8822,N_5994,N_3756);
nand U8823 (N_8823,N_5303,N_5154);
or U8824 (N_8824,N_4911,N_5383);
xnor U8825 (N_8825,N_5945,N_4629);
and U8826 (N_8826,N_4283,N_4335);
and U8827 (N_8827,N_3691,N_3829);
and U8828 (N_8828,N_5621,N_5094);
nor U8829 (N_8829,N_5187,N_3403);
nand U8830 (N_8830,N_4516,N_4000);
and U8831 (N_8831,N_5510,N_5192);
and U8832 (N_8832,N_5448,N_4308);
or U8833 (N_8833,N_5213,N_4944);
and U8834 (N_8834,N_5413,N_5460);
nor U8835 (N_8835,N_6083,N_3912);
nor U8836 (N_8836,N_3912,N_4152);
or U8837 (N_8837,N_3923,N_3659);
nor U8838 (N_8838,N_5491,N_5577);
or U8839 (N_8839,N_5571,N_5483);
xor U8840 (N_8840,N_3297,N_5195);
or U8841 (N_8841,N_3390,N_3845);
or U8842 (N_8842,N_4598,N_4313);
or U8843 (N_8843,N_4242,N_3793);
xor U8844 (N_8844,N_3812,N_4571);
nor U8845 (N_8845,N_3159,N_3201);
nor U8846 (N_8846,N_5336,N_5055);
nand U8847 (N_8847,N_4471,N_5129);
nand U8848 (N_8848,N_5128,N_6073);
nor U8849 (N_8849,N_3211,N_4076);
and U8850 (N_8850,N_5675,N_4460);
nand U8851 (N_8851,N_3258,N_4193);
or U8852 (N_8852,N_3530,N_5094);
and U8853 (N_8853,N_3298,N_4059);
nor U8854 (N_8854,N_4343,N_4649);
nand U8855 (N_8855,N_3703,N_5196);
nor U8856 (N_8856,N_5611,N_3522);
nand U8857 (N_8857,N_4904,N_4883);
nand U8858 (N_8858,N_6169,N_4359);
and U8859 (N_8859,N_5417,N_5323);
nor U8860 (N_8860,N_4205,N_5170);
nand U8861 (N_8861,N_4275,N_5856);
and U8862 (N_8862,N_4800,N_5935);
xnor U8863 (N_8863,N_3174,N_5632);
xnor U8864 (N_8864,N_5374,N_4671);
nand U8865 (N_8865,N_6140,N_5910);
nand U8866 (N_8866,N_4213,N_5587);
nand U8867 (N_8867,N_5669,N_4794);
nor U8868 (N_8868,N_3593,N_3545);
or U8869 (N_8869,N_6206,N_4369);
and U8870 (N_8870,N_3715,N_6135);
or U8871 (N_8871,N_3445,N_4710);
xor U8872 (N_8872,N_5332,N_4833);
nor U8873 (N_8873,N_4625,N_4879);
or U8874 (N_8874,N_5192,N_3508);
or U8875 (N_8875,N_4748,N_5258);
nor U8876 (N_8876,N_4275,N_4098);
nor U8877 (N_8877,N_5707,N_4471);
or U8878 (N_8878,N_4790,N_3552);
nor U8879 (N_8879,N_6139,N_5288);
xnor U8880 (N_8880,N_4179,N_4849);
nor U8881 (N_8881,N_3991,N_3194);
and U8882 (N_8882,N_5205,N_4690);
nand U8883 (N_8883,N_5697,N_3703);
and U8884 (N_8884,N_3982,N_3465);
nor U8885 (N_8885,N_4244,N_4378);
and U8886 (N_8886,N_5096,N_5160);
and U8887 (N_8887,N_3301,N_5000);
or U8888 (N_8888,N_3126,N_4467);
nand U8889 (N_8889,N_4192,N_5713);
nand U8890 (N_8890,N_4632,N_6166);
nand U8891 (N_8891,N_4998,N_3444);
xor U8892 (N_8892,N_3791,N_5698);
nand U8893 (N_8893,N_6096,N_3410);
or U8894 (N_8894,N_5448,N_6046);
nor U8895 (N_8895,N_5662,N_5637);
nand U8896 (N_8896,N_6114,N_6097);
and U8897 (N_8897,N_4839,N_4503);
nand U8898 (N_8898,N_5237,N_4272);
and U8899 (N_8899,N_4050,N_6041);
xnor U8900 (N_8900,N_6081,N_4076);
and U8901 (N_8901,N_5869,N_5732);
or U8902 (N_8902,N_3547,N_3142);
and U8903 (N_8903,N_6148,N_5096);
and U8904 (N_8904,N_4962,N_3785);
nor U8905 (N_8905,N_3353,N_4347);
or U8906 (N_8906,N_3253,N_6144);
and U8907 (N_8907,N_4199,N_4139);
nand U8908 (N_8908,N_3845,N_5192);
nand U8909 (N_8909,N_3509,N_5954);
nor U8910 (N_8910,N_5097,N_6166);
or U8911 (N_8911,N_3747,N_3206);
or U8912 (N_8912,N_3617,N_6048);
xor U8913 (N_8913,N_4709,N_5000);
and U8914 (N_8914,N_5959,N_3986);
nand U8915 (N_8915,N_5434,N_3721);
nand U8916 (N_8916,N_4082,N_5703);
xor U8917 (N_8917,N_5459,N_4402);
nor U8918 (N_8918,N_5288,N_3541);
nand U8919 (N_8919,N_3193,N_4574);
nand U8920 (N_8920,N_5165,N_4303);
and U8921 (N_8921,N_5822,N_5937);
and U8922 (N_8922,N_5939,N_5444);
or U8923 (N_8923,N_3553,N_3425);
or U8924 (N_8924,N_4552,N_3713);
nand U8925 (N_8925,N_4872,N_3956);
or U8926 (N_8926,N_3534,N_4109);
nand U8927 (N_8927,N_5566,N_4742);
and U8928 (N_8928,N_4447,N_5625);
and U8929 (N_8929,N_3321,N_3343);
or U8930 (N_8930,N_4707,N_6164);
nor U8931 (N_8931,N_4108,N_3867);
nor U8932 (N_8932,N_5743,N_4981);
nor U8933 (N_8933,N_4678,N_6042);
or U8934 (N_8934,N_5229,N_4724);
nand U8935 (N_8935,N_6049,N_3635);
nand U8936 (N_8936,N_6141,N_4708);
or U8937 (N_8937,N_5190,N_5164);
and U8938 (N_8938,N_6187,N_4349);
or U8939 (N_8939,N_5320,N_4469);
nand U8940 (N_8940,N_4887,N_3530);
xor U8941 (N_8941,N_5157,N_5091);
nand U8942 (N_8942,N_3260,N_3183);
and U8943 (N_8943,N_3878,N_5196);
and U8944 (N_8944,N_5964,N_3177);
nor U8945 (N_8945,N_3664,N_3927);
nor U8946 (N_8946,N_3928,N_5401);
nor U8947 (N_8947,N_4146,N_3848);
nor U8948 (N_8948,N_4768,N_3606);
or U8949 (N_8949,N_5768,N_3686);
xor U8950 (N_8950,N_4758,N_5454);
or U8951 (N_8951,N_3886,N_5949);
xor U8952 (N_8952,N_4527,N_4967);
or U8953 (N_8953,N_4256,N_4371);
nand U8954 (N_8954,N_5189,N_3358);
nand U8955 (N_8955,N_3292,N_4013);
nor U8956 (N_8956,N_3271,N_3888);
nor U8957 (N_8957,N_4243,N_3362);
or U8958 (N_8958,N_5911,N_5146);
or U8959 (N_8959,N_5055,N_3579);
or U8960 (N_8960,N_3675,N_4745);
or U8961 (N_8961,N_4410,N_5558);
nor U8962 (N_8962,N_3572,N_6062);
nor U8963 (N_8963,N_3320,N_4615);
nor U8964 (N_8964,N_4270,N_5271);
and U8965 (N_8965,N_5819,N_6247);
nor U8966 (N_8966,N_3882,N_5981);
nand U8967 (N_8967,N_4665,N_3333);
xor U8968 (N_8968,N_5375,N_3850);
and U8969 (N_8969,N_3794,N_5002);
nand U8970 (N_8970,N_5191,N_4932);
nor U8971 (N_8971,N_3780,N_3265);
and U8972 (N_8972,N_3768,N_4922);
nand U8973 (N_8973,N_6183,N_3955);
nor U8974 (N_8974,N_5948,N_4290);
nand U8975 (N_8975,N_4724,N_5804);
nand U8976 (N_8976,N_5129,N_5046);
and U8977 (N_8977,N_3126,N_5543);
or U8978 (N_8978,N_4886,N_5685);
or U8979 (N_8979,N_4148,N_4969);
xor U8980 (N_8980,N_5204,N_3395);
and U8981 (N_8981,N_5206,N_5786);
nor U8982 (N_8982,N_5030,N_5958);
nand U8983 (N_8983,N_4389,N_5692);
or U8984 (N_8984,N_5854,N_4661);
and U8985 (N_8985,N_5173,N_6002);
nand U8986 (N_8986,N_3876,N_3472);
and U8987 (N_8987,N_3880,N_3622);
nand U8988 (N_8988,N_4233,N_5368);
nand U8989 (N_8989,N_4835,N_4739);
or U8990 (N_8990,N_3883,N_4323);
xor U8991 (N_8991,N_3652,N_5542);
and U8992 (N_8992,N_3940,N_4128);
nor U8993 (N_8993,N_3203,N_3661);
xnor U8994 (N_8994,N_4387,N_3434);
and U8995 (N_8995,N_5745,N_4547);
nor U8996 (N_8996,N_5685,N_3152);
nand U8997 (N_8997,N_5987,N_3823);
nor U8998 (N_8998,N_3349,N_6148);
nand U8999 (N_8999,N_4990,N_6028);
or U9000 (N_9000,N_3686,N_6216);
and U9001 (N_9001,N_5503,N_5083);
and U9002 (N_9002,N_5447,N_5707);
xor U9003 (N_9003,N_5163,N_5547);
or U9004 (N_9004,N_4825,N_3245);
nand U9005 (N_9005,N_5308,N_4760);
nand U9006 (N_9006,N_3759,N_5903);
or U9007 (N_9007,N_4834,N_6098);
nor U9008 (N_9008,N_4086,N_5854);
nor U9009 (N_9009,N_5693,N_6042);
nand U9010 (N_9010,N_3470,N_4602);
and U9011 (N_9011,N_4951,N_5339);
and U9012 (N_9012,N_5776,N_4007);
xor U9013 (N_9013,N_4241,N_4743);
or U9014 (N_9014,N_5694,N_5097);
and U9015 (N_9015,N_3633,N_3202);
xnor U9016 (N_9016,N_3450,N_3157);
nand U9017 (N_9017,N_3996,N_4180);
or U9018 (N_9018,N_3585,N_4205);
nor U9019 (N_9019,N_6014,N_3970);
nand U9020 (N_9020,N_4784,N_4827);
or U9021 (N_9021,N_4881,N_3820);
nand U9022 (N_9022,N_5071,N_5973);
or U9023 (N_9023,N_6041,N_3509);
xnor U9024 (N_9024,N_4362,N_5224);
and U9025 (N_9025,N_4264,N_5891);
nand U9026 (N_9026,N_3758,N_6192);
and U9027 (N_9027,N_5986,N_6061);
nor U9028 (N_9028,N_3310,N_5539);
xnor U9029 (N_9029,N_3570,N_4229);
nand U9030 (N_9030,N_4638,N_5654);
nand U9031 (N_9031,N_3574,N_6224);
or U9032 (N_9032,N_5827,N_4334);
nand U9033 (N_9033,N_4795,N_3317);
nor U9034 (N_9034,N_4643,N_5731);
or U9035 (N_9035,N_4022,N_5294);
xor U9036 (N_9036,N_4816,N_3649);
xnor U9037 (N_9037,N_3190,N_5975);
nor U9038 (N_9038,N_5542,N_4023);
nand U9039 (N_9039,N_6131,N_5560);
and U9040 (N_9040,N_4589,N_5727);
or U9041 (N_9041,N_4295,N_4046);
nand U9042 (N_9042,N_3843,N_3373);
and U9043 (N_9043,N_4026,N_3942);
nand U9044 (N_9044,N_5886,N_4543);
and U9045 (N_9045,N_4821,N_4524);
or U9046 (N_9046,N_5517,N_5132);
nor U9047 (N_9047,N_4041,N_3875);
and U9048 (N_9048,N_4026,N_3946);
nand U9049 (N_9049,N_5987,N_4335);
and U9050 (N_9050,N_5353,N_3772);
and U9051 (N_9051,N_3837,N_3871);
and U9052 (N_9052,N_4495,N_6165);
nand U9053 (N_9053,N_3866,N_5420);
nand U9054 (N_9054,N_4381,N_5696);
nand U9055 (N_9055,N_3233,N_4251);
nand U9056 (N_9056,N_6146,N_4586);
or U9057 (N_9057,N_5261,N_4511);
and U9058 (N_9058,N_3205,N_5179);
and U9059 (N_9059,N_6214,N_5525);
xnor U9060 (N_9060,N_5361,N_4057);
and U9061 (N_9061,N_3649,N_4525);
xnor U9062 (N_9062,N_5929,N_4126);
or U9063 (N_9063,N_3843,N_4081);
or U9064 (N_9064,N_6140,N_5781);
nand U9065 (N_9065,N_3341,N_3167);
and U9066 (N_9066,N_5462,N_3322);
or U9067 (N_9067,N_4350,N_4897);
nor U9068 (N_9068,N_4110,N_4556);
nand U9069 (N_9069,N_4414,N_3433);
and U9070 (N_9070,N_4000,N_3723);
xor U9071 (N_9071,N_3534,N_5979);
nand U9072 (N_9072,N_4585,N_4841);
or U9073 (N_9073,N_5668,N_5276);
nor U9074 (N_9074,N_4861,N_3198);
and U9075 (N_9075,N_5250,N_3407);
nor U9076 (N_9076,N_4739,N_5386);
and U9077 (N_9077,N_3973,N_5331);
nor U9078 (N_9078,N_4099,N_4076);
or U9079 (N_9079,N_3371,N_5424);
nor U9080 (N_9080,N_3890,N_4376);
nor U9081 (N_9081,N_5410,N_3469);
nor U9082 (N_9082,N_4802,N_5376);
or U9083 (N_9083,N_3307,N_5066);
nor U9084 (N_9084,N_5339,N_3728);
nor U9085 (N_9085,N_4666,N_5557);
and U9086 (N_9086,N_5904,N_3661);
and U9087 (N_9087,N_5643,N_4212);
or U9088 (N_9088,N_4730,N_5530);
xnor U9089 (N_9089,N_4611,N_3748);
xor U9090 (N_9090,N_6084,N_5121);
nand U9091 (N_9091,N_4520,N_6144);
nor U9092 (N_9092,N_3981,N_5222);
xnor U9093 (N_9093,N_5701,N_5405);
nand U9094 (N_9094,N_4377,N_3723);
or U9095 (N_9095,N_4803,N_3262);
xnor U9096 (N_9096,N_3472,N_3369);
nand U9097 (N_9097,N_4899,N_3716);
nand U9098 (N_9098,N_5293,N_4179);
or U9099 (N_9099,N_5329,N_5159);
or U9100 (N_9100,N_5943,N_4118);
nand U9101 (N_9101,N_6040,N_3505);
nor U9102 (N_9102,N_6172,N_4405);
or U9103 (N_9103,N_4451,N_3786);
xor U9104 (N_9104,N_4875,N_5299);
and U9105 (N_9105,N_4493,N_3777);
nor U9106 (N_9106,N_5658,N_3889);
nand U9107 (N_9107,N_5949,N_3884);
xnor U9108 (N_9108,N_6021,N_4319);
nand U9109 (N_9109,N_5151,N_5999);
xnor U9110 (N_9110,N_5929,N_4330);
nand U9111 (N_9111,N_5842,N_4780);
and U9112 (N_9112,N_3321,N_4502);
and U9113 (N_9113,N_5779,N_3581);
nand U9114 (N_9114,N_4622,N_5839);
nand U9115 (N_9115,N_4240,N_3226);
nand U9116 (N_9116,N_3929,N_4366);
and U9117 (N_9117,N_4045,N_5458);
nand U9118 (N_9118,N_3801,N_3934);
and U9119 (N_9119,N_5064,N_3219);
or U9120 (N_9120,N_3803,N_4609);
nand U9121 (N_9121,N_5032,N_6139);
and U9122 (N_9122,N_4686,N_5098);
or U9123 (N_9123,N_4162,N_4621);
nor U9124 (N_9124,N_4836,N_3544);
nor U9125 (N_9125,N_5250,N_4206);
nand U9126 (N_9126,N_5400,N_3144);
nor U9127 (N_9127,N_3841,N_4177);
xnor U9128 (N_9128,N_4837,N_3172);
nand U9129 (N_9129,N_6032,N_3356);
nor U9130 (N_9130,N_5691,N_5273);
and U9131 (N_9131,N_4292,N_4545);
xnor U9132 (N_9132,N_4652,N_6117);
nand U9133 (N_9133,N_4491,N_4764);
nor U9134 (N_9134,N_3827,N_3286);
or U9135 (N_9135,N_3722,N_4242);
or U9136 (N_9136,N_5527,N_4873);
or U9137 (N_9137,N_5767,N_3498);
or U9138 (N_9138,N_5502,N_5349);
nor U9139 (N_9139,N_3563,N_5708);
nand U9140 (N_9140,N_4552,N_4881);
nand U9141 (N_9141,N_5359,N_3459);
or U9142 (N_9142,N_4362,N_3140);
nor U9143 (N_9143,N_5148,N_3439);
nor U9144 (N_9144,N_5771,N_4151);
and U9145 (N_9145,N_3185,N_4110);
nor U9146 (N_9146,N_5749,N_3706);
nand U9147 (N_9147,N_5489,N_5828);
and U9148 (N_9148,N_4495,N_4301);
nor U9149 (N_9149,N_4590,N_4469);
xor U9150 (N_9150,N_5183,N_3555);
and U9151 (N_9151,N_4374,N_5324);
or U9152 (N_9152,N_4890,N_3831);
nor U9153 (N_9153,N_5501,N_5199);
and U9154 (N_9154,N_4909,N_3851);
or U9155 (N_9155,N_6249,N_4192);
nand U9156 (N_9156,N_6018,N_5608);
nor U9157 (N_9157,N_3398,N_6064);
nand U9158 (N_9158,N_5590,N_4075);
nand U9159 (N_9159,N_3648,N_6142);
and U9160 (N_9160,N_3767,N_4358);
nand U9161 (N_9161,N_6116,N_3417);
and U9162 (N_9162,N_3742,N_5629);
xor U9163 (N_9163,N_4817,N_5161);
or U9164 (N_9164,N_5234,N_5876);
and U9165 (N_9165,N_4062,N_3429);
nand U9166 (N_9166,N_6168,N_5576);
and U9167 (N_9167,N_5188,N_3689);
and U9168 (N_9168,N_3939,N_3433);
xnor U9169 (N_9169,N_5470,N_6137);
nor U9170 (N_9170,N_5764,N_4814);
nor U9171 (N_9171,N_4521,N_4345);
or U9172 (N_9172,N_5351,N_5377);
nor U9173 (N_9173,N_4198,N_3720);
and U9174 (N_9174,N_5750,N_3932);
and U9175 (N_9175,N_5913,N_4555);
or U9176 (N_9176,N_5961,N_4215);
nand U9177 (N_9177,N_3163,N_4611);
and U9178 (N_9178,N_3526,N_5689);
nand U9179 (N_9179,N_5459,N_3314);
nand U9180 (N_9180,N_6249,N_3164);
nand U9181 (N_9181,N_5618,N_3587);
xor U9182 (N_9182,N_5311,N_5110);
or U9183 (N_9183,N_5868,N_3919);
nand U9184 (N_9184,N_6103,N_3230);
nand U9185 (N_9185,N_4101,N_5660);
and U9186 (N_9186,N_3371,N_4105);
or U9187 (N_9187,N_4627,N_3133);
nor U9188 (N_9188,N_4980,N_5328);
nor U9189 (N_9189,N_4704,N_5992);
nand U9190 (N_9190,N_4455,N_5506);
nor U9191 (N_9191,N_4708,N_3549);
nor U9192 (N_9192,N_3139,N_3977);
nor U9193 (N_9193,N_4749,N_5171);
nand U9194 (N_9194,N_5733,N_4068);
and U9195 (N_9195,N_5434,N_5425);
nor U9196 (N_9196,N_3215,N_5255);
xnor U9197 (N_9197,N_3439,N_3893);
nor U9198 (N_9198,N_3913,N_4907);
and U9199 (N_9199,N_5710,N_3949);
and U9200 (N_9200,N_5884,N_4868);
nand U9201 (N_9201,N_3987,N_4712);
and U9202 (N_9202,N_5973,N_5612);
and U9203 (N_9203,N_3760,N_4607);
and U9204 (N_9204,N_4064,N_6079);
xor U9205 (N_9205,N_5184,N_6149);
nor U9206 (N_9206,N_5738,N_4837);
nand U9207 (N_9207,N_4261,N_3866);
or U9208 (N_9208,N_5154,N_5928);
nor U9209 (N_9209,N_3535,N_4014);
nand U9210 (N_9210,N_5806,N_4158);
nand U9211 (N_9211,N_4340,N_4494);
nand U9212 (N_9212,N_4808,N_4269);
or U9213 (N_9213,N_4973,N_4512);
and U9214 (N_9214,N_3689,N_5472);
nor U9215 (N_9215,N_4541,N_5497);
and U9216 (N_9216,N_4781,N_6063);
nor U9217 (N_9217,N_3386,N_3414);
and U9218 (N_9218,N_5135,N_4691);
nor U9219 (N_9219,N_3882,N_5264);
or U9220 (N_9220,N_5851,N_3483);
xor U9221 (N_9221,N_6169,N_3469);
or U9222 (N_9222,N_5014,N_5132);
and U9223 (N_9223,N_4404,N_5312);
and U9224 (N_9224,N_3883,N_5659);
or U9225 (N_9225,N_3597,N_4278);
and U9226 (N_9226,N_4545,N_3527);
nor U9227 (N_9227,N_3194,N_5407);
or U9228 (N_9228,N_6235,N_5943);
nand U9229 (N_9229,N_4486,N_5956);
and U9230 (N_9230,N_3712,N_5127);
nand U9231 (N_9231,N_3230,N_3489);
or U9232 (N_9232,N_3479,N_3413);
or U9233 (N_9233,N_4425,N_3371);
nor U9234 (N_9234,N_4498,N_6166);
and U9235 (N_9235,N_3176,N_5832);
and U9236 (N_9236,N_5534,N_5270);
nor U9237 (N_9237,N_4360,N_4512);
or U9238 (N_9238,N_3323,N_5900);
or U9239 (N_9239,N_3343,N_3265);
nand U9240 (N_9240,N_5506,N_3765);
nor U9241 (N_9241,N_3170,N_4396);
or U9242 (N_9242,N_3467,N_5454);
and U9243 (N_9243,N_3285,N_5767);
and U9244 (N_9244,N_3583,N_4048);
or U9245 (N_9245,N_5659,N_6041);
and U9246 (N_9246,N_4568,N_3430);
nor U9247 (N_9247,N_4004,N_4710);
nand U9248 (N_9248,N_6240,N_5381);
and U9249 (N_9249,N_5511,N_4405);
and U9250 (N_9250,N_4210,N_5930);
nand U9251 (N_9251,N_3823,N_3609);
and U9252 (N_9252,N_3240,N_4765);
nor U9253 (N_9253,N_5030,N_6237);
and U9254 (N_9254,N_6006,N_3639);
nand U9255 (N_9255,N_5342,N_5358);
xnor U9256 (N_9256,N_4464,N_3822);
and U9257 (N_9257,N_3588,N_3150);
and U9258 (N_9258,N_4563,N_3653);
nor U9259 (N_9259,N_4727,N_6232);
nor U9260 (N_9260,N_4040,N_4732);
and U9261 (N_9261,N_5317,N_3966);
or U9262 (N_9262,N_4187,N_5280);
nand U9263 (N_9263,N_5858,N_5021);
or U9264 (N_9264,N_5024,N_4518);
nand U9265 (N_9265,N_3806,N_4371);
nor U9266 (N_9266,N_4514,N_6119);
xnor U9267 (N_9267,N_5177,N_3522);
nand U9268 (N_9268,N_5803,N_6203);
and U9269 (N_9269,N_4674,N_5228);
or U9270 (N_9270,N_5576,N_3758);
nor U9271 (N_9271,N_3611,N_4776);
nand U9272 (N_9272,N_3425,N_3362);
nand U9273 (N_9273,N_5152,N_5061);
nand U9274 (N_9274,N_3250,N_5448);
xnor U9275 (N_9275,N_3466,N_3697);
xnor U9276 (N_9276,N_4701,N_4732);
nor U9277 (N_9277,N_6107,N_4833);
nand U9278 (N_9278,N_6137,N_4614);
nor U9279 (N_9279,N_4900,N_4338);
and U9280 (N_9280,N_5125,N_3146);
and U9281 (N_9281,N_5611,N_5021);
or U9282 (N_9282,N_3520,N_5599);
and U9283 (N_9283,N_4029,N_5144);
and U9284 (N_9284,N_3469,N_5308);
nand U9285 (N_9285,N_5141,N_4592);
or U9286 (N_9286,N_4420,N_3981);
and U9287 (N_9287,N_3134,N_4829);
xnor U9288 (N_9288,N_4856,N_3756);
xnor U9289 (N_9289,N_5036,N_3658);
and U9290 (N_9290,N_3754,N_4481);
xnor U9291 (N_9291,N_6127,N_3395);
and U9292 (N_9292,N_4294,N_4970);
and U9293 (N_9293,N_4027,N_3308);
nand U9294 (N_9294,N_5573,N_5131);
nor U9295 (N_9295,N_4209,N_3277);
nand U9296 (N_9296,N_3763,N_4667);
nor U9297 (N_9297,N_4214,N_5349);
nand U9298 (N_9298,N_4295,N_4171);
or U9299 (N_9299,N_4437,N_4393);
nor U9300 (N_9300,N_3644,N_5569);
and U9301 (N_9301,N_3756,N_5805);
nor U9302 (N_9302,N_4318,N_5696);
and U9303 (N_9303,N_4230,N_5470);
nor U9304 (N_9304,N_5858,N_5056);
or U9305 (N_9305,N_4608,N_5250);
nand U9306 (N_9306,N_5360,N_4109);
xor U9307 (N_9307,N_6095,N_5459);
nand U9308 (N_9308,N_3618,N_3441);
nor U9309 (N_9309,N_3843,N_3922);
nor U9310 (N_9310,N_3978,N_5909);
and U9311 (N_9311,N_4359,N_3611);
or U9312 (N_9312,N_3890,N_5076);
nand U9313 (N_9313,N_4626,N_5584);
nor U9314 (N_9314,N_6221,N_4558);
and U9315 (N_9315,N_4933,N_3314);
and U9316 (N_9316,N_6231,N_4434);
and U9317 (N_9317,N_5675,N_6028);
nor U9318 (N_9318,N_4746,N_4614);
or U9319 (N_9319,N_3270,N_3417);
nand U9320 (N_9320,N_3264,N_4185);
nand U9321 (N_9321,N_5276,N_6068);
or U9322 (N_9322,N_5754,N_4300);
or U9323 (N_9323,N_4783,N_3826);
nor U9324 (N_9324,N_4076,N_6080);
and U9325 (N_9325,N_4515,N_4414);
or U9326 (N_9326,N_4684,N_5885);
nand U9327 (N_9327,N_4266,N_4979);
nand U9328 (N_9328,N_4175,N_3699);
and U9329 (N_9329,N_5846,N_6099);
and U9330 (N_9330,N_4929,N_5439);
and U9331 (N_9331,N_3946,N_5772);
nor U9332 (N_9332,N_5487,N_4307);
nor U9333 (N_9333,N_4215,N_5451);
or U9334 (N_9334,N_3639,N_3938);
and U9335 (N_9335,N_3296,N_4737);
or U9336 (N_9336,N_3488,N_5171);
or U9337 (N_9337,N_5496,N_5092);
nor U9338 (N_9338,N_3919,N_5600);
and U9339 (N_9339,N_4994,N_6077);
xnor U9340 (N_9340,N_5933,N_5294);
nor U9341 (N_9341,N_3133,N_3155);
nand U9342 (N_9342,N_3980,N_4822);
nand U9343 (N_9343,N_4429,N_4735);
nand U9344 (N_9344,N_3645,N_3632);
nand U9345 (N_9345,N_5150,N_4477);
nand U9346 (N_9346,N_3232,N_4749);
xnor U9347 (N_9347,N_5541,N_5157);
nor U9348 (N_9348,N_3999,N_5011);
or U9349 (N_9349,N_5350,N_5647);
nor U9350 (N_9350,N_3933,N_5836);
and U9351 (N_9351,N_4126,N_4586);
and U9352 (N_9352,N_4513,N_4950);
and U9353 (N_9353,N_3281,N_4107);
or U9354 (N_9354,N_5824,N_4357);
nand U9355 (N_9355,N_5621,N_3510);
or U9356 (N_9356,N_4724,N_5376);
nor U9357 (N_9357,N_3367,N_6238);
nand U9358 (N_9358,N_6203,N_5839);
and U9359 (N_9359,N_3872,N_5209);
or U9360 (N_9360,N_5500,N_4587);
xnor U9361 (N_9361,N_4625,N_4432);
nand U9362 (N_9362,N_3974,N_5960);
or U9363 (N_9363,N_6146,N_5403);
or U9364 (N_9364,N_3563,N_3206);
nand U9365 (N_9365,N_5860,N_3974);
nand U9366 (N_9366,N_4284,N_4204);
nor U9367 (N_9367,N_5622,N_4277);
nand U9368 (N_9368,N_5122,N_3858);
xor U9369 (N_9369,N_3647,N_3325);
nand U9370 (N_9370,N_3380,N_6090);
and U9371 (N_9371,N_3384,N_4307);
or U9372 (N_9372,N_5156,N_4043);
nand U9373 (N_9373,N_4553,N_5205);
nor U9374 (N_9374,N_4246,N_3861);
or U9375 (N_9375,N_6888,N_8820);
or U9376 (N_9376,N_9296,N_6575);
or U9377 (N_9377,N_6955,N_7624);
nor U9378 (N_9378,N_7880,N_6513);
and U9379 (N_9379,N_7046,N_8579);
or U9380 (N_9380,N_6407,N_8673);
nand U9381 (N_9381,N_6355,N_7061);
and U9382 (N_9382,N_8466,N_6889);
nand U9383 (N_9383,N_8189,N_7913);
xnor U9384 (N_9384,N_7720,N_6639);
and U9385 (N_9385,N_6844,N_8439);
nor U9386 (N_9386,N_7409,N_7645);
nor U9387 (N_9387,N_8505,N_6374);
xnor U9388 (N_9388,N_7738,N_6372);
and U9389 (N_9389,N_7454,N_7017);
and U9390 (N_9390,N_8352,N_6837);
or U9391 (N_9391,N_7415,N_7356);
or U9392 (N_9392,N_8855,N_6812);
nor U9393 (N_9393,N_8017,N_6700);
and U9394 (N_9394,N_7095,N_8784);
and U9395 (N_9395,N_9189,N_9312);
and U9396 (N_9396,N_7732,N_8679);
nor U9397 (N_9397,N_8378,N_7974);
and U9398 (N_9398,N_9138,N_6867);
nand U9399 (N_9399,N_6286,N_7243);
or U9400 (N_9400,N_9343,N_6787);
xor U9401 (N_9401,N_8893,N_8744);
or U9402 (N_9402,N_7040,N_6557);
and U9403 (N_9403,N_7188,N_9009);
nor U9404 (N_9404,N_8007,N_8083);
xnor U9405 (N_9405,N_8810,N_7097);
nand U9406 (N_9406,N_6265,N_6386);
xnor U9407 (N_9407,N_8989,N_7588);
or U9408 (N_9408,N_7165,N_7371);
or U9409 (N_9409,N_8792,N_9277);
nor U9410 (N_9410,N_6842,N_8490);
nor U9411 (N_9411,N_6493,N_7314);
nand U9412 (N_9412,N_7885,N_7685);
xor U9413 (N_9413,N_9227,N_8927);
and U9414 (N_9414,N_7080,N_6972);
or U9415 (N_9415,N_6761,N_7765);
or U9416 (N_9416,N_7386,N_8242);
or U9417 (N_9417,N_9246,N_8192);
or U9418 (N_9418,N_8484,N_8894);
nor U9419 (N_9419,N_8348,N_9339);
nand U9420 (N_9420,N_9030,N_9258);
or U9421 (N_9421,N_7241,N_7228);
nand U9422 (N_9422,N_8167,N_7033);
or U9423 (N_9423,N_8636,N_6278);
or U9424 (N_9424,N_6943,N_7769);
and U9425 (N_9425,N_6568,N_6976);
nor U9426 (N_9426,N_9336,N_8933);
and U9427 (N_9427,N_6417,N_8362);
nor U9428 (N_9428,N_8376,N_9156);
xnor U9429 (N_9429,N_6849,N_8476);
or U9430 (N_9430,N_7795,N_8285);
and U9431 (N_9431,N_7727,N_6318);
nand U9432 (N_9432,N_8351,N_8932);
or U9433 (N_9433,N_7195,N_8096);
nand U9434 (N_9434,N_8599,N_9232);
and U9435 (N_9435,N_7100,N_8848);
xor U9436 (N_9436,N_8994,N_8037);
nand U9437 (N_9437,N_7420,N_9207);
nand U9438 (N_9438,N_9025,N_7922);
and U9439 (N_9439,N_6928,N_6483);
nor U9440 (N_9440,N_7575,N_6786);
or U9441 (N_9441,N_8592,N_7231);
nand U9442 (N_9442,N_7341,N_8225);
or U9443 (N_9443,N_8394,N_7320);
nor U9444 (N_9444,N_9329,N_7150);
or U9445 (N_9445,N_8650,N_9095);
nand U9446 (N_9446,N_7625,N_7205);
nor U9447 (N_9447,N_6930,N_8906);
nor U9448 (N_9448,N_7107,N_7261);
xor U9449 (N_9449,N_8366,N_8545);
nand U9450 (N_9450,N_6688,N_6634);
and U9451 (N_9451,N_6670,N_8774);
and U9452 (N_9452,N_6971,N_6868);
and U9453 (N_9453,N_9283,N_7223);
and U9454 (N_9454,N_8067,N_8078);
nor U9455 (N_9455,N_8184,N_6910);
nor U9456 (N_9456,N_7013,N_6433);
nor U9457 (N_9457,N_8497,N_6498);
xor U9458 (N_9458,N_7042,N_9313);
nand U9459 (N_9459,N_8738,N_6940);
nor U9460 (N_9460,N_8682,N_8494);
xnor U9461 (N_9461,N_6830,N_7178);
nand U9462 (N_9462,N_8896,N_8972);
nor U9463 (N_9463,N_8742,N_8630);
nand U9464 (N_9464,N_8183,N_6739);
nand U9465 (N_9465,N_6313,N_7969);
nand U9466 (N_9466,N_8436,N_8216);
or U9467 (N_9467,N_7693,N_9174);
nor U9468 (N_9468,N_7764,N_7476);
nand U9469 (N_9469,N_7503,N_7888);
nor U9470 (N_9470,N_8332,N_8944);
nor U9471 (N_9471,N_7543,N_7418);
xor U9472 (N_9472,N_7545,N_9100);
nor U9473 (N_9473,N_6502,N_6469);
and U9474 (N_9474,N_7309,N_7316);
and U9475 (N_9475,N_8698,N_9289);
nor U9476 (N_9476,N_8125,N_7520);
or U9477 (N_9477,N_7036,N_8508);
nor U9478 (N_9478,N_8637,N_7681);
nand U9479 (N_9479,N_8945,N_7108);
xnor U9480 (N_9480,N_6798,N_8818);
nor U9481 (N_9481,N_7964,N_6749);
nor U9482 (N_9482,N_8176,N_6790);
xor U9483 (N_9483,N_7566,N_9021);
nand U9484 (N_9484,N_9228,N_6294);
and U9485 (N_9485,N_9007,N_7907);
and U9486 (N_9486,N_8209,N_7856);
and U9487 (N_9487,N_6695,N_7438);
xor U9488 (N_9488,N_9196,N_6587);
nand U9489 (N_9489,N_8547,N_7963);
or U9490 (N_9490,N_8261,N_7711);
or U9491 (N_9491,N_8008,N_8840);
nand U9492 (N_9492,N_8559,N_8799);
nand U9493 (N_9493,N_6655,N_7894);
and U9494 (N_9494,N_6295,N_9180);
and U9495 (N_9495,N_9182,N_7891);
or U9496 (N_9496,N_6298,N_8287);
nor U9497 (N_9497,N_6300,N_6906);
nor U9498 (N_9498,N_8375,N_9342);
or U9499 (N_9499,N_9347,N_8713);
nand U9500 (N_9500,N_6509,N_6991);
nand U9501 (N_9501,N_9082,N_8899);
nand U9502 (N_9502,N_8325,N_8883);
nor U9503 (N_9503,N_8942,N_6382);
nor U9504 (N_9504,N_6562,N_7069);
and U9505 (N_9505,N_9055,N_8835);
nor U9506 (N_9506,N_9241,N_8311);
nand U9507 (N_9507,N_7768,N_8664);
nor U9508 (N_9508,N_6327,N_7422);
and U9509 (N_9509,N_8863,N_6801);
nor U9510 (N_9510,N_9326,N_6452);
nand U9511 (N_9511,N_7130,N_6657);
and U9512 (N_9512,N_7020,N_9015);
nor U9513 (N_9513,N_6896,N_9224);
nand U9514 (N_9514,N_8521,N_8872);
or U9515 (N_9515,N_8589,N_7957);
nor U9516 (N_9516,N_7708,N_9051);
nand U9517 (N_9517,N_8905,N_8639);
nor U9518 (N_9518,N_8737,N_7351);
or U9519 (N_9519,N_6967,N_9341);
and U9520 (N_9520,N_8464,N_6361);
or U9521 (N_9521,N_8102,N_6503);
nand U9522 (N_9522,N_8361,N_8519);
or U9523 (N_9523,N_7073,N_8377);
or U9524 (N_9524,N_8718,N_8171);
and U9525 (N_9525,N_6561,N_8976);
or U9526 (N_9526,N_6863,N_6945);
nand U9527 (N_9527,N_6347,N_8526);
or U9528 (N_9528,N_6629,N_8719);
xnor U9529 (N_9529,N_6359,N_6291);
nor U9530 (N_9530,N_6907,N_7707);
and U9531 (N_9531,N_7583,N_6856);
nand U9532 (N_9532,N_8697,N_6258);
and U9533 (N_9533,N_7991,N_6846);
nand U9534 (N_9534,N_6541,N_6687);
nand U9535 (N_9535,N_7452,N_7971);
and U9536 (N_9536,N_7916,N_8875);
or U9537 (N_9537,N_9104,N_6705);
and U9538 (N_9538,N_7318,N_7290);
xnor U9539 (N_9539,N_6677,N_7235);
nor U9540 (N_9540,N_7984,N_8036);
and U9541 (N_9541,N_8758,N_7283);
or U9542 (N_9542,N_7267,N_8495);
and U9543 (N_9543,N_7983,N_8678);
nor U9544 (N_9544,N_8134,N_7799);
and U9545 (N_9545,N_8662,N_9158);
xnor U9546 (N_9546,N_7609,N_8728);
nor U9547 (N_9547,N_7372,N_6946);
or U9548 (N_9548,N_8703,N_7469);
and U9549 (N_9549,N_8540,N_6481);
and U9550 (N_9550,N_6693,N_9089);
and U9551 (N_9551,N_9344,N_9045);
nand U9552 (N_9552,N_9211,N_7004);
nand U9553 (N_9553,N_8132,N_6515);
or U9554 (N_9554,N_6752,N_8106);
nand U9555 (N_9555,N_9050,N_6444);
nand U9556 (N_9556,N_8239,N_8326);
or U9557 (N_9557,N_7110,N_6259);
or U9558 (N_9558,N_7676,N_8316);
or U9559 (N_9559,N_6485,N_8172);
nor U9560 (N_9560,N_7264,N_7380);
or U9561 (N_9561,N_6807,N_8460);
nor U9562 (N_9562,N_6684,N_8044);
or U9563 (N_9563,N_7849,N_7734);
or U9564 (N_9564,N_9357,N_7102);
xnor U9565 (N_9565,N_7162,N_7689);
nand U9566 (N_9566,N_7837,N_8836);
or U9567 (N_9567,N_6884,N_8343);
or U9568 (N_9568,N_9060,N_6722);
or U9569 (N_9569,N_7982,N_8983);
xor U9570 (N_9570,N_6305,N_6269);
and U9571 (N_9571,N_7389,N_8936);
or U9572 (N_9572,N_9190,N_7155);
nor U9573 (N_9573,N_6468,N_6385);
and U9574 (N_9574,N_7774,N_6252);
and U9575 (N_9575,N_6872,N_8122);
nor U9576 (N_9576,N_9194,N_7232);
nand U9577 (N_9577,N_8273,N_6584);
or U9578 (N_9578,N_7244,N_7749);
or U9579 (N_9579,N_9360,N_6900);
and U9580 (N_9580,N_7463,N_6766);
and U9581 (N_9581,N_7449,N_7801);
or U9582 (N_9582,N_8757,N_7462);
and U9583 (N_9583,N_8043,N_7035);
nand U9584 (N_9584,N_6741,N_8443);
nand U9585 (N_9585,N_8688,N_7759);
or U9586 (N_9586,N_8567,N_6559);
nand U9587 (N_9587,N_8969,N_6551);
nand U9588 (N_9588,N_7500,N_7120);
xnor U9589 (N_9589,N_7846,N_6263);
nor U9590 (N_9590,N_8564,N_7580);
or U9591 (N_9591,N_8309,N_8873);
and U9592 (N_9592,N_8594,N_8568);
or U9593 (N_9593,N_8203,N_7201);
nor U9594 (N_9594,N_8951,N_8667);
nor U9595 (N_9595,N_7074,N_8268);
nand U9596 (N_9596,N_9008,N_6949);
or U9597 (N_9597,N_8344,N_8197);
or U9598 (N_9598,N_7375,N_8014);
or U9599 (N_9599,N_8633,N_7519);
or U9600 (N_9600,N_8852,N_6979);
or U9601 (N_9601,N_7701,N_7174);
nand U9602 (N_9602,N_6871,N_8108);
or U9603 (N_9603,N_9003,N_7614);
nor U9604 (N_9604,N_7824,N_6886);
and U9605 (N_9605,N_6340,N_7731);
and U9606 (N_9606,N_8930,N_7972);
or U9607 (N_9607,N_8700,N_7426);
or U9608 (N_9608,N_6778,N_6637);
and U9609 (N_9609,N_6429,N_6609);
nand U9610 (N_9610,N_6363,N_7970);
and U9611 (N_9611,N_9142,N_7674);
nor U9612 (N_9612,N_8081,N_7822);
nor U9613 (N_9613,N_8024,N_7254);
nor U9614 (N_9614,N_6625,N_9058);
nand U9615 (N_9615,N_8558,N_8741);
nand U9616 (N_9616,N_8621,N_7112);
nor U9617 (N_9617,N_8339,N_8957);
nand U9618 (N_9618,N_6831,N_7159);
and U9619 (N_9619,N_6306,N_8919);
and U9620 (N_9620,N_7555,N_8860);
nor U9621 (N_9621,N_6572,N_7632);
and U9622 (N_9622,N_8004,N_7239);
and U9623 (N_9623,N_6658,N_7898);
nand U9624 (N_9624,N_6471,N_6708);
and U9625 (N_9625,N_6810,N_8958);
xnor U9626 (N_9626,N_8692,N_8337);
nor U9627 (N_9627,N_7412,N_6524);
nand U9628 (N_9628,N_7302,N_9144);
nand U9629 (N_9629,N_8033,N_7293);
or U9630 (N_9630,N_7180,N_6488);
nor U9631 (N_9631,N_7203,N_8626);
nor U9632 (N_9632,N_7639,N_7862);
nand U9633 (N_9633,N_6648,N_6343);
or U9634 (N_9634,N_6934,N_7820);
and U9635 (N_9635,N_8502,N_7581);
nor U9636 (N_9636,N_6999,N_7882);
and U9637 (N_9637,N_8350,N_7276);
nor U9638 (N_9638,N_7382,N_6475);
nand U9639 (N_9639,N_8072,N_8533);
nor U9640 (N_9640,N_6850,N_6839);
nand U9641 (N_9641,N_6342,N_7817);
xnor U9642 (N_9642,N_7604,N_9071);
nor U9643 (N_9643,N_8726,N_7712);
nor U9644 (N_9644,N_7656,N_8065);
or U9645 (N_9645,N_8243,N_7561);
and U9646 (N_9646,N_7401,N_7872);
nor U9647 (N_9647,N_6783,N_8303);
nand U9648 (N_9648,N_7474,N_6556);
nand U9649 (N_9649,N_8315,N_8995);
nor U9650 (N_9650,N_8949,N_8897);
nor U9651 (N_9651,N_6393,N_7027);
and U9652 (N_9652,N_6516,N_8885);
and U9653 (N_9653,N_8960,N_6765);
xor U9654 (N_9654,N_6462,N_7251);
nor U9655 (N_9655,N_8010,N_8890);
and U9656 (N_9656,N_7868,N_9185);
or U9657 (N_9657,N_7094,N_7839);
xor U9658 (N_9658,N_8272,N_9124);
nor U9659 (N_9659,N_8864,N_8405);
nor U9660 (N_9660,N_6354,N_8812);
nand U9661 (N_9661,N_8101,N_8003);
xor U9662 (N_9662,N_7496,N_8088);
nor U9663 (N_9663,N_7920,N_7410);
nor U9664 (N_9664,N_7168,N_8305);
or U9665 (N_9665,N_7870,N_7364);
and U9666 (N_9666,N_7976,N_9327);
or U9667 (N_9667,N_6998,N_8211);
nor U9668 (N_9668,N_9036,N_7746);
and U9669 (N_9669,N_6543,N_7833);
and U9670 (N_9670,N_7050,N_7640);
or U9671 (N_9671,N_6470,N_7941);
or U9672 (N_9672,N_7531,N_6627);
nor U9673 (N_9673,N_8259,N_7238);
nor U9674 (N_9674,N_6733,N_6981);
nand U9675 (N_9675,N_8605,N_6370);
xor U9676 (N_9676,N_7761,N_8665);
nor U9677 (N_9677,N_8298,N_7128);
or U9678 (N_9678,N_8373,N_9090);
xnor U9679 (N_9679,N_8838,N_7329);
nand U9680 (N_9680,N_8068,N_7446);
nor U9681 (N_9681,N_7284,N_7899);
or U9682 (N_9682,N_6893,N_8907);
nand U9683 (N_9683,N_6508,N_8821);
and U9684 (N_9684,N_7798,N_8583);
nand U9685 (N_9685,N_8510,N_8286);
and U9686 (N_9686,N_6995,N_6589);
nand U9687 (N_9687,N_6903,N_6299);
xor U9688 (N_9688,N_8485,N_6987);
and U9689 (N_9689,N_8137,N_6379);
nand U9690 (N_9690,N_8727,N_7395);
nor U9691 (N_9691,N_8996,N_7247);
or U9692 (N_9692,N_7842,N_6605);
and U9693 (N_9693,N_7925,N_9113);
and U9694 (N_9694,N_7751,N_8251);
or U9695 (N_9695,N_8699,N_7466);
and U9696 (N_9696,N_8593,N_8903);
or U9697 (N_9697,N_7047,N_9330);
and U9698 (N_9698,N_7439,N_6691);
xnor U9699 (N_9699,N_7631,N_7009);
nor U9700 (N_9700,N_7477,N_7910);
xor U9701 (N_9701,N_8246,N_6449);
nand U9702 (N_9702,N_7841,N_8180);
and U9703 (N_9703,N_9040,N_8961);
or U9704 (N_9704,N_8554,N_6970);
nand U9705 (N_9705,N_7657,N_9364);
nor U9706 (N_9706,N_8629,N_7758);
nand U9707 (N_9707,N_6740,N_7230);
nor U9708 (N_9708,N_8797,N_7305);
xor U9709 (N_9709,N_7266,N_9297);
nor U9710 (N_9710,N_8515,N_9168);
or U9711 (N_9711,N_9251,N_6496);
nand U9712 (N_9712,N_8914,N_7973);
and U9713 (N_9713,N_7537,N_6545);
nand U9714 (N_9714,N_8543,N_8837);
and U9715 (N_9715,N_9374,N_7608);
and U9716 (N_9716,N_6890,N_7958);
xnor U9717 (N_9717,N_8469,N_8159);
or U9718 (N_9718,N_7330,N_6679);
nor U9719 (N_9719,N_7687,N_8622);
or U9720 (N_9720,N_6885,N_8188);
or U9721 (N_9721,N_7343,N_7492);
and U9722 (N_9722,N_9022,N_7222);
and U9723 (N_9723,N_6579,N_8452);
and U9724 (N_9724,N_8981,N_6308);
and U9725 (N_9725,N_8028,N_8432);
or U9726 (N_9726,N_8750,N_8210);
or U9727 (N_9727,N_8206,N_7980);
nor U9728 (N_9728,N_9233,N_7427);
xor U9729 (N_9729,N_6350,N_8498);
nor U9730 (N_9730,N_7510,N_7381);
or U9731 (N_9731,N_9026,N_7664);
nand U9732 (N_9732,N_7863,N_9340);
or U9733 (N_9733,N_6757,N_7873);
nand U9734 (N_9734,N_7887,N_7357);
nand U9735 (N_9735,N_6391,N_8112);
and U9736 (N_9736,N_8631,N_9069);
or U9737 (N_9737,N_7985,N_7498);
and U9738 (N_9738,N_8710,N_6806);
and U9739 (N_9739,N_7805,N_6319);
nand U9740 (N_9740,N_7612,N_7124);
nor U9741 (N_9741,N_6723,N_8051);
nand U9742 (N_9742,N_6411,N_7635);
nor U9743 (N_9743,N_9331,N_7786);
or U9744 (N_9744,N_7179,N_7585);
and U9745 (N_9745,N_8947,N_7743);
nand U9746 (N_9746,N_7869,N_6768);
or U9747 (N_9747,N_7505,N_7258);
nor U9748 (N_9748,N_7425,N_7852);
or U9749 (N_9749,N_9114,N_6333);
nand U9750 (N_9750,N_6368,N_8098);
xnor U9751 (N_9751,N_7365,N_6915);
nand U9752 (N_9752,N_7391,N_6642);
or U9753 (N_9753,N_7806,N_8714);
nand U9754 (N_9754,N_9105,N_7298);
nand U9755 (N_9755,N_6732,N_8458);
nand U9756 (N_9756,N_9130,N_8548);
or U9757 (N_9757,N_8752,N_7045);
or U9758 (N_9758,N_6529,N_8552);
and U9759 (N_9759,N_7171,N_8217);
nand U9760 (N_9760,N_6489,N_7221);
xor U9761 (N_9761,N_7457,N_6977);
nand U9762 (N_9762,N_9188,N_8763);
or U9763 (N_9763,N_6989,N_9367);
and U9764 (N_9764,N_8623,N_8720);
nor U9765 (N_9765,N_7948,N_8089);
nor U9766 (N_9766,N_6951,N_7726);
nor U9767 (N_9767,N_6950,N_7952);
xor U9768 (N_9768,N_7650,N_6656);
or U9769 (N_9769,N_7661,N_9276);
nor U9770 (N_9770,N_7483,N_7029);
and U9771 (N_9771,N_8569,N_8668);
and U9772 (N_9772,N_7811,N_7131);
and U9773 (N_9773,N_6310,N_9333);
or U9774 (N_9774,N_7959,N_7953);
or U9775 (N_9775,N_6544,N_6501);
nand U9776 (N_9776,N_8321,N_8116);
nor U9777 (N_9777,N_9119,N_7603);
and U9778 (N_9778,N_8295,N_6709);
nor U9779 (N_9779,N_8620,N_9112);
or U9780 (N_9780,N_6344,N_7190);
and U9781 (N_9781,N_7993,N_7242);
and U9782 (N_9782,N_7549,N_6953);
xor U9783 (N_9783,N_9346,N_7400);
nor U9784 (N_9784,N_6957,N_6978);
nand U9785 (N_9785,N_6536,N_7554);
nand U9786 (N_9786,N_7350,N_6369);
or U9787 (N_9787,N_8114,N_6565);
or U9788 (N_9788,N_7197,N_6720);
or U9789 (N_9789,N_6577,N_9217);
xor U9790 (N_9790,N_7234,N_7473);
and U9791 (N_9791,N_7809,N_7481);
and U9792 (N_9792,N_6828,N_6861);
nand U9793 (N_9793,N_8479,N_8401);
and U9794 (N_9794,N_8222,N_6769);
nor U9795 (N_9795,N_8045,N_7023);
or U9796 (N_9796,N_8214,N_7275);
and U9797 (N_9797,N_7954,N_9239);
or U9798 (N_9798,N_7556,N_9024);
xnor U9799 (N_9799,N_8653,N_8560);
nor U9800 (N_9800,N_6985,N_7670);
or U9801 (N_9801,N_7838,N_9157);
or U9802 (N_9802,N_9369,N_7535);
or U9803 (N_9803,N_8909,N_6583);
nand U9804 (N_9804,N_6823,N_6459);
xor U9805 (N_9805,N_6659,N_8397);
and U9806 (N_9806,N_7273,N_8783);
and U9807 (N_9807,N_8470,N_7943);
nand U9808 (N_9808,N_8580,N_9193);
nand U9809 (N_9809,N_8025,N_9257);
or U9810 (N_9810,N_8590,N_8732);
or U9811 (N_9811,N_7792,N_8415);
and U9812 (N_9812,N_8975,N_9309);
nand U9813 (N_9813,N_6593,N_8091);
nand U9814 (N_9814,N_7643,N_8241);
nand U9815 (N_9815,N_7779,N_6697);
or U9816 (N_9816,N_6713,N_8127);
and U9817 (N_9817,N_8701,N_6833);
nor U9818 (N_9818,N_6388,N_7133);
nand U9819 (N_9819,N_9308,N_8227);
or U9820 (N_9820,N_7750,N_7123);
and U9821 (N_9821,N_8849,N_9147);
and U9822 (N_9822,N_7177,N_8787);
and U9823 (N_9823,N_8943,N_7630);
and U9824 (N_9824,N_8154,N_8634);
nand U9825 (N_9825,N_6824,N_7334);
nor U9826 (N_9826,N_6686,N_6865);
nor U9827 (N_9827,N_6647,N_7327);
xnor U9828 (N_9828,N_7667,N_8586);
nand U9829 (N_9829,N_7344,N_8293);
nand U9830 (N_9830,N_6406,N_8866);
nor U9831 (N_9831,N_9334,N_7960);
and U9832 (N_9832,N_7010,N_7877);
nor U9833 (N_9833,N_8765,N_7240);
nor U9834 (N_9834,N_8384,N_6307);
and U9835 (N_9835,N_6292,N_7928);
and U9836 (N_9836,N_6270,N_6706);
or U9837 (N_9837,N_7488,N_8511);
or U9838 (N_9838,N_6546,N_6698);
and U9839 (N_9839,N_9314,N_9290);
nand U9840 (N_9840,N_8959,N_8882);
xor U9841 (N_9841,N_8082,N_7099);
nand U9842 (N_9842,N_7840,N_6454);
nor U9843 (N_9843,N_7883,N_8483);
nand U9844 (N_9844,N_7186,N_8472);
nand U9845 (N_9845,N_7005,N_8212);
and U9846 (N_9846,N_6392,N_9181);
or U9847 (N_9847,N_7349,N_9295);
or U9848 (N_9848,N_9261,N_9213);
or U9849 (N_9849,N_6427,N_7724);
nand U9850 (N_9850,N_8912,N_6775);
nand U9851 (N_9851,N_8830,N_6415);
xnor U9852 (N_9852,N_8367,N_8674);
nand U9853 (N_9853,N_6604,N_7704);
nor U9854 (N_9854,N_8808,N_7596);
nand U9855 (N_9855,N_8473,N_7995);
or U9856 (N_9856,N_8754,N_7066);
nand U9857 (N_9857,N_9206,N_6814);
nor U9858 (N_9858,N_6821,N_6781);
nor U9859 (N_9859,N_8739,N_8607);
or U9860 (N_9860,N_6840,N_6378);
or U9861 (N_9861,N_8155,N_7270);
and U9862 (N_9862,N_6473,N_8111);
or U9863 (N_9863,N_8077,N_6699);
nand U9864 (N_9864,N_7695,N_7574);
nand U9865 (N_9865,N_6419,N_8652);
nor U9866 (N_9866,N_8874,N_6277);
xor U9867 (N_9867,N_9358,N_9153);
xor U9868 (N_9868,N_8953,N_8963);
nor U9869 (N_9869,N_9278,N_7322);
nand U9870 (N_9870,N_9315,N_7508);
and U9871 (N_9871,N_9264,N_6869);
or U9872 (N_9872,N_6395,N_6667);
or U9873 (N_9873,N_6377,N_7618);
nor U9874 (N_9874,N_6816,N_8115);
nand U9875 (N_9875,N_7699,N_7051);
or U9876 (N_9876,N_8709,N_7407);
nand U9877 (N_9877,N_8901,N_8048);
nand U9878 (N_9878,N_7363,N_6289);
nand U9879 (N_9879,N_8928,N_9222);
or U9880 (N_9880,N_8218,N_6811);
or U9881 (N_9881,N_8453,N_8815);
nor U9882 (N_9882,N_9099,N_7737);
or U9883 (N_9883,N_9267,N_7560);
nor U9884 (N_9884,N_8522,N_8409);
nand U9885 (N_9885,N_8121,N_6841);
xor U9886 (N_9886,N_7771,N_8926);
and U9887 (N_9887,N_9037,N_7855);
nand U9888 (N_9888,N_6923,N_7942);
nor U9889 (N_9889,N_7728,N_8382);
and U9890 (N_9890,N_8418,N_8990);
nor U9891 (N_9891,N_9120,N_7161);
nand U9892 (N_9892,N_8651,N_6439);
and U9893 (N_9893,N_7119,N_6570);
and U9894 (N_9894,N_7649,N_8721);
nor U9895 (N_9895,N_7878,N_7893);
nor U9896 (N_9896,N_8329,N_8603);
nand U9897 (N_9897,N_8313,N_9362);
xor U9898 (N_9898,N_8616,N_7536);
nor U9899 (N_9899,N_9205,N_9048);
xor U9900 (N_9900,N_9249,N_8435);
nand U9901 (N_9901,N_6624,N_6437);
xnor U9902 (N_9902,N_6754,N_7333);
xnor U9903 (N_9903,N_8284,N_8358);
nor U9904 (N_9904,N_9311,N_7722);
nor U9905 (N_9905,N_7886,N_6387);
xor U9906 (N_9906,N_9049,N_8060);
and U9907 (N_9907,N_6414,N_8266);
or U9908 (N_9908,N_7497,N_8788);
nand U9909 (N_9909,N_6283,N_8877);
nor U9910 (N_9910,N_9057,N_8807);
and U9911 (N_9911,N_6323,N_7039);
and U9912 (N_9912,N_7918,N_8465);
or U9913 (N_9913,N_7062,N_8841);
nand U9914 (N_9914,N_7166,N_7812);
nor U9915 (N_9915,N_7495,N_8398);
nor U9916 (N_9916,N_8643,N_6748);
nand U9917 (N_9917,N_8428,N_6360);
nor U9918 (N_9918,N_8130,N_8006);
or U9919 (N_9919,N_8878,N_7376);
xor U9920 (N_9920,N_7257,N_7458);
nor U9921 (N_9921,N_6826,N_8277);
xor U9922 (N_9922,N_8238,N_8451);
nor U9923 (N_9923,N_6933,N_8986);
and U9924 (N_9924,N_6472,N_6549);
nor U9925 (N_9925,N_7977,N_9352);
or U9926 (N_9926,N_9041,N_6610);
nand U9927 (N_9927,N_9067,N_6965);
or U9928 (N_9928,N_8563,N_9353);
nand U9929 (N_9929,N_7548,N_8123);
nand U9930 (N_9930,N_7815,N_6681);
nand U9931 (N_9931,N_7914,N_7299);
nand U9932 (N_9932,N_8880,N_6891);
or U9933 (N_9933,N_8759,N_8778);
or U9934 (N_9934,N_6262,N_9151);
nor U9935 (N_9935,N_9316,N_7992);
or U9936 (N_9936,N_8832,N_9125);
and U9937 (N_9937,N_8534,N_6398);
or U9938 (N_9938,N_6297,N_7530);
nand U9939 (N_9939,N_7544,N_7090);
nor U9940 (N_9940,N_8600,N_7271);
and U9941 (N_9941,N_6512,N_8300);
or U9942 (N_9942,N_7683,N_8263);
xnor U9943 (N_9943,N_6969,N_9317);
nand U9944 (N_9944,N_7434,N_8531);
or U9945 (N_9945,N_6389,N_7063);
nor U9946 (N_9946,N_8020,N_9046);
nand U9947 (N_9947,N_6399,N_8095);
and U9948 (N_9948,N_7633,N_7628);
nand U9949 (N_9949,N_6879,N_7307);
and U9950 (N_9950,N_7331,N_6808);
nor U9951 (N_9951,N_8440,N_7367);
nand U9952 (N_9952,N_9366,N_6980);
nor U9953 (N_9953,N_8798,N_8118);
nand U9954 (N_9954,N_7182,N_7291);
nor U9955 (N_9955,N_6357,N_6920);
xnor U9956 (N_9956,N_9092,N_7864);
xor U9957 (N_9957,N_7529,N_7834);
nand U9958 (N_9958,N_7101,N_7760);
and U9959 (N_9959,N_8179,N_8231);
xor U9960 (N_9960,N_7338,N_6615);
xor U9961 (N_9961,N_8092,N_6526);
or U9962 (N_9962,N_9014,N_6573);
nor U9963 (N_9963,N_6682,N_7219);
xor U9964 (N_9964,N_8196,N_7034);
xnor U9965 (N_9965,N_8320,N_6728);
nand U9966 (N_9966,N_8357,N_6416);
or U9967 (N_9967,N_7370,N_7002);
nor U9968 (N_9968,N_7807,N_8323);
nor U9969 (N_9969,N_6497,N_6925);
or U9970 (N_9970,N_7672,N_6371);
or U9971 (N_9971,N_7206,N_7443);
or U9972 (N_9972,N_9348,N_7605);
or U9973 (N_9973,N_8506,N_8421);
nor U9974 (N_9974,N_8071,N_7790);
or U9975 (N_9975,N_7646,N_8074);
nor U9976 (N_9976,N_8468,N_6422);
or U9977 (N_9977,N_7816,N_6796);
or U9978 (N_9978,N_7209,N_9132);
nand U9979 (N_9979,N_8480,N_7615);
nand U9980 (N_9980,N_6782,N_7310);
xnor U9981 (N_9981,N_7620,N_9098);
nor U9982 (N_9982,N_6866,N_7606);
and U9983 (N_9983,N_6607,N_7861);
nand U9984 (N_9984,N_8322,N_8555);
xor U9985 (N_9985,N_6533,N_7472);
or U9986 (N_9986,N_7086,N_6793);
and U9987 (N_9987,N_6435,N_7259);
or U9988 (N_9988,N_8696,N_6505);
or U9989 (N_9989,N_8867,N_8649);
or U9990 (N_9990,N_8185,N_8768);
nor U9991 (N_9991,N_8686,N_6675);
nand U9992 (N_9992,N_7280,N_9247);
xnor U9993 (N_9993,N_6663,N_8113);
nand U9994 (N_9994,N_7845,N_9121);
nor U9995 (N_9995,N_9097,N_7227);
xor U9996 (N_9996,N_7871,N_7153);
and U9997 (N_9997,N_6736,N_8638);
nand U9998 (N_9998,N_7589,N_7288);
and U9999 (N_9999,N_9225,N_8833);
or U10000 (N_10000,N_9106,N_7906);
or U10001 (N_10001,N_8794,N_8550);
nor U10002 (N_10002,N_9203,N_6820);
nor U10003 (N_10003,N_7460,N_8429);
nor U10004 (N_10004,N_8381,N_7929);
and U10005 (N_10005,N_7352,N_8399);
nand U10006 (N_10006,N_7319,N_8230);
nand U10007 (N_10007,N_8193,N_9361);
and U10008 (N_10008,N_8312,N_6804);
and U10009 (N_10009,N_7025,N_6702);
nand U10010 (N_10010,N_8086,N_9240);
nand U10011 (N_10011,N_8402,N_6514);
and U10012 (N_10012,N_7680,N_8891);
and U10013 (N_10013,N_8079,N_8481);
xnor U10014 (N_10014,N_7057,N_6302);
nor U10015 (N_10015,N_7301,N_6751);
xor U10016 (N_10016,N_9177,N_7105);
xnor U10017 (N_10017,N_7431,N_6538);
nand U10018 (N_10018,N_7818,N_8974);
nand U10019 (N_10019,N_7269,N_7602);
and U10020 (N_10020,N_6596,N_7173);
or U10021 (N_10021,N_9363,N_9354);
and U10022 (N_10022,N_8753,N_9281);
nor U10023 (N_10023,N_6446,N_7622);
xor U10024 (N_10024,N_6613,N_8582);
and U10025 (N_10025,N_7032,N_6491);
nor U10026 (N_10026,N_9135,N_7404);
nand U10027 (N_10027,N_6905,N_8151);
nand U10028 (N_10028,N_7595,N_6476);
or U10029 (N_10029,N_7467,N_7185);
nor U10030 (N_10030,N_9139,N_8734);
or U10031 (N_10031,N_8170,N_6747);
nor U10032 (N_10032,N_8748,N_7324);
nor U10033 (N_10033,N_6268,N_8174);
and U10034 (N_10034,N_8380,N_6982);
or U10035 (N_10035,N_6380,N_6986);
nor U10036 (N_10036,N_6803,N_7785);
and U10037 (N_10037,N_9013,N_6772);
nor U10038 (N_10038,N_8290,N_6582);
nor U10039 (N_10039,N_8057,N_7085);
nand U10040 (N_10040,N_7379,N_6346);
xor U10041 (N_10041,N_8107,N_9087);
and U10042 (N_10042,N_6852,N_8868);
nand U10043 (N_10043,N_6606,N_7937);
nor U10044 (N_10044,N_6598,N_6784);
or U10045 (N_10045,N_6770,N_6843);
nand U10046 (N_10046,N_7246,N_6959);
nor U10047 (N_10047,N_6956,N_6564);
and U10048 (N_10048,N_6540,N_8858);
xor U10049 (N_10049,N_6690,N_8161);
xor U10050 (N_10050,N_8064,N_8952);
nor U10051 (N_10051,N_7719,N_6311);
xor U10052 (N_10052,N_7600,N_8427);
nor U10053 (N_10053,N_6330,N_7773);
xnor U10054 (N_10054,N_8781,N_7865);
nor U10055 (N_10055,N_9145,N_7998);
nor U10056 (N_10056,N_8411,N_9218);
xor U10057 (N_10057,N_8984,N_6535);
or U10058 (N_10058,N_7456,N_8388);
nor U10059 (N_10059,N_7881,N_8887);
or U10060 (N_10060,N_8931,N_6486);
and U10061 (N_10061,N_8449,N_8328);
nor U10062 (N_10062,N_7511,N_8501);
xor U10063 (N_10063,N_8829,N_7994);
and U10064 (N_10064,N_6650,N_9002);
and U10065 (N_10065,N_7154,N_8201);
or U10066 (N_10066,N_7669,N_7064);
and U10067 (N_10067,N_7884,N_7528);
or U10068 (N_10068,N_7903,N_6458);
and U10069 (N_10069,N_8142,N_8881);
and U10070 (N_10070,N_9012,N_8632);
nor U10071 (N_10071,N_8624,N_8283);
nor U10072 (N_10072,N_8245,N_6936);
and U10073 (N_10073,N_8250,N_6902);
and U10074 (N_10074,N_7204,N_7579);
and U10075 (N_10075,N_7419,N_9118);
or U10076 (N_10076,N_9235,N_6964);
nor U10077 (N_10077,N_6576,N_6581);
nand U10078 (N_10078,N_8681,N_7076);
or U10079 (N_10079,N_6616,N_8827);
and U10080 (N_10080,N_7245,N_7393);
or U10081 (N_10081,N_6984,N_7706);
and U10082 (N_10082,N_6791,N_9043);
or U10083 (N_10083,N_6345,N_6621);
and U10084 (N_10084,N_7564,N_6952);
nand U10085 (N_10085,N_8516,N_8964);
and U10086 (N_10086,N_8918,N_8117);
and U10087 (N_10087,N_6255,N_8002);
nor U10088 (N_10088,N_8032,N_7482);
or U10089 (N_10089,N_7647,N_6394);
nor U10090 (N_10090,N_7850,N_7772);
nand U10091 (N_10091,N_6904,N_9328);
nand U10092 (N_10092,N_9059,N_6622);
nor U10093 (N_10093,N_8224,N_7858);
nor U10094 (N_10094,N_7491,N_8598);
nand U10095 (N_10095,N_7295,N_7136);
and U10096 (N_10096,N_6403,N_7041);
and U10097 (N_10097,N_8052,N_6316);
xnor U10098 (N_10098,N_7233,N_8715);
or U10099 (N_10099,N_7797,N_6281);
and U10100 (N_10100,N_8026,N_9053);
nand U10101 (N_10101,N_7569,N_6453);
or U10102 (N_10102,N_6595,N_9307);
nand U10103 (N_10103,N_7787,N_7317);
or U10104 (N_10104,N_7892,N_8542);
nor U10105 (N_10105,N_8450,N_7999);
nand U10106 (N_10106,N_7255,N_6287);
nand U10107 (N_10107,N_8400,N_8371);
and U10108 (N_10108,N_8455,N_6594);
nor U10109 (N_10109,N_9338,N_9072);
nand U10110 (N_10110,N_6390,N_7024);
or U10111 (N_10111,N_8302,N_7694);
or U10112 (N_10112,N_9163,N_8318);
and U10113 (N_10113,N_6992,N_7677);
or U10114 (N_10114,N_8257,N_6760);
nand U10115 (N_10115,N_7780,N_6467);
nor U10116 (N_10116,N_8165,N_7160);
and U10117 (N_10117,N_8946,N_7216);
nor U10118 (N_10118,N_7229,N_7022);
xor U10119 (N_10119,N_9062,N_6511);
nor U10120 (N_10120,N_8346,N_6618);
nand U10121 (N_10121,N_9356,N_6743);
and U10122 (N_10122,N_8143,N_9052);
xor U10123 (N_10123,N_6451,N_6948);
and U10124 (N_10124,N_9070,N_8767);
or U10125 (N_10125,N_8546,N_8746);
or U10126 (N_10126,N_7104,N_8140);
or U10127 (N_10127,N_6400,N_6701);
nor U10128 (N_10128,N_7277,N_6759);
nand U10129 (N_10129,N_6428,N_8488);
nor U10130 (N_10130,N_7691,N_7217);
nor U10131 (N_10131,N_7163,N_8910);
or U10132 (N_10132,N_9140,N_7804);
nor U10133 (N_10133,N_6410,N_7475);
nor U10134 (N_10134,N_8761,N_6431);
nor U10135 (N_10135,N_7782,N_6358);
nor U10136 (N_10136,N_8562,N_6954);
nand U10137 (N_10137,N_8379,N_7360);
nand U10138 (N_10138,N_8278,N_7098);
and U10139 (N_10139,N_6550,N_7028);
and U10140 (N_10140,N_7506,N_6799);
nand U10141 (N_10141,N_6617,N_7065);
and U10142 (N_10142,N_6874,N_6636);
and U10143 (N_10143,N_8570,N_7947);
and U10144 (N_10144,N_7684,N_7946);
or U10145 (N_10145,N_6296,N_8571);
or U10146 (N_10146,N_7175,N_8396);
and U10147 (N_10147,N_7208,N_7369);
or U10148 (N_10148,N_8487,N_9248);
and U10149 (N_10149,N_6555,N_6815);
or U10150 (N_10150,N_7279,N_7156);
xor U10151 (N_10151,N_8444,N_8208);
or U10152 (N_10152,N_6776,N_9167);
or U10153 (N_10153,N_6443,N_7459);
or U10154 (N_10154,N_8041,N_7796);
or U10155 (N_10155,N_7346,N_7923);
or U10156 (N_10156,N_6396,N_6336);
or U10157 (N_10157,N_7377,N_6937);
nand U10158 (N_10158,N_8162,N_8288);
nand U10159 (N_10159,N_9324,N_7917);
and U10160 (N_10160,N_9129,N_7089);
xor U10161 (N_10161,N_6669,N_6994);
or U10162 (N_10162,N_9038,N_6499);
nand U10163 (N_10163,N_7557,N_7829);
nor U10164 (N_10164,N_7844,N_6716);
nand U10165 (N_10165,N_8968,N_7905);
nand U10166 (N_10166,N_6795,N_6897);
or U10167 (N_10167,N_6825,N_8680);
nand U10168 (N_10168,N_7335,N_7311);
nor U10169 (N_10169,N_8528,N_8749);
nand U10170 (N_10170,N_7468,N_6895);
nor U10171 (N_10171,N_7617,N_6504);
nand U10172 (N_10172,N_9000,N_9065);
and U10173 (N_10173,N_8553,N_8731);
nor U10174 (N_10174,N_8149,N_7879);
and U10175 (N_10175,N_8707,N_8614);
nand U10176 (N_10176,N_7286,N_7587);
and U10177 (N_10177,N_8795,N_6894);
nor U10178 (N_10178,N_9073,N_6566);
or U10179 (N_10179,N_7705,N_7565);
nand U10180 (N_10180,N_8802,N_7149);
or U10181 (N_10181,N_9365,N_6334);
xnor U10182 (N_10182,N_8525,N_8751);
and U10183 (N_10183,N_8791,N_8390);
nor U10184 (N_10184,N_7437,N_7832);
and U10185 (N_10185,N_7026,N_8977);
and U10186 (N_10186,N_7675,N_6525);
or U10187 (N_10187,N_8722,N_8128);
or U10188 (N_10188,N_6478,N_6724);
and U10189 (N_10189,N_7736,N_8826);
nand U10190 (N_10190,N_7353,N_8198);
nor U10191 (N_10191,N_7781,N_8445);
and U10192 (N_10192,N_6721,N_6649);
nor U10193 (N_10193,N_7678,N_8999);
nor U10194 (N_10194,N_7436,N_7339);
nand U10195 (N_10195,N_8200,N_9200);
and U10196 (N_10196,N_7547,N_7196);
nand U10197 (N_10197,N_8053,N_7383);
nor U10198 (N_10198,N_9166,N_7610);
nand U10199 (N_10199,N_6780,N_8966);
xnor U10200 (N_10200,N_6993,N_7597);
nand U10201 (N_10201,N_7997,N_7590);
and U10202 (N_10202,N_8520,N_7702);
and U10203 (N_10203,N_8423,N_7814);
and U10204 (N_10204,N_9127,N_9280);
and U10205 (N_10205,N_8804,N_8035);
nor U10206 (N_10206,N_6530,N_9108);
xor U10207 (N_10207,N_9006,N_9063);
nand U10208 (N_10208,N_8578,N_9322);
and U10209 (N_10209,N_9284,N_7730);
nor U10210 (N_10210,N_9214,N_8462);
or U10211 (N_10211,N_7755,N_7810);
nor U10212 (N_10212,N_7770,N_6630);
or U10213 (N_10213,N_6266,N_7138);
nand U10214 (N_10214,N_9109,N_6640);
and U10215 (N_10215,N_7387,N_6672);
xnor U10216 (N_10216,N_8364,N_7740);
nor U10217 (N_10217,N_8034,N_7213);
xor U10218 (N_10218,N_7721,N_8066);
nor U10219 (N_10219,N_6689,N_9243);
nor U10220 (N_10220,N_9148,N_7433);
and U10221 (N_10221,N_6988,N_9094);
and U10222 (N_10222,N_8369,N_8493);
nor U10223 (N_10223,N_6597,N_7250);
nand U10224 (N_10224,N_8884,N_8587);
nor U10225 (N_10225,N_7679,N_8319);
nor U10226 (N_10226,N_7031,N_6731);
or U10227 (N_10227,N_9208,N_7202);
or U10228 (N_10228,N_8793,N_6883);
nand U10229 (N_10229,N_7312,N_8029);
or U10230 (N_10230,N_7800,N_7777);
nor U10231 (N_10231,N_7515,N_8886);
nand U10232 (N_10232,N_7388,N_8806);
nor U10233 (N_10233,N_8256,N_6764);
xnor U10234 (N_10234,N_7966,N_7532);
or U10235 (N_10235,N_6762,N_7874);
and U10236 (N_10236,N_8419,N_8956);
nor U10237 (N_10237,N_6938,N_8190);
or U10238 (N_10238,N_8747,N_8042);
nor U10239 (N_10239,N_8420,N_8187);
nand U10240 (N_10240,N_8645,N_6873);
nand U10241 (N_10241,N_6520,N_7791);
nor U10242 (N_10242,N_8046,N_8307);
and U10243 (N_10243,N_7374,N_6272);
or U10244 (N_10244,N_6465,N_6707);
nor U10245 (N_10245,N_8690,N_7830);
or U10246 (N_10246,N_8391,N_9355);
xor U10247 (N_10247,N_8892,N_7414);
or U10248 (N_10248,N_8948,N_9371);
or U10249 (N_10249,N_9101,N_9028);
nor U10250 (N_10250,N_6460,N_8084);
or U10251 (N_10251,N_7733,N_7634);
and U10252 (N_10252,N_7710,N_6918);
xor U10253 (N_10253,N_8012,N_6256);
or U10254 (N_10254,N_6264,N_7940);
xnor U10255 (N_10255,N_6680,N_8955);
and U10256 (N_10256,N_7499,N_9143);
or U10257 (N_10257,N_8478,N_6876);
or U10258 (N_10258,N_7875,N_7366);
nand U10259 (N_10259,N_7030,N_7576);
nor U10260 (N_10260,N_7986,N_9079);
and U10261 (N_10261,N_7808,N_8566);
nand U10262 (N_10262,N_7961,N_8131);
or U10263 (N_10263,N_7859,N_8608);
nor U10264 (N_10264,N_8437,N_7912);
or U10265 (N_10265,N_8076,N_9164);
xor U10266 (N_10266,N_7117,N_6619);
or U10267 (N_10267,N_8416,N_8022);
xnor U10268 (N_10268,N_9234,N_7577);
nand U10269 (N_10269,N_6326,N_6645);
nor U10270 (N_10270,N_8110,N_7453);
and U10271 (N_10271,N_8978,N_7249);
and U10272 (N_10272,N_6477,N_6983);
nand U10273 (N_10273,N_7616,N_9137);
nor U10274 (N_10274,N_8265,N_7866);
or U10275 (N_10275,N_9171,N_8430);
nand U10276 (N_10276,N_8387,N_9152);
nand U10277 (N_10277,N_7533,N_6523);
or U10278 (N_10278,N_7198,N_7142);
and U10279 (N_10279,N_6402,N_8503);
nor U10280 (N_10280,N_7642,N_8016);
nand U10281 (N_10281,N_8671,N_7753);
and U10282 (N_10282,N_8895,N_7037);
and U10283 (N_10283,N_6279,N_6580);
xnor U10284 (N_10284,N_9068,N_6662);
nand U10285 (N_10285,N_8666,N_8425);
or U10286 (N_10286,N_6789,N_8669);
and U10287 (N_10287,N_9083,N_9066);
or U10288 (N_10288,N_7573,N_7867);
and U10289 (N_10289,N_6494,N_7936);
nand U10290 (N_10290,N_8740,N_7794);
nand U10291 (N_10291,N_9117,N_8779);
nand U10292 (N_10292,N_8670,N_8627);
nor U10293 (N_10293,N_6608,N_7441);
nand U10294 (N_10294,N_6590,N_7486);
nor U10295 (N_10295,N_7692,N_8340);
and U10296 (N_10296,N_6282,N_8967);
and U10297 (N_10297,N_6916,N_6819);
nand U10298 (N_10298,N_8459,N_6932);
and U10299 (N_10299,N_8334,N_6563);
nand U10300 (N_10300,N_6714,N_6592);
nor U10301 (N_10301,N_6348,N_7975);
nand U10302 (N_10302,N_6750,N_9250);
and U10303 (N_10303,N_8980,N_8985);
and U10304 (N_10304,N_8276,N_8486);
and U10305 (N_10305,N_8342,N_6558);
nand U10306 (N_10306,N_9303,N_7145);
nor U10307 (N_10307,N_6321,N_7392);
nand U10308 (N_10308,N_6792,N_6696);
nand U10309 (N_10309,N_8921,N_9321);
nand U10310 (N_10310,N_9077,N_6668);
or U10311 (N_10311,N_6901,N_7200);
xnor U10312 (N_10312,N_7164,N_9074);
or U10313 (N_10313,N_7081,N_8935);
and U10314 (N_10314,N_6858,N_8523);
nand U10315 (N_10315,N_7494,N_7956);
and U10316 (N_10316,N_7078,N_8745);
nor U10317 (N_10317,N_8647,N_6254);
or U10318 (N_10318,N_8000,N_8040);
and U10319 (N_10319,N_8856,N_8279);
nor U10320 (N_10320,N_7927,N_7550);
or U10321 (N_10321,N_7408,N_6517);
or U10322 (N_10322,N_6408,N_8675);
and U10323 (N_10323,N_6926,N_8492);
nor U10324 (N_10324,N_9304,N_6973);
nor U10325 (N_10325,N_8796,N_8822);
xor U10326 (N_10326,N_7627,N_8672);
and U10327 (N_10327,N_6729,N_9282);
or U10328 (N_10328,N_7226,N_7594);
and U10329 (N_10329,N_9146,N_6644);
or U10330 (N_10330,N_8923,N_7783);
and U10331 (N_10331,N_8606,N_6588);
or U10332 (N_10332,N_7819,N_8904);
and U10333 (N_10333,N_7358,N_8920);
and U10334 (N_10334,N_7001,N_8998);
nor U10335 (N_10335,N_6641,N_7347);
and U10336 (N_10336,N_9286,N_6620);
nor U10337 (N_10337,N_7586,N_8870);
xor U10338 (N_10338,N_6963,N_8663);
or U10339 (N_10339,N_6939,N_8294);
nand U10340 (N_10340,N_9191,N_6805);
and U10341 (N_10341,N_9201,N_8572);
nor U10342 (N_10342,N_8640,N_8705);
or U10343 (N_10343,N_6284,N_8544);
and U10344 (N_10344,N_9110,N_8404);
nand U10345 (N_10345,N_7962,N_7666);
nand U10346 (N_10346,N_8433,N_8254);
or U10347 (N_10347,N_8144,N_7116);
and U10348 (N_10348,N_8139,N_8049);
and U10349 (N_10349,N_7442,N_8280);
or U10350 (N_10350,N_8965,N_6942);
and U10351 (N_10351,N_8442,N_7428);
nor U10352 (N_10352,N_7077,N_6466);
nor U10353 (N_10353,N_8597,N_7067);
nor U10354 (N_10354,N_8314,N_7789);
or U10355 (N_10355,N_9198,N_8766);
nor U10356 (N_10356,N_8805,N_7106);
nor U10357 (N_10357,N_8760,N_8158);
or U10358 (N_10358,N_8677,N_8687);
nand U10359 (N_10359,N_8056,N_8474);
or U10360 (N_10360,N_8275,N_8463);
xor U10361 (N_10361,N_6317,N_8454);
nor U10362 (N_10362,N_8496,N_8962);
nand U10363 (N_10363,N_8258,N_9220);
nand U10364 (N_10364,N_8789,N_8717);
and U10365 (N_10365,N_8865,N_8876);
or U10366 (N_10366,N_9231,N_6755);
nand U10367 (N_10367,N_6835,N_6548);
nor U10368 (N_10368,N_6974,N_7539);
xor U10369 (N_10369,N_7272,N_7570);
and U10370 (N_10370,N_8658,N_7741);
or U10371 (N_10371,N_7345,N_8085);
and U10372 (N_10372,N_8581,N_7825);
and U10373 (N_10373,N_8691,N_7084);
and U10374 (N_10374,N_9086,N_8297);
nor U10375 (N_10375,N_8019,N_7847);
nand U10376 (N_10376,N_7651,N_6875);
nor U10377 (N_10377,N_7435,N_7527);
or U10378 (N_10378,N_9319,N_7714);
nand U10379 (N_10379,N_9373,N_9287);
or U10380 (N_10380,N_7988,N_7541);
xor U10381 (N_10381,N_9044,N_8575);
xor U10382 (N_10382,N_8030,N_7285);
nand U10383 (N_10383,N_7072,N_7723);
or U10384 (N_10384,N_8306,N_6518);
nand U10385 (N_10385,N_7118,N_6779);
or U10386 (N_10386,N_8270,N_8228);
and U10387 (N_10387,N_7578,N_7626);
or U10388 (N_10388,N_6767,N_6975);
nor U10389 (N_10389,N_8551,N_8879);
or U10390 (N_10390,N_8370,N_7665);
nand U10391 (N_10391,N_8764,N_7263);
nand U10392 (N_10392,N_8178,N_8168);
nand U10393 (N_10393,N_7987,N_8308);
or U10394 (N_10394,N_6911,N_9223);
and U10395 (N_10395,N_8541,N_6822);
nand U10396 (N_10396,N_7487,N_7043);
nand U10397 (N_10397,N_7836,N_7396);
and U10398 (N_10398,N_8204,N_8413);
xnor U10399 (N_10399,N_8924,N_6290);
nand U10400 (N_10400,N_8221,N_7087);
nor U10401 (N_10401,N_7516,N_8610);
nand U10402 (N_10402,N_7748,N_8814);
nor U10403 (N_10403,N_7686,N_8099);
nor U10404 (N_10404,N_7015,N_6600);
and U10405 (N_10405,N_9136,N_7075);
nor U10406 (N_10406,N_6836,N_6756);
xor U10407 (N_10407,N_7757,N_6552);
nand U10408 (N_10408,N_8147,N_8602);
and U10409 (N_10409,N_8417,N_6404);
nand U10410 (N_10410,N_7007,N_7598);
nand U10411 (N_10411,N_8426,N_6463);
and U10412 (N_10412,N_9350,N_9237);
or U10413 (N_10413,N_7568,N_7187);
nand U10414 (N_10414,N_7336,N_9033);
xnor U10415 (N_10415,N_8129,N_8527);
xor U10416 (N_10416,N_7524,N_8491);
nand U10417 (N_10417,N_9031,N_8152);
nand U10418 (N_10418,N_7501,N_6519);
or U10419 (N_10419,N_7044,N_7793);
nor U10420 (N_10420,N_7038,N_9162);
nand U10421 (N_10421,N_7008,N_8916);
or U10422 (N_10422,N_7538,N_6746);
nor U10423 (N_10423,N_8090,N_9325);
and U10424 (N_10424,N_9202,N_6322);
nor U10425 (N_10425,N_7429,N_6434);
nor U10426 (N_10426,N_6742,N_6632);
nand U10427 (N_10427,N_9272,N_7522);
nand U10428 (N_10428,N_7079,N_7835);
nor U10429 (N_10429,N_8153,N_7328);
or U10430 (N_10430,N_7146,N_8431);
nor U10431 (N_10431,N_8509,N_7191);
or U10432 (N_10432,N_7148,N_7827);
xor U10433 (N_10433,N_8059,N_6878);
nor U10434 (N_10434,N_9056,N_6882);
nor U10435 (N_10435,N_7889,N_7700);
and U10436 (N_10436,N_9160,N_6860);
nor U10437 (N_10437,N_6560,N_7424);
or U10438 (N_10438,N_8817,N_7926);
or U10439 (N_10439,N_7430,N_8296);
or U10440 (N_10440,N_9154,N_8625);
nand U10441 (N_10441,N_6683,N_9293);
nand U10442 (N_10442,N_8094,N_8383);
and U10443 (N_10443,N_8001,N_7967);
or U10444 (N_10444,N_7003,N_7268);
or U10445 (N_10445,N_7049,N_9285);
nand U10446 (N_10446,N_6635,N_8517);
nand U10447 (N_10447,N_6809,N_6838);
and U10448 (N_10448,N_6813,N_7303);
nor U10449 (N_10449,N_9370,N_6338);
or U10450 (N_10450,N_9103,N_7945);
and U10451 (N_10451,N_6362,N_8424);
nand U10452 (N_10452,N_8565,N_6507);
nand U10453 (N_10453,N_7294,N_8133);
nor U10454 (N_10454,N_8612,N_7876);
nand U10455 (N_10455,N_7448,N_7053);
nand U10456 (N_10456,N_6864,N_8018);
or U10457 (N_10457,N_8557,N_8900);
and U10458 (N_10458,N_7304,N_9335);
and U10459 (N_10459,N_7464,N_9017);
and U10460 (N_10460,N_7176,N_9209);
and U10461 (N_10461,N_7896,N_8109);
and U10462 (N_10462,N_7542,N_6870);
and U10463 (N_10463,N_7070,N_6685);
or U10464 (N_10464,N_8857,N_9042);
nand U10465 (N_10465,N_8843,N_8786);
and U10466 (N_10466,N_8333,N_6818);
xnor U10467 (N_10467,N_7158,N_7521);
or U10468 (N_10468,N_9298,N_6328);
nor U10469 (N_10469,N_6854,N_7668);
nand U10470 (N_10470,N_6537,N_9175);
nand U10471 (N_10471,N_8937,N_7673);
nand U10472 (N_10472,N_8191,N_8743);
nand U10473 (N_10473,N_8385,N_7857);
and U10474 (N_10474,N_7648,N_6880);
or U10475 (N_10475,N_8138,N_7060);
and U10476 (N_10476,N_9351,N_8561);
and U10477 (N_10477,N_7210,N_6958);
nand U10478 (N_10478,N_8993,N_6908);
nor U10479 (N_10479,N_8823,N_8477);
and U10480 (N_10480,N_6425,N_6320);
or U10481 (N_10481,N_7282,N_6646);
nand U10482 (N_10482,N_6418,N_8839);
or U10483 (N_10483,N_8898,N_7509);
nor U10484 (N_10484,N_7109,N_6401);
nor U10485 (N_10485,N_8372,N_8889);
and U10486 (N_10486,N_6829,N_8861);
and U10487 (N_10487,N_6802,N_6734);
and U10488 (N_10488,N_7297,N_6464);
or U10489 (N_10489,N_9078,N_9245);
or U10490 (N_10490,N_7361,N_9301);
or U10491 (N_10491,N_9001,N_6851);
nand U10492 (N_10492,N_7152,N_8811);
nand U10493 (N_10493,N_8467,N_6941);
nand U10494 (N_10494,N_8164,N_8232);
nand U10495 (N_10495,N_7591,N_8226);
and U10496 (N_10496,N_8854,N_6643);
or U10497 (N_10497,N_8223,N_9275);
nor U10498 (N_10498,N_8403,N_7461);
or U10499 (N_10499,N_6966,N_7373);
nand U10500 (N_10500,N_8410,N_9155);
and U10501 (N_10501,N_9345,N_8215);
xnor U10502 (N_10502,N_9229,N_6913);
or U10503 (N_10503,N_6653,N_6929);
or U10504 (N_10504,N_6892,N_6257);
nor U10505 (N_10505,N_7644,N_9011);
nand U10506 (N_10506,N_6426,N_7014);
nand U10507 (N_10507,N_6881,N_6777);
or U10508 (N_10508,N_7979,N_8902);
and U10509 (N_10509,N_8406,N_6409);
nor U10510 (N_10510,N_8105,N_9178);
nand U10511 (N_10511,N_8126,N_7931);
nand U10512 (N_10512,N_9274,N_8327);
or U10513 (N_10513,N_7194,N_7103);
and U10514 (N_10514,N_8349,N_7512);
nand U10515 (N_10515,N_6692,N_9187);
xor U10516 (N_10516,N_8341,N_8824);
and U10517 (N_10517,N_7326,N_9096);
xor U10518 (N_10518,N_8950,N_8289);
or U10519 (N_10519,N_6329,N_8135);
nor U10520 (N_10520,N_8847,N_7021);
and U10521 (N_10521,N_6569,N_9126);
and U10522 (N_10522,N_8489,N_6712);
and U10523 (N_10523,N_7551,N_9027);
or U10524 (N_10524,N_8181,N_6753);
or U10525 (N_10525,N_7398,N_9107);
and U10526 (N_10526,N_6474,N_7274);
nand U10527 (N_10527,N_9035,N_7134);
xor U10528 (N_10528,N_9236,N_9244);
xnor U10529 (N_10529,N_6397,N_8207);
nand U10530 (N_10530,N_7068,N_6375);
or U10531 (N_10531,N_7584,N_8790);
nor U10532 (N_10532,N_8954,N_6671);
nand U10533 (N_10533,N_6276,N_6356);
or U10534 (N_10534,N_8708,N_8514);
nor U10535 (N_10535,N_9320,N_7248);
nand U10536 (N_10536,N_8938,N_7114);
nand U10537 (N_10537,N_7490,N_8846);
xnor U10538 (N_10538,N_7540,N_8233);
nor U10539 (N_10539,N_8195,N_8538);
nand U10540 (N_10540,N_8260,N_6542);
nor U10541 (N_10541,N_7127,N_7563);
xnor U10542 (N_10542,N_8365,N_6602);
nor U10543 (N_10543,N_7523,N_6717);
nor U10544 (N_10544,N_8475,N_6482);
xor U10545 (N_10545,N_7184,N_6349);
or U10546 (N_10546,N_6309,N_7621);
and U10547 (N_10547,N_6718,N_6506);
or U10548 (N_10548,N_7636,N_7144);
or U10549 (N_10549,N_8386,N_7183);
xor U10550 (N_10550,N_8368,N_6364);
nor U10551 (N_10551,N_9173,N_8353);
nand U10552 (N_10552,N_6710,N_6919);
and U10553 (N_10553,N_7725,N_6325);
and U10554 (N_10554,N_8628,N_9019);
and U10555 (N_10555,N_8706,N_8070);
or U10556 (N_10556,N_6628,N_9221);
or U10557 (N_10557,N_7900,N_8175);
and U10558 (N_10558,N_7996,N_7055);
and U10559 (N_10559,N_7934,N_7169);
or U10560 (N_10560,N_8619,N_8803);
nand U10561 (N_10561,N_8461,N_9080);
nand U10562 (N_10562,N_6611,N_6727);
and U10563 (N_10563,N_9294,N_9291);
nor U10564 (N_10564,N_6315,N_8729);
xor U10565 (N_10565,N_7752,N_7406);
nand U10566 (N_10566,N_6430,N_7915);
and U10567 (N_10567,N_8991,N_7890);
and U10568 (N_10568,N_6797,N_6436);
and U10569 (N_10569,N_8782,N_7413);
nor U10570 (N_10570,N_7613,N_7659);
and U10571 (N_10571,N_6788,N_9292);
nor U10572 (N_10572,N_8434,N_7745);
and U10573 (N_10573,N_8169,N_7821);
nand U10574 (N_10574,N_6405,N_6800);
nor U10575 (N_10575,N_6927,N_7278);
nor U10576 (N_10576,N_6626,N_8537);
and U10577 (N_10577,N_9332,N_9266);
and U10578 (N_10578,N_9254,N_8659);
xnor U10579 (N_10579,N_8317,N_6381);
nand U10580 (N_10580,N_7559,N_7315);
nor U10581 (N_10581,N_6603,N_8156);
and U10582 (N_10582,N_7059,N_7904);
and U10583 (N_10583,N_7308,N_6288);
and U10584 (N_10584,N_7016,N_8655);
nor U10585 (N_10585,N_6275,N_8530);
or U10586 (N_10586,N_9179,N_8075);
xnor U10587 (N_10587,N_8777,N_7504);
or U10588 (N_10588,N_8772,N_9263);
xnor U10589 (N_10589,N_6862,N_7911);
nand U10590 (N_10590,N_6450,N_7652);
or U10591 (N_10591,N_8087,N_8762);
nor U10592 (N_10592,N_7935,N_9271);
nor U10593 (N_10593,N_9064,N_7637);
or U10594 (N_10594,N_8499,N_6413);
and U10595 (N_10595,N_7951,N_7663);
nor U10596 (N_10596,N_7502,N_6424);
or U10597 (N_10597,N_8447,N_8576);
nand U10598 (N_10598,N_7742,N_7619);
or U10599 (N_10599,N_7655,N_8119);
nand U10600 (N_10600,N_7018,N_7716);
xor U10601 (N_10601,N_9230,N_7450);
xor U10602 (N_10602,N_7654,N_8145);
nand U10603 (N_10603,N_7362,N_7056);
nand U10604 (N_10604,N_9023,N_6898);
or U10605 (N_10605,N_7402,N_6633);
or U10606 (N_10606,N_7599,N_6745);
or U10607 (N_10607,N_8194,N_8809);
nor U10608 (N_10608,N_7147,N_9288);
xnor U10609 (N_10609,N_6456,N_7321);
nor U10610 (N_10610,N_8940,N_8512);
xor U10611 (N_10611,N_8163,N_8395);
nand U10612 (N_10612,N_7012,N_7908);
nand U10613 (N_10613,N_7141,N_7260);
or U10614 (N_10614,N_7132,N_8584);
and U10615 (N_10615,N_6365,N_7126);
and U10616 (N_10616,N_9302,N_6441);
nand U10617 (N_10617,N_8771,N_9204);
nand U10618 (N_10618,N_9159,N_6651);
nor U10619 (N_10619,N_8219,N_8695);
and U10620 (N_10620,N_8536,N_8693);
or U10621 (N_10621,N_9150,N_6521);
and U10622 (N_10622,N_7513,N_8229);
and U10623 (N_10623,N_8922,N_6271);
nand U10624 (N_10624,N_8100,N_7214);
and U10625 (N_10625,N_6531,N_7965);
or U10626 (N_10626,N_6585,N_8055);
nor U10627 (N_10627,N_6730,N_7921);
nor U10628 (N_10628,N_9306,N_9018);
or U10629 (N_10629,N_8657,N_7484);
nor U10630 (N_10630,N_8414,N_9122);
xor U10631 (N_10631,N_8009,N_7411);
nand U10632 (N_10632,N_8775,N_9170);
nand U10633 (N_10633,N_7083,N_6773);
nor U10634 (N_10634,N_8247,N_6440);
nand U10635 (N_10635,N_7989,N_7955);
nor U10636 (N_10636,N_8736,N_7006);
or U10637 (N_10637,N_8299,N_6578);
or U10638 (N_10638,N_8539,N_7729);
nor U10639 (N_10639,N_7518,N_7623);
or U10640 (N_10640,N_9165,N_8389);
nor U10641 (N_10641,N_7909,N_9172);
or U10642 (N_10642,N_9310,N_7826);
nand U10643 (N_10643,N_8712,N_6638);
and U10644 (N_10644,N_6857,N_9004);
and U10645 (N_10645,N_7167,N_8274);
nor U10646 (N_10646,N_8908,N_8825);
nor U10647 (N_10647,N_8363,N_7517);
and U10648 (N_10648,N_6704,N_7207);
nor U10649 (N_10649,N_6996,N_9149);
or U10650 (N_10650,N_7122,N_9273);
nor U10651 (N_10651,N_7924,N_8080);
or U10652 (N_10652,N_6301,N_9016);
nand U10653 (N_10653,N_8124,N_8660);
nor U10654 (N_10654,N_8199,N_6599);
or U10655 (N_10655,N_6931,N_8356);
or U10656 (N_10656,N_6774,N_8769);
nor U10657 (N_10657,N_7093,N_7129);
nand U10658 (N_10658,N_7340,N_7709);
or U10659 (N_10659,N_8262,N_9039);
and U10660 (N_10660,N_6711,N_6528);
or U10661 (N_10661,N_9216,N_7938);
xor U10662 (N_10662,N_7385,N_6253);
nand U10663 (N_10663,N_8103,N_9323);
nand U10664 (N_10664,N_6412,N_8611);
nand U10665 (N_10665,N_7778,N_8997);
nand U10666 (N_10666,N_6341,N_7000);
or U10667 (N_10667,N_8213,N_8588);
and U10668 (N_10668,N_6827,N_6914);
xnor U10669 (N_10669,N_9169,N_8988);
nand U10670 (N_10670,N_8973,N_8422);
nand U10671 (N_10671,N_8851,N_8683);
xor U10672 (N_10672,N_6674,N_9111);
xnor U10673 (N_10673,N_9253,N_7262);
or U10674 (N_10674,N_8816,N_8292);
nor U10675 (N_10675,N_8023,N_8711);
and U10676 (N_10676,N_6487,N_8005);
and U10677 (N_10677,N_9076,N_8393);
nor U10678 (N_10678,N_8330,N_6457);
or U10679 (N_10679,N_8097,N_6601);
nand U10680 (N_10680,N_7572,N_8780);
or U10681 (N_10681,N_9349,N_9305);
or U10682 (N_10682,N_8186,N_9215);
nand U10683 (N_10683,N_6366,N_9269);
and U10684 (N_10684,N_8456,N_7735);
and U10685 (N_10685,N_6273,N_7011);
nand U10686 (N_10686,N_8240,N_6676);
and U10687 (N_10687,N_6947,N_6703);
nand U10688 (N_10688,N_6960,N_8347);
nand U10689 (N_10689,N_8448,N_8408);
nor U10690 (N_10690,N_8235,N_6834);
nand U10691 (N_10691,N_8917,N_6654);
and U10692 (N_10692,N_7368,N_8500);
nor U10693 (N_10693,N_8831,N_6666);
and U10694 (N_10694,N_6591,N_8813);
nand U10695 (N_10695,N_7567,N_8441);
nand U10696 (N_10696,N_8971,N_7919);
nor U10697 (N_10697,N_8844,N_8054);
and U10698 (N_10698,N_7212,N_9047);
nand U10699 (N_10699,N_9238,N_7211);
nand U10700 (N_10700,N_6909,N_8596);
and U10701 (N_10701,N_8021,N_7558);
xnor U10702 (N_10702,N_7767,N_6853);
or U10703 (N_10703,N_8694,N_9255);
or U10704 (N_10704,N_6260,N_7143);
and U10705 (N_10705,N_9088,N_8282);
nand U10706 (N_10706,N_6335,N_8842);
nand U10707 (N_10707,N_6771,N_9268);
nand U10708 (N_10708,N_7092,N_8335);
nor U10709 (N_10709,N_6500,N_6574);
nand U10710 (N_10710,N_7480,N_6665);
or U10711 (N_10711,N_9116,N_6324);
xnor U10712 (N_10712,N_6461,N_7698);
nor U10713 (N_10713,N_8236,N_7470);
nor U10714 (N_10714,N_7287,N_6758);
xnor U10715 (N_10715,N_8120,N_8202);
nor U10716 (N_10716,N_6251,N_8819);
and U10717 (N_10717,N_6351,N_8617);
nor U10718 (N_10718,N_6660,N_7762);
nand U10719 (N_10719,N_7390,N_7224);
nor U10720 (N_10720,N_7713,N_7739);
xnor U10721 (N_10721,N_8013,N_7803);
and U10722 (N_10722,N_8457,N_9256);
and U10723 (N_10723,N_6859,N_8801);
and U10724 (N_10724,N_6887,N_8281);
or U10725 (N_10725,N_7289,N_9085);
or U10726 (N_10726,N_7776,N_7766);
nand U10727 (N_10727,N_8244,N_8929);
nor U10728 (N_10728,N_8331,N_7253);
nand U10729 (N_10729,N_6376,N_7189);
nand U10730 (N_10730,N_6432,N_8532);
nor U10731 (N_10731,N_8702,N_7641);
or U10732 (N_10732,N_8345,N_6847);
nand U10733 (N_10733,N_8635,N_9195);
or U10734 (N_10734,N_7638,N_8039);
nor U10735 (N_10735,N_8069,N_9212);
nand U10736 (N_10736,N_6832,N_7901);
nor U10737 (N_10737,N_7421,N_8136);
xnor U10738 (N_10738,N_7848,N_6492);
and U10739 (N_10739,N_6384,N_7747);
and U10740 (N_10740,N_8549,N_7236);
or U10741 (N_10741,N_7157,N_7525);
nor U10742 (N_10742,N_7851,N_9259);
xor U10743 (N_10743,N_6612,N_9081);
nor U10744 (N_10744,N_7592,N_8471);
nand U10745 (N_10745,N_7553,N_8939);
or U10746 (N_10746,N_7629,N_7493);
nand U10747 (N_10747,N_6961,N_8925);
nand U10748 (N_10748,N_7140,N_7135);
and U10749 (N_10749,N_9176,N_7902);
nand U10750 (N_10750,N_7088,N_7113);
nor U10751 (N_10751,N_8648,N_7082);
nand U10752 (N_10752,N_8093,N_6794);
nor U10753 (N_10753,N_7071,N_6737);
nor U10754 (N_10754,N_8716,N_7354);
nor U10755 (N_10755,N_8654,N_6673);
or U10756 (N_10756,N_7199,N_7788);
nand U10757 (N_10757,N_7843,N_9020);
nor U10758 (N_10758,N_7181,N_6652);
xnor U10759 (N_10759,N_9054,N_8656);
or U10760 (N_10760,N_6445,N_7514);
nor U10761 (N_10761,N_6726,N_8591);
nand U10762 (N_10762,N_7444,N_6367);
nand U10763 (N_10763,N_6490,N_8015);
nand U10764 (N_10764,N_8438,N_6261);
and U10765 (N_10765,N_7571,N_8338);
or U10766 (N_10766,N_6304,N_7096);
nor U10767 (N_10767,N_7930,N_8011);
nand U10768 (N_10768,N_6631,N_6990);
and U10769 (N_10769,N_9161,N_8324);
nand U10770 (N_10770,N_7823,N_7378);
nor U10771 (N_10771,N_6962,N_6735);
nor U10772 (N_10772,N_8205,N_7895);
nor U10773 (N_10773,N_8915,N_6293);
and U10774 (N_10774,N_7225,N_9123);
or U10775 (N_10775,N_8354,N_7281);
nor U10776 (N_10776,N_8724,N_7445);
and U10777 (N_10777,N_8061,N_6554);
nor U10778 (N_10778,N_7828,N_9093);
nor U10779 (N_10779,N_6845,N_8031);
nor U10780 (N_10780,N_9199,N_8723);
and U10781 (N_10781,N_8834,N_7939);
nand U10782 (N_10782,N_6678,N_9279);
nor U10783 (N_10783,N_7756,N_8535);
or U10784 (N_10784,N_9141,N_7048);
nor U10785 (N_10785,N_7485,N_7611);
nor U10786 (N_10786,N_7607,N_8504);
nand U10787 (N_10787,N_8157,N_7802);
xor U10788 (N_10788,N_6527,N_6586);
nor U10789 (N_10789,N_7052,N_7897);
nor U10790 (N_10790,N_8360,N_7342);
nor U10791 (N_10791,N_8301,N_7968);
and U10792 (N_10792,N_7688,N_8336);
xor U10793 (N_10793,N_8058,N_6480);
nor U10794 (N_10794,N_7121,N_7775);
nor U10795 (N_10795,N_8685,N_8828);
nor U10796 (N_10796,N_7860,N_9091);
xnor U10797 (N_10797,N_6510,N_8050);
nand U10798 (N_10798,N_7690,N_7671);
nand U10799 (N_10799,N_8182,N_9359);
nor U10800 (N_10800,N_6547,N_7653);
or U10801 (N_10801,N_8646,N_8853);
xor U10802 (N_10802,N_8676,N_7355);
or U10803 (N_10803,N_7394,N_8733);
and U10804 (N_10804,N_6715,N_7478);
nand U10805 (N_10805,N_6763,N_9368);
nor U10806 (N_10806,N_6855,N_9299);
nor U10807 (N_10807,N_8482,N_6922);
nor U10808 (N_10808,N_7682,N_7507);
or U10809 (N_10809,N_7601,N_7662);
or U10810 (N_10810,N_8027,N_8618);
nand U10811 (N_10811,N_8615,N_6479);
and U10812 (N_10812,N_9219,N_8220);
xnor U10813 (N_10813,N_8255,N_6420);
and U10814 (N_10814,N_7660,N_6785);
and U10815 (N_10815,N_8785,N_9131);
nand U10816 (N_10816,N_7054,N_7784);
and U10817 (N_10817,N_8291,N_8871);
or U10818 (N_10818,N_6438,N_7455);
xnor U10819 (N_10819,N_7981,N_7432);
or U10820 (N_10820,N_8518,N_7471);
nand U10821 (N_10821,N_8850,N_8845);
nor U10822 (N_10822,N_9184,N_6553);
nor U10823 (N_10823,N_7325,N_7091);
nor U10824 (N_10824,N_8237,N_8574);
nand U10825 (N_10825,N_7384,N_7348);
nand U10826 (N_10826,N_8604,N_6303);
and U10827 (N_10827,N_7696,N_8104);
and U10828 (N_10828,N_6944,N_6448);
and U10829 (N_10829,N_7763,N_9300);
or U10830 (N_10830,N_8577,N_6337);
or U10831 (N_10831,N_8934,N_8573);
or U10832 (N_10832,N_8595,N_9252);
nand U10833 (N_10833,N_8062,N_7479);
nor U10834 (N_10834,N_8609,N_8644);
or U10835 (N_10835,N_7323,N_7744);
and U10836 (N_10836,N_8063,N_7019);
nor U10837 (N_10837,N_9029,N_7125);
nor U10838 (N_10838,N_8253,N_7115);
nand U10839 (N_10839,N_6285,N_6495);
xor U10840 (N_10840,N_7215,N_6997);
or U10841 (N_10841,N_6383,N_8585);
or U10842 (N_10842,N_9226,N_7718);
nor U10843 (N_10843,N_9265,N_8756);
nor U10844 (N_10844,N_7831,N_9372);
nand U10845 (N_10845,N_7703,N_6312);
and U10846 (N_10846,N_7337,N_6623);
nand U10847 (N_10847,N_8987,N_8869);
and U10848 (N_10848,N_8529,N_6719);
nand U10849 (N_10849,N_8725,N_9134);
nand U10850 (N_10850,N_7990,N_8755);
and U10851 (N_10851,N_9128,N_6848);
and U10852 (N_10852,N_8166,N_9005);
and U10853 (N_10853,N_8141,N_6899);
or U10854 (N_10854,N_8735,N_8859);
nor U10855 (N_10855,N_7237,N_7754);
nor U10856 (N_10856,N_8252,N_8412);
or U10857 (N_10857,N_8911,N_8234);
and U10858 (N_10858,N_6267,N_7697);
nand U10859 (N_10859,N_6921,N_8601);
or U10860 (N_10860,N_7416,N_6353);
nand U10861 (N_10861,N_8177,N_8269);
nor U10862 (N_10862,N_9084,N_8770);
and U10863 (N_10863,N_6314,N_7170);
or U10864 (N_10864,N_9075,N_6917);
or U10865 (N_10865,N_7546,N_7582);
nor U10866 (N_10866,N_6442,N_6522);
xnor U10867 (N_10867,N_7715,N_7933);
nand U10868 (N_10868,N_6725,N_6447);
nand U10869 (N_10869,N_6421,N_7192);
nor U10870 (N_10870,N_8392,N_7397);
or U10871 (N_10871,N_8446,N_6614);
nor U10872 (N_10872,N_8146,N_7423);
nand U10873 (N_10873,N_7139,N_9061);
xor U10874 (N_10874,N_7440,N_8038);
nor U10875 (N_10875,N_6332,N_6877);
or U10876 (N_10876,N_9186,N_8888);
xor U10877 (N_10877,N_8047,N_6817);
xor U10878 (N_10878,N_9034,N_6738);
and U10879 (N_10879,N_9192,N_8982);
and U10880 (N_10880,N_8513,N_7256);
and U10881 (N_10881,N_9318,N_9197);
and U10882 (N_10882,N_8979,N_7854);
nor U10883 (N_10883,N_7944,N_9115);
nand U10884 (N_10884,N_8862,N_7658);
and U10885 (N_10885,N_6664,N_7151);
xor U10886 (N_10886,N_7111,N_8264);
and U10887 (N_10887,N_7932,N_7813);
xnor U10888 (N_10888,N_6250,N_8355);
xnor U10889 (N_10889,N_9337,N_7218);
nand U10890 (N_10890,N_6331,N_7950);
or U10891 (N_10891,N_8556,N_8150);
or U10892 (N_10892,N_6744,N_7552);
and U10893 (N_10893,N_8160,N_7399);
xor U10894 (N_10894,N_6532,N_6571);
and U10895 (N_10895,N_9010,N_7717);
xor U10896 (N_10896,N_7593,N_6968);
xor U10897 (N_10897,N_9032,N_8267);
and U10898 (N_10898,N_7949,N_7292);
and U10899 (N_10899,N_8689,N_8992);
and U10900 (N_10900,N_8800,N_8407);
nand U10901 (N_10901,N_7853,N_7220);
nor U10902 (N_10902,N_7403,N_8173);
xor U10903 (N_10903,N_8641,N_8970);
xor U10904 (N_10904,N_8730,N_8684);
and U10905 (N_10905,N_9270,N_9260);
nand U10906 (N_10906,N_6661,N_6567);
nor U10907 (N_10907,N_8507,N_7193);
or U10908 (N_10908,N_7252,N_8304);
and U10909 (N_10909,N_6280,N_8704);
and U10910 (N_10910,N_6423,N_6534);
xnor U10911 (N_10911,N_7405,N_9183);
and U10912 (N_10912,N_7451,N_7417);
or U10913 (N_10913,N_8773,N_7534);
or U10914 (N_10914,N_7465,N_8359);
and U10915 (N_10915,N_7058,N_7137);
and U10916 (N_10916,N_9210,N_6455);
or U10917 (N_10917,N_6484,N_8524);
xor U10918 (N_10918,N_8248,N_7313);
and U10919 (N_10919,N_6274,N_9102);
and U10920 (N_10920,N_7447,N_7172);
and U10921 (N_10921,N_8073,N_8941);
xnor U10922 (N_10922,N_8374,N_7489);
nor U10923 (N_10923,N_7978,N_8642);
nand U10924 (N_10924,N_6339,N_9242);
and U10925 (N_10925,N_7332,N_8613);
xnor U10926 (N_10926,N_7526,N_6924);
and U10927 (N_10927,N_7265,N_6694);
and U10928 (N_10928,N_7562,N_6352);
nor U10929 (N_10929,N_9262,N_8249);
nor U10930 (N_10930,N_7300,N_8776);
nand U10931 (N_10931,N_7296,N_6373);
and U10932 (N_10932,N_8661,N_6935);
nand U10933 (N_10933,N_7306,N_8271);
or U10934 (N_10934,N_8310,N_6539);
nor U10935 (N_10935,N_8913,N_9133);
nor U10936 (N_10936,N_8148,N_7359);
nand U10937 (N_10937,N_6912,N_7834);
xnor U10938 (N_10938,N_6859,N_6498);
xor U10939 (N_10939,N_8100,N_9088);
xor U10940 (N_10940,N_6670,N_8217);
and U10941 (N_10941,N_7312,N_7203);
or U10942 (N_10942,N_9342,N_6666);
or U10943 (N_10943,N_8029,N_7392);
and U10944 (N_10944,N_7761,N_7384);
or U10945 (N_10945,N_6299,N_8588);
xnor U10946 (N_10946,N_8479,N_6603);
nor U10947 (N_10947,N_7100,N_8728);
xor U10948 (N_10948,N_6825,N_6814);
nor U10949 (N_10949,N_7362,N_7015);
nand U10950 (N_10950,N_6937,N_6676);
nand U10951 (N_10951,N_6572,N_6906);
or U10952 (N_10952,N_6803,N_6373);
and U10953 (N_10953,N_8702,N_7087);
nor U10954 (N_10954,N_6583,N_7076);
nor U10955 (N_10955,N_7120,N_6372);
xor U10956 (N_10956,N_8160,N_8584);
nand U10957 (N_10957,N_7818,N_8115);
and U10958 (N_10958,N_6369,N_7863);
or U10959 (N_10959,N_7959,N_9089);
xnor U10960 (N_10960,N_7614,N_8044);
nand U10961 (N_10961,N_7268,N_8360);
nor U10962 (N_10962,N_7179,N_8360);
nand U10963 (N_10963,N_8731,N_6880);
nand U10964 (N_10964,N_6331,N_8415);
and U10965 (N_10965,N_6267,N_6274);
or U10966 (N_10966,N_8880,N_6772);
and U10967 (N_10967,N_9142,N_7511);
or U10968 (N_10968,N_6478,N_9052);
and U10969 (N_10969,N_9177,N_6596);
nor U10970 (N_10970,N_8662,N_8904);
and U10971 (N_10971,N_6641,N_7291);
nor U10972 (N_10972,N_9140,N_8568);
or U10973 (N_10973,N_6452,N_7424);
or U10974 (N_10974,N_6908,N_7844);
or U10975 (N_10975,N_9134,N_8729);
nor U10976 (N_10976,N_7760,N_8893);
xnor U10977 (N_10977,N_8191,N_6661);
and U10978 (N_10978,N_7791,N_7885);
xor U10979 (N_10979,N_6413,N_6741);
nor U10980 (N_10980,N_7395,N_8457);
nor U10981 (N_10981,N_7497,N_7584);
nor U10982 (N_10982,N_9304,N_8489);
nor U10983 (N_10983,N_8203,N_9147);
and U10984 (N_10984,N_6828,N_8571);
xnor U10985 (N_10985,N_8287,N_8254);
nand U10986 (N_10986,N_7457,N_8170);
or U10987 (N_10987,N_8230,N_6860);
and U10988 (N_10988,N_7178,N_6437);
nor U10989 (N_10989,N_7006,N_6873);
nor U10990 (N_10990,N_8716,N_9021);
or U10991 (N_10991,N_7087,N_6837);
nand U10992 (N_10992,N_8240,N_8685);
and U10993 (N_10993,N_9358,N_7348);
or U10994 (N_10994,N_6837,N_7368);
xnor U10995 (N_10995,N_7685,N_8582);
nor U10996 (N_10996,N_8175,N_7176);
nand U10997 (N_10997,N_7636,N_7352);
nor U10998 (N_10998,N_6257,N_8536);
and U10999 (N_10999,N_7972,N_8663);
and U11000 (N_11000,N_8400,N_8078);
nand U11001 (N_11001,N_9016,N_6316);
nand U11002 (N_11002,N_8593,N_8558);
or U11003 (N_11003,N_8549,N_7196);
nand U11004 (N_11004,N_7723,N_9063);
and U11005 (N_11005,N_8534,N_6670);
nand U11006 (N_11006,N_9355,N_8503);
nor U11007 (N_11007,N_8672,N_9200);
nor U11008 (N_11008,N_9148,N_9346);
or U11009 (N_11009,N_6523,N_8815);
or U11010 (N_11010,N_6936,N_9360);
nor U11011 (N_11011,N_8665,N_7610);
or U11012 (N_11012,N_9187,N_7562);
nand U11013 (N_11013,N_8096,N_8396);
nor U11014 (N_11014,N_8278,N_7386);
and U11015 (N_11015,N_6611,N_6865);
nand U11016 (N_11016,N_9154,N_7072);
or U11017 (N_11017,N_8712,N_7959);
xnor U11018 (N_11018,N_8337,N_8590);
nor U11019 (N_11019,N_7417,N_7596);
nand U11020 (N_11020,N_6953,N_7091);
nand U11021 (N_11021,N_7823,N_6548);
nand U11022 (N_11022,N_7643,N_7828);
and U11023 (N_11023,N_7927,N_6639);
nor U11024 (N_11024,N_8979,N_7803);
nand U11025 (N_11025,N_7535,N_8683);
nor U11026 (N_11026,N_8115,N_7652);
and U11027 (N_11027,N_7784,N_9086);
nor U11028 (N_11028,N_8177,N_6942);
nand U11029 (N_11029,N_7181,N_9020);
nand U11030 (N_11030,N_9066,N_8983);
nor U11031 (N_11031,N_8230,N_9266);
and U11032 (N_11032,N_8605,N_7653);
and U11033 (N_11033,N_7198,N_6435);
or U11034 (N_11034,N_8640,N_8587);
or U11035 (N_11035,N_6456,N_8994);
or U11036 (N_11036,N_7172,N_7243);
nand U11037 (N_11037,N_7197,N_7843);
xor U11038 (N_11038,N_6965,N_6481);
and U11039 (N_11039,N_7022,N_8137);
and U11040 (N_11040,N_6642,N_9069);
or U11041 (N_11041,N_6527,N_7415);
nand U11042 (N_11042,N_9347,N_6859);
nand U11043 (N_11043,N_6771,N_7743);
nor U11044 (N_11044,N_7581,N_8539);
or U11045 (N_11045,N_6929,N_8016);
or U11046 (N_11046,N_6285,N_6751);
and U11047 (N_11047,N_8252,N_7905);
nand U11048 (N_11048,N_8270,N_8547);
nand U11049 (N_11049,N_7406,N_7753);
or U11050 (N_11050,N_7204,N_8196);
nor U11051 (N_11051,N_8154,N_9303);
and U11052 (N_11052,N_7177,N_6724);
or U11053 (N_11053,N_7708,N_7659);
nand U11054 (N_11054,N_6537,N_6347);
nand U11055 (N_11055,N_8765,N_7372);
or U11056 (N_11056,N_9060,N_8937);
xnor U11057 (N_11057,N_7041,N_9312);
nor U11058 (N_11058,N_8303,N_7906);
xnor U11059 (N_11059,N_8767,N_9001);
and U11060 (N_11060,N_6574,N_7545);
nor U11061 (N_11061,N_8435,N_7762);
or U11062 (N_11062,N_8084,N_8847);
or U11063 (N_11063,N_6398,N_8313);
and U11064 (N_11064,N_7199,N_8516);
nand U11065 (N_11065,N_8918,N_9162);
and U11066 (N_11066,N_8859,N_7927);
and U11067 (N_11067,N_8643,N_9141);
and U11068 (N_11068,N_7459,N_7101);
nor U11069 (N_11069,N_9299,N_6347);
nand U11070 (N_11070,N_6544,N_6334);
or U11071 (N_11071,N_7541,N_7741);
nor U11072 (N_11072,N_8083,N_9213);
nand U11073 (N_11073,N_6422,N_8472);
or U11074 (N_11074,N_6810,N_8229);
or U11075 (N_11075,N_6602,N_9071);
nand U11076 (N_11076,N_7119,N_7679);
nand U11077 (N_11077,N_6394,N_8348);
nand U11078 (N_11078,N_7363,N_8182);
or U11079 (N_11079,N_8570,N_8631);
nand U11080 (N_11080,N_6914,N_7674);
nand U11081 (N_11081,N_8164,N_9305);
xnor U11082 (N_11082,N_8499,N_7185);
nor U11083 (N_11083,N_6888,N_6979);
and U11084 (N_11084,N_6938,N_8461);
nor U11085 (N_11085,N_6965,N_8603);
or U11086 (N_11086,N_6411,N_7455);
xnor U11087 (N_11087,N_7404,N_8780);
and U11088 (N_11088,N_7169,N_8798);
or U11089 (N_11089,N_7899,N_8223);
nor U11090 (N_11090,N_8200,N_8950);
or U11091 (N_11091,N_7421,N_7730);
nor U11092 (N_11092,N_8346,N_7826);
nor U11093 (N_11093,N_7153,N_6918);
and U11094 (N_11094,N_9238,N_6844);
xor U11095 (N_11095,N_8039,N_7346);
nand U11096 (N_11096,N_9190,N_8696);
nand U11097 (N_11097,N_8759,N_7858);
nor U11098 (N_11098,N_8070,N_9355);
xor U11099 (N_11099,N_7549,N_9048);
or U11100 (N_11100,N_7921,N_8673);
nand U11101 (N_11101,N_8041,N_6462);
xor U11102 (N_11102,N_7338,N_9198);
nor U11103 (N_11103,N_6996,N_7773);
nor U11104 (N_11104,N_9026,N_8863);
or U11105 (N_11105,N_7385,N_7846);
and U11106 (N_11106,N_7197,N_6530);
nor U11107 (N_11107,N_7722,N_6386);
or U11108 (N_11108,N_7189,N_7258);
or U11109 (N_11109,N_6282,N_8128);
and U11110 (N_11110,N_8534,N_9258);
or U11111 (N_11111,N_6572,N_8502);
or U11112 (N_11112,N_8668,N_8376);
xor U11113 (N_11113,N_7949,N_7071);
and U11114 (N_11114,N_7252,N_8335);
or U11115 (N_11115,N_7659,N_8326);
and U11116 (N_11116,N_6789,N_8196);
and U11117 (N_11117,N_6708,N_6725);
nor U11118 (N_11118,N_9010,N_6491);
nand U11119 (N_11119,N_7893,N_8636);
nand U11120 (N_11120,N_9149,N_8363);
and U11121 (N_11121,N_6743,N_7314);
xnor U11122 (N_11122,N_8701,N_8973);
nor U11123 (N_11123,N_9241,N_7365);
nor U11124 (N_11124,N_7787,N_7136);
and U11125 (N_11125,N_6754,N_8606);
and U11126 (N_11126,N_8878,N_7522);
or U11127 (N_11127,N_6890,N_7798);
nor U11128 (N_11128,N_8014,N_7677);
and U11129 (N_11129,N_8080,N_7788);
or U11130 (N_11130,N_7762,N_6255);
nand U11131 (N_11131,N_8671,N_8039);
xnor U11132 (N_11132,N_7182,N_8748);
or U11133 (N_11133,N_8057,N_8651);
or U11134 (N_11134,N_6440,N_7226);
or U11135 (N_11135,N_7940,N_8562);
xor U11136 (N_11136,N_7425,N_7909);
or U11137 (N_11137,N_6532,N_7642);
nor U11138 (N_11138,N_8695,N_7750);
or U11139 (N_11139,N_7459,N_7730);
nand U11140 (N_11140,N_8442,N_8609);
or U11141 (N_11141,N_8590,N_8822);
nand U11142 (N_11142,N_7378,N_7160);
nand U11143 (N_11143,N_7380,N_7538);
nor U11144 (N_11144,N_9327,N_9344);
nor U11145 (N_11145,N_9026,N_6641);
or U11146 (N_11146,N_7753,N_6415);
or U11147 (N_11147,N_8939,N_8190);
nand U11148 (N_11148,N_9160,N_8394);
nor U11149 (N_11149,N_7443,N_8335);
nand U11150 (N_11150,N_7624,N_8460);
and U11151 (N_11151,N_7835,N_8747);
and U11152 (N_11152,N_6331,N_8717);
nor U11153 (N_11153,N_6609,N_9069);
xnor U11154 (N_11154,N_8742,N_9025);
and U11155 (N_11155,N_8232,N_8908);
and U11156 (N_11156,N_7829,N_7135);
nand U11157 (N_11157,N_7509,N_9041);
nand U11158 (N_11158,N_8627,N_6361);
or U11159 (N_11159,N_6406,N_7905);
and U11160 (N_11160,N_7369,N_9088);
and U11161 (N_11161,N_8472,N_9030);
or U11162 (N_11162,N_8006,N_8151);
nor U11163 (N_11163,N_6738,N_9106);
nor U11164 (N_11164,N_7190,N_7803);
nand U11165 (N_11165,N_7180,N_8826);
nand U11166 (N_11166,N_7034,N_9302);
nand U11167 (N_11167,N_8897,N_7554);
and U11168 (N_11168,N_7652,N_9122);
nand U11169 (N_11169,N_7980,N_6414);
nand U11170 (N_11170,N_7436,N_9248);
nor U11171 (N_11171,N_7773,N_9111);
nand U11172 (N_11172,N_6770,N_8654);
or U11173 (N_11173,N_8612,N_8609);
nor U11174 (N_11174,N_6606,N_8291);
or U11175 (N_11175,N_8620,N_8268);
xnor U11176 (N_11176,N_6354,N_8769);
xor U11177 (N_11177,N_6797,N_8512);
nor U11178 (N_11178,N_8624,N_8146);
nand U11179 (N_11179,N_6926,N_7012);
and U11180 (N_11180,N_7613,N_6608);
and U11181 (N_11181,N_7844,N_8351);
nor U11182 (N_11182,N_7684,N_7905);
or U11183 (N_11183,N_8260,N_8626);
nor U11184 (N_11184,N_8575,N_7123);
or U11185 (N_11185,N_7222,N_8886);
nand U11186 (N_11186,N_7663,N_8991);
xnor U11187 (N_11187,N_6870,N_8279);
and U11188 (N_11188,N_7519,N_7410);
and U11189 (N_11189,N_6997,N_7119);
or U11190 (N_11190,N_6750,N_7310);
xor U11191 (N_11191,N_8580,N_6967);
nor U11192 (N_11192,N_7697,N_8283);
xor U11193 (N_11193,N_6974,N_8000);
xnor U11194 (N_11194,N_8129,N_8523);
or U11195 (N_11195,N_7633,N_8320);
and U11196 (N_11196,N_8600,N_7548);
or U11197 (N_11197,N_9240,N_7235);
or U11198 (N_11198,N_6858,N_8505);
nand U11199 (N_11199,N_6771,N_8386);
and U11200 (N_11200,N_7183,N_7429);
nor U11201 (N_11201,N_7086,N_9097);
nand U11202 (N_11202,N_7026,N_8599);
or U11203 (N_11203,N_7410,N_7994);
nand U11204 (N_11204,N_9034,N_9085);
nor U11205 (N_11205,N_8377,N_9011);
or U11206 (N_11206,N_8228,N_8678);
or U11207 (N_11207,N_8499,N_7820);
nand U11208 (N_11208,N_7366,N_8506);
and U11209 (N_11209,N_7749,N_7638);
xnor U11210 (N_11210,N_9061,N_6733);
nand U11211 (N_11211,N_7360,N_7262);
or U11212 (N_11212,N_8228,N_7349);
nand U11213 (N_11213,N_6371,N_6798);
or U11214 (N_11214,N_8617,N_7958);
or U11215 (N_11215,N_8926,N_8777);
nand U11216 (N_11216,N_7809,N_7878);
or U11217 (N_11217,N_6964,N_6801);
nor U11218 (N_11218,N_6852,N_7606);
nor U11219 (N_11219,N_8711,N_7420);
nor U11220 (N_11220,N_8289,N_8257);
and U11221 (N_11221,N_6542,N_8230);
or U11222 (N_11222,N_8193,N_7154);
nand U11223 (N_11223,N_8638,N_8063);
nand U11224 (N_11224,N_8128,N_6721);
nor U11225 (N_11225,N_7199,N_8768);
nand U11226 (N_11226,N_7319,N_6702);
or U11227 (N_11227,N_8955,N_7869);
nand U11228 (N_11228,N_8346,N_8085);
xor U11229 (N_11229,N_6263,N_8702);
nor U11230 (N_11230,N_6906,N_8144);
or U11231 (N_11231,N_7400,N_8826);
nor U11232 (N_11232,N_7903,N_9263);
or U11233 (N_11233,N_8265,N_6456);
nor U11234 (N_11234,N_6698,N_7849);
nand U11235 (N_11235,N_8962,N_8477);
xor U11236 (N_11236,N_7717,N_8812);
and U11237 (N_11237,N_6545,N_7363);
nor U11238 (N_11238,N_7624,N_6681);
and U11239 (N_11239,N_8599,N_7722);
or U11240 (N_11240,N_7780,N_7608);
nor U11241 (N_11241,N_7397,N_8438);
nand U11242 (N_11242,N_8747,N_9152);
nor U11243 (N_11243,N_8036,N_7607);
or U11244 (N_11244,N_8602,N_7214);
or U11245 (N_11245,N_7505,N_6830);
or U11246 (N_11246,N_7964,N_7932);
xnor U11247 (N_11247,N_9105,N_6664);
and U11248 (N_11248,N_8427,N_8429);
xor U11249 (N_11249,N_8449,N_6788);
or U11250 (N_11250,N_7429,N_9217);
and U11251 (N_11251,N_7064,N_8217);
nor U11252 (N_11252,N_7306,N_7579);
nand U11253 (N_11253,N_8172,N_6532);
nor U11254 (N_11254,N_7896,N_8509);
or U11255 (N_11255,N_8461,N_7122);
or U11256 (N_11256,N_8114,N_6422);
nand U11257 (N_11257,N_7073,N_8563);
or U11258 (N_11258,N_8802,N_9258);
nor U11259 (N_11259,N_7605,N_7472);
nand U11260 (N_11260,N_8416,N_8104);
xor U11261 (N_11261,N_7767,N_7294);
or U11262 (N_11262,N_8850,N_7409);
xnor U11263 (N_11263,N_7511,N_7651);
nand U11264 (N_11264,N_7246,N_8555);
nor U11265 (N_11265,N_7053,N_8515);
nand U11266 (N_11266,N_8206,N_6434);
nand U11267 (N_11267,N_7619,N_8006);
nand U11268 (N_11268,N_6413,N_8567);
and U11269 (N_11269,N_7601,N_6280);
and U11270 (N_11270,N_9045,N_7064);
or U11271 (N_11271,N_7316,N_8654);
xnor U11272 (N_11272,N_6350,N_8925);
or U11273 (N_11273,N_6882,N_7964);
or U11274 (N_11274,N_6307,N_9339);
and U11275 (N_11275,N_7034,N_7990);
and U11276 (N_11276,N_8198,N_6399);
nand U11277 (N_11277,N_7516,N_7848);
and U11278 (N_11278,N_6527,N_7682);
xnor U11279 (N_11279,N_7440,N_8173);
xor U11280 (N_11280,N_7752,N_8854);
or U11281 (N_11281,N_8005,N_6789);
nor U11282 (N_11282,N_8217,N_9349);
and U11283 (N_11283,N_6564,N_9053);
nor U11284 (N_11284,N_8101,N_6935);
or U11285 (N_11285,N_7680,N_7402);
or U11286 (N_11286,N_6964,N_8795);
and U11287 (N_11287,N_7264,N_8126);
nor U11288 (N_11288,N_8490,N_9335);
nand U11289 (N_11289,N_8334,N_8701);
nor U11290 (N_11290,N_8981,N_9007);
and U11291 (N_11291,N_9280,N_8828);
or U11292 (N_11292,N_7676,N_6539);
xnor U11293 (N_11293,N_6893,N_8979);
or U11294 (N_11294,N_7061,N_9209);
nand U11295 (N_11295,N_8042,N_6866);
and U11296 (N_11296,N_7527,N_6276);
nor U11297 (N_11297,N_6689,N_8426);
or U11298 (N_11298,N_7958,N_8706);
or U11299 (N_11299,N_6435,N_6759);
or U11300 (N_11300,N_6742,N_8907);
nor U11301 (N_11301,N_8070,N_8017);
nand U11302 (N_11302,N_8446,N_8473);
and U11303 (N_11303,N_6748,N_7059);
nor U11304 (N_11304,N_8399,N_8923);
and U11305 (N_11305,N_8484,N_6724);
xnor U11306 (N_11306,N_8996,N_6438);
and U11307 (N_11307,N_7203,N_8426);
nand U11308 (N_11308,N_7614,N_8960);
or U11309 (N_11309,N_9127,N_7579);
xnor U11310 (N_11310,N_7117,N_7109);
or U11311 (N_11311,N_9094,N_8966);
nor U11312 (N_11312,N_8659,N_8720);
nor U11313 (N_11313,N_7871,N_8976);
nand U11314 (N_11314,N_7596,N_8910);
nor U11315 (N_11315,N_8053,N_6665);
nor U11316 (N_11316,N_6321,N_6900);
nand U11317 (N_11317,N_7972,N_8118);
and U11318 (N_11318,N_6489,N_6680);
nor U11319 (N_11319,N_9189,N_6590);
and U11320 (N_11320,N_8593,N_6258);
nor U11321 (N_11321,N_6489,N_6479);
nor U11322 (N_11322,N_7836,N_7758);
and U11323 (N_11323,N_7698,N_8888);
xor U11324 (N_11324,N_8899,N_8054);
xnor U11325 (N_11325,N_6796,N_8019);
nand U11326 (N_11326,N_8659,N_8136);
nand U11327 (N_11327,N_6901,N_7368);
or U11328 (N_11328,N_7268,N_6965);
or U11329 (N_11329,N_8693,N_7624);
and U11330 (N_11330,N_8259,N_7928);
nand U11331 (N_11331,N_6487,N_7945);
and U11332 (N_11332,N_9078,N_6940);
xor U11333 (N_11333,N_9269,N_7491);
or U11334 (N_11334,N_6607,N_8599);
nor U11335 (N_11335,N_6393,N_7113);
nor U11336 (N_11336,N_8047,N_8892);
xor U11337 (N_11337,N_7718,N_7253);
and U11338 (N_11338,N_7418,N_8642);
xor U11339 (N_11339,N_6431,N_8705);
or U11340 (N_11340,N_9255,N_8247);
nor U11341 (N_11341,N_8227,N_9304);
nor U11342 (N_11342,N_9037,N_6748);
and U11343 (N_11343,N_8582,N_7617);
nor U11344 (N_11344,N_8332,N_7587);
and U11345 (N_11345,N_7242,N_7633);
xor U11346 (N_11346,N_9233,N_9354);
or U11347 (N_11347,N_8550,N_7646);
or U11348 (N_11348,N_9239,N_6520);
nor U11349 (N_11349,N_8462,N_9280);
nand U11350 (N_11350,N_7030,N_8830);
nor U11351 (N_11351,N_6424,N_8411);
nor U11352 (N_11352,N_7868,N_6548);
nor U11353 (N_11353,N_7673,N_8012);
and U11354 (N_11354,N_6634,N_9118);
or U11355 (N_11355,N_8284,N_8351);
xor U11356 (N_11356,N_9302,N_6554);
or U11357 (N_11357,N_7785,N_9024);
nor U11358 (N_11358,N_6600,N_8336);
nor U11359 (N_11359,N_7324,N_7779);
or U11360 (N_11360,N_8928,N_6945);
nor U11361 (N_11361,N_7122,N_8240);
or U11362 (N_11362,N_8369,N_9026);
xnor U11363 (N_11363,N_6814,N_9131);
nand U11364 (N_11364,N_7281,N_8241);
or U11365 (N_11365,N_7631,N_8511);
xor U11366 (N_11366,N_8063,N_7878);
or U11367 (N_11367,N_7231,N_7731);
or U11368 (N_11368,N_8453,N_8532);
and U11369 (N_11369,N_6394,N_6447);
or U11370 (N_11370,N_7944,N_6415);
or U11371 (N_11371,N_7609,N_7595);
and U11372 (N_11372,N_6346,N_8950);
nand U11373 (N_11373,N_6654,N_7530);
nor U11374 (N_11374,N_8128,N_8225);
nor U11375 (N_11375,N_7524,N_6817);
nand U11376 (N_11376,N_8119,N_9328);
nor U11377 (N_11377,N_8730,N_7245);
and U11378 (N_11378,N_7081,N_8450);
nand U11379 (N_11379,N_6618,N_6439);
and U11380 (N_11380,N_7314,N_8104);
nand U11381 (N_11381,N_8320,N_8252);
nor U11382 (N_11382,N_7207,N_7672);
and U11383 (N_11383,N_6526,N_6300);
nor U11384 (N_11384,N_7105,N_8977);
nand U11385 (N_11385,N_7057,N_8441);
xnor U11386 (N_11386,N_8460,N_7228);
nor U11387 (N_11387,N_7680,N_8980);
nor U11388 (N_11388,N_8359,N_7986);
or U11389 (N_11389,N_7992,N_7911);
or U11390 (N_11390,N_8242,N_8798);
or U11391 (N_11391,N_7859,N_6907);
and U11392 (N_11392,N_8620,N_8407);
or U11393 (N_11393,N_8065,N_7264);
xnor U11394 (N_11394,N_9084,N_7482);
nor U11395 (N_11395,N_8342,N_9337);
nand U11396 (N_11396,N_7544,N_6688);
or U11397 (N_11397,N_6955,N_8307);
nand U11398 (N_11398,N_6286,N_8428);
nand U11399 (N_11399,N_8028,N_6692);
nor U11400 (N_11400,N_8561,N_9353);
nand U11401 (N_11401,N_9274,N_6342);
and U11402 (N_11402,N_7347,N_8293);
nor U11403 (N_11403,N_8986,N_6723);
or U11404 (N_11404,N_6664,N_8515);
nand U11405 (N_11405,N_6657,N_8527);
nor U11406 (N_11406,N_8486,N_8417);
nand U11407 (N_11407,N_6484,N_7614);
nand U11408 (N_11408,N_6647,N_7338);
xnor U11409 (N_11409,N_6675,N_8673);
and U11410 (N_11410,N_6735,N_7766);
and U11411 (N_11411,N_8069,N_6630);
nor U11412 (N_11412,N_7682,N_8628);
nand U11413 (N_11413,N_8357,N_9029);
nor U11414 (N_11414,N_8773,N_8624);
and U11415 (N_11415,N_8083,N_7443);
nor U11416 (N_11416,N_9279,N_6409);
or U11417 (N_11417,N_7646,N_8948);
and U11418 (N_11418,N_7029,N_8985);
or U11419 (N_11419,N_8452,N_9063);
or U11420 (N_11420,N_6937,N_7256);
nand U11421 (N_11421,N_6441,N_8501);
nand U11422 (N_11422,N_6650,N_7960);
and U11423 (N_11423,N_6723,N_8413);
and U11424 (N_11424,N_7557,N_9306);
or U11425 (N_11425,N_9191,N_7455);
nor U11426 (N_11426,N_8558,N_8443);
nor U11427 (N_11427,N_8197,N_6921);
or U11428 (N_11428,N_9009,N_9309);
or U11429 (N_11429,N_7066,N_7904);
and U11430 (N_11430,N_6632,N_8198);
nor U11431 (N_11431,N_7851,N_9276);
or U11432 (N_11432,N_7474,N_9115);
or U11433 (N_11433,N_8536,N_6681);
or U11434 (N_11434,N_7133,N_7139);
nor U11435 (N_11435,N_8664,N_8444);
or U11436 (N_11436,N_7939,N_8978);
nor U11437 (N_11437,N_9269,N_8570);
or U11438 (N_11438,N_7747,N_8037);
nand U11439 (N_11439,N_8347,N_7022);
or U11440 (N_11440,N_7092,N_6698);
nor U11441 (N_11441,N_8629,N_7194);
nand U11442 (N_11442,N_8433,N_6854);
xnor U11443 (N_11443,N_6895,N_8905);
and U11444 (N_11444,N_8360,N_7971);
nor U11445 (N_11445,N_9358,N_9329);
nand U11446 (N_11446,N_6881,N_7134);
or U11447 (N_11447,N_7493,N_8446);
nor U11448 (N_11448,N_7631,N_6558);
nand U11449 (N_11449,N_6445,N_6485);
nand U11450 (N_11450,N_6278,N_8046);
nor U11451 (N_11451,N_8570,N_6753);
and U11452 (N_11452,N_7164,N_8917);
and U11453 (N_11453,N_8175,N_7734);
nor U11454 (N_11454,N_6598,N_7418);
nor U11455 (N_11455,N_7210,N_7212);
and U11456 (N_11456,N_7834,N_8438);
nand U11457 (N_11457,N_7186,N_8474);
nor U11458 (N_11458,N_7779,N_7868);
xor U11459 (N_11459,N_6894,N_7789);
and U11460 (N_11460,N_7885,N_6875);
nor U11461 (N_11461,N_8279,N_7981);
nand U11462 (N_11462,N_8345,N_7573);
and U11463 (N_11463,N_8272,N_7742);
nor U11464 (N_11464,N_6474,N_7462);
and U11465 (N_11465,N_8066,N_8756);
and U11466 (N_11466,N_8343,N_7804);
nand U11467 (N_11467,N_6283,N_7304);
or U11468 (N_11468,N_7329,N_6842);
nand U11469 (N_11469,N_9373,N_8213);
nor U11470 (N_11470,N_8675,N_7642);
nand U11471 (N_11471,N_7253,N_6938);
or U11472 (N_11472,N_8433,N_7756);
nand U11473 (N_11473,N_6323,N_6745);
nand U11474 (N_11474,N_8671,N_7534);
and U11475 (N_11475,N_6905,N_6298);
nor U11476 (N_11476,N_8139,N_6716);
and U11477 (N_11477,N_9359,N_8964);
and U11478 (N_11478,N_6401,N_8141);
and U11479 (N_11479,N_8606,N_6504);
or U11480 (N_11480,N_7629,N_7919);
xnor U11481 (N_11481,N_9349,N_8740);
xor U11482 (N_11482,N_6288,N_9312);
xnor U11483 (N_11483,N_7961,N_7017);
nor U11484 (N_11484,N_8302,N_8380);
xnor U11485 (N_11485,N_8742,N_7456);
and U11486 (N_11486,N_8218,N_7005);
nor U11487 (N_11487,N_7538,N_6488);
nand U11488 (N_11488,N_7350,N_6928);
or U11489 (N_11489,N_6740,N_7424);
nand U11490 (N_11490,N_7280,N_6278);
or U11491 (N_11491,N_7880,N_7388);
and U11492 (N_11492,N_9220,N_6536);
or U11493 (N_11493,N_7405,N_7683);
nor U11494 (N_11494,N_8871,N_7671);
or U11495 (N_11495,N_7979,N_8155);
or U11496 (N_11496,N_8790,N_7556);
or U11497 (N_11497,N_8090,N_6923);
and U11498 (N_11498,N_7393,N_7420);
nor U11499 (N_11499,N_7925,N_7973);
nor U11500 (N_11500,N_9354,N_7748);
and U11501 (N_11501,N_7416,N_8991);
nand U11502 (N_11502,N_9128,N_6809);
or U11503 (N_11503,N_8233,N_8516);
or U11504 (N_11504,N_6262,N_7277);
or U11505 (N_11505,N_6787,N_7886);
and U11506 (N_11506,N_6459,N_9261);
or U11507 (N_11507,N_8367,N_7117);
and U11508 (N_11508,N_7260,N_9115);
nand U11509 (N_11509,N_8510,N_8245);
xnor U11510 (N_11510,N_7766,N_8904);
or U11511 (N_11511,N_6631,N_8118);
nand U11512 (N_11512,N_8642,N_7354);
xnor U11513 (N_11513,N_8615,N_9215);
or U11514 (N_11514,N_7155,N_7393);
and U11515 (N_11515,N_7702,N_9284);
and U11516 (N_11516,N_7590,N_8112);
nor U11517 (N_11517,N_7822,N_9018);
nand U11518 (N_11518,N_8333,N_7252);
and U11519 (N_11519,N_7152,N_8553);
and U11520 (N_11520,N_7240,N_6765);
and U11521 (N_11521,N_6846,N_8760);
and U11522 (N_11522,N_6788,N_7724);
nand U11523 (N_11523,N_8721,N_8207);
and U11524 (N_11524,N_8722,N_9281);
nand U11525 (N_11525,N_7130,N_7981);
and U11526 (N_11526,N_6991,N_7910);
xor U11527 (N_11527,N_8854,N_8610);
nand U11528 (N_11528,N_7969,N_8771);
or U11529 (N_11529,N_8662,N_9223);
nand U11530 (N_11530,N_6639,N_7271);
nor U11531 (N_11531,N_8529,N_7372);
or U11532 (N_11532,N_6850,N_8643);
and U11533 (N_11533,N_8583,N_6430);
nand U11534 (N_11534,N_7939,N_6339);
nand U11535 (N_11535,N_6498,N_6370);
and U11536 (N_11536,N_7691,N_7423);
nand U11537 (N_11537,N_7222,N_7963);
and U11538 (N_11538,N_7221,N_7032);
or U11539 (N_11539,N_8491,N_9329);
xor U11540 (N_11540,N_8717,N_9063);
nand U11541 (N_11541,N_6938,N_7537);
nand U11542 (N_11542,N_8118,N_9341);
or U11543 (N_11543,N_8408,N_6826);
nor U11544 (N_11544,N_9261,N_7165);
and U11545 (N_11545,N_6446,N_6869);
xnor U11546 (N_11546,N_7898,N_6419);
nand U11547 (N_11547,N_9062,N_6582);
nand U11548 (N_11548,N_8656,N_6512);
xor U11549 (N_11549,N_6250,N_9253);
xnor U11550 (N_11550,N_6970,N_6955);
nand U11551 (N_11551,N_6507,N_8633);
nand U11552 (N_11552,N_6499,N_8782);
or U11553 (N_11553,N_8971,N_6939);
or U11554 (N_11554,N_8922,N_6810);
or U11555 (N_11555,N_8348,N_7335);
or U11556 (N_11556,N_8881,N_6657);
nor U11557 (N_11557,N_7372,N_7995);
nand U11558 (N_11558,N_6883,N_8532);
nand U11559 (N_11559,N_8638,N_7761);
or U11560 (N_11560,N_7530,N_8876);
nand U11561 (N_11561,N_6505,N_7033);
nor U11562 (N_11562,N_7518,N_7036);
nor U11563 (N_11563,N_8071,N_7294);
nand U11564 (N_11564,N_8173,N_7531);
or U11565 (N_11565,N_8425,N_7400);
nand U11566 (N_11566,N_7876,N_7257);
nor U11567 (N_11567,N_6283,N_8294);
and U11568 (N_11568,N_8173,N_7011);
nand U11569 (N_11569,N_8331,N_8826);
and U11570 (N_11570,N_8076,N_7576);
or U11571 (N_11571,N_8810,N_8417);
and U11572 (N_11572,N_6789,N_7970);
and U11573 (N_11573,N_6652,N_7385);
nor U11574 (N_11574,N_6905,N_8043);
or U11575 (N_11575,N_8242,N_6355);
nor U11576 (N_11576,N_8259,N_8130);
or U11577 (N_11577,N_6784,N_8255);
nand U11578 (N_11578,N_8786,N_9327);
nor U11579 (N_11579,N_7660,N_6659);
nor U11580 (N_11580,N_6553,N_7258);
nor U11581 (N_11581,N_7966,N_8719);
and U11582 (N_11582,N_7093,N_7081);
or U11583 (N_11583,N_9241,N_7264);
or U11584 (N_11584,N_6442,N_6267);
nor U11585 (N_11585,N_6812,N_9142);
nor U11586 (N_11586,N_7057,N_6332);
nor U11587 (N_11587,N_6797,N_8163);
xor U11588 (N_11588,N_7292,N_8531);
nand U11589 (N_11589,N_8544,N_7364);
nor U11590 (N_11590,N_7499,N_7283);
and U11591 (N_11591,N_9344,N_6512);
and U11592 (N_11592,N_7216,N_9361);
or U11593 (N_11593,N_6758,N_6543);
or U11594 (N_11594,N_8445,N_6388);
xor U11595 (N_11595,N_7982,N_8614);
nor U11596 (N_11596,N_8809,N_7889);
nor U11597 (N_11597,N_6795,N_7427);
nand U11598 (N_11598,N_7513,N_6851);
xnor U11599 (N_11599,N_9250,N_8416);
or U11600 (N_11600,N_6659,N_9369);
nor U11601 (N_11601,N_9033,N_8044);
nand U11602 (N_11602,N_7675,N_6315);
nor U11603 (N_11603,N_7101,N_8277);
nand U11604 (N_11604,N_6592,N_6827);
nor U11605 (N_11605,N_7743,N_8179);
and U11606 (N_11606,N_6618,N_7749);
nand U11607 (N_11607,N_6692,N_9075);
nor U11608 (N_11608,N_8815,N_8827);
or U11609 (N_11609,N_6844,N_7013);
nor U11610 (N_11610,N_6720,N_8193);
and U11611 (N_11611,N_8573,N_7575);
and U11612 (N_11612,N_9365,N_8234);
and U11613 (N_11613,N_7129,N_8332);
or U11614 (N_11614,N_7039,N_6669);
or U11615 (N_11615,N_8502,N_7012);
or U11616 (N_11616,N_7638,N_8116);
nor U11617 (N_11617,N_6714,N_7880);
or U11618 (N_11618,N_7063,N_6805);
and U11619 (N_11619,N_7439,N_8461);
and U11620 (N_11620,N_8560,N_8787);
nor U11621 (N_11621,N_6983,N_7343);
nand U11622 (N_11622,N_8619,N_8746);
nor U11623 (N_11623,N_9181,N_8694);
nand U11624 (N_11624,N_8873,N_6805);
nand U11625 (N_11625,N_9160,N_9229);
nor U11626 (N_11626,N_6800,N_8540);
nor U11627 (N_11627,N_7551,N_6744);
nand U11628 (N_11628,N_8653,N_8454);
nor U11629 (N_11629,N_6391,N_8424);
and U11630 (N_11630,N_7760,N_8028);
or U11631 (N_11631,N_7791,N_6938);
and U11632 (N_11632,N_6508,N_8757);
nand U11633 (N_11633,N_7612,N_6934);
and U11634 (N_11634,N_7116,N_7935);
nand U11635 (N_11635,N_6616,N_6741);
xor U11636 (N_11636,N_6502,N_7676);
xnor U11637 (N_11637,N_9017,N_6603);
nand U11638 (N_11638,N_7306,N_6293);
or U11639 (N_11639,N_8999,N_8359);
nor U11640 (N_11640,N_8615,N_8599);
nor U11641 (N_11641,N_6947,N_6407);
nand U11642 (N_11642,N_8616,N_7311);
and U11643 (N_11643,N_6961,N_7417);
or U11644 (N_11644,N_6960,N_6637);
nand U11645 (N_11645,N_6428,N_8656);
xnor U11646 (N_11646,N_7530,N_8843);
nand U11647 (N_11647,N_7521,N_6979);
and U11648 (N_11648,N_6450,N_6319);
nand U11649 (N_11649,N_7908,N_8651);
and U11650 (N_11650,N_8750,N_7164);
nand U11651 (N_11651,N_6454,N_8059);
and U11652 (N_11652,N_7669,N_7169);
or U11653 (N_11653,N_8624,N_9237);
nand U11654 (N_11654,N_8484,N_7399);
nor U11655 (N_11655,N_7741,N_6807);
nand U11656 (N_11656,N_8311,N_9216);
and U11657 (N_11657,N_8990,N_6759);
and U11658 (N_11658,N_6571,N_7384);
nor U11659 (N_11659,N_7056,N_7816);
nor U11660 (N_11660,N_8604,N_7808);
nor U11661 (N_11661,N_8073,N_7234);
nor U11662 (N_11662,N_8665,N_7237);
xnor U11663 (N_11663,N_7835,N_8021);
or U11664 (N_11664,N_9235,N_6714);
nor U11665 (N_11665,N_6749,N_8048);
nand U11666 (N_11666,N_9202,N_7294);
xnor U11667 (N_11667,N_9148,N_7626);
nand U11668 (N_11668,N_7739,N_6682);
nand U11669 (N_11669,N_7454,N_6519);
nand U11670 (N_11670,N_9090,N_7914);
and U11671 (N_11671,N_8789,N_7308);
nand U11672 (N_11672,N_7432,N_6412);
xor U11673 (N_11673,N_6688,N_9099);
and U11674 (N_11674,N_8269,N_7313);
xnor U11675 (N_11675,N_6981,N_8073);
nand U11676 (N_11676,N_8909,N_9001);
nand U11677 (N_11677,N_8610,N_9066);
xnor U11678 (N_11678,N_9195,N_8632);
or U11679 (N_11679,N_8301,N_8546);
and U11680 (N_11680,N_8360,N_7993);
or U11681 (N_11681,N_6807,N_8500);
nor U11682 (N_11682,N_6697,N_8868);
nor U11683 (N_11683,N_8138,N_8496);
nor U11684 (N_11684,N_8059,N_9193);
and U11685 (N_11685,N_6276,N_8598);
and U11686 (N_11686,N_6863,N_8272);
nand U11687 (N_11687,N_6838,N_8841);
nand U11688 (N_11688,N_6310,N_6915);
or U11689 (N_11689,N_7658,N_8646);
and U11690 (N_11690,N_7594,N_6731);
nand U11691 (N_11691,N_6735,N_7249);
nor U11692 (N_11692,N_7761,N_9278);
xor U11693 (N_11693,N_7967,N_7487);
xor U11694 (N_11694,N_7328,N_7471);
xnor U11695 (N_11695,N_8591,N_7325);
nand U11696 (N_11696,N_6383,N_7449);
and U11697 (N_11697,N_7463,N_7288);
nand U11698 (N_11698,N_7933,N_7544);
nand U11699 (N_11699,N_9246,N_7232);
nand U11700 (N_11700,N_7928,N_8049);
nand U11701 (N_11701,N_6350,N_8915);
xor U11702 (N_11702,N_6874,N_8742);
or U11703 (N_11703,N_7840,N_8815);
xor U11704 (N_11704,N_7026,N_8112);
and U11705 (N_11705,N_7102,N_6299);
and U11706 (N_11706,N_7154,N_7386);
nor U11707 (N_11707,N_7920,N_8314);
and U11708 (N_11708,N_6990,N_6729);
nor U11709 (N_11709,N_7471,N_6791);
or U11710 (N_11710,N_9282,N_9244);
or U11711 (N_11711,N_8927,N_6942);
or U11712 (N_11712,N_8860,N_8122);
xor U11713 (N_11713,N_6423,N_6722);
nand U11714 (N_11714,N_7284,N_7267);
nor U11715 (N_11715,N_9057,N_6625);
nand U11716 (N_11716,N_6973,N_6537);
and U11717 (N_11717,N_6835,N_8111);
and U11718 (N_11718,N_6414,N_7353);
nor U11719 (N_11719,N_6789,N_8467);
or U11720 (N_11720,N_8688,N_9077);
nand U11721 (N_11721,N_9256,N_9114);
and U11722 (N_11722,N_6431,N_7395);
nand U11723 (N_11723,N_6333,N_6574);
and U11724 (N_11724,N_8162,N_8831);
or U11725 (N_11725,N_7993,N_8537);
nand U11726 (N_11726,N_6523,N_6274);
nand U11727 (N_11727,N_6704,N_9282);
and U11728 (N_11728,N_8396,N_8036);
nor U11729 (N_11729,N_6952,N_6877);
nand U11730 (N_11730,N_7030,N_7235);
and U11731 (N_11731,N_7236,N_8943);
or U11732 (N_11732,N_6743,N_8038);
nor U11733 (N_11733,N_6867,N_8537);
nand U11734 (N_11734,N_8695,N_7229);
and U11735 (N_11735,N_9187,N_8242);
or U11736 (N_11736,N_9304,N_9261);
xor U11737 (N_11737,N_6836,N_6523);
nand U11738 (N_11738,N_6414,N_9201);
or U11739 (N_11739,N_8759,N_7394);
nand U11740 (N_11740,N_6424,N_9051);
or U11741 (N_11741,N_7906,N_7012);
xor U11742 (N_11742,N_8273,N_8789);
and U11743 (N_11743,N_7618,N_6369);
nand U11744 (N_11744,N_9333,N_8423);
and U11745 (N_11745,N_8208,N_9005);
and U11746 (N_11746,N_7863,N_8434);
nand U11747 (N_11747,N_7675,N_9182);
or U11748 (N_11748,N_6888,N_7869);
nor U11749 (N_11749,N_6278,N_8467);
nand U11750 (N_11750,N_6295,N_6468);
nor U11751 (N_11751,N_7956,N_7552);
nand U11752 (N_11752,N_8334,N_6716);
or U11753 (N_11753,N_6779,N_7813);
or U11754 (N_11754,N_7914,N_8976);
nand U11755 (N_11755,N_7002,N_9086);
and U11756 (N_11756,N_7358,N_6257);
or U11757 (N_11757,N_6650,N_7292);
and U11758 (N_11758,N_9040,N_8395);
and U11759 (N_11759,N_8677,N_7102);
or U11760 (N_11760,N_9105,N_8233);
nor U11761 (N_11761,N_6446,N_6852);
xor U11762 (N_11762,N_9221,N_8114);
nor U11763 (N_11763,N_9308,N_6566);
or U11764 (N_11764,N_8434,N_7281);
or U11765 (N_11765,N_7088,N_7758);
and U11766 (N_11766,N_7731,N_6763);
nor U11767 (N_11767,N_8739,N_7950);
and U11768 (N_11768,N_8240,N_8132);
nor U11769 (N_11769,N_7150,N_9186);
nand U11770 (N_11770,N_8448,N_7472);
xor U11771 (N_11771,N_7220,N_8407);
nand U11772 (N_11772,N_8810,N_8452);
or U11773 (N_11773,N_7759,N_7371);
nor U11774 (N_11774,N_9056,N_7482);
nand U11775 (N_11775,N_6778,N_7932);
nor U11776 (N_11776,N_7854,N_9050);
and U11777 (N_11777,N_8951,N_8911);
nor U11778 (N_11778,N_7809,N_8516);
and U11779 (N_11779,N_6583,N_7707);
nor U11780 (N_11780,N_6827,N_8276);
or U11781 (N_11781,N_7891,N_6310);
and U11782 (N_11782,N_6507,N_6762);
nor U11783 (N_11783,N_7854,N_8761);
nand U11784 (N_11784,N_9212,N_8745);
nor U11785 (N_11785,N_8016,N_6259);
nor U11786 (N_11786,N_7870,N_8910);
nor U11787 (N_11787,N_7956,N_8716);
or U11788 (N_11788,N_7630,N_8538);
nand U11789 (N_11789,N_7636,N_7281);
and U11790 (N_11790,N_6712,N_6422);
or U11791 (N_11791,N_8239,N_7548);
xnor U11792 (N_11792,N_9061,N_7427);
nor U11793 (N_11793,N_7135,N_8814);
nor U11794 (N_11794,N_8082,N_6592);
and U11795 (N_11795,N_7730,N_9309);
and U11796 (N_11796,N_6367,N_6386);
nor U11797 (N_11797,N_7409,N_7088);
nand U11798 (N_11798,N_7238,N_9092);
nand U11799 (N_11799,N_8302,N_9313);
or U11800 (N_11800,N_7356,N_7750);
nor U11801 (N_11801,N_9006,N_8424);
and U11802 (N_11802,N_8857,N_8183);
nor U11803 (N_11803,N_7119,N_6623);
nor U11804 (N_11804,N_8890,N_8459);
or U11805 (N_11805,N_6844,N_8739);
or U11806 (N_11806,N_7551,N_8303);
nand U11807 (N_11807,N_9341,N_8847);
nor U11808 (N_11808,N_8553,N_6534);
or U11809 (N_11809,N_7375,N_7187);
and U11810 (N_11810,N_8404,N_8715);
xnor U11811 (N_11811,N_8767,N_6870);
or U11812 (N_11812,N_7242,N_7406);
xnor U11813 (N_11813,N_6376,N_9278);
nor U11814 (N_11814,N_7442,N_8553);
nor U11815 (N_11815,N_7461,N_8750);
and U11816 (N_11816,N_7661,N_8529);
nor U11817 (N_11817,N_8225,N_7607);
nand U11818 (N_11818,N_7782,N_7146);
and U11819 (N_11819,N_7700,N_8188);
nor U11820 (N_11820,N_6714,N_7173);
and U11821 (N_11821,N_8576,N_6536);
nor U11822 (N_11822,N_8638,N_9304);
and U11823 (N_11823,N_7391,N_7685);
xnor U11824 (N_11824,N_6814,N_6842);
and U11825 (N_11825,N_8739,N_9123);
or U11826 (N_11826,N_7926,N_8375);
xnor U11827 (N_11827,N_8894,N_7963);
nand U11828 (N_11828,N_9033,N_8197);
and U11829 (N_11829,N_8048,N_8532);
or U11830 (N_11830,N_7427,N_7812);
and U11831 (N_11831,N_7267,N_7925);
nand U11832 (N_11832,N_8708,N_7552);
nand U11833 (N_11833,N_6670,N_8365);
xor U11834 (N_11834,N_6607,N_7331);
nor U11835 (N_11835,N_8494,N_8567);
and U11836 (N_11836,N_7349,N_6741);
or U11837 (N_11837,N_6358,N_7420);
and U11838 (N_11838,N_7459,N_9170);
nor U11839 (N_11839,N_9281,N_6462);
xnor U11840 (N_11840,N_8723,N_9318);
and U11841 (N_11841,N_8118,N_7865);
nand U11842 (N_11842,N_8753,N_8194);
and U11843 (N_11843,N_8509,N_6631);
and U11844 (N_11844,N_8378,N_7811);
or U11845 (N_11845,N_7573,N_8845);
xnor U11846 (N_11846,N_6488,N_6399);
nand U11847 (N_11847,N_8367,N_6573);
or U11848 (N_11848,N_8722,N_6399);
or U11849 (N_11849,N_7815,N_8427);
and U11850 (N_11850,N_7071,N_7280);
nor U11851 (N_11851,N_8719,N_6775);
and U11852 (N_11852,N_8402,N_8450);
nand U11853 (N_11853,N_8405,N_7499);
nand U11854 (N_11854,N_7504,N_6728);
nand U11855 (N_11855,N_8803,N_8623);
nand U11856 (N_11856,N_6909,N_7039);
and U11857 (N_11857,N_7019,N_7020);
nor U11858 (N_11858,N_7613,N_8452);
or U11859 (N_11859,N_6472,N_9244);
nor U11860 (N_11860,N_8844,N_8337);
or U11861 (N_11861,N_7530,N_9272);
nand U11862 (N_11862,N_7333,N_7250);
and U11863 (N_11863,N_8217,N_7354);
and U11864 (N_11864,N_8271,N_8605);
nand U11865 (N_11865,N_7484,N_6284);
nand U11866 (N_11866,N_8389,N_8924);
or U11867 (N_11867,N_7228,N_8701);
or U11868 (N_11868,N_8034,N_8979);
or U11869 (N_11869,N_7971,N_7514);
or U11870 (N_11870,N_7994,N_7254);
or U11871 (N_11871,N_8837,N_6593);
nand U11872 (N_11872,N_9023,N_8180);
nand U11873 (N_11873,N_7220,N_7470);
nor U11874 (N_11874,N_9171,N_6616);
nand U11875 (N_11875,N_7510,N_6376);
and U11876 (N_11876,N_6522,N_7496);
xor U11877 (N_11877,N_8035,N_8447);
nor U11878 (N_11878,N_6446,N_9239);
and U11879 (N_11879,N_7597,N_7377);
nand U11880 (N_11880,N_6615,N_9267);
nor U11881 (N_11881,N_8949,N_8802);
nor U11882 (N_11882,N_7913,N_8795);
nand U11883 (N_11883,N_6302,N_8393);
and U11884 (N_11884,N_6872,N_6499);
nand U11885 (N_11885,N_6254,N_7386);
nor U11886 (N_11886,N_8103,N_8937);
and U11887 (N_11887,N_8436,N_8952);
nor U11888 (N_11888,N_8293,N_8363);
nor U11889 (N_11889,N_6811,N_8856);
and U11890 (N_11890,N_8274,N_6956);
and U11891 (N_11891,N_8352,N_7366);
nor U11892 (N_11892,N_8643,N_9133);
nand U11893 (N_11893,N_8432,N_6775);
and U11894 (N_11894,N_9361,N_9241);
or U11895 (N_11895,N_8900,N_8732);
nor U11896 (N_11896,N_8939,N_7691);
and U11897 (N_11897,N_7703,N_7618);
nand U11898 (N_11898,N_8308,N_6659);
nand U11899 (N_11899,N_6605,N_7337);
nor U11900 (N_11900,N_6816,N_7200);
xnor U11901 (N_11901,N_9283,N_7621);
and U11902 (N_11902,N_8916,N_6297);
nand U11903 (N_11903,N_8256,N_6833);
nor U11904 (N_11904,N_6544,N_8832);
nand U11905 (N_11905,N_7297,N_8495);
nor U11906 (N_11906,N_9026,N_7576);
and U11907 (N_11907,N_7625,N_6992);
nor U11908 (N_11908,N_7616,N_8896);
nor U11909 (N_11909,N_6626,N_6630);
and U11910 (N_11910,N_7685,N_8024);
or U11911 (N_11911,N_6966,N_8962);
or U11912 (N_11912,N_6374,N_7804);
nor U11913 (N_11913,N_6524,N_8262);
nor U11914 (N_11914,N_8200,N_8239);
or U11915 (N_11915,N_8602,N_9314);
and U11916 (N_11916,N_8609,N_6778);
nor U11917 (N_11917,N_8878,N_6409);
nand U11918 (N_11918,N_7153,N_8000);
or U11919 (N_11919,N_8525,N_6673);
nand U11920 (N_11920,N_6719,N_6553);
nor U11921 (N_11921,N_7868,N_6709);
nand U11922 (N_11922,N_8320,N_8520);
nand U11923 (N_11923,N_7570,N_7974);
and U11924 (N_11924,N_7737,N_9132);
xor U11925 (N_11925,N_7154,N_8888);
and U11926 (N_11926,N_9048,N_9197);
xor U11927 (N_11927,N_8861,N_7637);
and U11928 (N_11928,N_6331,N_8194);
nor U11929 (N_11929,N_6455,N_6872);
nor U11930 (N_11930,N_7863,N_7479);
xnor U11931 (N_11931,N_6523,N_8437);
or U11932 (N_11932,N_8702,N_7256);
nor U11933 (N_11933,N_6252,N_7926);
or U11934 (N_11934,N_6481,N_6500);
or U11935 (N_11935,N_8511,N_7738);
nand U11936 (N_11936,N_8261,N_8185);
nor U11937 (N_11937,N_7140,N_8091);
nand U11938 (N_11938,N_8794,N_7156);
nor U11939 (N_11939,N_9111,N_6772);
or U11940 (N_11940,N_9072,N_9361);
xnor U11941 (N_11941,N_6337,N_9012);
and U11942 (N_11942,N_6643,N_7723);
and U11943 (N_11943,N_9346,N_6950);
xnor U11944 (N_11944,N_8272,N_8319);
nor U11945 (N_11945,N_7177,N_6937);
or U11946 (N_11946,N_6783,N_7936);
nand U11947 (N_11947,N_9345,N_9253);
and U11948 (N_11948,N_8854,N_6614);
xor U11949 (N_11949,N_7572,N_8209);
nor U11950 (N_11950,N_6689,N_8401);
nor U11951 (N_11951,N_7472,N_8790);
nor U11952 (N_11952,N_7776,N_9005);
nand U11953 (N_11953,N_6654,N_8613);
or U11954 (N_11954,N_8364,N_8467);
nand U11955 (N_11955,N_6987,N_8679);
xor U11956 (N_11956,N_9146,N_8312);
or U11957 (N_11957,N_7328,N_9345);
nor U11958 (N_11958,N_8717,N_9105);
or U11959 (N_11959,N_8923,N_7899);
and U11960 (N_11960,N_7486,N_9166);
nand U11961 (N_11961,N_7044,N_7535);
or U11962 (N_11962,N_6866,N_8268);
and U11963 (N_11963,N_7091,N_6307);
and U11964 (N_11964,N_6257,N_9202);
or U11965 (N_11965,N_7766,N_7791);
and U11966 (N_11966,N_8467,N_6950);
nand U11967 (N_11967,N_7511,N_9332);
nor U11968 (N_11968,N_6678,N_7308);
or U11969 (N_11969,N_7565,N_6374);
or U11970 (N_11970,N_8653,N_7394);
and U11971 (N_11971,N_7360,N_9139);
and U11972 (N_11972,N_7154,N_6981);
nand U11973 (N_11973,N_8001,N_6943);
xor U11974 (N_11974,N_7414,N_7374);
and U11975 (N_11975,N_7554,N_9283);
or U11976 (N_11976,N_8185,N_7415);
and U11977 (N_11977,N_8407,N_7323);
and U11978 (N_11978,N_8079,N_7687);
nor U11979 (N_11979,N_8734,N_7446);
xnor U11980 (N_11980,N_8291,N_6722);
nand U11981 (N_11981,N_7019,N_7458);
nor U11982 (N_11982,N_6509,N_6583);
nand U11983 (N_11983,N_7586,N_8572);
nor U11984 (N_11984,N_8303,N_7180);
xnor U11985 (N_11985,N_8696,N_7630);
and U11986 (N_11986,N_7623,N_8027);
nand U11987 (N_11987,N_8096,N_7076);
and U11988 (N_11988,N_7857,N_7136);
nand U11989 (N_11989,N_6975,N_6524);
and U11990 (N_11990,N_8059,N_7343);
or U11991 (N_11991,N_7191,N_9312);
nand U11992 (N_11992,N_9177,N_7283);
or U11993 (N_11993,N_6695,N_7709);
nand U11994 (N_11994,N_7877,N_8941);
and U11995 (N_11995,N_8493,N_8063);
or U11996 (N_11996,N_8125,N_8538);
xnor U11997 (N_11997,N_6688,N_7608);
or U11998 (N_11998,N_7448,N_8905);
and U11999 (N_11999,N_9266,N_8037);
nor U12000 (N_12000,N_6290,N_8787);
nor U12001 (N_12001,N_8757,N_6424);
nor U12002 (N_12002,N_6548,N_8462);
and U12003 (N_12003,N_8304,N_8250);
nand U12004 (N_12004,N_6431,N_6386);
nor U12005 (N_12005,N_6661,N_8490);
nand U12006 (N_12006,N_7649,N_8354);
nor U12007 (N_12007,N_6852,N_7152);
nor U12008 (N_12008,N_8702,N_8654);
and U12009 (N_12009,N_7431,N_6921);
nand U12010 (N_12010,N_8546,N_8216);
nand U12011 (N_12011,N_7585,N_8934);
nor U12012 (N_12012,N_8055,N_6924);
nand U12013 (N_12013,N_6600,N_7314);
nand U12014 (N_12014,N_7623,N_6746);
and U12015 (N_12015,N_7429,N_6768);
xor U12016 (N_12016,N_8206,N_8620);
and U12017 (N_12017,N_7922,N_7613);
nor U12018 (N_12018,N_9041,N_8887);
and U12019 (N_12019,N_8641,N_6557);
nor U12020 (N_12020,N_7517,N_8920);
xor U12021 (N_12021,N_6257,N_7647);
or U12022 (N_12022,N_7480,N_7338);
xor U12023 (N_12023,N_6610,N_8677);
nor U12024 (N_12024,N_8645,N_8567);
nor U12025 (N_12025,N_8501,N_7486);
and U12026 (N_12026,N_9168,N_8721);
nor U12027 (N_12027,N_6913,N_7060);
or U12028 (N_12028,N_9125,N_8168);
xnor U12029 (N_12029,N_7248,N_8470);
nor U12030 (N_12030,N_7995,N_7362);
nor U12031 (N_12031,N_6979,N_6878);
or U12032 (N_12032,N_7526,N_7653);
and U12033 (N_12033,N_7898,N_8977);
or U12034 (N_12034,N_7963,N_7928);
or U12035 (N_12035,N_7258,N_6819);
or U12036 (N_12036,N_6451,N_6686);
or U12037 (N_12037,N_6402,N_8288);
nor U12038 (N_12038,N_7158,N_7553);
or U12039 (N_12039,N_9272,N_9257);
xor U12040 (N_12040,N_6547,N_8023);
xnor U12041 (N_12041,N_7010,N_9197);
or U12042 (N_12042,N_8886,N_6773);
nand U12043 (N_12043,N_8718,N_6888);
xor U12044 (N_12044,N_8630,N_6312);
or U12045 (N_12045,N_7249,N_6844);
nand U12046 (N_12046,N_6904,N_7387);
or U12047 (N_12047,N_8374,N_8850);
nor U12048 (N_12048,N_6655,N_7051);
and U12049 (N_12049,N_8667,N_9017);
xor U12050 (N_12050,N_8456,N_6954);
nor U12051 (N_12051,N_8571,N_7777);
or U12052 (N_12052,N_9227,N_7463);
nor U12053 (N_12053,N_6250,N_6803);
or U12054 (N_12054,N_6909,N_8470);
nor U12055 (N_12055,N_9157,N_9301);
and U12056 (N_12056,N_7062,N_7125);
or U12057 (N_12057,N_8825,N_6772);
and U12058 (N_12058,N_8398,N_8457);
or U12059 (N_12059,N_6411,N_6404);
xnor U12060 (N_12060,N_8580,N_8111);
or U12061 (N_12061,N_8168,N_6885);
or U12062 (N_12062,N_6723,N_6685);
or U12063 (N_12063,N_6483,N_6976);
and U12064 (N_12064,N_7316,N_8978);
nor U12065 (N_12065,N_7349,N_7852);
xor U12066 (N_12066,N_6658,N_8888);
or U12067 (N_12067,N_6792,N_8600);
xor U12068 (N_12068,N_8810,N_6327);
or U12069 (N_12069,N_7006,N_8926);
and U12070 (N_12070,N_7414,N_7991);
and U12071 (N_12071,N_6700,N_7586);
nand U12072 (N_12072,N_8684,N_7107);
or U12073 (N_12073,N_6765,N_7707);
and U12074 (N_12074,N_6773,N_7132);
nand U12075 (N_12075,N_8003,N_7754);
or U12076 (N_12076,N_7587,N_9029);
nor U12077 (N_12077,N_6540,N_9078);
nand U12078 (N_12078,N_6726,N_7835);
and U12079 (N_12079,N_7174,N_7872);
and U12080 (N_12080,N_6573,N_6992);
or U12081 (N_12081,N_7849,N_6306);
or U12082 (N_12082,N_7684,N_9094);
nor U12083 (N_12083,N_8658,N_7902);
nor U12084 (N_12084,N_7701,N_6993);
and U12085 (N_12085,N_6913,N_7509);
nand U12086 (N_12086,N_7520,N_7680);
and U12087 (N_12087,N_6995,N_6389);
xnor U12088 (N_12088,N_7203,N_8827);
nand U12089 (N_12089,N_7749,N_8668);
or U12090 (N_12090,N_7888,N_6681);
and U12091 (N_12091,N_7391,N_6977);
nand U12092 (N_12092,N_6272,N_8822);
nand U12093 (N_12093,N_7310,N_6822);
nor U12094 (N_12094,N_7713,N_7697);
or U12095 (N_12095,N_7955,N_8114);
and U12096 (N_12096,N_8728,N_8575);
nor U12097 (N_12097,N_8964,N_7873);
or U12098 (N_12098,N_6290,N_7597);
nor U12099 (N_12099,N_6550,N_7008);
nor U12100 (N_12100,N_6862,N_8131);
or U12101 (N_12101,N_8827,N_8479);
or U12102 (N_12102,N_9233,N_8344);
xor U12103 (N_12103,N_7731,N_6442);
and U12104 (N_12104,N_8827,N_8538);
and U12105 (N_12105,N_9044,N_7138);
or U12106 (N_12106,N_7048,N_7128);
nor U12107 (N_12107,N_7918,N_6938);
and U12108 (N_12108,N_6631,N_7523);
xor U12109 (N_12109,N_8630,N_7208);
nand U12110 (N_12110,N_8059,N_7759);
nand U12111 (N_12111,N_9250,N_8307);
and U12112 (N_12112,N_7981,N_8583);
nand U12113 (N_12113,N_8532,N_8351);
or U12114 (N_12114,N_8894,N_9346);
nand U12115 (N_12115,N_6362,N_7178);
nor U12116 (N_12116,N_7390,N_8558);
and U12117 (N_12117,N_7828,N_7065);
nand U12118 (N_12118,N_6918,N_7178);
nand U12119 (N_12119,N_7991,N_8468);
nor U12120 (N_12120,N_6811,N_6267);
xor U12121 (N_12121,N_9340,N_6683);
xor U12122 (N_12122,N_7529,N_6312);
or U12123 (N_12123,N_9211,N_7162);
nor U12124 (N_12124,N_7191,N_6531);
or U12125 (N_12125,N_8164,N_8012);
nand U12126 (N_12126,N_7155,N_9143);
or U12127 (N_12127,N_6986,N_8689);
xnor U12128 (N_12128,N_6262,N_8535);
xor U12129 (N_12129,N_6967,N_7773);
and U12130 (N_12130,N_6934,N_8846);
or U12131 (N_12131,N_7822,N_6371);
xnor U12132 (N_12132,N_8065,N_6678);
or U12133 (N_12133,N_9366,N_6435);
xor U12134 (N_12134,N_8564,N_6261);
nand U12135 (N_12135,N_7969,N_8104);
xnor U12136 (N_12136,N_6621,N_7928);
nand U12137 (N_12137,N_8588,N_8207);
or U12138 (N_12138,N_6486,N_8394);
and U12139 (N_12139,N_6433,N_9103);
xnor U12140 (N_12140,N_9227,N_7918);
nor U12141 (N_12141,N_7601,N_7929);
and U12142 (N_12142,N_7993,N_6823);
nor U12143 (N_12143,N_6261,N_8539);
or U12144 (N_12144,N_9101,N_8001);
and U12145 (N_12145,N_8985,N_8593);
nor U12146 (N_12146,N_6278,N_7127);
xor U12147 (N_12147,N_7943,N_9292);
or U12148 (N_12148,N_8448,N_8208);
nand U12149 (N_12149,N_6679,N_7584);
nor U12150 (N_12150,N_7069,N_7113);
xor U12151 (N_12151,N_8620,N_6940);
nand U12152 (N_12152,N_8874,N_8489);
nand U12153 (N_12153,N_6333,N_6652);
or U12154 (N_12154,N_6314,N_6325);
nor U12155 (N_12155,N_6623,N_6691);
or U12156 (N_12156,N_8679,N_7570);
and U12157 (N_12157,N_8043,N_8449);
nor U12158 (N_12158,N_6560,N_7800);
and U12159 (N_12159,N_7659,N_8115);
nor U12160 (N_12160,N_7086,N_7794);
xor U12161 (N_12161,N_8437,N_9181);
nand U12162 (N_12162,N_8231,N_7421);
nand U12163 (N_12163,N_6904,N_7124);
or U12164 (N_12164,N_6495,N_6705);
nand U12165 (N_12165,N_8347,N_6307);
and U12166 (N_12166,N_7622,N_9021);
nand U12167 (N_12167,N_9078,N_6662);
and U12168 (N_12168,N_6493,N_6706);
or U12169 (N_12169,N_8425,N_7292);
nor U12170 (N_12170,N_6594,N_8145);
nor U12171 (N_12171,N_7473,N_8601);
nor U12172 (N_12172,N_6811,N_8033);
or U12173 (N_12173,N_6317,N_6759);
or U12174 (N_12174,N_8335,N_9352);
or U12175 (N_12175,N_8841,N_6855);
nor U12176 (N_12176,N_6981,N_8193);
nor U12177 (N_12177,N_8457,N_9034);
and U12178 (N_12178,N_9003,N_8503);
or U12179 (N_12179,N_6545,N_8395);
nor U12180 (N_12180,N_9356,N_7018);
nand U12181 (N_12181,N_8784,N_8588);
nand U12182 (N_12182,N_9026,N_6959);
or U12183 (N_12183,N_7547,N_6600);
or U12184 (N_12184,N_7398,N_8573);
nor U12185 (N_12185,N_6516,N_7473);
nand U12186 (N_12186,N_7920,N_8411);
nor U12187 (N_12187,N_7784,N_7359);
nor U12188 (N_12188,N_7274,N_8483);
and U12189 (N_12189,N_9124,N_8217);
and U12190 (N_12190,N_6287,N_6495);
or U12191 (N_12191,N_8354,N_7009);
xor U12192 (N_12192,N_7724,N_7534);
nor U12193 (N_12193,N_6412,N_6535);
nand U12194 (N_12194,N_6805,N_6411);
and U12195 (N_12195,N_8465,N_8336);
nand U12196 (N_12196,N_6660,N_7749);
or U12197 (N_12197,N_7106,N_6898);
nor U12198 (N_12198,N_8062,N_6882);
nand U12199 (N_12199,N_8356,N_7542);
and U12200 (N_12200,N_8889,N_6296);
or U12201 (N_12201,N_7279,N_8546);
or U12202 (N_12202,N_6851,N_6826);
nor U12203 (N_12203,N_6778,N_9343);
nor U12204 (N_12204,N_7686,N_6687);
or U12205 (N_12205,N_8305,N_8356);
and U12206 (N_12206,N_9047,N_7784);
or U12207 (N_12207,N_6420,N_6659);
or U12208 (N_12208,N_6599,N_8667);
or U12209 (N_12209,N_8533,N_7463);
and U12210 (N_12210,N_7523,N_6302);
or U12211 (N_12211,N_8494,N_8157);
and U12212 (N_12212,N_9011,N_7653);
and U12213 (N_12213,N_8751,N_8922);
or U12214 (N_12214,N_6501,N_7028);
and U12215 (N_12215,N_8773,N_6557);
nand U12216 (N_12216,N_9136,N_7800);
nand U12217 (N_12217,N_7146,N_8863);
nand U12218 (N_12218,N_6503,N_8740);
nor U12219 (N_12219,N_7600,N_7041);
nand U12220 (N_12220,N_7821,N_6879);
or U12221 (N_12221,N_7842,N_8993);
or U12222 (N_12222,N_8202,N_6780);
nand U12223 (N_12223,N_7965,N_8966);
and U12224 (N_12224,N_8467,N_6909);
xnor U12225 (N_12225,N_9270,N_9138);
nor U12226 (N_12226,N_7044,N_7691);
xnor U12227 (N_12227,N_7276,N_8983);
nor U12228 (N_12228,N_9206,N_8516);
nand U12229 (N_12229,N_6503,N_6391);
nand U12230 (N_12230,N_7184,N_6789);
nand U12231 (N_12231,N_6773,N_8493);
or U12232 (N_12232,N_6545,N_8310);
nand U12233 (N_12233,N_8900,N_9129);
nand U12234 (N_12234,N_6983,N_9329);
nand U12235 (N_12235,N_8761,N_6498);
nor U12236 (N_12236,N_8354,N_6518);
or U12237 (N_12237,N_7174,N_9183);
nor U12238 (N_12238,N_6250,N_6373);
nor U12239 (N_12239,N_8783,N_7036);
nand U12240 (N_12240,N_6900,N_8517);
or U12241 (N_12241,N_7701,N_6356);
nand U12242 (N_12242,N_9125,N_7636);
and U12243 (N_12243,N_6697,N_8296);
nor U12244 (N_12244,N_8120,N_6623);
xnor U12245 (N_12245,N_8410,N_6342);
or U12246 (N_12246,N_7889,N_7390);
and U12247 (N_12247,N_9286,N_6508);
or U12248 (N_12248,N_8308,N_8907);
and U12249 (N_12249,N_7525,N_6378);
nand U12250 (N_12250,N_7751,N_8527);
nand U12251 (N_12251,N_7137,N_8524);
nand U12252 (N_12252,N_8463,N_6661);
xor U12253 (N_12253,N_7421,N_8942);
nor U12254 (N_12254,N_7041,N_6667);
and U12255 (N_12255,N_7182,N_8432);
nand U12256 (N_12256,N_8711,N_6485);
nand U12257 (N_12257,N_7635,N_8886);
and U12258 (N_12258,N_6471,N_7462);
and U12259 (N_12259,N_8260,N_7550);
nand U12260 (N_12260,N_8408,N_6929);
nor U12261 (N_12261,N_6708,N_9172);
or U12262 (N_12262,N_9066,N_6450);
nor U12263 (N_12263,N_7576,N_6941);
or U12264 (N_12264,N_8139,N_7451);
nor U12265 (N_12265,N_7445,N_7482);
xor U12266 (N_12266,N_8847,N_7313);
nand U12267 (N_12267,N_9145,N_7538);
nand U12268 (N_12268,N_6472,N_7878);
nand U12269 (N_12269,N_7899,N_6357);
nor U12270 (N_12270,N_8433,N_9287);
and U12271 (N_12271,N_6925,N_6533);
or U12272 (N_12272,N_8761,N_8777);
xor U12273 (N_12273,N_9060,N_6976);
nand U12274 (N_12274,N_7777,N_8946);
and U12275 (N_12275,N_8808,N_7908);
and U12276 (N_12276,N_8425,N_9362);
or U12277 (N_12277,N_8837,N_6705);
or U12278 (N_12278,N_8363,N_8256);
xor U12279 (N_12279,N_8004,N_7684);
nor U12280 (N_12280,N_7940,N_6773);
or U12281 (N_12281,N_7905,N_7355);
or U12282 (N_12282,N_8288,N_7394);
or U12283 (N_12283,N_7870,N_6507);
and U12284 (N_12284,N_8009,N_8528);
and U12285 (N_12285,N_7536,N_7504);
and U12286 (N_12286,N_7267,N_6340);
and U12287 (N_12287,N_7972,N_7129);
or U12288 (N_12288,N_8702,N_8336);
and U12289 (N_12289,N_6831,N_7690);
nor U12290 (N_12290,N_6335,N_7155);
or U12291 (N_12291,N_6798,N_8255);
nand U12292 (N_12292,N_6478,N_7863);
or U12293 (N_12293,N_9310,N_8579);
nand U12294 (N_12294,N_7265,N_8220);
nand U12295 (N_12295,N_8821,N_8198);
nor U12296 (N_12296,N_8706,N_6904);
nor U12297 (N_12297,N_7524,N_7446);
nor U12298 (N_12298,N_6296,N_8038);
or U12299 (N_12299,N_8151,N_8689);
nor U12300 (N_12300,N_7992,N_6679);
nor U12301 (N_12301,N_8701,N_6959);
nand U12302 (N_12302,N_7987,N_8460);
xnor U12303 (N_12303,N_8198,N_6800);
and U12304 (N_12304,N_7675,N_8613);
nand U12305 (N_12305,N_6494,N_8813);
nor U12306 (N_12306,N_9370,N_7396);
nor U12307 (N_12307,N_7890,N_6456);
nand U12308 (N_12308,N_6761,N_6901);
nand U12309 (N_12309,N_8177,N_7451);
nor U12310 (N_12310,N_8614,N_8855);
nor U12311 (N_12311,N_8813,N_8709);
nand U12312 (N_12312,N_9263,N_6924);
nor U12313 (N_12313,N_6777,N_8913);
or U12314 (N_12314,N_6865,N_7936);
nor U12315 (N_12315,N_7684,N_8650);
nor U12316 (N_12316,N_8778,N_7520);
nand U12317 (N_12317,N_8335,N_6287);
nor U12318 (N_12318,N_9337,N_8944);
and U12319 (N_12319,N_7928,N_9150);
or U12320 (N_12320,N_7743,N_9201);
nor U12321 (N_12321,N_8440,N_7793);
and U12322 (N_12322,N_7402,N_8594);
and U12323 (N_12323,N_8074,N_9354);
nand U12324 (N_12324,N_8331,N_9144);
or U12325 (N_12325,N_6357,N_7005);
and U12326 (N_12326,N_6424,N_7113);
nor U12327 (N_12327,N_7513,N_6538);
nor U12328 (N_12328,N_8332,N_7392);
nand U12329 (N_12329,N_8849,N_8264);
nand U12330 (N_12330,N_9362,N_6766);
and U12331 (N_12331,N_7099,N_9203);
or U12332 (N_12332,N_6693,N_8478);
xor U12333 (N_12333,N_7790,N_7065);
xnor U12334 (N_12334,N_8578,N_8477);
nand U12335 (N_12335,N_8033,N_7688);
nor U12336 (N_12336,N_7294,N_6868);
or U12337 (N_12337,N_7981,N_7111);
or U12338 (N_12338,N_6764,N_7186);
and U12339 (N_12339,N_7480,N_9078);
or U12340 (N_12340,N_8181,N_9197);
or U12341 (N_12341,N_7023,N_7779);
nor U12342 (N_12342,N_9178,N_8453);
and U12343 (N_12343,N_6778,N_9025);
nand U12344 (N_12344,N_8719,N_7904);
or U12345 (N_12345,N_8479,N_7837);
nor U12346 (N_12346,N_8804,N_7280);
nor U12347 (N_12347,N_7427,N_6547);
nor U12348 (N_12348,N_8874,N_9220);
nor U12349 (N_12349,N_6925,N_8725);
nor U12350 (N_12350,N_9086,N_9220);
nand U12351 (N_12351,N_7108,N_6703);
or U12352 (N_12352,N_9357,N_6965);
nand U12353 (N_12353,N_6927,N_7785);
and U12354 (N_12354,N_9310,N_8611);
nor U12355 (N_12355,N_8349,N_8562);
nand U12356 (N_12356,N_6524,N_7855);
nor U12357 (N_12357,N_8485,N_7417);
and U12358 (N_12358,N_8234,N_8350);
nand U12359 (N_12359,N_7517,N_7632);
and U12360 (N_12360,N_8246,N_7560);
nor U12361 (N_12361,N_6518,N_7329);
xnor U12362 (N_12362,N_8637,N_7909);
nor U12363 (N_12363,N_8438,N_8829);
nor U12364 (N_12364,N_8550,N_6613);
and U12365 (N_12365,N_7540,N_6923);
and U12366 (N_12366,N_8593,N_8062);
or U12367 (N_12367,N_8038,N_7772);
nand U12368 (N_12368,N_7896,N_7624);
xor U12369 (N_12369,N_9365,N_6677);
nor U12370 (N_12370,N_8168,N_8813);
nor U12371 (N_12371,N_8277,N_6885);
or U12372 (N_12372,N_7479,N_8993);
nand U12373 (N_12373,N_7480,N_8027);
nand U12374 (N_12374,N_7454,N_6864);
or U12375 (N_12375,N_8397,N_7169);
and U12376 (N_12376,N_7694,N_6692);
nand U12377 (N_12377,N_6799,N_8525);
or U12378 (N_12378,N_8040,N_8087);
and U12379 (N_12379,N_7536,N_8129);
nand U12380 (N_12380,N_7689,N_8443);
xnor U12381 (N_12381,N_7399,N_9029);
xnor U12382 (N_12382,N_7241,N_8575);
nor U12383 (N_12383,N_7166,N_9365);
and U12384 (N_12384,N_9192,N_8725);
and U12385 (N_12385,N_8021,N_8291);
nor U12386 (N_12386,N_7163,N_8802);
nand U12387 (N_12387,N_7471,N_7559);
xnor U12388 (N_12388,N_8374,N_8352);
or U12389 (N_12389,N_8058,N_8111);
nand U12390 (N_12390,N_8342,N_8827);
nor U12391 (N_12391,N_8318,N_6928);
or U12392 (N_12392,N_7784,N_7106);
nor U12393 (N_12393,N_7990,N_7613);
nor U12394 (N_12394,N_8447,N_8488);
nand U12395 (N_12395,N_6832,N_7019);
or U12396 (N_12396,N_7828,N_6557);
or U12397 (N_12397,N_6385,N_7950);
or U12398 (N_12398,N_6364,N_7705);
nor U12399 (N_12399,N_7695,N_7974);
or U12400 (N_12400,N_8654,N_9113);
nor U12401 (N_12401,N_7446,N_7593);
nand U12402 (N_12402,N_6710,N_6650);
nor U12403 (N_12403,N_7483,N_8224);
nor U12404 (N_12404,N_7409,N_6287);
xor U12405 (N_12405,N_9292,N_6733);
and U12406 (N_12406,N_6683,N_7928);
nor U12407 (N_12407,N_6855,N_8985);
or U12408 (N_12408,N_7333,N_8312);
and U12409 (N_12409,N_6268,N_9085);
nand U12410 (N_12410,N_7015,N_7029);
nor U12411 (N_12411,N_6787,N_7462);
nor U12412 (N_12412,N_6469,N_8289);
and U12413 (N_12413,N_6872,N_8050);
nand U12414 (N_12414,N_6739,N_7246);
and U12415 (N_12415,N_7701,N_9087);
or U12416 (N_12416,N_8998,N_7202);
nor U12417 (N_12417,N_9370,N_9099);
nand U12418 (N_12418,N_6253,N_9194);
xor U12419 (N_12419,N_6464,N_7406);
nor U12420 (N_12420,N_7127,N_7710);
nand U12421 (N_12421,N_7394,N_7003);
xnor U12422 (N_12422,N_6916,N_8963);
nand U12423 (N_12423,N_8931,N_9171);
nor U12424 (N_12424,N_9321,N_6981);
nand U12425 (N_12425,N_7915,N_7424);
and U12426 (N_12426,N_7268,N_6822);
nand U12427 (N_12427,N_7574,N_8968);
xnor U12428 (N_12428,N_7974,N_6328);
nand U12429 (N_12429,N_6942,N_9228);
nor U12430 (N_12430,N_7140,N_7463);
nor U12431 (N_12431,N_7250,N_6495);
nand U12432 (N_12432,N_8191,N_8712);
nand U12433 (N_12433,N_7233,N_8540);
and U12434 (N_12434,N_6357,N_6808);
nand U12435 (N_12435,N_9017,N_9116);
and U12436 (N_12436,N_6322,N_7222);
or U12437 (N_12437,N_6955,N_8216);
and U12438 (N_12438,N_7176,N_9100);
or U12439 (N_12439,N_8469,N_7561);
or U12440 (N_12440,N_9352,N_6293);
or U12441 (N_12441,N_9089,N_8980);
nor U12442 (N_12442,N_8519,N_8270);
nor U12443 (N_12443,N_8226,N_8024);
or U12444 (N_12444,N_9285,N_8227);
xor U12445 (N_12445,N_8947,N_7339);
or U12446 (N_12446,N_7413,N_7114);
nand U12447 (N_12447,N_7540,N_8993);
nand U12448 (N_12448,N_8112,N_6499);
or U12449 (N_12449,N_7769,N_6933);
nor U12450 (N_12450,N_7369,N_6545);
nand U12451 (N_12451,N_8965,N_8003);
or U12452 (N_12452,N_7818,N_8301);
nand U12453 (N_12453,N_8066,N_7054);
or U12454 (N_12454,N_8700,N_6866);
nand U12455 (N_12455,N_6998,N_6288);
or U12456 (N_12456,N_9314,N_6706);
xor U12457 (N_12457,N_9091,N_6967);
nor U12458 (N_12458,N_6661,N_9129);
nor U12459 (N_12459,N_7582,N_8081);
or U12460 (N_12460,N_9345,N_6949);
xor U12461 (N_12461,N_6795,N_7829);
nor U12462 (N_12462,N_7835,N_7827);
nand U12463 (N_12463,N_6988,N_7029);
and U12464 (N_12464,N_8832,N_8018);
and U12465 (N_12465,N_6582,N_7272);
nand U12466 (N_12466,N_6486,N_7213);
nor U12467 (N_12467,N_8766,N_8623);
and U12468 (N_12468,N_8757,N_9372);
nor U12469 (N_12469,N_6742,N_8696);
and U12470 (N_12470,N_6678,N_7869);
nor U12471 (N_12471,N_6617,N_7988);
and U12472 (N_12472,N_8563,N_7089);
and U12473 (N_12473,N_6999,N_7987);
and U12474 (N_12474,N_6956,N_6398);
nand U12475 (N_12475,N_7139,N_9267);
nor U12476 (N_12476,N_8049,N_8754);
xnor U12477 (N_12477,N_8912,N_8155);
and U12478 (N_12478,N_9248,N_8759);
xor U12479 (N_12479,N_9136,N_8065);
and U12480 (N_12480,N_8076,N_8921);
nand U12481 (N_12481,N_6930,N_6817);
or U12482 (N_12482,N_7696,N_7610);
or U12483 (N_12483,N_7954,N_8140);
and U12484 (N_12484,N_8843,N_8751);
and U12485 (N_12485,N_6640,N_8215);
nand U12486 (N_12486,N_6939,N_8026);
nand U12487 (N_12487,N_7717,N_9349);
and U12488 (N_12488,N_8100,N_8145);
nand U12489 (N_12489,N_6307,N_8274);
or U12490 (N_12490,N_8532,N_9008);
and U12491 (N_12491,N_6676,N_8214);
xor U12492 (N_12492,N_8739,N_7070);
or U12493 (N_12493,N_8214,N_8919);
and U12494 (N_12494,N_6931,N_8063);
or U12495 (N_12495,N_6584,N_8105);
nand U12496 (N_12496,N_7836,N_6954);
xor U12497 (N_12497,N_6713,N_9338);
and U12498 (N_12498,N_8959,N_8099);
nor U12499 (N_12499,N_7554,N_9017);
xor U12500 (N_12500,N_10521,N_12095);
or U12501 (N_12501,N_11413,N_10574);
or U12502 (N_12502,N_10503,N_9432);
or U12503 (N_12503,N_9717,N_10101);
xor U12504 (N_12504,N_10341,N_11278);
nor U12505 (N_12505,N_11057,N_10776);
or U12506 (N_12506,N_10280,N_12047);
nand U12507 (N_12507,N_12169,N_10211);
nand U12508 (N_12508,N_10231,N_10508);
nor U12509 (N_12509,N_10668,N_10463);
xnor U12510 (N_12510,N_10781,N_12143);
or U12511 (N_12511,N_10836,N_11596);
nand U12512 (N_12512,N_11075,N_11222);
or U12513 (N_12513,N_9928,N_10262);
nor U12514 (N_12514,N_9534,N_10243);
nor U12515 (N_12515,N_12031,N_11181);
nand U12516 (N_12516,N_10009,N_12011);
nor U12517 (N_12517,N_10866,N_11091);
and U12518 (N_12518,N_11674,N_11831);
and U12519 (N_12519,N_10007,N_10838);
xnor U12520 (N_12520,N_11749,N_11484);
nand U12521 (N_12521,N_12294,N_11789);
nand U12522 (N_12522,N_12334,N_10891);
nand U12523 (N_12523,N_9981,N_11783);
nor U12524 (N_12524,N_9515,N_9995);
nand U12525 (N_12525,N_11073,N_11996);
xor U12526 (N_12526,N_12118,N_9689);
nand U12527 (N_12527,N_11244,N_10059);
xor U12528 (N_12528,N_10529,N_9488);
and U12529 (N_12529,N_10352,N_10098);
nand U12530 (N_12530,N_9606,N_9910);
xnor U12531 (N_12531,N_12416,N_10090);
nand U12532 (N_12532,N_11662,N_9621);
nand U12533 (N_12533,N_11800,N_10633);
and U12534 (N_12534,N_9588,N_12090);
and U12535 (N_12535,N_12459,N_11145);
xnor U12536 (N_12536,N_11387,N_10496);
and U12537 (N_12537,N_10702,N_9566);
nand U12538 (N_12538,N_9834,N_12193);
and U12539 (N_12539,N_9945,N_10543);
nor U12540 (N_12540,N_12432,N_10116);
nand U12541 (N_12541,N_10142,N_12002);
xnor U12542 (N_12542,N_9657,N_11345);
nor U12543 (N_12543,N_12166,N_9844);
and U12544 (N_12544,N_11464,N_12164);
or U12545 (N_12545,N_12151,N_9871);
and U12546 (N_12546,N_11129,N_12378);
nand U12547 (N_12547,N_11926,N_10322);
nand U12548 (N_12548,N_11884,N_10774);
nor U12549 (N_12549,N_11577,N_10136);
or U12550 (N_12550,N_12295,N_10381);
or U12551 (N_12551,N_10736,N_12240);
nor U12552 (N_12552,N_10636,N_9411);
nand U12553 (N_12553,N_11356,N_11742);
nand U12554 (N_12554,N_11786,N_11245);
and U12555 (N_12555,N_11794,N_12330);
or U12556 (N_12556,N_11530,N_10843);
nor U12557 (N_12557,N_9791,N_9642);
or U12558 (N_12558,N_11207,N_10871);
nor U12559 (N_12559,N_11955,N_10617);
or U12560 (N_12560,N_11127,N_9510);
and U12561 (N_12561,N_9692,N_10137);
and U12562 (N_12562,N_12313,N_10154);
nand U12563 (N_12563,N_10346,N_10439);
or U12564 (N_12564,N_11943,N_10414);
and U12565 (N_12565,N_12176,N_10740);
nand U12566 (N_12566,N_12403,N_10222);
xnor U12567 (N_12567,N_10292,N_10974);
xnor U12568 (N_12568,N_11133,N_12381);
xor U12569 (N_12569,N_10445,N_11552);
or U12570 (N_12570,N_10742,N_9448);
nand U12571 (N_12571,N_9568,N_12274);
xor U12572 (N_12572,N_11855,N_9915);
nor U12573 (N_12573,N_9982,N_9536);
and U12574 (N_12574,N_9636,N_11970);
nand U12575 (N_12575,N_10519,N_11515);
and U12576 (N_12576,N_9589,N_9545);
and U12577 (N_12577,N_11904,N_11443);
nor U12578 (N_12578,N_11374,N_12208);
or U12579 (N_12579,N_11286,N_9538);
nor U12580 (N_12580,N_11583,N_10818);
and U12581 (N_12581,N_11179,N_10797);
nand U12582 (N_12582,N_10255,N_11879);
and U12583 (N_12583,N_11924,N_11575);
and U12584 (N_12584,N_9394,N_9985);
nand U12585 (N_12585,N_12326,N_10491);
nand U12586 (N_12586,N_10535,N_11960);
or U12587 (N_12587,N_10450,N_11015);
nand U12588 (N_12588,N_11251,N_9397);
nor U12589 (N_12589,N_10965,N_11003);
nor U12590 (N_12590,N_11485,N_9919);
and U12591 (N_12591,N_11098,N_11185);
nor U12592 (N_12592,N_10763,N_9724);
or U12593 (N_12593,N_11937,N_10934);
and U12594 (N_12594,N_11110,N_9508);
and U12595 (N_12595,N_10865,N_9385);
nand U12596 (N_12596,N_10470,N_9709);
nand U12597 (N_12597,N_10822,N_11337);
or U12598 (N_12598,N_11574,N_10462);
nor U12599 (N_12599,N_10902,N_10619);
or U12600 (N_12600,N_10277,N_10706);
xor U12601 (N_12601,N_12037,N_12149);
nand U12602 (N_12602,N_12483,N_11467);
nand U12603 (N_12603,N_10783,N_11958);
xor U12604 (N_12604,N_10062,N_9728);
nand U12605 (N_12605,N_10817,N_11608);
nor U12606 (N_12606,N_10998,N_9810);
and U12607 (N_12607,N_9962,N_11232);
and U12608 (N_12608,N_11516,N_9492);
nor U12609 (N_12609,N_12191,N_11846);
and U12610 (N_12610,N_10741,N_11045);
nor U12611 (N_12611,N_11798,N_11657);
or U12612 (N_12612,N_10594,N_11947);
or U12613 (N_12613,N_12084,N_9529);
nand U12614 (N_12614,N_11827,N_10875);
or U12615 (N_12615,N_10613,N_12360);
nand U12616 (N_12616,N_10881,N_12324);
and U12617 (N_12617,N_9444,N_10933);
nand U12618 (N_12618,N_11494,N_10383);
nor U12619 (N_12619,N_10591,N_11806);
or U12620 (N_12620,N_11039,N_9680);
or U12621 (N_12621,N_11532,N_11055);
xnor U12622 (N_12622,N_10129,N_10584);
nand U12623 (N_12623,N_12484,N_11762);
nand U12624 (N_12624,N_9610,N_11673);
or U12625 (N_12625,N_11505,N_9922);
or U12626 (N_12626,N_10505,N_10523);
nor U12627 (N_12627,N_11314,N_11188);
nand U12628 (N_12628,N_11908,N_11991);
or U12629 (N_12629,N_11597,N_12343);
nor U12630 (N_12630,N_12203,N_12442);
or U12631 (N_12631,N_11711,N_11435);
xor U12632 (N_12632,N_9654,N_9384);
nor U12633 (N_12633,N_9990,N_9739);
or U12634 (N_12634,N_11343,N_11809);
and U12635 (N_12635,N_11441,N_11071);
nand U12636 (N_12636,N_12048,N_11650);
xnor U12637 (N_12637,N_10378,N_11829);
nand U12638 (N_12638,N_10180,N_10769);
xnor U12639 (N_12639,N_11945,N_11585);
or U12640 (N_12640,N_11121,N_11070);
and U12641 (N_12641,N_9929,N_10525);
xnor U12642 (N_12642,N_10812,N_12417);
nand U12643 (N_12643,N_10405,N_10995);
and U12644 (N_12644,N_11770,N_9651);
and U12645 (N_12645,N_10653,N_10206);
nor U12646 (N_12646,N_12289,N_11698);
nand U12647 (N_12647,N_11874,N_10249);
and U12648 (N_12648,N_11496,N_9874);
and U12649 (N_12649,N_9800,N_9644);
xor U12650 (N_12650,N_9404,N_10198);
nor U12651 (N_12651,N_12024,N_10607);
xor U12652 (N_12652,N_11400,N_12435);
or U12653 (N_12653,N_12448,N_10606);
or U12654 (N_12654,N_9480,N_11308);
nand U12655 (N_12655,N_11976,N_10885);
xnor U12656 (N_12656,N_11099,N_10828);
nand U12657 (N_12657,N_10560,N_9379);
nand U12658 (N_12658,N_11734,N_10155);
nor U12659 (N_12659,N_9387,N_10131);
xor U12660 (N_12660,N_10916,N_11940);
nor U12661 (N_12661,N_11439,N_9831);
xor U12662 (N_12662,N_10721,N_11566);
or U12663 (N_12663,N_10087,N_10404);
nand U12664 (N_12664,N_12056,N_10366);
nand U12665 (N_12665,N_11640,N_9599);
or U12666 (N_12666,N_12086,N_11281);
and U12667 (N_12667,N_10889,N_12280);
and U12668 (N_12668,N_10284,N_11270);
nor U12669 (N_12669,N_11171,N_11257);
and U12670 (N_12670,N_11229,N_12285);
or U12671 (N_12671,N_12434,N_10122);
or U12672 (N_12672,N_11214,N_10376);
nor U12673 (N_12673,N_9653,N_11396);
nor U12674 (N_12674,N_9400,N_11667);
xor U12675 (N_12675,N_11609,N_12113);
xor U12676 (N_12676,N_10458,N_9950);
and U12677 (N_12677,N_10796,N_10827);
nor U12678 (N_12678,N_10270,N_11157);
or U12679 (N_12679,N_9701,N_10273);
or U12680 (N_12680,N_10230,N_12019);
nor U12681 (N_12681,N_12287,N_11094);
nand U12682 (N_12682,N_11864,N_10791);
nor U12683 (N_12683,N_9509,N_11304);
nand U12684 (N_12684,N_12478,N_11436);
or U12685 (N_12685,N_10984,N_11856);
or U12686 (N_12686,N_9861,N_11573);
nand U12687 (N_12687,N_11042,N_9803);
and U12688 (N_12688,N_12254,N_10297);
or U12689 (N_12689,N_10616,N_11095);
or U12690 (N_12690,N_10219,N_10927);
or U12691 (N_12691,N_12440,N_10710);
and U12692 (N_12692,N_9482,N_9417);
nor U12693 (N_12693,N_9939,N_10005);
or U12694 (N_12694,N_10854,N_11663);
or U12695 (N_12695,N_9494,N_10054);
and U12696 (N_12696,N_11598,N_11366);
nor U12697 (N_12697,N_11194,N_10534);
or U12698 (N_12698,N_10247,N_12265);
xnor U12699 (N_12699,N_9434,N_11456);
nor U12700 (N_12700,N_10704,N_10072);
and U12701 (N_12701,N_11953,N_12135);
nand U12702 (N_12702,N_10430,N_11344);
and U12703 (N_12703,N_9814,N_10312);
or U12704 (N_12704,N_10127,N_11062);
nand U12705 (N_12705,N_10794,N_12430);
nor U12706 (N_12706,N_11932,N_11838);
and U12707 (N_12707,N_10202,N_10391);
and U12708 (N_12708,N_10406,N_10819);
and U12709 (N_12709,N_12137,N_10821);
and U12710 (N_12710,N_11192,N_9487);
or U12711 (N_12711,N_10799,N_10133);
nor U12712 (N_12712,N_11202,N_10217);
xor U12713 (N_12713,N_10055,N_11152);
nor U12714 (N_12714,N_11753,N_12490);
nor U12715 (N_12715,N_10354,N_9877);
nand U12716 (N_12716,N_9464,N_10325);
nand U12717 (N_12717,N_9907,N_10851);
nor U12718 (N_12718,N_10622,N_12229);
nand U12719 (N_12719,N_11537,N_12352);
nor U12720 (N_12720,N_10815,N_10402);
nand U12721 (N_12721,N_12312,N_10757);
and U12722 (N_12722,N_10333,N_11390);
and U12723 (N_12723,N_11318,N_10627);
or U12724 (N_12724,N_9825,N_10755);
xnor U12725 (N_12725,N_12277,N_11853);
and U12726 (N_12726,N_12241,N_11253);
nand U12727 (N_12727,N_11499,N_11148);
or U12728 (N_12728,N_9836,N_10811);
nor U12729 (N_12729,N_10259,N_9423);
and U12730 (N_12730,N_9638,N_10999);
and U12731 (N_12731,N_11747,N_11064);
nor U12732 (N_12732,N_10468,N_11466);
or U12733 (N_12733,N_10724,N_11733);
or U12734 (N_12734,N_11922,N_10629);
or U12735 (N_12735,N_10375,N_10513);
or U12736 (N_12736,N_9587,N_10729);
nand U12737 (N_12737,N_12069,N_9770);
and U12738 (N_12738,N_11891,N_11936);
nand U12739 (N_12739,N_11067,N_9410);
nor U12740 (N_12740,N_10960,N_11618);
nand U12741 (N_12741,N_10362,N_11842);
and U12742 (N_12742,N_9443,N_10532);
nand U12743 (N_12743,N_12181,N_11751);
nor U12744 (N_12744,N_11123,N_10530);
or U12745 (N_12745,N_11471,N_11427);
and U12746 (N_12746,N_11331,N_10514);
nand U12747 (N_12747,N_10688,N_10074);
nand U12748 (N_12748,N_9398,N_9532);
xor U12749 (N_12749,N_10477,N_11419);
or U12750 (N_12750,N_10476,N_11600);
and U12751 (N_12751,N_9513,N_11483);
and U12752 (N_12752,N_10052,N_10480);
or U12753 (N_12753,N_11927,N_11364);
nor U12754 (N_12754,N_12192,N_12060);
or U12755 (N_12755,N_12445,N_9595);
nand U12756 (N_12756,N_11275,N_10146);
and U12757 (N_12757,N_10245,N_11124);
nand U12758 (N_12758,N_10749,N_9745);
and U12759 (N_12759,N_12453,N_11754);
xor U12760 (N_12760,N_10303,N_10428);
xor U12761 (N_12761,N_9673,N_10631);
nor U12762 (N_12762,N_12014,N_11659);
and U12763 (N_12763,N_11323,N_12489);
xor U12764 (N_12764,N_9921,N_10380);
and U12765 (N_12765,N_9900,N_12177);
or U12766 (N_12766,N_9511,N_12346);
nor U12767 (N_12767,N_12171,N_10486);
and U12768 (N_12768,N_11558,N_12423);
xnor U12769 (N_12769,N_10319,N_10045);
and U12770 (N_12770,N_11590,N_11728);
xnor U12771 (N_12771,N_12027,N_10436);
nor U12772 (N_12772,N_9421,N_10909);
or U12773 (N_12773,N_10438,N_10913);
and U12774 (N_12774,N_10646,N_9547);
nand U12775 (N_12775,N_11085,N_12038);
nor U12776 (N_12776,N_12206,N_10343);
nor U12777 (N_12777,N_11902,N_10762);
xor U12778 (N_12778,N_10650,N_10566);
nor U12779 (N_12779,N_12260,N_10203);
or U12780 (N_12780,N_9548,N_11671);
xnor U12781 (N_12781,N_9389,N_10461);
nand U12782 (N_12782,N_9934,N_12405);
and U12783 (N_12783,N_9892,N_11226);
and U12784 (N_12784,N_10412,N_11658);
nor U12785 (N_12785,N_9878,N_12252);
nor U12786 (N_12786,N_10670,N_12369);
nor U12787 (N_12787,N_11163,N_10106);
nand U12788 (N_12788,N_12292,N_9808);
xor U12789 (N_12789,N_9375,N_9468);
and U12790 (N_12790,N_11812,N_12178);
xnor U12791 (N_12791,N_10326,N_9522);
and U12792 (N_12792,N_10469,N_11969);
xnor U12793 (N_12793,N_10077,N_10041);
or U12794 (N_12794,N_12134,N_10210);
nor U12795 (N_12795,N_12467,N_10390);
or U12796 (N_12796,N_11724,N_11804);
and U12797 (N_12797,N_9584,N_10835);
nand U12798 (N_12798,N_9996,N_10232);
nand U12799 (N_12799,N_10457,N_11028);
nor U12800 (N_12800,N_9899,N_11986);
xor U12801 (N_12801,N_11524,N_10361);
nand U12802 (N_12802,N_10531,N_9983);
or U12803 (N_12803,N_10795,N_11486);
and U12804 (N_12804,N_9806,N_11649);
nand U12805 (N_12805,N_12070,N_9794);
nand U12806 (N_12806,N_10658,N_10638);
and U12807 (N_12807,N_10618,N_9430);
nand U12808 (N_12808,N_10113,N_9751);
nand U12809 (N_12809,N_10242,N_12253);
xnor U12810 (N_12810,N_9916,N_9700);
nand U12811 (N_12811,N_11956,N_11588);
or U12812 (N_12812,N_11153,N_9987);
nand U12813 (N_12813,N_11433,N_11048);
nor U12814 (N_12814,N_10179,N_11495);
or U12815 (N_12815,N_11639,N_11973);
xor U12816 (N_12816,N_12126,N_11569);
or U12817 (N_12817,N_11688,N_12264);
or U12818 (N_12818,N_10895,N_10167);
and U12819 (N_12819,N_12407,N_10568);
or U12820 (N_12820,N_12349,N_11230);
nor U12821 (N_12821,N_10268,N_10315);
nor U12822 (N_12822,N_11665,N_9574);
nand U12823 (N_12823,N_11206,N_10360);
or U12824 (N_12824,N_11533,N_10845);
or U12825 (N_12825,N_11677,N_12245);
nor U12826 (N_12826,N_9440,N_10034);
or U12827 (N_12827,N_9821,N_9586);
nand U12828 (N_12828,N_9577,N_12148);
or U12829 (N_12829,N_11913,N_12234);
nand U12830 (N_12830,N_9670,N_9669);
and U12831 (N_12831,N_10806,N_12196);
and U12832 (N_12832,N_9879,N_11707);
nor U12833 (N_12833,N_10788,N_10642);
or U12834 (N_12834,N_9813,N_12398);
and U12835 (N_12835,N_12428,N_9965);
and U12836 (N_12836,N_9516,N_9390);
nand U12837 (N_12837,N_12498,N_12447);
nand U12838 (N_12838,N_12000,N_11033);
and U12839 (N_12839,N_10920,N_9695);
or U12840 (N_12840,N_10656,N_10425);
nand U12841 (N_12841,N_9714,N_9776);
nor U12842 (N_12842,N_11116,N_9467);
and U12843 (N_12843,N_10223,N_11412);
nand U12844 (N_12844,N_10302,N_10479);
and U12845 (N_12845,N_11981,N_11572);
nand U12846 (N_12846,N_10904,N_12074);
nand U12847 (N_12847,N_10169,N_11001);
nand U12848 (N_12848,N_10666,N_10388);
nor U12849 (N_12849,N_11604,N_11336);
nand U12850 (N_12850,N_10427,N_12081);
xor U12851 (N_12851,N_9761,N_10765);
and U12852 (N_12852,N_11426,N_12341);
nand U12853 (N_12853,N_10094,N_11289);
and U12854 (N_12854,N_12053,N_10538);
and U12855 (N_12855,N_10204,N_10421);
or U12856 (N_12856,N_10478,N_10161);
or U12857 (N_12857,N_10536,N_9852);
or U12858 (N_12858,N_10107,N_10082);
or U12859 (N_12859,N_10108,N_12362);
nand U12860 (N_12860,N_11545,N_10397);
nand U12861 (N_12861,N_11478,N_11288);
nand U12862 (N_12862,N_10334,N_9832);
nand U12863 (N_12863,N_10429,N_9426);
nor U12864 (N_12864,N_11404,N_11643);
or U12865 (N_12865,N_10067,N_11235);
and U12866 (N_12866,N_10024,N_10586);
nor U12867 (N_12867,N_12248,N_11617);
nand U12868 (N_12868,N_10582,N_10580);
xor U12869 (N_12869,N_9613,N_10569);
nand U12870 (N_12870,N_12474,N_11024);
nor U12871 (N_12871,N_10978,N_9740);
nand U12872 (N_12872,N_11005,N_11738);
nor U12873 (N_12873,N_9629,N_9446);
nor U12874 (N_12874,N_9958,N_10956);
or U12875 (N_12875,N_10473,N_11167);
nor U12876 (N_12876,N_11361,N_10598);
nor U12877 (N_12877,N_11046,N_11714);
nand U12878 (N_12878,N_11267,N_9531);
or U12879 (N_12879,N_11077,N_11131);
nand U12880 (N_12880,N_9957,N_12340);
nand U12881 (N_12881,N_11210,N_11186);
xnor U12882 (N_12882,N_10079,N_11303);
xnor U12883 (N_12883,N_10193,N_10677);
and U12884 (N_12884,N_11195,N_11900);
or U12885 (N_12885,N_12415,N_12227);
nand U12886 (N_12886,N_10570,N_11497);
nand U12887 (N_12887,N_11538,N_11136);
and U12888 (N_12888,N_10331,N_12470);
or U12889 (N_12889,N_10509,N_10780);
or U12890 (N_12890,N_10524,N_10683);
nor U12891 (N_12891,N_10951,N_9582);
and U12892 (N_12892,N_9935,N_9865);
xor U12893 (N_12893,N_11859,N_10571);
nor U12894 (N_12894,N_9683,N_12057);
nand U12895 (N_12895,N_10985,N_9817);
and U12896 (N_12896,N_12373,N_11790);
nor U12897 (N_12897,N_11138,N_9771);
and U12898 (N_12898,N_10981,N_11920);
and U12899 (N_12899,N_11542,N_11858);
nor U12900 (N_12900,N_10493,N_11009);
xnor U12901 (N_12901,N_9798,N_12243);
nor U12902 (N_12902,N_11114,N_9635);
nor U12903 (N_12903,N_12111,N_10112);
nor U12904 (N_12904,N_10792,N_11686);
nand U12905 (N_12905,N_10873,N_12043);
xor U12906 (N_12906,N_9783,N_12273);
or U12907 (N_12907,N_11462,N_11236);
and U12908 (N_12908,N_9895,N_11642);
and U12909 (N_12909,N_9399,N_10252);
nor U12910 (N_12910,N_10977,N_11508);
nand U12911 (N_12911,N_9540,N_9475);
and U12912 (N_12912,N_10737,N_10025);
nand U12913 (N_12913,N_10086,N_11013);
and U12914 (N_12914,N_11240,N_10639);
or U12915 (N_12915,N_9864,N_11810);
or U12916 (N_12916,N_12465,N_12282);
or U12917 (N_12917,N_9941,N_9696);
or U12918 (N_12918,N_10685,N_12046);
nor U12919 (N_12919,N_9604,N_11000);
and U12920 (N_12920,N_11815,N_10208);
or U12921 (N_12921,N_11784,N_12195);
and U12922 (N_12922,N_10182,N_12106);
nor U12923 (N_12923,N_11388,N_11634);
xnor U12924 (N_12924,N_11011,N_9615);
and U12925 (N_12925,N_11615,N_12197);
or U12926 (N_12926,N_10578,N_9526);
nand U12927 (N_12927,N_9827,N_11372);
nor U12928 (N_12928,N_10558,N_10400);
nand U12929 (N_12929,N_11654,N_12117);
and U12930 (N_12930,N_9503,N_12286);
nor U12931 (N_12931,N_11736,N_10660);
and U12932 (N_12932,N_11078,N_12220);
and U12933 (N_12933,N_12141,N_11249);
nand U12934 (N_12934,N_10426,N_11780);
xnor U12935 (N_12935,N_12123,N_10874);
and U12936 (N_12936,N_10810,N_11498);
or U12937 (N_12937,N_11962,N_9799);
nor U12938 (N_12938,N_11813,N_9512);
xor U12939 (N_12939,N_9969,N_10859);
nor U12940 (N_12940,N_9826,N_9691);
nand U12941 (N_12941,N_10042,N_9698);
nand U12942 (N_12942,N_9749,N_10968);
nor U12943 (N_12943,N_10922,N_11835);
nor U12944 (N_12944,N_12353,N_10733);
and U12945 (N_12945,N_10684,N_11370);
nand U12946 (N_12946,N_11151,N_10964);
nand U12947 (N_12947,N_9859,N_10745);
and U12948 (N_12948,N_10474,N_12354);
or U12949 (N_12949,N_9449,N_9930);
nand U12950 (N_12950,N_12144,N_10860);
or U12951 (N_12951,N_10526,N_10359);
and U12952 (N_12952,N_10184,N_9590);
nor U12953 (N_12953,N_10840,N_9413);
xor U12954 (N_12954,N_11579,N_11354);
and U12955 (N_12955,N_11389,N_11144);
or U12956 (N_12956,N_10471,N_10910);
and U12957 (N_12957,N_10948,N_10545);
or U12958 (N_12958,N_11823,N_9556);
and U12959 (N_12959,N_11213,N_10778);
and U12960 (N_12960,N_12455,N_12044);
nand U12961 (N_12961,N_10295,N_11872);
and U12962 (N_12962,N_10422,N_11887);
nor U12963 (N_12963,N_9773,N_11787);
and U12964 (N_12964,N_11215,N_12039);
and U12965 (N_12965,N_11043,N_10833);
or U12966 (N_12966,N_9893,N_12393);
or U12967 (N_12967,N_12482,N_10730);
or U12968 (N_12968,N_9578,N_9786);
or U12969 (N_12969,N_11239,N_11285);
nand U12970 (N_12970,N_11854,N_11126);
and U12971 (N_12971,N_12036,N_10393);
or U12972 (N_12972,N_11160,N_10092);
nand U12973 (N_12973,N_12250,N_12267);
and U12974 (N_12974,N_11442,N_10703);
nand U12975 (N_12975,N_11555,N_9793);
nor U12976 (N_12976,N_12358,N_10205);
nand U12977 (N_12977,N_11030,N_9386);
nor U12978 (N_12978,N_10275,N_11863);
nand U12979 (N_12979,N_12433,N_11549);
or U12980 (N_12980,N_12009,N_12230);
nor U12981 (N_12981,N_10111,N_10507);
nor U12982 (N_12982,N_10357,N_11966);
or U12983 (N_12983,N_11700,N_11529);
nor U12984 (N_12984,N_11432,N_9658);
nor U12985 (N_12985,N_12006,N_10465);
nor U12986 (N_12986,N_12439,N_11660);
and U12987 (N_12987,N_11358,N_9764);
nand U12988 (N_12988,N_9465,N_11694);
and U12989 (N_12989,N_11886,N_12159);
nand U12990 (N_12990,N_9447,N_12235);
nand U12991 (N_12991,N_12412,N_11273);
nor U12992 (N_12992,N_12266,N_11164);
xor U12993 (N_12993,N_10775,N_11403);
or U12994 (N_12994,N_12497,N_10058);
and U12995 (N_12995,N_11595,N_10192);
or U12996 (N_12996,N_10732,N_10171);
nor U12997 (N_12997,N_11755,N_9675);
nor U12998 (N_12998,N_12216,N_10038);
and U12999 (N_12999,N_9901,N_11265);
or U13000 (N_13000,N_11933,N_12058);
nor U13001 (N_13001,N_11717,N_12087);
or U13002 (N_13002,N_11571,N_12213);
nand U13003 (N_13003,N_10162,N_9868);
xnor U13004 (N_13004,N_9829,N_11802);
nand U13005 (N_13005,N_9439,N_11061);
and U13006 (N_13006,N_11102,N_10299);
nand U13007 (N_13007,N_9942,N_9473);
and U13008 (N_13008,N_10014,N_11567);
and U13009 (N_13009,N_9501,N_10298);
or U13010 (N_13010,N_12138,N_12444);
nor U13011 (N_13011,N_10564,N_12310);
or U13012 (N_13012,N_11238,N_10287);
nor U13013 (N_13013,N_9662,N_11105);
or U13014 (N_13014,N_10417,N_9484);
nand U13015 (N_13015,N_9550,N_11150);
nor U13016 (N_13016,N_11295,N_11935);
nor U13017 (N_13017,N_11279,N_11923);
and U13018 (N_13018,N_11948,N_12309);
nor U13019 (N_13019,N_10248,N_11627);
xor U13020 (N_13020,N_10118,N_10318);
nand U13021 (N_13021,N_9940,N_11851);
and U13022 (N_13022,N_12156,N_9737);
and U13023 (N_13023,N_12172,N_11221);
nor U13024 (N_13024,N_10748,N_10746);
and U13025 (N_13025,N_10516,N_11080);
nand U13026 (N_13026,N_11931,N_11557);
and U13027 (N_13027,N_10713,N_10164);
or U13028 (N_13028,N_12293,N_9616);
xnor U13029 (N_13029,N_10869,N_11862);
or U13030 (N_13030,N_10047,N_10499);
nor U13031 (N_13031,N_10831,N_9592);
xnor U13032 (N_13032,N_9570,N_12231);
or U13033 (N_13033,N_12210,N_12030);
xnor U13034 (N_13034,N_11301,N_9766);
nor U13035 (N_13035,N_11348,N_10973);
xor U13036 (N_13036,N_11601,N_12025);
or U13037 (N_13037,N_11705,N_10698);
nor U13038 (N_13038,N_11488,N_10576);
nand U13039 (N_13039,N_9648,N_9558);
or U13040 (N_13040,N_11952,N_10296);
nand U13041 (N_13041,N_12104,N_10990);
nand U13042 (N_13042,N_10829,N_11701);
or U13043 (N_13043,N_12325,N_10446);
nor U13044 (N_13044,N_10549,N_9876);
or U13045 (N_13045,N_11656,N_11704);
nor U13046 (N_13046,N_11402,N_10693);
and U13047 (N_13047,N_12270,N_10502);
xor U13048 (N_13048,N_11578,N_11875);
nand U13049 (N_13049,N_9530,N_9477);
and U13050 (N_13050,N_9624,N_12278);
nor U13051 (N_13051,N_11218,N_12102);
nand U13052 (N_13052,N_11541,N_12413);
or U13053 (N_13053,N_12202,N_10886);
or U13054 (N_13054,N_11584,N_11570);
nand U13055 (N_13055,N_9597,N_9795);
and U13056 (N_13056,N_11633,N_9883);
or U13057 (N_13057,N_10777,N_9971);
or U13058 (N_13058,N_12249,N_11299);
xor U13059 (N_13059,N_10738,N_10379);
or U13060 (N_13060,N_11108,N_12476);
nor U13061 (N_13061,N_9485,N_11964);
nor U13062 (N_13062,N_11290,N_11768);
nor U13063 (N_13063,N_11504,N_10879);
and U13064 (N_13064,N_12276,N_11599);
nand U13065 (N_13065,N_11769,N_12154);
nor U13066 (N_13066,N_11603,N_10751);
nand U13067 (N_13067,N_10274,N_10173);
nor U13068 (N_13068,N_11322,N_9445);
nor U13069 (N_13069,N_9567,N_10676);
nand U13070 (N_13070,N_10120,N_10100);
or U13071 (N_13071,N_10085,N_10768);
and U13072 (N_13072,N_11233,N_10288);
nor U13073 (N_13073,N_10553,N_10039);
nand U13074 (N_13074,N_9811,N_12480);
and U13075 (N_13075,N_11446,N_9726);
nand U13076 (N_13076,N_10991,N_11326);
nor U13077 (N_13077,N_10595,N_11018);
or U13078 (N_13078,N_11506,N_10528);
nor U13079 (N_13079,N_11149,N_11219);
or U13080 (N_13080,N_9627,N_11510);
nand U13081 (N_13081,N_10784,N_9666);
xor U13082 (N_13082,N_11772,N_11526);
nor U13083 (N_13083,N_10475,N_11522);
nand U13084 (N_13084,N_12397,N_11255);
nand U13085 (N_13085,N_12438,N_10856);
nand U13086 (N_13086,N_11894,N_11231);
nor U13087 (N_13087,N_9779,N_9422);
nand U13088 (N_13088,N_11375,N_11680);
and U13089 (N_13089,N_11187,N_11957);
and U13090 (N_13090,N_9456,N_10012);
or U13091 (N_13091,N_11104,N_10648);
xnor U13092 (N_13092,N_11616,N_12165);
xor U13093 (N_13093,N_10722,N_10573);
xor U13094 (N_13094,N_10218,N_11357);
and U13095 (N_13095,N_11074,N_10579);
nand U13096 (N_13096,N_11263,N_12368);
or U13097 (N_13097,N_9461,N_11010);
xnor U13098 (N_13098,N_10601,N_10770);
nor U13099 (N_13099,N_10893,N_10483);
nor U13100 (N_13100,N_11328,N_11685);
and U13101 (N_13101,N_10339,N_11170);
nand U13102 (N_13102,N_11444,N_11689);
or U13103 (N_13103,N_10065,N_9917);
nand U13104 (N_13104,N_11582,N_10345);
or U13105 (N_13105,N_11999,N_12115);
nand U13106 (N_13106,N_11089,N_12017);
nand U13107 (N_13107,N_10997,N_11468);
and U13108 (N_13108,N_9999,N_11420);
and U13109 (N_13109,N_10482,N_10267);
nor U13110 (N_13110,N_10278,N_10971);
nand U13111 (N_13111,N_10608,N_10864);
or U13112 (N_13112,N_11565,N_11371);
nand U13113 (N_13113,N_9782,N_9500);
and U13114 (N_13114,N_10369,N_12174);
and U13115 (N_13115,N_11293,N_12001);
and U13116 (N_13116,N_10719,N_10515);
or U13117 (N_13117,N_12365,N_11325);
or U13118 (N_13118,N_9967,N_9565);
nor U13119 (N_13119,N_11740,N_12363);
and U13120 (N_13120,N_11415,N_11543);
nand U13121 (N_13121,N_12182,N_10929);
or U13122 (N_13122,N_12064,N_10980);
and U13123 (N_13123,N_11036,N_11901);
nand U13124 (N_13124,N_10221,N_11416);
and U13125 (N_13125,N_9517,N_12488);
or U13126 (N_13126,N_11681,N_11172);
xor U13127 (N_13127,N_10061,N_11423);
or U13128 (N_13128,N_11072,N_10599);
and U13129 (N_13129,N_10027,N_9732);
and U13130 (N_13130,N_11053,N_10563);
and U13131 (N_13131,N_12098,N_11209);
nor U13132 (N_13132,N_10460,N_11775);
nand U13133 (N_13133,N_11369,N_10903);
nand U13134 (N_13134,N_11702,N_11076);
and U13135 (N_13135,N_12211,N_12464);
nand U13136 (N_13136,N_12350,N_11756);
or U13137 (N_13137,N_10177,N_11173);
and U13138 (N_13138,N_9991,N_11882);
or U13139 (N_13139,N_10805,N_12461);
nand U13140 (N_13140,N_9679,N_11843);
or U13141 (N_13141,N_9593,N_11873);
or U13142 (N_13142,N_9993,N_12212);
xnor U13143 (N_13143,N_10605,N_11176);
and U13144 (N_13144,N_12355,N_11735);
or U13145 (N_13145,N_10395,N_9551);
and U13146 (N_13146,N_10604,N_11216);
nor U13147 (N_13147,N_9992,N_9601);
or U13148 (N_13148,N_9789,N_11117);
or U13149 (N_13149,N_12020,N_12462);
and U13150 (N_13150,N_9472,N_10726);
and U13151 (N_13151,N_10782,N_10930);
and U13152 (N_13152,N_10644,N_9623);
and U13153 (N_13153,N_10870,N_12224);
nor U13154 (N_13154,N_11765,N_11561);
or U13155 (N_13155,N_10207,N_10178);
or U13156 (N_13156,N_10124,N_12145);
or U13157 (N_13157,N_12427,N_11118);
nand U13158 (N_13158,N_12458,N_10215);
nand U13159 (N_13159,N_9699,N_10286);
nand U13160 (N_13160,N_11830,N_11128);
and U13161 (N_13161,N_11367,N_11915);
nor U13162 (N_13162,N_11895,N_9442);
nand U13163 (N_13163,N_10244,N_10583);
and U13164 (N_13164,N_12242,N_10144);
xor U13165 (N_13165,N_10652,N_9618);
and U13166 (N_13166,N_11312,N_11386);
nand U13167 (N_13167,N_11531,N_10075);
or U13168 (N_13168,N_10091,N_10135);
xor U13169 (N_13169,N_10520,N_11675);
or U13170 (N_13170,N_10130,N_9481);
nand U13171 (N_13171,N_9759,N_10892);
nand U13172 (N_13172,N_12308,N_10143);
nand U13173 (N_13173,N_10423,N_10250);
and U13174 (N_13174,N_11338,N_9801);
or U13175 (N_13175,N_10804,N_9544);
and U13176 (N_13176,N_11315,N_10185);
and U13177 (N_13177,N_12395,N_11459);
nor U13178 (N_13178,N_11079,N_11134);
xnor U13179 (N_13179,N_9541,N_11154);
and U13180 (N_13180,N_9454,N_10308);
or U13181 (N_13181,N_12473,N_11132);
and U13182 (N_13182,N_10374,N_10444);
nand U13183 (N_13183,N_10753,N_10489);
nor U13184 (N_13184,N_11719,N_10541);
nor U13185 (N_13185,N_9415,N_9620);
or U13186 (N_13186,N_9838,N_9505);
or U13187 (N_13187,N_10687,N_9594);
nand U13188 (N_13188,N_10518,N_10976);
xor U13189 (N_13189,N_12186,N_11044);
and U13190 (N_13190,N_10276,N_9596);
nor U13191 (N_13191,N_9754,N_11059);
nor U13192 (N_13192,N_11399,N_10593);
or U13193 (N_13193,N_10050,N_11309);
and U13194 (N_13194,N_11540,N_11648);
or U13195 (N_13195,N_11276,N_9979);
nor U13196 (N_13196,N_9525,N_10689);
nand U13197 (N_13197,N_9750,N_11122);
and U13198 (N_13198,N_11612,N_12097);
and U13199 (N_13199,N_10880,N_11903);
nand U13200 (N_13200,N_10723,N_10963);
nand U13201 (N_13201,N_11818,N_12454);
nand U13202 (N_13202,N_11819,N_9377);
and U13203 (N_13203,N_12300,N_12263);
and U13204 (N_13204,N_11334,N_11083);
xor U13205 (N_13205,N_10905,N_11652);
nor U13206 (N_13206,N_10863,N_10044);
and U13207 (N_13207,N_11832,N_10080);
nor U13208 (N_13208,N_11696,N_11139);
and U13209 (N_13209,N_10675,N_11140);
nand U13210 (N_13210,N_11335,N_11280);
nand U13211 (N_13211,N_11208,N_9752);
nand U13212 (N_13212,N_12221,N_9742);
nand U13213 (N_13213,N_9837,N_11088);
and U13214 (N_13214,N_11834,N_10556);
nand U13215 (N_13215,N_9650,N_10335);
nand U13216 (N_13216,N_10336,N_10899);
nand U13217 (N_13217,N_10163,N_10271);
nand U13218 (N_13218,N_9453,N_9710);
or U13219 (N_13219,N_12251,N_11408);
nand U13220 (N_13220,N_10882,N_10898);
nand U13221 (N_13221,N_10305,N_10132);
nand U13222 (N_13222,N_10048,N_11454);
nor U13223 (N_13223,N_11672,N_11019);
or U13224 (N_13224,N_9402,N_9560);
and U13225 (N_13225,N_12139,N_11277);
and U13226 (N_13226,N_11824,N_11329);
nor U13227 (N_13227,N_10138,N_12431);
and U13228 (N_13228,N_10747,N_11125);
nand U13229 (N_13229,N_11562,N_9884);
nor U13230 (N_13230,N_12096,N_11180);
nand U13231 (N_13231,N_10624,N_10941);
nor U13232 (N_13232,N_10861,N_10253);
nor U13233 (N_13233,N_10790,N_9730);
and U13234 (N_13234,N_9671,N_10647);
nand U13235 (N_13235,N_12049,N_9533);
nor U13236 (N_13236,N_9455,N_11594);
xnor U13237 (N_13237,N_10682,N_9755);
or U13238 (N_13238,N_11737,N_11889);
nor U13239 (N_13239,N_9873,N_11930);
and U13240 (N_13240,N_10022,N_10187);
nand U13241 (N_13241,N_10907,N_10877);
nand U13242 (N_13242,N_11984,N_10533);
nor U13243 (N_13243,N_11646,N_11422);
xor U13244 (N_13244,N_9462,N_12045);
nand U13245 (N_13245,N_11474,N_11974);
nor U13246 (N_13246,N_11593,N_9406);
nand U13247 (N_13247,N_10081,N_12351);
nor U13248 (N_13248,N_10807,N_10832);
nand U13249 (N_13249,N_11189,N_11291);
nand U13250 (N_13250,N_9822,N_12281);
or U13251 (N_13251,N_10351,N_10989);
and U13252 (N_13252,N_11060,N_12079);
nor U13253 (N_13253,N_9802,N_11056);
and U13254 (N_13254,N_10170,N_11421);
or U13255 (N_13255,N_10718,N_10674);
nand U13256 (N_13256,N_10849,N_9918);
xnor U13257 (N_13257,N_12130,N_12379);
nor U13258 (N_13258,N_9643,N_12094);
and U13259 (N_13259,N_12255,N_11860);
and U13260 (N_13260,N_11298,N_10961);
xnor U13261 (N_13261,N_9830,N_10551);
nor U13262 (N_13262,N_12299,N_11625);
nand U13263 (N_13263,N_12335,N_10226);
nand U13264 (N_13264,N_11622,N_12258);
and U13265 (N_13265,N_11825,N_11473);
xor U13266 (N_13266,N_11792,N_10600);
nor U13267 (N_13267,N_11828,N_10897);
and U13268 (N_13268,N_11339,N_10166);
and U13269 (N_13269,N_11143,N_9414);
or U13270 (N_13270,N_11723,N_9820);
nand U13271 (N_13271,N_10823,N_10814);
and U13272 (N_13272,N_11844,N_11274);
xnor U13273 (N_13273,N_10443,N_12426);
xnor U13274 (N_13274,N_10216,N_9723);
or U13275 (N_13275,N_11869,N_9796);
nor U13276 (N_13276,N_9506,N_11961);
xnor U13277 (N_13277,N_10663,N_9520);
and U13278 (N_13278,N_11866,N_12410);
nor U13279 (N_13279,N_12466,N_10448);
nor U13280 (N_13280,N_12089,N_10615);
nor U13281 (N_13281,N_10969,N_11038);
nor U13282 (N_13282,N_9628,N_11980);
nand U13283 (N_13283,N_11259,N_10808);
and U13284 (N_13284,N_11012,N_11294);
nor U13285 (N_13285,N_9768,N_10156);
and U13286 (N_13286,N_12023,N_12205);
nor U13287 (N_13287,N_11401,N_9894);
nor U13288 (N_13288,N_12268,N_12256);
nor U13289 (N_13289,N_10952,N_11142);
nand U13290 (N_13290,N_10590,N_11165);
or U13291 (N_13291,N_11507,N_11576);
nand U13292 (N_13292,N_10236,N_12026);
nor U13293 (N_13293,N_11990,N_10890);
or U13294 (N_13294,N_10490,N_10585);
or U13295 (N_13295,N_10089,N_9812);
or U13296 (N_13296,N_11332,N_9583);
or U13297 (N_13297,N_12042,N_11949);
and U13298 (N_13298,N_11161,N_11284);
or U13299 (N_13299,N_11959,N_11636);
or U13300 (N_13300,N_12168,N_10645);
nor U13301 (N_13301,N_9600,N_9471);
nor U13302 (N_13302,N_11376,N_10767);
xnor U13303 (N_13303,N_12339,N_11447);
and U13304 (N_13304,N_12279,N_9605);
and U13305 (N_13305,N_10695,N_10938);
nor U13306 (N_13306,N_10589,N_10289);
xor U13307 (N_13307,N_11746,N_11978);
or U13308 (N_13308,N_9535,N_10867);
nand U13309 (N_13309,N_9504,N_9632);
nor U13310 (N_13310,N_11896,N_10386);
or U13311 (N_13311,N_9772,N_10678);
and U13312 (N_13312,N_10800,N_11007);
and U13313 (N_13313,N_11385,N_9641);
nor U13314 (N_13314,N_10347,N_12013);
nand U13315 (N_13315,N_9713,N_11353);
or U13316 (N_13316,N_9619,N_10610);
nor U13317 (N_13317,N_11632,N_9507);
nand U13318 (N_13318,N_10015,N_12124);
nand U13319 (N_13319,N_11501,N_11528);
nand U13320 (N_13320,N_12066,N_11086);
nand U13321 (N_13321,N_10611,N_11023);
and U13322 (N_13322,N_10141,N_10442);
nand U13323 (N_13323,N_9933,N_10988);
nor U13324 (N_13324,N_11405,N_11349);
nand U13325 (N_13325,N_10004,N_11821);
or U13326 (N_13326,N_10492,N_11035);
nand U13327 (N_13327,N_10011,N_10200);
nand U13328 (N_13328,N_11977,N_11807);
nand U13329 (N_13329,N_11096,N_9502);
or U13330 (N_13330,N_10398,N_10172);
or U13331 (N_13331,N_9977,N_11242);
nor U13332 (N_13332,N_10754,N_10572);
nand U13333 (N_13333,N_9519,N_9756);
nor U13334 (N_13334,N_12194,N_12155);
xnor U13335 (N_13335,N_12114,N_10517);
and U13336 (N_13336,N_12450,N_11317);
nor U13337 (N_13337,N_12377,N_11112);
or U13338 (N_13338,N_12493,N_9479);
or U13339 (N_13339,N_9514,N_11330);
or U13340 (N_13340,N_9949,N_10150);
nand U13341 (N_13341,N_10294,N_10057);
xnor U13342 (N_13342,N_12336,N_11968);
xnor U13343 (N_13343,N_12063,N_10434);
nand U13344 (N_13344,N_10000,N_9652);
nand U13345 (N_13345,N_11411,N_10850);
nand U13346 (N_13346,N_11087,N_10355);
nand U13347 (N_13347,N_11141,N_9974);
and U13348 (N_13348,N_9622,N_11264);
nor U13349 (N_13349,N_10233,N_9937);
and U13350 (N_13350,N_9660,N_10149);
and U13351 (N_13351,N_10076,N_10389);
nor U13352 (N_13352,N_10725,N_12406);
or U13353 (N_13353,N_11460,N_11752);
nand U13354 (N_13354,N_9483,N_11103);
nand U13355 (N_13355,N_12322,N_10189);
xor U13356 (N_13356,N_10269,N_11475);
and U13357 (N_13357,N_10407,N_11287);
or U13358 (N_13358,N_11147,N_10735);
and U13359 (N_13359,N_9807,N_10119);
nor U13360 (N_13360,N_11224,N_11758);
nand U13361 (N_13361,N_12261,N_11697);
or U13362 (N_13362,N_11260,N_11168);
nor U13363 (N_13363,N_11503,N_11365);
nand U13364 (N_13364,N_11006,N_9867);
xnor U13365 (N_13365,N_11398,N_11919);
and U13366 (N_13366,N_12239,N_10887);
xnor U13367 (N_13367,N_10739,N_9781);
nand U13368 (N_13368,N_9712,N_11084);
or U13369 (N_13369,N_10377,N_10970);
nor U13370 (N_13370,N_11418,N_10816);
nor U13371 (N_13371,N_11799,N_11776);
xor U13372 (N_13372,N_10550,N_11852);
nand U13373 (N_13373,N_10323,N_9816);
and U13374 (N_13374,N_12173,N_9640);
nand U13375 (N_13375,N_9729,N_11355);
nand U13376 (N_13376,N_9603,N_10168);
and U13377 (N_13377,N_9978,N_10623);
nor U13378 (N_13378,N_11509,N_11888);
nor U13379 (N_13379,N_10945,N_9678);
nand U13380 (N_13380,N_11269,N_11282);
xnor U13381 (N_13381,N_10454,N_10307);
nor U13382 (N_13382,N_11607,N_11695);
nor U13383 (N_13383,N_9753,N_9470);
nor U13384 (N_13384,N_9956,N_9452);
or U13385 (N_13385,N_9612,N_10368);
nor U13386 (N_13386,N_11368,N_10979);
xnor U13387 (N_13387,N_11022,N_12472);
xor U13388 (N_13388,N_9787,N_9889);
or U13389 (N_13389,N_11693,N_9735);
nand U13390 (N_13390,N_11341,N_10241);
nand U13391 (N_13391,N_10959,N_10587);
or U13392 (N_13392,N_11183,N_11941);
and U13393 (N_13393,N_10010,N_9579);
nand U13394 (N_13394,N_12323,N_10160);
and U13395 (N_13395,N_10411,N_11254);
nand U13396 (N_13396,N_10826,N_10878);
xnor U13397 (N_13397,N_11031,N_10466);
and U13398 (N_13398,N_11745,N_9674);
xor U13399 (N_13399,N_10321,N_11967);
nor U13400 (N_13400,N_12028,N_10040);
nand U13401 (N_13401,N_11158,N_12179);
and U13402 (N_13402,N_10640,N_10035);
and U13403 (N_13403,N_12401,N_12329);
or U13404 (N_13404,N_12032,N_10300);
nand U13405 (N_13405,N_9848,N_9655);
or U13406 (N_13406,N_10196,N_10152);
nand U13407 (N_13407,N_11306,N_10030);
xor U13408 (N_13408,N_12337,N_9378);
xor U13409 (N_13409,N_11635,N_12457);
nor U13410 (N_13410,N_9707,N_10575);
nand U13411 (N_13411,N_10918,N_11921);
or U13412 (N_13412,N_10254,N_10209);
nand U13413 (N_13413,N_9711,N_11766);
and U13414 (N_13414,N_12018,N_11431);
and U13415 (N_13415,N_9944,N_12232);
or U13416 (N_13416,N_10068,N_10157);
or U13417 (N_13417,N_10717,N_11822);
nand U13418 (N_13418,N_10021,N_11519);
xor U13419 (N_13419,N_9738,N_11169);
or U13420 (N_13420,N_11987,N_9469);
xnor U13421 (N_13421,N_10962,N_12160);
and U13422 (N_13422,N_11272,N_10327);
nand U13423 (N_13423,N_11025,N_10264);
nor U13424 (N_13424,N_12316,N_11761);
nor U13425 (N_13425,N_10199,N_12328);
nand U13426 (N_13426,N_10914,N_11606);
nand U13427 (N_13427,N_11382,N_9885);
and U13428 (N_13428,N_11063,N_10134);
or U13429 (N_13429,N_10972,N_9380);
nand U13430 (N_13430,N_10620,N_9706);
and U13431 (N_13431,N_10708,N_11564);
nor U13432 (N_13432,N_11384,N_11156);
nor U13433 (N_13433,N_10338,N_12348);
or U13434 (N_13434,N_11430,N_11111);
xnor U13435 (N_13435,N_11909,N_9722);
and U13436 (N_13436,N_11455,N_11744);
nor U13437 (N_13437,N_11417,N_9682);
and U13438 (N_13438,N_11081,N_10437);
nor U13439 (N_13439,N_10752,N_10053);
xor U13440 (N_13440,N_9569,N_11360);
nand U13441 (N_13441,N_10527,N_11052);
and U13442 (N_13442,N_10256,N_10123);
nand U13443 (N_13443,N_10175,N_10396);
nor U13444 (N_13444,N_11767,N_12471);
nor U13445 (N_13445,N_9748,N_9746);
or U13446 (N_13446,N_9984,N_10802);
xnor U13447 (N_13447,N_9734,N_9554);
nand U13448 (N_13448,N_9493,N_11177);
or U13449 (N_13449,N_10911,N_12010);
and U13450 (N_13450,N_10522,N_10992);
and U13451 (N_13451,N_10756,N_11397);
nand U13452 (N_13452,N_10858,N_9382);
nor U13453 (N_13453,N_10416,N_11928);
or U13454 (N_13454,N_11623,N_11771);
nor U13455 (N_13455,N_11850,N_9664);
nor U13456 (N_13456,N_11493,N_9835);
or U13457 (N_13457,N_12315,N_9425);
or U13458 (N_13458,N_11898,N_12127);
and U13459 (N_13459,N_9954,N_12468);
nor U13460 (N_13460,N_9736,N_11893);
or U13461 (N_13461,N_9823,N_11720);
nor U13462 (N_13462,N_11544,N_11175);
xor U13463 (N_13463,N_10559,N_10953);
or U13464 (N_13464,N_12306,N_9904);
nand U13465 (N_13465,N_9546,N_9686);
nand U13466 (N_13466,N_12065,N_10117);
and U13467 (N_13467,N_12262,N_12384);
or U13468 (N_13468,N_11106,N_10213);
and U13469 (N_13469,N_10651,N_9747);
and U13470 (N_13470,N_9804,N_10671);
nor U13471 (N_13471,N_10174,N_11983);
nor U13472 (N_13472,N_11811,N_10420);
nor U13473 (N_13473,N_12332,N_11305);
and U13474 (N_13474,N_10096,N_9961);
and U13475 (N_13475,N_9886,N_12386);
nand U13476 (N_13476,N_10228,N_9855);
or U13477 (N_13477,N_10908,N_10609);
nor U13478 (N_13478,N_10996,N_9902);
or U13479 (N_13479,N_10453,N_10484);
and U13480 (N_13480,N_10285,N_9788);
or U13481 (N_13481,N_12437,N_10309);
nand U13482 (N_13482,N_11611,N_12361);
or U13483 (N_13483,N_9896,N_12284);
and U13484 (N_13484,N_11520,N_9775);
and U13485 (N_13485,N_10201,N_10744);
and U13486 (N_13486,N_12175,N_9765);
nor U13487 (N_13487,N_9824,N_11989);
or U13488 (N_13488,N_11434,N_10026);
or U13489 (N_13489,N_11002,N_9913);
nor U13490 (N_13490,N_12121,N_10387);
nand U13491 (N_13491,N_12008,N_10626);
nand U13492 (N_13492,N_10419,N_10239);
and U13493 (N_13493,N_11380,N_11197);
or U13494 (N_13494,N_11200,N_11041);
nand U13495 (N_13495,N_11548,N_10839);
nand U13496 (N_13496,N_11993,N_9408);
and U13497 (N_13497,N_12091,N_9860);
or U13498 (N_13498,N_9872,N_11020);
nor U13499 (N_13499,N_10760,N_11795);
nor U13500 (N_13500,N_9630,N_12420);
and U13501 (N_13501,N_10825,N_9920);
nor U13502 (N_13502,N_10924,N_10188);
nand U13503 (N_13503,N_12272,N_10669);
or U13504 (N_13504,N_9391,N_10488);
nor U13505 (N_13505,N_11190,N_10926);
and U13506 (N_13506,N_12083,N_11651);
and U13507 (N_13507,N_11452,N_9498);
or U13508 (N_13508,N_11377,N_12418);
or U13509 (N_13509,N_11392,N_9458);
or U13510 (N_13510,N_10635,N_10643);
and U13511 (N_13511,N_12050,N_10709);
nand U13512 (N_13512,N_11848,N_9809);
nor U13513 (N_13513,N_11586,N_10008);
or U13514 (N_13514,N_9880,N_9489);
xnor U13515 (N_13515,N_12198,N_9986);
nor U13516 (N_13516,N_9441,N_9790);
nand U13517 (N_13517,N_12307,N_11997);
or U13518 (N_13518,N_11820,N_9862);
and U13519 (N_13519,N_12120,N_11414);
nand U13520 (N_13520,N_11130,N_11319);
xnor U13521 (N_13521,N_10432,N_11311);
nor U13522 (N_13522,N_9976,N_10194);
nand U13523 (N_13523,N_10281,N_10649);
or U13524 (N_13524,N_11655,N_12225);
nand U13525 (N_13525,N_11324,N_10716);
and U13526 (N_13526,N_9741,N_9785);
and U13527 (N_13527,N_11359,N_9964);
and U13528 (N_13528,N_12185,N_11346);
xor U13529 (N_13529,N_12247,N_11985);
and U13530 (N_13530,N_10906,N_10066);
nand U13531 (N_13531,N_11166,N_9688);
nor U13532 (N_13532,N_10554,N_9659);
nand U13533 (N_13533,N_11004,N_12101);
and U13534 (N_13534,N_12218,N_11135);
and U13535 (N_13535,N_11313,N_10310);
and U13536 (N_13536,N_11589,N_9718);
nand U13537 (N_13537,N_12073,N_10872);
nor U13538 (N_13538,N_12259,N_11605);
nor U13539 (N_13539,N_10919,N_11876);
nand U13540 (N_13540,N_11739,N_12305);
and U13541 (N_13541,N_12345,N_11992);
or U13542 (N_13542,N_9524,N_10121);
xor U13543 (N_13543,N_10565,N_11217);
and U13544 (N_13544,N_12357,N_10158);
nand U13545 (N_13545,N_9611,N_12366);
nor U13546 (N_13546,N_10441,N_9758);
nand U13547 (N_13547,N_11410,N_10279);
or U13548 (N_13548,N_12072,N_12237);
and U13549 (N_13549,N_12215,N_11845);
nor U13550 (N_13550,N_12429,N_11512);
or U13551 (N_13551,N_11362,N_10145);
nand U13552 (N_13552,N_11069,N_9926);
nand U13553 (N_13553,N_10095,N_12119);
xnor U13554 (N_13554,N_12222,N_10006);
and U13555 (N_13555,N_9637,N_9973);
nand U13556 (N_13556,N_9960,N_10342);
nor U13557 (N_13557,N_11227,N_11741);
nor U13558 (N_13558,N_10701,N_9598);
xor U13559 (N_13559,N_11511,N_9975);
or U13560 (N_13560,N_11699,N_9457);
or U13561 (N_13561,N_12136,N_10344);
nor U13562 (N_13562,N_9792,N_9539);
nor U13563 (N_13563,N_9438,N_10501);
and U13564 (N_13564,N_12494,N_9875);
nor U13565 (N_13565,N_12452,N_11614);
or U13566 (N_13566,N_11712,N_9537);
or U13567 (N_13567,N_11547,N_11234);
nor U13568 (N_13568,N_9866,N_10410);
nor U13569 (N_13569,N_10547,N_10139);
nand U13570 (N_13570,N_10596,N_11630);
or U13571 (N_13571,N_12233,N_12385);
and U13572 (N_13572,N_11748,N_10935);
and U13573 (N_13573,N_11929,N_9581);
or U13574 (N_13574,N_11706,N_12317);
nor U13575 (N_13575,N_11743,N_10942);
nand U13576 (N_13576,N_11523,N_9805);
and U13577 (N_13577,N_11491,N_9528);
xnor U13578 (N_13578,N_10857,N_10328);
nand U13579 (N_13579,N_9925,N_11808);
and U13580 (N_13580,N_10126,N_11692);
nand U13581 (N_13581,N_10766,N_12109);
nand U13582 (N_13582,N_10415,N_10110);
or U13583 (N_13583,N_11407,N_12297);
or U13584 (N_13584,N_11068,N_12344);
and U13585 (N_13585,N_11527,N_12321);
or U13586 (N_13586,N_10542,N_9614);
xnor U13587 (N_13587,N_12116,N_11199);
and U13588 (N_13588,N_10104,N_12085);
nor U13589 (N_13589,N_9731,N_9727);
or U13590 (N_13590,N_11292,N_11817);
or U13591 (N_13591,N_9424,N_9863);
or U13592 (N_13592,N_11979,N_9609);
nor U13593 (N_13593,N_10449,N_11490);
nor U13594 (N_13594,N_10282,N_10506);
and U13595 (N_13595,N_10181,N_11793);
or U13596 (N_13596,N_9966,N_10686);
or U13597 (N_13597,N_9708,N_11050);
or U13598 (N_13598,N_11258,N_9496);
nor U13599 (N_13599,N_12246,N_9851);
and U13600 (N_13600,N_10301,N_12481);
nor U13601 (N_13601,N_10940,N_11205);
or U13602 (N_13602,N_11687,N_11679);
or U13603 (N_13603,N_9914,N_12485);
and U13604 (N_13604,N_10680,N_11546);
nand U13605 (N_13605,N_10692,N_10176);
and U13606 (N_13606,N_10673,N_11082);
nor U13607 (N_13607,N_11097,N_12436);
and U13608 (N_13608,N_11971,N_12446);
nand U13609 (N_13609,N_11518,N_11716);
nand U13610 (N_13610,N_11196,N_10824);
or U13611 (N_13611,N_11560,N_9909);
xnor U13612 (N_13612,N_11320,N_9626);
and U13613 (N_13613,N_10088,N_12167);
and U13614 (N_13614,N_12180,N_10950);
and U13615 (N_13615,N_10771,N_9932);
xor U13616 (N_13616,N_9677,N_10212);
or U13617 (N_13617,N_11965,N_9870);
and U13618 (N_13618,N_9575,N_10820);
nand U13619 (N_13619,N_11619,N_10562);
xor U13620 (N_13620,N_10097,N_11951);
nor U13621 (N_13621,N_11912,N_10225);
or U13622 (N_13622,N_11351,N_11890);
nor U13623 (N_13623,N_10409,N_11892);
nand U13624 (N_13624,N_12238,N_9576);
and U13625 (N_13625,N_12059,N_11861);
nand U13626 (N_13626,N_12376,N_11797);
nand U13627 (N_13627,N_11914,N_9672);
or U13628 (N_13628,N_9774,N_9431);
nand U13629 (N_13629,N_11034,N_12040);
or U13630 (N_13630,N_11703,N_11395);
xnor U13631 (N_13631,N_12303,N_11801);
and U13632 (N_13632,N_9463,N_11521);
nand U13633 (N_13633,N_11722,N_11910);
or U13634 (N_13634,N_11090,N_11982);
or U13635 (N_13635,N_9955,N_10955);
nand U13636 (N_13636,N_9828,N_9543);
or U13637 (N_13637,N_9585,N_9407);
nor U13638 (N_13638,N_10628,N_10340);
xnor U13639 (N_13639,N_11877,N_9757);
xnor U13640 (N_13640,N_9602,N_11867);
nand U13641 (N_13641,N_11204,N_10720);
or U13642 (N_13642,N_12441,N_11220);
xor U13643 (N_13643,N_9777,N_10662);
xnor U13644 (N_13644,N_9697,N_11729);
nor U13645 (N_13645,N_11481,N_9553);
nand U13646 (N_13646,N_10148,N_11774);
or U13647 (N_13647,N_12062,N_10392);
nand U13648 (N_13648,N_11626,N_12244);
or U13649 (N_13649,N_11449,N_10070);
or U13650 (N_13650,N_9721,N_11155);
and U13651 (N_13651,N_9767,N_9947);
or U13652 (N_13652,N_10862,N_12078);
nor U13653 (N_13653,N_10313,N_10043);
nand U13654 (N_13654,N_9646,N_11228);
and U13655 (N_13655,N_11256,N_9690);
nand U13656 (N_13656,N_9891,N_11378);
or U13657 (N_13657,N_9912,N_9946);
or U13658 (N_13658,N_10987,N_9931);
and U13659 (N_13659,N_12236,N_9842);
and U13660 (N_13660,N_10846,N_10539);
and U13661 (N_13661,N_10033,N_12492);
and U13662 (N_13662,N_9846,N_11243);
xor U13663 (N_13663,N_9557,N_12152);
nand U13664 (N_13664,N_9478,N_11833);
nand U13665 (N_13665,N_11262,N_12331);
or U13666 (N_13666,N_10588,N_10023);
nand U13667 (N_13667,N_11669,N_10504);
xnor U13668 (N_13668,N_10946,N_11472);
and U13669 (N_13669,N_9392,N_10712);
nand U13670 (N_13670,N_11725,N_10734);
or U13671 (N_13671,N_12409,N_11342);
nor U13672 (N_13672,N_10621,N_9853);
or U13673 (N_13673,N_9495,N_10238);
or U13674 (N_13674,N_9684,N_10020);
nand U13675 (N_13675,N_12147,N_12304);
or U13676 (N_13676,N_9784,N_11178);
nand U13677 (N_13677,N_10364,N_12422);
nand U13678 (N_13678,N_11458,N_11049);
or U13679 (N_13679,N_10921,N_11917);
and U13680 (N_13680,N_9561,N_10592);
nand U13681 (N_13681,N_9608,N_11316);
and U13682 (N_13682,N_9665,N_12414);
nand U13683 (N_13683,N_11223,N_12190);
and U13684 (N_13684,N_10102,N_11938);
and U13685 (N_13685,N_12375,N_11539);
and U13686 (N_13686,N_10051,N_11796);
and U13687 (N_13687,N_9661,N_10031);
nand U13688 (N_13688,N_10868,N_12204);
nand U13689 (N_13689,N_10511,N_11461);
and U13690 (N_13690,N_10147,N_12364);
nor U13691 (N_13691,N_11710,N_11137);
nor U13692 (N_13692,N_12209,N_12153);
or U13693 (N_13693,N_10917,N_11054);
nand U13694 (N_13694,N_10659,N_11268);
nand U13695 (N_13695,N_11109,N_12132);
nand U13696 (N_13696,N_9936,N_11517);
nand U13697 (N_13697,N_9451,N_10727);
nand U13698 (N_13698,N_10761,N_11998);
xnor U13699 (N_13699,N_9815,N_10577);
nand U13700 (N_13700,N_9563,N_10966);
xnor U13701 (N_13701,N_10373,N_10672);
or U13702 (N_13702,N_12499,N_12475);
nand U13703 (N_13703,N_10944,N_12016);
or U13704 (N_13704,N_10841,N_9419);
or U13705 (N_13705,N_10046,N_11620);
nand U13706 (N_13706,N_9625,N_9845);
and U13707 (N_13707,N_12383,N_11429);
nor U13708 (N_13708,N_11682,N_11757);
xor U13709 (N_13709,N_11047,N_11246);
and U13710 (N_13710,N_11641,N_10787);
nand U13711 (N_13711,N_12479,N_9943);
xor U13712 (N_13712,N_10332,N_12183);
nor U13713 (N_13713,N_12200,N_9649);
and U13714 (N_13714,N_10548,N_11437);
nor U13715 (N_13715,N_10125,N_9849);
nand U13716 (N_13716,N_12217,N_11805);
and U13717 (N_13717,N_10291,N_10001);
xor U13718 (N_13718,N_10084,N_11448);
xnor U13719 (N_13719,N_12290,N_10809);
xnor U13720 (N_13720,N_11212,N_12093);
xor U13721 (N_13721,N_12400,N_12219);
and U13722 (N_13722,N_9376,N_12071);
or U13723 (N_13723,N_11092,N_11477);
nand U13724 (N_13724,N_12443,N_12314);
nor U13725 (N_13725,N_11847,N_9841);
and U13726 (N_13726,N_10447,N_9898);
or U13727 (N_13727,N_10637,N_9667);
and U13728 (N_13728,N_12275,N_10367);
nor U13729 (N_13729,N_11489,N_11553);
and U13730 (N_13730,N_11638,N_11906);
nor U13731 (N_13731,N_12496,N_12041);
and U13732 (N_13732,N_9840,N_10064);
or U13733 (N_13733,N_11394,N_9562);
nor U13734 (N_13734,N_10801,N_12469);
xnor U13735 (N_13735,N_9634,N_10099);
or U13736 (N_13736,N_10353,N_11668);
and U13737 (N_13737,N_10372,N_11631);
xor U13738 (N_13738,N_11283,N_11841);
xor U13739 (N_13739,N_10151,N_10510);
and U13740 (N_13740,N_12301,N_11451);
or U13741 (N_13741,N_10440,N_10707);
and U13742 (N_13742,N_12269,N_10190);
nor U13743 (N_13743,N_10456,N_12157);
nor U13744 (N_13744,N_10049,N_10283);
or U13745 (N_13745,N_12054,N_10842);
xor U13746 (N_13746,N_10358,N_9988);
or U13747 (N_13747,N_9656,N_12319);
or U13748 (N_13748,N_11568,N_11925);
and U13749 (N_13749,N_9908,N_9819);
nor U13750 (N_13750,N_12380,N_10433);
xor U13751 (N_13751,N_10237,N_9694);
and U13752 (N_13752,N_11629,N_9938);
or U13753 (N_13753,N_12140,N_10691);
or U13754 (N_13754,N_11785,N_12133);
or U13755 (N_13755,N_10855,N_9416);
or U13756 (N_13756,N_12125,N_9383);
nor U13757 (N_13757,N_10632,N_10191);
or U13758 (N_13758,N_12080,N_11911);
nor U13759 (N_13759,N_12228,N_12271);
and U13760 (N_13760,N_12077,N_12161);
or U13761 (N_13761,N_11065,N_9743);
nand U13762 (N_13762,N_12201,N_12392);
nand U13763 (N_13763,N_10017,N_11211);
nand U13764 (N_13764,N_11592,N_10888);
nor U13765 (N_13765,N_11551,N_10348);
nor U13766 (N_13766,N_11465,N_10246);
xnor U13767 (N_13767,N_12007,N_10773);
nand U13768 (N_13768,N_11248,N_11536);
and U13769 (N_13769,N_10261,N_12291);
nor U13770 (N_13770,N_11021,N_11297);
nand U13771 (N_13771,N_11857,N_10758);
or U13772 (N_13772,N_10853,N_9998);
or U13773 (N_13773,N_9704,N_11107);
nor U13774 (N_13774,N_10696,N_12034);
nor U13775 (N_13775,N_12311,N_9778);
xor U13776 (N_13776,N_12372,N_11816);
and U13777 (N_13777,N_11424,N_9564);
nand U13778 (N_13778,N_10664,N_10324);
nand U13779 (N_13779,N_10567,N_12425);
nand U13780 (N_13780,N_9970,N_11406);
and U13781 (N_13781,N_11839,N_12207);
or U13782 (N_13782,N_9676,N_10884);
or U13783 (N_13783,N_10224,N_9491);
nand U13784 (N_13784,N_10083,N_11198);
nor U13785 (N_13785,N_10290,N_9405);
or U13786 (N_13786,N_11040,N_11463);
or U13787 (N_13787,N_10785,N_11352);
nor U13788 (N_13788,N_11944,N_10813);
nor U13789 (N_13789,N_11788,N_12108);
nand U13790 (N_13790,N_11995,N_10109);
nor U13791 (N_13791,N_11934,N_11731);
or U13792 (N_13792,N_10093,N_11708);
nand U13793 (N_13793,N_11779,N_11782);
and U13794 (N_13794,N_9733,N_11373);
nor U13795 (N_13795,N_9591,N_12318);
or U13796 (N_13796,N_9702,N_10258);
nor U13797 (N_13797,N_10700,N_11814);
and U13798 (N_13798,N_11610,N_11525);
or U13799 (N_13799,N_10263,N_11653);
and U13800 (N_13800,N_10018,N_12187);
nand U13801 (N_13801,N_11514,N_9542);
xnor U13802 (N_13802,N_9906,N_9381);
nor U13803 (N_13803,N_10634,N_11836);
nor U13804 (N_13804,N_9617,N_11730);
and U13805 (N_13805,N_11803,N_9923);
and U13806 (N_13806,N_9663,N_9980);
xnor U13807 (N_13807,N_11051,N_10597);
xnor U13808 (N_13808,N_11027,N_12404);
or U13809 (N_13809,N_11587,N_11942);
or U13810 (N_13810,N_10431,N_10002);
nand U13811 (N_13811,N_10019,N_12411);
nand U13812 (N_13812,N_12342,N_12004);
nor U13813 (N_13813,N_11016,N_10552);
and U13814 (N_13814,N_10467,N_11100);
nand U13815 (N_13815,N_12302,N_10037);
or U13816 (N_13816,N_10272,N_9571);
and U13817 (N_13817,N_11773,N_11691);
or U13818 (N_13818,N_11162,N_11470);
nand U13819 (N_13819,N_10371,N_12359);
and U13820 (N_13820,N_11645,N_11445);
and U13821 (N_13821,N_11383,N_10764);
nand U13822 (N_13822,N_10495,N_11678);
nand U13823 (N_13823,N_11487,N_12067);
nand U13824 (N_13824,N_11300,N_12399);
or U13825 (N_13825,N_11905,N_11241);
xnor U13826 (N_13826,N_11261,N_11482);
nor U13827 (N_13827,N_11760,N_12347);
xor U13828 (N_13828,N_9401,N_12100);
or U13829 (N_13829,N_11492,N_10786);
nor U13830 (N_13830,N_10498,N_10464);
xor U13831 (N_13831,N_10901,N_10186);
nand U13832 (N_13832,N_12055,N_11307);
and U13833 (N_13833,N_10837,N_9716);
xnor U13834 (N_13834,N_11870,N_10852);
nor U13835 (N_13835,N_9720,N_11878);
and U13836 (N_13836,N_11428,N_11918);
nor U13837 (N_13837,N_12075,N_10731);
nor U13838 (N_13838,N_12029,N_12170);
xnor U13839 (N_13839,N_12327,N_10983);
nor U13840 (N_13840,N_12092,N_9890);
nor U13841 (N_13841,N_12320,N_11513);
or U13842 (N_13842,N_12257,N_10544);
and U13843 (N_13843,N_9521,N_12356);
nor U13844 (N_13844,N_9857,N_9460);
and U13845 (N_13845,N_12389,N_12402);
or U13846 (N_13846,N_11554,N_11534);
xnor U13847 (N_13847,N_10016,N_9762);
nor U13848 (N_13848,N_10485,N_9573);
xor U13849 (N_13849,N_11469,N_10793);
nand U13850 (N_13850,N_10500,N_9466);
nand U13851 (N_13851,N_10954,N_10265);
and U13852 (N_13852,N_10894,N_12146);
nand U13853 (N_13853,N_11119,N_10779);
nor U13854 (N_13854,N_10435,N_11184);
and U13855 (N_13855,N_10728,N_12333);
nor U13856 (N_13856,N_11182,N_11193);
nand U13857 (N_13857,N_10408,N_10183);
nor U13858 (N_13858,N_11994,N_9497);
or U13859 (N_13859,N_11440,N_12188);
or U13860 (N_13860,N_11791,N_11871);
or U13861 (N_13861,N_12456,N_11637);
or U13862 (N_13862,N_12463,N_11146);
or U13863 (N_13863,N_10394,N_11954);
and U13864 (N_13864,N_12112,N_11438);
xnor U13865 (N_13865,N_9607,N_11113);
nand U13866 (N_13866,N_9403,N_10711);
or U13867 (N_13867,N_9972,N_11333);
or U13868 (N_13868,N_12122,N_11975);
xnor U13869 (N_13869,N_12107,N_11916);
nor U13870 (N_13870,N_12371,N_9580);
nand U13871 (N_13871,N_10986,N_9459);
or U13872 (N_13872,N_11726,N_11849);
and U13873 (N_13873,N_9797,N_11750);
or U13874 (N_13874,N_11581,N_11266);
or U13875 (N_13875,N_10013,N_10694);
nor U13876 (N_13876,N_9703,N_9959);
nand U13877 (N_13877,N_9388,N_9486);
nor U13878 (N_13878,N_12158,N_10003);
nor U13879 (N_13879,N_10316,N_10063);
nor U13880 (N_13880,N_10512,N_9427);
nand U13881 (N_13881,N_11115,N_9780);
xnor U13882 (N_13882,N_10830,N_12131);
nor U13883 (N_13883,N_9433,N_9499);
nand U13884 (N_13884,N_10234,N_10915);
nor U13885 (N_13885,N_11718,N_11379);
nor U13886 (N_13886,N_12288,N_11310);
nor U13887 (N_13887,N_11664,N_10798);
nor U13888 (N_13888,N_10943,N_12338);
nand U13889 (N_13889,N_9549,N_11683);
nor U13890 (N_13890,N_12491,N_10370);
or U13891 (N_13891,N_9645,N_10481);
nand U13892 (N_13892,N_12150,N_12283);
nand U13893 (N_13893,N_9856,N_11058);
nand U13894 (N_13894,N_12298,N_10382);
or U13895 (N_13895,N_9474,N_10140);
or U13896 (N_13896,N_10365,N_10690);
or U13897 (N_13897,N_12394,N_10128);
or U13898 (N_13898,N_11613,N_11450);
nand U13899 (N_13899,N_11237,N_10399);
nor U13900 (N_13900,N_9843,N_10028);
nand U13901 (N_13901,N_9435,N_10715);
xnor U13902 (N_13902,N_11101,N_11727);
nor U13903 (N_13903,N_11950,N_9647);
nor U13904 (N_13904,N_12367,N_10561);
nor U13905 (N_13905,N_11093,N_9854);
and U13906 (N_13906,N_9555,N_9948);
xor U13907 (N_13907,N_12051,N_11759);
and U13908 (N_13908,N_12022,N_10330);
and U13909 (N_13909,N_10260,N_10602);
or U13910 (N_13910,N_11014,N_12082);
nand U13911 (N_13911,N_11621,N_10967);
or U13912 (N_13912,N_9393,N_10681);
nor U13913 (N_13913,N_10876,N_10403);
nor U13914 (N_13914,N_10195,N_9911);
xor U13915 (N_13915,N_10667,N_10665);
or U13916 (N_13916,N_10925,N_11391);
or U13917 (N_13917,N_12199,N_10975);
nand U13918 (N_13918,N_9437,N_10958);
and U13919 (N_13919,N_11159,N_11017);
xnor U13920 (N_13920,N_12486,N_11963);
nor U13921 (N_13921,N_10105,N_9951);
or U13922 (N_13922,N_11972,N_9850);
or U13923 (N_13923,N_11425,N_12035);
nor U13924 (N_13924,N_12487,N_12390);
or U13925 (N_13925,N_9887,N_10654);
xor U13926 (N_13926,N_11120,N_11363);
and U13927 (N_13927,N_10699,N_9693);
and U13928 (N_13928,N_10883,N_9409);
nand U13929 (N_13929,N_11066,N_12142);
and U13930 (N_13930,N_12015,N_11480);
or U13931 (N_13931,N_10494,N_10540);
nand U13932 (N_13932,N_11409,N_10641);
xnor U13933 (N_13933,N_12110,N_12099);
and U13934 (N_13934,N_10317,N_11988);
or U13935 (N_13935,N_10413,N_12129);
and U13936 (N_13936,N_12382,N_10847);
xor U13937 (N_13937,N_9769,N_10844);
or U13938 (N_13938,N_9559,N_12460);
nand U13939 (N_13939,N_11453,N_11865);
and U13940 (N_13940,N_11946,N_11252);
xnor U13941 (N_13941,N_12068,N_9420);
nor U13942 (N_13942,N_9989,N_11302);
xor U13943 (N_13943,N_12449,N_10947);
nand U13944 (N_13944,N_12012,N_10957);
or U13945 (N_13945,N_10337,N_10384);
and U13946 (N_13946,N_11721,N_10661);
nor U13947 (N_13947,N_9744,N_12408);
or U13948 (N_13948,N_9527,N_12021);
nor U13949 (N_13949,N_10418,N_10114);
or U13950 (N_13950,N_10912,N_10537);
nand U13951 (N_13951,N_9395,N_12495);
or U13952 (N_13952,N_11225,N_11883);
or U13953 (N_13953,N_10939,N_9839);
xor U13954 (N_13954,N_11713,N_11563);
or U13955 (N_13955,N_9523,N_11777);
or U13956 (N_13956,N_9685,N_11250);
nand U13957 (N_13957,N_10320,N_10329);
xnor U13958 (N_13958,N_12226,N_9725);
nor U13959 (N_13959,N_10472,N_11347);
and U13960 (N_13960,N_12424,N_10546);
or U13961 (N_13961,N_10197,N_12052);
and U13962 (N_13962,N_9412,N_10928);
nand U13963 (N_13963,N_12189,N_9994);
nand U13964 (N_13964,N_11868,N_10459);
or U13965 (N_13965,N_10401,N_11666);
and U13966 (N_13966,N_10153,N_10834);
nand U13967 (N_13967,N_11500,N_9715);
xor U13968 (N_13968,N_11676,N_10424);
and U13969 (N_13969,N_11559,N_11350);
or U13970 (N_13970,N_11381,N_9760);
and U13971 (N_13971,N_9396,N_9924);
nand U13972 (N_13972,N_11029,N_10069);
or U13973 (N_13973,N_10452,N_9963);
or U13974 (N_13974,N_12477,N_10071);
xor U13975 (N_13975,N_10772,N_11479);
nand U13976 (N_13976,N_11899,N_11939);
and U13977 (N_13977,N_9818,N_12005);
and U13978 (N_13978,N_9490,N_9881);
or U13979 (N_13979,N_11644,N_9903);
nand U13980 (N_13980,N_10900,N_11327);
nand U13981 (N_13981,N_12391,N_10625);
nand U13982 (N_13982,N_9668,N_11670);
xor U13983 (N_13983,N_11732,N_10349);
nand U13984 (N_13984,N_10657,N_10497);
nand U13985 (N_13985,N_10235,N_11763);
nand U13986 (N_13986,N_9639,N_11174);
nor U13987 (N_13987,N_10789,N_12374);
and U13988 (N_13988,N_10078,N_10311);
nor U13989 (N_13989,N_10251,N_11781);
nor U13990 (N_13990,N_11661,N_12214);
or U13991 (N_13991,N_11897,N_11837);
or U13992 (N_13992,N_10451,N_11591);
or U13993 (N_13993,N_10705,N_9952);
and U13994 (N_13994,N_9968,N_10227);
or U13995 (N_13995,N_11826,N_10487);
nor U13996 (N_13996,N_11556,N_10455);
nand U13997 (N_13997,N_12419,N_10029);
and U13998 (N_13998,N_11647,N_10356);
and U13999 (N_13999,N_10555,N_10714);
or U14000 (N_14000,N_10073,N_11037);
nor U14001 (N_14001,N_10363,N_11502);
nor U14002 (N_14002,N_11340,N_11535);
or U14003 (N_14003,N_12076,N_12033);
nor U14004 (N_14004,N_10655,N_11907);
nor U14005 (N_14005,N_10159,N_10697);
xnor U14006 (N_14006,N_9450,N_11296);
or U14007 (N_14007,N_10994,N_10032);
or U14008 (N_14008,N_9633,N_9847);
or U14009 (N_14009,N_9953,N_10350);
nand U14010 (N_14010,N_11778,N_10385);
nor U14011 (N_14011,N_10306,N_12003);
nor U14012 (N_14012,N_10614,N_10923);
and U14013 (N_14013,N_11580,N_10581);
or U14014 (N_14014,N_9858,N_12163);
and U14015 (N_14015,N_9518,N_9897);
and U14016 (N_14016,N_10679,N_9763);
or U14017 (N_14017,N_11271,N_11247);
nor U14018 (N_14018,N_10304,N_12105);
nand U14019 (N_14019,N_11628,N_10936);
or U14020 (N_14020,N_9572,N_9997);
and U14021 (N_14021,N_12451,N_9719);
and U14022 (N_14022,N_9705,N_11690);
and U14023 (N_14023,N_12103,N_10257);
and U14024 (N_14024,N_9429,N_9888);
and U14025 (N_14025,N_9552,N_11476);
and U14026 (N_14026,N_10293,N_11201);
xor U14027 (N_14027,N_11885,N_11715);
nor U14028 (N_14028,N_10229,N_10743);
nor U14029 (N_14029,N_12387,N_10220);
nand U14030 (N_14030,N_11191,N_12296);
or U14031 (N_14031,N_9428,N_11032);
or U14032 (N_14032,N_9631,N_9882);
nor U14033 (N_14033,N_10982,N_12223);
nor U14034 (N_14034,N_10803,N_11764);
nor U14035 (N_14035,N_10848,N_10314);
xnor U14036 (N_14036,N_10896,N_12396);
or U14037 (N_14037,N_9681,N_10103);
nand U14038 (N_14038,N_10036,N_9833);
nor U14039 (N_14039,N_10240,N_9476);
and U14040 (N_14040,N_10759,N_12162);
nand U14041 (N_14041,N_11840,N_9905);
or U14042 (N_14042,N_11880,N_9436);
and U14043 (N_14043,N_10115,N_12370);
xor U14044 (N_14044,N_11602,N_11709);
or U14045 (N_14045,N_10932,N_10060);
or U14046 (N_14046,N_10630,N_12088);
nand U14047 (N_14047,N_10056,N_9687);
and U14048 (N_14048,N_10557,N_10937);
or U14049 (N_14049,N_11550,N_12184);
xor U14050 (N_14050,N_11457,N_9927);
or U14051 (N_14051,N_9869,N_11008);
nand U14052 (N_14052,N_11026,N_10993);
nand U14053 (N_14053,N_10266,N_12421);
nand U14054 (N_14054,N_10214,N_11624);
nand U14055 (N_14055,N_10612,N_9418);
nor U14056 (N_14056,N_11321,N_10603);
nand U14057 (N_14057,N_11881,N_10750);
nand U14058 (N_14058,N_12061,N_10165);
or U14059 (N_14059,N_12128,N_11203);
or U14060 (N_14060,N_11393,N_12388);
or U14061 (N_14061,N_10931,N_11684);
nor U14062 (N_14062,N_10949,N_12012);
and U14063 (N_14063,N_12339,N_11865);
or U14064 (N_14064,N_11172,N_10312);
nor U14065 (N_14065,N_10487,N_10017);
nor U14066 (N_14066,N_12237,N_9989);
or U14067 (N_14067,N_10014,N_11852);
or U14068 (N_14068,N_9375,N_10321);
or U14069 (N_14069,N_9945,N_9817);
nand U14070 (N_14070,N_12293,N_12494);
or U14071 (N_14071,N_9443,N_11477);
and U14072 (N_14072,N_11217,N_12477);
nand U14073 (N_14073,N_9919,N_12333);
or U14074 (N_14074,N_10860,N_11832);
nor U14075 (N_14075,N_11210,N_11765);
xnor U14076 (N_14076,N_10743,N_11302);
or U14077 (N_14077,N_9876,N_10029);
nor U14078 (N_14078,N_10339,N_11596);
nand U14079 (N_14079,N_12231,N_10456);
and U14080 (N_14080,N_12324,N_11526);
or U14081 (N_14081,N_11610,N_11905);
xor U14082 (N_14082,N_11005,N_11979);
xor U14083 (N_14083,N_9754,N_11794);
nand U14084 (N_14084,N_10112,N_12375);
nand U14085 (N_14085,N_11487,N_11290);
nor U14086 (N_14086,N_9377,N_12364);
nor U14087 (N_14087,N_11508,N_10483);
nor U14088 (N_14088,N_12157,N_10251);
xnor U14089 (N_14089,N_11348,N_11850);
nand U14090 (N_14090,N_10246,N_11318);
nand U14091 (N_14091,N_9665,N_9774);
nor U14092 (N_14092,N_12169,N_9778);
and U14093 (N_14093,N_9982,N_12425);
nand U14094 (N_14094,N_11150,N_9642);
or U14095 (N_14095,N_10717,N_10681);
xnor U14096 (N_14096,N_11324,N_10841);
or U14097 (N_14097,N_10101,N_12303);
and U14098 (N_14098,N_10786,N_10167);
and U14099 (N_14099,N_9850,N_12201);
and U14100 (N_14100,N_10705,N_11971);
xor U14101 (N_14101,N_10378,N_11369);
nor U14102 (N_14102,N_11177,N_11689);
and U14103 (N_14103,N_12246,N_12374);
nor U14104 (N_14104,N_10816,N_11781);
or U14105 (N_14105,N_12091,N_12296);
and U14106 (N_14106,N_11680,N_11071);
and U14107 (N_14107,N_12076,N_9523);
and U14108 (N_14108,N_11577,N_9573);
nor U14109 (N_14109,N_11128,N_10773);
nand U14110 (N_14110,N_10533,N_9617);
and U14111 (N_14111,N_10069,N_10316);
and U14112 (N_14112,N_12058,N_11215);
or U14113 (N_14113,N_12073,N_12074);
and U14114 (N_14114,N_12135,N_12445);
nor U14115 (N_14115,N_12429,N_10609);
and U14116 (N_14116,N_11029,N_11968);
and U14117 (N_14117,N_9526,N_10148);
nor U14118 (N_14118,N_9546,N_11988);
nand U14119 (N_14119,N_11133,N_10089);
or U14120 (N_14120,N_11796,N_9657);
nand U14121 (N_14121,N_11734,N_11364);
or U14122 (N_14122,N_12125,N_9663);
or U14123 (N_14123,N_11581,N_12493);
or U14124 (N_14124,N_9686,N_10833);
nand U14125 (N_14125,N_11048,N_9488);
nand U14126 (N_14126,N_11542,N_10384);
and U14127 (N_14127,N_12288,N_10158);
nand U14128 (N_14128,N_9599,N_10045);
and U14129 (N_14129,N_11251,N_10346);
or U14130 (N_14130,N_9450,N_12011);
nor U14131 (N_14131,N_9423,N_12406);
nor U14132 (N_14132,N_10207,N_9638);
or U14133 (N_14133,N_11094,N_12101);
nor U14134 (N_14134,N_10384,N_10088);
nor U14135 (N_14135,N_10377,N_10381);
and U14136 (N_14136,N_12234,N_11520);
or U14137 (N_14137,N_10656,N_10698);
and U14138 (N_14138,N_9846,N_11104);
nand U14139 (N_14139,N_9404,N_11054);
or U14140 (N_14140,N_9884,N_11923);
nand U14141 (N_14141,N_9590,N_11746);
nand U14142 (N_14142,N_11951,N_9574);
nand U14143 (N_14143,N_9722,N_11068);
nor U14144 (N_14144,N_9477,N_10105);
or U14145 (N_14145,N_12164,N_9868);
or U14146 (N_14146,N_11306,N_11593);
nor U14147 (N_14147,N_10389,N_10868);
and U14148 (N_14148,N_9699,N_10907);
nand U14149 (N_14149,N_11400,N_10927);
or U14150 (N_14150,N_12258,N_11143);
and U14151 (N_14151,N_11069,N_10752);
nand U14152 (N_14152,N_11967,N_10967);
nor U14153 (N_14153,N_10343,N_11649);
and U14154 (N_14154,N_10594,N_11808);
nor U14155 (N_14155,N_11768,N_11185);
and U14156 (N_14156,N_10943,N_10803);
or U14157 (N_14157,N_9734,N_12227);
or U14158 (N_14158,N_10107,N_11692);
nor U14159 (N_14159,N_12103,N_10632);
and U14160 (N_14160,N_10601,N_11642);
nor U14161 (N_14161,N_11549,N_9559);
nor U14162 (N_14162,N_10347,N_10213);
nor U14163 (N_14163,N_12094,N_10851);
nand U14164 (N_14164,N_11826,N_10689);
or U14165 (N_14165,N_11789,N_10407);
nand U14166 (N_14166,N_11270,N_10486);
or U14167 (N_14167,N_10436,N_11085);
or U14168 (N_14168,N_11385,N_11051);
nand U14169 (N_14169,N_12107,N_10818);
or U14170 (N_14170,N_9951,N_11897);
nand U14171 (N_14171,N_10849,N_11776);
and U14172 (N_14172,N_11006,N_12254);
nor U14173 (N_14173,N_11030,N_9440);
or U14174 (N_14174,N_11696,N_10038);
or U14175 (N_14175,N_12078,N_9505);
or U14176 (N_14176,N_10006,N_9592);
and U14177 (N_14177,N_9466,N_9779);
nor U14178 (N_14178,N_11233,N_10649);
or U14179 (N_14179,N_9420,N_11492);
or U14180 (N_14180,N_12097,N_11783);
nor U14181 (N_14181,N_10645,N_11916);
nand U14182 (N_14182,N_9822,N_11597);
nand U14183 (N_14183,N_9534,N_10895);
or U14184 (N_14184,N_12068,N_11573);
and U14185 (N_14185,N_10098,N_11605);
xor U14186 (N_14186,N_10131,N_12153);
and U14187 (N_14187,N_10419,N_9859);
nand U14188 (N_14188,N_10290,N_12378);
nand U14189 (N_14189,N_10031,N_11158);
nor U14190 (N_14190,N_11691,N_10104);
nor U14191 (N_14191,N_10573,N_11830);
and U14192 (N_14192,N_11422,N_11193);
and U14193 (N_14193,N_11052,N_12207);
nor U14194 (N_14194,N_9504,N_11831);
and U14195 (N_14195,N_10587,N_9910);
xor U14196 (N_14196,N_12001,N_11591);
and U14197 (N_14197,N_11493,N_11918);
nor U14198 (N_14198,N_10275,N_9481);
and U14199 (N_14199,N_9732,N_12078);
and U14200 (N_14200,N_10382,N_10911);
nand U14201 (N_14201,N_11634,N_10297);
nor U14202 (N_14202,N_12377,N_9499);
or U14203 (N_14203,N_11558,N_12021);
nor U14204 (N_14204,N_12238,N_10612);
nand U14205 (N_14205,N_9558,N_10345);
nand U14206 (N_14206,N_10324,N_10991);
or U14207 (N_14207,N_11696,N_10637);
nor U14208 (N_14208,N_11015,N_9842);
nor U14209 (N_14209,N_10008,N_12302);
xnor U14210 (N_14210,N_9468,N_11976);
or U14211 (N_14211,N_10197,N_12334);
and U14212 (N_14212,N_9577,N_9627);
nor U14213 (N_14213,N_10995,N_9998);
nand U14214 (N_14214,N_11038,N_12460);
nor U14215 (N_14215,N_9806,N_11628);
xor U14216 (N_14216,N_9562,N_12047);
xnor U14217 (N_14217,N_12241,N_11451);
xnor U14218 (N_14218,N_9535,N_9740);
nor U14219 (N_14219,N_10204,N_11179);
nor U14220 (N_14220,N_11558,N_11312);
and U14221 (N_14221,N_10236,N_10992);
nor U14222 (N_14222,N_10781,N_9868);
xnor U14223 (N_14223,N_10615,N_12178);
nand U14224 (N_14224,N_11847,N_12023);
or U14225 (N_14225,N_9986,N_11172);
and U14226 (N_14226,N_11938,N_10368);
or U14227 (N_14227,N_9800,N_12378);
nor U14228 (N_14228,N_10792,N_10908);
nor U14229 (N_14229,N_11930,N_11448);
nand U14230 (N_14230,N_11755,N_10850);
nand U14231 (N_14231,N_12222,N_10323);
or U14232 (N_14232,N_11370,N_11554);
or U14233 (N_14233,N_11336,N_11275);
nand U14234 (N_14234,N_10404,N_11367);
nor U14235 (N_14235,N_10957,N_10476);
and U14236 (N_14236,N_11871,N_10455);
nand U14237 (N_14237,N_11710,N_10606);
or U14238 (N_14238,N_10837,N_11363);
or U14239 (N_14239,N_9570,N_11988);
nor U14240 (N_14240,N_12478,N_9383);
and U14241 (N_14241,N_9979,N_9808);
and U14242 (N_14242,N_11135,N_12211);
nand U14243 (N_14243,N_12021,N_12113);
or U14244 (N_14244,N_11329,N_9488);
or U14245 (N_14245,N_10427,N_12269);
or U14246 (N_14246,N_9951,N_9518);
nand U14247 (N_14247,N_10320,N_11517);
nor U14248 (N_14248,N_11322,N_9652);
and U14249 (N_14249,N_9848,N_12129);
nand U14250 (N_14250,N_9665,N_11367);
nand U14251 (N_14251,N_11678,N_12416);
and U14252 (N_14252,N_11722,N_9696);
nor U14253 (N_14253,N_11571,N_12420);
nor U14254 (N_14254,N_9803,N_12084);
nand U14255 (N_14255,N_11695,N_9749);
and U14256 (N_14256,N_11652,N_10524);
or U14257 (N_14257,N_12240,N_9592);
nor U14258 (N_14258,N_11847,N_9812);
and U14259 (N_14259,N_11881,N_9624);
nor U14260 (N_14260,N_12497,N_10527);
nand U14261 (N_14261,N_9915,N_11526);
or U14262 (N_14262,N_11966,N_11316);
nand U14263 (N_14263,N_10612,N_10115);
and U14264 (N_14264,N_9532,N_11700);
nand U14265 (N_14265,N_9623,N_12205);
xnor U14266 (N_14266,N_10443,N_12459);
and U14267 (N_14267,N_11215,N_10057);
nand U14268 (N_14268,N_10776,N_9749);
nand U14269 (N_14269,N_10600,N_11663);
nor U14270 (N_14270,N_9744,N_11919);
nor U14271 (N_14271,N_9868,N_11545);
and U14272 (N_14272,N_11921,N_10928);
or U14273 (N_14273,N_11936,N_12096);
nor U14274 (N_14274,N_9432,N_12264);
xor U14275 (N_14275,N_9992,N_12243);
nor U14276 (N_14276,N_11949,N_9749);
xnor U14277 (N_14277,N_12063,N_9781);
and U14278 (N_14278,N_10407,N_10745);
or U14279 (N_14279,N_11458,N_9609);
nor U14280 (N_14280,N_9771,N_11845);
or U14281 (N_14281,N_12181,N_10838);
and U14282 (N_14282,N_11727,N_10356);
xor U14283 (N_14283,N_10783,N_12022);
nor U14284 (N_14284,N_9376,N_12165);
or U14285 (N_14285,N_12100,N_12395);
and U14286 (N_14286,N_10809,N_12426);
and U14287 (N_14287,N_10525,N_9697);
nand U14288 (N_14288,N_9651,N_11608);
xor U14289 (N_14289,N_10792,N_9811);
and U14290 (N_14290,N_10717,N_11844);
nand U14291 (N_14291,N_12327,N_10556);
or U14292 (N_14292,N_11084,N_9866);
or U14293 (N_14293,N_11076,N_11891);
nor U14294 (N_14294,N_12185,N_9402);
nor U14295 (N_14295,N_11631,N_10962);
nor U14296 (N_14296,N_10955,N_11477);
or U14297 (N_14297,N_11179,N_10861);
xor U14298 (N_14298,N_12055,N_10243);
and U14299 (N_14299,N_12356,N_11887);
or U14300 (N_14300,N_11224,N_11416);
or U14301 (N_14301,N_11660,N_12032);
xnor U14302 (N_14302,N_10484,N_10206);
nor U14303 (N_14303,N_12479,N_12130);
xor U14304 (N_14304,N_12479,N_11426);
nand U14305 (N_14305,N_9779,N_11072);
nand U14306 (N_14306,N_11538,N_10017);
xnor U14307 (N_14307,N_12265,N_11313);
or U14308 (N_14308,N_9856,N_9866);
xnor U14309 (N_14309,N_12327,N_11917);
or U14310 (N_14310,N_11242,N_12052);
nand U14311 (N_14311,N_11128,N_11885);
or U14312 (N_14312,N_9817,N_12078);
or U14313 (N_14313,N_10414,N_12029);
or U14314 (N_14314,N_10940,N_11135);
nand U14315 (N_14315,N_11655,N_12498);
nor U14316 (N_14316,N_9914,N_9475);
nand U14317 (N_14317,N_11962,N_9727);
and U14318 (N_14318,N_9380,N_11961);
or U14319 (N_14319,N_11503,N_11471);
or U14320 (N_14320,N_9572,N_11247);
or U14321 (N_14321,N_11168,N_10001);
nand U14322 (N_14322,N_11340,N_12123);
nor U14323 (N_14323,N_10894,N_10749);
nor U14324 (N_14324,N_10173,N_12474);
or U14325 (N_14325,N_10509,N_10229);
nand U14326 (N_14326,N_11742,N_9726);
or U14327 (N_14327,N_10134,N_10348);
nor U14328 (N_14328,N_12118,N_11476);
nor U14329 (N_14329,N_12225,N_11316);
or U14330 (N_14330,N_12292,N_10859);
and U14331 (N_14331,N_11011,N_11663);
xnor U14332 (N_14332,N_10776,N_11089);
or U14333 (N_14333,N_9674,N_9939);
and U14334 (N_14334,N_9947,N_10670);
or U14335 (N_14335,N_11135,N_9495);
or U14336 (N_14336,N_9781,N_12447);
and U14337 (N_14337,N_9666,N_12072);
nor U14338 (N_14338,N_10675,N_9653);
xnor U14339 (N_14339,N_10477,N_9799);
nand U14340 (N_14340,N_9697,N_11266);
and U14341 (N_14341,N_12226,N_11742);
or U14342 (N_14342,N_12394,N_11595);
or U14343 (N_14343,N_10230,N_9769);
nor U14344 (N_14344,N_12398,N_12263);
or U14345 (N_14345,N_10928,N_11143);
and U14346 (N_14346,N_10796,N_10094);
and U14347 (N_14347,N_10986,N_11933);
or U14348 (N_14348,N_10514,N_10853);
and U14349 (N_14349,N_9412,N_11908);
or U14350 (N_14350,N_10564,N_11726);
or U14351 (N_14351,N_9939,N_9388);
and U14352 (N_14352,N_10965,N_10013);
nor U14353 (N_14353,N_11280,N_9911);
nand U14354 (N_14354,N_9989,N_11428);
or U14355 (N_14355,N_9613,N_10061);
and U14356 (N_14356,N_12471,N_11008);
and U14357 (N_14357,N_10490,N_9666);
or U14358 (N_14358,N_10806,N_12264);
nand U14359 (N_14359,N_10330,N_12359);
nand U14360 (N_14360,N_9798,N_11841);
nand U14361 (N_14361,N_10715,N_12089);
xnor U14362 (N_14362,N_11385,N_10906);
or U14363 (N_14363,N_10361,N_10930);
and U14364 (N_14364,N_10488,N_11962);
nor U14365 (N_14365,N_11040,N_10035);
nor U14366 (N_14366,N_11926,N_12092);
or U14367 (N_14367,N_11874,N_11057);
nand U14368 (N_14368,N_9897,N_9445);
and U14369 (N_14369,N_9559,N_12108);
or U14370 (N_14370,N_9422,N_9484);
nand U14371 (N_14371,N_9876,N_9989);
and U14372 (N_14372,N_10972,N_11193);
nor U14373 (N_14373,N_9981,N_12407);
and U14374 (N_14374,N_9572,N_9916);
xor U14375 (N_14375,N_10938,N_10857);
and U14376 (N_14376,N_11276,N_11407);
xnor U14377 (N_14377,N_10067,N_9417);
or U14378 (N_14378,N_9587,N_10508);
or U14379 (N_14379,N_12434,N_12355);
or U14380 (N_14380,N_11040,N_11332);
nor U14381 (N_14381,N_11104,N_11095);
xor U14382 (N_14382,N_9951,N_12038);
xor U14383 (N_14383,N_11878,N_11602);
nor U14384 (N_14384,N_9417,N_12063);
nand U14385 (N_14385,N_10175,N_10980);
and U14386 (N_14386,N_9423,N_10816);
and U14387 (N_14387,N_9924,N_11460);
nand U14388 (N_14388,N_9691,N_12478);
and U14389 (N_14389,N_12409,N_11537);
and U14390 (N_14390,N_10188,N_10915);
and U14391 (N_14391,N_10037,N_11812);
nor U14392 (N_14392,N_11715,N_12257);
xnor U14393 (N_14393,N_11757,N_10495);
nand U14394 (N_14394,N_12082,N_11421);
and U14395 (N_14395,N_9613,N_10264);
xor U14396 (N_14396,N_10782,N_10929);
nand U14397 (N_14397,N_12018,N_10565);
nor U14398 (N_14398,N_12047,N_10557);
nor U14399 (N_14399,N_9902,N_12443);
nand U14400 (N_14400,N_9494,N_11264);
and U14401 (N_14401,N_10705,N_11779);
xor U14402 (N_14402,N_11888,N_10794);
and U14403 (N_14403,N_12420,N_10158);
nor U14404 (N_14404,N_12341,N_10815);
nor U14405 (N_14405,N_12372,N_10285);
nand U14406 (N_14406,N_9837,N_12052);
and U14407 (N_14407,N_11001,N_11858);
xnor U14408 (N_14408,N_10121,N_11559);
nor U14409 (N_14409,N_9553,N_10871);
nor U14410 (N_14410,N_10704,N_10259);
xor U14411 (N_14411,N_11231,N_11270);
nand U14412 (N_14412,N_10716,N_9859);
or U14413 (N_14413,N_10851,N_10866);
or U14414 (N_14414,N_11192,N_10998);
nand U14415 (N_14415,N_10767,N_11398);
nor U14416 (N_14416,N_11714,N_9512);
nand U14417 (N_14417,N_10542,N_11050);
and U14418 (N_14418,N_12415,N_9993);
or U14419 (N_14419,N_10116,N_11059);
nand U14420 (N_14420,N_10655,N_12489);
nand U14421 (N_14421,N_12197,N_9936);
nand U14422 (N_14422,N_11889,N_10689);
or U14423 (N_14423,N_9520,N_9763);
nor U14424 (N_14424,N_11274,N_11974);
nand U14425 (N_14425,N_11966,N_9765);
and U14426 (N_14426,N_9480,N_12436);
nor U14427 (N_14427,N_10563,N_12082);
nor U14428 (N_14428,N_10964,N_11272);
nor U14429 (N_14429,N_10167,N_9415);
xor U14430 (N_14430,N_10558,N_10037);
nand U14431 (N_14431,N_9759,N_12355);
nand U14432 (N_14432,N_11952,N_9810);
or U14433 (N_14433,N_9804,N_12301);
nor U14434 (N_14434,N_12050,N_9611);
and U14435 (N_14435,N_10269,N_9417);
nand U14436 (N_14436,N_11977,N_12232);
nor U14437 (N_14437,N_9426,N_10983);
and U14438 (N_14438,N_11137,N_11364);
nor U14439 (N_14439,N_11211,N_11464);
or U14440 (N_14440,N_11578,N_10755);
nor U14441 (N_14441,N_10736,N_11740);
nor U14442 (N_14442,N_11980,N_11214);
or U14443 (N_14443,N_9476,N_11452);
or U14444 (N_14444,N_9621,N_11744);
nor U14445 (N_14445,N_11768,N_10198);
or U14446 (N_14446,N_10526,N_10449);
or U14447 (N_14447,N_11650,N_10184);
nand U14448 (N_14448,N_9849,N_12251);
nor U14449 (N_14449,N_9565,N_10105);
nand U14450 (N_14450,N_10926,N_10420);
or U14451 (N_14451,N_12049,N_10211);
or U14452 (N_14452,N_11842,N_10483);
nor U14453 (N_14453,N_11417,N_10289);
nand U14454 (N_14454,N_11830,N_11285);
nor U14455 (N_14455,N_11807,N_11833);
or U14456 (N_14456,N_11186,N_9645);
nor U14457 (N_14457,N_9494,N_10138);
or U14458 (N_14458,N_12205,N_9680);
or U14459 (N_14459,N_10519,N_10159);
or U14460 (N_14460,N_12165,N_10804);
or U14461 (N_14461,N_9919,N_10939);
and U14462 (N_14462,N_9981,N_11657);
or U14463 (N_14463,N_10402,N_10726);
nor U14464 (N_14464,N_12320,N_12310);
nand U14465 (N_14465,N_11964,N_9801);
nor U14466 (N_14466,N_11026,N_11260);
nor U14467 (N_14467,N_10886,N_11383);
nor U14468 (N_14468,N_9998,N_10197);
nor U14469 (N_14469,N_12390,N_12241);
nor U14470 (N_14470,N_10221,N_11464);
or U14471 (N_14471,N_9670,N_11466);
or U14472 (N_14472,N_12443,N_11121);
nor U14473 (N_14473,N_9913,N_10002);
nand U14474 (N_14474,N_10310,N_9878);
and U14475 (N_14475,N_10173,N_9585);
xnor U14476 (N_14476,N_11806,N_12178);
or U14477 (N_14477,N_10723,N_10330);
and U14478 (N_14478,N_11530,N_9973);
or U14479 (N_14479,N_10567,N_11594);
nor U14480 (N_14480,N_9670,N_12186);
nand U14481 (N_14481,N_11252,N_10587);
and U14482 (N_14482,N_12285,N_10840);
nor U14483 (N_14483,N_11325,N_9855);
and U14484 (N_14484,N_11128,N_12069);
nand U14485 (N_14485,N_10098,N_11771);
and U14486 (N_14486,N_11489,N_11240);
nor U14487 (N_14487,N_11171,N_12301);
and U14488 (N_14488,N_11762,N_10024);
nand U14489 (N_14489,N_10678,N_12402);
or U14490 (N_14490,N_11150,N_9633);
and U14491 (N_14491,N_12473,N_11458);
and U14492 (N_14492,N_12446,N_10373);
nand U14493 (N_14493,N_11019,N_9688);
xnor U14494 (N_14494,N_12158,N_11074);
nor U14495 (N_14495,N_10504,N_10521);
and U14496 (N_14496,N_10160,N_10333);
and U14497 (N_14497,N_10515,N_11153);
or U14498 (N_14498,N_10919,N_12013);
or U14499 (N_14499,N_10517,N_10867);
or U14500 (N_14500,N_10265,N_9873);
and U14501 (N_14501,N_9793,N_10450);
nand U14502 (N_14502,N_10515,N_10922);
nor U14503 (N_14503,N_12335,N_11043);
and U14504 (N_14504,N_9807,N_10782);
xnor U14505 (N_14505,N_12078,N_10212);
nor U14506 (N_14506,N_11626,N_10248);
or U14507 (N_14507,N_9813,N_11453);
nand U14508 (N_14508,N_12154,N_11644);
and U14509 (N_14509,N_9520,N_11027);
and U14510 (N_14510,N_11234,N_9725);
and U14511 (N_14511,N_10128,N_9548);
or U14512 (N_14512,N_10030,N_11725);
nand U14513 (N_14513,N_12294,N_12263);
nor U14514 (N_14514,N_9404,N_10495);
or U14515 (N_14515,N_12251,N_11475);
xor U14516 (N_14516,N_11949,N_12496);
and U14517 (N_14517,N_11419,N_10274);
or U14518 (N_14518,N_11076,N_11991);
nor U14519 (N_14519,N_12356,N_11271);
or U14520 (N_14520,N_10287,N_10687);
nand U14521 (N_14521,N_9869,N_12265);
or U14522 (N_14522,N_9386,N_10273);
or U14523 (N_14523,N_11701,N_11736);
nor U14524 (N_14524,N_9529,N_11278);
nor U14525 (N_14525,N_11114,N_12161);
and U14526 (N_14526,N_10907,N_9981);
and U14527 (N_14527,N_10930,N_10210);
or U14528 (N_14528,N_11220,N_12031);
nand U14529 (N_14529,N_12199,N_12305);
nand U14530 (N_14530,N_10946,N_10271);
and U14531 (N_14531,N_9464,N_10135);
nor U14532 (N_14532,N_11137,N_9679);
xor U14533 (N_14533,N_12062,N_11454);
nor U14534 (N_14534,N_12404,N_10256);
or U14535 (N_14535,N_11878,N_10866);
nor U14536 (N_14536,N_11517,N_11286);
nand U14537 (N_14537,N_11585,N_12478);
or U14538 (N_14538,N_11440,N_11558);
or U14539 (N_14539,N_10472,N_10795);
nand U14540 (N_14540,N_9502,N_11101);
or U14541 (N_14541,N_9471,N_10372);
nor U14542 (N_14542,N_10494,N_9818);
and U14543 (N_14543,N_10627,N_9602);
or U14544 (N_14544,N_12498,N_10565);
or U14545 (N_14545,N_9882,N_10977);
or U14546 (N_14546,N_10198,N_10121);
nor U14547 (N_14547,N_12209,N_10882);
nor U14548 (N_14548,N_12009,N_11969);
nor U14549 (N_14549,N_11569,N_10067);
or U14550 (N_14550,N_9535,N_9935);
nand U14551 (N_14551,N_12242,N_9545);
xor U14552 (N_14552,N_10719,N_11991);
xor U14553 (N_14553,N_11175,N_10074);
and U14554 (N_14554,N_9721,N_11464);
nor U14555 (N_14555,N_12369,N_10382);
nand U14556 (N_14556,N_9962,N_9740);
and U14557 (N_14557,N_11154,N_10452);
nor U14558 (N_14558,N_10291,N_11012);
nand U14559 (N_14559,N_11913,N_9833);
nand U14560 (N_14560,N_12183,N_12318);
or U14561 (N_14561,N_11645,N_12378);
xor U14562 (N_14562,N_11524,N_12064);
nand U14563 (N_14563,N_12196,N_12377);
nand U14564 (N_14564,N_10273,N_11750);
nor U14565 (N_14565,N_11753,N_9973);
or U14566 (N_14566,N_10835,N_11146);
nand U14567 (N_14567,N_11673,N_11701);
nor U14568 (N_14568,N_11120,N_12348);
xnor U14569 (N_14569,N_12486,N_9599);
xor U14570 (N_14570,N_9900,N_10716);
nand U14571 (N_14571,N_11824,N_10985);
and U14572 (N_14572,N_9747,N_10515);
nor U14573 (N_14573,N_9699,N_11590);
nand U14574 (N_14574,N_12188,N_11782);
nand U14575 (N_14575,N_10011,N_11747);
xnor U14576 (N_14576,N_9832,N_11154);
nor U14577 (N_14577,N_12438,N_11347);
or U14578 (N_14578,N_11677,N_11823);
and U14579 (N_14579,N_9770,N_12140);
or U14580 (N_14580,N_9932,N_11146);
or U14581 (N_14581,N_10739,N_12489);
or U14582 (N_14582,N_11195,N_12461);
or U14583 (N_14583,N_10784,N_11880);
nor U14584 (N_14584,N_10822,N_11370);
nor U14585 (N_14585,N_11098,N_9771);
nor U14586 (N_14586,N_11073,N_11745);
xor U14587 (N_14587,N_10701,N_10505);
nor U14588 (N_14588,N_10568,N_10597);
xnor U14589 (N_14589,N_10304,N_10076);
nor U14590 (N_14590,N_10084,N_9452);
nand U14591 (N_14591,N_11151,N_12417);
or U14592 (N_14592,N_10564,N_10959);
nor U14593 (N_14593,N_11692,N_11584);
nor U14594 (N_14594,N_10342,N_11257);
nor U14595 (N_14595,N_9778,N_10279);
and U14596 (N_14596,N_10998,N_12451);
or U14597 (N_14597,N_10285,N_11712);
nand U14598 (N_14598,N_10811,N_9924);
nand U14599 (N_14599,N_11528,N_10574);
nor U14600 (N_14600,N_9836,N_11633);
nand U14601 (N_14601,N_11364,N_9452);
and U14602 (N_14602,N_10028,N_10098);
nand U14603 (N_14603,N_10591,N_9405);
or U14604 (N_14604,N_12000,N_10333);
nand U14605 (N_14605,N_11587,N_9629);
nand U14606 (N_14606,N_9859,N_11829);
or U14607 (N_14607,N_10829,N_9382);
or U14608 (N_14608,N_12477,N_11713);
xnor U14609 (N_14609,N_11564,N_12364);
xor U14610 (N_14610,N_9464,N_11373);
nor U14611 (N_14611,N_12446,N_12486);
xnor U14612 (N_14612,N_12364,N_10384);
nor U14613 (N_14613,N_10054,N_10838);
nor U14614 (N_14614,N_10244,N_9912);
nand U14615 (N_14615,N_12154,N_11148);
nand U14616 (N_14616,N_10309,N_11950);
nand U14617 (N_14617,N_11580,N_12095);
and U14618 (N_14618,N_10426,N_12472);
and U14619 (N_14619,N_11080,N_11597);
nand U14620 (N_14620,N_11366,N_12293);
nand U14621 (N_14621,N_10263,N_11278);
xor U14622 (N_14622,N_11864,N_11135);
and U14623 (N_14623,N_10866,N_9835);
nor U14624 (N_14624,N_9467,N_10370);
xnor U14625 (N_14625,N_12453,N_9470);
nor U14626 (N_14626,N_10675,N_12369);
nor U14627 (N_14627,N_11982,N_12157);
or U14628 (N_14628,N_12436,N_11110);
nor U14629 (N_14629,N_11574,N_12251);
nand U14630 (N_14630,N_11286,N_9749);
nand U14631 (N_14631,N_10002,N_10980);
or U14632 (N_14632,N_11207,N_10789);
xnor U14633 (N_14633,N_11917,N_9390);
or U14634 (N_14634,N_10480,N_11205);
nor U14635 (N_14635,N_9993,N_10325);
nand U14636 (N_14636,N_12350,N_10940);
xor U14637 (N_14637,N_9916,N_9995);
and U14638 (N_14638,N_11481,N_11161);
or U14639 (N_14639,N_11384,N_12396);
nor U14640 (N_14640,N_9915,N_11514);
and U14641 (N_14641,N_10468,N_12178);
and U14642 (N_14642,N_9954,N_10990);
and U14643 (N_14643,N_11069,N_11345);
or U14644 (N_14644,N_9515,N_10329);
or U14645 (N_14645,N_11916,N_9514);
nor U14646 (N_14646,N_10978,N_9902);
nor U14647 (N_14647,N_11356,N_11351);
or U14648 (N_14648,N_9431,N_9622);
or U14649 (N_14649,N_10780,N_11596);
and U14650 (N_14650,N_12378,N_10293);
and U14651 (N_14651,N_11856,N_11298);
and U14652 (N_14652,N_10574,N_11289);
xnor U14653 (N_14653,N_9382,N_10372);
nor U14654 (N_14654,N_12287,N_11489);
nand U14655 (N_14655,N_11955,N_9479);
nor U14656 (N_14656,N_10672,N_11855);
nor U14657 (N_14657,N_11898,N_11370);
nor U14658 (N_14658,N_9823,N_11222);
nor U14659 (N_14659,N_11176,N_11411);
and U14660 (N_14660,N_10241,N_9695);
nand U14661 (N_14661,N_12217,N_11177);
or U14662 (N_14662,N_10843,N_11456);
and U14663 (N_14663,N_10884,N_9643);
nor U14664 (N_14664,N_9684,N_12450);
and U14665 (N_14665,N_10525,N_11946);
nor U14666 (N_14666,N_12199,N_10697);
and U14667 (N_14667,N_9566,N_10146);
nand U14668 (N_14668,N_10424,N_9818);
nor U14669 (N_14669,N_11820,N_10916);
and U14670 (N_14670,N_11379,N_10541);
xnor U14671 (N_14671,N_11745,N_9682);
and U14672 (N_14672,N_10657,N_10817);
or U14673 (N_14673,N_9604,N_11390);
nor U14674 (N_14674,N_10225,N_10431);
or U14675 (N_14675,N_11346,N_9727);
nand U14676 (N_14676,N_11636,N_10686);
nor U14677 (N_14677,N_9929,N_12105);
or U14678 (N_14678,N_10315,N_9406);
and U14679 (N_14679,N_12385,N_11657);
nor U14680 (N_14680,N_9949,N_10890);
nand U14681 (N_14681,N_9610,N_9993);
or U14682 (N_14682,N_10591,N_11613);
or U14683 (N_14683,N_11856,N_11031);
nand U14684 (N_14684,N_11733,N_9924);
nor U14685 (N_14685,N_11870,N_10058);
or U14686 (N_14686,N_9521,N_10376);
nand U14687 (N_14687,N_9605,N_11631);
nor U14688 (N_14688,N_12177,N_11201);
and U14689 (N_14689,N_9915,N_11908);
or U14690 (N_14690,N_9555,N_10186);
nor U14691 (N_14691,N_11969,N_11300);
or U14692 (N_14692,N_10902,N_10085);
nand U14693 (N_14693,N_10710,N_9419);
nor U14694 (N_14694,N_11405,N_10229);
or U14695 (N_14695,N_11660,N_9940);
and U14696 (N_14696,N_12220,N_11591);
nor U14697 (N_14697,N_10515,N_12015);
xnor U14698 (N_14698,N_12434,N_11013);
nand U14699 (N_14699,N_9528,N_11485);
nor U14700 (N_14700,N_11227,N_11926);
and U14701 (N_14701,N_10862,N_9442);
nand U14702 (N_14702,N_9985,N_11642);
xor U14703 (N_14703,N_10921,N_9507);
nand U14704 (N_14704,N_9722,N_10783);
nor U14705 (N_14705,N_12025,N_10775);
or U14706 (N_14706,N_11358,N_9493);
and U14707 (N_14707,N_9786,N_10711);
nor U14708 (N_14708,N_10197,N_9878);
nand U14709 (N_14709,N_12051,N_12231);
and U14710 (N_14710,N_10389,N_10624);
nand U14711 (N_14711,N_9492,N_10649);
nand U14712 (N_14712,N_12291,N_12303);
nor U14713 (N_14713,N_10440,N_11000);
or U14714 (N_14714,N_12322,N_11101);
and U14715 (N_14715,N_11350,N_10057);
xor U14716 (N_14716,N_11136,N_9406);
xor U14717 (N_14717,N_9379,N_12211);
xnor U14718 (N_14718,N_11382,N_10376);
nor U14719 (N_14719,N_10438,N_9401);
or U14720 (N_14720,N_12429,N_11068);
xor U14721 (N_14721,N_11353,N_9614);
and U14722 (N_14722,N_11472,N_9484);
or U14723 (N_14723,N_9948,N_11760);
xnor U14724 (N_14724,N_9882,N_10948);
and U14725 (N_14725,N_10459,N_11016);
or U14726 (N_14726,N_9784,N_11077);
nor U14727 (N_14727,N_9650,N_10472);
nor U14728 (N_14728,N_11257,N_11658);
and U14729 (N_14729,N_10634,N_11630);
nand U14730 (N_14730,N_10182,N_12045);
and U14731 (N_14731,N_11871,N_12371);
or U14732 (N_14732,N_10019,N_9673);
nor U14733 (N_14733,N_11916,N_9402);
and U14734 (N_14734,N_9997,N_12100);
nand U14735 (N_14735,N_11714,N_12282);
nand U14736 (N_14736,N_10644,N_11086);
nor U14737 (N_14737,N_12417,N_12328);
or U14738 (N_14738,N_9403,N_10013);
or U14739 (N_14739,N_12236,N_11541);
nor U14740 (N_14740,N_9428,N_10235);
and U14741 (N_14741,N_10119,N_10411);
or U14742 (N_14742,N_11315,N_10796);
nand U14743 (N_14743,N_10747,N_11603);
or U14744 (N_14744,N_10095,N_12087);
xnor U14745 (N_14745,N_9583,N_12132);
nor U14746 (N_14746,N_11354,N_10323);
and U14747 (N_14747,N_11349,N_11264);
nand U14748 (N_14748,N_10324,N_10343);
xnor U14749 (N_14749,N_10895,N_11633);
or U14750 (N_14750,N_10792,N_11366);
nor U14751 (N_14751,N_11512,N_11002);
or U14752 (N_14752,N_9577,N_11098);
or U14753 (N_14753,N_11389,N_11590);
nor U14754 (N_14754,N_9527,N_12306);
nand U14755 (N_14755,N_10887,N_9661);
and U14756 (N_14756,N_9920,N_11304);
nor U14757 (N_14757,N_11786,N_12222);
nand U14758 (N_14758,N_9650,N_12388);
nand U14759 (N_14759,N_11338,N_11546);
and U14760 (N_14760,N_11278,N_12399);
and U14761 (N_14761,N_11562,N_12435);
nand U14762 (N_14762,N_11288,N_12235);
xor U14763 (N_14763,N_9985,N_9711);
nand U14764 (N_14764,N_11666,N_11205);
or U14765 (N_14765,N_11541,N_11057);
or U14766 (N_14766,N_10456,N_9872);
nor U14767 (N_14767,N_10189,N_12253);
or U14768 (N_14768,N_9974,N_10002);
and U14769 (N_14769,N_11551,N_9955);
or U14770 (N_14770,N_9901,N_10009);
nand U14771 (N_14771,N_9868,N_10491);
or U14772 (N_14772,N_11681,N_9618);
xor U14773 (N_14773,N_12179,N_9445);
or U14774 (N_14774,N_12056,N_12295);
nand U14775 (N_14775,N_9874,N_9946);
and U14776 (N_14776,N_10509,N_11429);
xor U14777 (N_14777,N_12193,N_10135);
nand U14778 (N_14778,N_10763,N_11410);
nor U14779 (N_14779,N_10292,N_12422);
or U14780 (N_14780,N_11733,N_10818);
nand U14781 (N_14781,N_10698,N_9458);
and U14782 (N_14782,N_9899,N_11375);
and U14783 (N_14783,N_11500,N_12215);
and U14784 (N_14784,N_11709,N_10907);
nand U14785 (N_14785,N_11848,N_11831);
xnor U14786 (N_14786,N_12342,N_9558);
and U14787 (N_14787,N_11596,N_12253);
xor U14788 (N_14788,N_10566,N_10738);
or U14789 (N_14789,N_11664,N_11626);
and U14790 (N_14790,N_11855,N_12345);
and U14791 (N_14791,N_11586,N_10439);
nor U14792 (N_14792,N_12481,N_12248);
xnor U14793 (N_14793,N_10051,N_9555);
nor U14794 (N_14794,N_11283,N_9462);
or U14795 (N_14795,N_12448,N_10490);
nand U14796 (N_14796,N_10860,N_10592);
nand U14797 (N_14797,N_9476,N_10294);
nor U14798 (N_14798,N_9889,N_9767);
nand U14799 (N_14799,N_11337,N_11692);
nand U14800 (N_14800,N_10038,N_11033);
and U14801 (N_14801,N_12037,N_10926);
nand U14802 (N_14802,N_9847,N_11712);
and U14803 (N_14803,N_12272,N_11597);
or U14804 (N_14804,N_12220,N_11005);
nor U14805 (N_14805,N_12466,N_9996);
nand U14806 (N_14806,N_10488,N_12419);
nand U14807 (N_14807,N_10548,N_11074);
and U14808 (N_14808,N_10497,N_11177);
and U14809 (N_14809,N_9975,N_12222);
nand U14810 (N_14810,N_10136,N_12290);
and U14811 (N_14811,N_9766,N_11596);
and U14812 (N_14812,N_10963,N_10365);
and U14813 (N_14813,N_12047,N_9407);
nand U14814 (N_14814,N_12371,N_9897);
and U14815 (N_14815,N_9659,N_11294);
nor U14816 (N_14816,N_10100,N_9750);
nand U14817 (N_14817,N_11068,N_12421);
nor U14818 (N_14818,N_11787,N_10168);
nor U14819 (N_14819,N_10060,N_9383);
and U14820 (N_14820,N_9737,N_9456);
nand U14821 (N_14821,N_10558,N_10355);
and U14822 (N_14822,N_12074,N_11151);
and U14823 (N_14823,N_12423,N_10127);
nor U14824 (N_14824,N_9558,N_11764);
nor U14825 (N_14825,N_11517,N_9749);
nor U14826 (N_14826,N_12341,N_11361);
nor U14827 (N_14827,N_10956,N_12099);
nand U14828 (N_14828,N_9413,N_12481);
or U14829 (N_14829,N_12238,N_10915);
or U14830 (N_14830,N_9772,N_12092);
nand U14831 (N_14831,N_10070,N_10429);
nand U14832 (N_14832,N_10104,N_12423);
or U14833 (N_14833,N_12423,N_10656);
and U14834 (N_14834,N_12019,N_11851);
nor U14835 (N_14835,N_9416,N_9629);
and U14836 (N_14836,N_11124,N_11432);
and U14837 (N_14837,N_10666,N_11708);
nand U14838 (N_14838,N_11392,N_9482);
or U14839 (N_14839,N_10009,N_10269);
nor U14840 (N_14840,N_12448,N_9851);
and U14841 (N_14841,N_12430,N_11592);
and U14842 (N_14842,N_11288,N_9777);
nand U14843 (N_14843,N_9476,N_12302);
or U14844 (N_14844,N_11003,N_10584);
and U14845 (N_14845,N_10309,N_9969);
or U14846 (N_14846,N_10324,N_12162);
nor U14847 (N_14847,N_11231,N_10940);
or U14848 (N_14848,N_9827,N_12113);
or U14849 (N_14849,N_10588,N_11452);
xnor U14850 (N_14850,N_10128,N_12358);
xnor U14851 (N_14851,N_12161,N_9385);
nand U14852 (N_14852,N_10058,N_9395);
and U14853 (N_14853,N_11502,N_11728);
and U14854 (N_14854,N_11790,N_9523);
or U14855 (N_14855,N_10076,N_10501);
nand U14856 (N_14856,N_10419,N_12463);
and U14857 (N_14857,N_11602,N_11362);
or U14858 (N_14858,N_10400,N_10253);
nand U14859 (N_14859,N_12005,N_10049);
and U14860 (N_14860,N_12353,N_11616);
nor U14861 (N_14861,N_10304,N_9891);
nand U14862 (N_14862,N_12374,N_12104);
nor U14863 (N_14863,N_9921,N_10446);
xnor U14864 (N_14864,N_10614,N_10848);
and U14865 (N_14865,N_11861,N_10470);
xnor U14866 (N_14866,N_10578,N_11121);
and U14867 (N_14867,N_10731,N_11689);
or U14868 (N_14868,N_9390,N_12138);
xor U14869 (N_14869,N_10184,N_10522);
nand U14870 (N_14870,N_10269,N_11318);
or U14871 (N_14871,N_9572,N_10240);
nor U14872 (N_14872,N_9829,N_9390);
nand U14873 (N_14873,N_12245,N_10374);
nor U14874 (N_14874,N_11920,N_10483);
nand U14875 (N_14875,N_12006,N_10685);
nor U14876 (N_14876,N_11018,N_10664);
and U14877 (N_14877,N_11906,N_9552);
and U14878 (N_14878,N_12284,N_9860);
xnor U14879 (N_14879,N_10017,N_11937);
or U14880 (N_14880,N_11027,N_11124);
or U14881 (N_14881,N_11345,N_10970);
nand U14882 (N_14882,N_9560,N_11710);
and U14883 (N_14883,N_10375,N_10108);
xor U14884 (N_14884,N_12472,N_11611);
or U14885 (N_14885,N_10724,N_11176);
and U14886 (N_14886,N_12437,N_10906);
or U14887 (N_14887,N_11592,N_10100);
or U14888 (N_14888,N_12283,N_10641);
or U14889 (N_14889,N_12027,N_11882);
or U14890 (N_14890,N_10806,N_10910);
nor U14891 (N_14891,N_10649,N_12458);
xnor U14892 (N_14892,N_11230,N_9790);
nor U14893 (N_14893,N_9582,N_10417);
nor U14894 (N_14894,N_11255,N_12429);
nor U14895 (N_14895,N_11440,N_10522);
nand U14896 (N_14896,N_12470,N_11651);
nor U14897 (N_14897,N_10244,N_12114);
xnor U14898 (N_14898,N_12148,N_10269);
or U14899 (N_14899,N_10426,N_12493);
xor U14900 (N_14900,N_10971,N_11857);
nand U14901 (N_14901,N_9504,N_9386);
nor U14902 (N_14902,N_11204,N_9559);
nor U14903 (N_14903,N_10639,N_9933);
nand U14904 (N_14904,N_9964,N_12244);
or U14905 (N_14905,N_10663,N_11923);
or U14906 (N_14906,N_10093,N_10881);
nand U14907 (N_14907,N_10375,N_9607);
xnor U14908 (N_14908,N_10233,N_11711);
and U14909 (N_14909,N_10308,N_11295);
nand U14910 (N_14910,N_10970,N_9952);
nand U14911 (N_14911,N_9950,N_11788);
nand U14912 (N_14912,N_10074,N_9549);
or U14913 (N_14913,N_12472,N_11545);
or U14914 (N_14914,N_11887,N_9945);
nor U14915 (N_14915,N_10201,N_9670);
nor U14916 (N_14916,N_11042,N_10128);
or U14917 (N_14917,N_11055,N_11398);
nor U14918 (N_14918,N_10682,N_9967);
and U14919 (N_14919,N_10185,N_12305);
nand U14920 (N_14920,N_11820,N_10650);
and U14921 (N_14921,N_10580,N_9840);
nor U14922 (N_14922,N_9574,N_10338);
nor U14923 (N_14923,N_11068,N_9761);
xor U14924 (N_14924,N_10536,N_10508);
nand U14925 (N_14925,N_11069,N_10756);
nand U14926 (N_14926,N_10543,N_10575);
nor U14927 (N_14927,N_9446,N_12374);
and U14928 (N_14928,N_12176,N_10760);
nor U14929 (N_14929,N_10936,N_9548);
nor U14930 (N_14930,N_11386,N_10184);
or U14931 (N_14931,N_9646,N_10460);
xor U14932 (N_14932,N_12190,N_10527);
or U14933 (N_14933,N_9820,N_10500);
or U14934 (N_14934,N_10815,N_11019);
nand U14935 (N_14935,N_10818,N_9746);
xnor U14936 (N_14936,N_9764,N_10011);
nor U14937 (N_14937,N_12153,N_11612);
or U14938 (N_14938,N_10113,N_12239);
and U14939 (N_14939,N_10420,N_12238);
nor U14940 (N_14940,N_10121,N_10666);
and U14941 (N_14941,N_11389,N_12313);
nor U14942 (N_14942,N_10959,N_9882);
and U14943 (N_14943,N_11053,N_10520);
nor U14944 (N_14944,N_9989,N_10986);
or U14945 (N_14945,N_10539,N_12489);
nand U14946 (N_14946,N_11440,N_11444);
nand U14947 (N_14947,N_9767,N_10600);
xnor U14948 (N_14948,N_10488,N_9697);
nand U14949 (N_14949,N_11990,N_11404);
nand U14950 (N_14950,N_12041,N_9442);
xnor U14951 (N_14951,N_9757,N_10776);
nand U14952 (N_14952,N_9687,N_11302);
and U14953 (N_14953,N_10102,N_12368);
or U14954 (N_14954,N_11890,N_9910);
and U14955 (N_14955,N_11437,N_10432);
and U14956 (N_14956,N_10361,N_11615);
xor U14957 (N_14957,N_10779,N_11554);
nand U14958 (N_14958,N_10078,N_10111);
nand U14959 (N_14959,N_9587,N_9796);
nor U14960 (N_14960,N_11626,N_10149);
or U14961 (N_14961,N_11669,N_10590);
or U14962 (N_14962,N_10874,N_12143);
or U14963 (N_14963,N_10858,N_11101);
nand U14964 (N_14964,N_10480,N_11626);
or U14965 (N_14965,N_9911,N_10304);
xor U14966 (N_14966,N_11669,N_10824);
or U14967 (N_14967,N_11581,N_9720);
and U14968 (N_14968,N_10363,N_10045);
nor U14969 (N_14969,N_12318,N_11191);
or U14970 (N_14970,N_9455,N_11398);
and U14971 (N_14971,N_10125,N_11107);
xor U14972 (N_14972,N_11423,N_12190);
xor U14973 (N_14973,N_9944,N_9994);
or U14974 (N_14974,N_11306,N_11094);
and U14975 (N_14975,N_11897,N_9682);
nand U14976 (N_14976,N_11003,N_11684);
or U14977 (N_14977,N_12384,N_12428);
and U14978 (N_14978,N_10572,N_10019);
and U14979 (N_14979,N_11170,N_9905);
or U14980 (N_14980,N_11260,N_10007);
or U14981 (N_14981,N_12479,N_10480);
nor U14982 (N_14982,N_11226,N_9963);
nor U14983 (N_14983,N_11487,N_10962);
and U14984 (N_14984,N_9408,N_10859);
nor U14985 (N_14985,N_11364,N_10287);
nand U14986 (N_14986,N_12149,N_9533);
nand U14987 (N_14987,N_9911,N_11369);
or U14988 (N_14988,N_11354,N_12448);
nor U14989 (N_14989,N_12111,N_10650);
nor U14990 (N_14990,N_10814,N_10562);
or U14991 (N_14991,N_12342,N_10542);
or U14992 (N_14992,N_10562,N_11848);
and U14993 (N_14993,N_9391,N_12179);
and U14994 (N_14994,N_11314,N_11300);
and U14995 (N_14995,N_9600,N_12371);
nor U14996 (N_14996,N_11068,N_10905);
or U14997 (N_14997,N_12153,N_12178);
and U14998 (N_14998,N_9558,N_11496);
xnor U14999 (N_14999,N_10068,N_12308);
nand U15000 (N_15000,N_9456,N_11375);
or U15001 (N_15001,N_9794,N_10384);
or U15002 (N_15002,N_12284,N_11405);
nor U15003 (N_15003,N_10622,N_12322);
and U15004 (N_15004,N_10777,N_11787);
or U15005 (N_15005,N_12102,N_9550);
or U15006 (N_15006,N_11353,N_11671);
and U15007 (N_15007,N_10466,N_9898);
and U15008 (N_15008,N_10882,N_10911);
nor U15009 (N_15009,N_10962,N_11231);
and U15010 (N_15010,N_10757,N_11590);
or U15011 (N_15011,N_9655,N_12273);
nand U15012 (N_15012,N_10355,N_11555);
nor U15013 (N_15013,N_12372,N_11067);
or U15014 (N_15014,N_11927,N_12359);
and U15015 (N_15015,N_11071,N_12111);
nor U15016 (N_15016,N_11743,N_12322);
or U15017 (N_15017,N_10188,N_10292);
or U15018 (N_15018,N_11775,N_9432);
nand U15019 (N_15019,N_10551,N_9397);
nor U15020 (N_15020,N_12419,N_12183);
nand U15021 (N_15021,N_10191,N_11022);
nor U15022 (N_15022,N_10662,N_11586);
and U15023 (N_15023,N_9972,N_10083);
nor U15024 (N_15024,N_9991,N_11588);
nor U15025 (N_15025,N_11502,N_10771);
nand U15026 (N_15026,N_11680,N_9496);
nor U15027 (N_15027,N_9641,N_9496);
nor U15028 (N_15028,N_11193,N_12182);
nand U15029 (N_15029,N_12022,N_11533);
nor U15030 (N_15030,N_10243,N_10467);
nand U15031 (N_15031,N_10679,N_10064);
or U15032 (N_15032,N_10561,N_9500);
and U15033 (N_15033,N_9689,N_10152);
nand U15034 (N_15034,N_10818,N_12322);
or U15035 (N_15035,N_10583,N_10779);
nor U15036 (N_15036,N_9491,N_10697);
nand U15037 (N_15037,N_9389,N_9427);
nor U15038 (N_15038,N_9765,N_9657);
xnor U15039 (N_15039,N_9375,N_11402);
nor U15040 (N_15040,N_12097,N_9816);
xor U15041 (N_15041,N_10148,N_10834);
xor U15042 (N_15042,N_9921,N_10264);
nand U15043 (N_15043,N_10285,N_12452);
nand U15044 (N_15044,N_9407,N_10865);
nor U15045 (N_15045,N_11850,N_10635);
and U15046 (N_15046,N_10851,N_9656);
or U15047 (N_15047,N_10683,N_11118);
and U15048 (N_15048,N_12074,N_10627);
nand U15049 (N_15049,N_10229,N_12092);
nand U15050 (N_15050,N_10668,N_9941);
nand U15051 (N_15051,N_10203,N_10260);
or U15052 (N_15052,N_10187,N_10556);
or U15053 (N_15053,N_11622,N_9626);
nand U15054 (N_15054,N_10462,N_10225);
or U15055 (N_15055,N_10136,N_11119);
nand U15056 (N_15056,N_9451,N_12384);
and U15057 (N_15057,N_11521,N_11572);
xor U15058 (N_15058,N_10926,N_9386);
and U15059 (N_15059,N_9806,N_9735);
xnor U15060 (N_15060,N_12440,N_12405);
nor U15061 (N_15061,N_12465,N_10756);
nor U15062 (N_15062,N_10440,N_9950);
xnor U15063 (N_15063,N_9551,N_9449);
and U15064 (N_15064,N_12049,N_10153);
and U15065 (N_15065,N_11263,N_10734);
nor U15066 (N_15066,N_10287,N_11602);
or U15067 (N_15067,N_9637,N_9724);
nor U15068 (N_15068,N_10079,N_11519);
nor U15069 (N_15069,N_11392,N_10690);
nor U15070 (N_15070,N_9573,N_11982);
or U15071 (N_15071,N_9637,N_11520);
nand U15072 (N_15072,N_10949,N_12381);
nand U15073 (N_15073,N_12210,N_11458);
nor U15074 (N_15074,N_11209,N_10949);
or U15075 (N_15075,N_9931,N_11603);
nor U15076 (N_15076,N_11231,N_9975);
nor U15077 (N_15077,N_11677,N_11466);
nor U15078 (N_15078,N_10121,N_10298);
nor U15079 (N_15079,N_9534,N_10129);
xor U15080 (N_15080,N_10090,N_10166);
nor U15081 (N_15081,N_11017,N_9882);
or U15082 (N_15082,N_10412,N_11203);
or U15083 (N_15083,N_10076,N_10328);
and U15084 (N_15084,N_9604,N_10829);
nor U15085 (N_15085,N_10625,N_11010);
and U15086 (N_15086,N_11263,N_11514);
and U15087 (N_15087,N_11838,N_11840);
or U15088 (N_15088,N_10364,N_10171);
xnor U15089 (N_15089,N_10277,N_9977);
or U15090 (N_15090,N_12110,N_10358);
or U15091 (N_15091,N_9532,N_10030);
nand U15092 (N_15092,N_9694,N_10268);
nor U15093 (N_15093,N_11064,N_12118);
or U15094 (N_15094,N_9765,N_10475);
nor U15095 (N_15095,N_11092,N_10298);
nand U15096 (N_15096,N_9490,N_12240);
nor U15097 (N_15097,N_9788,N_9860);
nand U15098 (N_15098,N_9777,N_12332);
nand U15099 (N_15099,N_9452,N_9903);
nand U15100 (N_15100,N_9562,N_11708);
and U15101 (N_15101,N_12064,N_10700);
nand U15102 (N_15102,N_10808,N_12474);
nand U15103 (N_15103,N_10800,N_12205);
nor U15104 (N_15104,N_12236,N_10916);
or U15105 (N_15105,N_9620,N_10707);
and U15106 (N_15106,N_10431,N_11875);
xor U15107 (N_15107,N_10979,N_11325);
and U15108 (N_15108,N_11035,N_11765);
xnor U15109 (N_15109,N_12193,N_11237);
and U15110 (N_15110,N_9760,N_10679);
or U15111 (N_15111,N_10548,N_9460);
nand U15112 (N_15112,N_10621,N_12085);
nor U15113 (N_15113,N_11778,N_9391);
and U15114 (N_15114,N_12279,N_11779);
or U15115 (N_15115,N_11543,N_11973);
or U15116 (N_15116,N_11441,N_9412);
nand U15117 (N_15117,N_11295,N_9951);
nand U15118 (N_15118,N_10015,N_12151);
nor U15119 (N_15119,N_11663,N_12024);
xor U15120 (N_15120,N_10666,N_10860);
nor U15121 (N_15121,N_10173,N_9773);
nand U15122 (N_15122,N_11285,N_9699);
nor U15123 (N_15123,N_11710,N_11521);
nand U15124 (N_15124,N_9758,N_11326);
and U15125 (N_15125,N_9494,N_11703);
xor U15126 (N_15126,N_9774,N_9776);
and U15127 (N_15127,N_11686,N_10080);
xnor U15128 (N_15128,N_10004,N_10720);
or U15129 (N_15129,N_10930,N_10912);
xor U15130 (N_15130,N_10538,N_10219);
nor U15131 (N_15131,N_11275,N_9502);
nor U15132 (N_15132,N_10922,N_12040);
xnor U15133 (N_15133,N_11069,N_11321);
or U15134 (N_15134,N_11911,N_11864);
nor U15135 (N_15135,N_9406,N_10865);
xor U15136 (N_15136,N_10706,N_12080);
and U15137 (N_15137,N_11660,N_9978);
or U15138 (N_15138,N_12175,N_9818);
or U15139 (N_15139,N_9519,N_11028);
or U15140 (N_15140,N_11891,N_12086);
nand U15141 (N_15141,N_11797,N_10640);
nor U15142 (N_15142,N_11354,N_10487);
nand U15143 (N_15143,N_10746,N_12126);
nor U15144 (N_15144,N_11430,N_9927);
nand U15145 (N_15145,N_10224,N_11541);
or U15146 (N_15146,N_9869,N_12322);
nor U15147 (N_15147,N_11386,N_11811);
nand U15148 (N_15148,N_10419,N_11036);
and U15149 (N_15149,N_12497,N_11132);
and U15150 (N_15150,N_12404,N_11469);
nor U15151 (N_15151,N_11989,N_10952);
nand U15152 (N_15152,N_12469,N_11844);
and U15153 (N_15153,N_11445,N_9998);
and U15154 (N_15154,N_12483,N_11101);
or U15155 (N_15155,N_10367,N_11319);
nor U15156 (N_15156,N_9722,N_10952);
xor U15157 (N_15157,N_10607,N_11040);
and U15158 (N_15158,N_12285,N_11701);
nor U15159 (N_15159,N_12368,N_9526);
nand U15160 (N_15160,N_11435,N_10595);
or U15161 (N_15161,N_12189,N_10125);
xnor U15162 (N_15162,N_11718,N_12339);
or U15163 (N_15163,N_10270,N_11519);
and U15164 (N_15164,N_12075,N_9770);
xnor U15165 (N_15165,N_12353,N_10932);
nand U15166 (N_15166,N_12152,N_9605);
nor U15167 (N_15167,N_9583,N_10376);
or U15168 (N_15168,N_11275,N_11430);
or U15169 (N_15169,N_9406,N_10612);
or U15170 (N_15170,N_11337,N_11420);
and U15171 (N_15171,N_12191,N_10219);
xnor U15172 (N_15172,N_11068,N_10115);
and U15173 (N_15173,N_10372,N_10877);
and U15174 (N_15174,N_12268,N_9837);
or U15175 (N_15175,N_9848,N_9671);
or U15176 (N_15176,N_11610,N_11541);
or U15177 (N_15177,N_9410,N_12410);
or U15178 (N_15178,N_9566,N_11791);
xnor U15179 (N_15179,N_10933,N_9375);
and U15180 (N_15180,N_10129,N_11665);
nand U15181 (N_15181,N_10399,N_9494);
or U15182 (N_15182,N_10087,N_12371);
nand U15183 (N_15183,N_12216,N_10747);
or U15184 (N_15184,N_10954,N_9446);
and U15185 (N_15185,N_10043,N_11507);
nand U15186 (N_15186,N_9461,N_10334);
and U15187 (N_15187,N_10391,N_9511);
or U15188 (N_15188,N_10061,N_12113);
nor U15189 (N_15189,N_9935,N_10657);
and U15190 (N_15190,N_10906,N_11325);
nor U15191 (N_15191,N_11754,N_10093);
nor U15192 (N_15192,N_9862,N_10408);
nor U15193 (N_15193,N_10192,N_12018);
and U15194 (N_15194,N_10842,N_10871);
and U15195 (N_15195,N_11397,N_10553);
nor U15196 (N_15196,N_9442,N_12084);
and U15197 (N_15197,N_10657,N_10321);
nor U15198 (N_15198,N_9902,N_10173);
and U15199 (N_15199,N_11826,N_11895);
nor U15200 (N_15200,N_11701,N_10203);
nor U15201 (N_15201,N_11546,N_11483);
or U15202 (N_15202,N_9661,N_11703);
nand U15203 (N_15203,N_10967,N_9601);
nor U15204 (N_15204,N_12227,N_10681);
and U15205 (N_15205,N_11045,N_10850);
and U15206 (N_15206,N_9931,N_10489);
and U15207 (N_15207,N_11875,N_10939);
and U15208 (N_15208,N_10224,N_11542);
or U15209 (N_15209,N_10519,N_11633);
or U15210 (N_15210,N_11577,N_11022);
xor U15211 (N_15211,N_11748,N_9742);
or U15212 (N_15212,N_12323,N_11194);
nor U15213 (N_15213,N_9961,N_12328);
nor U15214 (N_15214,N_10584,N_12225);
nand U15215 (N_15215,N_10097,N_11463);
nor U15216 (N_15216,N_11566,N_10272);
or U15217 (N_15217,N_10068,N_11420);
or U15218 (N_15218,N_11766,N_12165);
nor U15219 (N_15219,N_9812,N_11556);
nor U15220 (N_15220,N_12141,N_10573);
nor U15221 (N_15221,N_10335,N_11796);
and U15222 (N_15222,N_9566,N_10700);
or U15223 (N_15223,N_10114,N_12097);
nor U15224 (N_15224,N_10378,N_9940);
and U15225 (N_15225,N_10449,N_10952);
nand U15226 (N_15226,N_9893,N_12004);
nor U15227 (N_15227,N_11708,N_10812);
xor U15228 (N_15228,N_10860,N_12296);
nand U15229 (N_15229,N_10402,N_10811);
nor U15230 (N_15230,N_11999,N_9506);
or U15231 (N_15231,N_12497,N_11854);
nor U15232 (N_15232,N_10292,N_9958);
or U15233 (N_15233,N_9596,N_10907);
nand U15234 (N_15234,N_12338,N_11135);
or U15235 (N_15235,N_11115,N_9895);
xor U15236 (N_15236,N_12153,N_10949);
or U15237 (N_15237,N_9771,N_9709);
nand U15238 (N_15238,N_11615,N_11371);
nand U15239 (N_15239,N_9919,N_10796);
nor U15240 (N_15240,N_12379,N_12264);
nand U15241 (N_15241,N_9537,N_10437);
nor U15242 (N_15242,N_10376,N_10305);
nand U15243 (N_15243,N_12136,N_12114);
or U15244 (N_15244,N_11762,N_11615);
nor U15245 (N_15245,N_9962,N_12189);
or U15246 (N_15246,N_11992,N_9753);
nor U15247 (N_15247,N_9854,N_9889);
nor U15248 (N_15248,N_10627,N_10133);
nor U15249 (N_15249,N_12455,N_11592);
nand U15250 (N_15250,N_11350,N_9822);
or U15251 (N_15251,N_11023,N_12495);
nand U15252 (N_15252,N_9527,N_11095);
nor U15253 (N_15253,N_10060,N_10371);
and U15254 (N_15254,N_10790,N_10000);
nor U15255 (N_15255,N_10389,N_9794);
nand U15256 (N_15256,N_10270,N_10449);
or U15257 (N_15257,N_12348,N_9869);
nand U15258 (N_15258,N_11969,N_9443);
or U15259 (N_15259,N_12419,N_11398);
and U15260 (N_15260,N_10324,N_12403);
nor U15261 (N_15261,N_10514,N_9702);
nor U15262 (N_15262,N_10404,N_12374);
or U15263 (N_15263,N_9773,N_11386);
nor U15264 (N_15264,N_9727,N_12066);
nand U15265 (N_15265,N_12225,N_10065);
or U15266 (N_15266,N_11528,N_12335);
and U15267 (N_15267,N_11555,N_10298);
nand U15268 (N_15268,N_12200,N_9889);
nand U15269 (N_15269,N_11121,N_11424);
and U15270 (N_15270,N_11689,N_10157);
nand U15271 (N_15271,N_10837,N_9997);
nand U15272 (N_15272,N_12435,N_11458);
and U15273 (N_15273,N_12133,N_10868);
or U15274 (N_15274,N_10703,N_11475);
or U15275 (N_15275,N_11929,N_9795);
and U15276 (N_15276,N_10659,N_11202);
and U15277 (N_15277,N_10314,N_11761);
nor U15278 (N_15278,N_9952,N_9960);
xor U15279 (N_15279,N_11754,N_9584);
nand U15280 (N_15280,N_11078,N_12092);
nand U15281 (N_15281,N_10915,N_10886);
or U15282 (N_15282,N_12317,N_9488);
or U15283 (N_15283,N_11170,N_9892);
nand U15284 (N_15284,N_10704,N_9804);
nand U15285 (N_15285,N_11920,N_10445);
and U15286 (N_15286,N_11332,N_9939);
and U15287 (N_15287,N_9754,N_10176);
xnor U15288 (N_15288,N_11683,N_11112);
nand U15289 (N_15289,N_11528,N_12485);
nand U15290 (N_15290,N_10135,N_12070);
nor U15291 (N_15291,N_11760,N_12357);
or U15292 (N_15292,N_12198,N_9473);
and U15293 (N_15293,N_11612,N_12368);
or U15294 (N_15294,N_10550,N_10087);
nand U15295 (N_15295,N_10406,N_11153);
nand U15296 (N_15296,N_10047,N_9866);
and U15297 (N_15297,N_9535,N_12475);
xor U15298 (N_15298,N_11658,N_9458);
nor U15299 (N_15299,N_11323,N_11531);
and U15300 (N_15300,N_11065,N_10287);
or U15301 (N_15301,N_11844,N_12368);
and U15302 (N_15302,N_11402,N_10584);
and U15303 (N_15303,N_10227,N_9844);
and U15304 (N_15304,N_11997,N_10391);
nand U15305 (N_15305,N_9961,N_10323);
xor U15306 (N_15306,N_10313,N_9655);
or U15307 (N_15307,N_9979,N_12035);
nor U15308 (N_15308,N_10646,N_11870);
or U15309 (N_15309,N_12451,N_12309);
nand U15310 (N_15310,N_9539,N_12122);
or U15311 (N_15311,N_10085,N_12404);
nor U15312 (N_15312,N_11597,N_12245);
or U15313 (N_15313,N_11046,N_9377);
nor U15314 (N_15314,N_11881,N_10427);
nand U15315 (N_15315,N_11219,N_12081);
nand U15316 (N_15316,N_9446,N_9862);
nor U15317 (N_15317,N_10928,N_10006);
or U15318 (N_15318,N_10433,N_12333);
nor U15319 (N_15319,N_12080,N_11214);
or U15320 (N_15320,N_11815,N_10275);
nand U15321 (N_15321,N_10437,N_11121);
and U15322 (N_15322,N_11617,N_12059);
and U15323 (N_15323,N_10805,N_10058);
nor U15324 (N_15324,N_9536,N_12404);
nor U15325 (N_15325,N_10966,N_10310);
nor U15326 (N_15326,N_12499,N_10114);
and U15327 (N_15327,N_9828,N_11256);
and U15328 (N_15328,N_9870,N_11313);
xor U15329 (N_15329,N_9902,N_10726);
xnor U15330 (N_15330,N_10849,N_9750);
xnor U15331 (N_15331,N_10299,N_11825);
or U15332 (N_15332,N_11849,N_10667);
nand U15333 (N_15333,N_12134,N_11171);
and U15334 (N_15334,N_10372,N_10042);
nand U15335 (N_15335,N_10028,N_11629);
or U15336 (N_15336,N_11962,N_10290);
and U15337 (N_15337,N_10619,N_11493);
nor U15338 (N_15338,N_10558,N_11143);
nor U15339 (N_15339,N_12003,N_9973);
nand U15340 (N_15340,N_10160,N_12065);
nor U15341 (N_15341,N_10318,N_10321);
or U15342 (N_15342,N_11595,N_9972);
or U15343 (N_15343,N_11894,N_10346);
nor U15344 (N_15344,N_10536,N_9683);
nor U15345 (N_15345,N_10573,N_10662);
or U15346 (N_15346,N_9587,N_11659);
xnor U15347 (N_15347,N_10567,N_11841);
nand U15348 (N_15348,N_10696,N_10659);
nor U15349 (N_15349,N_11623,N_9546);
nand U15350 (N_15350,N_12153,N_11865);
xnor U15351 (N_15351,N_10791,N_11883);
and U15352 (N_15352,N_10707,N_9578);
nor U15353 (N_15353,N_12300,N_9693);
or U15354 (N_15354,N_9710,N_9746);
and U15355 (N_15355,N_11741,N_9375);
and U15356 (N_15356,N_11092,N_11522);
nand U15357 (N_15357,N_12054,N_12318);
nand U15358 (N_15358,N_10167,N_9452);
and U15359 (N_15359,N_11207,N_11606);
or U15360 (N_15360,N_10368,N_9513);
and U15361 (N_15361,N_12044,N_10211);
nand U15362 (N_15362,N_9560,N_9903);
nor U15363 (N_15363,N_11506,N_10351);
nand U15364 (N_15364,N_9403,N_12252);
nor U15365 (N_15365,N_10379,N_12322);
nand U15366 (N_15366,N_11658,N_9420);
and U15367 (N_15367,N_11664,N_9877);
nand U15368 (N_15368,N_11829,N_9883);
and U15369 (N_15369,N_9440,N_11844);
nand U15370 (N_15370,N_11293,N_12081);
or U15371 (N_15371,N_9452,N_9513);
or U15372 (N_15372,N_9977,N_12161);
and U15373 (N_15373,N_10478,N_10808);
nor U15374 (N_15374,N_11570,N_10511);
and U15375 (N_15375,N_11251,N_10182);
nand U15376 (N_15376,N_10544,N_10295);
xor U15377 (N_15377,N_10436,N_10798);
or U15378 (N_15378,N_9718,N_11122);
nor U15379 (N_15379,N_9464,N_11408);
nor U15380 (N_15380,N_10133,N_10267);
nand U15381 (N_15381,N_12051,N_10452);
nand U15382 (N_15382,N_10967,N_11037);
nand U15383 (N_15383,N_11565,N_11609);
or U15384 (N_15384,N_10941,N_10442);
nand U15385 (N_15385,N_11977,N_12287);
or U15386 (N_15386,N_11628,N_10493);
nor U15387 (N_15387,N_9398,N_10494);
and U15388 (N_15388,N_10228,N_12064);
or U15389 (N_15389,N_11152,N_12310);
or U15390 (N_15390,N_10549,N_9834);
and U15391 (N_15391,N_12193,N_11274);
or U15392 (N_15392,N_9842,N_10837);
nand U15393 (N_15393,N_11926,N_11083);
and U15394 (N_15394,N_10097,N_9821);
or U15395 (N_15395,N_10795,N_11813);
or U15396 (N_15396,N_10070,N_10353);
or U15397 (N_15397,N_11538,N_9569);
xor U15398 (N_15398,N_10089,N_11241);
and U15399 (N_15399,N_10984,N_11202);
or U15400 (N_15400,N_10165,N_9642);
nand U15401 (N_15401,N_12378,N_9419);
or U15402 (N_15402,N_11828,N_11613);
or U15403 (N_15403,N_10084,N_11193);
or U15404 (N_15404,N_9695,N_12271);
or U15405 (N_15405,N_10840,N_12477);
or U15406 (N_15406,N_12172,N_12379);
nor U15407 (N_15407,N_10698,N_11725);
nor U15408 (N_15408,N_11246,N_9627);
and U15409 (N_15409,N_10849,N_10411);
nand U15410 (N_15410,N_11086,N_12060);
nor U15411 (N_15411,N_9503,N_12232);
or U15412 (N_15412,N_9430,N_11711);
xor U15413 (N_15413,N_12155,N_10144);
nand U15414 (N_15414,N_9727,N_9617);
or U15415 (N_15415,N_10676,N_11216);
nor U15416 (N_15416,N_9472,N_9625);
and U15417 (N_15417,N_9454,N_12213);
and U15418 (N_15418,N_10330,N_9396);
nand U15419 (N_15419,N_11776,N_11426);
nand U15420 (N_15420,N_11133,N_11509);
and U15421 (N_15421,N_11943,N_12368);
or U15422 (N_15422,N_10487,N_9701);
and U15423 (N_15423,N_12296,N_9935);
or U15424 (N_15424,N_10154,N_10631);
and U15425 (N_15425,N_9543,N_11175);
and U15426 (N_15426,N_9755,N_10664);
nor U15427 (N_15427,N_9600,N_9636);
and U15428 (N_15428,N_11993,N_10745);
xnor U15429 (N_15429,N_10300,N_9854);
and U15430 (N_15430,N_12061,N_11401);
and U15431 (N_15431,N_9645,N_10858);
and U15432 (N_15432,N_11441,N_10782);
nor U15433 (N_15433,N_9503,N_10007);
and U15434 (N_15434,N_12422,N_12378);
or U15435 (N_15435,N_12033,N_10139);
and U15436 (N_15436,N_10580,N_10470);
and U15437 (N_15437,N_10078,N_11372);
and U15438 (N_15438,N_10850,N_9810);
nand U15439 (N_15439,N_10705,N_11288);
nand U15440 (N_15440,N_10198,N_11756);
nor U15441 (N_15441,N_11054,N_10879);
or U15442 (N_15442,N_11585,N_10450);
nand U15443 (N_15443,N_10497,N_10923);
or U15444 (N_15444,N_12290,N_11799);
nand U15445 (N_15445,N_12466,N_9445);
nor U15446 (N_15446,N_9512,N_11918);
or U15447 (N_15447,N_10743,N_12275);
and U15448 (N_15448,N_9829,N_11300);
nand U15449 (N_15449,N_11337,N_9419);
and U15450 (N_15450,N_10040,N_11364);
nor U15451 (N_15451,N_11049,N_10192);
nand U15452 (N_15452,N_10373,N_10407);
nand U15453 (N_15453,N_9462,N_9903);
nor U15454 (N_15454,N_11006,N_9427);
and U15455 (N_15455,N_9900,N_11468);
nand U15456 (N_15456,N_11975,N_11785);
or U15457 (N_15457,N_10705,N_11536);
nor U15458 (N_15458,N_11368,N_11444);
nand U15459 (N_15459,N_9516,N_10777);
nand U15460 (N_15460,N_9682,N_10098);
xor U15461 (N_15461,N_11629,N_9375);
and U15462 (N_15462,N_10675,N_12318);
or U15463 (N_15463,N_10673,N_12472);
nand U15464 (N_15464,N_12480,N_9480);
nor U15465 (N_15465,N_12013,N_10804);
or U15466 (N_15466,N_12190,N_11298);
and U15467 (N_15467,N_9988,N_12121);
nor U15468 (N_15468,N_10173,N_10878);
or U15469 (N_15469,N_11492,N_10456);
and U15470 (N_15470,N_11323,N_10531);
nand U15471 (N_15471,N_10075,N_12258);
nand U15472 (N_15472,N_11884,N_11075);
and U15473 (N_15473,N_10047,N_9617);
nor U15474 (N_15474,N_11031,N_9643);
and U15475 (N_15475,N_11453,N_9550);
and U15476 (N_15476,N_11038,N_10857);
and U15477 (N_15477,N_9774,N_12234);
xnor U15478 (N_15478,N_12220,N_10652);
or U15479 (N_15479,N_10342,N_11884);
nand U15480 (N_15480,N_9757,N_11215);
or U15481 (N_15481,N_10300,N_12213);
or U15482 (N_15482,N_10579,N_11161);
nand U15483 (N_15483,N_10115,N_10854);
nand U15484 (N_15484,N_9451,N_11200);
nor U15485 (N_15485,N_10018,N_9741);
nor U15486 (N_15486,N_12068,N_11238);
or U15487 (N_15487,N_10557,N_10870);
or U15488 (N_15488,N_10183,N_12364);
nand U15489 (N_15489,N_10766,N_10948);
nor U15490 (N_15490,N_12471,N_10282);
nor U15491 (N_15491,N_12362,N_10135);
or U15492 (N_15492,N_10975,N_11263);
or U15493 (N_15493,N_11979,N_11112);
or U15494 (N_15494,N_9774,N_12194);
or U15495 (N_15495,N_11235,N_12116);
nor U15496 (N_15496,N_11465,N_10035);
nand U15497 (N_15497,N_11909,N_10126);
and U15498 (N_15498,N_10305,N_10233);
nor U15499 (N_15499,N_11474,N_10676);
xor U15500 (N_15500,N_10439,N_10428);
xor U15501 (N_15501,N_10080,N_10724);
or U15502 (N_15502,N_11785,N_9619);
nand U15503 (N_15503,N_10474,N_9960);
nand U15504 (N_15504,N_11155,N_11094);
nand U15505 (N_15505,N_10103,N_10447);
and U15506 (N_15506,N_10142,N_10272);
and U15507 (N_15507,N_9534,N_9414);
nor U15508 (N_15508,N_10875,N_11818);
nand U15509 (N_15509,N_10291,N_9683);
nor U15510 (N_15510,N_11297,N_10770);
nand U15511 (N_15511,N_11707,N_12381);
nand U15512 (N_15512,N_12337,N_11358);
and U15513 (N_15513,N_10692,N_9834);
or U15514 (N_15514,N_10350,N_9952);
nand U15515 (N_15515,N_11414,N_10588);
and U15516 (N_15516,N_11067,N_12079);
nor U15517 (N_15517,N_10685,N_10012);
nand U15518 (N_15518,N_11670,N_11451);
nor U15519 (N_15519,N_12050,N_11469);
xnor U15520 (N_15520,N_10993,N_11338);
and U15521 (N_15521,N_10063,N_10533);
or U15522 (N_15522,N_10985,N_9539);
nor U15523 (N_15523,N_9834,N_10629);
nor U15524 (N_15524,N_9998,N_9870);
and U15525 (N_15525,N_12298,N_12407);
nor U15526 (N_15526,N_11467,N_11081);
or U15527 (N_15527,N_11613,N_11146);
or U15528 (N_15528,N_10167,N_11764);
and U15529 (N_15529,N_11764,N_11135);
nand U15530 (N_15530,N_11282,N_10063);
nor U15531 (N_15531,N_11286,N_12044);
xnor U15532 (N_15532,N_12466,N_11148);
or U15533 (N_15533,N_11735,N_11228);
and U15534 (N_15534,N_10734,N_9444);
and U15535 (N_15535,N_10189,N_9717);
nor U15536 (N_15536,N_9701,N_10904);
nand U15537 (N_15537,N_9906,N_10553);
and U15538 (N_15538,N_12234,N_11129);
nor U15539 (N_15539,N_12199,N_12051);
or U15540 (N_15540,N_10728,N_9865);
nand U15541 (N_15541,N_10765,N_11275);
and U15542 (N_15542,N_12192,N_11369);
and U15543 (N_15543,N_11516,N_9533);
and U15544 (N_15544,N_10424,N_9574);
or U15545 (N_15545,N_11246,N_10153);
nor U15546 (N_15546,N_9922,N_11705);
nand U15547 (N_15547,N_11007,N_9862);
or U15548 (N_15548,N_9881,N_10140);
and U15549 (N_15549,N_9939,N_11004);
xnor U15550 (N_15550,N_11930,N_10633);
nor U15551 (N_15551,N_11932,N_10512);
nor U15552 (N_15552,N_11061,N_10214);
nand U15553 (N_15553,N_10655,N_11984);
or U15554 (N_15554,N_12085,N_11391);
or U15555 (N_15555,N_10540,N_12118);
nand U15556 (N_15556,N_9477,N_9718);
and U15557 (N_15557,N_9918,N_9392);
or U15558 (N_15558,N_12327,N_9804);
nand U15559 (N_15559,N_11753,N_11372);
xor U15560 (N_15560,N_11694,N_10123);
nand U15561 (N_15561,N_11953,N_11726);
or U15562 (N_15562,N_11778,N_11751);
and U15563 (N_15563,N_9562,N_10921);
or U15564 (N_15564,N_9769,N_11137);
nand U15565 (N_15565,N_9472,N_9591);
or U15566 (N_15566,N_9968,N_11996);
or U15567 (N_15567,N_10511,N_12148);
or U15568 (N_15568,N_10256,N_10923);
xnor U15569 (N_15569,N_9870,N_9539);
and U15570 (N_15570,N_10631,N_11319);
nor U15571 (N_15571,N_10710,N_9673);
nand U15572 (N_15572,N_9805,N_11049);
and U15573 (N_15573,N_11778,N_12313);
or U15574 (N_15574,N_10499,N_11388);
nor U15575 (N_15575,N_11476,N_10106);
nand U15576 (N_15576,N_10215,N_11987);
nor U15577 (N_15577,N_10996,N_11039);
xor U15578 (N_15578,N_10225,N_12298);
and U15579 (N_15579,N_11323,N_9637);
or U15580 (N_15580,N_10539,N_10726);
or U15581 (N_15581,N_10696,N_11992);
nor U15582 (N_15582,N_11465,N_10217);
nand U15583 (N_15583,N_10507,N_12085);
and U15584 (N_15584,N_12061,N_10596);
and U15585 (N_15585,N_11231,N_10434);
and U15586 (N_15586,N_9843,N_11396);
nor U15587 (N_15587,N_9746,N_11591);
nand U15588 (N_15588,N_11409,N_9395);
and U15589 (N_15589,N_10328,N_10421);
or U15590 (N_15590,N_9406,N_11170);
nor U15591 (N_15591,N_9932,N_11355);
or U15592 (N_15592,N_10672,N_11052);
nor U15593 (N_15593,N_11643,N_9460);
and U15594 (N_15594,N_12221,N_11027);
nor U15595 (N_15595,N_12051,N_9468);
and U15596 (N_15596,N_11036,N_11506);
nand U15597 (N_15597,N_12476,N_9954);
nor U15598 (N_15598,N_10302,N_11493);
nand U15599 (N_15599,N_12124,N_10740);
nand U15600 (N_15600,N_10940,N_10589);
and U15601 (N_15601,N_11612,N_12158);
nand U15602 (N_15602,N_11148,N_10083);
or U15603 (N_15603,N_10375,N_9415);
nor U15604 (N_15604,N_10069,N_10930);
nand U15605 (N_15605,N_12344,N_12161);
or U15606 (N_15606,N_11778,N_10635);
nor U15607 (N_15607,N_9846,N_11006);
or U15608 (N_15608,N_10711,N_10256);
nand U15609 (N_15609,N_12174,N_9779);
or U15610 (N_15610,N_10861,N_10938);
nor U15611 (N_15611,N_11126,N_10765);
nor U15612 (N_15612,N_9613,N_11727);
and U15613 (N_15613,N_11127,N_9719);
nand U15614 (N_15614,N_10287,N_9794);
or U15615 (N_15615,N_9823,N_12098);
nor U15616 (N_15616,N_9469,N_11387);
or U15617 (N_15617,N_9945,N_10801);
nand U15618 (N_15618,N_10629,N_10785);
or U15619 (N_15619,N_11630,N_11365);
nand U15620 (N_15620,N_11231,N_10184);
or U15621 (N_15621,N_11673,N_12218);
nor U15622 (N_15622,N_11891,N_10767);
or U15623 (N_15623,N_9672,N_9522);
and U15624 (N_15624,N_11260,N_11152);
nand U15625 (N_15625,N_12813,N_15030);
nor U15626 (N_15626,N_14603,N_13153);
and U15627 (N_15627,N_14594,N_14573);
xnor U15628 (N_15628,N_15558,N_15287);
or U15629 (N_15629,N_12512,N_15512);
and U15630 (N_15630,N_13337,N_12577);
nand U15631 (N_15631,N_12574,N_14254);
and U15632 (N_15632,N_14045,N_14305);
nor U15633 (N_15633,N_14734,N_12689);
nand U15634 (N_15634,N_15484,N_14372);
xnor U15635 (N_15635,N_13742,N_12620);
nand U15636 (N_15636,N_12593,N_13871);
or U15637 (N_15637,N_15439,N_14685);
or U15638 (N_15638,N_12985,N_14286);
nand U15639 (N_15639,N_14808,N_13213);
nor U15640 (N_15640,N_14052,N_15070);
and U15641 (N_15641,N_15243,N_14447);
nor U15642 (N_15642,N_12789,N_14561);
or U15643 (N_15643,N_12629,N_14905);
xnor U15644 (N_15644,N_14716,N_13204);
and U15645 (N_15645,N_12876,N_15379);
nand U15646 (N_15646,N_14966,N_14066);
or U15647 (N_15647,N_13293,N_15536);
xnor U15648 (N_15648,N_14365,N_13815);
or U15649 (N_15649,N_14710,N_14773);
nor U15650 (N_15650,N_14162,N_12653);
and U15651 (N_15651,N_13238,N_13864);
nor U15652 (N_15652,N_13068,N_15338);
nor U15653 (N_15653,N_14706,N_13459);
and U15654 (N_15654,N_12909,N_14415);
nand U15655 (N_15655,N_12527,N_15072);
or U15656 (N_15656,N_12896,N_12592);
nor U15657 (N_15657,N_15275,N_14761);
nand U15658 (N_15658,N_13217,N_14376);
nor U15659 (N_15659,N_12646,N_13012);
nor U15660 (N_15660,N_12591,N_15292);
nand U15661 (N_15661,N_15028,N_15541);
and U15662 (N_15662,N_15443,N_12524);
xnor U15663 (N_15663,N_13946,N_15180);
nor U15664 (N_15664,N_14221,N_14770);
nor U15665 (N_15665,N_14641,N_13721);
xnor U15666 (N_15666,N_13673,N_15010);
nor U15667 (N_15667,N_14965,N_13906);
nor U15668 (N_15668,N_14954,N_14334);
and U15669 (N_15669,N_14512,N_14886);
and U15670 (N_15670,N_14395,N_15083);
xnor U15671 (N_15671,N_15502,N_15049);
or U15672 (N_15672,N_13642,N_14830);
nor U15673 (N_15673,N_13967,N_15055);
and U15674 (N_15674,N_12709,N_12777);
or U15675 (N_15675,N_14549,N_15378);
xor U15676 (N_15676,N_13802,N_12587);
nor U15677 (N_15677,N_15493,N_12768);
nor U15678 (N_15678,N_14633,N_12585);
nor U15679 (N_15679,N_14950,N_13892);
and U15680 (N_15680,N_13001,N_15230);
nand U15681 (N_15681,N_12847,N_15510);
or U15682 (N_15682,N_12949,N_14592);
nand U15683 (N_15683,N_15377,N_14064);
or U15684 (N_15684,N_12690,N_13912);
xnor U15685 (N_15685,N_15468,N_14956);
nand U15686 (N_15686,N_13395,N_14964);
or U15687 (N_15687,N_12866,N_15156);
nor U15688 (N_15688,N_14851,N_14374);
or U15689 (N_15689,N_14361,N_15426);
or U15690 (N_15690,N_15238,N_13883);
or U15691 (N_15691,N_13242,N_14292);
xor U15692 (N_15692,N_12739,N_14308);
and U15693 (N_15693,N_13463,N_15508);
nand U15694 (N_15694,N_13273,N_14503);
nor U15695 (N_15695,N_12658,N_15556);
or U15696 (N_15696,N_14417,N_13179);
xnor U15697 (N_15697,N_13531,N_13415);
and U15698 (N_15698,N_14547,N_14164);
nand U15699 (N_15699,N_14607,N_15150);
and U15700 (N_15700,N_13552,N_14934);
xnor U15701 (N_15701,N_13438,N_12517);
nor U15702 (N_15702,N_14586,N_14514);
nand U15703 (N_15703,N_13601,N_12553);
xor U15704 (N_15704,N_14195,N_14980);
nand U15705 (N_15705,N_15020,N_12693);
and U15706 (N_15706,N_15600,N_13882);
nand U15707 (N_15707,N_14459,N_13482);
nand U15708 (N_15708,N_12586,N_13466);
and U15709 (N_15709,N_14754,N_12819);
nand U15710 (N_15710,N_15285,N_13751);
or U15711 (N_15711,N_14914,N_13465);
and U15712 (N_15712,N_13903,N_14590);
nor U15713 (N_15713,N_15572,N_15110);
and U15714 (N_15714,N_14485,N_12665);
and U15715 (N_15715,N_13738,N_14461);
nand U15716 (N_15716,N_14427,N_13306);
nand U15717 (N_15717,N_13402,N_15181);
and U15718 (N_15718,N_14546,N_13890);
or U15719 (N_15719,N_13403,N_15056);
and U15720 (N_15720,N_12976,N_14733);
or U15721 (N_15721,N_14071,N_12862);
or U15722 (N_15722,N_15267,N_15463);
or U15723 (N_15723,N_15079,N_13959);
or U15724 (N_15724,N_13610,N_12856);
nand U15725 (N_15725,N_14917,N_12661);
nor U15726 (N_15726,N_13520,N_14139);
nand U15727 (N_15727,N_13763,N_15179);
or U15728 (N_15728,N_14516,N_14029);
nor U15729 (N_15729,N_13231,N_13176);
nand U15730 (N_15730,N_15245,N_14636);
and U15731 (N_15731,N_13529,N_12990);
nand U15732 (N_15732,N_14741,N_12506);
xnor U15733 (N_15733,N_14036,N_13362);
or U15734 (N_15734,N_13343,N_14751);
and U15735 (N_15735,N_14337,N_15337);
xor U15736 (N_15736,N_14253,N_12897);
and U15737 (N_15737,N_12830,N_14588);
and U15738 (N_15738,N_14882,N_14656);
or U15739 (N_15739,N_15399,N_13135);
nand U15740 (N_15740,N_13447,N_13506);
or U15741 (N_15741,N_12817,N_13338);
nand U15742 (N_15742,N_14646,N_14405);
and U15743 (N_15743,N_14853,N_14082);
or U15744 (N_15744,N_15587,N_15575);
and U15745 (N_15745,N_13521,N_13608);
nor U15746 (N_15746,N_13858,N_14236);
nand U15747 (N_15747,N_14911,N_15196);
nand U15748 (N_15748,N_12843,N_13874);
or U15749 (N_15749,N_14432,N_14113);
and U15750 (N_15750,N_14739,N_15359);
and U15751 (N_15751,N_12511,N_14868);
xor U15752 (N_15752,N_13487,N_15316);
and U15753 (N_15753,N_14524,N_13114);
or U15754 (N_15754,N_15246,N_12718);
nand U15755 (N_15755,N_14217,N_13455);
nand U15756 (N_15756,N_13607,N_12628);
or U15757 (N_15757,N_13046,N_12598);
or U15758 (N_15758,N_14848,N_15041);
nor U15759 (N_15759,N_14854,N_14540);
xnor U15760 (N_15760,N_15244,N_14347);
xor U15761 (N_15761,N_13593,N_14210);
and U15762 (N_15762,N_13619,N_13299);
xnor U15763 (N_15763,N_15325,N_14811);
xor U15764 (N_15764,N_13737,N_13060);
and U15765 (N_15765,N_13232,N_14428);
nand U15766 (N_15766,N_12713,N_13705);
nand U15767 (N_15767,N_15237,N_12853);
and U15768 (N_15768,N_15423,N_12998);
nand U15769 (N_15769,N_15547,N_12963);
xor U15770 (N_15770,N_14765,N_13988);
xnor U15771 (N_15771,N_13128,N_13361);
nor U15772 (N_15772,N_15159,N_12699);
nor U15773 (N_15773,N_15405,N_14440);
nor U15774 (N_15774,N_12670,N_14198);
nand U15775 (N_15775,N_12698,N_12980);
and U15776 (N_15776,N_14789,N_15537);
nor U15777 (N_15777,N_14595,N_14898);
or U15778 (N_15778,N_13308,N_13494);
xnor U15779 (N_15779,N_15226,N_15097);
or U15780 (N_15780,N_13430,N_15622);
nor U15781 (N_15781,N_15497,N_14916);
or U15782 (N_15782,N_12618,N_12924);
nor U15783 (N_15783,N_12728,N_14431);
and U15784 (N_15784,N_12735,N_12773);
nand U15785 (N_15785,N_12941,N_15217);
nor U15786 (N_15786,N_14842,N_13022);
nor U15787 (N_15787,N_14460,N_13781);
nand U15788 (N_15788,N_13160,N_15099);
nand U15789 (N_15789,N_12951,N_13942);
xor U15790 (N_15790,N_15588,N_15216);
and U15791 (N_15791,N_14653,N_14631);
xor U15792 (N_15792,N_14737,N_14904);
xor U15793 (N_15793,N_15323,N_15438);
xor U15794 (N_15794,N_15569,N_15074);
xor U15795 (N_15795,N_13687,N_13212);
or U15796 (N_15796,N_13066,N_12855);
nand U15797 (N_15797,N_12624,N_12991);
or U15798 (N_15798,N_13765,N_14609);
nor U15799 (N_15799,N_15584,N_12753);
and U15800 (N_15800,N_12903,N_13379);
or U15801 (N_15801,N_15094,N_13806);
nor U15802 (N_15802,N_13331,N_13196);
or U15803 (N_15803,N_12717,N_15448);
or U15804 (N_15804,N_13978,N_14368);
xor U15805 (N_15805,N_14735,N_15123);
nand U15806 (N_15806,N_12549,N_13834);
nor U15807 (N_15807,N_12759,N_12799);
and U15808 (N_15808,N_15040,N_15376);
or U15809 (N_15809,N_14475,N_13477);
and U15810 (N_15810,N_13905,N_14795);
or U15811 (N_15811,N_14785,N_15224);
nand U15812 (N_15812,N_13023,N_14130);
or U15813 (N_15813,N_15103,N_13002);
xor U15814 (N_15814,N_12548,N_12842);
or U15815 (N_15815,N_13872,N_12883);
nor U15816 (N_15816,N_14004,N_14788);
and U15817 (N_15817,N_13827,N_13382);
nand U15818 (N_15818,N_14065,N_14200);
nor U15819 (N_15819,N_12934,N_12617);
nand U15820 (N_15820,N_14570,N_15252);
nor U15821 (N_15821,N_13021,N_13133);
or U15822 (N_15822,N_13790,N_15520);
and U15823 (N_15823,N_15501,N_14274);
or U15824 (N_15824,N_12938,N_14659);
and U15825 (N_15825,N_15551,N_14304);
nand U15826 (N_15826,N_14243,N_13836);
and U15827 (N_15827,N_14942,N_14939);
nor U15828 (N_15828,N_14907,N_13869);
or U15829 (N_15829,N_15225,N_12541);
nand U15830 (N_15830,N_13649,N_12810);
nand U15831 (N_15831,N_15539,N_13678);
nor U15832 (N_15832,N_14426,N_13537);
or U15833 (N_15833,N_15073,N_13983);
xnor U15834 (N_15834,N_14801,N_15190);
nand U15835 (N_15835,N_13569,N_14507);
or U15836 (N_15836,N_14324,N_12892);
or U15837 (N_15837,N_15619,N_13853);
xnor U15838 (N_15838,N_13694,N_12737);
and U15839 (N_15839,N_14193,N_13436);
nor U15840 (N_15840,N_13107,N_12879);
nor U15841 (N_15841,N_13211,N_12751);
nand U15842 (N_15842,N_14545,N_13434);
and U15843 (N_15843,N_13604,N_12516);
and U15844 (N_15844,N_14229,N_13165);
or U15845 (N_15845,N_15606,N_15249);
and U15846 (N_15846,N_15408,N_13252);
nand U15847 (N_15847,N_13230,N_15404);
and U15848 (N_15848,N_14348,N_14976);
or U15849 (N_15849,N_12568,N_15467);
nor U15850 (N_15850,N_15290,N_13750);
nand U15851 (N_15851,N_14060,N_13258);
or U15852 (N_15852,N_12956,N_14177);
nor U15853 (N_15853,N_14730,N_14430);
nand U15854 (N_15854,N_12555,N_13224);
xor U15855 (N_15855,N_12538,N_14564);
nand U15856 (N_15856,N_13866,N_14975);
and U15857 (N_15857,N_13507,N_14552);
nor U15858 (N_15858,N_14600,N_14419);
or U15859 (N_15859,N_13198,N_12543);
xnor U15860 (N_15860,N_15057,N_12796);
nand U15861 (N_15861,N_13123,N_13683);
nor U15862 (N_15862,N_14894,N_13691);
nand U15863 (N_15863,N_14481,N_13272);
nor U15864 (N_15864,N_12521,N_15415);
and U15865 (N_15865,N_14682,N_13805);
xnor U15866 (N_15866,N_14100,N_13907);
or U15867 (N_15867,N_15223,N_13227);
nand U15868 (N_15868,N_14483,N_15340);
or U15869 (N_15869,N_14442,N_12657);
nor U15870 (N_15870,N_15349,N_15106);
nand U15871 (N_15871,N_15276,N_15478);
xor U15872 (N_15872,N_14208,N_14913);
nor U15873 (N_15873,N_14157,N_13077);
and U15874 (N_15874,N_14703,N_15436);
and U15875 (N_15875,N_15117,N_12943);
or U15876 (N_15876,N_13398,N_13072);
nand U15877 (N_15877,N_14783,N_15538);
xor U15878 (N_15878,N_13894,N_15042);
and U15879 (N_15879,N_13467,N_14420);
and U15880 (N_15880,N_13911,N_12684);
and U15881 (N_15881,N_13154,N_15362);
and U15882 (N_15882,N_13980,N_13734);
nand U15883 (N_15883,N_14194,N_12958);
nor U15884 (N_15884,N_12864,N_15194);
nand U15885 (N_15885,N_13847,N_13645);
or U15886 (N_15886,N_13784,N_15026);
or U15887 (N_15887,N_14138,N_13510);
nand U15888 (N_15888,N_14018,N_14434);
nand U15889 (N_15889,N_14252,N_15477);
and U15890 (N_15890,N_13711,N_13860);
xor U15891 (N_15891,N_15603,N_15534);
and U15892 (N_15892,N_14903,N_13208);
nand U15893 (N_15893,N_12845,N_15302);
nor U15894 (N_15894,N_14134,N_12588);
nor U15895 (N_15895,N_14127,N_13307);
nand U15896 (N_15896,N_13798,N_14617);
nand U15897 (N_15897,N_14445,N_14694);
nor U15898 (N_15898,N_15431,N_13084);
or U15899 (N_15899,N_15419,N_14167);
nor U15900 (N_15900,N_14019,N_12584);
or U15901 (N_15901,N_12606,N_13950);
nor U15902 (N_15902,N_14081,N_13803);
nand U15903 (N_15903,N_14862,N_14798);
nor U15904 (N_15904,N_13493,N_14152);
nand U15905 (N_15905,N_13662,N_13094);
nor U15906 (N_15906,N_15367,N_13096);
or U15907 (N_15907,N_15183,N_15453);
or U15908 (N_15908,N_14794,N_15108);
and U15909 (N_15909,N_14335,N_13536);
or U15910 (N_15910,N_14443,N_15071);
or U15911 (N_15911,N_13178,N_13939);
or U15912 (N_15912,N_15387,N_14363);
or U15913 (N_15913,N_15372,N_14743);
or U15914 (N_15914,N_13106,N_14073);
nand U15915 (N_15915,N_12576,N_14836);
nor U15916 (N_15916,N_14380,N_14366);
and U15917 (N_15917,N_13615,N_14752);
nor U15918 (N_15918,N_13885,N_14702);
nand U15919 (N_15919,N_15457,N_12659);
nand U15920 (N_15920,N_13666,N_14247);
xor U15921 (N_15921,N_12560,N_13443);
or U15922 (N_15922,N_13342,N_14323);
or U15923 (N_15923,N_15332,N_13192);
nand U15924 (N_15924,N_13201,N_12723);
xnor U15925 (N_15925,N_15229,N_14952);
or U15926 (N_15926,N_13508,N_14206);
or U15927 (N_15927,N_12849,N_13358);
and U15928 (N_15928,N_13605,N_14557);
nand U15929 (N_15929,N_12989,N_13914);
and U15930 (N_15930,N_14762,N_15442);
xnor U15931 (N_15931,N_13136,N_14989);
and U15932 (N_15932,N_13512,N_12614);
and U15933 (N_15933,N_13100,N_15413);
and U15934 (N_15934,N_14992,N_13356);
or U15935 (N_15935,N_14303,N_13938);
and U15936 (N_15936,N_13093,N_14606);
or U15937 (N_15937,N_13731,N_14219);
nor U15938 (N_15938,N_14930,N_15096);
or U15939 (N_15939,N_12904,N_13281);
xor U15940 (N_15940,N_15218,N_14963);
and U15941 (N_15941,N_13902,N_13219);
nand U15942 (N_15942,N_14471,N_14054);
nor U15943 (N_15943,N_14046,N_15306);
or U15944 (N_15944,N_12537,N_14926);
and U15945 (N_15945,N_15578,N_13164);
nor U15946 (N_15946,N_13053,N_14076);
and U15947 (N_15947,N_13011,N_14291);
or U15948 (N_15948,N_15565,N_13530);
nor U15949 (N_15949,N_13057,N_12884);
nand U15950 (N_15950,N_13524,N_13188);
and U15951 (N_15951,N_13652,N_14259);
nand U15952 (N_15952,N_12979,N_14556);
nor U15953 (N_15953,N_13071,N_15441);
nand U15954 (N_15954,N_14387,N_12877);
nand U15955 (N_15955,N_13875,N_14179);
and U15956 (N_15956,N_14297,N_15585);
or U15957 (N_15957,N_15164,N_13714);
nor U15958 (N_15958,N_12762,N_14007);
nand U15959 (N_15959,N_15045,N_13899);
nand U15960 (N_15960,N_13915,N_13909);
xor U15961 (N_15961,N_12935,N_14790);
nand U15962 (N_15962,N_12615,N_12542);
nor U15963 (N_15963,N_13326,N_14016);
xnor U15964 (N_15964,N_13701,N_14643);
xnor U15965 (N_15965,N_14627,N_13920);
nand U15966 (N_15966,N_13376,N_12836);
or U15967 (N_15967,N_13410,N_15490);
or U15968 (N_15968,N_13103,N_14355);
or U15969 (N_15969,N_13565,N_12695);
nor U15970 (N_15970,N_13868,N_13431);
nand U15971 (N_15971,N_15552,N_15014);
or U15972 (N_15972,N_13095,N_13218);
or U15973 (N_15973,N_12648,N_13809);
or U15974 (N_15974,N_14978,N_13743);
nand U15975 (N_15975,N_14448,N_13378);
or U15976 (N_15976,N_13917,N_15345);
nor U15977 (N_15977,N_13474,N_14924);
or U15978 (N_15978,N_15261,N_14920);
nand U15979 (N_15979,N_13172,N_13710);
or U15980 (N_15980,N_12716,N_13413);
nand U15981 (N_15981,N_13586,N_14698);
nand U15982 (N_15982,N_14186,N_12922);
and U15983 (N_15983,N_14791,N_14002);
or U15984 (N_15984,N_14116,N_14582);
nor U15985 (N_15985,N_13774,N_14213);
nor U15986 (N_15986,N_13086,N_12525);
nor U15987 (N_15987,N_13045,N_12507);
or U15988 (N_15988,N_15235,N_15432);
and U15989 (N_15989,N_12895,N_13500);
nor U15990 (N_15990,N_13812,N_14784);
xor U15991 (N_15991,N_12596,N_12707);
nand U15992 (N_15992,N_14820,N_14416);
nand U15993 (N_15993,N_13274,N_13458);
nor U15994 (N_15994,N_15182,N_12748);
nor U15995 (N_15995,N_13703,N_13748);
or U15996 (N_15996,N_13422,N_15564);
nor U15997 (N_15997,N_13177,N_13654);
and U15998 (N_15998,N_13202,N_14386);
nand U15999 (N_15999,N_13729,N_13193);
or U16000 (N_16000,N_14940,N_14639);
nand U16001 (N_16001,N_14747,N_15589);
nand U16002 (N_16002,N_13638,N_14185);
and U16003 (N_16003,N_12993,N_14893);
or U16004 (N_16004,N_14285,N_13304);
nor U16005 (N_16005,N_14970,N_12582);
nor U16006 (N_16006,N_15250,N_15595);
and U16007 (N_16007,N_14439,N_14424);
nand U16008 (N_16008,N_13736,N_13725);
and U16009 (N_16009,N_13837,N_15416);
xnor U16010 (N_16010,N_14038,N_14080);
or U16011 (N_16011,N_15029,N_14539);
nand U16012 (N_16012,N_12656,N_13291);
and U16013 (N_16013,N_14981,N_12552);
nand U16014 (N_16014,N_13576,N_14035);
nor U16015 (N_16015,N_12821,N_14345);
nand U16016 (N_16016,N_12678,N_14482);
nor U16017 (N_16017,N_13928,N_12832);
nor U16018 (N_16018,N_13419,N_15363);
and U16019 (N_16019,N_15168,N_13541);
xor U16020 (N_16020,N_13375,N_13665);
and U16021 (N_16021,N_13448,N_14070);
and U16022 (N_16022,N_15279,N_14377);
nor U16023 (N_16023,N_12686,N_13637);
and U16024 (N_16024,N_14068,N_14296);
nor U16025 (N_16025,N_15100,N_14937);
nor U16026 (N_16026,N_13561,N_15483);
and U16027 (N_16027,N_15059,N_13795);
and U16028 (N_16028,N_12929,N_14040);
and U16029 (N_16029,N_15315,N_12936);
nand U16030 (N_16030,N_12633,N_13492);
nor U16031 (N_16031,N_15128,N_12634);
nand U16032 (N_16032,N_14768,N_14147);
and U16033 (N_16033,N_14159,N_15195);
or U16034 (N_16034,N_14585,N_14058);
xnor U16035 (N_16035,N_13515,N_12974);
or U16036 (N_16036,N_13570,N_14536);
and U16037 (N_16037,N_12649,N_12581);
nand U16038 (N_16038,N_13782,N_12679);
xor U16039 (N_16039,N_14776,N_13689);
xnor U16040 (N_16040,N_13149,N_13733);
xnor U16041 (N_16041,N_14425,N_12613);
or U16042 (N_16042,N_13353,N_12824);
xnor U16043 (N_16043,N_14771,N_14227);
and U16044 (N_16044,N_13651,N_14034);
and U16045 (N_16045,N_14654,N_15360);
or U16046 (N_16046,N_15215,N_15482);
or U16047 (N_16047,N_13083,N_12607);
or U16048 (N_16048,N_14568,N_12964);
and U16049 (N_16049,N_15308,N_15104);
xnor U16050 (N_16050,N_13594,N_13505);
nor U16051 (N_16051,N_13157,N_13420);
or U16052 (N_16052,N_13551,N_15139);
nand U16053 (N_16053,N_14928,N_12962);
and U16054 (N_16054,N_14072,N_12988);
and U16055 (N_16055,N_12816,N_15339);
nand U16056 (N_16056,N_14490,N_13937);
or U16057 (N_16057,N_13648,N_14199);
and U16058 (N_16058,N_14182,N_13363);
nand U16059 (N_16059,N_13706,N_13484);
nor U16060 (N_16060,N_15444,N_13377);
nor U16061 (N_16061,N_12647,N_15007);
xor U16062 (N_16062,N_13661,N_14091);
nor U16063 (N_16063,N_13502,N_14088);
nor U16064 (N_16064,N_14242,N_15371);
and U16065 (N_16065,N_12966,N_14156);
and U16066 (N_16066,N_13409,N_15296);
nand U16067 (N_16067,N_13617,N_14013);
or U16068 (N_16068,N_14745,N_12928);
and U16069 (N_16069,N_13519,N_13181);
nand U16070 (N_16070,N_13264,N_13813);
nor U16071 (N_16071,N_14676,N_13089);
and U16072 (N_16072,N_13854,N_12960);
or U16073 (N_16073,N_14878,N_13295);
and U16074 (N_16074,N_15003,N_13732);
nand U16075 (N_16075,N_15260,N_14844);
nand U16076 (N_16076,N_14406,N_15542);
nor U16077 (N_16077,N_12975,N_14160);
or U16078 (N_16078,N_14895,N_13595);
nor U16079 (N_16079,N_15544,N_13807);
or U16080 (N_16080,N_14810,N_13048);
or U16081 (N_16081,N_14418,N_14095);
or U16082 (N_16082,N_15177,N_14458);
nor U16083 (N_16083,N_13047,N_12688);
and U16084 (N_16084,N_13488,N_14083);
nor U16085 (N_16085,N_15178,N_14257);
nor U16086 (N_16086,N_15105,N_14067);
nor U16087 (N_16087,N_14959,N_13779);
or U16088 (N_16088,N_14909,N_13063);
and U16089 (N_16089,N_13609,N_14566);
and U16090 (N_16090,N_14670,N_13414);
nor U16091 (N_16091,N_15035,N_13539);
nand U16092 (N_16092,N_13191,N_13630);
or U16093 (N_16093,N_15594,N_14936);
and U16094 (N_16094,N_13040,N_15219);
nand U16095 (N_16095,N_14850,N_14097);
nor U16096 (N_16096,N_15370,N_14339);
nor U16097 (N_16097,N_13104,N_14779);
nand U16098 (N_16098,N_12765,N_14102);
or U16099 (N_16099,N_12890,N_15268);
and U16100 (N_16100,N_12800,N_13457);
nor U16101 (N_16101,N_13628,N_14875);
nor U16102 (N_16102,N_12520,N_12575);
nor U16103 (N_16103,N_14581,N_15596);
nor U16104 (N_16104,N_13931,N_13940);
nor U16105 (N_16105,N_13052,N_12891);
or U16106 (N_16106,N_13453,N_12808);
or U16107 (N_16107,N_14849,N_13117);
nand U16108 (N_16108,N_13995,N_12860);
nand U16109 (N_16109,N_13087,N_14329);
or U16110 (N_16110,N_14881,N_14558);
nand U16111 (N_16111,N_14697,N_15580);
and U16112 (N_16112,N_15452,N_13125);
or U16113 (N_16113,N_14542,N_14319);
nor U16114 (N_16114,N_13064,N_13334);
and U16115 (N_16115,N_13333,N_14350);
or U16116 (N_16116,N_13489,N_14772);
or U16117 (N_16117,N_14718,N_14003);
nor U16118 (N_16118,N_14378,N_12802);
or U16119 (N_16119,N_12942,N_15211);
nand U16120 (N_16120,N_12732,N_15522);
nand U16121 (N_16121,N_13282,N_13567);
nor U16122 (N_16122,N_15529,N_14841);
nand U16123 (N_16123,N_14401,N_12921);
and U16124 (N_16124,N_14449,N_14946);
and U16125 (N_16125,N_14488,N_14379);
or U16126 (N_16126,N_13166,N_15507);
nand U16127 (N_16127,N_14262,N_14945);
nor U16128 (N_16128,N_13268,N_14574);
nor U16129 (N_16129,N_13934,N_14094);
or U16130 (N_16130,N_15602,N_13599);
nor U16131 (N_16131,N_13055,N_13206);
or U16132 (N_16132,N_13540,N_15621);
nand U16133 (N_16133,N_12996,N_13473);
and U16134 (N_16134,N_15231,N_13367);
nor U16135 (N_16135,N_14859,N_12920);
nand U16136 (N_16136,N_14352,N_13116);
or U16137 (N_16137,N_13354,N_14051);
xnor U16138 (N_16138,N_13384,N_12812);
and U16139 (N_16139,N_15327,N_14642);
and U16140 (N_16140,N_13468,N_14370);
nor U16141 (N_16141,N_12734,N_13677);
or U16142 (N_16142,N_13461,N_15418);
nor U16143 (N_16143,N_14283,N_14518);
or U16144 (N_16144,N_15022,N_15446);
or U16145 (N_16145,N_13532,N_14728);
nor U16146 (N_16146,N_13014,N_15456);
nand U16147 (N_16147,N_13161,N_13325);
nor U16148 (N_16148,N_13111,N_15165);
and U16149 (N_16149,N_12594,N_13069);
nor U16150 (N_16150,N_14467,N_12823);
nor U16151 (N_16151,N_12888,N_14689);
nor U16152 (N_16152,N_14867,N_14021);
nor U16153 (N_16153,N_14822,N_12769);
nor U16154 (N_16154,N_15465,N_12886);
or U16155 (N_16155,N_13623,N_12700);
nor U16156 (N_16156,N_15384,N_15500);
nor U16157 (N_16157,N_13766,N_12605);
nor U16158 (N_16158,N_12815,N_12589);
or U16159 (N_16159,N_14126,N_13697);
nor U16160 (N_16160,N_13696,N_12968);
and U16161 (N_16161,N_14958,N_15562);
and U16162 (N_16162,N_13932,N_13659);
nand U16163 (N_16163,N_15012,N_13838);
or U16164 (N_16164,N_14465,N_13880);
and U16165 (N_16165,N_14373,N_12795);
and U16166 (N_16166,N_13265,N_15274);
or U16167 (N_16167,N_15118,N_15425);
and U16168 (N_16168,N_15318,N_14342);
nand U16169 (N_16169,N_14663,N_14110);
and U16170 (N_16170,N_14315,N_15598);
nor U16171 (N_16171,N_14807,N_12910);
nor U16172 (N_16172,N_13221,N_14349);
nand U16173 (N_16173,N_14629,N_14321);
nand U16174 (N_16174,N_15188,N_13749);
and U16175 (N_16175,N_14421,N_13483);
xnor U16176 (N_16176,N_13810,N_13244);
and U16177 (N_16177,N_13433,N_12515);
nand U16178 (N_16178,N_15460,N_15382);
nand U16179 (N_16179,N_13921,N_14457);
nand U16180 (N_16180,N_14560,N_13989);
nor U16181 (N_16181,N_13708,N_12818);
nand U16182 (N_16182,N_14883,N_12714);
nand U16183 (N_16183,N_14205,N_14915);
nand U16184 (N_16184,N_13298,N_14897);
nor U16185 (N_16185,N_12639,N_14244);
nor U16186 (N_16186,N_13476,N_12887);
nor U16187 (N_16187,N_13222,N_14207);
and U16188 (N_16188,N_13392,N_14026);
nand U16189 (N_16189,N_14388,N_14249);
xnor U16190 (N_16190,N_13590,N_15175);
nand U16191 (N_16191,N_12913,N_14695);
and U16192 (N_16192,N_13229,N_14829);
nand U16193 (N_16193,N_12595,N_14864);
nand U16194 (N_16194,N_13913,N_14828);
nor U16195 (N_16195,N_15269,N_13740);
xnor U16196 (N_16196,N_14327,N_14515);
or U16197 (N_16197,N_15033,N_14533);
and U16198 (N_16198,N_14278,N_14197);
and U16199 (N_16199,N_15076,N_14775);
nand U16200 (N_16200,N_14128,N_14055);
and U16201 (N_16201,N_13143,N_15604);
or U16202 (N_16202,N_14154,N_13851);
xnor U16203 (N_16203,N_13092,N_14112);
and U16204 (N_16204,N_14403,N_13772);
nand U16205 (N_16205,N_15400,N_13563);
nor U16206 (N_16206,N_13050,N_13626);
or U16207 (N_16207,N_13017,N_15515);
and U16208 (N_16208,N_14429,N_14103);
nand U16209 (N_16209,N_15491,N_13097);
and U16210 (N_16210,N_13792,N_13372);
nand U16211 (N_16211,N_12833,N_12889);
nand U16212 (N_16212,N_12914,N_14027);
nand U16213 (N_16213,N_14392,N_12530);
nand U16214 (N_16214,N_15282,N_12874);
nor U16215 (N_16215,N_14456,N_13424);
or U16216 (N_16216,N_14993,N_12880);
nand U16217 (N_16217,N_14583,N_14042);
and U16218 (N_16218,N_12740,N_14645);
nand U16219 (N_16219,N_14662,N_15263);
and U16220 (N_16220,N_13119,N_12676);
or U16221 (N_16221,N_13856,N_13789);
and U16222 (N_16222,N_13585,N_13776);
xnor U16223 (N_16223,N_15374,N_12850);
nand U16224 (N_16224,N_15391,N_15044);
nand U16225 (N_16225,N_15494,N_14188);
nand U16226 (N_16226,N_13826,N_13970);
and U16227 (N_16227,N_13501,N_13393);
or U16228 (N_16228,N_14865,N_12756);
nand U16229 (N_16229,N_13927,N_13236);
nor U16230 (N_16230,N_12846,N_15498);
xnor U16231 (N_16231,N_15506,N_15011);
or U16232 (N_16232,N_15364,N_15333);
nand U16233 (N_16233,N_13110,N_14548);
and U16234 (N_16234,N_14423,N_14559);
and U16235 (N_16235,N_15077,N_15264);
nand U16236 (N_16236,N_13692,N_15169);
and U16237 (N_16237,N_12953,N_13335);
nand U16238 (N_16238,N_12727,N_14133);
xnor U16239 (N_16239,N_14272,N_14340);
xnor U16240 (N_16240,N_14932,N_13396);
or U16241 (N_16241,N_14832,N_13526);
and U16242 (N_16242,N_12997,N_14122);
nor U16243 (N_16243,N_13550,N_14121);
or U16244 (N_16244,N_13113,N_12971);
nand U16245 (N_16245,N_12801,N_13724);
nand U16246 (N_16246,N_13771,N_15385);
nor U16247 (N_16247,N_15523,N_15293);
nor U16248 (N_16248,N_12508,N_15336);
and U16249 (N_16249,N_12898,N_13112);
and U16250 (N_16250,N_14999,N_14202);
nand U16251 (N_16251,N_14140,N_14687);
or U16252 (N_16252,N_12518,N_13098);
or U16253 (N_16253,N_13132,N_12803);
and U16254 (N_16254,N_14351,N_13075);
and U16255 (N_16255,N_14118,N_13879);
and U16256 (N_16256,N_13562,N_14371);
xor U16257 (N_16257,N_13877,N_12504);
or U16258 (N_16258,N_12619,N_13993);
xnor U16259 (N_16259,N_12708,N_15002);
or U16260 (N_16260,N_15084,N_14322);
nand U16261 (N_16261,N_12757,N_15098);
nor U16262 (N_16262,N_13583,N_12566);
nand U16263 (N_16263,N_14504,N_14647);
nor U16264 (N_16264,N_13241,N_14738);
or U16265 (N_16265,N_14664,N_13058);
or U16266 (N_16266,N_14555,N_13962);
xnor U16267 (N_16267,N_12797,N_14693);
and U16268 (N_16268,N_15582,N_14887);
nor U16269 (N_16269,N_14671,N_14667);
or U16270 (N_16270,N_14151,N_14983);
nand U16271 (N_16271,N_13321,N_13728);
or U16272 (N_16272,N_13690,N_15095);
or U16273 (N_16273,N_13292,N_13067);
or U16274 (N_16274,N_14753,N_13958);
nor U16275 (N_16275,N_12701,N_14384);
and U16276 (N_16276,N_13770,N_12513);
nor U16277 (N_16277,N_13139,N_14537);
and U16278 (N_16278,N_15198,N_13209);
or U16279 (N_16279,N_14024,N_13670);
xnor U16280 (N_16280,N_14681,N_12631);
nor U16281 (N_16281,N_14037,N_13210);
nor U16282 (N_16282,N_15329,N_14393);
or U16283 (N_16283,N_14700,N_14234);
or U16284 (N_16284,N_13043,N_14782);
xnor U16285 (N_16285,N_12644,N_14890);
or U16286 (N_16286,N_14264,N_14888);
and U16287 (N_16287,N_14677,N_13464);
and U16288 (N_16288,N_13412,N_14527);
nor U16289 (N_16289,N_12528,N_13848);
or U16290 (N_16290,N_13657,N_14927);
nand U16291 (N_16291,N_13945,N_12840);
xor U16292 (N_16292,N_15102,N_13888);
nand U16293 (N_16293,N_13033,N_14263);
and U16294 (N_16294,N_13622,N_15081);
nor U16295 (N_16295,N_14620,N_14587);
and U16296 (N_16296,N_13975,N_12683);
or U16297 (N_16297,N_13175,N_12531);
nand U16298 (N_16298,N_13625,N_15623);
nor U16299 (N_16299,N_15530,N_15047);
or U16300 (N_16300,N_13303,N_13624);
or U16301 (N_16301,N_12563,N_14129);
or U16302 (N_16302,N_13686,N_14861);
and U16303 (N_16303,N_13324,N_13544);
nor U16304 (N_16304,N_15570,N_13785);
and U16305 (N_16305,N_12715,N_14093);
nand U16306 (N_16306,N_14271,N_15549);
nor U16307 (N_16307,N_12859,N_15228);
nor U16308 (N_16308,N_12779,N_13831);
and U16309 (N_16309,N_14686,N_12663);
xnor U16310 (N_16310,N_12919,N_14241);
or U16311 (N_16311,N_12782,N_13965);
or U16312 (N_16312,N_13754,N_13700);
nor U16313 (N_16313,N_13364,N_15350);
nand U16314 (N_16314,N_12784,N_12685);
or U16315 (N_16315,N_13320,N_12556);
xor U16316 (N_16316,N_13102,N_13237);
and U16317 (N_16317,N_12710,N_13712);
nand U16318 (N_16318,N_15006,N_13491);
and U16319 (N_16319,N_15140,N_13280);
nand U16320 (N_16320,N_14466,N_12783);
nor U16321 (N_16321,N_14131,N_15531);
or U16322 (N_16322,N_15469,N_13758);
or U16323 (N_16323,N_15034,N_12807);
and U16324 (N_16324,N_14521,N_13346);
nand U16325 (N_16325,N_12626,N_15064);
or U16326 (N_16326,N_15021,N_14211);
nor U16327 (N_16327,N_12680,N_15486);
xnor U16328 (N_16328,N_14982,N_14099);
xor U16329 (N_16329,N_15601,N_13256);
and U16330 (N_16330,N_12940,N_15273);
and U16331 (N_16331,N_13254,N_15069);
and U16332 (N_16332,N_15334,N_14800);
and U16333 (N_16333,N_15430,N_13462);
or U16334 (N_16334,N_14623,N_12851);
nand U16335 (N_16335,N_13828,N_14591);
and U16336 (N_16336,N_13949,N_13134);
nand U16337 (N_16337,N_13251,N_13881);
nand U16338 (N_16338,N_13832,N_13456);
nand U16339 (N_16339,N_15624,N_15597);
or U16340 (N_16340,N_15304,N_13759);
nand U16341 (N_16341,N_14672,N_14683);
nor U16342 (N_16342,N_15398,N_13301);
nand U16343 (N_16343,N_13034,N_14455);
nand U16344 (N_16344,N_13401,N_12822);
or U16345 (N_16345,N_13640,N_12609);
or U16346 (N_16346,N_15514,N_15277);
or U16347 (N_16347,N_13355,N_12798);
or U16348 (N_16348,N_14892,N_13639);
xnor U16349 (N_16349,N_12557,N_14990);
and U16350 (N_16350,N_15496,N_15616);
xnor U16351 (N_16351,N_14707,N_14929);
nor U16352 (N_16352,N_13155,N_13704);
xor U16353 (N_16353,N_15116,N_14496);
nor U16354 (N_16354,N_12827,N_15058);
nand U16355 (N_16355,N_14971,N_13036);
xnor U16356 (N_16356,N_15204,N_12820);
and U16357 (N_16357,N_13844,N_14577);
or U16358 (N_16358,N_15127,N_13373);
nor U16359 (N_16359,N_14528,N_15132);
xor U16360 (N_16360,N_12771,N_14411);
or U16361 (N_16361,N_12632,N_14290);
or U16362 (N_16362,N_14691,N_14367);
and U16363 (N_16363,N_13240,N_15472);
xor U16364 (N_16364,N_15236,N_12583);
and U16365 (N_16365,N_14028,N_13963);
nand U16366 (N_16366,N_14612,N_15533);
nand U16367 (N_16367,N_13006,N_12792);
and U16368 (N_16368,N_13118,N_14270);
nand U16369 (N_16369,N_14008,N_14793);
nand U16370 (N_16370,N_14502,N_13796);
and U16371 (N_16371,N_14218,N_15298);
nor U16372 (N_16372,N_12579,N_14412);
nor U16373 (N_16373,N_12703,N_15200);
nand U16374 (N_16374,N_14214,N_12533);
nand U16375 (N_16375,N_15036,N_13719);
or U16376 (N_16376,N_13170,N_13350);
nor U16377 (N_16377,N_13284,N_13340);
and U16378 (N_16378,N_14724,N_13073);
nand U16379 (N_16379,N_14077,N_13542);
or U16380 (N_16380,N_13310,N_14541);
and U16381 (N_16381,N_15341,N_13819);
or U16382 (N_16382,N_12752,N_14341);
and U16383 (N_16383,N_14565,N_13986);
and U16384 (N_16384,N_13644,N_13873);
and U16385 (N_16385,N_14299,N_12671);
xnor U16386 (N_16386,N_14684,N_15212);
nor U16387 (N_16387,N_14125,N_12599);
or U16388 (N_16388,N_13215,N_13248);
nor U16389 (N_16389,N_13745,N_14522);
or U16390 (N_16390,N_15167,N_15152);
nor U16391 (N_16391,N_14326,N_13602);
or U16392 (N_16392,N_13974,N_13031);
or U16393 (N_16393,N_14005,N_14608);
or U16394 (N_16394,N_15122,N_14006);
nor U16395 (N_16395,N_14692,N_13517);
or U16396 (N_16396,N_14089,N_12731);
and U16397 (N_16397,N_15561,N_15004);
or U16398 (N_16398,N_13269,N_14260);
and U16399 (N_16399,N_13560,N_13990);
or U16400 (N_16400,N_15031,N_14579);
nor U16401 (N_16401,N_13821,N_14834);
or U16402 (N_16402,N_15417,N_13279);
nor U16403 (N_16403,N_13028,N_13523);
nand U16404 (N_16404,N_12932,N_15324);
xor U16405 (N_16405,N_14957,N_13311);
nor U16406 (N_16406,N_13070,N_15234);
or U16407 (N_16407,N_15473,N_15357);
xor U16408 (N_16408,N_14935,N_14974);
or U16409 (N_16409,N_14106,N_13956);
or U16410 (N_16410,N_12662,N_12861);
xnor U16411 (N_16411,N_14385,N_13893);
nand U16412 (N_16412,N_14996,N_13936);
and U16413 (N_16413,N_14847,N_15048);
or U16414 (N_16414,N_14995,N_13889);
xor U16415 (N_16415,N_13568,N_15172);
nand U16416 (N_16416,N_14450,N_13614);
nand U16417 (N_16417,N_14148,N_14806);
xor U16418 (N_16418,N_13611,N_13985);
and U16419 (N_16419,N_12681,N_12722);
nand U16420 (N_16420,N_12697,N_12501);
xnor U16421 (N_16421,N_14941,N_14307);
and U16422 (N_16422,N_15346,N_12721);
or U16423 (N_16423,N_15023,N_12559);
nor U16424 (N_16424,N_15543,N_15476);
or U16425 (N_16425,N_15401,N_13223);
or U16426 (N_16426,N_15153,N_13144);
nor U16427 (N_16427,N_13416,N_13397);
or U16428 (N_16428,N_15259,N_15221);
nand U16429 (N_16429,N_13952,N_12829);
and U16430 (N_16430,N_14059,N_12746);
and U16431 (N_16431,N_14613,N_15289);
nor U16432 (N_16432,N_14827,N_13435);
nand U16433 (N_16433,N_13004,N_13564);
and U16434 (N_16434,N_14619,N_15088);
nor U16435 (N_16435,N_13091,N_12623);
nand U16436 (N_16436,N_15344,N_14709);
nor U16437 (N_16437,N_12545,N_13478);
or U16438 (N_16438,N_15414,N_14023);
and U16439 (N_16439,N_14719,N_15052);
and U16440 (N_16440,N_15256,N_12858);
nor U16441 (N_16441,N_12712,N_15242);
nand U16442 (N_16442,N_12775,N_13385);
or U16443 (N_16443,N_15136,N_13976);
nor U16444 (N_16444,N_13723,N_14166);
or U16445 (N_16445,N_13336,N_15424);
and U16446 (N_16446,N_14597,N_15008);
and U16447 (N_16447,N_15025,N_15017);
nand U16448 (N_16448,N_13981,N_14948);
and U16449 (N_16449,N_15458,N_13328);
or U16450 (N_16450,N_14404,N_15009);
xnor U16451 (N_16451,N_13777,N_15051);
or U16452 (N_16452,N_13850,N_12602);
and U16453 (N_16453,N_14919,N_12503);
nand U16454 (N_16454,N_13460,N_14863);
nand U16455 (N_16455,N_15365,N_13833);
xnor U16456 (N_16456,N_13820,N_15618);
and U16457 (N_16457,N_12972,N_14979);
or U16458 (N_16458,N_13318,N_14962);
nor U16459 (N_16459,N_13315,N_13480);
nor U16460 (N_16460,N_15024,N_15232);
nand U16461 (N_16461,N_13835,N_14033);
nand U16462 (N_16462,N_12655,N_14022);
and U16463 (N_16463,N_14543,N_13341);
xor U16464 (N_16464,N_14838,N_12580);
nor U16465 (N_16465,N_14938,N_14835);
nor U16466 (N_16466,N_15210,N_15342);
and U16467 (N_16467,N_15410,N_15248);
and U16468 (N_16468,N_12597,N_13582);
xor U16469 (N_16469,N_14550,N_14750);
nor U16470 (N_16470,N_12603,N_13613);
nand U16471 (N_16471,N_14433,N_14410);
or U16472 (N_16472,N_14804,N_12848);
or U16473 (N_16473,N_15470,N_13793);
or U16474 (N_16474,N_14756,N_14985);
nor U16475 (N_16475,N_14517,N_13538);
or U16476 (N_16476,N_13015,N_15255);
nor U16477 (N_16477,N_13718,N_13452);
nand U16478 (N_16478,N_15310,N_15620);
xnor U16479 (N_16479,N_14451,N_15487);
nor U16480 (N_16480,N_12675,N_14871);
nor U16481 (N_16481,N_13257,N_13589);
nand U16482 (N_16482,N_13636,N_15109);
and U16483 (N_16483,N_12669,N_13518);
and U16484 (N_16484,N_13549,N_12500);
nand U16485 (N_16485,N_14390,N_15450);
xnor U16486 (N_16486,N_14120,N_13472);
nor U16487 (N_16487,N_14187,N_14525);
xnor U16488 (N_16488,N_14650,N_14215);
nand U16489 (N_16489,N_12621,N_13194);
and U16490 (N_16490,N_12758,N_13744);
nor U16491 (N_16491,N_13099,N_12611);
xor U16492 (N_16492,N_15402,N_14599);
nor U16493 (N_16493,N_14997,N_15202);
xnor U16494 (N_16494,N_15107,N_15142);
nand U16495 (N_16495,N_15532,N_13451);
nand U16496 (N_16496,N_14576,N_15421);
nand U16497 (N_16497,N_14544,N_14731);
and U16498 (N_16498,N_13124,N_15207);
or U16499 (N_16499,N_13579,N_13953);
nor U16500 (N_16500,N_13887,N_14843);
and U16501 (N_16501,N_15309,N_13716);
nor U16502 (N_16502,N_14312,N_14748);
or U16503 (N_16503,N_15068,N_14947);
and U16504 (N_16504,N_12604,N_14749);
nand U16505 (N_16505,N_12747,N_13470);
or U16506 (N_16506,N_13016,N_15347);
and U16507 (N_16507,N_12906,N_13406);
and U16508 (N_16508,N_15266,N_15396);
nor U16509 (N_16509,N_14889,N_13260);
nor U16510 (N_16510,N_14531,N_14396);
or U16511 (N_16511,N_14666,N_15065);
or U16512 (N_16512,N_14261,N_12939);
and U16513 (N_16513,N_13249,N_15160);
nand U16514 (N_16514,N_13998,N_15015);
nor U16515 (N_16515,N_15201,N_12725);
and U16516 (N_16516,N_14269,N_14141);
nand U16517 (N_16517,N_13261,N_14175);
or U16518 (N_16518,N_13049,N_15437);
xnor U16519 (N_16519,N_14505,N_12720);
nand U16520 (N_16520,N_15086,N_15361);
nor U16521 (N_16521,N_12704,N_14726);
and U16522 (N_16522,N_13263,N_13297);
and U16523 (N_16523,N_14057,N_15173);
and U16524 (N_16524,N_12826,N_15573);
nand U16525 (N_16525,N_14593,N_15614);
or U16526 (N_16526,N_14831,N_15001);
nand U16527 (N_16527,N_13559,N_13533);
nor U16528 (N_16528,N_15571,N_15427);
and U16529 (N_16529,N_12630,N_15550);
nor U16530 (N_16530,N_13522,N_14852);
nor U16531 (N_16531,N_15591,N_14397);
xor U16532 (N_16532,N_13259,N_13186);
xor U16533 (N_16533,N_13870,N_12878);
nand U16534 (N_16534,N_14722,N_14711);
nor U16535 (N_16535,N_15191,N_12729);
nand U16536 (N_16536,N_13078,N_15174);
or U16537 (N_16537,N_14857,N_14354);
nand U16538 (N_16538,N_14618,N_14086);
and U16539 (N_16539,N_12660,N_13994);
xnor U16540 (N_16540,N_15511,N_14438);
and U16541 (N_16541,N_13799,N_14235);
and U16542 (N_16542,N_14858,N_14203);
and U16543 (N_16543,N_12835,N_14353);
and U16544 (N_16544,N_14124,N_15233);
xnor U16545 (N_16545,N_12749,N_15321);
and U16546 (N_16546,N_12863,N_13987);
xor U16547 (N_16547,N_13672,N_13753);
or U16548 (N_16548,N_12645,N_14899);
and U16549 (N_16549,N_13421,N_15488);
or U16550 (N_16550,N_12554,N_13020);
nand U16551 (N_16551,N_14553,N_13368);
nor U16552 (N_16552,N_15032,N_12805);
nand U16553 (N_16553,N_14640,N_15554);
xnor U16554 (N_16554,N_14096,N_15082);
nand U16555 (N_16555,N_12637,N_14812);
nand U16556 (N_16556,N_13039,N_13088);
or U16557 (N_16557,N_15540,N_14282);
or U16558 (N_16558,N_15288,N_12691);
nand U16559 (N_16559,N_14673,N_14563);
nor U16560 (N_16560,N_13158,N_14201);
nor U16561 (N_16561,N_14567,N_13197);
nand U16562 (N_16562,N_13922,N_13527);
and U16563 (N_16563,N_15599,N_15158);
xnor U16564 (N_16564,N_13982,N_15208);
xor U16565 (N_16565,N_13747,N_13891);
nand U16566 (N_16566,N_13190,N_14382);
nand U16567 (N_16567,N_13167,N_14325);
nand U16568 (N_16568,N_15583,N_12933);
nand U16569 (N_16569,N_13553,N_14237);
nor U16570 (N_16570,N_14074,N_15409);
nand U16571 (N_16571,N_14444,N_14343);
nor U16572 (N_16572,N_13653,N_15265);
nor U16573 (N_16573,N_13855,N_13830);
or U16574 (N_16574,N_13817,N_12610);
nand U16575 (N_16575,N_12711,N_15505);
xor U16576 (N_16576,N_13698,N_13788);
xnor U16577 (N_16577,N_15567,N_13216);
and U16578 (N_16578,N_13159,N_14727);
xnor U16579 (N_16579,N_13908,N_14923);
or U16580 (N_16580,N_13741,N_14632);
nor U16581 (N_16581,N_13005,N_13713);
or U16582 (N_16582,N_13171,N_14107);
or U16583 (N_16583,N_12760,N_14053);
and U16584 (N_16584,N_12952,N_14289);
and U16585 (N_16585,N_14280,N_13184);
nor U16586 (N_16586,N_15019,N_12999);
or U16587 (N_16587,N_12870,N_15375);
nand U16588 (N_16588,N_14150,N_14226);
or U16589 (N_16589,N_14961,N_14250);
and U16590 (N_16590,N_13943,N_13148);
xor U16591 (N_16591,N_13896,N_13405);
and U16592 (N_16592,N_13577,N_13919);
nand U16593 (N_16593,N_13575,N_12741);
nor U16594 (N_16594,N_14494,N_13029);
or U16595 (N_16595,N_14369,N_14258);
or U16596 (N_16596,N_13109,N_14248);
nor U16597 (N_16597,N_12917,N_13818);
nor U16598 (N_16598,N_15356,N_13715);
or U16599 (N_16599,N_12854,N_13105);
xnor U16600 (N_16600,N_13146,N_14869);
nor U16601 (N_16601,N_14153,N_12930);
and U16602 (N_16602,N_13695,N_14398);
nor U16603 (N_16603,N_14301,N_12923);
nor U16604 (N_16604,N_12995,N_15577);
xor U16605 (N_16605,N_14240,N_12811);
or U16606 (N_16606,N_12608,N_14885);
nor U16607 (N_16607,N_14601,N_14435);
and U16608 (N_16608,N_12916,N_13228);
nand U16609 (N_16609,N_12642,N_15609);
and U16610 (N_16610,N_15149,N_12677);
xnor U16611 (N_16611,N_12944,N_14479);
or U16612 (N_16612,N_14821,N_12540);
nand U16613 (N_16613,N_14309,N_13026);
nor U16614 (N_16614,N_14657,N_14955);
xnor U16615 (N_16615,N_14209,N_13366);
nor U16616 (N_16616,N_13314,N_14357);
nor U16617 (N_16617,N_13137,N_13574);
nor U16618 (N_16618,N_13773,N_15061);
nor U16619 (N_16619,N_15155,N_14611);
and U16620 (N_16620,N_15101,N_14845);
nand U16621 (N_16621,N_13122,N_14062);
or U16622 (N_16622,N_14098,N_13044);
or U16623 (N_16623,N_13054,N_13840);
or U16624 (N_16624,N_13090,N_14409);
nand U16625 (N_16625,N_14364,N_15131);
nand U16626 (N_16626,N_14781,N_12873);
nor U16627 (N_16627,N_12776,N_12546);
nor U16628 (N_16628,N_15525,N_13348);
nor U16629 (N_16629,N_13925,N_14602);
xnor U16630 (N_16630,N_13003,N_12793);
nor U16631 (N_16631,N_13768,N_15495);
and U16632 (N_16632,N_12643,N_14399);
and U16633 (N_16633,N_13235,N_13612);
nor U16634 (N_16634,N_14196,N_13323);
xnor U16635 (N_16635,N_15271,N_12900);
or U16636 (N_16636,N_15566,N_14774);
or U16637 (N_16637,N_12857,N_13621);
nand U16638 (N_16638,N_15043,N_14918);
xor U16639 (N_16639,N_13895,N_14520);
xnor U16640 (N_16640,N_14000,N_14910);
nand U16641 (N_16641,N_14562,N_14079);
or U16642 (N_16642,N_15018,N_15555);
nand U16643 (N_16643,N_14661,N_13082);
nor U16644 (N_16644,N_13332,N_15270);
nor U16645 (N_16645,N_13682,N_13829);
nand U16646 (N_16646,N_15559,N_13535);
nor U16647 (N_16647,N_12937,N_13591);
nand U16648 (N_16648,N_13580,N_14872);
nand U16649 (N_16649,N_14491,N_12967);
nand U16650 (N_16650,N_15297,N_13278);
xnor U16651 (N_16651,N_15138,N_14715);
and U16652 (N_16652,N_12562,N_13357);
xor U16653 (N_16653,N_14394,N_15617);
or U16654 (N_16654,N_15369,N_13862);
xor U16655 (N_16655,N_14346,N_14294);
or U16656 (N_16656,N_14736,N_14212);
or U16657 (N_16657,N_14189,N_13059);
or U16658 (N_16658,N_15206,N_13878);
and U16659 (N_16659,N_13702,N_12636);
nor U16660 (N_16660,N_15027,N_14284);
and U16661 (N_16661,N_15433,N_12766);
nand U16662 (N_16662,N_12558,N_12547);
or U16663 (N_16663,N_12915,N_13352);
nand U16664 (N_16664,N_12925,N_14705);
nor U16665 (N_16665,N_14300,N_13693);
and U16666 (N_16666,N_12744,N_13543);
or U16667 (N_16667,N_14176,N_13450);
xor U16668 (N_16668,N_15354,N_14625);
nor U16669 (N_16669,N_13930,N_12526);
nand U16670 (N_16670,N_13498,N_12622);
or U16671 (N_16671,N_14204,N_13239);
or U16672 (N_16672,N_14760,N_13147);
or U16673 (N_16673,N_14884,N_14012);
xor U16674 (N_16674,N_13162,N_14306);
and U16675 (N_16675,N_14758,N_14267);
or U16676 (N_16676,N_15563,N_14506);
and U16677 (N_16677,N_14819,N_15394);
nand U16678 (N_16678,N_12973,N_15120);
and U16679 (N_16679,N_15492,N_13992);
nor U16680 (N_16680,N_14061,N_15335);
and U16681 (N_16681,N_15134,N_14786);
or U16682 (N_16682,N_14987,N_14183);
and U16683 (N_16683,N_15358,N_13426);
nand U16684 (N_16684,N_14090,N_13449);
nor U16685 (N_16685,N_14519,N_12696);
and U16686 (N_16686,N_12667,N_12899);
nand U16687 (N_16687,N_14713,N_15479);
or U16688 (N_16688,N_14763,N_12806);
nand U16689 (N_16689,N_12745,N_13951);
nor U16690 (N_16690,N_14714,N_13680);
or U16691 (N_16691,N_13018,N_12987);
nand U16692 (N_16692,N_12901,N_13794);
and U16693 (N_16693,N_14056,N_14402);
xnor U16694 (N_16694,N_12565,N_14764);
or U16695 (N_16695,N_13646,N_13360);
nor U16696 (N_16696,N_13739,N_14803);
nand U16697 (N_16697,N_15294,N_14817);
xnor U16698 (N_16698,N_15311,N_12668);
nor U16699 (N_16699,N_15314,N_13032);
or U16700 (N_16700,N_13296,N_14610);
and U16701 (N_16701,N_13145,N_14413);
nor U16702 (N_16702,N_13446,N_14114);
nor U16703 (N_16703,N_14408,N_13347);
nor U16704 (N_16704,N_14922,N_15146);
xnor U16705 (N_16705,N_13699,N_13141);
and U16706 (N_16706,N_15471,N_13400);
and U16707 (N_16707,N_12905,N_15330);
and U16708 (N_16708,N_13816,N_13481);
nor U16709 (N_16709,N_14757,N_14359);
nor U16710 (N_16710,N_14191,N_14181);
xnor U16711 (N_16711,N_13961,N_12673);
or U16712 (N_16712,N_13929,N_14295);
nor U16713 (N_16713,N_14630,N_15038);
and U16714 (N_16714,N_14320,N_12912);
and U16715 (N_16715,N_15141,N_14638);
nor U16716 (N_16716,N_13183,N_14473);
or U16717 (N_16717,N_12841,N_13150);
and U16718 (N_16718,N_14031,N_13441);
nor U16719 (N_16719,N_14422,N_13955);
nand U16720 (N_16720,N_12788,N_12666);
nand U16721 (N_16721,N_15054,N_12767);
or U16722 (N_16722,N_14017,N_13220);
or U16723 (N_16723,N_14720,N_14510);
nor U16724 (N_16724,N_15305,N_13634);
nand U16725 (N_16725,N_14108,N_14085);
or U16726 (N_16726,N_14462,N_13080);
and U16727 (N_16727,N_13010,N_13746);
nand U16728 (N_16728,N_14767,N_14344);
or U16729 (N_16729,N_14192,N_15392);
nor U16730 (N_16730,N_15067,N_15395);
nor U16731 (N_16731,N_13007,N_14414);
nor U16732 (N_16732,N_13247,N_14799);
xor U16733 (N_16733,N_13557,N_13189);
xnor U16734 (N_16734,N_15053,N_15129);
or U16735 (N_16735,N_14446,N_12733);
nor U16736 (N_16736,N_15517,N_13329);
nor U16737 (N_16737,N_14538,N_14866);
nor U16738 (N_16738,N_13627,N_12961);
nand U16739 (N_16739,N_14879,N_13085);
xnor U16740 (N_16740,N_14584,N_15608);
nor U16741 (N_16741,N_13606,N_12872);
nor U16742 (N_16742,N_14011,N_15521);
nor U16743 (N_16743,N_15464,N_13783);
xor U16744 (N_16744,N_14049,N_13650);
and U16745 (N_16745,N_12786,N_12907);
nor U16746 (N_16746,N_13972,N_14047);
or U16747 (N_16747,N_12627,N_15454);
nand U16748 (N_16748,N_13656,N_12954);
and U16749 (N_16749,N_13769,N_13852);
or U16750 (N_16750,N_14674,N_13344);
nor U16751 (N_16751,N_14158,N_15066);
nand U16752 (N_16752,N_13074,N_13631);
and U16753 (N_16753,N_13418,N_15557);
nor U16754 (N_16754,N_12529,N_14972);
nand U16755 (N_16755,N_15130,N_15247);
or U16756 (N_16756,N_14908,N_15258);
nor U16757 (N_16757,N_12948,N_15091);
or U16758 (N_16758,N_14604,N_15343);
and U16759 (N_16759,N_12778,N_13283);
nor U16760 (N_16760,N_12977,N_12844);
or U16761 (N_16761,N_13174,N_13300);
nand U16762 (N_16762,N_14498,N_12534);
nand U16763 (N_16763,N_13486,N_13685);
or U16764 (N_16764,N_13270,N_14977);
xnor U16765 (N_16765,N_13926,N_13234);
or U16766 (N_16766,N_14816,N_15184);
and U16767 (N_16767,N_13966,N_14165);
nand U16768 (N_16768,N_14030,N_15605);
nand U16769 (N_16769,N_14530,N_12672);
and U16770 (N_16770,N_13991,N_13427);
or U16771 (N_16771,N_12838,N_13439);
nand U16772 (N_16772,N_12571,N_13381);
nor U16773 (N_16773,N_12502,N_15581);
or U16774 (N_16774,N_13814,N_14605);
and U16775 (N_16775,N_15474,N_15504);
or U16776 (N_16776,N_13061,N_15114);
or U16777 (N_16777,N_12947,N_14991);
and U16778 (N_16778,N_15192,N_14900);
and U16779 (N_16779,N_15176,N_14084);
nand U16780 (N_16780,N_14598,N_13954);
nor U16781 (N_16781,N_12550,N_14360);
and U16782 (N_16782,N_12902,N_13205);
and U16783 (N_16783,N_13008,N_12885);
nand U16784 (N_16784,N_14805,N_14614);
nor U16785 (N_16785,N_13632,N_14497);
and U16786 (N_16786,N_14453,N_12804);
nor U16787 (N_16787,N_13019,N_15428);
and U16788 (N_16788,N_14472,N_13664);
and U16789 (N_16789,N_15489,N_14644);
or U16790 (N_16790,N_14624,N_14043);
or U16791 (N_16791,N_13823,N_12983);
nor U16792 (N_16792,N_14437,N_15085);
and U16793 (N_16793,N_15397,N_13558);
nor U16794 (N_16794,N_14276,N_13129);
nor U16795 (N_16795,N_12931,N_15145);
nand U16796 (N_16796,N_14232,N_13035);
nand U16797 (N_16797,N_15411,N_12523);
and U16798 (N_16798,N_12781,N_12724);
xor U16799 (N_16799,N_15112,N_14572);
and U16800 (N_16800,N_14949,N_13778);
xor U16801 (N_16801,N_13675,N_12791);
or U16802 (N_16802,N_14658,N_14231);
xnor U16803 (N_16803,N_14220,N_13516);
and U16804 (N_16804,N_15278,N_12635);
nand U16805 (N_16805,N_14511,N_12828);
or U16806 (N_16806,N_14277,N_15574);
and U16807 (N_16807,N_15331,N_14144);
nor U16808 (N_16808,N_13511,N_13121);
nor U16809 (N_16809,N_15560,N_14998);
nor U16810 (N_16810,N_14333,N_13056);
nand U16811 (N_16811,N_14824,N_13025);
and U16812 (N_16812,N_13169,N_13801);
nor U16813 (N_16813,N_13390,N_13076);
or U16814 (N_16814,N_13180,N_14796);
nand U16815 (N_16815,N_14626,N_14075);
nor U16816 (N_16816,N_13255,N_13534);
or U16817 (N_16817,N_14943,N_14480);
and U16818 (N_16818,N_12950,N_13581);
xor U16819 (N_16819,N_13163,N_13545);
nor U16820 (N_16820,N_12825,N_12754);
nor U16821 (N_16821,N_13548,N_13081);
nor U16822 (N_16822,N_15166,N_14902);
nor U16823 (N_16823,N_14474,N_13761);
nor U16824 (N_16824,N_14275,N_15462);
nor U16825 (N_16825,N_14712,N_14837);
nor U16826 (N_16826,N_13030,N_14571);
nand U16827 (N_16827,N_13933,N_12719);
or U16828 (N_16828,N_13101,N_13757);
or U16829 (N_16829,N_12650,N_13598);
or U16830 (N_16830,N_14172,N_14452);
and U16831 (N_16831,N_14044,N_15213);
and U16832 (N_16832,N_14223,N_14696);
and U16833 (N_16833,N_13641,N_15548);
or U16834 (N_16834,N_15475,N_15144);
nand U16835 (N_16835,N_14025,N_15197);
nor U16836 (N_16836,N_15135,N_14174);
nand U16837 (N_16837,N_15060,N_13276);
and U16838 (N_16838,N_14891,N_14149);
nand U16839 (N_16839,N_12539,N_15480);
xor U16840 (N_16840,N_14622,N_13138);
and U16841 (N_16841,N_12750,N_12834);
nor U16842 (N_16842,N_12908,N_14487);
nand U16843 (N_16843,N_13843,N_13437);
xor U16844 (N_16844,N_13062,N_14508);
xnor U16845 (N_16845,N_12969,N_14596);
nor U16846 (N_16846,N_13720,N_13944);
and U16847 (N_16847,N_14245,N_15280);
and U16848 (N_16848,N_12774,N_14143);
xor U16849 (N_16849,N_15209,N_14877);
and U16850 (N_16850,N_15189,N_14014);
nor U16851 (N_16851,N_13825,N_15449);
and U16852 (N_16852,N_14041,N_15576);
or U16853 (N_16853,N_15251,N_14233);
and U16854 (N_16854,N_12544,N_12770);
and U16855 (N_16855,N_14651,N_13432);
and U16856 (N_16856,N_15170,N_12572);
xnor U16857 (N_16857,N_12865,N_14759);
nand U16858 (N_16858,N_14818,N_15351);
nor U16859 (N_16859,N_14792,N_14896);
nor U16860 (N_16860,N_12946,N_15412);
nand U16861 (N_16861,N_15124,N_14787);
or U16862 (N_16862,N_15113,N_12514);
and U16863 (N_16863,N_14463,N_14224);
and U16864 (N_16864,N_14953,N_14222);
or U16865 (N_16865,N_12787,N_13151);
nor U16866 (N_16866,N_14701,N_14814);
nor U16867 (N_16867,N_15254,N_13287);
and U16868 (N_16868,N_12532,N_15613);
and U16869 (N_16869,N_14273,N_14256);
nand U16870 (N_16870,N_13663,N_14015);
nor U16871 (N_16871,N_14870,N_14575);
or U16872 (N_16872,N_14901,N_15388);
or U16873 (N_16873,N_14680,N_14328);
or U16874 (N_16874,N_13667,N_13200);
nand U16875 (N_16875,N_13475,N_14375);
or U16876 (N_16876,N_15447,N_13996);
nor U16877 (N_16877,N_14986,N_12868);
nor U16878 (N_16878,N_13867,N_13442);
nand U16879 (N_16879,N_15121,N_13152);
xnor U16880 (N_16880,N_14302,N_14755);
and U16881 (N_16881,N_13262,N_13620);
nand U16882 (N_16882,N_14925,N_14876);
or U16883 (N_16883,N_15281,N_14634);
nor U16884 (N_16884,N_13918,N_12867);
xor U16885 (N_16885,N_13762,N_14994);
and U16886 (N_16886,N_13245,N_15313);
nor U16887 (N_16887,N_13824,N_12839);
nor U16888 (N_16888,N_13013,N_13302);
or U16889 (N_16889,N_13369,N_14840);
and U16890 (N_16890,N_13142,N_14168);
nand U16891 (N_16891,N_13726,N_15516);
and U16892 (N_16892,N_13207,N_13140);
and U16893 (N_16893,N_15612,N_14331);
and U16894 (N_16894,N_15163,N_14660);
xor U16895 (N_16895,N_14356,N_14318);
or U16896 (N_16896,N_14500,N_12682);
and U16897 (N_16897,N_13380,N_12674);
nor U16898 (N_16898,N_14554,N_14279);
nand U16899 (N_16899,N_14391,N_13399);
nor U16900 (N_16900,N_13471,N_13275);
and U16901 (N_16901,N_13288,N_12505);
nor U16902 (N_16902,N_14495,N_14648);
nand U16903 (N_16903,N_15240,N_13115);
or U16904 (N_16904,N_13709,N_15013);
or U16905 (N_16905,N_13578,N_14266);
or U16906 (N_16906,N_15610,N_14802);
and U16907 (N_16907,N_12927,N_15607);
nor U16908 (N_16908,N_13485,N_13173);
nor U16909 (N_16909,N_13865,N_15291);
and U16910 (N_16910,N_15093,N_13643);
and U16911 (N_16911,N_13964,N_13547);
or U16912 (N_16912,N_14529,N_12535);
or U16913 (N_16913,N_15253,N_12742);
nor U16914 (N_16914,N_12882,N_14255);
and U16915 (N_16915,N_12982,N_13797);
and U16916 (N_16916,N_13592,N_13756);
nor U16917 (N_16917,N_13676,N_13499);
and U16918 (N_16918,N_15046,N_13496);
and U16919 (N_16919,N_13168,N_14839);
or U16920 (N_16920,N_12651,N_12706);
and U16921 (N_16921,N_14313,N_15455);
nor U16922 (N_16922,N_14535,N_14469);
or U16923 (N_16923,N_15193,N_13999);
nand U16924 (N_16924,N_13635,N_15185);
or U16925 (N_16925,N_14690,N_13941);
nand U16926 (N_16926,N_13546,N_12957);
and U16927 (N_16927,N_15147,N_13041);
or U16928 (N_16928,N_15390,N_12654);
and U16929 (N_16929,N_13633,N_13185);
and U16930 (N_16930,N_12869,N_14137);
or U16931 (N_16931,N_14383,N_13897);
and U16932 (N_16932,N_12692,N_12790);
or U16933 (N_16933,N_15301,N_15262);
and U16934 (N_16934,N_15239,N_13120);
and U16935 (N_16935,N_14039,N_12616);
nor U16936 (N_16936,N_15322,N_12831);
nand U16937 (N_16937,N_14287,N_14740);
nand U16938 (N_16938,N_13600,N_13389);
xor U16939 (N_16939,N_12763,N_13065);
or U16940 (N_16940,N_13425,N_13130);
nand U16941 (N_16941,N_14628,N_14101);
and U16942 (N_16942,N_15526,N_15429);
or U16943 (N_16943,N_12573,N_13886);
nor U16944 (N_16944,N_12959,N_14721);
and U16945 (N_16945,N_14216,N_12612);
nand U16946 (N_16946,N_15286,N_14441);
nor U16947 (N_16947,N_14001,N_14251);
or U16948 (N_16948,N_13780,N_14723);
xor U16949 (N_16949,N_13671,N_15199);
nor U16950 (N_16950,N_15553,N_13444);
nor U16951 (N_16951,N_14230,N_15406);
or U16952 (N_16952,N_14668,N_13786);
nand U16953 (N_16953,N_14960,N_14744);
nand U16954 (N_16954,N_14381,N_13979);
or U16955 (N_16955,N_14968,N_13775);
nand U16956 (N_16956,N_15227,N_14969);
xor U16957 (N_16957,N_13730,N_15518);
or U16958 (N_16958,N_14678,N_12590);
or U16959 (N_16959,N_13000,N_13901);
and U16960 (N_16960,N_13935,N_13127);
and U16961 (N_16961,N_15039,N_14860);
xor U16962 (N_16962,N_13681,N_14136);
nor U16963 (N_16963,N_13811,N_15137);
nand U16964 (N_16964,N_15373,N_12601);
nand U16965 (N_16965,N_14778,N_13588);
or U16966 (N_16966,N_13973,N_14513);
and U16967 (N_16967,N_13910,N_13411);
and U16968 (N_16968,N_14358,N_14050);
xor U16969 (N_16969,N_15317,N_15434);
nor U16970 (N_16970,N_14180,N_14856);
nand U16971 (N_16971,N_12736,N_15348);
and U16972 (N_16972,N_13977,N_15389);
and U16973 (N_16973,N_13327,N_12687);
and U16974 (N_16974,N_13042,N_12726);
nand U16975 (N_16975,N_14020,N_15499);
nand U16976 (N_16976,N_14161,N_15407);
and U16977 (N_16977,N_15257,N_13417);
and U16978 (N_16978,N_15241,N_14155);
or U16979 (N_16979,N_14967,N_15451);
nand U16980 (N_16980,N_15545,N_13126);
nor U16981 (N_16981,N_13948,N_14717);
nor U16982 (N_16982,N_13108,N_12772);
nand U16983 (N_16983,N_13947,N_14145);
nand U16984 (N_16984,N_13365,N_13305);
nand U16985 (N_16985,N_14826,N_15063);
nand U16986 (N_16986,N_15154,N_13309);
nand U16987 (N_16987,N_13423,N_15151);
nor U16988 (N_16988,N_14665,N_13727);
nand U16989 (N_16989,N_13971,N_14239);
or U16990 (N_16990,N_14336,N_13312);
nand U16991 (N_16991,N_14163,N_13408);
or U16992 (N_16992,N_15037,N_14489);
nand U16993 (N_16993,N_13243,N_14228);
or U16994 (N_16994,N_13764,N_13371);
nor U16995 (N_16995,N_13573,N_15485);
or U16996 (N_16996,N_12638,N_15461);
nand U16997 (N_16997,N_13497,N_12981);
and U16998 (N_16998,N_14704,N_14281);
or U16999 (N_16999,N_14069,N_14509);
xor U17000 (N_17000,N_13655,N_13968);
or U17001 (N_17001,N_12509,N_12965);
nor U17002 (N_17002,N_13846,N_13688);
and U17003 (N_17003,N_14815,N_13233);
nor U17004 (N_17004,N_14746,N_14288);
nand U17005 (N_17005,N_13984,N_14637);
nand U17006 (N_17006,N_14470,N_12510);
nand U17007 (N_17007,N_14766,N_14298);
and U17008 (N_17008,N_13760,N_12536);
and U17009 (N_17009,N_13509,N_12809);
or U17010 (N_17010,N_12945,N_13440);
and U17011 (N_17011,N_13513,N_12738);
and U17012 (N_17012,N_13647,N_15615);
or U17013 (N_17013,N_12970,N_12871);
nand U17014 (N_17014,N_13597,N_13479);
nor U17015 (N_17015,N_13717,N_15162);
or U17016 (N_17016,N_14855,N_14311);
and U17017 (N_17017,N_12852,N_15466);
nand U17018 (N_17018,N_13555,N_13388);
nor U17019 (N_17019,N_13587,N_14238);
or U17020 (N_17020,N_13969,N_13253);
nand U17021 (N_17021,N_13394,N_12894);
and U17022 (N_17022,N_13669,N_12694);
and U17023 (N_17023,N_12814,N_14104);
xnor U17024 (N_17024,N_13900,N_15111);
or U17025 (N_17025,N_14493,N_14464);
nor U17026 (N_17026,N_13572,N_13800);
nand U17027 (N_17027,N_15381,N_14809);
or U17028 (N_17028,N_13226,N_13250);
nor U17029 (N_17029,N_15000,N_14616);
nand U17030 (N_17030,N_14190,N_14825);
nand U17031 (N_17031,N_14486,N_14407);
and U17032 (N_17032,N_13503,N_14117);
and U17033 (N_17033,N_12625,N_15509);
nand U17034 (N_17034,N_14010,N_15320);
or U17035 (N_17035,N_14135,N_14777);
nor U17036 (N_17036,N_15393,N_14580);
nand U17037 (N_17037,N_14984,N_14310);
nor U17038 (N_17038,N_13267,N_13495);
or U17039 (N_17039,N_15080,N_13957);
or U17040 (N_17040,N_13131,N_13469);
or U17041 (N_17041,N_13266,N_15125);
nor U17042 (N_17042,N_12664,N_12702);
or U17043 (N_17043,N_15090,N_13554);
xor U17044 (N_17044,N_12794,N_13359);
or U17045 (N_17045,N_15459,N_14655);
nor U17046 (N_17046,N_15214,N_14111);
or U17047 (N_17047,N_12564,N_14246);
nor U17048 (N_17048,N_12567,N_13156);
nor U17049 (N_17049,N_12978,N_12519);
or U17050 (N_17050,N_12780,N_15300);
xor U17051 (N_17051,N_13571,N_14921);
nor U17052 (N_17052,N_13668,N_15092);
nor U17053 (N_17053,N_15283,N_13319);
nor U17054 (N_17054,N_14087,N_15481);
and U17055 (N_17055,N_12926,N_13735);
nand U17056 (N_17056,N_13679,N_13556);
or U17057 (N_17057,N_14314,N_15078);
and U17058 (N_17058,N_13214,N_13195);
nand U17059 (N_17059,N_13528,N_13861);
nand U17060 (N_17060,N_14142,N_14906);
or U17061 (N_17061,N_14769,N_14635);
nor U17062 (N_17062,N_15368,N_12640);
nor U17063 (N_17063,N_13884,N_15171);
or U17064 (N_17064,N_14813,N_14823);
nand U17065 (N_17065,N_13707,N_13199);
and U17066 (N_17066,N_13841,N_13349);
nor U17067 (N_17067,N_12705,N_15328);
and U17068 (N_17068,N_13504,N_13454);
nand U17069 (N_17069,N_15089,N_15353);
and U17070 (N_17070,N_13317,N_15284);
and U17071 (N_17071,N_14400,N_15383);
nand U17072 (N_17072,N_14729,N_13658);
nor U17073 (N_17073,N_13386,N_13038);
and U17074 (N_17074,N_14436,N_14933);
and U17075 (N_17075,N_15075,N_12641);
and U17076 (N_17076,N_14330,N_14742);
or U17077 (N_17077,N_14675,N_12837);
and U17078 (N_17078,N_13490,N_12755);
and U17079 (N_17079,N_13445,N_13629);
or U17080 (N_17080,N_15513,N_14063);
nand U17081 (N_17081,N_15143,N_14268);
nand U17082 (N_17082,N_14708,N_13024);
nor U17083 (N_17083,N_15422,N_13339);
or U17084 (N_17084,N_13842,N_13182);
nand U17085 (N_17085,N_15546,N_13674);
nand U17086 (N_17086,N_13857,N_13684);
nand U17087 (N_17087,N_13923,N_13808);
or U17088 (N_17088,N_13383,N_12578);
nand U17089 (N_17089,N_13660,N_15386);
and U17090 (N_17090,N_13271,N_14389);
or U17091 (N_17091,N_13289,N_14526);
and U17092 (N_17092,N_13566,N_14316);
nor U17093 (N_17093,N_13051,N_13351);
and U17094 (N_17094,N_13407,N_15590);
nand U17095 (N_17095,N_15592,N_14873);
nand U17096 (N_17096,N_14184,N_12730);
nor U17097 (N_17097,N_14652,N_15319);
and U17098 (N_17098,N_12570,N_15611);
nand U17099 (N_17099,N_12522,N_14944);
nand U17100 (N_17100,N_14732,N_15203);
nor U17101 (N_17101,N_14119,N_14109);
nand U17102 (N_17102,N_15535,N_14338);
or U17103 (N_17103,N_14679,N_13313);
and U17104 (N_17104,N_13374,N_14649);
nand U17105 (N_17105,N_15326,N_14332);
or U17106 (N_17106,N_15568,N_14589);
nand U17107 (N_17107,N_13863,N_15115);
or U17108 (N_17108,N_14615,N_13285);
nor U17109 (N_17109,N_13584,N_14578);
nor U17110 (N_17110,N_15503,N_12764);
nand U17111 (N_17111,N_14146,N_12785);
or U17112 (N_17112,N_14115,N_13822);
nand U17113 (N_17113,N_15187,N_14492);
and U17114 (N_17114,N_14478,N_15519);
or U17115 (N_17115,N_13767,N_13791);
xnor U17116 (N_17116,N_13618,N_13027);
xor U17117 (N_17117,N_14170,N_14569);
xnor U17118 (N_17118,N_13839,N_13845);
nand U17119 (N_17119,N_15220,N_13596);
nor U17120 (N_17120,N_13387,N_14988);
or U17121 (N_17121,N_15272,N_13616);
and U17122 (N_17122,N_14912,N_14846);
nand U17123 (N_17123,N_15126,N_12992);
nor U17124 (N_17124,N_12761,N_12569);
nor U17125 (N_17125,N_13722,N_14009);
nand U17126 (N_17126,N_15205,N_14476);
or U17127 (N_17127,N_13316,N_13037);
or U17128 (N_17128,N_14032,N_12875);
or U17129 (N_17129,N_15312,N_12652);
or U17130 (N_17130,N_12986,N_15403);
and U17131 (N_17131,N_14092,N_13294);
or U17132 (N_17132,N_14225,N_15420);
nand U17133 (N_17133,N_14171,N_14105);
nor U17134 (N_17134,N_13009,N_14874);
nand U17135 (N_17135,N_13277,N_13924);
nor U17136 (N_17136,N_12994,N_13286);
nand U17137 (N_17137,N_15005,N_13290);
nand U17138 (N_17138,N_13345,N_13079);
nor U17139 (N_17139,N_15161,N_14265);
or U17140 (N_17140,N_14178,N_12893);
or U17141 (N_17141,N_14048,N_13849);
or U17142 (N_17142,N_14699,N_13859);
or U17143 (N_17143,N_12600,N_13187);
or U17144 (N_17144,N_13370,N_13404);
or U17145 (N_17145,N_13755,N_15366);
xor U17146 (N_17146,N_12743,N_14123);
or U17147 (N_17147,N_14931,N_14293);
and U17148 (N_17148,N_13916,N_13804);
or U17149 (N_17149,N_13225,N_13997);
and U17150 (N_17150,N_14833,N_13391);
nor U17151 (N_17151,N_15222,N_15307);
or U17152 (N_17152,N_14173,N_15295);
and U17153 (N_17153,N_13514,N_13428);
xor U17154 (N_17154,N_14973,N_14551);
and U17155 (N_17155,N_14688,N_12955);
or U17156 (N_17156,N_12551,N_14621);
or U17157 (N_17157,N_14362,N_13752);
nor U17158 (N_17158,N_13787,N_15527);
or U17159 (N_17159,N_13429,N_14523);
xnor U17160 (N_17160,N_15435,N_13330);
xor U17161 (N_17161,N_13203,N_15352);
xnor U17162 (N_17162,N_12561,N_15062);
nor U17163 (N_17163,N_15593,N_13322);
or U17164 (N_17164,N_14534,N_13876);
nand U17165 (N_17165,N_15119,N_15087);
nand U17166 (N_17166,N_15445,N_14532);
nand U17167 (N_17167,N_14880,N_14169);
or U17168 (N_17168,N_15148,N_12984);
nor U17169 (N_17169,N_15528,N_14797);
and U17170 (N_17170,N_15157,N_14078);
nand U17171 (N_17171,N_13904,N_14780);
nand U17172 (N_17172,N_15299,N_15133);
nor U17173 (N_17173,N_15016,N_12881);
nand U17174 (N_17174,N_15303,N_15186);
xor U17175 (N_17175,N_15586,N_15579);
or U17176 (N_17176,N_14317,N_13525);
xor U17177 (N_17177,N_13246,N_15380);
or U17178 (N_17178,N_12911,N_14468);
nand U17179 (N_17179,N_14484,N_15524);
or U17180 (N_17180,N_14951,N_12918);
nand U17181 (N_17181,N_14725,N_14501);
and U17182 (N_17182,N_14669,N_14454);
nor U17183 (N_17183,N_15440,N_13898);
nand U17184 (N_17184,N_15355,N_15050);
or U17185 (N_17185,N_14477,N_14132);
or U17186 (N_17186,N_13603,N_13960);
nor U17187 (N_17187,N_14499,N_12823);
and U17188 (N_17188,N_15390,N_13129);
nor U17189 (N_17189,N_15227,N_15225);
nand U17190 (N_17190,N_15553,N_14329);
nand U17191 (N_17191,N_13037,N_14876);
and U17192 (N_17192,N_14691,N_13163);
nor U17193 (N_17193,N_15340,N_13017);
and U17194 (N_17194,N_13701,N_14848);
or U17195 (N_17195,N_13425,N_14763);
or U17196 (N_17196,N_15015,N_12680);
xor U17197 (N_17197,N_14239,N_13427);
and U17198 (N_17198,N_14924,N_13148);
and U17199 (N_17199,N_13942,N_14921);
nand U17200 (N_17200,N_14999,N_13056);
and U17201 (N_17201,N_13161,N_14338);
and U17202 (N_17202,N_15555,N_14021);
and U17203 (N_17203,N_12929,N_13852);
and U17204 (N_17204,N_13025,N_13391);
and U17205 (N_17205,N_12843,N_15465);
nand U17206 (N_17206,N_14671,N_13535);
and U17207 (N_17207,N_12815,N_12527);
or U17208 (N_17208,N_15264,N_15527);
or U17209 (N_17209,N_12780,N_14354);
and U17210 (N_17210,N_14023,N_13450);
nand U17211 (N_17211,N_13690,N_14717);
xor U17212 (N_17212,N_15174,N_14076);
nor U17213 (N_17213,N_12591,N_15424);
xor U17214 (N_17214,N_12744,N_12832);
nand U17215 (N_17215,N_12763,N_15425);
or U17216 (N_17216,N_12531,N_12861);
and U17217 (N_17217,N_13681,N_12729);
nand U17218 (N_17218,N_15205,N_13285);
nand U17219 (N_17219,N_12673,N_13872);
and U17220 (N_17220,N_15432,N_15042);
or U17221 (N_17221,N_14168,N_14005);
or U17222 (N_17222,N_12741,N_13382);
or U17223 (N_17223,N_14159,N_14431);
nor U17224 (N_17224,N_14906,N_13806);
nand U17225 (N_17225,N_13918,N_15283);
nand U17226 (N_17226,N_12868,N_13587);
or U17227 (N_17227,N_13970,N_13384);
and U17228 (N_17228,N_14864,N_15004);
nand U17229 (N_17229,N_12771,N_13517);
or U17230 (N_17230,N_15121,N_14332);
xnor U17231 (N_17231,N_14815,N_13389);
and U17232 (N_17232,N_13761,N_14301);
nand U17233 (N_17233,N_15098,N_12546);
nand U17234 (N_17234,N_12549,N_13357);
or U17235 (N_17235,N_14950,N_13990);
or U17236 (N_17236,N_13741,N_13584);
and U17237 (N_17237,N_13236,N_14514);
nand U17238 (N_17238,N_13160,N_14826);
nand U17239 (N_17239,N_12956,N_15576);
nor U17240 (N_17240,N_15031,N_15479);
or U17241 (N_17241,N_14508,N_12761);
nor U17242 (N_17242,N_13893,N_13065);
or U17243 (N_17243,N_14394,N_14585);
nor U17244 (N_17244,N_13060,N_12999);
xnor U17245 (N_17245,N_12829,N_13145);
nor U17246 (N_17246,N_14864,N_14136);
and U17247 (N_17247,N_13113,N_15448);
nor U17248 (N_17248,N_15195,N_14559);
nor U17249 (N_17249,N_13576,N_12598);
and U17250 (N_17250,N_13842,N_12756);
or U17251 (N_17251,N_15260,N_15316);
nor U17252 (N_17252,N_13450,N_14598);
and U17253 (N_17253,N_14601,N_13581);
nand U17254 (N_17254,N_15217,N_13411);
nand U17255 (N_17255,N_15195,N_13934);
or U17256 (N_17256,N_15436,N_13763);
and U17257 (N_17257,N_15469,N_12901);
nor U17258 (N_17258,N_13560,N_14474);
nor U17259 (N_17259,N_14702,N_14582);
and U17260 (N_17260,N_12899,N_14908);
or U17261 (N_17261,N_14030,N_13283);
and U17262 (N_17262,N_15234,N_13636);
or U17263 (N_17263,N_13333,N_15082);
and U17264 (N_17264,N_14764,N_15510);
xnor U17265 (N_17265,N_13992,N_13383);
and U17266 (N_17266,N_15392,N_13778);
and U17267 (N_17267,N_13846,N_13789);
and U17268 (N_17268,N_15248,N_14471);
nor U17269 (N_17269,N_14388,N_14345);
and U17270 (N_17270,N_12927,N_14982);
nor U17271 (N_17271,N_14011,N_15062);
and U17272 (N_17272,N_13749,N_15236);
nor U17273 (N_17273,N_12506,N_14074);
nor U17274 (N_17274,N_13667,N_13081);
and U17275 (N_17275,N_14656,N_14383);
or U17276 (N_17276,N_13498,N_12963);
nor U17277 (N_17277,N_14546,N_13396);
and U17278 (N_17278,N_12894,N_13123);
nand U17279 (N_17279,N_14585,N_14884);
and U17280 (N_17280,N_14932,N_14986);
or U17281 (N_17281,N_12500,N_13419);
or U17282 (N_17282,N_14086,N_14659);
nand U17283 (N_17283,N_14359,N_15441);
xnor U17284 (N_17284,N_12800,N_13479);
nand U17285 (N_17285,N_13841,N_14152);
or U17286 (N_17286,N_13176,N_15514);
and U17287 (N_17287,N_12629,N_14491);
nor U17288 (N_17288,N_13614,N_15161);
nand U17289 (N_17289,N_14075,N_14679);
nor U17290 (N_17290,N_15613,N_12810);
nand U17291 (N_17291,N_13679,N_12879);
or U17292 (N_17292,N_14450,N_13604);
or U17293 (N_17293,N_14754,N_12522);
or U17294 (N_17294,N_13339,N_13993);
nand U17295 (N_17295,N_12962,N_12920);
and U17296 (N_17296,N_13265,N_15020);
nand U17297 (N_17297,N_14950,N_13374);
and U17298 (N_17298,N_14598,N_13885);
nand U17299 (N_17299,N_13230,N_13637);
or U17300 (N_17300,N_15036,N_12589);
nor U17301 (N_17301,N_15485,N_14327);
or U17302 (N_17302,N_15142,N_15339);
or U17303 (N_17303,N_13752,N_15569);
nor U17304 (N_17304,N_14321,N_14078);
nand U17305 (N_17305,N_14634,N_15610);
nand U17306 (N_17306,N_13146,N_14320);
and U17307 (N_17307,N_13475,N_14441);
nor U17308 (N_17308,N_15471,N_15037);
nor U17309 (N_17309,N_15469,N_14020);
nand U17310 (N_17310,N_13476,N_13033);
nor U17311 (N_17311,N_14996,N_15142);
and U17312 (N_17312,N_14240,N_12831);
nor U17313 (N_17313,N_13994,N_13031);
or U17314 (N_17314,N_15260,N_13952);
and U17315 (N_17315,N_13350,N_12954);
xnor U17316 (N_17316,N_13325,N_13338);
nor U17317 (N_17317,N_13961,N_14296);
nand U17318 (N_17318,N_13982,N_14963);
or U17319 (N_17319,N_14246,N_13912);
nand U17320 (N_17320,N_15287,N_14232);
or U17321 (N_17321,N_15254,N_14790);
nand U17322 (N_17322,N_13227,N_15483);
and U17323 (N_17323,N_14676,N_12637);
nor U17324 (N_17324,N_14723,N_13669);
and U17325 (N_17325,N_13785,N_14183);
nand U17326 (N_17326,N_13891,N_13516);
or U17327 (N_17327,N_13309,N_13728);
xnor U17328 (N_17328,N_15299,N_13800);
nor U17329 (N_17329,N_14024,N_12872);
nand U17330 (N_17330,N_15358,N_15519);
nand U17331 (N_17331,N_14806,N_12701);
nand U17332 (N_17332,N_15431,N_13557);
nor U17333 (N_17333,N_13565,N_15362);
nor U17334 (N_17334,N_14621,N_12690);
xor U17335 (N_17335,N_14353,N_15059);
nand U17336 (N_17336,N_15492,N_15546);
xor U17337 (N_17337,N_12749,N_13516);
nand U17338 (N_17338,N_15421,N_12645);
nor U17339 (N_17339,N_14951,N_13890);
nor U17340 (N_17340,N_13436,N_13246);
or U17341 (N_17341,N_13287,N_14452);
nor U17342 (N_17342,N_14682,N_15122);
nand U17343 (N_17343,N_13184,N_14631);
nand U17344 (N_17344,N_14560,N_12954);
and U17345 (N_17345,N_13701,N_15603);
nand U17346 (N_17346,N_12504,N_14033);
or U17347 (N_17347,N_13744,N_13466);
xor U17348 (N_17348,N_15413,N_14301);
and U17349 (N_17349,N_13294,N_14511);
or U17350 (N_17350,N_15379,N_12803);
nor U17351 (N_17351,N_13382,N_15078);
or U17352 (N_17352,N_13092,N_14634);
nand U17353 (N_17353,N_13346,N_13794);
and U17354 (N_17354,N_15531,N_14263);
nand U17355 (N_17355,N_12562,N_15245);
nand U17356 (N_17356,N_15596,N_13139);
or U17357 (N_17357,N_13891,N_13097);
nor U17358 (N_17358,N_13914,N_14405);
or U17359 (N_17359,N_15437,N_15155);
or U17360 (N_17360,N_15074,N_12680);
nand U17361 (N_17361,N_15176,N_13068);
nor U17362 (N_17362,N_15568,N_15575);
and U17363 (N_17363,N_14723,N_14324);
or U17364 (N_17364,N_13197,N_15410);
nor U17365 (N_17365,N_15015,N_13969);
or U17366 (N_17366,N_14940,N_13629);
and U17367 (N_17367,N_15100,N_13533);
and U17368 (N_17368,N_15449,N_14459);
and U17369 (N_17369,N_14271,N_12612);
nand U17370 (N_17370,N_13848,N_14161);
and U17371 (N_17371,N_13239,N_15058);
and U17372 (N_17372,N_15099,N_14546);
and U17373 (N_17373,N_14701,N_15414);
and U17374 (N_17374,N_12553,N_12795);
nor U17375 (N_17375,N_14661,N_14054);
and U17376 (N_17376,N_12568,N_13566);
nor U17377 (N_17377,N_12705,N_14925);
xor U17378 (N_17378,N_13427,N_14465);
nand U17379 (N_17379,N_15085,N_13130);
or U17380 (N_17380,N_14913,N_14980);
or U17381 (N_17381,N_15582,N_15004);
and U17382 (N_17382,N_15449,N_13279);
and U17383 (N_17383,N_13327,N_14818);
or U17384 (N_17384,N_14694,N_14433);
nand U17385 (N_17385,N_14024,N_14072);
or U17386 (N_17386,N_13297,N_14875);
and U17387 (N_17387,N_13479,N_13993);
and U17388 (N_17388,N_13699,N_14804);
and U17389 (N_17389,N_13032,N_13444);
nor U17390 (N_17390,N_15143,N_13645);
nor U17391 (N_17391,N_13354,N_15431);
nand U17392 (N_17392,N_13922,N_12920);
nand U17393 (N_17393,N_15473,N_14387);
and U17394 (N_17394,N_14748,N_14282);
or U17395 (N_17395,N_12594,N_13890);
or U17396 (N_17396,N_14850,N_14630);
or U17397 (N_17397,N_12558,N_13188);
nand U17398 (N_17398,N_14322,N_13128);
and U17399 (N_17399,N_12802,N_14083);
and U17400 (N_17400,N_13132,N_15255);
xor U17401 (N_17401,N_14439,N_12611);
nor U17402 (N_17402,N_14186,N_14655);
xnor U17403 (N_17403,N_14776,N_15088);
nand U17404 (N_17404,N_14455,N_15435);
xnor U17405 (N_17405,N_14686,N_14208);
nor U17406 (N_17406,N_14666,N_12731);
and U17407 (N_17407,N_14870,N_14327);
or U17408 (N_17408,N_12917,N_13567);
or U17409 (N_17409,N_13394,N_12674);
or U17410 (N_17410,N_14262,N_14411);
nor U17411 (N_17411,N_15373,N_15454);
and U17412 (N_17412,N_14016,N_14720);
xor U17413 (N_17413,N_13927,N_14589);
xor U17414 (N_17414,N_14059,N_13267);
nand U17415 (N_17415,N_12779,N_14090);
nor U17416 (N_17416,N_14163,N_13441);
or U17417 (N_17417,N_12892,N_14668);
nand U17418 (N_17418,N_14299,N_13906);
nor U17419 (N_17419,N_13446,N_15345);
and U17420 (N_17420,N_14171,N_14474);
and U17421 (N_17421,N_13359,N_15033);
and U17422 (N_17422,N_13163,N_15103);
or U17423 (N_17423,N_14000,N_14689);
nor U17424 (N_17424,N_13897,N_12633);
nand U17425 (N_17425,N_15065,N_15277);
and U17426 (N_17426,N_15442,N_14670);
nand U17427 (N_17427,N_13256,N_14145);
and U17428 (N_17428,N_14661,N_13492);
xor U17429 (N_17429,N_14608,N_12550);
xnor U17430 (N_17430,N_14484,N_13004);
or U17431 (N_17431,N_13026,N_13250);
nand U17432 (N_17432,N_15483,N_12536);
and U17433 (N_17433,N_14814,N_13675);
nor U17434 (N_17434,N_15567,N_15180);
nand U17435 (N_17435,N_13317,N_15613);
or U17436 (N_17436,N_15129,N_14107);
and U17437 (N_17437,N_14338,N_13870);
nor U17438 (N_17438,N_13409,N_14955);
or U17439 (N_17439,N_14425,N_14109);
and U17440 (N_17440,N_14193,N_13327);
or U17441 (N_17441,N_13926,N_13656);
nand U17442 (N_17442,N_15222,N_14270);
nand U17443 (N_17443,N_13380,N_13425);
or U17444 (N_17444,N_12686,N_14726);
or U17445 (N_17445,N_15530,N_14826);
and U17446 (N_17446,N_14206,N_12951);
nand U17447 (N_17447,N_14423,N_12590);
and U17448 (N_17448,N_13461,N_13904);
nand U17449 (N_17449,N_13273,N_13542);
nand U17450 (N_17450,N_14729,N_14587);
nor U17451 (N_17451,N_12512,N_15589);
nand U17452 (N_17452,N_13454,N_12955);
nor U17453 (N_17453,N_14385,N_14306);
and U17454 (N_17454,N_13544,N_15361);
xor U17455 (N_17455,N_14856,N_13937);
and U17456 (N_17456,N_14569,N_13824);
or U17457 (N_17457,N_14244,N_13880);
nand U17458 (N_17458,N_12792,N_13928);
nand U17459 (N_17459,N_14183,N_13169);
nor U17460 (N_17460,N_13127,N_13265);
nand U17461 (N_17461,N_15531,N_12781);
and U17462 (N_17462,N_14587,N_13462);
nand U17463 (N_17463,N_14672,N_15048);
xnor U17464 (N_17464,N_13881,N_14405);
or U17465 (N_17465,N_15194,N_12688);
nor U17466 (N_17466,N_14375,N_14548);
or U17467 (N_17467,N_13580,N_14757);
xor U17468 (N_17468,N_15088,N_14200);
nor U17469 (N_17469,N_14869,N_13790);
nor U17470 (N_17470,N_14543,N_13657);
and U17471 (N_17471,N_13934,N_14458);
xor U17472 (N_17472,N_13402,N_13632);
nand U17473 (N_17473,N_12969,N_14191);
nor U17474 (N_17474,N_13947,N_12834);
and U17475 (N_17475,N_14821,N_14732);
nand U17476 (N_17476,N_13922,N_12795);
nand U17477 (N_17477,N_14566,N_14627);
nand U17478 (N_17478,N_14758,N_13803);
xnor U17479 (N_17479,N_15359,N_12847);
or U17480 (N_17480,N_13239,N_14026);
nor U17481 (N_17481,N_12800,N_14511);
nand U17482 (N_17482,N_12992,N_12870);
or U17483 (N_17483,N_14490,N_15427);
or U17484 (N_17484,N_14062,N_13067);
nand U17485 (N_17485,N_14226,N_13639);
or U17486 (N_17486,N_13272,N_14152);
nand U17487 (N_17487,N_12786,N_15582);
and U17488 (N_17488,N_14572,N_14914);
nor U17489 (N_17489,N_13321,N_13483);
nor U17490 (N_17490,N_14505,N_14196);
xnor U17491 (N_17491,N_15205,N_12878);
nor U17492 (N_17492,N_14145,N_12759);
or U17493 (N_17493,N_14534,N_13895);
and U17494 (N_17494,N_14837,N_15332);
or U17495 (N_17495,N_13292,N_15552);
xor U17496 (N_17496,N_14962,N_15288);
and U17497 (N_17497,N_13194,N_13221);
xor U17498 (N_17498,N_15566,N_15248);
nor U17499 (N_17499,N_13797,N_13941);
xor U17500 (N_17500,N_12767,N_12725);
nand U17501 (N_17501,N_14960,N_13277);
nand U17502 (N_17502,N_14176,N_14671);
nor U17503 (N_17503,N_14765,N_13665);
or U17504 (N_17504,N_15373,N_13697);
nor U17505 (N_17505,N_13134,N_15617);
xnor U17506 (N_17506,N_15080,N_14590);
nor U17507 (N_17507,N_15162,N_14146);
and U17508 (N_17508,N_13408,N_14098);
or U17509 (N_17509,N_14194,N_15108);
or U17510 (N_17510,N_14991,N_13712);
xnor U17511 (N_17511,N_14364,N_13347);
or U17512 (N_17512,N_15192,N_12791);
or U17513 (N_17513,N_14042,N_12765);
xor U17514 (N_17514,N_12643,N_14142);
nor U17515 (N_17515,N_13563,N_14707);
nor U17516 (N_17516,N_14238,N_13529);
nand U17517 (N_17517,N_13833,N_13739);
or U17518 (N_17518,N_13920,N_14608);
or U17519 (N_17519,N_15229,N_14133);
and U17520 (N_17520,N_15454,N_13741);
nand U17521 (N_17521,N_13977,N_13852);
nor U17522 (N_17522,N_13637,N_14210);
xor U17523 (N_17523,N_14285,N_15010);
nand U17524 (N_17524,N_13344,N_15482);
nand U17525 (N_17525,N_15173,N_14587);
nand U17526 (N_17526,N_14449,N_15116);
or U17527 (N_17527,N_13474,N_13735);
nor U17528 (N_17528,N_14326,N_15605);
nand U17529 (N_17529,N_15468,N_13563);
or U17530 (N_17530,N_13848,N_13750);
and U17531 (N_17531,N_13470,N_15108);
and U17532 (N_17532,N_13597,N_14715);
nor U17533 (N_17533,N_14190,N_13093);
and U17534 (N_17534,N_13660,N_13943);
or U17535 (N_17535,N_14832,N_15053);
and U17536 (N_17536,N_14387,N_13831);
nor U17537 (N_17537,N_15377,N_14584);
or U17538 (N_17538,N_14041,N_15603);
nor U17539 (N_17539,N_13861,N_14325);
or U17540 (N_17540,N_12946,N_13485);
nand U17541 (N_17541,N_13644,N_15225);
nand U17542 (N_17542,N_12875,N_12614);
nand U17543 (N_17543,N_13192,N_13639);
and U17544 (N_17544,N_13082,N_12626);
and U17545 (N_17545,N_13006,N_14297);
nand U17546 (N_17546,N_13542,N_13708);
or U17547 (N_17547,N_15150,N_14786);
and U17548 (N_17548,N_13704,N_15057);
or U17549 (N_17549,N_12860,N_14872);
nor U17550 (N_17550,N_14389,N_13067);
nor U17551 (N_17551,N_14719,N_12953);
and U17552 (N_17552,N_14063,N_12772);
xor U17553 (N_17553,N_13504,N_12863);
nor U17554 (N_17554,N_12925,N_13871);
or U17555 (N_17555,N_14825,N_14351);
nand U17556 (N_17556,N_12914,N_15125);
nand U17557 (N_17557,N_13444,N_14859);
nor U17558 (N_17558,N_12812,N_12927);
nor U17559 (N_17559,N_14833,N_13986);
and U17560 (N_17560,N_12789,N_13194);
nor U17561 (N_17561,N_15547,N_13426);
nor U17562 (N_17562,N_13991,N_15318);
nand U17563 (N_17563,N_12787,N_14305);
and U17564 (N_17564,N_14656,N_13995);
or U17565 (N_17565,N_12751,N_14031);
xnor U17566 (N_17566,N_15318,N_13876);
nor U17567 (N_17567,N_12964,N_14094);
nor U17568 (N_17568,N_14212,N_14912);
or U17569 (N_17569,N_13120,N_13659);
nor U17570 (N_17570,N_13630,N_14206);
nor U17571 (N_17571,N_13087,N_13711);
nor U17572 (N_17572,N_13043,N_15285);
and U17573 (N_17573,N_13003,N_15482);
nor U17574 (N_17574,N_14341,N_13030);
and U17575 (N_17575,N_14691,N_14581);
or U17576 (N_17576,N_15513,N_14593);
nand U17577 (N_17577,N_13591,N_13828);
nand U17578 (N_17578,N_12853,N_15333);
and U17579 (N_17579,N_13965,N_15196);
nand U17580 (N_17580,N_14864,N_13612);
and U17581 (N_17581,N_13569,N_13726);
nor U17582 (N_17582,N_14572,N_12971);
nand U17583 (N_17583,N_15039,N_15404);
nor U17584 (N_17584,N_14969,N_15496);
or U17585 (N_17585,N_12659,N_14253);
xnor U17586 (N_17586,N_15069,N_14180);
or U17587 (N_17587,N_14465,N_15549);
and U17588 (N_17588,N_12921,N_15129);
or U17589 (N_17589,N_12894,N_13255);
or U17590 (N_17590,N_15465,N_13035);
and U17591 (N_17591,N_12966,N_15418);
or U17592 (N_17592,N_14627,N_12739);
nor U17593 (N_17593,N_15540,N_14416);
nor U17594 (N_17594,N_13671,N_14165);
nand U17595 (N_17595,N_13462,N_14926);
or U17596 (N_17596,N_14866,N_13186);
nor U17597 (N_17597,N_14164,N_12562);
nor U17598 (N_17598,N_12807,N_14804);
xnor U17599 (N_17599,N_15530,N_12757);
or U17600 (N_17600,N_15354,N_14258);
or U17601 (N_17601,N_14391,N_13579);
xor U17602 (N_17602,N_15560,N_15310);
and U17603 (N_17603,N_12743,N_15557);
and U17604 (N_17604,N_14221,N_14923);
nor U17605 (N_17605,N_15553,N_14838);
or U17606 (N_17606,N_14414,N_15486);
nor U17607 (N_17607,N_12842,N_13947);
nor U17608 (N_17608,N_15073,N_13195);
nand U17609 (N_17609,N_12505,N_14341);
nor U17610 (N_17610,N_14844,N_12798);
nor U17611 (N_17611,N_15094,N_12751);
xnor U17612 (N_17612,N_15483,N_14766);
nor U17613 (N_17613,N_14944,N_12813);
and U17614 (N_17614,N_14136,N_15562);
nor U17615 (N_17615,N_14469,N_12674);
or U17616 (N_17616,N_15143,N_13769);
xnor U17617 (N_17617,N_14589,N_13069);
nor U17618 (N_17618,N_13499,N_12796);
nor U17619 (N_17619,N_13782,N_14032);
nand U17620 (N_17620,N_13540,N_12860);
nand U17621 (N_17621,N_12928,N_13846);
and U17622 (N_17622,N_13636,N_15530);
and U17623 (N_17623,N_13927,N_14208);
or U17624 (N_17624,N_14375,N_14478);
and U17625 (N_17625,N_13180,N_13732);
or U17626 (N_17626,N_12609,N_15151);
or U17627 (N_17627,N_13140,N_12989);
xor U17628 (N_17628,N_13477,N_15465);
nor U17629 (N_17629,N_14425,N_13638);
nand U17630 (N_17630,N_12573,N_15200);
and U17631 (N_17631,N_13514,N_15209);
xnor U17632 (N_17632,N_12711,N_15604);
nand U17633 (N_17633,N_12991,N_14484);
and U17634 (N_17634,N_12514,N_15011);
nor U17635 (N_17635,N_14577,N_15207);
nand U17636 (N_17636,N_13424,N_15073);
or U17637 (N_17637,N_14173,N_12814);
nor U17638 (N_17638,N_13014,N_14275);
or U17639 (N_17639,N_13724,N_13100);
nor U17640 (N_17640,N_14891,N_14375);
nand U17641 (N_17641,N_14528,N_13445);
and U17642 (N_17642,N_14346,N_13703);
nand U17643 (N_17643,N_13743,N_12508);
nand U17644 (N_17644,N_15568,N_15291);
nand U17645 (N_17645,N_12739,N_13322);
xor U17646 (N_17646,N_12534,N_15198);
nor U17647 (N_17647,N_12731,N_14305);
xnor U17648 (N_17648,N_13377,N_13141);
nor U17649 (N_17649,N_13512,N_15431);
or U17650 (N_17650,N_15125,N_12968);
and U17651 (N_17651,N_15011,N_15199);
nor U17652 (N_17652,N_15437,N_15067);
nor U17653 (N_17653,N_14325,N_14364);
nor U17654 (N_17654,N_13204,N_13200);
nor U17655 (N_17655,N_14773,N_14086);
or U17656 (N_17656,N_13169,N_13122);
and U17657 (N_17657,N_14266,N_12527);
and U17658 (N_17658,N_15286,N_14201);
nor U17659 (N_17659,N_13889,N_13181);
xor U17660 (N_17660,N_14523,N_14581);
and U17661 (N_17661,N_13731,N_14622);
and U17662 (N_17662,N_15065,N_12637);
nand U17663 (N_17663,N_13230,N_15468);
nand U17664 (N_17664,N_15230,N_12952);
nand U17665 (N_17665,N_13093,N_14389);
nor U17666 (N_17666,N_13824,N_14875);
nor U17667 (N_17667,N_14619,N_14104);
nor U17668 (N_17668,N_13361,N_14214);
nor U17669 (N_17669,N_14995,N_14618);
nand U17670 (N_17670,N_15262,N_15383);
or U17671 (N_17671,N_13528,N_14776);
nor U17672 (N_17672,N_14308,N_14557);
nor U17673 (N_17673,N_12717,N_13999);
and U17674 (N_17674,N_13360,N_13640);
nand U17675 (N_17675,N_14585,N_14356);
nand U17676 (N_17676,N_13385,N_13603);
or U17677 (N_17677,N_14368,N_15492);
or U17678 (N_17678,N_14540,N_13611);
and U17679 (N_17679,N_13059,N_13567);
nand U17680 (N_17680,N_13873,N_15181);
nand U17681 (N_17681,N_13229,N_14700);
nand U17682 (N_17682,N_13697,N_12782);
nor U17683 (N_17683,N_13048,N_14733);
and U17684 (N_17684,N_13535,N_15052);
nand U17685 (N_17685,N_13450,N_14830);
nor U17686 (N_17686,N_13208,N_13759);
or U17687 (N_17687,N_14106,N_12664);
xor U17688 (N_17688,N_12622,N_13914);
nor U17689 (N_17689,N_12789,N_14816);
and U17690 (N_17690,N_14733,N_13579);
and U17691 (N_17691,N_14216,N_13750);
nand U17692 (N_17692,N_13945,N_14900);
or U17693 (N_17693,N_13541,N_13609);
or U17694 (N_17694,N_15176,N_14517);
or U17695 (N_17695,N_13252,N_15271);
nor U17696 (N_17696,N_14225,N_15001);
and U17697 (N_17697,N_12860,N_15361);
nand U17698 (N_17698,N_14486,N_13026);
nand U17699 (N_17699,N_13956,N_15233);
or U17700 (N_17700,N_13071,N_14463);
or U17701 (N_17701,N_15348,N_14367);
nor U17702 (N_17702,N_13339,N_15102);
xnor U17703 (N_17703,N_13248,N_14278);
xnor U17704 (N_17704,N_15523,N_13032);
or U17705 (N_17705,N_12878,N_14937);
and U17706 (N_17706,N_13850,N_13202);
or U17707 (N_17707,N_15326,N_15300);
or U17708 (N_17708,N_15176,N_13544);
or U17709 (N_17709,N_13191,N_15619);
nor U17710 (N_17710,N_12928,N_15121);
nor U17711 (N_17711,N_14047,N_14046);
or U17712 (N_17712,N_14975,N_14279);
nand U17713 (N_17713,N_13140,N_12900);
and U17714 (N_17714,N_14799,N_13463);
nor U17715 (N_17715,N_12569,N_12660);
or U17716 (N_17716,N_13904,N_12992);
xnor U17717 (N_17717,N_13831,N_14156);
nor U17718 (N_17718,N_13068,N_15315);
nand U17719 (N_17719,N_14876,N_14284);
and U17720 (N_17720,N_15261,N_15020);
nand U17721 (N_17721,N_13142,N_14917);
nor U17722 (N_17722,N_13215,N_14042);
and U17723 (N_17723,N_14637,N_12761);
or U17724 (N_17724,N_14467,N_14922);
nand U17725 (N_17725,N_14858,N_14549);
nand U17726 (N_17726,N_14933,N_13439);
and U17727 (N_17727,N_12684,N_13438);
xor U17728 (N_17728,N_15316,N_15617);
and U17729 (N_17729,N_12600,N_15524);
and U17730 (N_17730,N_14593,N_15130);
and U17731 (N_17731,N_14027,N_14494);
nor U17732 (N_17732,N_13279,N_14862);
or U17733 (N_17733,N_12918,N_15130);
or U17734 (N_17734,N_14220,N_13319);
or U17735 (N_17735,N_13954,N_14088);
or U17736 (N_17736,N_14338,N_14557);
nor U17737 (N_17737,N_13440,N_13509);
nor U17738 (N_17738,N_12756,N_14811);
and U17739 (N_17739,N_13476,N_13228);
nand U17740 (N_17740,N_13107,N_13973);
or U17741 (N_17741,N_15340,N_12785);
nor U17742 (N_17742,N_15426,N_13356);
and U17743 (N_17743,N_14593,N_12901);
nand U17744 (N_17744,N_12982,N_12510);
nand U17745 (N_17745,N_15467,N_13173);
nor U17746 (N_17746,N_13823,N_14349);
and U17747 (N_17747,N_14760,N_12561);
and U17748 (N_17748,N_15565,N_13301);
nand U17749 (N_17749,N_13530,N_15386);
and U17750 (N_17750,N_15611,N_14105);
xor U17751 (N_17751,N_13557,N_14259);
nand U17752 (N_17752,N_13055,N_14798);
nor U17753 (N_17753,N_13731,N_14157);
and U17754 (N_17754,N_15028,N_14186);
or U17755 (N_17755,N_13288,N_12581);
nand U17756 (N_17756,N_13155,N_15063);
or U17757 (N_17757,N_14960,N_13522);
nor U17758 (N_17758,N_14140,N_13926);
xor U17759 (N_17759,N_13710,N_12825);
and U17760 (N_17760,N_13030,N_15021);
and U17761 (N_17761,N_14937,N_14522);
nand U17762 (N_17762,N_15456,N_14612);
nor U17763 (N_17763,N_15605,N_13946);
xor U17764 (N_17764,N_13471,N_14545);
or U17765 (N_17765,N_14428,N_14646);
nor U17766 (N_17766,N_13404,N_14637);
or U17767 (N_17767,N_14703,N_15299);
and U17768 (N_17768,N_15577,N_13806);
and U17769 (N_17769,N_12759,N_13776);
or U17770 (N_17770,N_12954,N_12866);
or U17771 (N_17771,N_15099,N_13657);
or U17772 (N_17772,N_14487,N_13670);
nor U17773 (N_17773,N_13799,N_14767);
or U17774 (N_17774,N_12989,N_13066);
or U17775 (N_17775,N_12911,N_13472);
xnor U17776 (N_17776,N_12948,N_14307);
nand U17777 (N_17777,N_15315,N_14027);
xnor U17778 (N_17778,N_12714,N_13892);
nor U17779 (N_17779,N_15441,N_15604);
nand U17780 (N_17780,N_14892,N_13629);
xor U17781 (N_17781,N_15006,N_14838);
xnor U17782 (N_17782,N_13641,N_13201);
nor U17783 (N_17783,N_15172,N_13749);
or U17784 (N_17784,N_14710,N_14972);
or U17785 (N_17785,N_14745,N_15416);
nand U17786 (N_17786,N_15125,N_14441);
or U17787 (N_17787,N_15240,N_12557);
xnor U17788 (N_17788,N_14472,N_12899);
nor U17789 (N_17789,N_14533,N_14128);
or U17790 (N_17790,N_14388,N_15177);
nand U17791 (N_17791,N_13017,N_15179);
nor U17792 (N_17792,N_14031,N_12789);
nand U17793 (N_17793,N_12776,N_13759);
nand U17794 (N_17794,N_12543,N_13077);
nand U17795 (N_17795,N_13388,N_12830);
nor U17796 (N_17796,N_13125,N_15343);
nand U17797 (N_17797,N_14546,N_12886);
and U17798 (N_17798,N_12858,N_13579);
nand U17799 (N_17799,N_14970,N_14358);
nand U17800 (N_17800,N_14709,N_14259);
nor U17801 (N_17801,N_13112,N_14113);
nand U17802 (N_17802,N_15038,N_14074);
or U17803 (N_17803,N_15514,N_13432);
and U17804 (N_17804,N_13526,N_12515);
nand U17805 (N_17805,N_14420,N_14231);
nor U17806 (N_17806,N_12665,N_13412);
or U17807 (N_17807,N_14870,N_14768);
or U17808 (N_17808,N_13978,N_13036);
or U17809 (N_17809,N_12964,N_13146);
nor U17810 (N_17810,N_13465,N_13765);
or U17811 (N_17811,N_15290,N_12577);
or U17812 (N_17812,N_13001,N_14474);
xnor U17813 (N_17813,N_12837,N_13152);
or U17814 (N_17814,N_14843,N_12794);
and U17815 (N_17815,N_15197,N_14820);
nor U17816 (N_17816,N_15370,N_12926);
or U17817 (N_17817,N_14989,N_13201);
and U17818 (N_17818,N_14819,N_12778);
nor U17819 (N_17819,N_13245,N_13964);
nor U17820 (N_17820,N_15242,N_14828);
and U17821 (N_17821,N_15369,N_15622);
nand U17822 (N_17822,N_15557,N_13524);
nand U17823 (N_17823,N_13619,N_13525);
xor U17824 (N_17824,N_15180,N_14305);
or U17825 (N_17825,N_14003,N_13931);
and U17826 (N_17826,N_12710,N_13900);
nor U17827 (N_17827,N_13991,N_14914);
or U17828 (N_17828,N_14149,N_14146);
xnor U17829 (N_17829,N_13811,N_15076);
nor U17830 (N_17830,N_12955,N_13506);
xor U17831 (N_17831,N_13472,N_12802);
or U17832 (N_17832,N_14612,N_13154);
nor U17833 (N_17833,N_12794,N_13412);
and U17834 (N_17834,N_13884,N_14680);
nand U17835 (N_17835,N_15247,N_15423);
nand U17836 (N_17836,N_15024,N_15316);
and U17837 (N_17837,N_13173,N_14278);
nor U17838 (N_17838,N_14359,N_13438);
and U17839 (N_17839,N_13796,N_12931);
or U17840 (N_17840,N_14271,N_14112);
or U17841 (N_17841,N_14908,N_14696);
or U17842 (N_17842,N_15463,N_15162);
or U17843 (N_17843,N_15262,N_14208);
and U17844 (N_17844,N_15434,N_12909);
nand U17845 (N_17845,N_13629,N_14540);
nand U17846 (N_17846,N_14278,N_13399);
nor U17847 (N_17847,N_13184,N_13278);
nand U17848 (N_17848,N_12656,N_14042);
nand U17849 (N_17849,N_13465,N_12772);
nand U17850 (N_17850,N_12678,N_14400);
and U17851 (N_17851,N_12706,N_13250);
nor U17852 (N_17852,N_15059,N_13988);
or U17853 (N_17853,N_13778,N_13371);
xor U17854 (N_17854,N_12779,N_14117);
and U17855 (N_17855,N_14111,N_14232);
or U17856 (N_17856,N_12940,N_13767);
nor U17857 (N_17857,N_14393,N_14849);
or U17858 (N_17858,N_14966,N_13518);
or U17859 (N_17859,N_14988,N_12900);
and U17860 (N_17860,N_13698,N_14205);
nor U17861 (N_17861,N_12568,N_13389);
nor U17862 (N_17862,N_13526,N_13139);
nand U17863 (N_17863,N_13529,N_14698);
nor U17864 (N_17864,N_15498,N_13498);
or U17865 (N_17865,N_13016,N_13410);
nor U17866 (N_17866,N_13551,N_14067);
nand U17867 (N_17867,N_12901,N_14282);
nand U17868 (N_17868,N_14566,N_14822);
nor U17869 (N_17869,N_15545,N_14002);
nand U17870 (N_17870,N_13280,N_14387);
nand U17871 (N_17871,N_15428,N_14448);
nand U17872 (N_17872,N_15269,N_14427);
and U17873 (N_17873,N_13068,N_13466);
nand U17874 (N_17874,N_15554,N_15372);
or U17875 (N_17875,N_15352,N_14039);
nand U17876 (N_17876,N_12714,N_14841);
and U17877 (N_17877,N_14471,N_12503);
or U17878 (N_17878,N_14791,N_13870);
nand U17879 (N_17879,N_15400,N_15534);
nand U17880 (N_17880,N_14977,N_15590);
and U17881 (N_17881,N_15570,N_13156);
xor U17882 (N_17882,N_15192,N_13035);
nand U17883 (N_17883,N_12944,N_12812);
nor U17884 (N_17884,N_14431,N_14865);
xnor U17885 (N_17885,N_13362,N_14542);
or U17886 (N_17886,N_12981,N_13481);
and U17887 (N_17887,N_15460,N_15293);
nor U17888 (N_17888,N_15212,N_15605);
and U17889 (N_17889,N_13281,N_15619);
nand U17890 (N_17890,N_13590,N_13559);
nor U17891 (N_17891,N_13032,N_14110);
nand U17892 (N_17892,N_12842,N_15409);
nand U17893 (N_17893,N_14008,N_13862);
and U17894 (N_17894,N_12796,N_12837);
nor U17895 (N_17895,N_13826,N_14320);
nand U17896 (N_17896,N_15546,N_13686);
or U17897 (N_17897,N_12680,N_13133);
and U17898 (N_17898,N_13573,N_13693);
xnor U17899 (N_17899,N_12741,N_13433);
and U17900 (N_17900,N_15084,N_14560);
nor U17901 (N_17901,N_15615,N_13095);
and U17902 (N_17902,N_15515,N_14154);
xor U17903 (N_17903,N_13390,N_14019);
nor U17904 (N_17904,N_13515,N_13803);
and U17905 (N_17905,N_12637,N_12900);
nand U17906 (N_17906,N_15089,N_13222);
or U17907 (N_17907,N_12543,N_15394);
and U17908 (N_17908,N_13760,N_13942);
xor U17909 (N_17909,N_14038,N_12677);
or U17910 (N_17910,N_13192,N_15197);
or U17911 (N_17911,N_15465,N_15560);
nand U17912 (N_17912,N_14453,N_13476);
nor U17913 (N_17913,N_12544,N_14401);
nor U17914 (N_17914,N_14731,N_13410);
and U17915 (N_17915,N_14493,N_13249);
nor U17916 (N_17916,N_13550,N_12808);
xor U17917 (N_17917,N_14674,N_15175);
xor U17918 (N_17918,N_13251,N_14885);
nor U17919 (N_17919,N_14576,N_13282);
nor U17920 (N_17920,N_14087,N_14603);
nand U17921 (N_17921,N_15102,N_15159);
or U17922 (N_17922,N_15162,N_13020);
xor U17923 (N_17923,N_12507,N_14380);
nor U17924 (N_17924,N_13123,N_14574);
and U17925 (N_17925,N_13880,N_12997);
and U17926 (N_17926,N_15591,N_13809);
and U17927 (N_17927,N_12610,N_15208);
xnor U17928 (N_17928,N_12619,N_13460);
nor U17929 (N_17929,N_13406,N_15224);
nand U17930 (N_17930,N_13156,N_14234);
and U17931 (N_17931,N_13313,N_15270);
or U17932 (N_17932,N_13021,N_13017);
nand U17933 (N_17933,N_13697,N_15345);
nand U17934 (N_17934,N_14146,N_12936);
nand U17935 (N_17935,N_15098,N_13903);
nor U17936 (N_17936,N_15323,N_12933);
nor U17937 (N_17937,N_12690,N_14756);
nor U17938 (N_17938,N_14043,N_14840);
nor U17939 (N_17939,N_13511,N_15384);
nand U17940 (N_17940,N_14664,N_13340);
and U17941 (N_17941,N_14965,N_14545);
nor U17942 (N_17942,N_15581,N_15245);
nand U17943 (N_17943,N_14382,N_12536);
nor U17944 (N_17944,N_15073,N_14308);
or U17945 (N_17945,N_13219,N_12912);
and U17946 (N_17946,N_12899,N_15576);
xnor U17947 (N_17947,N_15544,N_12958);
and U17948 (N_17948,N_14725,N_14752);
and U17949 (N_17949,N_12986,N_15356);
nor U17950 (N_17950,N_13856,N_14900);
or U17951 (N_17951,N_14573,N_15215);
and U17952 (N_17952,N_14810,N_14006);
or U17953 (N_17953,N_15103,N_15358);
nor U17954 (N_17954,N_15034,N_13184);
or U17955 (N_17955,N_13296,N_13482);
xor U17956 (N_17956,N_14707,N_15428);
or U17957 (N_17957,N_14533,N_15215);
nand U17958 (N_17958,N_12671,N_15594);
nand U17959 (N_17959,N_14164,N_15417);
and U17960 (N_17960,N_13518,N_15421);
xnor U17961 (N_17961,N_13609,N_15116);
or U17962 (N_17962,N_13558,N_14060);
nand U17963 (N_17963,N_15379,N_13822);
nor U17964 (N_17964,N_12535,N_15575);
nand U17965 (N_17965,N_14767,N_15086);
or U17966 (N_17966,N_13205,N_13582);
or U17967 (N_17967,N_15212,N_14827);
and U17968 (N_17968,N_13745,N_12756);
and U17969 (N_17969,N_13484,N_15475);
nand U17970 (N_17970,N_13372,N_12583);
and U17971 (N_17971,N_14264,N_13753);
or U17972 (N_17972,N_12917,N_14226);
nor U17973 (N_17973,N_14752,N_14444);
nand U17974 (N_17974,N_14194,N_15129);
nor U17975 (N_17975,N_13680,N_14121);
xnor U17976 (N_17976,N_15060,N_13815);
or U17977 (N_17977,N_12770,N_12631);
nand U17978 (N_17978,N_13368,N_12546);
and U17979 (N_17979,N_13242,N_15424);
or U17980 (N_17980,N_14689,N_14513);
and U17981 (N_17981,N_14374,N_13813);
or U17982 (N_17982,N_13821,N_15542);
and U17983 (N_17983,N_14318,N_13985);
or U17984 (N_17984,N_13196,N_13153);
and U17985 (N_17985,N_14602,N_14799);
and U17986 (N_17986,N_14450,N_12532);
or U17987 (N_17987,N_15586,N_13145);
and U17988 (N_17988,N_12577,N_13682);
nand U17989 (N_17989,N_14124,N_14578);
xnor U17990 (N_17990,N_13094,N_14848);
nor U17991 (N_17991,N_14262,N_14016);
and U17992 (N_17992,N_12870,N_14401);
nand U17993 (N_17993,N_14832,N_14756);
nor U17994 (N_17994,N_14130,N_14423);
xor U17995 (N_17995,N_15102,N_13098);
and U17996 (N_17996,N_13719,N_13670);
or U17997 (N_17997,N_15234,N_14442);
or U17998 (N_17998,N_13670,N_12524);
or U17999 (N_17999,N_15020,N_13593);
or U18000 (N_18000,N_14532,N_15191);
or U18001 (N_18001,N_15031,N_15391);
or U18002 (N_18002,N_14627,N_15484);
and U18003 (N_18003,N_14076,N_13581);
or U18004 (N_18004,N_14053,N_14758);
or U18005 (N_18005,N_13281,N_15299);
or U18006 (N_18006,N_13644,N_14065);
xor U18007 (N_18007,N_15401,N_12598);
or U18008 (N_18008,N_13891,N_13244);
or U18009 (N_18009,N_13548,N_13018);
and U18010 (N_18010,N_15367,N_13567);
nand U18011 (N_18011,N_12535,N_14918);
or U18012 (N_18012,N_12872,N_15086);
nor U18013 (N_18013,N_12859,N_14389);
nand U18014 (N_18014,N_14823,N_14893);
nand U18015 (N_18015,N_14112,N_14304);
or U18016 (N_18016,N_12571,N_12819);
nor U18017 (N_18017,N_15036,N_13392);
nor U18018 (N_18018,N_12652,N_14988);
or U18019 (N_18019,N_14688,N_14568);
and U18020 (N_18020,N_14883,N_13467);
nand U18021 (N_18021,N_14190,N_14323);
and U18022 (N_18022,N_15410,N_12720);
nor U18023 (N_18023,N_14541,N_12932);
nor U18024 (N_18024,N_14277,N_13904);
nor U18025 (N_18025,N_13229,N_13799);
xor U18026 (N_18026,N_14789,N_12880);
xnor U18027 (N_18027,N_15040,N_14183);
nand U18028 (N_18028,N_13576,N_14547);
and U18029 (N_18029,N_14305,N_14237);
or U18030 (N_18030,N_14192,N_15380);
or U18031 (N_18031,N_13037,N_13176);
nor U18032 (N_18032,N_12770,N_13501);
nand U18033 (N_18033,N_14725,N_13017);
or U18034 (N_18034,N_13425,N_12720);
nand U18035 (N_18035,N_14710,N_14626);
nand U18036 (N_18036,N_15196,N_12764);
nand U18037 (N_18037,N_13794,N_14952);
xor U18038 (N_18038,N_12649,N_14586);
or U18039 (N_18039,N_13043,N_14425);
nand U18040 (N_18040,N_13973,N_13559);
and U18041 (N_18041,N_15205,N_15578);
xnor U18042 (N_18042,N_13508,N_13809);
or U18043 (N_18043,N_14861,N_13674);
and U18044 (N_18044,N_13548,N_13731);
nor U18045 (N_18045,N_14955,N_13942);
nor U18046 (N_18046,N_15119,N_13487);
or U18047 (N_18047,N_15317,N_14313);
nor U18048 (N_18048,N_13884,N_15484);
or U18049 (N_18049,N_12836,N_12998);
xor U18050 (N_18050,N_13767,N_14828);
or U18051 (N_18051,N_14295,N_15396);
nor U18052 (N_18052,N_15042,N_13489);
and U18053 (N_18053,N_13752,N_14292);
nor U18054 (N_18054,N_13976,N_14460);
nand U18055 (N_18055,N_13789,N_15260);
and U18056 (N_18056,N_14780,N_12545);
nor U18057 (N_18057,N_13564,N_13339);
or U18058 (N_18058,N_14410,N_12533);
nand U18059 (N_18059,N_15372,N_12622);
nand U18060 (N_18060,N_13125,N_14411);
and U18061 (N_18061,N_12763,N_14557);
and U18062 (N_18062,N_15131,N_13024);
and U18063 (N_18063,N_14144,N_12951);
nor U18064 (N_18064,N_14405,N_15446);
xnor U18065 (N_18065,N_13081,N_14011);
or U18066 (N_18066,N_15334,N_14553);
nand U18067 (N_18067,N_15432,N_12774);
nand U18068 (N_18068,N_13008,N_13767);
nor U18069 (N_18069,N_14404,N_13436);
xnor U18070 (N_18070,N_13107,N_12792);
and U18071 (N_18071,N_13127,N_13501);
and U18072 (N_18072,N_15613,N_12602);
and U18073 (N_18073,N_15108,N_15426);
or U18074 (N_18074,N_12792,N_13486);
and U18075 (N_18075,N_14435,N_14229);
nand U18076 (N_18076,N_13021,N_13333);
nand U18077 (N_18077,N_12786,N_13234);
or U18078 (N_18078,N_12824,N_13189);
or U18079 (N_18079,N_12568,N_12626);
nand U18080 (N_18080,N_15442,N_13533);
nand U18081 (N_18081,N_12924,N_14013);
nor U18082 (N_18082,N_13884,N_13637);
nor U18083 (N_18083,N_14354,N_15329);
or U18084 (N_18084,N_14607,N_14307);
nand U18085 (N_18085,N_14600,N_14798);
xor U18086 (N_18086,N_13765,N_15237);
nor U18087 (N_18087,N_13464,N_15028);
and U18088 (N_18088,N_14065,N_14988);
or U18089 (N_18089,N_12541,N_13503);
or U18090 (N_18090,N_14357,N_12736);
nor U18091 (N_18091,N_13584,N_13847);
and U18092 (N_18092,N_15089,N_13998);
xor U18093 (N_18093,N_14698,N_13207);
nor U18094 (N_18094,N_14742,N_13986);
nor U18095 (N_18095,N_12653,N_14879);
and U18096 (N_18096,N_13697,N_15290);
and U18097 (N_18097,N_12917,N_14554);
nor U18098 (N_18098,N_13983,N_12737);
nand U18099 (N_18099,N_12859,N_12938);
nand U18100 (N_18100,N_14522,N_14449);
and U18101 (N_18101,N_13546,N_12503);
and U18102 (N_18102,N_12753,N_13302);
nor U18103 (N_18103,N_14973,N_15423);
xnor U18104 (N_18104,N_13490,N_15195);
or U18105 (N_18105,N_12863,N_13919);
nand U18106 (N_18106,N_15598,N_14413);
nor U18107 (N_18107,N_13397,N_14851);
or U18108 (N_18108,N_12986,N_13785);
xnor U18109 (N_18109,N_13331,N_12948);
xor U18110 (N_18110,N_15242,N_13862);
nand U18111 (N_18111,N_13799,N_14282);
nand U18112 (N_18112,N_12512,N_13784);
nor U18113 (N_18113,N_14161,N_15052);
nand U18114 (N_18114,N_13291,N_15396);
and U18115 (N_18115,N_13661,N_13852);
nand U18116 (N_18116,N_14172,N_13590);
nand U18117 (N_18117,N_13891,N_12578);
and U18118 (N_18118,N_13097,N_15102);
or U18119 (N_18119,N_13154,N_13218);
or U18120 (N_18120,N_12547,N_13301);
nor U18121 (N_18121,N_13271,N_14759);
nand U18122 (N_18122,N_13118,N_14828);
xnor U18123 (N_18123,N_14176,N_14098);
nor U18124 (N_18124,N_14421,N_15293);
and U18125 (N_18125,N_13151,N_13780);
xor U18126 (N_18126,N_14380,N_13450);
nand U18127 (N_18127,N_14148,N_14454);
or U18128 (N_18128,N_15510,N_14115);
or U18129 (N_18129,N_13224,N_13566);
nand U18130 (N_18130,N_14357,N_12633);
nor U18131 (N_18131,N_14272,N_12645);
and U18132 (N_18132,N_13998,N_14298);
or U18133 (N_18133,N_12659,N_12822);
nand U18134 (N_18134,N_13401,N_15262);
or U18135 (N_18135,N_15247,N_14554);
nand U18136 (N_18136,N_13362,N_12549);
or U18137 (N_18137,N_14901,N_14135);
nor U18138 (N_18138,N_14896,N_12521);
xnor U18139 (N_18139,N_15502,N_12870);
and U18140 (N_18140,N_13804,N_14605);
or U18141 (N_18141,N_13210,N_13592);
xor U18142 (N_18142,N_13725,N_12979);
nor U18143 (N_18143,N_12572,N_12718);
and U18144 (N_18144,N_12874,N_12981);
nand U18145 (N_18145,N_13936,N_13994);
and U18146 (N_18146,N_13019,N_12688);
or U18147 (N_18147,N_13061,N_15245);
or U18148 (N_18148,N_13691,N_13140);
nand U18149 (N_18149,N_13944,N_14287);
xor U18150 (N_18150,N_13271,N_15344);
nor U18151 (N_18151,N_14723,N_15079);
xor U18152 (N_18152,N_14807,N_15591);
nand U18153 (N_18153,N_15375,N_15591);
and U18154 (N_18154,N_13714,N_13765);
and U18155 (N_18155,N_14784,N_12963);
xnor U18156 (N_18156,N_15329,N_14958);
nand U18157 (N_18157,N_14239,N_14874);
nand U18158 (N_18158,N_13654,N_14689);
nor U18159 (N_18159,N_15453,N_13304);
nor U18160 (N_18160,N_14020,N_13936);
nor U18161 (N_18161,N_13833,N_13660);
nand U18162 (N_18162,N_15287,N_13559);
nor U18163 (N_18163,N_15319,N_14922);
or U18164 (N_18164,N_13510,N_14940);
nand U18165 (N_18165,N_14312,N_14860);
and U18166 (N_18166,N_12906,N_12974);
nand U18167 (N_18167,N_15339,N_15122);
or U18168 (N_18168,N_14145,N_14111);
and U18169 (N_18169,N_14679,N_14845);
and U18170 (N_18170,N_15127,N_15394);
or U18171 (N_18171,N_12911,N_14590);
nor U18172 (N_18172,N_13657,N_15535);
nand U18173 (N_18173,N_15086,N_13992);
nand U18174 (N_18174,N_15244,N_14607);
nor U18175 (N_18175,N_14143,N_15173);
and U18176 (N_18176,N_14003,N_13563);
xnor U18177 (N_18177,N_13994,N_12508);
xor U18178 (N_18178,N_14263,N_14204);
nand U18179 (N_18179,N_14580,N_15251);
nor U18180 (N_18180,N_13198,N_12532);
and U18181 (N_18181,N_15451,N_12782);
and U18182 (N_18182,N_13279,N_14196);
nor U18183 (N_18183,N_15359,N_15146);
or U18184 (N_18184,N_14462,N_13553);
nand U18185 (N_18185,N_14270,N_15249);
and U18186 (N_18186,N_15190,N_14777);
or U18187 (N_18187,N_15115,N_14374);
nand U18188 (N_18188,N_15220,N_15444);
or U18189 (N_18189,N_14295,N_13267);
nand U18190 (N_18190,N_15511,N_15611);
nand U18191 (N_18191,N_13267,N_15417);
and U18192 (N_18192,N_14839,N_14120);
and U18193 (N_18193,N_12530,N_13796);
and U18194 (N_18194,N_13258,N_14394);
nor U18195 (N_18195,N_12874,N_13922);
nor U18196 (N_18196,N_12731,N_12722);
nand U18197 (N_18197,N_14959,N_14875);
or U18198 (N_18198,N_15024,N_12929);
or U18199 (N_18199,N_13468,N_12913);
nor U18200 (N_18200,N_13187,N_13730);
and U18201 (N_18201,N_13442,N_12625);
and U18202 (N_18202,N_14175,N_13585);
nand U18203 (N_18203,N_14682,N_13818);
and U18204 (N_18204,N_15466,N_14764);
nand U18205 (N_18205,N_15280,N_14549);
xnor U18206 (N_18206,N_15274,N_13013);
nor U18207 (N_18207,N_15501,N_14179);
and U18208 (N_18208,N_15420,N_14978);
or U18209 (N_18209,N_15576,N_14113);
or U18210 (N_18210,N_12828,N_14321);
nor U18211 (N_18211,N_14628,N_14163);
xor U18212 (N_18212,N_13760,N_14879);
xnor U18213 (N_18213,N_12943,N_12662);
xor U18214 (N_18214,N_14416,N_13878);
and U18215 (N_18215,N_13621,N_15572);
nand U18216 (N_18216,N_13405,N_14510);
and U18217 (N_18217,N_13140,N_13107);
and U18218 (N_18218,N_14866,N_14940);
nand U18219 (N_18219,N_15341,N_14133);
and U18220 (N_18220,N_15070,N_15516);
xnor U18221 (N_18221,N_14418,N_13309);
and U18222 (N_18222,N_14513,N_12979);
nor U18223 (N_18223,N_12815,N_12681);
nor U18224 (N_18224,N_14641,N_13458);
nor U18225 (N_18225,N_15460,N_12984);
nor U18226 (N_18226,N_15002,N_13303);
nand U18227 (N_18227,N_13168,N_14154);
and U18228 (N_18228,N_14612,N_13328);
and U18229 (N_18229,N_14921,N_13952);
nor U18230 (N_18230,N_13726,N_14002);
xor U18231 (N_18231,N_15217,N_15454);
xor U18232 (N_18232,N_15193,N_13508);
nor U18233 (N_18233,N_14034,N_12802);
nand U18234 (N_18234,N_13418,N_12530);
xor U18235 (N_18235,N_13025,N_13537);
and U18236 (N_18236,N_12799,N_13810);
or U18237 (N_18237,N_14290,N_14471);
nand U18238 (N_18238,N_14306,N_13277);
and U18239 (N_18239,N_14226,N_13581);
xnor U18240 (N_18240,N_13484,N_13885);
nor U18241 (N_18241,N_12645,N_12711);
nand U18242 (N_18242,N_15411,N_12800);
or U18243 (N_18243,N_13229,N_13675);
nor U18244 (N_18244,N_13598,N_14512);
or U18245 (N_18245,N_15502,N_14119);
nor U18246 (N_18246,N_12940,N_14522);
or U18247 (N_18247,N_14623,N_15101);
nand U18248 (N_18248,N_13051,N_13510);
and U18249 (N_18249,N_14083,N_14792);
nand U18250 (N_18250,N_14008,N_14326);
nand U18251 (N_18251,N_15209,N_13439);
and U18252 (N_18252,N_14573,N_12520);
nor U18253 (N_18253,N_15259,N_14840);
or U18254 (N_18254,N_14030,N_13275);
and U18255 (N_18255,N_12722,N_13777);
and U18256 (N_18256,N_12836,N_13789);
nor U18257 (N_18257,N_13833,N_12505);
nand U18258 (N_18258,N_14709,N_12787);
or U18259 (N_18259,N_15466,N_15300);
or U18260 (N_18260,N_13280,N_12868);
xnor U18261 (N_18261,N_15463,N_12896);
and U18262 (N_18262,N_13397,N_15440);
nor U18263 (N_18263,N_14341,N_14068);
nor U18264 (N_18264,N_15020,N_14913);
nand U18265 (N_18265,N_13545,N_12516);
nor U18266 (N_18266,N_12564,N_14550);
xor U18267 (N_18267,N_14062,N_15460);
nor U18268 (N_18268,N_15208,N_14460);
or U18269 (N_18269,N_14142,N_14220);
nand U18270 (N_18270,N_13505,N_14628);
nand U18271 (N_18271,N_13614,N_13020);
nand U18272 (N_18272,N_15361,N_14560);
or U18273 (N_18273,N_13805,N_13078);
nor U18274 (N_18274,N_13801,N_14604);
nand U18275 (N_18275,N_13404,N_12802);
and U18276 (N_18276,N_14424,N_14800);
and U18277 (N_18277,N_13028,N_14798);
and U18278 (N_18278,N_14126,N_14379);
nand U18279 (N_18279,N_15610,N_12637);
nand U18280 (N_18280,N_12988,N_14094);
nand U18281 (N_18281,N_13527,N_13024);
xor U18282 (N_18282,N_14013,N_14356);
nor U18283 (N_18283,N_13765,N_15041);
and U18284 (N_18284,N_14107,N_13628);
or U18285 (N_18285,N_13568,N_14560);
xor U18286 (N_18286,N_13023,N_13535);
nor U18287 (N_18287,N_12840,N_13761);
nand U18288 (N_18288,N_12668,N_15129);
nor U18289 (N_18289,N_14000,N_14485);
or U18290 (N_18290,N_15532,N_13447);
or U18291 (N_18291,N_13534,N_12750);
nand U18292 (N_18292,N_14775,N_14667);
or U18293 (N_18293,N_14756,N_12910);
or U18294 (N_18294,N_15332,N_13029);
and U18295 (N_18295,N_15101,N_14334);
and U18296 (N_18296,N_14177,N_14134);
and U18297 (N_18297,N_12531,N_12991);
xor U18298 (N_18298,N_12553,N_13167);
and U18299 (N_18299,N_12935,N_14749);
nand U18300 (N_18300,N_13341,N_13503);
nor U18301 (N_18301,N_14322,N_14327);
and U18302 (N_18302,N_13865,N_15493);
nor U18303 (N_18303,N_12711,N_14483);
or U18304 (N_18304,N_13213,N_13988);
or U18305 (N_18305,N_14473,N_12913);
and U18306 (N_18306,N_14519,N_15371);
and U18307 (N_18307,N_15611,N_12770);
and U18308 (N_18308,N_12660,N_14716);
nor U18309 (N_18309,N_14938,N_14595);
nor U18310 (N_18310,N_12900,N_12889);
or U18311 (N_18311,N_14722,N_13428);
nor U18312 (N_18312,N_13055,N_13401);
and U18313 (N_18313,N_15121,N_12635);
nand U18314 (N_18314,N_13808,N_14823);
nor U18315 (N_18315,N_13984,N_13246);
or U18316 (N_18316,N_14586,N_14327);
nor U18317 (N_18317,N_13262,N_14075);
or U18318 (N_18318,N_15561,N_13549);
nor U18319 (N_18319,N_15256,N_13260);
nand U18320 (N_18320,N_15207,N_12556);
nand U18321 (N_18321,N_13065,N_13869);
xnor U18322 (N_18322,N_13351,N_14972);
nand U18323 (N_18323,N_14726,N_14280);
nand U18324 (N_18324,N_12834,N_14855);
nor U18325 (N_18325,N_15466,N_12821);
nor U18326 (N_18326,N_13368,N_15581);
nand U18327 (N_18327,N_13722,N_15287);
xnor U18328 (N_18328,N_14507,N_15549);
and U18329 (N_18329,N_14811,N_14439);
nor U18330 (N_18330,N_14015,N_13682);
or U18331 (N_18331,N_14200,N_14911);
nor U18332 (N_18332,N_12730,N_15599);
nor U18333 (N_18333,N_12724,N_13540);
nand U18334 (N_18334,N_14824,N_12746);
and U18335 (N_18335,N_14984,N_13961);
nand U18336 (N_18336,N_13807,N_15155);
or U18337 (N_18337,N_15049,N_14101);
nand U18338 (N_18338,N_14157,N_13580);
or U18339 (N_18339,N_13185,N_14192);
or U18340 (N_18340,N_13658,N_13332);
xnor U18341 (N_18341,N_15600,N_14176);
or U18342 (N_18342,N_12865,N_12576);
nor U18343 (N_18343,N_13429,N_13670);
nor U18344 (N_18344,N_15080,N_12576);
and U18345 (N_18345,N_15289,N_13021);
and U18346 (N_18346,N_13452,N_13660);
and U18347 (N_18347,N_15152,N_14624);
and U18348 (N_18348,N_13882,N_15326);
xnor U18349 (N_18349,N_15020,N_13396);
nand U18350 (N_18350,N_13612,N_13631);
xor U18351 (N_18351,N_15135,N_14457);
xor U18352 (N_18352,N_14776,N_14670);
and U18353 (N_18353,N_13807,N_14196);
nor U18354 (N_18354,N_13802,N_15209);
and U18355 (N_18355,N_15260,N_12989);
and U18356 (N_18356,N_15038,N_12692);
and U18357 (N_18357,N_13877,N_14463);
nand U18358 (N_18358,N_15005,N_14646);
nor U18359 (N_18359,N_13316,N_15428);
and U18360 (N_18360,N_14894,N_14641);
or U18361 (N_18361,N_13785,N_15120);
nand U18362 (N_18362,N_12981,N_13633);
nand U18363 (N_18363,N_12806,N_14158);
nor U18364 (N_18364,N_14581,N_13066);
xnor U18365 (N_18365,N_13671,N_14284);
and U18366 (N_18366,N_12500,N_13489);
xnor U18367 (N_18367,N_15248,N_13698);
xnor U18368 (N_18368,N_12898,N_15595);
or U18369 (N_18369,N_14014,N_15371);
nor U18370 (N_18370,N_13286,N_14137);
or U18371 (N_18371,N_13168,N_13881);
and U18372 (N_18372,N_15372,N_15229);
nor U18373 (N_18373,N_13972,N_15083);
nand U18374 (N_18374,N_13876,N_15015);
and U18375 (N_18375,N_15048,N_12972);
or U18376 (N_18376,N_14427,N_13608);
nor U18377 (N_18377,N_14291,N_13556);
xnor U18378 (N_18378,N_15093,N_12554);
nor U18379 (N_18379,N_14017,N_13757);
or U18380 (N_18380,N_13507,N_13328);
nand U18381 (N_18381,N_13805,N_14261);
nor U18382 (N_18382,N_12571,N_14766);
or U18383 (N_18383,N_14337,N_15054);
nor U18384 (N_18384,N_13549,N_13390);
or U18385 (N_18385,N_15027,N_14256);
and U18386 (N_18386,N_13866,N_15124);
nor U18387 (N_18387,N_14353,N_12538);
nor U18388 (N_18388,N_15300,N_15412);
nand U18389 (N_18389,N_15448,N_14648);
and U18390 (N_18390,N_13529,N_13301);
nor U18391 (N_18391,N_12570,N_13511);
xor U18392 (N_18392,N_14833,N_12820);
nand U18393 (N_18393,N_12578,N_13780);
xnor U18394 (N_18394,N_14877,N_15569);
nand U18395 (N_18395,N_13240,N_14150);
or U18396 (N_18396,N_12849,N_14721);
nand U18397 (N_18397,N_14039,N_13141);
and U18398 (N_18398,N_15304,N_13646);
or U18399 (N_18399,N_15291,N_13796);
and U18400 (N_18400,N_13715,N_14261);
or U18401 (N_18401,N_14362,N_13837);
nand U18402 (N_18402,N_14533,N_12693);
and U18403 (N_18403,N_13679,N_14315);
and U18404 (N_18404,N_13750,N_13069);
nand U18405 (N_18405,N_14303,N_12590);
and U18406 (N_18406,N_13684,N_12638);
nand U18407 (N_18407,N_14166,N_14294);
or U18408 (N_18408,N_14684,N_15601);
nand U18409 (N_18409,N_13282,N_13738);
nand U18410 (N_18410,N_13410,N_12860);
nand U18411 (N_18411,N_15352,N_15462);
and U18412 (N_18412,N_14527,N_15127);
nor U18413 (N_18413,N_14544,N_14456);
and U18414 (N_18414,N_14852,N_13811);
nor U18415 (N_18415,N_13024,N_14041);
xnor U18416 (N_18416,N_12501,N_12737);
and U18417 (N_18417,N_14049,N_15390);
or U18418 (N_18418,N_13331,N_13281);
or U18419 (N_18419,N_14389,N_13859);
or U18420 (N_18420,N_15582,N_14587);
nor U18421 (N_18421,N_14905,N_13384);
nor U18422 (N_18422,N_14634,N_14170);
nand U18423 (N_18423,N_13915,N_13082);
nor U18424 (N_18424,N_14982,N_14840);
xor U18425 (N_18425,N_12868,N_15171);
and U18426 (N_18426,N_13057,N_15375);
xor U18427 (N_18427,N_14904,N_15515);
nand U18428 (N_18428,N_13720,N_14442);
xnor U18429 (N_18429,N_13900,N_13069);
nand U18430 (N_18430,N_15218,N_14991);
xor U18431 (N_18431,N_13174,N_14900);
and U18432 (N_18432,N_12732,N_13285);
xor U18433 (N_18433,N_12838,N_13671);
nor U18434 (N_18434,N_14891,N_12519);
or U18435 (N_18435,N_13311,N_13337);
or U18436 (N_18436,N_13907,N_15045);
xnor U18437 (N_18437,N_13601,N_14722);
nand U18438 (N_18438,N_14411,N_15527);
nor U18439 (N_18439,N_12529,N_12565);
nand U18440 (N_18440,N_13602,N_14117);
nor U18441 (N_18441,N_15294,N_14833);
nand U18442 (N_18442,N_13252,N_15153);
xnor U18443 (N_18443,N_13522,N_15401);
or U18444 (N_18444,N_13242,N_14857);
and U18445 (N_18445,N_13816,N_14336);
or U18446 (N_18446,N_14712,N_15080);
nand U18447 (N_18447,N_13625,N_13344);
nand U18448 (N_18448,N_14145,N_13623);
and U18449 (N_18449,N_14861,N_13229);
xor U18450 (N_18450,N_14736,N_13433);
and U18451 (N_18451,N_13008,N_15401);
and U18452 (N_18452,N_14254,N_14219);
nor U18453 (N_18453,N_12941,N_14755);
and U18454 (N_18454,N_13637,N_12598);
xor U18455 (N_18455,N_15372,N_15495);
nand U18456 (N_18456,N_13176,N_14445);
or U18457 (N_18457,N_15101,N_14946);
xnor U18458 (N_18458,N_13808,N_14625);
nor U18459 (N_18459,N_12779,N_15037);
nand U18460 (N_18460,N_14382,N_12791);
and U18461 (N_18461,N_12523,N_13704);
or U18462 (N_18462,N_14500,N_13124);
nand U18463 (N_18463,N_13082,N_13203);
nor U18464 (N_18464,N_12595,N_13914);
nand U18465 (N_18465,N_13516,N_14826);
nor U18466 (N_18466,N_14708,N_13004);
or U18467 (N_18467,N_12790,N_15081);
nand U18468 (N_18468,N_13754,N_12518);
and U18469 (N_18469,N_14388,N_13643);
nand U18470 (N_18470,N_13966,N_12544);
nand U18471 (N_18471,N_14103,N_12631);
nor U18472 (N_18472,N_13872,N_13053);
nand U18473 (N_18473,N_13953,N_14748);
nor U18474 (N_18474,N_12790,N_13139);
or U18475 (N_18475,N_14397,N_13931);
nor U18476 (N_18476,N_14803,N_13722);
or U18477 (N_18477,N_12667,N_15401);
nor U18478 (N_18478,N_14905,N_15615);
nor U18479 (N_18479,N_15287,N_15007);
or U18480 (N_18480,N_14511,N_15121);
or U18481 (N_18481,N_15260,N_14039);
nand U18482 (N_18482,N_13578,N_14415);
nand U18483 (N_18483,N_12966,N_14045);
and U18484 (N_18484,N_15464,N_12603);
nor U18485 (N_18485,N_14259,N_12776);
nor U18486 (N_18486,N_13588,N_14624);
nand U18487 (N_18487,N_13767,N_14786);
nor U18488 (N_18488,N_12903,N_12681);
nand U18489 (N_18489,N_15178,N_13238);
nor U18490 (N_18490,N_13887,N_15421);
nor U18491 (N_18491,N_13627,N_13009);
nand U18492 (N_18492,N_14589,N_14438);
nor U18493 (N_18493,N_13108,N_15010);
and U18494 (N_18494,N_15009,N_14995);
nand U18495 (N_18495,N_15503,N_14317);
or U18496 (N_18496,N_14591,N_14323);
or U18497 (N_18497,N_14589,N_13564);
nand U18498 (N_18498,N_15212,N_12984);
nor U18499 (N_18499,N_13872,N_15153);
nor U18500 (N_18500,N_15083,N_13588);
or U18501 (N_18501,N_13749,N_14370);
and U18502 (N_18502,N_15174,N_12778);
and U18503 (N_18503,N_13286,N_13473);
nand U18504 (N_18504,N_14281,N_12870);
nand U18505 (N_18505,N_15254,N_14187);
nand U18506 (N_18506,N_14919,N_13937);
nand U18507 (N_18507,N_12567,N_14680);
and U18508 (N_18508,N_14454,N_12951);
and U18509 (N_18509,N_15416,N_15005);
nand U18510 (N_18510,N_14390,N_14117);
and U18511 (N_18511,N_15046,N_13887);
and U18512 (N_18512,N_15066,N_14488);
or U18513 (N_18513,N_13778,N_14080);
nand U18514 (N_18514,N_12960,N_13724);
nand U18515 (N_18515,N_15167,N_12531);
and U18516 (N_18516,N_12777,N_14072);
and U18517 (N_18517,N_14773,N_13418);
nand U18518 (N_18518,N_15017,N_14088);
and U18519 (N_18519,N_13576,N_15235);
nand U18520 (N_18520,N_14166,N_12559);
nor U18521 (N_18521,N_15294,N_15535);
nand U18522 (N_18522,N_14587,N_14131);
nand U18523 (N_18523,N_14271,N_13060);
or U18524 (N_18524,N_13302,N_14584);
xnor U18525 (N_18525,N_13462,N_13477);
xnor U18526 (N_18526,N_15528,N_14052);
xor U18527 (N_18527,N_13088,N_15187);
or U18528 (N_18528,N_13102,N_13844);
nand U18529 (N_18529,N_14897,N_13897);
or U18530 (N_18530,N_13054,N_13871);
or U18531 (N_18531,N_14856,N_13147);
nand U18532 (N_18532,N_15069,N_12533);
and U18533 (N_18533,N_12624,N_14799);
or U18534 (N_18534,N_14013,N_13075);
or U18535 (N_18535,N_13813,N_13864);
nand U18536 (N_18536,N_13606,N_12717);
nand U18537 (N_18537,N_14533,N_13036);
nor U18538 (N_18538,N_15368,N_14760);
or U18539 (N_18539,N_13084,N_14980);
nor U18540 (N_18540,N_13584,N_14756);
nand U18541 (N_18541,N_13716,N_14115);
nor U18542 (N_18542,N_15327,N_14692);
and U18543 (N_18543,N_14820,N_14342);
nand U18544 (N_18544,N_14725,N_12597);
and U18545 (N_18545,N_13766,N_14841);
nor U18546 (N_18546,N_15084,N_13450);
or U18547 (N_18547,N_14401,N_14033);
nand U18548 (N_18548,N_13564,N_15124);
nor U18549 (N_18549,N_14319,N_13131);
nand U18550 (N_18550,N_13215,N_13415);
nand U18551 (N_18551,N_13856,N_12533);
or U18552 (N_18552,N_13101,N_14637);
and U18553 (N_18553,N_13528,N_15300);
nor U18554 (N_18554,N_12983,N_13077);
nor U18555 (N_18555,N_14242,N_13161);
or U18556 (N_18556,N_14136,N_13226);
nor U18557 (N_18557,N_15234,N_14608);
nor U18558 (N_18558,N_14795,N_15406);
nand U18559 (N_18559,N_13297,N_15493);
or U18560 (N_18560,N_13966,N_13726);
nand U18561 (N_18561,N_13414,N_14477);
or U18562 (N_18562,N_15564,N_13228);
nor U18563 (N_18563,N_15137,N_14223);
nor U18564 (N_18564,N_12859,N_14498);
and U18565 (N_18565,N_12520,N_13725);
and U18566 (N_18566,N_14821,N_12792);
nor U18567 (N_18567,N_13236,N_14324);
nor U18568 (N_18568,N_12719,N_12842);
nand U18569 (N_18569,N_15438,N_15091);
nor U18570 (N_18570,N_14395,N_14891);
and U18571 (N_18571,N_15272,N_13898);
or U18572 (N_18572,N_13263,N_12555);
xor U18573 (N_18573,N_14740,N_14181);
or U18574 (N_18574,N_12610,N_13429);
and U18575 (N_18575,N_14572,N_15559);
nand U18576 (N_18576,N_13147,N_14252);
nor U18577 (N_18577,N_14609,N_13647);
or U18578 (N_18578,N_12994,N_15490);
nand U18579 (N_18579,N_13660,N_14197);
or U18580 (N_18580,N_14900,N_13062);
nand U18581 (N_18581,N_12549,N_12619);
nand U18582 (N_18582,N_15044,N_14003);
and U18583 (N_18583,N_12940,N_14191);
nand U18584 (N_18584,N_13997,N_14380);
nand U18585 (N_18585,N_14563,N_13231);
xnor U18586 (N_18586,N_14743,N_13145);
and U18587 (N_18587,N_13334,N_13053);
nor U18588 (N_18588,N_13843,N_14775);
and U18589 (N_18589,N_13937,N_15524);
or U18590 (N_18590,N_14465,N_14183);
nand U18591 (N_18591,N_14165,N_15027);
or U18592 (N_18592,N_14675,N_12823);
xnor U18593 (N_18593,N_13716,N_13051);
and U18594 (N_18594,N_14501,N_14212);
xor U18595 (N_18595,N_14991,N_12964);
nand U18596 (N_18596,N_14602,N_14784);
and U18597 (N_18597,N_15366,N_13277);
xnor U18598 (N_18598,N_14710,N_13905);
nand U18599 (N_18599,N_14836,N_13072);
nor U18600 (N_18600,N_14171,N_13851);
xnor U18601 (N_18601,N_12632,N_15092);
nor U18602 (N_18602,N_12509,N_14241);
or U18603 (N_18603,N_15487,N_14445);
nand U18604 (N_18604,N_13108,N_15487);
xor U18605 (N_18605,N_14495,N_13177);
nor U18606 (N_18606,N_14289,N_13847);
and U18607 (N_18607,N_15279,N_13816);
and U18608 (N_18608,N_12960,N_14845);
nor U18609 (N_18609,N_15530,N_15120);
or U18610 (N_18610,N_14793,N_14994);
and U18611 (N_18611,N_14794,N_14780);
and U18612 (N_18612,N_13154,N_14961);
or U18613 (N_18613,N_14946,N_15091);
nor U18614 (N_18614,N_15578,N_15064);
or U18615 (N_18615,N_13577,N_13880);
xor U18616 (N_18616,N_13383,N_15123);
nor U18617 (N_18617,N_15021,N_13307);
or U18618 (N_18618,N_13809,N_15382);
nand U18619 (N_18619,N_15045,N_14909);
xor U18620 (N_18620,N_15459,N_13764);
or U18621 (N_18621,N_15562,N_14689);
nor U18622 (N_18622,N_12875,N_15147);
nand U18623 (N_18623,N_13991,N_14289);
nor U18624 (N_18624,N_14285,N_13594);
or U18625 (N_18625,N_12847,N_14827);
nand U18626 (N_18626,N_14959,N_15616);
xnor U18627 (N_18627,N_14959,N_12751);
nand U18628 (N_18628,N_13894,N_13553);
and U18629 (N_18629,N_12869,N_14057);
nor U18630 (N_18630,N_15265,N_12530);
nand U18631 (N_18631,N_15273,N_12621);
or U18632 (N_18632,N_12512,N_12983);
nor U18633 (N_18633,N_14597,N_13694);
nand U18634 (N_18634,N_15031,N_13154);
nand U18635 (N_18635,N_15133,N_13897);
nor U18636 (N_18636,N_12740,N_12897);
and U18637 (N_18637,N_14901,N_13604);
or U18638 (N_18638,N_14790,N_14289);
nor U18639 (N_18639,N_13453,N_14665);
nand U18640 (N_18640,N_12989,N_15251);
or U18641 (N_18641,N_12663,N_13355);
xor U18642 (N_18642,N_14882,N_13840);
nand U18643 (N_18643,N_13209,N_12574);
nand U18644 (N_18644,N_13353,N_14752);
nor U18645 (N_18645,N_15091,N_13974);
and U18646 (N_18646,N_15556,N_13992);
or U18647 (N_18647,N_13447,N_14628);
and U18648 (N_18648,N_13805,N_15547);
or U18649 (N_18649,N_15523,N_14338);
nand U18650 (N_18650,N_14288,N_12515);
nand U18651 (N_18651,N_14316,N_13756);
or U18652 (N_18652,N_13350,N_14275);
nand U18653 (N_18653,N_13974,N_14719);
and U18654 (N_18654,N_14266,N_13597);
nor U18655 (N_18655,N_13444,N_12863);
nand U18656 (N_18656,N_13717,N_13275);
nand U18657 (N_18657,N_13838,N_13703);
and U18658 (N_18658,N_15058,N_12672);
nor U18659 (N_18659,N_14452,N_13530);
nor U18660 (N_18660,N_14779,N_12724);
nor U18661 (N_18661,N_13283,N_14265);
and U18662 (N_18662,N_13465,N_13513);
and U18663 (N_18663,N_14586,N_15102);
nand U18664 (N_18664,N_12794,N_12693);
nand U18665 (N_18665,N_12591,N_12975);
nand U18666 (N_18666,N_13208,N_15252);
nor U18667 (N_18667,N_14066,N_13531);
xor U18668 (N_18668,N_14392,N_14586);
nand U18669 (N_18669,N_13538,N_13498);
nand U18670 (N_18670,N_14636,N_14254);
nand U18671 (N_18671,N_12827,N_13015);
or U18672 (N_18672,N_14636,N_14403);
or U18673 (N_18673,N_15373,N_13213);
or U18674 (N_18674,N_15354,N_14433);
xor U18675 (N_18675,N_13414,N_15583);
and U18676 (N_18676,N_13021,N_14876);
nand U18677 (N_18677,N_14685,N_15189);
nand U18678 (N_18678,N_13088,N_13636);
nand U18679 (N_18679,N_13517,N_14217);
or U18680 (N_18680,N_13039,N_12902);
nor U18681 (N_18681,N_12599,N_13802);
xor U18682 (N_18682,N_13630,N_14221);
or U18683 (N_18683,N_14758,N_13405);
or U18684 (N_18684,N_13948,N_13833);
and U18685 (N_18685,N_15169,N_13562);
or U18686 (N_18686,N_14280,N_13639);
and U18687 (N_18687,N_13623,N_15087);
or U18688 (N_18688,N_13163,N_14360);
nand U18689 (N_18689,N_14154,N_14075);
nand U18690 (N_18690,N_14631,N_14451);
and U18691 (N_18691,N_14972,N_14868);
or U18692 (N_18692,N_15585,N_14083);
or U18693 (N_18693,N_12550,N_13635);
nor U18694 (N_18694,N_15164,N_12812);
xor U18695 (N_18695,N_13184,N_12592);
or U18696 (N_18696,N_14630,N_15223);
or U18697 (N_18697,N_12579,N_14257);
and U18698 (N_18698,N_14085,N_15278);
nand U18699 (N_18699,N_14752,N_14302);
and U18700 (N_18700,N_12873,N_12666);
or U18701 (N_18701,N_14645,N_13268);
nor U18702 (N_18702,N_13277,N_13854);
nor U18703 (N_18703,N_14345,N_15383);
or U18704 (N_18704,N_13582,N_15048);
xor U18705 (N_18705,N_13384,N_14707);
and U18706 (N_18706,N_12690,N_12684);
nor U18707 (N_18707,N_13431,N_13447);
and U18708 (N_18708,N_14880,N_13565);
and U18709 (N_18709,N_12950,N_12955);
nor U18710 (N_18710,N_14318,N_13559);
nor U18711 (N_18711,N_14058,N_13686);
and U18712 (N_18712,N_14372,N_14875);
and U18713 (N_18713,N_12806,N_15061);
xnor U18714 (N_18714,N_12904,N_14566);
or U18715 (N_18715,N_14915,N_15042);
nand U18716 (N_18716,N_14706,N_13572);
nand U18717 (N_18717,N_13915,N_13801);
nand U18718 (N_18718,N_15559,N_14382);
nand U18719 (N_18719,N_14220,N_15484);
and U18720 (N_18720,N_14646,N_13812);
xor U18721 (N_18721,N_15317,N_13546);
and U18722 (N_18722,N_14628,N_12915);
and U18723 (N_18723,N_14385,N_14030);
or U18724 (N_18724,N_15336,N_14858);
xnor U18725 (N_18725,N_13618,N_12524);
or U18726 (N_18726,N_14017,N_14138);
or U18727 (N_18727,N_15256,N_13595);
nand U18728 (N_18728,N_13853,N_13367);
nor U18729 (N_18729,N_13293,N_13542);
nand U18730 (N_18730,N_14770,N_15199);
nor U18731 (N_18731,N_13508,N_13607);
or U18732 (N_18732,N_14590,N_14871);
xnor U18733 (N_18733,N_15283,N_14750);
or U18734 (N_18734,N_14538,N_13635);
nor U18735 (N_18735,N_13296,N_13567);
nand U18736 (N_18736,N_14292,N_13593);
or U18737 (N_18737,N_13528,N_14232);
or U18738 (N_18738,N_13781,N_15493);
and U18739 (N_18739,N_15545,N_12898);
nor U18740 (N_18740,N_15356,N_13014);
or U18741 (N_18741,N_13176,N_13640);
nor U18742 (N_18742,N_12612,N_13274);
and U18743 (N_18743,N_14497,N_12691);
and U18744 (N_18744,N_12983,N_13129);
nand U18745 (N_18745,N_13242,N_13925);
nor U18746 (N_18746,N_12740,N_12693);
and U18747 (N_18747,N_12642,N_15376);
nand U18748 (N_18748,N_14245,N_13066);
or U18749 (N_18749,N_12801,N_13443);
nor U18750 (N_18750,N_17265,N_16292);
or U18751 (N_18751,N_16821,N_15854);
nor U18752 (N_18752,N_16765,N_15715);
and U18753 (N_18753,N_15711,N_16317);
nand U18754 (N_18754,N_17044,N_16053);
or U18755 (N_18755,N_17455,N_18186);
nand U18756 (N_18756,N_17055,N_16699);
or U18757 (N_18757,N_17373,N_18104);
or U18758 (N_18758,N_18103,N_16008);
nand U18759 (N_18759,N_17108,N_18215);
nor U18760 (N_18760,N_17681,N_18107);
and U18761 (N_18761,N_17129,N_16675);
nor U18762 (N_18762,N_17920,N_17814);
xor U18763 (N_18763,N_16243,N_18260);
and U18764 (N_18764,N_17513,N_16749);
xnor U18765 (N_18765,N_18580,N_17783);
nor U18766 (N_18766,N_17665,N_18172);
nand U18767 (N_18767,N_18737,N_17710);
nor U18768 (N_18768,N_17519,N_17145);
nor U18769 (N_18769,N_16543,N_18445);
and U18770 (N_18770,N_16278,N_18306);
and U18771 (N_18771,N_17235,N_17307);
xor U18772 (N_18772,N_18018,N_17153);
xnor U18773 (N_18773,N_15996,N_16493);
and U18774 (N_18774,N_15877,N_15732);
nand U18775 (N_18775,N_18575,N_15763);
nand U18776 (N_18776,N_15923,N_16143);
and U18777 (N_18777,N_16003,N_15810);
nor U18778 (N_18778,N_18224,N_16990);
nand U18779 (N_18779,N_16970,N_18377);
and U18780 (N_18780,N_15859,N_16922);
and U18781 (N_18781,N_16721,N_18257);
and U18782 (N_18782,N_16342,N_17975);
and U18783 (N_18783,N_16147,N_16888);
or U18784 (N_18784,N_17175,N_17105);
nand U18785 (N_18785,N_15644,N_16792);
nand U18786 (N_18786,N_17002,N_16748);
and U18787 (N_18787,N_17270,N_16426);
or U18788 (N_18788,N_17994,N_16898);
or U18789 (N_18789,N_16827,N_16183);
nand U18790 (N_18790,N_16529,N_17887);
xor U18791 (N_18791,N_15892,N_16957);
nand U18792 (N_18792,N_18493,N_18508);
nor U18793 (N_18793,N_17817,N_17979);
nand U18794 (N_18794,N_17846,N_17532);
nand U18795 (N_18795,N_18604,N_17928);
nand U18796 (N_18796,N_18342,N_18500);
nor U18797 (N_18797,N_15856,N_17346);
and U18798 (N_18798,N_17323,N_17177);
xnor U18799 (N_18799,N_15782,N_16715);
and U18800 (N_18800,N_18683,N_18219);
and U18801 (N_18801,N_18139,N_15946);
and U18802 (N_18802,N_18328,N_17734);
nor U18803 (N_18803,N_18441,N_18541);
nand U18804 (N_18804,N_18372,N_15991);
or U18805 (N_18805,N_16286,N_16691);
nor U18806 (N_18806,N_17220,N_17913);
or U18807 (N_18807,N_16073,N_17892);
nand U18808 (N_18808,N_16451,N_18271);
nand U18809 (N_18809,N_17831,N_17308);
and U18810 (N_18810,N_16343,N_15640);
nor U18811 (N_18811,N_17758,N_16218);
nor U18812 (N_18812,N_16519,N_16695);
and U18813 (N_18813,N_18557,N_17878);
nand U18814 (N_18814,N_17061,N_17049);
and U18815 (N_18815,N_17833,N_17964);
or U18816 (N_18816,N_16461,N_18705);
nand U18817 (N_18817,N_15866,N_16945);
and U18818 (N_18818,N_16518,N_16041);
xor U18819 (N_18819,N_18221,N_16639);
or U18820 (N_18820,N_17343,N_18619);
or U18821 (N_18821,N_17406,N_16573);
and U18822 (N_18822,N_16754,N_16714);
nor U18823 (N_18823,N_18471,N_16668);
and U18824 (N_18824,N_16681,N_16415);
xor U18825 (N_18825,N_18533,N_17868);
or U18826 (N_18826,N_16522,N_17836);
nor U18827 (N_18827,N_16058,N_16804);
and U18828 (N_18828,N_16410,N_17171);
and U18829 (N_18829,N_18719,N_17355);
nand U18830 (N_18830,N_17820,N_16188);
and U18831 (N_18831,N_17518,N_17938);
nand U18832 (N_18832,N_16967,N_15950);
xor U18833 (N_18833,N_18634,N_18448);
or U18834 (N_18834,N_15900,N_15825);
or U18835 (N_18835,N_16829,N_16021);
and U18836 (N_18836,N_15977,N_18243);
or U18837 (N_18837,N_17617,N_17179);
nor U18838 (N_18838,N_16732,N_16355);
and U18839 (N_18839,N_18661,N_17219);
and U18840 (N_18840,N_17349,N_16806);
or U18841 (N_18841,N_17637,N_18147);
nor U18842 (N_18842,N_16365,N_16197);
nor U18843 (N_18843,N_17092,N_15673);
xor U18844 (N_18844,N_15933,N_17239);
and U18845 (N_18845,N_18376,N_16880);
nor U18846 (N_18846,N_16788,N_18418);
or U18847 (N_18847,N_17487,N_17863);
nor U18848 (N_18848,N_17860,N_17223);
xor U18849 (N_18849,N_18483,N_16348);
nand U18850 (N_18850,N_16314,N_16448);
and U18851 (N_18851,N_17871,N_16986);
nor U18852 (N_18852,N_17752,N_17114);
nand U18853 (N_18853,N_17340,N_16545);
and U18854 (N_18854,N_17301,N_18343);
and U18855 (N_18855,N_18542,N_17855);
nand U18856 (N_18856,N_17462,N_17038);
and U18857 (N_18857,N_18280,N_18349);
nor U18858 (N_18858,N_18539,N_16574);
and U18859 (N_18859,N_16981,N_15981);
nand U18860 (N_18860,N_16859,N_18276);
nand U18861 (N_18861,N_16568,N_15738);
xor U18862 (N_18862,N_16293,N_15742);
nand U18863 (N_18863,N_15870,N_16747);
nor U18864 (N_18864,N_17150,N_17800);
nor U18865 (N_18865,N_16395,N_18430);
nor U18866 (N_18866,N_17312,N_18347);
nand U18867 (N_18867,N_17375,N_18019);
or U18868 (N_18868,N_16905,N_17656);
and U18869 (N_18869,N_17910,N_17282);
or U18870 (N_18870,N_17001,N_18509);
and U18871 (N_18871,N_17254,N_18436);
nand U18872 (N_18872,N_18151,N_17216);
nand U18873 (N_18873,N_15997,N_18395);
nor U18874 (N_18874,N_17821,N_16576);
and U18875 (N_18875,N_17309,N_17715);
xor U18876 (N_18876,N_15862,N_16347);
nor U18877 (N_18877,N_17012,N_17556);
nor U18878 (N_18878,N_17830,N_17537);
and U18879 (N_18879,N_15941,N_16995);
and U18880 (N_18880,N_18079,N_17670);
or U18881 (N_18881,N_18292,N_17023);
and U18882 (N_18882,N_17541,N_16787);
nand U18883 (N_18883,N_18022,N_18055);
nor U18884 (N_18884,N_16835,N_16614);
nor U18885 (N_18885,N_15757,N_16130);
xor U18886 (N_18886,N_15649,N_15826);
nor U18887 (N_18887,N_16264,N_17588);
or U18888 (N_18888,N_17377,N_16772);
nand U18889 (N_18889,N_16737,N_17799);
and U18890 (N_18890,N_16902,N_16036);
or U18891 (N_18891,N_18077,N_17545);
or U18892 (N_18892,N_17082,N_18248);
nor U18893 (N_18893,N_16931,N_17371);
and U18894 (N_18894,N_18563,N_16359);
nor U18895 (N_18895,N_18529,N_16734);
nor U18896 (N_18896,N_18236,N_18031);
nor U18897 (N_18897,N_17087,N_17168);
xnor U18898 (N_18898,N_17768,N_18053);
or U18899 (N_18899,N_17692,N_17492);
nand U18900 (N_18900,N_18339,N_18534);
nand U18901 (N_18901,N_18459,N_18318);
nand U18902 (N_18902,N_18703,N_16217);
xnor U18903 (N_18903,N_17891,N_18662);
and U18904 (N_18904,N_16839,N_16066);
or U18905 (N_18905,N_18733,N_17350);
nand U18906 (N_18906,N_18262,N_17103);
nor U18907 (N_18907,N_18222,N_18659);
nor U18908 (N_18908,N_16273,N_18470);
nand U18909 (N_18909,N_18621,N_16467);
and U18910 (N_18910,N_16151,N_16024);
nor U18911 (N_18911,N_16847,N_15984);
nand U18912 (N_18912,N_15967,N_18142);
xor U18913 (N_18913,N_17929,N_16156);
and U18914 (N_18914,N_16775,N_15785);
nand U18915 (N_18915,N_17304,N_18497);
and U18916 (N_18916,N_18253,N_18013);
and U18917 (N_18917,N_16297,N_15897);
or U18918 (N_18918,N_16165,N_18289);
and U18919 (N_18919,N_15724,N_16756);
nor U18920 (N_18920,N_18035,N_18657);
and U18921 (N_18921,N_16996,N_18614);
xor U18922 (N_18922,N_17744,N_17751);
and U18923 (N_18923,N_16688,N_16299);
nand U18924 (N_18924,N_16750,N_17077);
or U18925 (N_18925,N_16527,N_16113);
nand U18926 (N_18926,N_17682,N_15807);
and U18927 (N_18927,N_18281,N_17774);
or U18928 (N_18928,N_17969,N_18417);
and U18929 (N_18929,N_17428,N_16603);
and U18930 (N_18930,N_15894,N_17008);
nor U18931 (N_18931,N_18279,N_16540);
nand U18932 (N_18932,N_17828,N_16776);
and U18933 (N_18933,N_15822,N_16846);
nor U18934 (N_18934,N_17769,N_17474);
or U18935 (N_18935,N_18184,N_17629);
nor U18936 (N_18936,N_16369,N_17745);
nor U18937 (N_18937,N_18736,N_18071);
and U18938 (N_18938,N_17066,N_16917);
and U18939 (N_18939,N_15809,N_16757);
or U18940 (N_18940,N_16163,N_17847);
nor U18941 (N_18941,N_16785,N_17740);
nor U18942 (N_18942,N_16020,N_18105);
or U18943 (N_18943,N_16731,N_16786);
or U18944 (N_18944,N_16488,N_17865);
xnor U18945 (N_18945,N_18299,N_15642);
or U18946 (N_18946,N_15638,N_16660);
and U18947 (N_18947,N_17251,N_16943);
nand U18948 (N_18948,N_18605,N_18729);
nand U18949 (N_18949,N_17596,N_15920);
and U18950 (N_18950,N_17572,N_18679);
and U18951 (N_18951,N_16248,N_17881);
or U18952 (N_18952,N_16659,N_15794);
or U18953 (N_18953,N_16009,N_16795);
nor U18954 (N_18954,N_16896,N_16012);
or U18955 (N_18955,N_18331,N_18183);
or U18956 (N_18956,N_16629,N_18370);
nand U18957 (N_18957,N_16865,N_16242);
nand U18958 (N_18958,N_16051,N_15907);
or U18959 (N_18959,N_18210,N_17542);
or U18960 (N_18960,N_18261,N_17527);
or U18961 (N_18961,N_17595,N_18157);
nor U18962 (N_18962,N_17586,N_16592);
xnor U18963 (N_18963,N_18174,N_16532);
nor U18964 (N_18964,N_16949,N_16460);
and U18965 (N_18965,N_15998,N_16298);
nand U18966 (N_18966,N_17845,N_18389);
or U18967 (N_18967,N_16126,N_18636);
xor U18968 (N_18968,N_16812,N_17893);
nand U18969 (N_18969,N_16239,N_16594);
nand U18970 (N_18970,N_17227,N_16068);
nor U18971 (N_18971,N_17389,N_17628);
nand U18972 (N_18972,N_17658,N_17674);
nand U18973 (N_18973,N_16762,N_15974);
and U18974 (N_18974,N_16857,N_17784);
xnor U18975 (N_18975,N_16071,N_17042);
xor U18976 (N_18976,N_18622,N_16475);
nand U18977 (N_18977,N_18660,N_16977);
nand U18978 (N_18978,N_17361,N_17184);
or U18979 (N_18979,N_18173,N_17719);
and U18980 (N_18980,N_18738,N_18096);
or U18981 (N_18981,N_15883,N_17263);
nor U18982 (N_18982,N_16556,N_16251);
and U18983 (N_18983,N_15891,N_18066);
or U18984 (N_18984,N_16627,N_15949);
or U18985 (N_18985,N_18642,N_18411);
or U18986 (N_18986,N_18637,N_18199);
and U18987 (N_18987,N_15820,N_16958);
xnor U18988 (N_18988,N_16149,N_16559);
or U18989 (N_18989,N_16083,N_17829);
and U18990 (N_18990,N_18405,N_16667);
nor U18991 (N_18991,N_18327,N_15700);
nand U18992 (N_18992,N_18582,N_18064);
nand U18993 (N_18993,N_17151,N_18536);
xnor U18994 (N_18994,N_17456,N_16032);
nand U18995 (N_18995,N_16483,N_18295);
xor U18996 (N_18996,N_17224,N_16783);
or U18997 (N_18997,N_17449,N_16005);
nand U18998 (N_18998,N_18177,N_18695);
and U18999 (N_18999,N_17515,N_18698);
nor U19000 (N_19000,N_15966,N_17926);
and U19001 (N_19001,N_16712,N_17050);
or U19002 (N_19002,N_15698,N_17030);
xor U19003 (N_19003,N_17159,N_16878);
nand U19004 (N_19004,N_18095,N_17494);
or U19005 (N_19005,N_16457,N_15959);
or U19006 (N_19006,N_15741,N_16561);
nor U19007 (N_19007,N_18606,N_17621);
xor U19008 (N_19008,N_17423,N_17712);
and U19009 (N_19009,N_16599,N_17507);
xnor U19010 (N_19010,N_18348,N_16102);
or U19011 (N_19011,N_17036,N_16209);
nor U19012 (N_19012,N_17512,N_15861);
nand U19013 (N_19013,N_17269,N_16136);
nand U19014 (N_19014,N_17095,N_18190);
and U19015 (N_19015,N_16105,N_17260);
nor U19016 (N_19016,N_17411,N_17936);
and U19017 (N_19017,N_17877,N_17508);
or U19018 (N_19018,N_16796,N_17037);
or U19019 (N_19019,N_17089,N_15683);
nor U19020 (N_19020,N_17679,N_16729);
or U19021 (N_19021,N_17162,N_15725);
or U19022 (N_19022,N_18450,N_17286);
nand U19023 (N_19023,N_18531,N_18152);
and U19024 (N_19024,N_16399,N_17320);
and U19025 (N_19025,N_18048,N_17345);
nor U19026 (N_19026,N_17778,N_18340);
or U19027 (N_19027,N_18229,N_17854);
nand U19028 (N_19028,N_16307,N_16572);
nand U19029 (N_19029,N_16541,N_16505);
nand U19030 (N_19030,N_17869,N_18181);
or U19031 (N_19031,N_17764,N_16368);
nand U19032 (N_19032,N_16429,N_16707);
nand U19033 (N_19033,N_18457,N_17400);
nor U19034 (N_19034,N_15790,N_17464);
nor U19035 (N_19035,N_17732,N_18093);
or U19036 (N_19036,N_18523,N_15918);
nor U19037 (N_19037,N_17544,N_15654);
nor U19038 (N_19038,N_17170,N_17000);
or U19039 (N_19039,N_18629,N_16418);
or U19040 (N_19040,N_16863,N_16887);
nor U19041 (N_19041,N_17683,N_18685);
xor U19042 (N_19042,N_16075,N_18435);
or U19043 (N_19043,N_17660,N_16271);
and U19044 (N_19044,N_17017,N_16029);
or U19045 (N_19045,N_16081,N_18643);
and U19046 (N_19046,N_15818,N_15860);
or U19047 (N_19047,N_17738,N_17761);
nor U19048 (N_19048,N_16980,N_16069);
xor U19049 (N_19049,N_15761,N_16442);
nor U19050 (N_19050,N_18029,N_16496);
and U19051 (N_19051,N_18314,N_16841);
and U19052 (N_19052,N_15786,N_18119);
and U19053 (N_19053,N_16112,N_16685);
nand U19054 (N_19054,N_18598,N_17779);
nand U19055 (N_19055,N_15755,N_17480);
nand U19056 (N_19056,N_16890,N_15645);
and U19057 (N_19057,N_17046,N_18042);
or U19058 (N_19058,N_17298,N_18240);
xor U19059 (N_19059,N_16489,N_17790);
and U19060 (N_19060,N_17146,N_17634);
nand U19061 (N_19061,N_16913,N_18136);
and U19062 (N_19062,N_17627,N_17991);
nor U19063 (N_19063,N_18625,N_17294);
and U19064 (N_19064,N_15789,N_17957);
nor U19065 (N_19065,N_15960,N_16587);
xnor U19066 (N_19066,N_16553,N_16172);
nor U19067 (N_19067,N_17945,N_18302);
nor U19068 (N_19068,N_15922,N_17798);
and U19069 (N_19069,N_18036,N_18412);
or U19070 (N_19070,N_15871,N_16909);
xnor U19071 (N_19071,N_15727,N_17873);
nor U19072 (N_19072,N_16015,N_18034);
and U19073 (N_19073,N_16588,N_18016);
xnor U19074 (N_19074,N_18192,N_17217);
and U19075 (N_19075,N_17385,N_16868);
xnor U19076 (N_19076,N_16598,N_17249);
and U19077 (N_19077,N_16246,N_16413);
nand U19078 (N_19078,N_16612,N_16345);
nand U19079 (N_19079,N_15989,N_18682);
nand U19080 (N_19080,N_15844,N_17574);
xor U19081 (N_19081,N_16692,N_15952);
or U19082 (N_19082,N_16915,N_16414);
nand U19083 (N_19083,N_16974,N_18701);
or U19084 (N_19084,N_18658,N_16928);
nand U19085 (N_19085,N_18713,N_18081);
xor U19086 (N_19086,N_18148,N_18454);
nand U19087 (N_19087,N_18254,N_18266);
nor U19088 (N_19088,N_17418,N_16690);
and U19089 (N_19089,N_16296,N_15913);
or U19090 (N_19090,N_15679,N_17052);
xnor U19091 (N_19091,N_16316,N_17927);
and U19092 (N_19092,N_18004,N_17376);
and U19093 (N_19093,N_16159,N_16708);
xnor U19094 (N_19094,N_18649,N_17404);
or U19095 (N_19095,N_16830,N_18021);
and U19096 (N_19096,N_17906,N_16050);
nand U19097 (N_19097,N_18425,N_18490);
and U19098 (N_19098,N_16084,N_18489);
nor U19099 (N_19099,N_17677,N_17959);
or U19100 (N_19100,N_17721,N_18562);
nor U19101 (N_19101,N_16118,N_16774);
or U19102 (N_19102,N_18728,N_17417);
and U19103 (N_19103,N_16164,N_18294);
or U19104 (N_19104,N_17491,N_18718);
nand U19105 (N_19105,N_15695,N_17231);
nand U19106 (N_19106,N_15756,N_17398);
or U19107 (N_19107,N_18206,N_17693);
nor U19108 (N_19108,N_18163,N_17198);
nand U19109 (N_19109,N_15955,N_16360);
and U19110 (N_19110,N_16648,N_17576);
nand U19111 (N_19111,N_17668,N_16027);
and U19112 (N_19112,N_18125,N_17652);
nand U19113 (N_19113,N_16910,N_16508);
and U19114 (N_19114,N_16760,N_17318);
nor U19115 (N_19115,N_16212,N_18491);
and U19116 (N_19116,N_17787,N_17181);
and U19117 (N_19117,N_18403,N_16422);
nand U19118 (N_19118,N_17946,N_18707);
and U19119 (N_19119,N_15689,N_15690);
xnor U19120 (N_19120,N_15990,N_16528);
nand U19121 (N_19121,N_15863,N_15963);
nor U19122 (N_19122,N_16304,N_17930);
and U19123 (N_19123,N_16144,N_16644);
nor U19124 (N_19124,N_17422,N_16275);
nor U19125 (N_19125,N_17180,N_16727);
or U19126 (N_19126,N_18650,N_18486);
and U19127 (N_19127,N_17438,N_17594);
nor U19128 (N_19128,N_18118,N_17503);
and U19129 (N_19129,N_17288,N_15704);
and U19130 (N_19130,N_17954,N_16790);
or U19131 (N_19131,N_15935,N_18182);
nor U19132 (N_19132,N_18058,N_15671);
nand U19133 (N_19133,N_17033,N_18715);
or U19134 (N_19134,N_16769,N_16551);
and U19135 (N_19135,N_17671,N_18724);
or U19136 (N_19136,N_18675,N_16019);
and U19137 (N_19137,N_17213,N_16434);
nor U19138 (N_19138,N_15992,N_15694);
or U19139 (N_19139,N_17070,N_18185);
nor U19140 (N_19140,N_16499,N_17993);
nor U19141 (N_19141,N_16595,N_17702);
xor U19142 (N_19142,N_16552,N_16398);
nand U19143 (N_19143,N_16613,N_18002);
nor U19144 (N_19144,N_17923,N_17718);
nand U19145 (N_19145,N_16641,N_16745);
nand U19146 (N_19146,N_17148,N_17357);
or U19147 (N_19147,N_17090,N_16874);
nor U19148 (N_19148,N_17965,N_16328);
or U19149 (N_19149,N_16454,N_16570);
and U19150 (N_19150,N_17447,N_16184);
nand U19151 (N_19151,N_18160,N_16103);
nor U19152 (N_19152,N_17981,N_17207);
nor U19153 (N_19153,N_16263,N_15627);
and U19154 (N_19154,N_16070,N_17773);
and U19155 (N_19155,N_17540,N_18460);
and U19156 (N_19156,N_16131,N_17673);
or U19157 (N_19157,N_16884,N_17822);
or U19158 (N_19158,N_16471,N_17706);
nor U19159 (N_19159,N_17604,N_16617);
nor U19160 (N_19160,N_17086,N_16975);
or U19161 (N_19161,N_16352,N_17306);
or U19162 (N_19162,N_17238,N_16445);
nor U19163 (N_19163,N_18094,N_16274);
nand U19164 (N_19164,N_18218,N_18068);
and U19165 (N_19165,N_18646,N_16329);
xor U19166 (N_19166,N_15719,N_18524);
nor U19167 (N_19167,N_17533,N_17463);
or U19168 (N_19168,N_16386,N_18145);
and U19169 (N_19169,N_18566,N_17395);
and U19170 (N_19170,N_18296,N_17071);
and U19171 (N_19171,N_18083,N_16767);
or U19172 (N_19172,N_16632,N_17996);
xnor U19173 (N_19173,N_18012,N_16989);
and U19174 (N_19174,N_17293,N_17021);
or U19175 (N_19175,N_18739,N_18074);
or U19176 (N_19176,N_16336,N_16906);
xor U19177 (N_19177,N_18242,N_18478);
or U19178 (N_19178,N_17290,N_17497);
xor U19179 (N_19179,N_16844,N_16758);
nor U19180 (N_19180,N_16230,N_16831);
and U19181 (N_19181,N_16052,N_17765);
and U19182 (N_19182,N_16826,N_17210);
nor U19183 (N_19183,N_16635,N_17128);
nand U19184 (N_19184,N_17642,N_18134);
or U19185 (N_19185,N_15655,N_17059);
nand U19186 (N_19186,N_18278,N_16309);
or U19187 (N_19187,N_18080,N_16375);
and U19188 (N_19188,N_17484,N_16214);
and U19189 (N_19189,N_18426,N_18416);
nand U19190 (N_19190,N_18421,N_16807);
and U19191 (N_19191,N_16881,N_18522);
nor U19192 (N_19192,N_17362,N_18609);
xor U19193 (N_19193,N_16301,N_15857);
nor U19194 (N_19194,N_17748,N_18298);
or U19195 (N_19195,N_15767,N_15819);
or U19196 (N_19196,N_15969,N_15985);
xnor U19197 (N_19197,N_15631,N_18267);
or U19198 (N_19198,N_18284,N_17026);
xnor U19199 (N_19199,N_18115,N_17949);
or U19200 (N_19200,N_15657,N_16222);
or U19201 (N_19201,N_17788,N_17454);
nor U19202 (N_19202,N_17669,N_17271);
nand U19203 (N_19203,N_18131,N_18312);
or U19204 (N_19204,N_15751,N_17027);
nor U19205 (N_19205,N_17546,N_18390);
nand U19206 (N_19206,N_17248,N_16033);
and U19207 (N_19207,N_16190,N_18513);
and U19208 (N_19208,N_17164,N_16971);
and U19209 (N_19209,N_15916,N_17316);
nor U19210 (N_19210,N_15867,N_17025);
or U19211 (N_19211,N_18357,N_16268);
xor U19212 (N_19212,N_16199,N_18571);
and U19213 (N_19213,N_15958,N_17502);
and U19214 (N_19214,N_17908,N_16463);
nor U19215 (N_19215,N_16179,N_18359);
nor U19216 (N_19216,N_16104,N_17205);
nor U19217 (N_19217,N_16408,N_15869);
or U19218 (N_19218,N_17880,N_17195);
nor U19219 (N_19219,N_17427,N_16057);
and U19220 (N_19220,N_17470,N_16167);
xnor U19221 (N_19221,N_16658,N_18256);
nand U19222 (N_19222,N_18585,N_17971);
or U19223 (N_19223,N_17559,N_18545);
nand U19224 (N_19224,N_16446,N_17172);
and U19225 (N_19225,N_16469,N_17522);
nand U19226 (N_19226,N_17232,N_16261);
or U19227 (N_19227,N_18102,N_17757);
nor U19228 (N_19228,N_16140,N_16723);
and U19229 (N_19229,N_16099,N_16139);
xor U19230 (N_19230,N_17735,N_18270);
nand U19231 (N_19231,N_18400,N_16649);
and U19232 (N_19232,N_18439,N_16662);
nand U19233 (N_19233,N_15729,N_18335);
and U19234 (N_19234,N_16120,N_16349);
nor U19235 (N_19235,N_16354,N_17806);
and U19236 (N_19236,N_18717,N_16206);
and U19237 (N_19237,N_16082,N_16150);
nor U19238 (N_19238,N_16982,N_18154);
or U19239 (N_19239,N_15639,N_17348);
and U19240 (N_19240,N_15678,N_16280);
or U19241 (N_19241,N_17529,N_16575);
xor U19242 (N_19242,N_17912,N_18607);
nor U19243 (N_19243,N_17775,N_15750);
or U19244 (N_19244,N_17818,N_16877);
nand U19245 (N_19245,N_15972,N_18656);
or U19246 (N_19246,N_17193,N_18087);
nor U19247 (N_19247,N_18462,N_17112);
nand U19248 (N_19248,N_16655,N_17713);
or U19249 (N_19249,N_16234,N_16929);
nor U19250 (N_19250,N_18166,N_18503);
nand U19251 (N_19251,N_16391,N_17281);
nor U19252 (N_19252,N_18409,N_18225);
xnor U19253 (N_19253,N_17486,N_17552);
and U19254 (N_19254,N_16064,N_16236);
or U19255 (N_19255,N_18211,N_17756);
nand U19256 (N_19256,N_17022,N_16432);
nor U19257 (N_19257,N_17875,N_16135);
or U19258 (N_19258,N_17606,N_16702);
xor U19259 (N_19259,N_16738,N_16327);
nand U19260 (N_19260,N_17292,N_15656);
nor U19261 (N_19261,N_18355,N_17941);
nand U19262 (N_19262,N_17514,N_16262);
and U19263 (N_19263,N_18516,N_15708);
nor U19264 (N_19264,N_18525,N_18250);
nand U19265 (N_19265,N_16312,N_18162);
xnor U19266 (N_19266,N_17565,N_17152);
nor U19267 (N_19267,N_16773,N_17018);
nand U19268 (N_19268,N_15968,N_17253);
nand U19269 (N_19269,N_17261,N_16946);
and U19270 (N_19270,N_17394,N_16646);
nand U19271 (N_19271,N_17791,N_16152);
and U19272 (N_19272,N_16194,N_15864);
and U19273 (N_19273,N_16193,N_16539);
or U19274 (N_19274,N_17085,N_16417);
and U19275 (N_19275,N_16564,N_17097);
nand U19276 (N_19276,N_16610,N_18671);
nor U19277 (N_19277,N_16728,N_18749);
or U19278 (N_19278,N_15791,N_17344);
or U19279 (N_19279,N_16498,N_18602);
or U19280 (N_19280,N_17897,N_15722);
xnor U19281 (N_19281,N_16963,N_18721);
or U19282 (N_19282,N_17183,N_15976);
or U19283 (N_19283,N_17431,N_15728);
xor U19284 (N_19284,N_17084,N_16578);
and U19285 (N_19285,N_17113,N_18052);
nand U19286 (N_19286,N_17214,N_16889);
nor U19287 (N_19287,N_17460,N_17551);
and U19288 (N_19288,N_17031,N_18601);
xnor U19289 (N_19289,N_16824,N_17974);
nor U19290 (N_19290,N_17924,N_18114);
nor U19291 (N_19291,N_15910,N_17384);
or U19292 (N_19292,N_18677,N_15927);
or U19293 (N_19293,N_17130,N_16621);
or U19294 (N_19294,N_16208,N_15834);
xnor U19295 (N_19295,N_17367,N_18220);
nand U19296 (N_19296,N_16438,N_15780);
xnor U19297 (N_19297,N_17663,N_17351);
or U19298 (N_19298,N_16921,N_16536);
or U19299 (N_19299,N_17743,N_16110);
or U19300 (N_19300,N_18008,N_17624);
nor U19301 (N_19301,N_16856,N_18692);
nand U19302 (N_19302,N_17792,N_17136);
nand U19303 (N_19303,N_17589,N_16547);
nand U19304 (N_19304,N_18710,N_16870);
nor U19305 (N_19305,N_15664,N_18325);
nor U19306 (N_19306,N_17358,N_15630);
or U19307 (N_19307,N_16622,N_16866);
or U19308 (N_19308,N_15957,N_17646);
or U19309 (N_19309,N_18203,N_18383);
or U19310 (N_19310,N_17319,N_17940);
nor U19311 (N_19311,N_17921,N_16801);
nor U19312 (N_19312,N_15886,N_16755);
nor U19313 (N_19313,N_16378,N_15693);
or U19314 (N_19314,N_18442,N_15954);
or U19315 (N_19315,N_16407,N_18526);
and U19316 (N_19316,N_17703,N_16011);
and U19317 (N_19317,N_15801,N_17158);
or U19318 (N_19318,N_18101,N_17325);
nand U19319 (N_19319,N_16596,N_15999);
or U19320 (N_19320,N_15709,N_16406);
nor U19321 (N_19321,N_16470,N_16249);
nor U19322 (N_19322,N_18309,N_17688);
or U19323 (N_19323,N_15939,N_16441);
and U19324 (N_19324,N_16148,N_15851);
and U19325 (N_19325,N_16606,N_18039);
nand U19326 (N_19326,N_17689,N_16340);
nor U19327 (N_19327,N_17610,N_16999);
or U19328 (N_19328,N_16953,N_16367);
or U19329 (N_19329,N_18086,N_17888);
or U19330 (N_19330,N_18530,N_15736);
nor U19331 (N_19331,N_18456,N_17083);
nand U19332 (N_19332,N_18444,N_17562);
nand U19333 (N_19333,N_15815,N_16843);
or U19334 (N_19334,N_18097,N_17909);
and U19335 (N_19335,N_17063,N_17832);
or U19336 (N_19336,N_17573,N_15914);
or U19337 (N_19337,N_16972,N_17206);
or U19338 (N_19338,N_17771,N_18560);
nand U19339 (N_19339,N_16224,N_17980);
nor U19340 (N_19340,N_16630,N_18124);
or U19341 (N_19341,N_17616,N_18578);
or U19342 (N_19342,N_16624,N_18747);
and U19343 (N_19343,N_17415,N_17997);
nand U19344 (N_19344,N_15665,N_16607);
nor U19345 (N_19345,N_15769,N_16031);
nor U19346 (N_19346,N_18088,N_17433);
nor U19347 (N_19347,N_18090,N_17737);
or U19348 (N_19348,N_16512,N_17274);
nor U19349 (N_19349,N_15872,N_18615);
xnor U19350 (N_19350,N_16948,N_18482);
or U19351 (N_19351,N_17468,N_17388);
or U19352 (N_19352,N_18406,N_18123);
nand U19353 (N_19353,N_18334,N_15707);
and U19354 (N_19354,N_16531,N_17592);
nand U19355 (N_19355,N_15912,N_16014);
xor U19356 (N_19356,N_16816,N_16371);
nor U19357 (N_19357,N_17283,N_16397);
and U19358 (N_19358,N_18479,N_18583);
xor U19359 (N_19359,N_16238,N_17419);
nand U19360 (N_19360,N_18251,N_17747);
or U19361 (N_19361,N_16191,N_16108);
nand U19362 (N_19362,N_16048,N_15658);
nor U19363 (N_19363,N_17125,N_16959);
nand U19364 (N_19364,N_18408,N_17032);
nor U19365 (N_19365,N_16026,N_17165);
or U19366 (N_19366,N_18399,N_16363);
or U19367 (N_19367,N_16952,N_15758);
or U19368 (N_19368,N_17983,N_17905);
nand U19369 (N_19369,N_16666,N_17709);
nand U19370 (N_19370,N_17287,N_17074);
nor U19371 (N_19371,N_17899,N_15687);
nand U19372 (N_19372,N_17313,N_16382);
nor U19373 (N_19373,N_17228,N_18388);
nor U19374 (N_19374,N_16894,N_17440);
xor U19375 (N_19375,N_17155,N_17958);
nor U19376 (N_19376,N_16683,N_16653);
xor U19377 (N_19377,N_17808,N_15848);
or U19378 (N_19378,N_15936,N_17583);
or U19379 (N_19379,N_17127,N_18492);
or U19380 (N_19380,N_16387,N_16513);
nor U19381 (N_19381,N_15797,N_17619);
nand U19382 (N_19382,N_17843,N_18098);
nor U19383 (N_19383,N_17230,N_16942);
xnor U19384 (N_19384,N_18742,N_18555);
nor U19385 (N_19385,N_18063,N_17222);
xor U19386 (N_19386,N_16951,N_15651);
and U19387 (N_19387,N_17901,N_15944);
nor U19388 (N_19388,N_16993,N_18075);
or U19389 (N_19389,N_16007,N_18363);
nor U19390 (N_19390,N_18073,N_17566);
or U19391 (N_19391,N_18005,N_16997);
or U19392 (N_19392,N_16169,N_16341);
and U19393 (N_19393,N_18085,N_18393);
nor U19394 (N_19394,N_17795,N_15926);
nand U19395 (N_19395,N_15779,N_17457);
xor U19396 (N_19396,N_17708,N_16034);
and U19397 (N_19397,N_17133,N_17276);
nor U19398 (N_19398,N_18702,N_16231);
and U19399 (N_19399,N_17215,N_17311);
and U19400 (N_19400,N_18252,N_18392);
xor U19401 (N_19401,N_17884,N_18538);
and U19402 (N_19402,N_16563,N_18588);
xnor U19403 (N_19403,N_16569,N_17056);
nor U19404 (N_19404,N_18589,N_17203);
nand U19405 (N_19405,N_16674,N_17387);
and U19406 (N_19406,N_17973,N_15833);
nand U19407 (N_19407,N_16439,N_17684);
nand U19408 (N_19408,N_18431,N_15669);
and U19409 (N_19409,N_16751,N_15803);
nand U19410 (N_19410,N_15684,N_15938);
nand U19411 (N_19411,N_16704,N_16916);
nand U19412 (N_19412,N_17401,N_17020);
and U19413 (N_19413,N_15928,N_18324);
nor U19414 (N_19414,N_17317,N_16615);
nand U19415 (N_19415,N_16459,N_15643);
nand U19416 (N_19416,N_17553,N_17520);
nand U19417 (N_19417,N_17898,N_18572);
nor U19418 (N_19418,N_16250,N_17856);
nor U19419 (N_19419,N_17644,N_16586);
nor U19420 (N_19420,N_16601,N_15768);
nor U19421 (N_19421,N_17720,N_17612);
and U19422 (N_19422,N_16046,N_17439);
xnor U19423 (N_19423,N_16049,N_15983);
nand U19424 (N_19424,N_16591,N_18089);
nor U19425 (N_19425,N_16456,N_17436);
and U19426 (N_19426,N_16247,N_17984);
nor U19427 (N_19427,N_17166,N_16710);
or U19428 (N_19428,N_17733,N_17332);
or U19429 (N_19429,N_18310,N_17243);
and U19430 (N_19430,N_17391,N_17648);
xnor U19431 (N_19431,N_18504,N_16279);
nand U19432 (N_19432,N_15971,N_17755);
nand U19433 (N_19433,N_16554,N_18099);
and U19434 (N_19434,N_16364,N_15668);
and U19435 (N_19435,N_17465,N_16828);
or U19436 (N_19436,N_17707,N_15762);
or U19437 (N_19437,N_16966,N_17521);
and U19438 (N_19438,N_18543,N_16383);
nand U19439 (N_19439,N_17711,N_18477);
or U19440 (N_19440,N_17339,N_17914);
and U19441 (N_19441,N_16092,N_18237);
nor U19442 (N_19442,N_17850,N_16926);
nor U19443 (N_19443,N_16736,N_18593);
xnor U19444 (N_19444,N_16813,N_18367);
nand U19445 (N_19445,N_16852,N_17730);
and U19446 (N_19446,N_16252,N_18263);
nand U19447 (N_19447,N_15893,N_15843);
nor U19448 (N_19448,N_15965,N_15850);
nor U19449 (N_19449,N_18332,N_16869);
nand U19450 (N_19450,N_17432,N_15713);
nand U19451 (N_19451,N_16908,N_18170);
nand U19452 (N_19452,N_18510,N_16484);
or U19453 (N_19453,N_17157,N_18268);
nand U19454 (N_19454,N_18150,N_17504);
or U19455 (N_19455,N_16741,N_17607);
nand U19456 (N_19456,N_17186,N_17121);
nand U19457 (N_19457,N_17685,N_18360);
nand U19458 (N_19458,N_18505,N_18193);
nand U19459 (N_19459,N_17359,N_18466);
nand U19460 (N_19460,N_18592,N_16893);
xnor U19461 (N_19461,N_16381,N_17722);
nor U19462 (N_19462,N_17051,N_15846);
nor U19463 (N_19463,N_18286,N_17539);
and U19464 (N_19464,N_16892,N_17322);
and U19465 (N_19465,N_15962,N_18429);
or U19466 (N_19466,N_17876,N_16435);
nand U19467 (N_19467,N_16361,N_16628);
nor U19468 (N_19468,N_17314,N_16078);
nor U19469 (N_19469,N_18587,N_16223);
xor U19470 (N_19470,N_17870,N_18394);
nand U19471 (N_19471,N_16694,N_16955);
nand U19472 (N_19472,N_16254,N_18610);
nand U19473 (N_19473,N_17262,N_18570);
xor U19474 (N_19474,N_15740,N_17807);
xnor U19475 (N_19475,N_17804,N_16423);
and U19476 (N_19476,N_18617,N_15675);
xnor U19477 (N_19477,N_17054,N_17842);
xnor U19478 (N_19478,N_15730,N_16855);
or U19479 (N_19479,N_18300,N_17421);
or U19480 (N_19480,N_17329,N_16815);
nor U19481 (N_19481,N_17995,N_17568);
nand U19482 (N_19482,N_17029,N_16039);
nor U19483 (N_19483,N_17950,N_16733);
nor U19484 (N_19484,N_18704,N_17353);
xnor U19485 (N_19485,N_18726,N_18351);
xnor U19486 (N_19486,N_15821,N_16514);
and U19487 (N_19487,N_16722,N_17493);
or U19488 (N_19488,N_17200,N_18386);
nand U19489 (N_19489,N_15744,N_17776);
nand U19490 (N_19490,N_16346,N_18374);
or U19491 (N_19491,N_16322,N_17264);
nor U19492 (N_19492,N_15925,N_17191);
xor U19493 (N_19493,N_17506,N_16706);
nor U19494 (N_19494,N_16836,N_17879);
xnor U19495 (N_19495,N_17495,N_16619);
xor U19496 (N_19496,N_15737,N_16160);
or U19497 (N_19497,N_16285,N_17111);
and U19498 (N_19498,N_18461,N_17444);
nor U19499 (N_19499,N_16525,N_18110);
nor U19500 (N_19500,N_17058,N_17937);
nor U19501 (N_19501,N_16719,N_16960);
or U19502 (N_19502,N_16241,N_15934);
or U19503 (N_19503,N_17258,N_18716);
and U19504 (N_19504,N_18440,N_16609);
or U19505 (N_19505,N_16725,N_16651);
xor U19506 (N_19506,N_16132,N_17862);
nand U19507 (N_19507,N_17109,N_17963);
and U19508 (N_19508,N_17947,N_17190);
or U19509 (N_19509,N_18401,N_16335);
nand U19510 (N_19510,N_15975,N_17990);
or U19511 (N_19511,N_16043,N_18020);
xor U19512 (N_19512,N_15765,N_16107);
nor U19513 (N_19513,N_16353,N_17782);
nor U19514 (N_19514,N_16507,N_18207);
and U19515 (N_19515,N_16991,N_18573);
and U19516 (N_19516,N_18049,N_18201);
nor U19517 (N_19517,N_17245,N_17102);
or U19518 (N_19518,N_16411,N_16567);
or U19519 (N_19519,N_18574,N_15633);
or U19520 (N_19520,N_17016,N_16060);
xnor U19521 (N_19521,N_18313,N_17424);
nor U19522 (N_19522,N_17766,N_16584);
nor U19523 (N_19523,N_17982,N_17458);
nand U19524 (N_19524,N_18277,N_18596);
nand U19525 (N_19525,N_18164,N_17866);
and U19526 (N_19526,N_15717,N_16805);
nand U19527 (N_19527,N_17091,N_16618);
nand U19528 (N_19528,N_16452,N_17336);
or U19529 (N_19529,N_18485,N_17386);
nand U19530 (N_19530,N_17101,N_16215);
or U19531 (N_19531,N_18670,N_17107);
or U19532 (N_19532,N_18169,N_17620);
or U19533 (N_19533,N_16602,N_15760);
nand U19534 (N_19534,N_18501,N_16511);
or U19535 (N_19535,N_17690,N_15637);
nand U19536 (N_19536,N_17173,N_18269);
xnor U19537 (N_19537,N_18507,N_17485);
or U19538 (N_19538,N_16526,N_17483);
or U19539 (N_19539,N_15772,N_18344);
and U19540 (N_19540,N_17372,N_18212);
or U19541 (N_19541,N_17429,N_17277);
xnor U19542 (N_19542,N_17844,N_15882);
or U19543 (N_19543,N_15828,N_16186);
and U19544 (N_19544,N_17366,N_16431);
xnor U19545 (N_19545,N_16474,N_17582);
nand U19546 (N_19546,N_16087,N_16941);
and U19547 (N_19547,N_17931,N_16142);
and U19548 (N_19548,N_16037,N_18633);
nor U19549 (N_19549,N_16670,N_18714);
xnor U19550 (N_19550,N_17197,N_16061);
nor U19551 (N_19551,N_16121,N_18216);
and U19552 (N_19552,N_17475,N_16845);
nand U19553 (N_19553,N_16492,N_17867);
xor U19554 (N_19554,N_16797,N_16510);
xnor U19555 (N_19555,N_17334,N_17280);
nand U19556 (N_19556,N_18106,N_17667);
nand U19557 (N_19557,N_17434,N_17057);
nor U19558 (N_19558,N_16782,N_17966);
xnor U19559 (N_19559,N_18341,N_18228);
nor U19560 (N_19560,N_18307,N_17726);
and U19561 (N_19561,N_16326,N_18438);
nor U19562 (N_19562,N_18259,N_16100);
or U19563 (N_19563,N_16196,N_15796);
and U19564 (N_19564,N_17079,N_16173);
and U19565 (N_19565,N_17781,N_16582);
xnor U19566 (N_19566,N_17368,N_18057);
nor U19567 (N_19567,N_17135,N_18686);
or U19568 (N_19568,N_17379,N_16671);
nand U19569 (N_19569,N_18155,N_17202);
nand U19570 (N_19570,N_17895,N_16311);
xor U19571 (N_19571,N_18452,N_17305);
or U19572 (N_19572,N_17498,N_18535);
or U19573 (N_19573,N_15901,N_15838);
or U19574 (N_19574,N_17392,N_17139);
and U19575 (N_19575,N_18641,N_16244);
and U19576 (N_19576,N_17137,N_17789);
xnor U19577 (N_19577,N_16357,N_18067);
nor U19578 (N_19578,N_17119,N_16823);
or U19579 (N_19579,N_18553,N_17837);
and U19580 (N_19580,N_16315,N_16211);
nor U19581 (N_19581,N_18565,N_17188);
nand U19582 (N_19582,N_16739,N_17809);
nand U19583 (N_19583,N_18159,N_15806);
or U19584 (N_19584,N_18451,N_15800);
or U19585 (N_19585,N_16010,N_16178);
nand U19586 (N_19586,N_16777,N_18480);
nand U19587 (N_19587,N_17916,N_16466);
or U19588 (N_19588,N_18202,N_16356);
xor U19589 (N_19589,N_17407,N_17729);
and U19590 (N_19590,N_18178,N_18515);
nand U19591 (N_19591,N_18072,N_17241);
nand U19592 (N_19592,N_18043,N_18161);
xor U19593 (N_19593,N_15906,N_17383);
and U19594 (N_19594,N_17643,N_18709);
nor U19595 (N_19595,N_17805,N_18584);
or U19596 (N_19596,N_15739,N_15816);
nor U19597 (N_19597,N_18653,N_18205);
or U19598 (N_19598,N_17934,N_17695);
nor U19599 (N_19599,N_16409,N_17147);
nor U19600 (N_19600,N_15699,N_17933);
nand U19601 (N_19601,N_18655,N_17645);
nor U19602 (N_19602,N_18744,N_17696);
and U19603 (N_19603,N_18467,N_15887);
and U19604 (N_19604,N_16427,N_18168);
and U19605 (N_19605,N_16793,N_16481);
and U19606 (N_19606,N_17007,N_15632);
and U19607 (N_19607,N_16740,N_17956);
nor U19608 (N_19608,N_18336,N_16825);
and U19609 (N_19609,N_17413,N_16396);
nor U19610 (N_19610,N_16089,N_17578);
or U19611 (N_19611,N_16430,N_16800);
and U19612 (N_19612,N_15799,N_18196);
nand U19613 (N_19613,N_17793,N_16875);
nor U19614 (N_19614,N_18265,N_16389);
and U19615 (N_19615,N_17338,N_18745);
xor U19616 (N_19616,N_16123,N_16611);
nor U19617 (N_19617,N_16742,N_17655);
or U19618 (N_19618,N_16465,N_18371);
nand U19619 (N_19619,N_16485,N_15743);
and U19620 (N_19620,N_15646,N_17547);
xnor U19621 (N_19621,N_18640,N_17686);
nor U19622 (N_19622,N_18567,N_17330);
xnor U19623 (N_19623,N_18249,N_17526);
nor U19624 (N_19624,N_18594,N_18472);
nand U19625 (N_19625,N_16323,N_17678);
and U19626 (N_19626,N_16302,N_15781);
nor U19627 (N_19627,N_16530,N_18647);
nand U19628 (N_19628,N_18627,N_15879);
xnor U19629 (N_19629,N_17041,N_16634);
nor U19630 (N_19630,N_16393,N_18264);
and U19631 (N_19631,N_17742,N_15710);
or U19632 (N_19632,N_16558,N_16111);
xor U19633 (N_19633,N_17272,N_15840);
nor U19634 (N_19634,N_15837,N_15853);
and U19635 (N_19635,N_16056,N_16129);
and U19636 (N_19636,N_15691,N_17196);
or U19637 (N_19637,N_17072,N_18648);
nand U19638 (N_19638,N_16324,N_17068);
and U19639 (N_19639,N_17252,N_17110);
nor U19640 (N_19640,N_15953,N_18137);
and U19641 (N_19641,N_17848,N_18046);
nand U19642 (N_19642,N_17864,N_15688);
xnor U19643 (N_19643,N_18428,N_16283);
or U19644 (N_19644,N_16161,N_16337);
and U19645 (N_19645,N_17767,N_18130);
nand U19646 (N_19646,N_16437,N_17701);
and U19647 (N_19647,N_16930,N_16180);
xnor U19648 (N_19648,N_17561,N_17450);
and U19649 (N_19649,N_18069,N_17894);
nor U19650 (N_19650,N_18496,N_17661);
nor U19651 (N_19651,N_18195,N_17236);
nand U19652 (N_19652,N_15956,N_17581);
nand U19653 (N_19653,N_16903,N_16520);
nand U19654 (N_19654,N_18521,N_16701);
nor U19655 (N_19655,N_16939,N_16577);
nand U19656 (N_19656,N_18132,N_18551);
nor U19657 (N_19657,N_16077,N_17570);
or U19658 (N_19658,N_15784,N_18586);
or U19659 (N_19659,N_18320,N_17812);
nand U19660 (N_19660,N_15888,N_16004);
nor U19661 (N_19661,N_15899,N_17698);
or U19662 (N_19662,N_16002,N_15749);
nand U19663 (N_19663,N_15885,N_17510);
and U19664 (N_19664,N_16693,N_17374);
or U19665 (N_19665,N_15832,N_16331);
and U19666 (N_19666,N_17525,N_18100);
nor U19667 (N_19667,N_16665,N_16428);
and U19668 (N_19668,N_17635,N_17488);
nor U19669 (N_19669,N_15682,N_18238);
and U19670 (N_19670,N_18511,N_18117);
or U19671 (N_19671,N_16203,N_17099);
nor U19672 (N_19672,N_16486,N_17469);
xnor U19673 (N_19673,N_16055,N_18419);
or U19674 (N_19674,N_18693,N_16080);
or U19675 (N_19675,N_16192,N_17654);
nor U19676 (N_19676,N_17777,N_17961);
and U19677 (N_19677,N_16810,N_17801);
nand U19678 (N_19678,N_16886,N_17567);
and U19679 (N_19679,N_18475,N_18198);
and U19680 (N_19680,N_16550,N_16281);
nand U19681 (N_19681,N_17615,N_18413);
nand U19682 (N_19682,N_15845,N_17605);
and U19683 (N_19683,N_17459,N_16849);
xnor U19684 (N_19684,N_16837,N_16677);
nand U19685 (N_19685,N_18631,N_15849);
and U19686 (N_19686,N_18652,N_16287);
nand U19687 (N_19687,N_17378,N_16380);
and U19688 (N_19688,N_18514,N_16978);
or U19689 (N_19689,N_18293,N_15766);
xor U19690 (N_19690,N_18179,N_18549);
or U19691 (N_19691,N_17505,N_17902);
and U19692 (N_19692,N_17609,N_18180);
nor U19693 (N_19693,N_16158,N_17310);
and U19694 (N_19694,N_16820,N_16318);
and U19695 (N_19695,N_15931,N_16235);
xor U19696 (N_19696,N_15855,N_16643);
nor U19697 (N_19697,N_17024,N_16022);
nor U19698 (N_19698,N_16932,N_16818);
nor U19699 (N_19699,N_18084,N_16969);
and U19700 (N_19700,N_18568,N_18455);
and U19701 (N_19701,N_16900,N_17749);
nand U19702 (N_19702,N_17229,N_18398);
nand U19703 (N_19703,N_17549,N_18517);
nand U19704 (N_19704,N_18423,N_17649);
nand U19705 (N_19705,N_15874,N_18556);
nand U19706 (N_19706,N_17794,N_18291);
or U19707 (N_19707,N_16689,N_17250);
or U19708 (N_19708,N_16711,N_18076);
nor U19709 (N_19709,N_16202,N_16883);
xnor U19710 (N_19710,N_16637,N_18708);
nor U19711 (N_19711,N_18600,N_17240);
and U19712 (N_19712,N_18364,N_16509);
nor U19713 (N_19713,N_15813,N_18528);
nand U19714 (N_19714,N_17989,N_17580);
nand U19715 (N_19715,N_16501,N_18558);
and U19716 (N_19716,N_18473,N_16743);
and U19717 (N_19717,N_16090,N_17341);
xor U19718 (N_19718,N_16730,N_15676);
or U19719 (N_19719,N_18285,N_18375);
nand U19720 (N_19720,N_17770,N_17499);
and U19721 (N_19721,N_18247,N_17244);
nand U19722 (N_19722,N_18697,N_16403);
nor U19723 (N_19723,N_17536,N_17986);
and U19724 (N_19724,N_18006,N_15625);
or U19725 (N_19725,N_16549,N_17221);
nor U19726 (N_19726,N_15947,N_16047);
and U19727 (N_19727,N_16647,N_16109);
and U19728 (N_19728,N_17786,N_15714);
and U19729 (N_19729,N_16237,N_15746);
or U19730 (N_19730,N_17347,N_16735);
and U19731 (N_19731,N_18165,N_17813);
or U19732 (N_19732,N_16663,N_15917);
and U19733 (N_19733,N_16778,N_18023);
nor U19734 (N_19734,N_17811,N_17819);
or U19735 (N_19735,N_16625,N_16185);
and U19736 (N_19736,N_18191,N_15629);
or U19737 (N_19737,N_16330,N_17987);
or U19738 (N_19738,N_17939,N_17448);
and U19739 (N_19739,N_16284,N_15964);
nor U19740 (N_19740,N_16705,N_15674);
xor U19741 (N_19741,N_18000,N_15747);
nand U19742 (N_19742,N_15880,N_16487);
nor U19743 (N_19743,N_18402,N_16300);
or U19744 (N_19744,N_18144,N_18208);
nand U19745 (N_19745,N_16901,N_18748);
or U19746 (N_19746,N_15753,N_16157);
and U19747 (N_19747,N_16781,N_17299);
nand U19748 (N_19748,N_16809,N_17614);
nor U19749 (N_19749,N_16654,N_17952);
nand U19750 (N_19750,N_17040,N_15940);
nand U19751 (N_19751,N_17824,N_18330);
xnor U19752 (N_19752,N_18616,N_17826);
nor U19753 (N_19753,N_17472,N_17857);
nand U19754 (N_19754,N_16515,N_16566);
and U19755 (N_19755,N_17948,N_17587);
xor U19756 (N_19756,N_17785,N_18434);
and U19757 (N_19757,N_16272,N_17543);
xnor U19758 (N_19758,N_17124,N_17257);
and U19759 (N_19759,N_17657,N_16524);
and U19760 (N_19760,N_15875,N_18499);
or U19761 (N_19761,N_17237,N_15626);
nand U19762 (N_19762,N_18146,N_18630);
or U19763 (N_19763,N_15686,N_16833);
nand U19764 (N_19764,N_18414,N_17922);
nor U19765 (N_19765,N_17883,N_16716);
and U19766 (N_19766,N_18432,N_18612);
nor U19767 (N_19767,N_16421,N_15718);
nand U19768 (N_19768,N_16789,N_18437);
nor U19769 (N_19769,N_15680,N_18564);
or U19770 (N_19770,N_17078,N_18030);
nor U19771 (N_19771,N_18690,N_17088);
nor U19772 (N_19772,N_18415,N_17516);
or U19773 (N_19773,N_15685,N_18015);
or U19774 (N_19774,N_17998,N_16482);
or U19775 (N_19775,N_16600,N_16992);
or U19776 (N_19776,N_18577,N_18322);
and U19777 (N_19777,N_15878,N_16128);
nand U19778 (N_19778,N_17563,N_18611);
and U19779 (N_19779,N_15759,N_16814);
or U19780 (N_19780,N_17838,N_16885);
nand U19781 (N_19781,N_15835,N_18187);
and U19782 (N_19782,N_17968,N_18167);
and U19783 (N_19783,N_17496,N_16453);
nand U19784 (N_19784,N_17571,N_18397);
nor U19785 (N_19785,N_18581,N_16645);
nor U19786 (N_19786,N_16226,N_18214);
xnor U19787 (N_19787,N_16664,N_15987);
nor U19788 (N_19788,N_17174,N_16088);
nor U19789 (N_19789,N_15908,N_16956);
and U19790 (N_19790,N_16779,N_16907);
xor U19791 (N_19791,N_16288,N_16858);
nor U19792 (N_19792,N_17352,N_16571);
nor U19793 (N_19793,N_18007,N_18010);
and U19794 (N_19794,N_15881,N_18735);
and U19795 (N_19795,N_18044,N_17278);
nand U19796 (N_19796,N_18311,N_16752);
xor U19797 (N_19797,N_18734,N_16923);
nand U19798 (N_19798,N_18082,N_18223);
and U19799 (N_19799,N_17106,N_18033);
and U19800 (N_19800,N_17490,N_15808);
or U19801 (N_19801,N_16998,N_16848);
nor U19802 (N_19802,N_17841,N_17978);
and U19803 (N_19803,N_17204,N_18591);
nor U19804 (N_19804,N_16682,N_17246);
nand U19805 (N_19805,N_16678,N_18128);
and U19806 (N_19806,N_16794,N_17441);
and U19807 (N_19807,N_16650,N_16817);
xnor U19808 (N_19808,N_18696,N_15748);
or U19809 (N_19809,N_16450,N_18038);
xor U19810 (N_19810,N_15876,N_17641);
or U19811 (N_19811,N_16291,N_16044);
and U19812 (N_19812,N_16761,N_16425);
nor U19813 (N_19813,N_15937,N_18333);
nor U19814 (N_19814,N_17907,N_17028);
or U19815 (N_19815,N_17569,N_16181);
nor U19816 (N_19816,N_17851,N_18576);
or U19817 (N_19817,N_18639,N_15788);
nand U19818 (N_19818,N_16744,N_18684);
or U19819 (N_19819,N_18463,N_16388);
xor U19820 (N_19820,N_18424,N_17622);
and U19821 (N_19821,N_15770,N_18156);
and U19822 (N_19822,N_17705,N_17212);
or U19823 (N_19823,N_15805,N_17187);
nand U19824 (N_19824,N_18056,N_18338);
nor U19825 (N_19825,N_18378,N_18138);
nor U19826 (N_19826,N_18352,N_18373);
nor U19827 (N_19827,N_16636,N_18111);
or U19828 (N_19828,N_17900,N_17015);
or U19829 (N_19829,N_17697,N_16266);
or U19830 (N_19830,N_17466,N_15948);
nor U19831 (N_19831,N_17759,N_18458);
and U19832 (N_19832,N_16700,N_18315);
or U19833 (N_19833,N_17999,N_15696);
xnor U19834 (N_19834,N_17356,N_18387);
and U19835 (N_19835,N_17955,N_17396);
or U19836 (N_19836,N_16174,N_16270);
or U19837 (N_19837,N_17076,N_18469);
or U19838 (N_19838,N_16987,N_16497);
or U19839 (N_19839,N_18427,N_18546);
xor U19840 (N_19840,N_15647,N_17279);
xor U19841 (N_19841,N_16376,N_17116);
or U19842 (N_19842,N_18540,N_17426);
nand U19843 (N_19843,N_16122,N_15988);
nand U19844 (N_19844,N_18443,N_17266);
nand U19845 (N_19845,N_17618,N_18209);
or U19846 (N_19846,N_15706,N_18040);
or U19847 (N_19847,N_18484,N_18544);
nor U19848 (N_19848,N_15754,N_18283);
nor U19849 (N_19849,N_18689,N_17636);
xor U19850 (N_19850,N_18691,N_15776);
and U19851 (N_19851,N_16419,N_18603);
and U19852 (N_19852,N_16867,N_16228);
nor U19853 (N_19853,N_17861,N_16189);
or U19854 (N_19854,N_17716,N_17369);
or U19855 (N_19855,N_15652,N_16227);
or U19856 (N_19856,N_17853,N_17736);
nand U19857 (N_19857,N_16565,N_15924);
nand U19858 (N_19858,N_18624,N_16145);
nor U19859 (N_19859,N_17623,N_18527);
and U19860 (N_19860,N_18062,N_16259);
nand U19861 (N_19861,N_16679,N_17535);
nand U19862 (N_19862,N_16616,N_17192);
nand U19863 (N_19863,N_17461,N_18628);
nand U19864 (N_19864,N_17531,N_17815);
and U19865 (N_19865,N_16940,N_18644);
and U19866 (N_19866,N_16726,N_17035);
nand U19867 (N_19867,N_18078,N_16822);
or U19868 (N_19868,N_17326,N_17672);
or U19869 (N_19869,N_17953,N_16768);
nand U19870 (N_19870,N_16947,N_17226);
or U19871 (N_19871,N_17797,N_18465);
nand U19872 (N_19872,N_17639,N_17481);
and U19873 (N_19873,N_17013,N_18537);
or U19874 (N_19874,N_18116,N_15836);
nor U19875 (N_19875,N_17523,N_17399);
or U19876 (N_19876,N_15787,N_16170);
and U19877 (N_19877,N_16811,N_18273);
and U19878 (N_19878,N_16557,N_16455);
xnor U19879 (N_19879,N_18051,N_15911);
nand U19880 (N_19880,N_18599,N_17014);
nor U19881 (N_19881,N_16153,N_15868);
or U19882 (N_19882,N_17268,N_16784);
and U19883 (N_19883,N_17081,N_17919);
nand U19884 (N_19884,N_15932,N_17117);
xnor U19885 (N_19885,N_16560,N_17482);
and U19886 (N_19886,N_16934,N_17680);
nor U19887 (N_19887,N_16860,N_18112);
nand U19888 (N_19888,N_17163,N_16253);
nor U19889 (N_19889,N_15663,N_18645);
nor U19890 (N_19890,N_18017,N_18356);
and U19891 (N_19891,N_15723,N_18669);
and U19892 (N_19892,N_16661,N_17810);
nor U19893 (N_19893,N_17410,N_16404);
nor U19894 (N_19894,N_17275,N_15733);
and U19895 (N_19895,N_15915,N_16334);
xnor U19896 (N_19896,N_16095,N_17694);
and U19897 (N_19897,N_16195,N_15660);
nor U19898 (N_19898,N_15659,N_16798);
and U19899 (N_19899,N_15865,N_17597);
and U19900 (N_19900,N_15775,N_18727);
and U19901 (N_19901,N_18321,N_16303);
and U19902 (N_19902,N_16620,N_18618);
nand U19903 (N_19903,N_18453,N_17425);
or U19904 (N_19904,N_17772,N_17140);
or U19905 (N_19905,N_17123,N_18666);
xnor U19906 (N_19906,N_18561,N_18502);
and U19907 (N_19907,N_15635,N_17903);
or U19908 (N_19908,N_16684,N_17451);
or U19909 (N_19909,N_16766,N_16920);
xnor U19910 (N_19910,N_16000,N_16623);
nand U19911 (N_19911,N_16580,N_18688);
or U19912 (N_19912,N_17331,N_18548);
nor U19913 (N_19913,N_15982,N_18032);
and U19914 (N_19914,N_18474,N_18706);
or U19915 (N_19915,N_17069,N_17835);
or U19916 (N_19916,N_18595,N_16791);
and U19917 (N_19917,N_16313,N_17992);
nor U19918 (N_19918,N_17796,N_16366);
xor U19919 (N_19919,N_15661,N_17557);
and U19920 (N_19920,N_16904,N_18135);
and U19921 (N_19921,N_17303,N_18552);
nor U19922 (N_19922,N_16072,N_18274);
xnor U19923 (N_19923,N_18133,N_17144);
nand U19924 (N_19924,N_18381,N_18213);
or U19925 (N_19925,N_16067,N_16534);
and U19926 (N_19926,N_15921,N_18143);
nand U19927 (N_19927,N_16332,N_17004);
nor U19928 (N_19928,N_17289,N_17558);
or U19929 (N_19929,N_17154,N_18326);
or U19930 (N_19930,N_18700,N_17285);
or U19931 (N_19931,N_17445,N_17725);
nand U19932 (N_19932,N_17189,N_16984);
xnor U19933 (N_19933,N_15980,N_17010);
or U19934 (N_19934,N_18358,N_16555);
nand U19935 (N_19935,N_18410,N_17872);
and U19936 (N_19936,N_18014,N_18009);
nand U19937 (N_19937,N_16965,N_17599);
and U19938 (N_19938,N_15662,N_17530);
and U19939 (N_19939,N_17896,N_17651);
and U19940 (N_19940,N_16379,N_17943);
nand U19941 (N_19941,N_17131,N_17478);
nor U19942 (N_19942,N_16325,N_16842);
and U19943 (N_19943,N_17988,N_18176);
nand U19944 (N_19944,N_16045,N_16687);
and U19945 (N_19945,N_18422,N_17632);
or U19946 (N_19946,N_16862,N_18687);
nand U19947 (N_19947,N_18730,N_18694);
nand U19948 (N_19948,N_15703,N_15811);
or U19949 (N_19949,N_17600,N_18512);
nand U19950 (N_19950,N_18447,N_16771);
nand U19951 (N_19951,N_16101,N_15830);
nand U19952 (N_19952,N_17548,N_18345);
or U19953 (N_19953,N_18361,N_17630);
or U19954 (N_19954,N_17169,N_18620);
or U19955 (N_19955,N_17700,N_17442);
nand U19956 (N_19956,N_17062,N_18024);
and U19957 (N_19957,N_17960,N_17354);
or U19958 (N_19958,N_16476,N_16968);
nand U19959 (N_19959,N_18244,N_17723);
and U19960 (N_19960,N_16074,N_17763);
or U19961 (N_19961,N_16579,N_16521);
nand U19962 (N_19962,N_15702,N_17185);
xor U19963 (N_19963,N_17073,N_16871);
xor U19964 (N_19964,N_18255,N_16799);
or U19965 (N_19965,N_18673,N_16538);
nor U19966 (N_19966,N_16720,N_17590);
or U19967 (N_19967,N_15890,N_16229);
nor U19968 (N_19968,N_18109,N_17538);
and U19969 (N_19969,N_16834,N_15942);
or U19970 (N_19970,N_16402,N_15793);
and U19971 (N_19971,N_16374,N_16523);
nand U19972 (N_19972,N_17208,N_16604);
xnor U19973 (N_19973,N_16517,N_16676);
nand U19974 (N_19974,N_16503,N_18141);
and U19975 (N_19975,N_17328,N_16038);
and U19976 (N_19976,N_17664,N_16593);
and U19977 (N_19977,N_18672,N_18317);
or U19978 (N_19978,N_16924,N_18391);
or U19979 (N_19979,N_16724,N_16936);
xor U19980 (N_19980,N_16861,N_17284);
xor U19981 (N_19981,N_15852,N_17047);
xor U19982 (N_19982,N_15905,N_17134);
or U19983 (N_19983,N_17467,N_16490);
or U19984 (N_19984,N_16116,N_16405);
nor U19985 (N_19985,N_16424,N_16988);
or U19986 (N_19986,N_16891,N_18613);
nor U19987 (N_19987,N_16468,N_16962);
or U19988 (N_19988,N_17650,N_16686);
or U19989 (N_19989,N_16065,N_16320);
nand U19990 (N_19990,N_17602,N_16276);
nand U19991 (N_19991,N_16447,N_18129);
xnor U19992 (N_19992,N_16401,N_15667);
nand U19993 (N_19993,N_17194,N_17452);
and U19994 (N_19994,N_18001,N_17647);
nand U19995 (N_19995,N_15812,N_16819);
nand U19996 (N_19996,N_16295,N_17840);
nor U19997 (N_19997,N_17633,N_17904);
nand U19998 (N_19998,N_16124,N_17370);
xnor U19999 (N_19999,N_15792,N_17944);
or U20000 (N_20000,N_17443,N_16310);
xor U20001 (N_20001,N_16176,N_16516);
nand U20002 (N_20002,N_18047,N_18743);
nor U20003 (N_20003,N_18316,N_16473);
and U20004 (N_20004,N_15650,N_17209);
nor U20005 (N_20005,N_17402,N_17477);
and U20006 (N_20006,N_17849,N_18731);
and U20007 (N_20007,N_15909,N_17327);
or U20008 (N_20008,N_16182,N_18158);
nand U20009 (N_20009,N_16764,N_16091);
nor U20010 (N_20010,N_15930,N_16808);
and U20011 (N_20011,N_17100,N_16680);
nand U20012 (N_20012,N_15842,N_16207);
nand U20013 (N_20013,N_17942,N_17291);
and U20014 (N_20014,N_17064,N_15945);
nand U20015 (N_20015,N_16373,N_18746);
xnor U20016 (N_20016,N_18723,N_18231);
xor U20017 (N_20017,N_17201,N_18449);
and U20018 (N_20018,N_18626,N_16927);
or U20019 (N_20019,N_15795,N_16840);
and U20020 (N_20020,N_18232,N_17762);
and U20021 (N_20021,N_16333,N_18272);
or U20022 (N_20022,N_16581,N_16697);
nor U20023 (N_20023,N_16265,N_16672);
or U20024 (N_20024,N_18676,N_17471);
nor U20025 (N_20025,N_17302,N_16240);
nor U20026 (N_20026,N_17827,N_17096);
and U20027 (N_20027,N_17802,N_17704);
nor U20028 (N_20028,N_18275,N_18365);
nor U20029 (N_20029,N_16477,N_16085);
nand U20030 (N_20030,N_15681,N_17601);
nor U20031 (N_20031,N_17080,N_15929);
nand U20032 (N_20032,N_18059,N_16097);
nor U20033 (N_20033,N_15771,N_16631);
xor U20034 (N_20034,N_15986,N_18126);
and U20035 (N_20035,N_16392,N_18122);
and U20036 (N_20036,N_18420,N_16321);
nand U20037 (N_20037,N_15745,N_16076);
nor U20038 (N_20038,N_16168,N_17143);
xor U20039 (N_20039,N_17653,N_18194);
nor U20040 (N_20040,N_18550,N_18288);
or U20041 (N_20041,N_18651,N_18396);
nand U20042 (N_20042,N_15752,N_15973);
and U20043 (N_20043,N_16976,N_18241);
and U20044 (N_20044,N_18153,N_16308);
nor U20045 (N_20045,N_17585,N_15735);
nor U20046 (N_20046,N_18346,N_17935);
and U20047 (N_20047,N_17337,N_18635);
nand U20048 (N_20048,N_17393,N_15829);
and U20049 (N_20049,N_15978,N_17625);
nor U20050 (N_20050,N_15720,N_15898);
nor U20051 (N_20051,N_17724,N_16879);
and U20052 (N_20052,N_17380,N_17803);
nand U20053 (N_20053,N_17019,N_15778);
nor U20054 (N_20054,N_16933,N_18041);
nor U20055 (N_20055,N_16377,N_17501);
and U20056 (N_20056,N_16433,N_16638);
nor U20057 (N_20057,N_17932,N_17666);
and U20058 (N_20058,N_16137,N_17094);
and U20059 (N_20059,N_18027,N_18446);
or U20060 (N_20060,N_16713,N_17675);
and U20061 (N_20061,N_15995,N_17739);
or U20062 (N_20062,N_18654,N_17408);
xnor U20063 (N_20063,N_17687,N_17517);
or U20064 (N_20064,N_15804,N_16420);
nor U20065 (N_20065,N_16533,N_16198);
nor U20066 (N_20066,N_17593,N_16054);
nand U20067 (N_20067,N_18230,N_18385);
nor U20068 (N_20068,N_17178,N_16696);
or U20069 (N_20069,N_16961,N_17554);
nor U20070 (N_20070,N_16017,N_18061);
nor U20071 (N_20071,N_15831,N_16753);
nand U20072 (N_20072,N_18569,N_16155);
and U20073 (N_20073,N_15701,N_18407);
xnor U20074 (N_20074,N_16370,N_17149);
nand U20075 (N_20075,N_16656,N_18037);
and U20076 (N_20076,N_15666,N_16200);
nand U20077 (N_20077,N_18404,N_16362);
and U20078 (N_20078,N_15712,N_15823);
nor U20079 (N_20079,N_17405,N_17885);
nand U20080 (N_20080,N_16838,N_16220);
nor U20081 (N_20081,N_17397,N_16232);
nand U20082 (N_20082,N_16171,N_17420);
or U20083 (N_20083,N_16746,N_15970);
or U20084 (N_20084,N_16597,N_16854);
nor U20085 (N_20085,N_17120,N_15774);
and U20086 (N_20086,N_17626,N_18234);
nand U20087 (N_20087,N_16269,N_17918);
nor U20088 (N_20088,N_17247,N_17006);
nand U20089 (N_20089,N_18204,N_17409);
nor U20090 (N_20090,N_16944,N_17524);
or U20091 (N_20091,N_16850,N_15716);
nand U20092 (N_20092,N_16954,N_16718);
nand U20093 (N_20093,N_15783,N_17575);
and U20094 (N_20094,N_15979,N_16305);
nand U20095 (N_20095,N_16918,N_16673);
xnor U20096 (N_20096,N_16462,N_16025);
nand U20097 (N_20097,N_18741,N_17611);
or U20098 (N_20098,N_17259,N_17416);
xnor U20099 (N_20099,N_15814,N_16319);
nor U20100 (N_20100,N_16562,N_17577);
xnor U20101 (N_20101,N_16919,N_17741);
and U20102 (N_20102,N_18045,N_16282);
nand U20103 (N_20103,N_17233,N_17699);
nor U20104 (N_20104,N_15697,N_17613);
or U20105 (N_20105,N_15773,N_16914);
nand U20106 (N_20106,N_16127,N_16506);
or U20107 (N_20107,N_18354,N_16882);
nor U20108 (N_20108,N_16277,N_17300);
nand U20109 (N_20109,N_18547,N_18590);
or U20110 (N_20110,N_16458,N_18287);
or U20111 (N_20111,N_17098,N_17753);
nor U20112 (N_20112,N_16133,N_16216);
and U20113 (N_20113,N_16138,N_17234);
nor U20114 (N_20114,N_17075,N_18175);
nor U20115 (N_20115,N_16925,N_15902);
nor U20116 (N_20116,N_16205,N_17714);
nand U20117 (N_20117,N_16400,N_18050);
nor U20118 (N_20118,N_16204,N_18384);
or U20119 (N_20119,N_16028,N_16983);
and U20120 (N_20120,N_16079,N_16210);
nor U20121 (N_20121,N_16780,N_16098);
nand U20122 (N_20122,N_15993,N_18498);
nor U20123 (N_20123,N_17886,N_18665);
and U20124 (N_20124,N_16384,N_16023);
nor U20125 (N_20125,N_18506,N_17717);
nand U20126 (N_20126,N_18664,N_17048);
xnor U20127 (N_20127,N_17534,N_15798);
nor U20128 (N_20128,N_16640,N_17412);
nor U20129 (N_20129,N_16201,N_18638);
nand U20130 (N_20130,N_15858,N_16233);
or U20131 (N_20131,N_16657,N_16899);
and U20132 (N_20132,N_17874,N_17608);
xor U20133 (N_20133,N_17446,N_17390);
nand U20134 (N_20134,N_16187,N_17972);
or U20135 (N_20135,N_18495,N_17437);
nor U20136 (N_20136,N_17479,N_16864);
or U20137 (N_20137,N_16717,N_15726);
xnor U20138 (N_20138,N_17182,N_17161);
and U20139 (N_20139,N_16698,N_18632);
or U20140 (N_20140,N_17045,N_18189);
nand U20141 (N_20141,N_18487,N_18519);
and U20142 (N_20142,N_18108,N_16221);
or U20143 (N_20143,N_16001,N_18297);
and U20144 (N_20144,N_18623,N_15648);
nand U20145 (N_20145,N_17005,N_17065);
nand U20146 (N_20146,N_17640,N_17067);
and U20147 (N_20147,N_18382,N_18488);
and U20148 (N_20148,N_17970,N_17476);
and U20149 (N_20149,N_15731,N_15884);
or U20150 (N_20150,N_16608,N_17489);
and U20151 (N_20151,N_18597,N_16979);
or U20152 (N_20152,N_18369,N_15896);
xor U20153 (N_20153,N_15672,N_17603);
or U20154 (N_20154,N_15847,N_18667);
and U20155 (N_20155,N_16642,N_16985);
nor U20156 (N_20156,N_17296,N_17060);
or U20157 (N_20157,N_18674,N_16895);
nor U20158 (N_20158,N_16770,N_16585);
nand U20159 (N_20159,N_18217,N_16537);
nand U20160 (N_20160,N_16258,N_18518);
xor U20161 (N_20161,N_15636,N_16175);
and U20162 (N_20162,N_15628,N_18026);
nand U20163 (N_20163,N_16935,N_17138);
nor U20164 (N_20164,N_17560,N_17917);
nand U20165 (N_20165,N_17043,N_16042);
or U20166 (N_20166,N_16119,N_16260);
nand U20167 (N_20167,N_15994,N_17132);
or U20168 (N_20168,N_17333,N_17727);
or U20169 (N_20169,N_18362,N_16449);
and U20170 (N_20170,N_16040,N_16548);
nor U20171 (N_20171,N_15670,N_16162);
xnor U20172 (N_20172,N_18060,N_16294);
xor U20173 (N_20173,N_16535,N_16478);
nor U20174 (N_20174,N_16938,N_17156);
and U20175 (N_20175,N_18239,N_18120);
or U20176 (N_20176,N_16106,N_17403);
nand U20177 (N_20177,N_16479,N_17760);
nor U20178 (N_20178,N_16832,N_15802);
and U20179 (N_20179,N_18003,N_18663);
nand U20180 (N_20180,N_16290,N_17528);
or U20181 (N_20181,N_17834,N_17211);
nand U20182 (N_20182,N_18121,N_17951);
xor U20183 (N_20183,N_17315,N_18329);
nand U20184 (N_20184,N_16344,N_17218);
nor U20185 (N_20185,N_17473,N_17911);
nand U20186 (N_20186,N_16134,N_17579);
nor U20187 (N_20187,N_18337,N_17962);
nand U20188 (N_20188,N_17342,N_17564);
nor U20189 (N_20189,N_17659,N_17591);
xnor U20190 (N_20190,N_18245,N_17381);
and U20191 (N_20191,N_18520,N_18579);
and U20192 (N_20192,N_17754,N_17126);
or U20193 (N_20193,N_17167,N_16117);
and U20194 (N_20194,N_17267,N_18380);
xor U20195 (N_20195,N_17555,N_16937);
or U20196 (N_20196,N_17511,N_17780);
nor U20197 (N_20197,N_17731,N_16213);
nor U20198 (N_20198,N_16436,N_17638);
and U20199 (N_20199,N_17176,N_18476);
and U20200 (N_20200,N_16633,N_16245);
nand U20201 (N_20201,N_15839,N_18559);
nand U20202 (N_20202,N_18554,N_17662);
or U20203 (N_20203,N_18681,N_18732);
nor U20204 (N_20204,N_16372,N_16590);
or U20205 (N_20205,N_15889,N_16086);
or U20206 (N_20206,N_16542,N_17199);
and U20207 (N_20207,N_17889,N_17500);
and U20208 (N_20208,N_18353,N_16166);
nand U20209 (N_20209,N_15951,N_18481);
nor U20210 (N_20210,N_16096,N_16964);
xor U20211 (N_20211,N_17141,N_16141);
and U20212 (N_20212,N_16443,N_16876);
or U20213 (N_20213,N_16546,N_16440);
nand U20214 (N_20214,N_16177,N_18725);
and U20215 (N_20215,N_15943,N_18197);
nand U20216 (N_20216,N_18305,N_16013);
nand U20217 (N_20217,N_16219,N_16289);
or U20218 (N_20218,N_18113,N_17816);
nor U20219 (N_20219,N_15841,N_18319);
and U20220 (N_20220,N_18699,N_16030);
and U20221 (N_20221,N_16950,N_16853);
and U20222 (N_20222,N_18065,N_18092);
nor U20223 (N_20223,N_17631,N_15961);
or U20224 (N_20224,N_18711,N_17256);
nand U20225 (N_20225,N_18532,N_17011);
and U20226 (N_20226,N_18494,N_18171);
and U20227 (N_20227,N_16256,N_17364);
and U20228 (N_20228,N_18227,N_18323);
or U20229 (N_20229,N_16385,N_16146);
nor U20230 (N_20230,N_18468,N_16464);
and U20231 (N_20231,N_18290,N_15817);
or U20232 (N_20232,N_17365,N_17360);
nor U20233 (N_20233,N_18303,N_18720);
nand U20234 (N_20234,N_16872,N_17825);
nand U20235 (N_20235,N_17890,N_17142);
xor U20236 (N_20236,N_15692,N_16495);
or U20237 (N_20237,N_16544,N_16006);
and U20238 (N_20238,N_17009,N_17273);
and U20239 (N_20239,N_17034,N_15705);
nand U20240 (N_20240,N_16257,N_16154);
xor U20241 (N_20241,N_16358,N_15895);
nor U20242 (N_20242,N_16589,N_18366);
xnor U20243 (N_20243,N_17750,N_18350);
nand U20244 (N_20244,N_16016,N_18200);
and U20245 (N_20245,N_16502,N_16851);
nor U20246 (N_20246,N_18680,N_17118);
nor U20247 (N_20247,N_16626,N_15641);
or U20248 (N_20248,N_16763,N_18304);
nor U20249 (N_20249,N_18301,N_17324);
nand U20250 (N_20250,N_17160,N_17295);
nor U20251 (N_20251,N_17852,N_18188);
nand U20252 (N_20252,N_17882,N_16583);
xnor U20253 (N_20253,N_17584,N_16669);
nand U20254 (N_20254,N_16351,N_16472);
nand U20255 (N_20255,N_16225,N_17225);
and U20256 (N_20256,N_16973,N_16255);
nand U20257 (N_20257,N_16350,N_16605);
and U20258 (N_20258,N_17363,N_16652);
xor U20259 (N_20259,N_17122,N_17242);
and U20260 (N_20260,N_17435,N_17976);
or U20261 (N_20261,N_17509,N_17003);
nor U20262 (N_20262,N_17967,N_18668);
or U20263 (N_20263,N_17321,N_16125);
or U20264 (N_20264,N_18226,N_18149);
and U20265 (N_20265,N_17453,N_15764);
and U20266 (N_20266,N_16267,N_16873);
nor U20267 (N_20267,N_17985,N_17414);
nand U20268 (N_20268,N_18740,N_15827);
nand U20269 (N_20269,N_16306,N_17823);
and U20270 (N_20270,N_15873,N_15919);
and U20271 (N_20271,N_16803,N_18368);
nand U20272 (N_20272,N_18233,N_17925);
nand U20273 (N_20273,N_16911,N_16491);
xor U20274 (N_20274,N_15653,N_16115);
and U20275 (N_20275,N_16062,N_18140);
and U20276 (N_20276,N_15824,N_17858);
nand U20277 (N_20277,N_18246,N_16897);
xnor U20278 (N_20278,N_16094,N_18091);
or U20279 (N_20279,N_17859,N_16339);
or U20280 (N_20280,N_18433,N_16494);
nand U20281 (N_20281,N_16416,N_16018);
and U20282 (N_20282,N_16338,N_16709);
or U20283 (N_20283,N_16802,N_18464);
xnor U20284 (N_20284,N_17839,N_18011);
nor U20285 (N_20285,N_16390,N_15677);
nand U20286 (N_20286,N_18282,N_17255);
nand U20287 (N_20287,N_16480,N_16394);
or U20288 (N_20288,N_16412,N_16059);
nor U20289 (N_20289,N_16504,N_17093);
nand U20290 (N_20290,N_17691,N_16912);
nor U20291 (N_20291,N_17297,N_17104);
or U20292 (N_20292,N_17550,N_17430);
or U20293 (N_20293,N_17335,N_17039);
nor U20294 (N_20294,N_17977,N_17728);
nand U20295 (N_20295,N_18379,N_18722);
nor U20296 (N_20296,N_18025,N_17746);
nand U20297 (N_20297,N_18712,N_15721);
nand U20298 (N_20298,N_18235,N_17382);
nand U20299 (N_20299,N_17115,N_16444);
and U20300 (N_20300,N_18127,N_17053);
nor U20301 (N_20301,N_16703,N_18028);
nand U20302 (N_20302,N_15903,N_15777);
xnor U20303 (N_20303,N_17598,N_16500);
and U20304 (N_20304,N_16759,N_17676);
and U20305 (N_20305,N_16063,N_18054);
or U20306 (N_20306,N_18308,N_18678);
and U20307 (N_20307,N_16035,N_17915);
nor U20308 (N_20308,N_15904,N_15734);
and U20309 (N_20309,N_16093,N_16994);
and U20310 (N_20310,N_18608,N_16114);
xnor U20311 (N_20311,N_15634,N_18070);
xnor U20312 (N_20312,N_18258,N_16684);
nor U20313 (N_20313,N_17181,N_17635);
or U20314 (N_20314,N_17428,N_15912);
xnor U20315 (N_20315,N_16761,N_16892);
nand U20316 (N_20316,N_18680,N_17874);
nor U20317 (N_20317,N_16161,N_18195);
nor U20318 (N_20318,N_17836,N_15857);
and U20319 (N_20319,N_16442,N_17307);
and U20320 (N_20320,N_17319,N_17710);
and U20321 (N_20321,N_15654,N_16325);
nor U20322 (N_20322,N_18637,N_17420);
and U20323 (N_20323,N_17157,N_17438);
nand U20324 (N_20324,N_16429,N_17113);
or U20325 (N_20325,N_17021,N_16620);
or U20326 (N_20326,N_16479,N_18622);
or U20327 (N_20327,N_16717,N_18569);
xor U20328 (N_20328,N_16636,N_16424);
nor U20329 (N_20329,N_15843,N_16008);
nand U20330 (N_20330,N_16605,N_17298);
nand U20331 (N_20331,N_17284,N_18341);
nand U20332 (N_20332,N_16286,N_18393);
nor U20333 (N_20333,N_16076,N_18216);
nor U20334 (N_20334,N_16994,N_17744);
nor U20335 (N_20335,N_15738,N_17988);
nor U20336 (N_20336,N_18491,N_16420);
or U20337 (N_20337,N_16158,N_16729);
nor U20338 (N_20338,N_16515,N_15660);
nand U20339 (N_20339,N_16418,N_15986);
nor U20340 (N_20340,N_16574,N_18668);
and U20341 (N_20341,N_16435,N_16244);
or U20342 (N_20342,N_17258,N_16024);
nor U20343 (N_20343,N_16607,N_15708);
or U20344 (N_20344,N_17290,N_17458);
nand U20345 (N_20345,N_18243,N_16071);
nor U20346 (N_20346,N_18662,N_16788);
nor U20347 (N_20347,N_15815,N_16131);
nor U20348 (N_20348,N_18353,N_18588);
and U20349 (N_20349,N_18525,N_16285);
and U20350 (N_20350,N_15818,N_18554);
nor U20351 (N_20351,N_16685,N_15907);
nor U20352 (N_20352,N_16439,N_17797);
and U20353 (N_20353,N_18223,N_17417);
and U20354 (N_20354,N_16068,N_18318);
and U20355 (N_20355,N_18586,N_18651);
or U20356 (N_20356,N_17813,N_16969);
nor U20357 (N_20357,N_16725,N_15739);
nand U20358 (N_20358,N_17332,N_17073);
nor U20359 (N_20359,N_16433,N_16083);
nand U20360 (N_20360,N_18229,N_16691);
nor U20361 (N_20361,N_17510,N_18689);
nand U20362 (N_20362,N_17806,N_17092);
or U20363 (N_20363,N_16766,N_17274);
and U20364 (N_20364,N_15703,N_18198);
and U20365 (N_20365,N_18271,N_17734);
or U20366 (N_20366,N_18703,N_16608);
or U20367 (N_20367,N_18412,N_15991);
nor U20368 (N_20368,N_17577,N_15809);
nand U20369 (N_20369,N_18251,N_16243);
and U20370 (N_20370,N_17697,N_15871);
xnor U20371 (N_20371,N_17137,N_16393);
nor U20372 (N_20372,N_18378,N_15770);
xnor U20373 (N_20373,N_17542,N_17705);
xor U20374 (N_20374,N_16274,N_16153);
and U20375 (N_20375,N_17023,N_16770);
and U20376 (N_20376,N_16537,N_16561);
or U20377 (N_20377,N_17396,N_16546);
or U20378 (N_20378,N_16261,N_18307);
nor U20379 (N_20379,N_18358,N_17033);
nor U20380 (N_20380,N_16705,N_17852);
and U20381 (N_20381,N_18054,N_16074);
and U20382 (N_20382,N_16183,N_16487);
nand U20383 (N_20383,N_16802,N_17535);
and U20384 (N_20384,N_16989,N_18612);
xor U20385 (N_20385,N_18563,N_18056);
and U20386 (N_20386,N_17747,N_16243);
and U20387 (N_20387,N_16759,N_15789);
or U20388 (N_20388,N_18311,N_16408);
nand U20389 (N_20389,N_15731,N_17813);
and U20390 (N_20390,N_18428,N_17585);
or U20391 (N_20391,N_18715,N_16446);
or U20392 (N_20392,N_16037,N_16831);
or U20393 (N_20393,N_16902,N_16061);
nor U20394 (N_20394,N_18696,N_17755);
and U20395 (N_20395,N_18112,N_18291);
nand U20396 (N_20396,N_17446,N_17086);
nor U20397 (N_20397,N_16235,N_17548);
and U20398 (N_20398,N_15778,N_18234);
xnor U20399 (N_20399,N_17983,N_15738);
and U20400 (N_20400,N_16194,N_16674);
and U20401 (N_20401,N_16677,N_18656);
nand U20402 (N_20402,N_17569,N_17089);
nand U20403 (N_20403,N_16428,N_17066);
nand U20404 (N_20404,N_17949,N_16385);
nand U20405 (N_20405,N_18047,N_17526);
nand U20406 (N_20406,N_18668,N_16631);
or U20407 (N_20407,N_17142,N_16929);
xor U20408 (N_20408,N_17646,N_15785);
and U20409 (N_20409,N_17256,N_17301);
nand U20410 (N_20410,N_16517,N_18603);
and U20411 (N_20411,N_15723,N_17507);
or U20412 (N_20412,N_16683,N_18334);
or U20413 (N_20413,N_15979,N_15726);
or U20414 (N_20414,N_16536,N_15999);
nand U20415 (N_20415,N_17949,N_16180);
nor U20416 (N_20416,N_18497,N_16591);
and U20417 (N_20417,N_16827,N_18351);
nor U20418 (N_20418,N_16847,N_16494);
and U20419 (N_20419,N_15652,N_16612);
nand U20420 (N_20420,N_17440,N_16556);
nor U20421 (N_20421,N_16349,N_16799);
nand U20422 (N_20422,N_17829,N_16115);
or U20423 (N_20423,N_18487,N_17347);
or U20424 (N_20424,N_18713,N_17412);
or U20425 (N_20425,N_18631,N_17223);
nor U20426 (N_20426,N_17176,N_18729);
nor U20427 (N_20427,N_15855,N_17616);
nor U20428 (N_20428,N_17491,N_16841);
nand U20429 (N_20429,N_17711,N_16078);
or U20430 (N_20430,N_16427,N_18369);
and U20431 (N_20431,N_15968,N_18248);
nor U20432 (N_20432,N_15645,N_16225);
or U20433 (N_20433,N_17226,N_16503);
nand U20434 (N_20434,N_17699,N_17135);
xnor U20435 (N_20435,N_16414,N_15626);
and U20436 (N_20436,N_15838,N_15654);
xnor U20437 (N_20437,N_16387,N_17620);
nand U20438 (N_20438,N_15878,N_17654);
nand U20439 (N_20439,N_18152,N_15992);
and U20440 (N_20440,N_16273,N_15919);
nand U20441 (N_20441,N_18192,N_17024);
nand U20442 (N_20442,N_18719,N_16101);
and U20443 (N_20443,N_17648,N_17401);
and U20444 (N_20444,N_16816,N_17531);
or U20445 (N_20445,N_18717,N_16097);
or U20446 (N_20446,N_17498,N_18267);
nor U20447 (N_20447,N_16729,N_18372);
and U20448 (N_20448,N_17604,N_16207);
or U20449 (N_20449,N_17492,N_16213);
nor U20450 (N_20450,N_18435,N_16875);
and U20451 (N_20451,N_16461,N_18618);
nor U20452 (N_20452,N_18319,N_17368);
xnor U20453 (N_20453,N_18565,N_17208);
nor U20454 (N_20454,N_16277,N_15729);
nand U20455 (N_20455,N_18455,N_16481);
or U20456 (N_20456,N_16404,N_18648);
nor U20457 (N_20457,N_16299,N_16068);
nor U20458 (N_20458,N_15655,N_18590);
and U20459 (N_20459,N_18595,N_17980);
nand U20460 (N_20460,N_17399,N_17840);
xor U20461 (N_20461,N_18745,N_16664);
and U20462 (N_20462,N_16143,N_17576);
nor U20463 (N_20463,N_16997,N_17605);
nor U20464 (N_20464,N_16799,N_17767);
xor U20465 (N_20465,N_18264,N_17900);
or U20466 (N_20466,N_18054,N_18294);
nand U20467 (N_20467,N_18015,N_16011);
or U20468 (N_20468,N_18396,N_17657);
xnor U20469 (N_20469,N_16254,N_15867);
or U20470 (N_20470,N_17233,N_15833);
nor U20471 (N_20471,N_15650,N_16881);
and U20472 (N_20472,N_18623,N_17869);
nor U20473 (N_20473,N_16498,N_16224);
nor U20474 (N_20474,N_16849,N_18337);
nor U20475 (N_20475,N_16907,N_18468);
nand U20476 (N_20476,N_15732,N_18303);
xnor U20477 (N_20477,N_16844,N_16665);
nand U20478 (N_20478,N_16663,N_15641);
and U20479 (N_20479,N_17517,N_18466);
nor U20480 (N_20480,N_17935,N_16367);
or U20481 (N_20481,N_18599,N_17774);
and U20482 (N_20482,N_18355,N_17132);
nand U20483 (N_20483,N_16363,N_17910);
nor U20484 (N_20484,N_18166,N_18379);
or U20485 (N_20485,N_17224,N_17390);
nor U20486 (N_20486,N_16038,N_17630);
xor U20487 (N_20487,N_15856,N_17639);
nor U20488 (N_20488,N_18450,N_18749);
nor U20489 (N_20489,N_17601,N_17755);
nor U20490 (N_20490,N_18501,N_16487);
nor U20491 (N_20491,N_17997,N_15916);
or U20492 (N_20492,N_16877,N_16184);
or U20493 (N_20493,N_15862,N_18269);
or U20494 (N_20494,N_17219,N_15740);
and U20495 (N_20495,N_16744,N_17647);
or U20496 (N_20496,N_18075,N_16658);
nor U20497 (N_20497,N_16650,N_17483);
xor U20498 (N_20498,N_18560,N_17925);
xor U20499 (N_20499,N_17107,N_18191);
nor U20500 (N_20500,N_16358,N_18374);
nand U20501 (N_20501,N_17943,N_15924);
or U20502 (N_20502,N_17416,N_16027);
and U20503 (N_20503,N_15890,N_15976);
and U20504 (N_20504,N_16908,N_15993);
nand U20505 (N_20505,N_15710,N_16779);
and U20506 (N_20506,N_16286,N_16189);
and U20507 (N_20507,N_18122,N_18002);
and U20508 (N_20508,N_17822,N_18329);
or U20509 (N_20509,N_17843,N_16180);
or U20510 (N_20510,N_18164,N_16035);
nor U20511 (N_20511,N_18181,N_15903);
and U20512 (N_20512,N_17858,N_16367);
or U20513 (N_20513,N_16101,N_18386);
nor U20514 (N_20514,N_16273,N_18358);
nor U20515 (N_20515,N_16522,N_18015);
and U20516 (N_20516,N_17886,N_16011);
or U20517 (N_20517,N_18486,N_15736);
or U20518 (N_20518,N_16425,N_18153);
nand U20519 (N_20519,N_18127,N_15936);
and U20520 (N_20520,N_17952,N_16500);
and U20521 (N_20521,N_17874,N_16067);
and U20522 (N_20522,N_17539,N_17119);
nor U20523 (N_20523,N_16910,N_15719);
and U20524 (N_20524,N_15639,N_17427);
nor U20525 (N_20525,N_15881,N_16532);
nand U20526 (N_20526,N_17525,N_17032);
nand U20527 (N_20527,N_17063,N_18666);
nand U20528 (N_20528,N_17604,N_18502);
or U20529 (N_20529,N_16952,N_17337);
or U20530 (N_20530,N_15759,N_17205);
nand U20531 (N_20531,N_17687,N_17321);
or U20532 (N_20532,N_15848,N_17203);
or U20533 (N_20533,N_15897,N_18360);
and U20534 (N_20534,N_18211,N_15941);
nor U20535 (N_20535,N_15803,N_16428);
or U20536 (N_20536,N_16583,N_17837);
and U20537 (N_20537,N_16334,N_15866);
nand U20538 (N_20538,N_18708,N_16318);
or U20539 (N_20539,N_16545,N_16151);
nor U20540 (N_20540,N_16388,N_17612);
nand U20541 (N_20541,N_15828,N_16189);
xnor U20542 (N_20542,N_17810,N_15947);
nor U20543 (N_20543,N_17367,N_17619);
nand U20544 (N_20544,N_15897,N_17565);
nor U20545 (N_20545,N_18492,N_18630);
and U20546 (N_20546,N_18403,N_16823);
or U20547 (N_20547,N_17154,N_16646);
nor U20548 (N_20548,N_16062,N_16750);
and U20549 (N_20549,N_17400,N_16991);
and U20550 (N_20550,N_18029,N_17369);
nand U20551 (N_20551,N_16917,N_17860);
nor U20552 (N_20552,N_15947,N_16522);
nor U20553 (N_20553,N_16525,N_15773);
or U20554 (N_20554,N_17365,N_16552);
or U20555 (N_20555,N_16695,N_16541);
nor U20556 (N_20556,N_16639,N_18746);
and U20557 (N_20557,N_18180,N_18056);
nand U20558 (N_20558,N_16613,N_16422);
or U20559 (N_20559,N_18385,N_16230);
nor U20560 (N_20560,N_17371,N_18411);
or U20561 (N_20561,N_18418,N_16016);
nor U20562 (N_20562,N_18288,N_16118);
or U20563 (N_20563,N_16973,N_16066);
nor U20564 (N_20564,N_17915,N_18015);
xor U20565 (N_20565,N_16759,N_18164);
or U20566 (N_20566,N_16274,N_16555);
and U20567 (N_20567,N_16251,N_17540);
nor U20568 (N_20568,N_15937,N_18517);
or U20569 (N_20569,N_16659,N_15741);
nand U20570 (N_20570,N_17679,N_17722);
or U20571 (N_20571,N_16653,N_15667);
nand U20572 (N_20572,N_17491,N_17717);
nand U20573 (N_20573,N_16346,N_16627);
nor U20574 (N_20574,N_15690,N_16728);
nor U20575 (N_20575,N_16975,N_16282);
nand U20576 (N_20576,N_17803,N_17498);
nor U20577 (N_20577,N_17132,N_15821);
xor U20578 (N_20578,N_16759,N_16057);
and U20579 (N_20579,N_17769,N_18114);
or U20580 (N_20580,N_16576,N_18118);
and U20581 (N_20581,N_15795,N_16875);
and U20582 (N_20582,N_17577,N_17996);
and U20583 (N_20583,N_16511,N_17020);
nand U20584 (N_20584,N_16099,N_18605);
and U20585 (N_20585,N_17642,N_16287);
xnor U20586 (N_20586,N_16946,N_18097);
or U20587 (N_20587,N_16237,N_17701);
or U20588 (N_20588,N_16862,N_17412);
nand U20589 (N_20589,N_16741,N_16047);
nand U20590 (N_20590,N_18265,N_16575);
and U20591 (N_20591,N_17917,N_17482);
nand U20592 (N_20592,N_15826,N_16800);
or U20593 (N_20593,N_16253,N_18391);
nor U20594 (N_20594,N_18307,N_17553);
or U20595 (N_20595,N_18357,N_17455);
nand U20596 (N_20596,N_16185,N_15725);
xnor U20597 (N_20597,N_15933,N_17807);
nand U20598 (N_20598,N_17344,N_17035);
and U20599 (N_20599,N_15797,N_18100);
nand U20600 (N_20600,N_17321,N_17550);
nand U20601 (N_20601,N_18050,N_16692);
nand U20602 (N_20602,N_17913,N_17651);
or U20603 (N_20603,N_17914,N_18096);
nor U20604 (N_20604,N_17371,N_16373);
xnor U20605 (N_20605,N_17869,N_17419);
or U20606 (N_20606,N_17110,N_17767);
nand U20607 (N_20607,N_18417,N_17792);
nor U20608 (N_20608,N_16508,N_15721);
nor U20609 (N_20609,N_16653,N_18594);
xor U20610 (N_20610,N_17080,N_16220);
or U20611 (N_20611,N_15774,N_16808);
and U20612 (N_20612,N_15984,N_16925);
nor U20613 (N_20613,N_16278,N_16090);
or U20614 (N_20614,N_16860,N_17111);
or U20615 (N_20615,N_17601,N_16033);
or U20616 (N_20616,N_17976,N_16123);
and U20617 (N_20617,N_18199,N_16446);
nand U20618 (N_20618,N_16782,N_16412);
nor U20619 (N_20619,N_17660,N_18244);
nand U20620 (N_20620,N_18559,N_17289);
nor U20621 (N_20621,N_17818,N_17949);
nor U20622 (N_20622,N_16494,N_15958);
or U20623 (N_20623,N_17296,N_17539);
or U20624 (N_20624,N_18084,N_16342);
and U20625 (N_20625,N_18247,N_16636);
and U20626 (N_20626,N_17380,N_16610);
or U20627 (N_20627,N_15739,N_16228);
nor U20628 (N_20628,N_18460,N_16120);
and U20629 (N_20629,N_17805,N_18202);
and U20630 (N_20630,N_16773,N_18647);
or U20631 (N_20631,N_15794,N_17825);
or U20632 (N_20632,N_17162,N_15812);
nor U20633 (N_20633,N_16180,N_16679);
and U20634 (N_20634,N_16099,N_16277);
and U20635 (N_20635,N_17851,N_18059);
nor U20636 (N_20636,N_17390,N_18250);
or U20637 (N_20637,N_16453,N_17499);
xnor U20638 (N_20638,N_17712,N_15716);
nand U20639 (N_20639,N_16642,N_18154);
or U20640 (N_20640,N_17425,N_18530);
nand U20641 (N_20641,N_18113,N_17616);
nor U20642 (N_20642,N_15942,N_15864);
and U20643 (N_20643,N_17781,N_18287);
and U20644 (N_20644,N_16685,N_16792);
and U20645 (N_20645,N_18305,N_15967);
or U20646 (N_20646,N_16224,N_18144);
nand U20647 (N_20647,N_15638,N_15976);
nand U20648 (N_20648,N_18276,N_16053);
and U20649 (N_20649,N_15811,N_15671);
nor U20650 (N_20650,N_17570,N_18107);
or U20651 (N_20651,N_18190,N_18168);
or U20652 (N_20652,N_18429,N_18648);
or U20653 (N_20653,N_16790,N_16589);
and U20654 (N_20654,N_18441,N_18422);
xor U20655 (N_20655,N_18195,N_18413);
xnor U20656 (N_20656,N_16692,N_17059);
or U20657 (N_20657,N_17311,N_17946);
or U20658 (N_20658,N_17866,N_16827);
or U20659 (N_20659,N_17373,N_18681);
or U20660 (N_20660,N_18736,N_15790);
nor U20661 (N_20661,N_17974,N_17820);
or U20662 (N_20662,N_17355,N_16262);
or U20663 (N_20663,N_15905,N_17534);
nor U20664 (N_20664,N_16224,N_17503);
and U20665 (N_20665,N_15800,N_18280);
and U20666 (N_20666,N_18243,N_16999);
nor U20667 (N_20667,N_18216,N_15909);
or U20668 (N_20668,N_18727,N_17419);
nor U20669 (N_20669,N_16652,N_16380);
nand U20670 (N_20670,N_15727,N_15668);
nand U20671 (N_20671,N_15754,N_18607);
nand U20672 (N_20672,N_18711,N_17861);
or U20673 (N_20673,N_15631,N_16544);
and U20674 (N_20674,N_18657,N_17019);
nor U20675 (N_20675,N_16842,N_17983);
nor U20676 (N_20676,N_17408,N_17438);
or U20677 (N_20677,N_18534,N_15861);
nor U20678 (N_20678,N_17724,N_15976);
nand U20679 (N_20679,N_17757,N_17361);
nand U20680 (N_20680,N_17454,N_17057);
and U20681 (N_20681,N_18351,N_18447);
nor U20682 (N_20682,N_17720,N_16683);
and U20683 (N_20683,N_16613,N_17560);
or U20684 (N_20684,N_17008,N_17457);
nor U20685 (N_20685,N_17725,N_17524);
or U20686 (N_20686,N_16452,N_16320);
nor U20687 (N_20687,N_17862,N_16994);
xor U20688 (N_20688,N_16206,N_16372);
and U20689 (N_20689,N_16864,N_16725);
nand U20690 (N_20690,N_18066,N_18401);
and U20691 (N_20691,N_17568,N_15733);
and U20692 (N_20692,N_16425,N_17617);
and U20693 (N_20693,N_17617,N_16072);
xnor U20694 (N_20694,N_17214,N_18178);
or U20695 (N_20695,N_17305,N_18575);
nand U20696 (N_20696,N_16355,N_16382);
nor U20697 (N_20697,N_16355,N_18005);
nor U20698 (N_20698,N_16886,N_18440);
and U20699 (N_20699,N_16850,N_17836);
nor U20700 (N_20700,N_18448,N_18358);
nor U20701 (N_20701,N_16006,N_18644);
nor U20702 (N_20702,N_18472,N_16660);
nand U20703 (N_20703,N_15981,N_17288);
nor U20704 (N_20704,N_16545,N_18669);
and U20705 (N_20705,N_18232,N_18692);
nor U20706 (N_20706,N_16051,N_16665);
or U20707 (N_20707,N_17395,N_16206);
nor U20708 (N_20708,N_17087,N_16315);
nand U20709 (N_20709,N_17897,N_17881);
nand U20710 (N_20710,N_18535,N_18628);
or U20711 (N_20711,N_17679,N_16306);
and U20712 (N_20712,N_16265,N_16058);
nand U20713 (N_20713,N_17401,N_17912);
xnor U20714 (N_20714,N_18672,N_15749);
nand U20715 (N_20715,N_17477,N_16244);
nand U20716 (N_20716,N_16974,N_15696);
or U20717 (N_20717,N_18030,N_17562);
nor U20718 (N_20718,N_18633,N_16706);
xnor U20719 (N_20719,N_15763,N_17839);
and U20720 (N_20720,N_17274,N_16295);
nand U20721 (N_20721,N_18324,N_18307);
and U20722 (N_20722,N_16401,N_17000);
nand U20723 (N_20723,N_18282,N_18535);
nor U20724 (N_20724,N_16337,N_16804);
or U20725 (N_20725,N_18275,N_15646);
and U20726 (N_20726,N_15822,N_16017);
or U20727 (N_20727,N_17838,N_16635);
and U20728 (N_20728,N_17671,N_16893);
nand U20729 (N_20729,N_15780,N_15954);
nand U20730 (N_20730,N_17151,N_16096);
or U20731 (N_20731,N_15714,N_15966);
or U20732 (N_20732,N_16870,N_17033);
nor U20733 (N_20733,N_17079,N_15800);
nand U20734 (N_20734,N_16033,N_15847);
or U20735 (N_20735,N_17889,N_16928);
nand U20736 (N_20736,N_15712,N_18163);
nand U20737 (N_20737,N_17615,N_17493);
nor U20738 (N_20738,N_17900,N_15921);
or U20739 (N_20739,N_16284,N_18727);
nand U20740 (N_20740,N_17115,N_17587);
nor U20741 (N_20741,N_17554,N_18297);
and U20742 (N_20742,N_17507,N_18349);
nor U20743 (N_20743,N_16158,N_16922);
nand U20744 (N_20744,N_17510,N_18729);
and U20745 (N_20745,N_16135,N_17771);
and U20746 (N_20746,N_15720,N_16080);
nand U20747 (N_20747,N_17614,N_18050);
nor U20748 (N_20748,N_17587,N_17318);
nor U20749 (N_20749,N_15882,N_17391);
and U20750 (N_20750,N_17205,N_16401);
nor U20751 (N_20751,N_17452,N_17274);
nand U20752 (N_20752,N_15898,N_16994);
nand U20753 (N_20753,N_17646,N_18295);
or U20754 (N_20754,N_16590,N_16392);
nand U20755 (N_20755,N_18438,N_16763);
nor U20756 (N_20756,N_17009,N_16393);
and U20757 (N_20757,N_17906,N_15909);
and U20758 (N_20758,N_17891,N_15626);
nand U20759 (N_20759,N_17351,N_16590);
or U20760 (N_20760,N_16216,N_17168);
nor U20761 (N_20761,N_18315,N_18533);
nor U20762 (N_20762,N_16120,N_16392);
xnor U20763 (N_20763,N_16734,N_18655);
nor U20764 (N_20764,N_16593,N_15650);
or U20765 (N_20765,N_18675,N_17808);
nor U20766 (N_20766,N_17623,N_16164);
and U20767 (N_20767,N_17353,N_16485);
nor U20768 (N_20768,N_15914,N_16817);
and U20769 (N_20769,N_17069,N_16451);
nor U20770 (N_20770,N_17360,N_18670);
nand U20771 (N_20771,N_15835,N_18312);
nor U20772 (N_20772,N_18072,N_18284);
nand U20773 (N_20773,N_15840,N_17706);
nand U20774 (N_20774,N_16794,N_18314);
nor U20775 (N_20775,N_17116,N_16944);
nor U20776 (N_20776,N_17682,N_18262);
or U20777 (N_20777,N_18647,N_17088);
or U20778 (N_20778,N_16454,N_18338);
and U20779 (N_20779,N_17239,N_15633);
or U20780 (N_20780,N_18550,N_15719);
and U20781 (N_20781,N_18425,N_17608);
and U20782 (N_20782,N_17342,N_17809);
nand U20783 (N_20783,N_17924,N_17455);
nor U20784 (N_20784,N_17602,N_17485);
and U20785 (N_20785,N_15673,N_17361);
nor U20786 (N_20786,N_17115,N_17708);
or U20787 (N_20787,N_16820,N_18294);
and U20788 (N_20788,N_16115,N_18717);
xnor U20789 (N_20789,N_16908,N_16580);
and U20790 (N_20790,N_15953,N_16661);
and U20791 (N_20791,N_17663,N_16267);
nand U20792 (N_20792,N_15680,N_16733);
nor U20793 (N_20793,N_18583,N_18297);
nand U20794 (N_20794,N_15949,N_18488);
nand U20795 (N_20795,N_18502,N_16224);
nor U20796 (N_20796,N_18720,N_15847);
nand U20797 (N_20797,N_18126,N_18674);
or U20798 (N_20798,N_15735,N_18428);
nand U20799 (N_20799,N_18213,N_16494);
and U20800 (N_20800,N_15891,N_16076);
and U20801 (N_20801,N_18738,N_17068);
nor U20802 (N_20802,N_16907,N_16321);
xnor U20803 (N_20803,N_17889,N_15901);
nand U20804 (N_20804,N_17936,N_17629);
or U20805 (N_20805,N_16507,N_17323);
xor U20806 (N_20806,N_15682,N_18618);
nor U20807 (N_20807,N_17908,N_18611);
xor U20808 (N_20808,N_18215,N_18365);
nor U20809 (N_20809,N_17728,N_16412);
and U20810 (N_20810,N_18163,N_17658);
or U20811 (N_20811,N_16558,N_18559);
nand U20812 (N_20812,N_17603,N_18659);
nand U20813 (N_20813,N_18457,N_17572);
or U20814 (N_20814,N_17661,N_17099);
nor U20815 (N_20815,N_15916,N_18106);
xnor U20816 (N_20816,N_18491,N_16549);
nor U20817 (N_20817,N_16008,N_16795);
or U20818 (N_20818,N_17958,N_17722);
and U20819 (N_20819,N_17092,N_15788);
and U20820 (N_20820,N_16107,N_16392);
or U20821 (N_20821,N_18706,N_17087);
and U20822 (N_20822,N_16775,N_16831);
or U20823 (N_20823,N_18162,N_17208);
and U20824 (N_20824,N_18107,N_17703);
nor U20825 (N_20825,N_17558,N_16735);
and U20826 (N_20826,N_17969,N_18290);
nor U20827 (N_20827,N_18214,N_16793);
xnor U20828 (N_20828,N_16748,N_17322);
and U20829 (N_20829,N_17441,N_16619);
xnor U20830 (N_20830,N_16544,N_15822);
nor U20831 (N_20831,N_16079,N_18514);
nand U20832 (N_20832,N_16086,N_16242);
nor U20833 (N_20833,N_16856,N_18447);
nand U20834 (N_20834,N_17730,N_18208);
or U20835 (N_20835,N_17066,N_16382);
and U20836 (N_20836,N_17369,N_16127);
nor U20837 (N_20837,N_16659,N_17265);
and U20838 (N_20838,N_18506,N_16867);
nor U20839 (N_20839,N_16239,N_16742);
or U20840 (N_20840,N_18011,N_17269);
nor U20841 (N_20841,N_17756,N_17494);
nor U20842 (N_20842,N_15742,N_16206);
or U20843 (N_20843,N_18298,N_17787);
xor U20844 (N_20844,N_17609,N_16360);
or U20845 (N_20845,N_16208,N_16632);
nand U20846 (N_20846,N_16929,N_16652);
xor U20847 (N_20847,N_16163,N_17186);
or U20848 (N_20848,N_16793,N_17479);
nor U20849 (N_20849,N_17503,N_16912);
xnor U20850 (N_20850,N_18026,N_15929);
nor U20851 (N_20851,N_17321,N_17740);
and U20852 (N_20852,N_17166,N_15915);
nand U20853 (N_20853,N_18288,N_17794);
nand U20854 (N_20854,N_18362,N_17368);
nand U20855 (N_20855,N_16954,N_17917);
nor U20856 (N_20856,N_17937,N_18732);
and U20857 (N_20857,N_16869,N_17269);
nand U20858 (N_20858,N_17160,N_17729);
or U20859 (N_20859,N_17027,N_15632);
nand U20860 (N_20860,N_17841,N_17921);
or U20861 (N_20861,N_16500,N_17792);
nor U20862 (N_20862,N_15636,N_18009);
nand U20863 (N_20863,N_17010,N_18310);
nand U20864 (N_20864,N_17003,N_15967);
or U20865 (N_20865,N_18105,N_16597);
and U20866 (N_20866,N_17698,N_17621);
nor U20867 (N_20867,N_17723,N_18206);
or U20868 (N_20868,N_17521,N_16540);
and U20869 (N_20869,N_16260,N_18423);
nor U20870 (N_20870,N_17489,N_16458);
nand U20871 (N_20871,N_16089,N_15932);
nor U20872 (N_20872,N_16442,N_16127);
and U20873 (N_20873,N_18424,N_17421);
nor U20874 (N_20874,N_16211,N_16006);
and U20875 (N_20875,N_17678,N_17105);
nand U20876 (N_20876,N_17002,N_15863);
nor U20877 (N_20877,N_18697,N_16441);
or U20878 (N_20878,N_15686,N_16784);
or U20879 (N_20879,N_17526,N_17287);
or U20880 (N_20880,N_18194,N_16744);
nand U20881 (N_20881,N_17101,N_16628);
nor U20882 (N_20882,N_17874,N_15762);
nor U20883 (N_20883,N_18441,N_16804);
and U20884 (N_20884,N_17915,N_16427);
nor U20885 (N_20885,N_17174,N_15699);
or U20886 (N_20886,N_18604,N_16893);
nor U20887 (N_20887,N_17214,N_17674);
xnor U20888 (N_20888,N_18487,N_18469);
or U20889 (N_20889,N_16555,N_16941);
and U20890 (N_20890,N_17581,N_17550);
nor U20891 (N_20891,N_16573,N_17628);
or U20892 (N_20892,N_16695,N_16230);
or U20893 (N_20893,N_16500,N_17083);
nor U20894 (N_20894,N_17640,N_16713);
xor U20895 (N_20895,N_17550,N_16951);
nor U20896 (N_20896,N_17877,N_16005);
nor U20897 (N_20897,N_18515,N_16828);
and U20898 (N_20898,N_18580,N_16103);
nand U20899 (N_20899,N_16500,N_16612);
nand U20900 (N_20900,N_18076,N_16927);
nand U20901 (N_20901,N_17569,N_16843);
and U20902 (N_20902,N_17387,N_16225);
nand U20903 (N_20903,N_16448,N_15694);
and U20904 (N_20904,N_17435,N_15770);
xnor U20905 (N_20905,N_17120,N_16606);
or U20906 (N_20906,N_18545,N_18068);
and U20907 (N_20907,N_15704,N_18229);
nand U20908 (N_20908,N_17790,N_17610);
and U20909 (N_20909,N_16192,N_17280);
or U20910 (N_20910,N_18081,N_18119);
and U20911 (N_20911,N_16416,N_17898);
or U20912 (N_20912,N_17162,N_16606);
nand U20913 (N_20913,N_16409,N_17913);
nand U20914 (N_20914,N_17490,N_18374);
nor U20915 (N_20915,N_16037,N_16454);
nand U20916 (N_20916,N_18282,N_18429);
and U20917 (N_20917,N_17115,N_18072);
or U20918 (N_20918,N_18267,N_18260);
or U20919 (N_20919,N_17013,N_18023);
and U20920 (N_20920,N_16866,N_18129);
nand U20921 (N_20921,N_17448,N_17395);
nor U20922 (N_20922,N_17384,N_17766);
nor U20923 (N_20923,N_16426,N_17379);
or U20924 (N_20924,N_16334,N_18103);
nor U20925 (N_20925,N_17844,N_16495);
and U20926 (N_20926,N_17792,N_17453);
nor U20927 (N_20927,N_15801,N_16178);
nor U20928 (N_20928,N_18075,N_17113);
or U20929 (N_20929,N_16132,N_16432);
nor U20930 (N_20930,N_18379,N_17074);
xnor U20931 (N_20931,N_16636,N_16782);
nand U20932 (N_20932,N_18087,N_17397);
nand U20933 (N_20933,N_15924,N_17291);
nor U20934 (N_20934,N_16426,N_18178);
xor U20935 (N_20935,N_16127,N_17414);
nor U20936 (N_20936,N_17070,N_17989);
nor U20937 (N_20937,N_16472,N_18264);
or U20938 (N_20938,N_17066,N_18583);
or U20939 (N_20939,N_16116,N_17742);
xnor U20940 (N_20940,N_18020,N_17461);
and U20941 (N_20941,N_16454,N_17491);
and U20942 (N_20942,N_16302,N_16359);
nor U20943 (N_20943,N_16346,N_15993);
and U20944 (N_20944,N_18532,N_18099);
nor U20945 (N_20945,N_16621,N_17381);
nand U20946 (N_20946,N_16089,N_16282);
nand U20947 (N_20947,N_17472,N_16530);
and U20948 (N_20948,N_18081,N_16256);
nor U20949 (N_20949,N_16802,N_17839);
nand U20950 (N_20950,N_17684,N_15688);
nor U20951 (N_20951,N_17599,N_15693);
nor U20952 (N_20952,N_16058,N_18158);
nand U20953 (N_20953,N_17992,N_17358);
nand U20954 (N_20954,N_18634,N_16174);
or U20955 (N_20955,N_15707,N_17428);
xnor U20956 (N_20956,N_16825,N_17123);
nor U20957 (N_20957,N_16043,N_16432);
xnor U20958 (N_20958,N_16223,N_16884);
xnor U20959 (N_20959,N_15946,N_18068);
or U20960 (N_20960,N_15889,N_17918);
nand U20961 (N_20961,N_17846,N_18224);
or U20962 (N_20962,N_15774,N_18148);
nand U20963 (N_20963,N_17126,N_16309);
nor U20964 (N_20964,N_17560,N_18532);
or U20965 (N_20965,N_18016,N_16083);
nor U20966 (N_20966,N_17456,N_15670);
and U20967 (N_20967,N_18722,N_18050);
xor U20968 (N_20968,N_16885,N_17535);
or U20969 (N_20969,N_16346,N_17239);
or U20970 (N_20970,N_17409,N_17625);
or U20971 (N_20971,N_17946,N_16023);
and U20972 (N_20972,N_15647,N_18242);
nor U20973 (N_20973,N_16656,N_15939);
nor U20974 (N_20974,N_17599,N_17161);
nand U20975 (N_20975,N_17763,N_16590);
and U20976 (N_20976,N_16995,N_16810);
or U20977 (N_20977,N_15876,N_17286);
and U20978 (N_20978,N_16950,N_17340);
or U20979 (N_20979,N_16507,N_18609);
xor U20980 (N_20980,N_18356,N_17781);
nand U20981 (N_20981,N_18320,N_15966);
nand U20982 (N_20982,N_15891,N_17016);
and U20983 (N_20983,N_17688,N_15654);
nor U20984 (N_20984,N_18186,N_18546);
and U20985 (N_20985,N_18158,N_15938);
and U20986 (N_20986,N_17054,N_18017);
nor U20987 (N_20987,N_18495,N_17570);
nor U20988 (N_20988,N_16599,N_17032);
nor U20989 (N_20989,N_15822,N_18259);
nand U20990 (N_20990,N_17739,N_16713);
and U20991 (N_20991,N_16991,N_18311);
and U20992 (N_20992,N_15870,N_17429);
nor U20993 (N_20993,N_16005,N_16944);
and U20994 (N_20994,N_17356,N_18166);
nor U20995 (N_20995,N_18405,N_16353);
nand U20996 (N_20996,N_16229,N_18023);
nand U20997 (N_20997,N_16115,N_18334);
xor U20998 (N_20998,N_18636,N_15744);
or U20999 (N_20999,N_15920,N_17329);
xor U21000 (N_21000,N_18036,N_16155);
nand U21001 (N_21001,N_15765,N_16438);
and U21002 (N_21002,N_18689,N_15992);
nor U21003 (N_21003,N_15717,N_18115);
nor U21004 (N_21004,N_18033,N_18597);
nand U21005 (N_21005,N_18287,N_18221);
and U21006 (N_21006,N_17501,N_16002);
or U21007 (N_21007,N_17694,N_17489);
nand U21008 (N_21008,N_17186,N_16824);
and U21009 (N_21009,N_17051,N_18488);
or U21010 (N_21010,N_15920,N_17809);
nand U21011 (N_21011,N_17676,N_15763);
or U21012 (N_21012,N_16231,N_17364);
nand U21013 (N_21013,N_18494,N_17947);
or U21014 (N_21014,N_17933,N_16944);
nor U21015 (N_21015,N_15955,N_17745);
nand U21016 (N_21016,N_17257,N_17845);
or U21017 (N_21017,N_17863,N_17116);
or U21018 (N_21018,N_17703,N_18685);
xnor U21019 (N_21019,N_18090,N_15847);
or U21020 (N_21020,N_16351,N_16438);
nor U21021 (N_21021,N_17664,N_16917);
nand U21022 (N_21022,N_18114,N_18509);
and U21023 (N_21023,N_18127,N_18300);
nor U21024 (N_21024,N_17472,N_18577);
xor U21025 (N_21025,N_17083,N_18326);
or U21026 (N_21026,N_18465,N_18665);
xnor U21027 (N_21027,N_15687,N_15754);
nand U21028 (N_21028,N_15915,N_16164);
nor U21029 (N_21029,N_16272,N_17932);
nor U21030 (N_21030,N_18387,N_17907);
nand U21031 (N_21031,N_18587,N_18579);
nand U21032 (N_21032,N_16213,N_16772);
or U21033 (N_21033,N_18077,N_16730);
nor U21034 (N_21034,N_16053,N_17173);
nor U21035 (N_21035,N_17856,N_18581);
xor U21036 (N_21036,N_18087,N_17276);
and U21037 (N_21037,N_18549,N_17436);
and U21038 (N_21038,N_15636,N_16705);
nand U21039 (N_21039,N_16530,N_15883);
and U21040 (N_21040,N_16130,N_16325);
and U21041 (N_21041,N_18126,N_17851);
nand U21042 (N_21042,N_17545,N_17277);
and U21043 (N_21043,N_17626,N_15752);
nor U21044 (N_21044,N_18327,N_17119);
nand U21045 (N_21045,N_17382,N_15966);
nor U21046 (N_21046,N_16806,N_16395);
or U21047 (N_21047,N_16532,N_16486);
and U21048 (N_21048,N_16514,N_18577);
nand U21049 (N_21049,N_15806,N_16440);
and U21050 (N_21050,N_16106,N_16807);
xor U21051 (N_21051,N_17017,N_15894);
xor U21052 (N_21052,N_17678,N_16994);
xor U21053 (N_21053,N_17089,N_15733);
nand U21054 (N_21054,N_18575,N_16370);
nor U21055 (N_21055,N_17130,N_17564);
nor U21056 (N_21056,N_17407,N_16797);
or U21057 (N_21057,N_16825,N_18194);
nand U21058 (N_21058,N_16199,N_15683);
and U21059 (N_21059,N_16631,N_18683);
or U21060 (N_21060,N_16961,N_18452);
nand U21061 (N_21061,N_16473,N_17833);
xnor U21062 (N_21062,N_18333,N_18503);
and U21063 (N_21063,N_15649,N_17706);
nor U21064 (N_21064,N_16758,N_16200);
and U21065 (N_21065,N_16149,N_16009);
or U21066 (N_21066,N_17213,N_15931);
and U21067 (N_21067,N_16540,N_16978);
and U21068 (N_21068,N_17379,N_18453);
or U21069 (N_21069,N_16593,N_17525);
or U21070 (N_21070,N_15877,N_16763);
or U21071 (N_21071,N_16868,N_16435);
nor U21072 (N_21072,N_18363,N_16598);
nand U21073 (N_21073,N_15792,N_17650);
nor U21074 (N_21074,N_17866,N_17118);
or U21075 (N_21075,N_17981,N_16816);
and U21076 (N_21076,N_17772,N_16324);
xnor U21077 (N_21077,N_16135,N_18052);
nand U21078 (N_21078,N_16103,N_16133);
xor U21079 (N_21079,N_16950,N_17113);
nor U21080 (N_21080,N_15973,N_18331);
or U21081 (N_21081,N_17843,N_17683);
and U21082 (N_21082,N_16527,N_17090);
or U21083 (N_21083,N_18453,N_17190);
xor U21084 (N_21084,N_18656,N_16564);
and U21085 (N_21085,N_15656,N_16741);
xnor U21086 (N_21086,N_17125,N_16962);
and U21087 (N_21087,N_17886,N_16682);
nand U21088 (N_21088,N_16887,N_18023);
nand U21089 (N_21089,N_17024,N_17190);
nand U21090 (N_21090,N_17529,N_18189);
nand U21091 (N_21091,N_17277,N_18458);
nand U21092 (N_21092,N_17050,N_16333);
and U21093 (N_21093,N_16786,N_16142);
nand U21094 (N_21094,N_15979,N_17871);
or U21095 (N_21095,N_17792,N_17120);
nand U21096 (N_21096,N_17734,N_16540);
nand U21097 (N_21097,N_17745,N_16751);
and U21098 (N_21098,N_17998,N_17780);
nor U21099 (N_21099,N_15891,N_17999);
and U21100 (N_21100,N_17806,N_18609);
and U21101 (N_21101,N_16437,N_16833);
nor U21102 (N_21102,N_16204,N_18107);
nand U21103 (N_21103,N_18618,N_18450);
or U21104 (N_21104,N_18062,N_17388);
xnor U21105 (N_21105,N_17703,N_15709);
nor U21106 (N_21106,N_17651,N_17966);
nand U21107 (N_21107,N_17765,N_17634);
nand U21108 (N_21108,N_16076,N_17356);
nand U21109 (N_21109,N_17108,N_17285);
and U21110 (N_21110,N_18289,N_16791);
nand U21111 (N_21111,N_17061,N_18451);
nand U21112 (N_21112,N_15682,N_15884);
or U21113 (N_21113,N_18316,N_15768);
or U21114 (N_21114,N_16036,N_18120);
or U21115 (N_21115,N_16620,N_15775);
nand U21116 (N_21116,N_16964,N_18177);
xor U21117 (N_21117,N_17689,N_16565);
xnor U21118 (N_21118,N_15969,N_16848);
nor U21119 (N_21119,N_16694,N_17579);
or U21120 (N_21120,N_17404,N_16780);
nor U21121 (N_21121,N_18283,N_17846);
nor U21122 (N_21122,N_16533,N_18577);
nand U21123 (N_21123,N_16668,N_18437);
nor U21124 (N_21124,N_17434,N_17188);
and U21125 (N_21125,N_18248,N_17257);
or U21126 (N_21126,N_16107,N_16517);
or U21127 (N_21127,N_16075,N_16179);
or U21128 (N_21128,N_16015,N_17731);
nor U21129 (N_21129,N_17643,N_18124);
xnor U21130 (N_21130,N_16719,N_16173);
nand U21131 (N_21131,N_16885,N_18208);
and U21132 (N_21132,N_15935,N_17742);
nand U21133 (N_21133,N_17695,N_16814);
or U21134 (N_21134,N_18428,N_16070);
xnor U21135 (N_21135,N_16148,N_15653);
nor U21136 (N_21136,N_17909,N_16526);
nand U21137 (N_21137,N_18514,N_16459);
or U21138 (N_21138,N_16775,N_18138);
nor U21139 (N_21139,N_15969,N_17554);
and U21140 (N_21140,N_17654,N_16494);
and U21141 (N_21141,N_16309,N_18112);
and U21142 (N_21142,N_16402,N_17385);
or U21143 (N_21143,N_18285,N_16245);
nor U21144 (N_21144,N_17490,N_18008);
nor U21145 (N_21145,N_17531,N_16517);
nand U21146 (N_21146,N_18640,N_17979);
or U21147 (N_21147,N_15859,N_17087);
or U21148 (N_21148,N_17285,N_16939);
nor U21149 (N_21149,N_16238,N_18258);
nand U21150 (N_21150,N_17905,N_18153);
and U21151 (N_21151,N_17956,N_16692);
nand U21152 (N_21152,N_18203,N_18046);
nand U21153 (N_21153,N_17204,N_16560);
nor U21154 (N_21154,N_17980,N_17561);
nor U21155 (N_21155,N_18232,N_16937);
and U21156 (N_21156,N_18204,N_17998);
nor U21157 (N_21157,N_16791,N_17539);
nor U21158 (N_21158,N_17336,N_15951);
nand U21159 (N_21159,N_16180,N_17182);
or U21160 (N_21160,N_16189,N_16222);
nand U21161 (N_21161,N_16995,N_17754);
nor U21162 (N_21162,N_17639,N_18375);
nand U21163 (N_21163,N_16774,N_15660);
or U21164 (N_21164,N_18556,N_18466);
and U21165 (N_21165,N_16358,N_17498);
or U21166 (N_21166,N_16467,N_17812);
nor U21167 (N_21167,N_17109,N_17795);
or U21168 (N_21168,N_16858,N_18571);
nor U21169 (N_21169,N_16130,N_18245);
or U21170 (N_21170,N_16344,N_15843);
or U21171 (N_21171,N_17670,N_15902);
nand U21172 (N_21172,N_16000,N_17924);
nor U21173 (N_21173,N_16753,N_18129);
or U21174 (N_21174,N_17509,N_16219);
nor U21175 (N_21175,N_17662,N_16737);
nand U21176 (N_21176,N_17407,N_17778);
nor U21177 (N_21177,N_16601,N_17547);
and U21178 (N_21178,N_16151,N_17029);
nand U21179 (N_21179,N_16143,N_18554);
nor U21180 (N_21180,N_18652,N_16289);
xor U21181 (N_21181,N_17926,N_15930);
and U21182 (N_21182,N_15807,N_16030);
nor U21183 (N_21183,N_17786,N_17199);
or U21184 (N_21184,N_17924,N_17951);
and U21185 (N_21185,N_18513,N_16019);
or U21186 (N_21186,N_17281,N_16051);
or U21187 (N_21187,N_18405,N_18571);
and U21188 (N_21188,N_18321,N_16880);
nor U21189 (N_21189,N_16645,N_16027);
nand U21190 (N_21190,N_17600,N_16363);
nor U21191 (N_21191,N_16571,N_16038);
and U21192 (N_21192,N_18070,N_17243);
or U21193 (N_21193,N_15986,N_16177);
nand U21194 (N_21194,N_17598,N_17578);
or U21195 (N_21195,N_15887,N_17265);
nor U21196 (N_21196,N_16705,N_16711);
and U21197 (N_21197,N_18577,N_18119);
and U21198 (N_21198,N_16753,N_16012);
nand U21199 (N_21199,N_18285,N_16553);
nand U21200 (N_21200,N_16552,N_16544);
nand U21201 (N_21201,N_17014,N_18595);
and U21202 (N_21202,N_18271,N_18244);
nand U21203 (N_21203,N_18028,N_18232);
nor U21204 (N_21204,N_15835,N_15836);
xor U21205 (N_21205,N_17461,N_15799);
nand U21206 (N_21206,N_18311,N_16664);
nor U21207 (N_21207,N_18339,N_16823);
or U21208 (N_21208,N_16852,N_16659);
nand U21209 (N_21209,N_16635,N_17017);
nand U21210 (N_21210,N_16789,N_16703);
nand U21211 (N_21211,N_17496,N_18135);
nor U21212 (N_21212,N_15940,N_16861);
nand U21213 (N_21213,N_17580,N_15807);
and U21214 (N_21214,N_15825,N_18636);
or U21215 (N_21215,N_18596,N_16136);
xor U21216 (N_21216,N_18269,N_16558);
nor U21217 (N_21217,N_17420,N_16911);
and U21218 (N_21218,N_18340,N_15989);
nor U21219 (N_21219,N_18143,N_16188);
nand U21220 (N_21220,N_18095,N_15956);
nor U21221 (N_21221,N_18431,N_16218);
nor U21222 (N_21222,N_18487,N_16693);
nand U21223 (N_21223,N_18679,N_16070);
nor U21224 (N_21224,N_16875,N_18606);
nor U21225 (N_21225,N_18285,N_16578);
nor U21226 (N_21226,N_15749,N_18430);
or U21227 (N_21227,N_18629,N_17357);
nand U21228 (N_21228,N_17438,N_17295);
nand U21229 (N_21229,N_18029,N_18698);
nand U21230 (N_21230,N_15772,N_16393);
or U21231 (N_21231,N_16836,N_17019);
nand U21232 (N_21232,N_18373,N_15636);
nand U21233 (N_21233,N_18069,N_16322);
and U21234 (N_21234,N_16674,N_15780);
nand U21235 (N_21235,N_18341,N_17370);
nor U21236 (N_21236,N_18418,N_18377);
or U21237 (N_21237,N_18496,N_16119);
nand U21238 (N_21238,N_18731,N_17215);
nand U21239 (N_21239,N_17533,N_18713);
nand U21240 (N_21240,N_18276,N_17713);
or U21241 (N_21241,N_16593,N_17528);
nand U21242 (N_21242,N_18323,N_16153);
xnor U21243 (N_21243,N_17939,N_16037);
or U21244 (N_21244,N_16467,N_17326);
or U21245 (N_21245,N_16780,N_15639);
or U21246 (N_21246,N_17788,N_16706);
nand U21247 (N_21247,N_17164,N_17921);
or U21248 (N_21248,N_16678,N_17220);
nor U21249 (N_21249,N_18107,N_16479);
xnor U21250 (N_21250,N_17944,N_17221);
or U21251 (N_21251,N_16557,N_15685);
xor U21252 (N_21252,N_18191,N_17353);
or U21253 (N_21253,N_17628,N_17716);
nor U21254 (N_21254,N_16228,N_16990);
nand U21255 (N_21255,N_17357,N_18339);
nor U21256 (N_21256,N_17335,N_18010);
and U21257 (N_21257,N_16653,N_16548);
or U21258 (N_21258,N_15645,N_17905);
or U21259 (N_21259,N_17983,N_16847);
or U21260 (N_21260,N_16483,N_16639);
and U21261 (N_21261,N_17064,N_18161);
nor U21262 (N_21262,N_17262,N_16413);
or U21263 (N_21263,N_15884,N_16985);
or U21264 (N_21264,N_18503,N_18443);
and U21265 (N_21265,N_18134,N_15933);
or U21266 (N_21266,N_18280,N_18302);
nor U21267 (N_21267,N_16659,N_15696);
or U21268 (N_21268,N_18245,N_18064);
nand U21269 (N_21269,N_17275,N_16086);
and U21270 (N_21270,N_15808,N_18135);
and U21271 (N_21271,N_18648,N_16270);
and U21272 (N_21272,N_15993,N_16168);
nor U21273 (N_21273,N_17983,N_16505);
nor U21274 (N_21274,N_18449,N_16049);
nand U21275 (N_21275,N_17024,N_17039);
and U21276 (N_21276,N_16000,N_18350);
nand U21277 (N_21277,N_17428,N_17564);
nand U21278 (N_21278,N_15935,N_18042);
or U21279 (N_21279,N_17041,N_17902);
nand U21280 (N_21280,N_18692,N_17927);
and U21281 (N_21281,N_17852,N_16875);
and U21282 (N_21282,N_15827,N_17965);
or U21283 (N_21283,N_16712,N_16616);
nand U21284 (N_21284,N_18520,N_16065);
and U21285 (N_21285,N_17591,N_17439);
nor U21286 (N_21286,N_16436,N_17187);
nor U21287 (N_21287,N_17833,N_18110);
or U21288 (N_21288,N_16219,N_17562);
or U21289 (N_21289,N_16531,N_18720);
nand U21290 (N_21290,N_15711,N_18434);
nand U21291 (N_21291,N_16430,N_17928);
nand U21292 (N_21292,N_16270,N_18159);
xnor U21293 (N_21293,N_17309,N_17601);
or U21294 (N_21294,N_16691,N_18327);
nand U21295 (N_21295,N_16665,N_17150);
or U21296 (N_21296,N_15749,N_16399);
or U21297 (N_21297,N_17106,N_18503);
and U21298 (N_21298,N_18328,N_16085);
nand U21299 (N_21299,N_17605,N_18610);
or U21300 (N_21300,N_18328,N_16118);
nand U21301 (N_21301,N_17861,N_16664);
nor U21302 (N_21302,N_17214,N_16966);
and U21303 (N_21303,N_18306,N_17166);
or U21304 (N_21304,N_17531,N_16036);
nor U21305 (N_21305,N_15689,N_18016);
and U21306 (N_21306,N_17463,N_18161);
or U21307 (N_21307,N_18110,N_15836);
and U21308 (N_21308,N_16730,N_18744);
nand U21309 (N_21309,N_16205,N_17339);
nor U21310 (N_21310,N_15679,N_15673);
xor U21311 (N_21311,N_15978,N_17333);
xor U21312 (N_21312,N_17457,N_18373);
and U21313 (N_21313,N_17634,N_17868);
nor U21314 (N_21314,N_15665,N_18729);
and U21315 (N_21315,N_18141,N_18740);
nand U21316 (N_21316,N_18524,N_18276);
nor U21317 (N_21317,N_16671,N_15917);
nor U21318 (N_21318,N_16529,N_18504);
nand U21319 (N_21319,N_16536,N_18109);
or U21320 (N_21320,N_18473,N_18377);
and U21321 (N_21321,N_18555,N_17809);
and U21322 (N_21322,N_16526,N_16550);
xor U21323 (N_21323,N_17740,N_17003);
nand U21324 (N_21324,N_17152,N_17269);
or U21325 (N_21325,N_18686,N_18177);
or U21326 (N_21326,N_17819,N_16909);
or U21327 (N_21327,N_15918,N_17604);
nand U21328 (N_21328,N_17834,N_18039);
nand U21329 (N_21329,N_17475,N_18556);
or U21330 (N_21330,N_15703,N_16639);
nand U21331 (N_21331,N_16492,N_15845);
nor U21332 (N_21332,N_16869,N_18552);
or U21333 (N_21333,N_16782,N_16735);
xor U21334 (N_21334,N_17451,N_18290);
or U21335 (N_21335,N_16791,N_16172);
and U21336 (N_21336,N_15783,N_18414);
nand U21337 (N_21337,N_16919,N_17942);
nor U21338 (N_21338,N_17194,N_18324);
nor U21339 (N_21339,N_16924,N_17830);
nand U21340 (N_21340,N_18125,N_16696);
nor U21341 (N_21341,N_17351,N_16421);
or U21342 (N_21342,N_17016,N_18415);
nand U21343 (N_21343,N_18460,N_17656);
nor U21344 (N_21344,N_17065,N_15888);
and U21345 (N_21345,N_15735,N_16400);
nor U21346 (N_21346,N_16801,N_15678);
or U21347 (N_21347,N_17666,N_16665);
and U21348 (N_21348,N_16759,N_16079);
and U21349 (N_21349,N_17245,N_18045);
nor U21350 (N_21350,N_16167,N_15932);
and U21351 (N_21351,N_18200,N_16444);
or U21352 (N_21352,N_17523,N_15980);
and U21353 (N_21353,N_18327,N_17687);
and U21354 (N_21354,N_16805,N_18326);
xnor U21355 (N_21355,N_15904,N_16509);
and U21356 (N_21356,N_18273,N_17078);
and U21357 (N_21357,N_16261,N_17676);
or U21358 (N_21358,N_16604,N_17344);
and U21359 (N_21359,N_17742,N_16758);
nor U21360 (N_21360,N_17426,N_16321);
or U21361 (N_21361,N_18129,N_17368);
and U21362 (N_21362,N_16205,N_17561);
nand U21363 (N_21363,N_17207,N_16883);
nor U21364 (N_21364,N_16705,N_18457);
and U21365 (N_21365,N_16330,N_16335);
nand U21366 (N_21366,N_18223,N_18053);
nand U21367 (N_21367,N_16598,N_16652);
nor U21368 (N_21368,N_16307,N_16102);
and U21369 (N_21369,N_15900,N_16374);
and U21370 (N_21370,N_16097,N_16261);
or U21371 (N_21371,N_17676,N_18238);
and U21372 (N_21372,N_16911,N_16011);
nand U21373 (N_21373,N_18302,N_18040);
xor U21374 (N_21374,N_17043,N_17279);
or U21375 (N_21375,N_18614,N_17768);
nor U21376 (N_21376,N_15918,N_17181);
nor U21377 (N_21377,N_15947,N_18374);
nor U21378 (N_21378,N_15724,N_16061);
nand U21379 (N_21379,N_15988,N_16530);
and U21380 (N_21380,N_17186,N_17361);
or U21381 (N_21381,N_16839,N_17259);
or U21382 (N_21382,N_15759,N_18234);
nand U21383 (N_21383,N_17022,N_17680);
xor U21384 (N_21384,N_18292,N_17857);
nand U21385 (N_21385,N_18206,N_18481);
nand U21386 (N_21386,N_17590,N_15703);
or U21387 (N_21387,N_15937,N_18271);
xor U21388 (N_21388,N_17668,N_17307);
and U21389 (N_21389,N_15856,N_17985);
nor U21390 (N_21390,N_16638,N_15659);
or U21391 (N_21391,N_16762,N_16670);
or U21392 (N_21392,N_16921,N_16049);
nor U21393 (N_21393,N_16801,N_17512);
nand U21394 (N_21394,N_16766,N_16092);
nor U21395 (N_21395,N_18328,N_18408);
nor U21396 (N_21396,N_17903,N_16336);
or U21397 (N_21397,N_16614,N_16104);
nand U21398 (N_21398,N_17660,N_18083);
nand U21399 (N_21399,N_17863,N_15786);
nor U21400 (N_21400,N_17506,N_16501);
nand U21401 (N_21401,N_18569,N_17502);
nor U21402 (N_21402,N_15862,N_17498);
nor U21403 (N_21403,N_16766,N_15635);
or U21404 (N_21404,N_18150,N_17707);
or U21405 (N_21405,N_16655,N_18229);
xnor U21406 (N_21406,N_16286,N_16323);
nor U21407 (N_21407,N_18703,N_16293);
nor U21408 (N_21408,N_18634,N_15662);
and U21409 (N_21409,N_17330,N_16774);
nand U21410 (N_21410,N_18124,N_16855);
nand U21411 (N_21411,N_18021,N_18219);
and U21412 (N_21412,N_17976,N_18428);
and U21413 (N_21413,N_16339,N_18390);
nor U21414 (N_21414,N_18401,N_17130);
or U21415 (N_21415,N_18708,N_18117);
and U21416 (N_21416,N_17582,N_15869);
nand U21417 (N_21417,N_18487,N_18576);
or U21418 (N_21418,N_18284,N_16405);
or U21419 (N_21419,N_16741,N_17398);
xnor U21420 (N_21420,N_16505,N_17865);
nor U21421 (N_21421,N_17110,N_16701);
or U21422 (N_21422,N_16503,N_17644);
and U21423 (N_21423,N_17859,N_16252);
nand U21424 (N_21424,N_18475,N_18366);
nand U21425 (N_21425,N_16324,N_16899);
or U21426 (N_21426,N_18576,N_18089);
or U21427 (N_21427,N_18467,N_17957);
xnor U21428 (N_21428,N_16037,N_16485);
or U21429 (N_21429,N_16958,N_17010);
nand U21430 (N_21430,N_18216,N_18489);
or U21431 (N_21431,N_17958,N_16262);
nor U21432 (N_21432,N_17825,N_18679);
and U21433 (N_21433,N_18632,N_17493);
or U21434 (N_21434,N_17253,N_17885);
nor U21435 (N_21435,N_16504,N_17480);
nand U21436 (N_21436,N_16080,N_17446);
and U21437 (N_21437,N_16552,N_16801);
xnor U21438 (N_21438,N_17467,N_18057);
and U21439 (N_21439,N_17775,N_17923);
and U21440 (N_21440,N_18020,N_18135);
and U21441 (N_21441,N_17655,N_18385);
nor U21442 (N_21442,N_15636,N_18171);
nor U21443 (N_21443,N_17646,N_16362);
nand U21444 (N_21444,N_16419,N_16282);
nor U21445 (N_21445,N_17656,N_16976);
xnor U21446 (N_21446,N_16590,N_15988);
and U21447 (N_21447,N_16057,N_16764);
nor U21448 (N_21448,N_17232,N_17214);
nor U21449 (N_21449,N_16519,N_18206);
or U21450 (N_21450,N_16814,N_18690);
nor U21451 (N_21451,N_17733,N_16287);
or U21452 (N_21452,N_16530,N_17363);
nand U21453 (N_21453,N_18390,N_16287);
and U21454 (N_21454,N_18143,N_16747);
nand U21455 (N_21455,N_17956,N_16295);
and U21456 (N_21456,N_16686,N_16047);
and U21457 (N_21457,N_17431,N_17461);
and U21458 (N_21458,N_16526,N_16379);
nand U21459 (N_21459,N_16864,N_18308);
nor U21460 (N_21460,N_15752,N_16038);
nor U21461 (N_21461,N_17108,N_18670);
nand U21462 (N_21462,N_17978,N_18142);
xnor U21463 (N_21463,N_17721,N_18176);
and U21464 (N_21464,N_17750,N_15943);
or U21465 (N_21465,N_18513,N_17694);
or U21466 (N_21466,N_17428,N_17201);
nand U21467 (N_21467,N_15628,N_15785);
and U21468 (N_21468,N_16114,N_15851);
xor U21469 (N_21469,N_17596,N_17431);
or U21470 (N_21470,N_18595,N_18706);
and U21471 (N_21471,N_15892,N_15941);
and U21472 (N_21472,N_18715,N_15923);
and U21473 (N_21473,N_18024,N_16204);
or U21474 (N_21474,N_17655,N_17915);
nor U21475 (N_21475,N_16564,N_15890);
nand U21476 (N_21476,N_17184,N_18653);
and U21477 (N_21477,N_18458,N_15754);
nor U21478 (N_21478,N_17940,N_16723);
and U21479 (N_21479,N_18111,N_17963);
and U21480 (N_21480,N_16235,N_18022);
and U21481 (N_21481,N_16098,N_17581);
xnor U21482 (N_21482,N_15850,N_15951);
xor U21483 (N_21483,N_16319,N_16130);
nor U21484 (N_21484,N_17402,N_17416);
or U21485 (N_21485,N_17890,N_16941);
or U21486 (N_21486,N_15850,N_15925);
nor U21487 (N_21487,N_15983,N_16925);
nand U21488 (N_21488,N_16221,N_16831);
xnor U21489 (N_21489,N_18157,N_16769);
nand U21490 (N_21490,N_16997,N_18539);
or U21491 (N_21491,N_18231,N_15848);
nor U21492 (N_21492,N_16381,N_18649);
nand U21493 (N_21493,N_16113,N_16213);
or U21494 (N_21494,N_17632,N_15993);
nor U21495 (N_21495,N_18543,N_18482);
or U21496 (N_21496,N_15857,N_16472);
nand U21497 (N_21497,N_15781,N_16329);
nor U21498 (N_21498,N_16425,N_17690);
nand U21499 (N_21499,N_17579,N_17166);
and U21500 (N_21500,N_16257,N_16935);
or U21501 (N_21501,N_18731,N_18225);
nor U21502 (N_21502,N_16785,N_17235);
or U21503 (N_21503,N_18211,N_16159);
and U21504 (N_21504,N_16401,N_15869);
nor U21505 (N_21505,N_17653,N_17744);
and U21506 (N_21506,N_18675,N_16930);
and U21507 (N_21507,N_15810,N_17336);
or U21508 (N_21508,N_18152,N_16463);
or U21509 (N_21509,N_17301,N_17705);
and U21510 (N_21510,N_18576,N_16612);
or U21511 (N_21511,N_17439,N_17500);
nand U21512 (N_21512,N_17082,N_16556);
nor U21513 (N_21513,N_17094,N_16046);
or U21514 (N_21514,N_17477,N_15799);
nand U21515 (N_21515,N_16160,N_18693);
or U21516 (N_21516,N_16298,N_17237);
nor U21517 (N_21517,N_18111,N_17512);
and U21518 (N_21518,N_17690,N_16086);
nor U21519 (N_21519,N_18531,N_18498);
nand U21520 (N_21520,N_15958,N_18015);
or U21521 (N_21521,N_17492,N_17517);
xnor U21522 (N_21522,N_16453,N_18728);
nor U21523 (N_21523,N_16615,N_16406);
xnor U21524 (N_21524,N_15638,N_18032);
or U21525 (N_21525,N_18245,N_17463);
xor U21526 (N_21526,N_17320,N_17205);
or U21527 (N_21527,N_16168,N_18394);
and U21528 (N_21528,N_16172,N_16983);
nand U21529 (N_21529,N_16037,N_18639);
and U21530 (N_21530,N_18369,N_17613);
and U21531 (N_21531,N_17426,N_15983);
or U21532 (N_21532,N_18076,N_16160);
nor U21533 (N_21533,N_18401,N_17182);
xnor U21534 (N_21534,N_17808,N_17661);
and U21535 (N_21535,N_15687,N_16427);
nand U21536 (N_21536,N_17874,N_17168);
or U21537 (N_21537,N_17623,N_17768);
nor U21538 (N_21538,N_16525,N_17154);
nand U21539 (N_21539,N_17596,N_16567);
or U21540 (N_21540,N_16662,N_17599);
nand U21541 (N_21541,N_17584,N_18589);
or U21542 (N_21542,N_17092,N_17271);
or U21543 (N_21543,N_17591,N_16452);
and U21544 (N_21544,N_15790,N_16275);
and U21545 (N_21545,N_17660,N_18422);
nand U21546 (N_21546,N_16865,N_16237);
and U21547 (N_21547,N_15762,N_16113);
and U21548 (N_21548,N_17124,N_17399);
nor U21549 (N_21549,N_18362,N_18503);
nand U21550 (N_21550,N_18602,N_16789);
or U21551 (N_21551,N_16066,N_17348);
nor U21552 (N_21552,N_15800,N_16457);
nor U21553 (N_21553,N_17892,N_16277);
or U21554 (N_21554,N_18072,N_17380);
nor U21555 (N_21555,N_18314,N_18576);
nor U21556 (N_21556,N_16077,N_15927);
nand U21557 (N_21557,N_15968,N_18580);
and U21558 (N_21558,N_16330,N_17691);
and U21559 (N_21559,N_17493,N_17562);
and U21560 (N_21560,N_17761,N_18307);
nor U21561 (N_21561,N_17704,N_17005);
xnor U21562 (N_21562,N_16125,N_18171);
nand U21563 (N_21563,N_16805,N_16331);
nor U21564 (N_21564,N_17131,N_17297);
and U21565 (N_21565,N_18335,N_15937);
nand U21566 (N_21566,N_16027,N_16861);
nor U21567 (N_21567,N_17316,N_16685);
nor U21568 (N_21568,N_18423,N_15661);
and U21569 (N_21569,N_15747,N_16316);
nor U21570 (N_21570,N_17834,N_17375);
nand U21571 (N_21571,N_18355,N_17714);
or U21572 (N_21572,N_18121,N_16798);
nand U21573 (N_21573,N_16117,N_16517);
and U21574 (N_21574,N_17005,N_16942);
nand U21575 (N_21575,N_15987,N_15940);
nand U21576 (N_21576,N_17860,N_15793);
nand U21577 (N_21577,N_17156,N_18022);
xor U21578 (N_21578,N_18092,N_15657);
nor U21579 (N_21579,N_15921,N_16026);
nor U21580 (N_21580,N_16896,N_17535);
or U21581 (N_21581,N_16498,N_18331);
or U21582 (N_21582,N_16343,N_16948);
or U21583 (N_21583,N_17905,N_17005);
xnor U21584 (N_21584,N_16004,N_16760);
nor U21585 (N_21585,N_17092,N_16651);
nor U21586 (N_21586,N_17989,N_18116);
or U21587 (N_21587,N_15868,N_16898);
and U21588 (N_21588,N_16656,N_17599);
nor U21589 (N_21589,N_18713,N_16774);
nor U21590 (N_21590,N_18284,N_16251);
nand U21591 (N_21591,N_18256,N_16162);
nand U21592 (N_21592,N_16634,N_17892);
and U21593 (N_21593,N_17328,N_15878);
nand U21594 (N_21594,N_17329,N_17386);
and U21595 (N_21595,N_18200,N_17896);
or U21596 (N_21596,N_17562,N_18464);
nand U21597 (N_21597,N_16230,N_18473);
or U21598 (N_21598,N_17680,N_17332);
nor U21599 (N_21599,N_18264,N_18229);
and U21600 (N_21600,N_17897,N_16900);
or U21601 (N_21601,N_18734,N_18248);
or U21602 (N_21602,N_18494,N_18375);
and U21603 (N_21603,N_18695,N_17196);
nand U21604 (N_21604,N_17511,N_15860);
and U21605 (N_21605,N_18531,N_18659);
nor U21606 (N_21606,N_16575,N_16201);
and U21607 (N_21607,N_18373,N_18547);
nand U21608 (N_21608,N_15911,N_16537);
nor U21609 (N_21609,N_18132,N_15737);
and U21610 (N_21610,N_18595,N_15910);
and U21611 (N_21611,N_17870,N_16419);
and U21612 (N_21612,N_17254,N_16877);
nand U21613 (N_21613,N_17772,N_17019);
nor U21614 (N_21614,N_15770,N_17867);
or U21615 (N_21615,N_16754,N_18273);
or U21616 (N_21616,N_17209,N_15857);
nor U21617 (N_21617,N_17849,N_18625);
and U21618 (N_21618,N_16107,N_16995);
and U21619 (N_21619,N_16035,N_16529);
or U21620 (N_21620,N_18586,N_17316);
xnor U21621 (N_21621,N_18192,N_17458);
and U21622 (N_21622,N_16332,N_16022);
nand U21623 (N_21623,N_17966,N_18412);
and U21624 (N_21624,N_16124,N_16250);
and U21625 (N_21625,N_18345,N_16129);
nand U21626 (N_21626,N_15716,N_18649);
nand U21627 (N_21627,N_17849,N_18557);
and U21628 (N_21628,N_16157,N_18569);
nor U21629 (N_21629,N_15939,N_17006);
nor U21630 (N_21630,N_17860,N_17154);
and U21631 (N_21631,N_16490,N_16994);
nor U21632 (N_21632,N_16137,N_17658);
nor U21633 (N_21633,N_16258,N_17326);
xnor U21634 (N_21634,N_15847,N_18063);
and U21635 (N_21635,N_17351,N_17852);
nand U21636 (N_21636,N_17432,N_17328);
and U21637 (N_21637,N_18208,N_17710);
xor U21638 (N_21638,N_16201,N_17859);
nand U21639 (N_21639,N_17033,N_18408);
and U21640 (N_21640,N_16978,N_17885);
and U21641 (N_21641,N_17702,N_15915);
and U21642 (N_21642,N_17842,N_18683);
nand U21643 (N_21643,N_18707,N_18114);
and U21644 (N_21644,N_16035,N_17580);
and U21645 (N_21645,N_16800,N_16544);
and U21646 (N_21646,N_16909,N_15765);
nand U21647 (N_21647,N_18258,N_18251);
nand U21648 (N_21648,N_16028,N_18005);
and U21649 (N_21649,N_18092,N_16497);
nor U21650 (N_21650,N_17917,N_17070);
nor U21651 (N_21651,N_16168,N_17500);
and U21652 (N_21652,N_16020,N_17049);
or U21653 (N_21653,N_16488,N_18140);
and U21654 (N_21654,N_15964,N_17877);
nor U21655 (N_21655,N_18612,N_16411);
nor U21656 (N_21656,N_17443,N_18340);
nand U21657 (N_21657,N_18085,N_17386);
and U21658 (N_21658,N_15915,N_17509);
and U21659 (N_21659,N_18436,N_17932);
nand U21660 (N_21660,N_15741,N_15798);
or U21661 (N_21661,N_16218,N_16036);
and U21662 (N_21662,N_18674,N_16417);
and U21663 (N_21663,N_16356,N_18051);
nand U21664 (N_21664,N_17256,N_16782);
xnor U21665 (N_21665,N_16737,N_17555);
nand U21666 (N_21666,N_17993,N_16853);
nor U21667 (N_21667,N_17813,N_15924);
nand U21668 (N_21668,N_18626,N_17452);
nand U21669 (N_21669,N_17915,N_15727);
nand U21670 (N_21670,N_17544,N_17604);
nor U21671 (N_21671,N_16247,N_17256);
or U21672 (N_21672,N_18699,N_16844);
nand U21673 (N_21673,N_15932,N_17688);
nor U21674 (N_21674,N_17521,N_16868);
and U21675 (N_21675,N_18560,N_18523);
and U21676 (N_21676,N_17213,N_15816);
or U21677 (N_21677,N_16790,N_18538);
nor U21678 (N_21678,N_18509,N_17389);
nor U21679 (N_21679,N_15991,N_18618);
nand U21680 (N_21680,N_15869,N_16141);
nor U21681 (N_21681,N_18729,N_17932);
or U21682 (N_21682,N_15961,N_17387);
nor U21683 (N_21683,N_16397,N_17710);
or U21684 (N_21684,N_16505,N_18665);
or U21685 (N_21685,N_16270,N_16315);
nor U21686 (N_21686,N_15769,N_18315);
or U21687 (N_21687,N_15844,N_18245);
xor U21688 (N_21688,N_17984,N_18357);
or U21689 (N_21689,N_15918,N_16158);
nor U21690 (N_21690,N_17549,N_17713);
nand U21691 (N_21691,N_18538,N_16234);
and U21692 (N_21692,N_15752,N_17507);
and U21693 (N_21693,N_18163,N_16829);
xnor U21694 (N_21694,N_16850,N_17138);
nand U21695 (N_21695,N_16580,N_15934);
or U21696 (N_21696,N_18210,N_16790);
or U21697 (N_21697,N_18288,N_18690);
and U21698 (N_21698,N_17055,N_17572);
nor U21699 (N_21699,N_17053,N_16369);
or U21700 (N_21700,N_16681,N_18222);
xor U21701 (N_21701,N_18714,N_17831);
nand U21702 (N_21702,N_17212,N_16687);
and U21703 (N_21703,N_17659,N_16251);
xor U21704 (N_21704,N_16797,N_15749);
or U21705 (N_21705,N_16937,N_17039);
nor U21706 (N_21706,N_16852,N_16809);
and U21707 (N_21707,N_15976,N_15866);
and U21708 (N_21708,N_18732,N_17780);
nor U21709 (N_21709,N_16184,N_16843);
nor U21710 (N_21710,N_18243,N_18013);
nor U21711 (N_21711,N_16059,N_18370);
nor U21712 (N_21712,N_17580,N_16433);
nor U21713 (N_21713,N_15734,N_17631);
xnor U21714 (N_21714,N_16566,N_17134);
nor U21715 (N_21715,N_17275,N_17220);
and U21716 (N_21716,N_16602,N_17962);
and U21717 (N_21717,N_16782,N_17241);
or U21718 (N_21718,N_17958,N_15723);
or U21719 (N_21719,N_17952,N_18467);
or U21720 (N_21720,N_17741,N_16274);
nand U21721 (N_21721,N_15950,N_16692);
nor U21722 (N_21722,N_18432,N_18138);
or U21723 (N_21723,N_16984,N_18704);
and U21724 (N_21724,N_17349,N_17969);
nor U21725 (N_21725,N_17590,N_15871);
and U21726 (N_21726,N_18151,N_16010);
nand U21727 (N_21727,N_17020,N_18279);
or U21728 (N_21728,N_17521,N_15703);
xor U21729 (N_21729,N_18699,N_16469);
and U21730 (N_21730,N_18158,N_18630);
or U21731 (N_21731,N_15792,N_17664);
xor U21732 (N_21732,N_16757,N_18369);
xor U21733 (N_21733,N_18176,N_18371);
and U21734 (N_21734,N_17916,N_17001);
nor U21735 (N_21735,N_17862,N_17614);
or U21736 (N_21736,N_18003,N_16703);
xnor U21737 (N_21737,N_16900,N_15678);
and U21738 (N_21738,N_18514,N_17805);
or U21739 (N_21739,N_17658,N_17342);
nand U21740 (N_21740,N_16447,N_16588);
and U21741 (N_21741,N_17323,N_17063);
and U21742 (N_21742,N_17523,N_16761);
and U21743 (N_21743,N_15783,N_18362);
and U21744 (N_21744,N_16028,N_18003);
xnor U21745 (N_21745,N_16314,N_16473);
xnor U21746 (N_21746,N_17915,N_16475);
nand U21747 (N_21747,N_16062,N_17606);
nand U21748 (N_21748,N_18515,N_17865);
xnor U21749 (N_21749,N_16076,N_18729);
or U21750 (N_21750,N_16841,N_15865);
nand U21751 (N_21751,N_16028,N_17727);
nand U21752 (N_21752,N_17479,N_17749);
nor U21753 (N_21753,N_15814,N_17430);
nor U21754 (N_21754,N_17139,N_18164);
nand U21755 (N_21755,N_16065,N_17075);
or U21756 (N_21756,N_17040,N_17896);
or U21757 (N_21757,N_17375,N_17582);
nor U21758 (N_21758,N_15857,N_16564);
xnor U21759 (N_21759,N_16732,N_16426);
or U21760 (N_21760,N_16263,N_18503);
or U21761 (N_21761,N_18628,N_16694);
xor U21762 (N_21762,N_17845,N_16008);
and U21763 (N_21763,N_18007,N_18146);
nor U21764 (N_21764,N_16465,N_17874);
and U21765 (N_21765,N_16476,N_17261);
or U21766 (N_21766,N_15946,N_17658);
or U21767 (N_21767,N_15859,N_17095);
nand U21768 (N_21768,N_17208,N_17947);
xor U21769 (N_21769,N_18290,N_18743);
and U21770 (N_21770,N_17318,N_17935);
nand U21771 (N_21771,N_18262,N_16252);
nor U21772 (N_21772,N_18409,N_16497);
or U21773 (N_21773,N_16258,N_18336);
nand U21774 (N_21774,N_16467,N_18726);
nand U21775 (N_21775,N_17667,N_18143);
and U21776 (N_21776,N_16555,N_17586);
and U21777 (N_21777,N_16264,N_17116);
or U21778 (N_21778,N_17074,N_17590);
or U21779 (N_21779,N_18208,N_18481);
and U21780 (N_21780,N_15744,N_15739);
nand U21781 (N_21781,N_18705,N_18247);
nor U21782 (N_21782,N_18226,N_17579);
and U21783 (N_21783,N_17661,N_17507);
and U21784 (N_21784,N_18323,N_17988);
and U21785 (N_21785,N_16874,N_16071);
xor U21786 (N_21786,N_16538,N_16445);
or U21787 (N_21787,N_18344,N_15627);
nor U21788 (N_21788,N_18481,N_15650);
nor U21789 (N_21789,N_18675,N_16682);
or U21790 (N_21790,N_16934,N_17683);
nand U21791 (N_21791,N_16246,N_17933);
nand U21792 (N_21792,N_16474,N_17785);
xor U21793 (N_21793,N_17944,N_16775);
nand U21794 (N_21794,N_16360,N_15906);
nand U21795 (N_21795,N_17244,N_17120);
nand U21796 (N_21796,N_16252,N_15737);
xnor U21797 (N_21797,N_17969,N_17904);
nand U21798 (N_21798,N_16481,N_16515);
or U21799 (N_21799,N_17589,N_18664);
or U21800 (N_21800,N_17737,N_16420);
nor U21801 (N_21801,N_15661,N_15650);
nor U21802 (N_21802,N_17718,N_15744);
nor U21803 (N_21803,N_18598,N_17141);
or U21804 (N_21804,N_18257,N_18714);
nor U21805 (N_21805,N_17332,N_17099);
nand U21806 (N_21806,N_17577,N_17058);
and U21807 (N_21807,N_18162,N_18665);
nand U21808 (N_21808,N_18066,N_16430);
or U21809 (N_21809,N_15899,N_18506);
and U21810 (N_21810,N_16500,N_18175);
or U21811 (N_21811,N_16887,N_18431);
nor U21812 (N_21812,N_16278,N_16251);
or U21813 (N_21813,N_17686,N_16493);
and U21814 (N_21814,N_18082,N_16113);
nor U21815 (N_21815,N_18235,N_17402);
nand U21816 (N_21816,N_18199,N_17981);
nor U21817 (N_21817,N_18664,N_17863);
nand U21818 (N_21818,N_17903,N_18595);
and U21819 (N_21819,N_16884,N_17222);
nor U21820 (N_21820,N_17524,N_16852);
nand U21821 (N_21821,N_16490,N_18253);
and U21822 (N_21822,N_17972,N_17358);
nand U21823 (N_21823,N_17686,N_16270);
nor U21824 (N_21824,N_16432,N_15711);
and U21825 (N_21825,N_16078,N_16262);
and U21826 (N_21826,N_15935,N_16907);
or U21827 (N_21827,N_18537,N_16813);
nor U21828 (N_21828,N_17595,N_16395);
or U21829 (N_21829,N_17634,N_17025);
and U21830 (N_21830,N_17707,N_17782);
or U21831 (N_21831,N_16768,N_16199);
nand U21832 (N_21832,N_17547,N_16823);
and U21833 (N_21833,N_18399,N_17197);
and U21834 (N_21834,N_16866,N_16259);
nor U21835 (N_21835,N_15630,N_18162);
nand U21836 (N_21836,N_18603,N_18356);
or U21837 (N_21837,N_17403,N_16300);
and U21838 (N_21838,N_18173,N_17375);
and U21839 (N_21839,N_18196,N_17666);
and U21840 (N_21840,N_16422,N_18485);
or U21841 (N_21841,N_17369,N_18736);
and U21842 (N_21842,N_17191,N_16057);
or U21843 (N_21843,N_16148,N_17930);
and U21844 (N_21844,N_16644,N_18482);
nor U21845 (N_21845,N_16294,N_16956);
nand U21846 (N_21846,N_16835,N_17364);
or U21847 (N_21847,N_17297,N_16825);
nand U21848 (N_21848,N_16785,N_15789);
or U21849 (N_21849,N_18438,N_17244);
xnor U21850 (N_21850,N_16583,N_18604);
nor U21851 (N_21851,N_16002,N_17294);
nand U21852 (N_21852,N_15996,N_16425);
nand U21853 (N_21853,N_17973,N_18100);
or U21854 (N_21854,N_16664,N_17877);
nor U21855 (N_21855,N_17240,N_17397);
nand U21856 (N_21856,N_15850,N_16086);
nor U21857 (N_21857,N_15650,N_17661);
or U21858 (N_21858,N_15930,N_16054);
or U21859 (N_21859,N_16995,N_17656);
xnor U21860 (N_21860,N_16078,N_16402);
and U21861 (N_21861,N_16525,N_15634);
nor U21862 (N_21862,N_17036,N_16406);
nand U21863 (N_21863,N_17205,N_16680);
nand U21864 (N_21864,N_16035,N_18045);
and U21865 (N_21865,N_17669,N_18704);
nand U21866 (N_21866,N_16640,N_16578);
nand U21867 (N_21867,N_17173,N_18553);
and U21868 (N_21868,N_17949,N_15708);
xor U21869 (N_21869,N_15849,N_17701);
nor U21870 (N_21870,N_16133,N_18520);
or U21871 (N_21871,N_18704,N_16560);
nand U21872 (N_21872,N_17707,N_16371);
or U21873 (N_21873,N_18367,N_16729);
or U21874 (N_21874,N_16364,N_17068);
or U21875 (N_21875,N_19335,N_18813);
nand U21876 (N_21876,N_19741,N_21563);
nand U21877 (N_21877,N_18773,N_21735);
nor U21878 (N_21878,N_20014,N_20065);
nor U21879 (N_21879,N_19547,N_19431);
xor U21880 (N_21880,N_20497,N_20339);
or U21881 (N_21881,N_21360,N_21095);
xnor U21882 (N_21882,N_19743,N_19871);
and U21883 (N_21883,N_21315,N_20624);
xor U21884 (N_21884,N_20763,N_20131);
and U21885 (N_21885,N_21460,N_19237);
nor U21886 (N_21886,N_20224,N_20464);
or U21887 (N_21887,N_20778,N_19200);
and U21888 (N_21888,N_19816,N_20284);
or U21889 (N_21889,N_19725,N_20445);
nand U21890 (N_21890,N_21854,N_21545);
and U21891 (N_21891,N_19705,N_21367);
xnor U21892 (N_21892,N_21321,N_18764);
or U21893 (N_21893,N_20851,N_20407);
nor U21894 (N_21894,N_20831,N_20936);
nor U21895 (N_21895,N_20958,N_19793);
nor U21896 (N_21896,N_20174,N_21217);
xnor U21897 (N_21897,N_20058,N_20678);
and U21898 (N_21898,N_19569,N_19825);
nor U21899 (N_21899,N_21813,N_21323);
nand U21900 (N_21900,N_20708,N_21422);
nor U21901 (N_21901,N_20033,N_21814);
or U21902 (N_21902,N_21757,N_18783);
and U21903 (N_21903,N_18986,N_19722);
nor U21904 (N_21904,N_21288,N_20453);
or U21905 (N_21905,N_19154,N_19105);
xor U21906 (N_21906,N_20069,N_19817);
and U21907 (N_21907,N_21615,N_19144);
and U21908 (N_21908,N_21358,N_19690);
nor U21909 (N_21909,N_18852,N_19985);
or U21910 (N_21910,N_20122,N_21281);
and U21911 (N_21911,N_19808,N_19076);
nand U21912 (N_21912,N_20452,N_20773);
or U21913 (N_21913,N_18921,N_19776);
and U21914 (N_21914,N_19242,N_20027);
and U21915 (N_21915,N_19671,N_20351);
nand U21916 (N_21916,N_20682,N_21684);
or U21917 (N_21917,N_20366,N_19266);
and U21918 (N_21918,N_19914,N_20162);
xor U21919 (N_21919,N_20946,N_20079);
nor U21920 (N_21920,N_21830,N_21825);
nand U21921 (N_21921,N_21183,N_19605);
nor U21922 (N_21922,N_19185,N_20455);
xor U21923 (N_21923,N_21478,N_20603);
nor U21924 (N_21924,N_20051,N_21595);
nand U21925 (N_21925,N_20769,N_21754);
nand U21926 (N_21926,N_19410,N_19572);
and U21927 (N_21927,N_21463,N_20211);
nor U21928 (N_21928,N_20276,N_18928);
and U21929 (N_21929,N_20722,N_20903);
and U21930 (N_21930,N_19901,N_21466);
or U21931 (N_21931,N_18846,N_19870);
or U21932 (N_21932,N_19933,N_21429);
xor U21933 (N_21933,N_19460,N_19486);
and U21934 (N_21934,N_20371,N_20290);
and U21935 (N_21935,N_19481,N_19639);
nand U21936 (N_21936,N_19786,N_20743);
and U21937 (N_21937,N_21715,N_20871);
and U21938 (N_21938,N_21448,N_21574);
nand U21939 (N_21939,N_20706,N_19523);
and U21940 (N_21940,N_21761,N_19413);
nor U21941 (N_21941,N_20039,N_19094);
and U21942 (N_21942,N_19361,N_20578);
nand U21943 (N_21943,N_21285,N_19804);
nor U21944 (N_21944,N_19762,N_21052);
nor U21945 (N_21945,N_20654,N_20320);
and U21946 (N_21946,N_21704,N_19658);
nand U21947 (N_21947,N_20523,N_19283);
xnor U21948 (N_21948,N_19442,N_20103);
nor U21949 (N_21949,N_20471,N_20726);
and U21950 (N_21950,N_21257,N_20280);
nor U21951 (N_21951,N_18835,N_20228);
nand U21952 (N_21952,N_19814,N_20525);
nand U21953 (N_21953,N_21708,N_20089);
nor U21954 (N_21954,N_20856,N_19982);
nand U21955 (N_21955,N_19840,N_21197);
xnor U21956 (N_21956,N_20929,N_19192);
or U21957 (N_21957,N_19432,N_18924);
nand U21958 (N_21958,N_19924,N_20244);
xnor U21959 (N_21959,N_19554,N_20776);
and U21960 (N_21960,N_20943,N_20234);
xnor U21961 (N_21961,N_21393,N_21407);
nand U21962 (N_21962,N_18810,N_20101);
nand U21963 (N_21963,N_20202,N_21071);
or U21964 (N_21964,N_20976,N_20710);
or U21965 (N_21965,N_19541,N_19699);
nor U21966 (N_21966,N_18858,N_21439);
nand U21967 (N_21967,N_19249,N_21192);
and U21968 (N_21968,N_19909,N_20006);
xnor U21969 (N_21969,N_21032,N_18757);
and U21970 (N_21970,N_21055,N_20309);
and U21971 (N_21971,N_20792,N_20558);
xor U21972 (N_21972,N_19204,N_19519);
xnor U21973 (N_21973,N_21173,N_19517);
and U21974 (N_21974,N_19995,N_21792);
and U21975 (N_21975,N_19222,N_20233);
nor U21976 (N_21976,N_21536,N_20590);
nor U21977 (N_21977,N_21331,N_20466);
nor U21978 (N_21978,N_20119,N_19856);
or U21979 (N_21979,N_21234,N_21420);
or U21980 (N_21980,N_19300,N_20826);
or U21981 (N_21981,N_19221,N_21230);
and U21982 (N_21982,N_19846,N_20697);
and U21983 (N_21983,N_21620,N_21293);
nand U21984 (N_21984,N_21001,N_19451);
nand U21985 (N_21985,N_19411,N_21289);
and U21986 (N_21986,N_18899,N_21558);
nor U21987 (N_21987,N_21828,N_18784);
nor U21988 (N_21988,N_21568,N_19838);
nor U21989 (N_21989,N_21622,N_20198);
nand U21990 (N_21990,N_19594,N_19456);
nand U21991 (N_21991,N_20696,N_20306);
and U21992 (N_21992,N_18867,N_20670);
xnor U21993 (N_21993,N_20388,N_20510);
nor U21994 (N_21994,N_19683,N_20095);
or U21995 (N_21995,N_19157,N_21324);
nor U21996 (N_21996,N_20744,N_21572);
or U21997 (N_21997,N_21824,N_20865);
and U21998 (N_21998,N_19966,N_21273);
nand U21999 (N_21999,N_19674,N_21734);
nor U22000 (N_22000,N_19781,N_20611);
nor U22001 (N_22001,N_19219,N_21397);
and U22002 (N_22002,N_18808,N_19708);
nor U22003 (N_22003,N_19498,N_21566);
nand U22004 (N_22004,N_18789,N_19503);
or U22005 (N_22005,N_19224,N_19977);
and U22006 (N_22006,N_20379,N_21596);
nor U22007 (N_22007,N_21798,N_21077);
and U22008 (N_22008,N_21581,N_19390);
nand U22009 (N_22009,N_19796,N_21712);
nor U22010 (N_22010,N_20334,N_21274);
nor U22011 (N_22011,N_21379,N_19975);
nand U22012 (N_22012,N_21800,N_18972);
nor U22013 (N_22013,N_20934,N_21503);
nand U22014 (N_22014,N_19152,N_18929);
nor U22015 (N_22015,N_19060,N_19891);
and U22016 (N_22016,N_19533,N_19401);
nand U22017 (N_22017,N_19007,N_19499);
and U22018 (N_22018,N_20702,N_19593);
xor U22019 (N_22019,N_19120,N_20256);
or U22020 (N_22020,N_21441,N_21416);
nand U22021 (N_22021,N_21056,N_21258);
and U22022 (N_22022,N_21635,N_21510);
nand U22023 (N_22023,N_20362,N_20998);
or U22024 (N_22024,N_19961,N_19435);
nand U22025 (N_22025,N_21755,N_21455);
nor U22026 (N_22026,N_21205,N_20272);
and U22027 (N_22027,N_19555,N_19339);
xor U22028 (N_22028,N_20022,N_20960);
nand U22029 (N_22029,N_20567,N_20389);
or U22030 (N_22030,N_21191,N_20410);
or U22031 (N_22031,N_21085,N_19761);
and U22032 (N_22032,N_20004,N_18876);
and U22033 (N_22033,N_21041,N_20532);
nor U22034 (N_22034,N_21580,N_21674);
xnor U22035 (N_22035,N_20031,N_20323);
nand U22036 (N_22036,N_21725,N_20994);
nor U22037 (N_22037,N_21599,N_21625);
xor U22038 (N_22038,N_20528,N_21264);
nor U22039 (N_22039,N_21256,N_18787);
xnor U22040 (N_22040,N_21844,N_21556);
and U22041 (N_22041,N_20250,N_19057);
xor U22042 (N_22042,N_20199,N_19052);
or U22043 (N_22043,N_20693,N_20335);
and U22044 (N_22044,N_18973,N_18957);
and U22045 (N_22045,N_21294,N_21352);
and U22046 (N_22046,N_19617,N_19501);
nor U22047 (N_22047,N_21817,N_21683);
nor U22048 (N_22048,N_19385,N_19272);
or U22049 (N_22049,N_21202,N_21243);
nor U22050 (N_22050,N_20349,N_21035);
nor U22051 (N_22051,N_20206,N_20788);
and U22052 (N_22052,N_19061,N_18829);
and U22053 (N_22053,N_20917,N_21337);
or U22054 (N_22054,N_20660,N_21790);
and U22055 (N_22055,N_18934,N_19245);
nor U22056 (N_22056,N_19780,N_20922);
xnor U22057 (N_22057,N_20341,N_20952);
or U22058 (N_22058,N_21851,N_21014);
xnor U22059 (N_22059,N_20220,N_21210);
and U22060 (N_22060,N_20164,N_18913);
nand U22061 (N_22061,N_19608,N_19999);
nor U22062 (N_22062,N_19751,N_21401);
or U22063 (N_22063,N_19552,N_21030);
or U22064 (N_22064,N_21768,N_19243);
nand U22065 (N_22065,N_19186,N_21451);
and U22066 (N_22066,N_21506,N_20397);
and U22067 (N_22067,N_20935,N_18833);
and U22068 (N_22068,N_19679,N_20519);
nor U22069 (N_22069,N_20003,N_21189);
nand U22070 (N_22070,N_20085,N_20391);
nand U22071 (N_22071,N_20905,N_21370);
nand U22072 (N_22072,N_19710,N_20138);
or U22073 (N_22073,N_21349,N_19673);
nand U22074 (N_22074,N_21396,N_18756);
nand U22075 (N_22075,N_19175,N_20026);
nand U22076 (N_22076,N_20919,N_20880);
or U22077 (N_22077,N_20734,N_18998);
or U22078 (N_22078,N_20633,N_20277);
nor U22079 (N_22079,N_20313,N_21547);
or U22080 (N_22080,N_19469,N_19286);
or U22081 (N_22081,N_20091,N_20945);
or U22082 (N_22082,N_21533,N_21414);
or U22083 (N_22083,N_19281,N_20368);
or U22084 (N_22084,N_19349,N_21729);
and U22085 (N_22085,N_20983,N_20414);
nor U22086 (N_22086,N_20484,N_21665);
and U22087 (N_22087,N_19027,N_20154);
or U22088 (N_22088,N_21485,N_20714);
and U22089 (N_22089,N_21618,N_19691);
or U22090 (N_22090,N_19806,N_21312);
and U22091 (N_22091,N_19675,N_21788);
xor U22092 (N_22092,N_21650,N_21594);
nor U22093 (N_22093,N_18926,N_19306);
and U22094 (N_22094,N_19903,N_21124);
nor U22095 (N_22095,N_21314,N_20017);
xor U22096 (N_22096,N_20582,N_21526);
nand U22097 (N_22097,N_19884,N_19827);
xor U22098 (N_22098,N_21659,N_21562);
nand U22099 (N_22099,N_19034,N_20894);
xor U22100 (N_22100,N_18753,N_20166);
and U22101 (N_22101,N_20443,N_21190);
or U22102 (N_22102,N_18982,N_19942);
and U22103 (N_22103,N_20949,N_19558);
nand U22104 (N_22104,N_21653,N_21473);
or U22105 (N_22105,N_20648,N_20915);
and U22106 (N_22106,N_21789,N_20802);
nor U22107 (N_22107,N_20360,N_19275);
and U22108 (N_22108,N_19146,N_21428);
nor U22109 (N_22109,N_21421,N_19527);
and U22110 (N_22110,N_20193,N_20786);
or U22111 (N_22111,N_21573,N_21706);
nor U22112 (N_22112,N_20757,N_19201);
nand U22113 (N_22113,N_19291,N_19086);
and U22114 (N_22114,N_19858,N_21647);
nor U22115 (N_22115,N_20900,N_20442);
or U22116 (N_22116,N_20692,N_21468);
or U22117 (N_22117,N_20892,N_19434);
and U22118 (N_22118,N_21799,N_21797);
or U22119 (N_22119,N_20562,N_21039);
and U22120 (N_22120,N_20668,N_19173);
nor U22121 (N_22121,N_20090,N_19923);
and U22122 (N_22122,N_20476,N_19399);
and U22123 (N_22123,N_19386,N_20308);
nand U22124 (N_22124,N_18960,N_18911);
or U22125 (N_22125,N_19998,N_18977);
or U22126 (N_22126,N_20762,N_20437);
and U22127 (N_22127,N_19987,N_18827);
and U22128 (N_22128,N_19574,N_21476);
or U22129 (N_22129,N_20376,N_18875);
and U22130 (N_22130,N_19676,N_19158);
nand U22131 (N_22131,N_20655,N_21053);
and U22132 (N_22132,N_21120,N_21181);
nand U22133 (N_22133,N_21626,N_19643);
nor U22134 (N_22134,N_18888,N_20752);
nand U22135 (N_22135,N_20132,N_20585);
nand U22136 (N_22136,N_20275,N_20651);
xnor U22137 (N_22137,N_20719,N_19647);
and U22138 (N_22138,N_21597,N_20404);
nand U22139 (N_22139,N_19313,N_19700);
nand U22140 (N_22140,N_20429,N_19788);
and U22141 (N_22141,N_19338,N_19402);
xnor U22142 (N_22142,N_20487,N_18919);
nor U22143 (N_22143,N_19444,N_21554);
xor U22144 (N_22144,N_20171,N_19794);
nand U22145 (N_22145,N_21749,N_21459);
or U22146 (N_22146,N_20395,N_20517);
and U22147 (N_22147,N_19641,N_19782);
nor U22148 (N_22148,N_19564,N_21376);
nand U22149 (N_22149,N_19315,N_19910);
or U22150 (N_22150,N_19769,N_21802);
or U22151 (N_22151,N_20238,N_19180);
and U22152 (N_22152,N_21710,N_19461);
and U22153 (N_22153,N_21458,N_20677);
nand U22154 (N_22154,N_19654,N_19379);
nor U22155 (N_22155,N_18836,N_20288);
nand U22156 (N_22156,N_21097,N_21801);
and U22157 (N_22157,N_21224,N_21872);
and U22158 (N_22158,N_20842,N_18799);
nor U22159 (N_22159,N_20814,N_19150);
or U22160 (N_22160,N_21447,N_21366);
and U22161 (N_22161,N_20819,N_21187);
or U22162 (N_22162,N_19409,N_18984);
nor U22163 (N_22163,N_19848,N_20216);
or U22164 (N_22164,N_21200,N_19602);
xor U22165 (N_22165,N_20327,N_20036);
and U22166 (N_22166,N_18906,N_18798);
nand U22167 (N_22167,N_18751,N_19248);
xnor U22168 (N_22168,N_20314,N_21592);
and U22169 (N_22169,N_19970,N_20966);
and U22170 (N_22170,N_20390,N_21320);
nor U22171 (N_22171,N_20032,N_20302);
nand U22172 (N_22172,N_19849,N_20113);
xnor U22173 (N_22173,N_20215,N_19745);
or U22174 (N_22174,N_21100,N_20870);
nor U22175 (N_22175,N_19203,N_18905);
or U22176 (N_22176,N_19509,N_20850);
and U22177 (N_22177,N_21380,N_21643);
and U22178 (N_22178,N_20088,N_19785);
nor U22179 (N_22179,N_20249,N_19025);
nand U22180 (N_22180,N_19474,N_19960);
nand U22181 (N_22181,N_21291,N_20972);
nand U22182 (N_22182,N_21544,N_21316);
xnor U22183 (N_22183,N_21021,N_20765);
nand U22184 (N_22184,N_20106,N_20687);
nor U22185 (N_22185,N_20685,N_20526);
nand U22186 (N_22186,N_19013,N_19592);
or U22187 (N_22187,N_21279,N_20398);
nand U22188 (N_22188,N_21237,N_21275);
nor U22189 (N_22189,N_19163,N_19738);
nand U22190 (N_22190,N_21411,N_19889);
nand U22191 (N_22191,N_20980,N_19104);
and U22192 (N_22192,N_19866,N_20533);
nand U22193 (N_22193,N_19270,N_21318);
nor U22194 (N_22194,N_21450,N_18995);
nand U22195 (N_22195,N_21483,N_20638);
and U22196 (N_22196,N_21386,N_20649);
nand U22197 (N_22197,N_19562,N_20964);
xnor U22198 (N_22198,N_19988,N_19131);
nor U22199 (N_22199,N_21481,N_19459);
nand U22200 (N_22200,N_20068,N_19491);
or U22201 (N_22201,N_20522,N_21410);
or U22202 (N_22202,N_21541,N_21128);
or U22203 (N_22203,N_21303,N_19707);
nor U22204 (N_22204,N_21390,N_19121);
and U22205 (N_22205,N_20770,N_20640);
or U22206 (N_22206,N_19189,N_21247);
xnor U22207 (N_22207,N_21513,N_20286);
and U22208 (N_22208,N_19199,N_21054);
or U22209 (N_22209,N_20781,N_20427);
or U22210 (N_22210,N_19718,N_20486);
or U22211 (N_22211,N_19102,N_19984);
nor U22212 (N_22212,N_19778,N_19755);
or U22213 (N_22213,N_21751,N_20899);
or U22214 (N_22214,N_20890,N_20963);
nor U22215 (N_22215,N_20185,N_18932);
and U22216 (N_22216,N_21131,N_20543);
or U22217 (N_22217,N_20385,N_21613);
nand U22218 (N_22218,N_21023,N_20779);
or U22219 (N_22219,N_19630,N_20183);
nor U22220 (N_22220,N_21559,N_20634);
nor U22221 (N_22221,N_18993,N_19397);
nor U22222 (N_22222,N_21859,N_20159);
and U22223 (N_22223,N_20503,N_21110);
nor U22224 (N_22224,N_19099,N_19916);
nor U22225 (N_22225,N_20337,N_19515);
and U22226 (N_22226,N_20712,N_19118);
nand U22227 (N_22227,N_19114,N_18979);
and U22228 (N_22228,N_20570,N_18850);
and U22229 (N_22229,N_20959,N_19832);
nand U22230 (N_22230,N_19305,N_19067);
and U22231 (N_22231,N_21076,N_20598);
nand U22232 (N_22232,N_21848,N_19318);
xnor U22233 (N_22233,N_20579,N_21186);
nor U22234 (N_22234,N_19472,N_21863);
nor U22235 (N_22235,N_20645,N_21424);
and U22236 (N_22236,N_19749,N_21748);
and U22237 (N_22237,N_20575,N_20264);
nand U22238 (N_22238,N_21204,N_21296);
nor U22239 (N_22239,N_20248,N_19370);
nand U22240 (N_22240,N_18897,N_19495);
nand U22241 (N_22241,N_21272,N_19904);
or U22242 (N_22242,N_20573,N_20008);
nand U22243 (N_22243,N_19588,N_18927);
and U22244 (N_22244,N_19075,N_21730);
nor U22245 (N_22245,N_20797,N_21013);
xor U22246 (N_22246,N_19792,N_20424);
or U22247 (N_22247,N_20644,N_21654);
or U22248 (N_22248,N_21027,N_21645);
nand U22249 (N_22249,N_20730,N_20107);
or U22250 (N_22250,N_20067,N_20176);
nor U22251 (N_22251,N_19967,N_20357);
or U22252 (N_22252,N_20156,N_18840);
nor U22253 (N_22253,N_19920,N_19068);
nand U22254 (N_22254,N_18944,N_19947);
nand U22255 (N_22255,N_20255,N_19578);
and U22256 (N_22256,N_20681,N_19160);
and U22257 (N_22257,N_18885,N_21302);
nand U22258 (N_22258,N_20109,N_19570);
and U22259 (N_22259,N_20260,N_19862);
and U22260 (N_22260,N_19557,N_21675);
nor U22261 (N_22261,N_20785,N_20015);
nor U22262 (N_22262,N_19005,N_21619);
nor U22263 (N_22263,N_20242,N_19747);
nand U22264 (N_22264,N_19303,N_19770);
xnor U22265 (N_22265,N_21836,N_21514);
xor U22266 (N_22266,N_20285,N_18775);
and U22267 (N_22267,N_20877,N_20086);
nor U22268 (N_22268,N_20419,N_20435);
nand U22269 (N_22269,N_20396,N_19191);
nand U22270 (N_22270,N_20953,N_21660);
xor U22271 (N_22271,N_20612,N_21214);
and U22272 (N_22272,N_19886,N_19805);
nor U22273 (N_22273,N_21866,N_20035);
nand U22274 (N_22274,N_20843,N_21261);
and U22275 (N_22275,N_20020,N_20933);
nand U22276 (N_22276,N_19065,N_21387);
nor U22277 (N_22277,N_19276,N_20214);
nor U22278 (N_22278,N_21691,N_19545);
nand U22279 (N_22279,N_20804,N_20992);
nor U22280 (N_22280,N_21145,N_20204);
xnor U22281 (N_22281,N_18881,N_21443);
nand U22282 (N_22282,N_21377,N_20135);
nor U22283 (N_22283,N_20321,N_20173);
nor U22284 (N_22284,N_19391,N_21771);
nand U22285 (N_22285,N_20705,N_19513);
nor U22286 (N_22286,N_20147,N_21837);
and U22287 (N_22287,N_20918,N_21709);
nor U22288 (N_22288,N_20704,N_21538);
and U22289 (N_22289,N_19056,N_19353);
and U22290 (N_22290,N_20988,N_18803);
nor U22291 (N_22291,N_18990,N_19583);
nor U22292 (N_22292,N_19626,N_20237);
or U22293 (N_22293,N_21348,N_20616);
nor U22294 (N_22294,N_20669,N_18768);
nand U22295 (N_22295,N_21456,N_19069);
nor U22296 (N_22296,N_21511,N_20910);
or U22297 (N_22297,N_20354,N_21278);
nor U22298 (N_22298,N_18989,N_20673);
xor U22299 (N_22299,N_21591,N_21781);
nand U22300 (N_22300,N_19278,N_21765);
nor U22301 (N_22301,N_20557,N_19208);
nor U22302 (N_22302,N_18893,N_19352);
or U22303 (N_22303,N_19615,N_20326);
nor U22304 (N_22304,N_19994,N_21164);
nand U22305 (N_22305,N_20699,N_19818);
nand U22306 (N_22306,N_19255,N_20394);
and U22307 (N_22307,N_19990,N_18978);
nor U22308 (N_22308,N_18814,N_20686);
nor U22309 (N_22309,N_21283,N_21433);
and U22310 (N_22310,N_18853,N_18806);
and U22311 (N_22311,N_19869,N_21767);
or U22312 (N_22312,N_21539,N_21327);
nand U22313 (N_22313,N_19321,N_19763);
or U22314 (N_22314,N_21342,N_19484);
or U22315 (N_22315,N_19271,N_21676);
xor U22316 (N_22316,N_21508,N_21577);
or U22317 (N_22317,N_20563,N_19326);
and U22318 (N_22318,N_21385,N_19071);
or U22319 (N_22319,N_19600,N_19528);
nor U22320 (N_22320,N_19081,N_21336);
and U22321 (N_22321,N_19797,N_20071);
and U22322 (N_22322,N_18788,N_19378);
and U22323 (N_22323,N_20140,N_19418);
nand U22324 (N_22324,N_21185,N_19599);
xnor U22325 (N_22325,N_20745,N_19396);
nand U22326 (N_22326,N_19845,N_19876);
nor U22327 (N_22327,N_21492,N_21699);
or U22328 (N_22328,N_19346,N_21856);
nor U22329 (N_22329,N_19277,N_20583);
and U22330 (N_22330,N_20646,N_20967);
nand U22331 (N_22331,N_21438,N_21585);
or U22332 (N_22332,N_19325,N_19865);
or U22333 (N_22333,N_19991,N_19724);
xor U22334 (N_22334,N_18950,N_19363);
nor U22335 (N_22335,N_21542,N_19412);
or U22336 (N_22336,N_20000,N_20495);
xnor U22337 (N_22337,N_21028,N_20521);
nor U22338 (N_22338,N_21168,N_21713);
or U22339 (N_22339,N_19803,N_19293);
or U22340 (N_22340,N_20798,N_21091);
nand U22341 (N_22341,N_21354,N_19965);
nor U22342 (N_22342,N_20145,N_19742);
nand U22343 (N_22343,N_21663,N_21417);
and U22344 (N_22344,N_20430,N_18801);
nand U22345 (N_22345,N_20767,N_19801);
nor U22346 (N_22346,N_20913,N_20733);
nand U22347 (N_22347,N_21717,N_20811);
or U22348 (N_22348,N_19726,N_19508);
nor U22349 (N_22349,N_19149,N_21807);
and U22350 (N_22350,N_19427,N_19324);
or U22351 (N_22351,N_21157,N_19807);
nor U22352 (N_22352,N_19854,N_19666);
or U22353 (N_22353,N_21122,N_21227);
or U22354 (N_22354,N_19753,N_21738);
or U22355 (N_22355,N_21022,N_21112);
and U22356 (N_22356,N_19715,N_19016);
and U22357 (N_22357,N_21284,N_21504);
nor U22358 (N_22358,N_19717,N_21242);
or U22359 (N_22359,N_21861,N_21834);
nand U22360 (N_22360,N_21048,N_21226);
nand U22361 (N_22361,N_19502,N_20904);
and U22362 (N_22362,N_20393,N_21821);
or U22363 (N_22363,N_18965,N_18761);
and U22364 (N_22364,N_20760,N_20540);
or U22365 (N_22365,N_19047,N_18878);
nor U22366 (N_22366,N_21078,N_19760);
or U22367 (N_22367,N_19127,N_20999);
nand U22368 (N_22368,N_19359,N_21195);
nor U22369 (N_22369,N_20955,N_19811);
nand U22370 (N_22370,N_21576,N_19168);
nor U22371 (N_22371,N_21335,N_20230);
and U22372 (N_22372,N_19310,N_20097);
nand U22373 (N_22373,N_19454,N_19100);
and U22374 (N_22374,N_21090,N_20561);
or U22375 (N_22375,N_19627,N_18959);
nand U22376 (N_22376,N_20110,N_20488);
nand U22377 (N_22377,N_20609,N_19669);
and U22378 (N_22378,N_21644,N_21306);
nor U22379 (N_22379,N_20283,N_18868);
or U22380 (N_22380,N_21793,N_19584);
nor U22381 (N_22381,N_19441,N_19360);
nor U22382 (N_22382,N_19228,N_19744);
nand U22383 (N_22383,N_20845,N_20023);
xnor U22384 (N_22384,N_18922,N_20623);
or U22385 (N_22385,N_19620,N_21846);
nor U22386 (N_22386,N_20184,N_19119);
nand U22387 (N_22387,N_20566,N_20888);
nand U22388 (N_22388,N_19055,N_21125);
nand U22389 (N_22389,N_20675,N_21426);
nor U22390 (N_22390,N_20329,N_21398);
nand U22391 (N_22391,N_21156,N_18882);
nand U22392 (N_22392,N_20690,N_19633);
and U22393 (N_22393,N_20278,N_19332);
xnor U22394 (N_22394,N_19134,N_19695);
nand U22395 (N_22395,N_20011,N_21018);
xnor U22396 (N_22396,N_19380,N_20492);
nor U22397 (N_22397,N_20434,N_19252);
nor U22398 (N_22398,N_19116,N_18851);
and U22399 (N_22399,N_21843,N_20262);
nand U22400 (N_22400,N_20217,N_21561);
nand U22401 (N_22401,N_21682,N_20075);
nor U22402 (N_22402,N_20218,N_20549);
nor U22403 (N_22403,N_21003,N_21040);
nor U22404 (N_22404,N_18974,N_18898);
and U22405 (N_22405,N_19038,N_19684);
nor U22406 (N_22406,N_19458,N_20318);
xor U22407 (N_22407,N_20854,N_20587);
and U22408 (N_22408,N_20725,N_20021);
and U22409 (N_22409,N_20187,N_20296);
or U22410 (N_22410,N_19176,N_19980);
nand U22411 (N_22411,N_21494,N_21140);
nor U22412 (N_22412,N_20996,N_21098);
or U22413 (N_22413,N_20787,N_18884);
nand U22414 (N_22414,N_21305,N_21529);
nor U22415 (N_22415,N_19049,N_21031);
xnor U22416 (N_22416,N_21490,N_21701);
xor U22417 (N_22417,N_19453,N_19230);
xnor U22418 (N_22418,N_19188,N_20083);
or U22419 (N_22419,N_20127,N_20034);
nand U22420 (N_22420,N_21732,N_19568);
nor U22421 (N_22421,N_19392,N_19648);
and U22422 (N_22422,N_19476,N_19981);
nand U22423 (N_22423,N_19032,N_20319);
nand U22424 (N_22424,N_20062,N_20775);
xnor U22425 (N_22425,N_21368,N_21364);
nor U22426 (N_22426,N_21182,N_19522);
nor U22427 (N_22427,N_20592,N_19422);
nand U22428 (N_22428,N_21394,N_19962);
and U22429 (N_22429,N_19095,N_19927);
nor U22430 (N_22430,N_19177,N_21139);
nand U22431 (N_22431,N_21346,N_21718);
or U22432 (N_22432,N_21655,N_19155);
nor U22433 (N_22433,N_20691,N_21829);
nand U22434 (N_22434,N_18886,N_20082);
and U22435 (N_22435,N_18983,N_18980);
nor U22436 (N_22436,N_21196,N_19539);
and U22437 (N_22437,N_19946,N_19416);
and U22438 (N_22438,N_20399,N_19489);
nand U22439 (N_22439,N_20783,N_20251);
nand U22440 (N_22440,N_20507,N_19750);
or U22441 (N_22441,N_19622,N_21808);
nor U22442 (N_22442,N_19447,N_20791);
or U22443 (N_22443,N_18863,N_21002);
and U22444 (N_22444,N_21067,N_19419);
or U22445 (N_22445,N_21498,N_19768);
or U22446 (N_22446,N_19772,N_21629);
or U22447 (N_22447,N_19012,N_19170);
or U22448 (N_22448,N_18797,N_21220);
nor U22449 (N_22449,N_21250,N_21286);
nor U22450 (N_22450,N_19790,N_20087);
nand U22451 (N_22451,N_18908,N_20608);
and U22452 (N_22452,N_20663,N_20560);
nor U22453 (N_22453,N_21059,N_19651);
and U22454 (N_22454,N_20363,N_20350);
or U22455 (N_22455,N_19455,N_20081);
and U22456 (N_22456,N_18755,N_20149);
and U22457 (N_22457,N_21330,N_19462);
nor U22458 (N_22458,N_21070,N_18780);
nor U22459 (N_22459,N_21025,N_21741);
nor U22460 (N_22460,N_19193,N_18776);
or U22461 (N_22461,N_20055,N_19008);
or U22462 (N_22462,N_19253,N_21482);
xor U22463 (N_22463,N_21109,N_19628);
or U22464 (N_22464,N_20333,N_19948);
nand U22465 (N_22465,N_20300,N_18758);
nor U22466 (N_22466,N_20859,N_21785);
nor U22467 (N_22467,N_20190,N_19124);
and U22468 (N_22468,N_18946,N_19939);
xor U22469 (N_22469,N_21118,N_19467);
and U22470 (N_22470,N_19220,N_20530);
and U22471 (N_22471,N_21493,N_19408);
or U22472 (N_22472,N_19692,N_18778);
and U22473 (N_22473,N_19883,N_18883);
or U22474 (N_22474,N_20985,N_20456);
nor U22475 (N_22475,N_18849,N_18765);
nand U22476 (N_22476,N_18992,N_21745);
nand U22477 (N_22477,N_19542,N_19563);
xnor U22478 (N_22478,N_19404,N_19837);
xor U22479 (N_22479,N_21126,N_21672);
nor U22480 (N_22480,N_21780,N_21188);
nand U22481 (N_22481,N_19694,N_19873);
nor U22482 (N_22482,N_20105,N_21764);
and U22483 (N_22483,N_21199,N_20045);
and U22484 (N_22484,N_20200,N_21301);
nand U22485 (N_22485,N_20485,N_19440);
xnor U22486 (N_22486,N_21499,N_19575);
nand U22487 (N_22487,N_21431,N_19993);
and U22488 (N_22488,N_20887,N_20157);
and U22489 (N_22489,N_19686,N_20665);
nand U22490 (N_22490,N_19443,N_19954);
nor U22491 (N_22491,N_20990,N_18845);
nand U22492 (N_22492,N_20271,N_19014);
nor U22493 (N_22493,N_18805,N_19952);
xor U22494 (N_22494,N_21791,N_19510);
nor U22495 (N_22495,N_20451,N_20117);
nand U22496 (N_22496,N_20152,N_21773);
nand U22497 (N_22497,N_20377,N_21277);
or U22498 (N_22498,N_21203,N_20405);
nor U22499 (N_22499,N_20160,N_18951);
and U22500 (N_22500,N_19108,N_20191);
nand U22501 (N_22501,N_20595,N_21759);
nor U22502 (N_22502,N_19892,N_19126);
nand U22503 (N_22503,N_21642,N_20862);
and U22504 (N_22504,N_21123,N_20459);
nor U22505 (N_22505,N_20951,N_21252);
or U22506 (N_22506,N_20828,N_20954);
or U22507 (N_22507,N_19907,N_21611);
nand U22508 (N_22508,N_21606,N_19436);
and U22509 (N_22509,N_19577,N_19340);
and U22510 (N_22510,N_21462,N_21117);
nor U22511 (N_22511,N_21746,N_20891);
or U22512 (N_22512,N_19777,N_21512);
xnor U22513 (N_22513,N_19516,N_18880);
xor U22514 (N_22514,N_19637,N_20846);
nand U22515 (N_22515,N_19598,N_20969);
nor U22516 (N_22516,N_19682,N_20838);
and U22517 (N_22517,N_19009,N_20239);
or U22518 (N_22518,N_21149,N_20576);
nor U22519 (N_22519,N_19111,N_21582);
xor U22520 (N_22520,N_19162,N_21038);
nand U22521 (N_22521,N_18781,N_19347);
nand U22522 (N_22522,N_21206,N_20736);
nor U22523 (N_22523,N_19247,N_20968);
nand U22524 (N_22524,N_19330,N_19537);
or U22525 (N_22525,N_20550,N_20151);
or U22526 (N_22526,N_20243,N_20737);
or U22527 (N_22527,N_20835,N_21617);
and U22528 (N_22528,N_18879,N_20970);
or U22529 (N_22529,N_21826,N_19706);
or U22530 (N_22530,N_20641,N_21811);
nand U22531 (N_22531,N_21475,N_19989);
nor U22532 (N_22532,N_20993,N_21339);
and U22533 (N_22533,N_20294,N_19064);
xnor U22534 (N_22534,N_21739,N_20615);
and U22535 (N_22535,N_20209,N_20144);
or U22536 (N_22536,N_21111,N_19194);
nand U22537 (N_22537,N_21233,N_20601);
nand U22538 (N_22538,N_19113,N_20458);
and U22539 (N_22539,N_20529,N_18759);
nor U22540 (N_22540,N_20282,N_19290);
nand U22541 (N_22541,N_21222,N_20825);
and U22542 (N_22542,N_20676,N_18985);
xor U22543 (N_22543,N_19492,N_21669);
xor U22544 (N_22544,N_21216,N_21778);
or U22545 (N_22545,N_20772,N_20864);
xnor U22546 (N_22546,N_19802,N_19329);
nand U22547 (N_22547,N_19015,N_20662);
or U22548 (N_22548,N_21266,N_19141);
nand U22549 (N_22549,N_19490,N_19670);
nor U22550 (N_22550,N_19934,N_20768);
and U22551 (N_22551,N_19258,N_20077);
and U22552 (N_22552,N_19531,N_19799);
xnor U22553 (N_22553,N_20246,N_20975);
and U22554 (N_22554,N_21108,N_19004);
nand U22555 (N_22555,N_21467,N_19576);
or U22556 (N_22556,N_19895,N_21664);
nor U22557 (N_22557,N_19727,N_20426);
or U22558 (N_22558,N_20475,N_20254);
nor U22559 (N_22559,N_19137,N_19551);
or U22560 (N_22560,N_21480,N_19024);
or U22561 (N_22561,N_21593,N_20552);
or U22562 (N_22562,N_20431,N_21865);
and U22563 (N_22563,N_19296,N_19740);
and U22564 (N_22564,N_20581,N_21624);
or U22565 (N_22565,N_21361,N_19159);
and U22566 (N_22566,N_19018,N_21365);
nand U22567 (N_22567,N_20473,N_18940);
and U22568 (N_22568,N_19216,N_19003);
nor U22569 (N_22569,N_19259,N_21418);
and U22570 (N_22570,N_20343,N_19446);
nor U22571 (N_22571,N_19139,N_20053);
nor U22572 (N_22572,N_19784,N_19766);
nor U22573 (N_22573,N_20661,N_19308);
nand U22574 (N_22574,N_21497,N_20627);
and U22575 (N_22575,N_20931,N_21723);
and U22576 (N_22576,N_20416,N_20468);
or U22577 (N_22577,N_20724,N_19257);
and U22578 (N_22578,N_20301,N_18942);
and U22579 (N_22579,N_21560,N_21372);
or U22580 (N_22580,N_20729,N_20099);
nand U22581 (N_22581,N_21446,N_21453);
nor U22582 (N_22582,N_18782,N_20514);
or U22583 (N_22583,N_21171,N_20659);
nor U22584 (N_22584,N_21698,N_19587);
and U22585 (N_22585,N_20358,N_18873);
nor U22586 (N_22586,N_18967,N_19333);
or U22587 (N_22587,N_18804,N_19059);
and U22588 (N_22588,N_19655,N_21029);
or U22589 (N_22589,N_21425,N_21138);
nand U22590 (N_22590,N_21638,N_19696);
and U22591 (N_22591,N_19549,N_21383);
nor U22592 (N_22592,N_20914,N_20924);
or U22593 (N_22593,N_19093,N_19376);
nor U22594 (N_22594,N_19546,N_20867);
and U22595 (N_22595,N_20428,N_20133);
nand U22596 (N_22596,N_19423,N_19285);
or U22597 (N_22597,N_20766,N_21860);
or U22598 (N_22598,N_19240,N_20534);
nor U22599 (N_22599,N_21435,N_21062);
xnor U22600 (N_22600,N_19915,N_19714);
nand U22601 (N_22601,N_18994,N_20515);
nand U22602 (N_22602,N_19941,N_20060);
and U22603 (N_22603,N_21535,N_20784);
nor U22604 (N_22604,N_20709,N_18938);
nor U22605 (N_22605,N_21464,N_21340);
nor U22606 (N_22606,N_19868,N_20128);
nor U22607 (N_22607,N_20213,N_19297);
nand U22608 (N_22608,N_19500,N_20417);
nor U22609 (N_22609,N_19430,N_20057);
nand U22610 (N_22610,N_21760,N_20520);
nand U22611 (N_22611,N_19581,N_20538);
and U22612 (N_22612,N_20738,N_20324);
or U22613 (N_22613,N_21548,N_20016);
xor U22614 (N_22614,N_20369,N_21549);
nand U22615 (N_22615,N_19899,N_19097);
and U22616 (N_22616,N_19125,N_20666);
and U22617 (N_22617,N_19468,N_19051);
nor U22618 (N_22618,N_19721,N_21101);
and U22619 (N_22619,N_19078,N_21341);
or U22620 (N_22620,N_19044,N_21391);
nor U22621 (N_22621,N_20279,N_20818);
xnor U22622 (N_22622,N_20626,N_20799);
nand U22623 (N_22623,N_19215,N_19709);
nand U22624 (N_22624,N_19872,N_21641);
and U22625 (N_22625,N_21831,N_19087);
nor U22626 (N_22626,N_20273,N_19616);
nor U22627 (N_22627,N_20232,N_20436);
or U22628 (N_22628,N_19839,N_20630);
nand U22629 (N_22629,N_19206,N_20042);
and U22630 (N_22630,N_20801,N_20444);
or U22631 (N_22631,N_21044,N_19613);
and U22632 (N_22632,N_21630,N_19614);
and U22633 (N_22633,N_21835,N_20297);
or U22634 (N_22634,N_21491,N_21686);
nor U22635 (N_22635,N_19393,N_19917);
xor U22636 (N_22636,N_18958,N_19550);
nand U22637 (N_22637,N_19036,N_19765);
and U22638 (N_22638,N_19767,N_21384);
nand U22639 (N_22639,N_19579,N_18931);
xnor U22640 (N_22640,N_18918,N_21228);
or U22641 (N_22641,N_20111,N_21721);
nor U22642 (N_22642,N_20172,N_21375);
nor U22643 (N_22643,N_21132,N_19986);
xor U22644 (N_22644,N_20413,N_21590);
nor U22645 (N_22645,N_19507,N_19701);
nor U22646 (N_22646,N_20555,N_18914);
or U22647 (N_22647,N_21371,N_20137);
and U22648 (N_22648,N_18866,N_19795);
nand U22649 (N_22649,N_20267,N_19142);
nand U22650 (N_22650,N_19595,N_19752);
or U22651 (N_22651,N_21488,N_21614);
nor U22652 (N_22652,N_21119,N_19530);
xor U22653 (N_22653,N_20169,N_21649);
nor U22654 (N_22654,N_18821,N_20860);
nand U22655 (N_22655,N_20259,N_18847);
xnor U22656 (N_22656,N_21005,N_21167);
and U22657 (N_22657,N_21406,N_20916);
nand U22658 (N_22658,N_21007,N_19774);
nor U22659 (N_22659,N_21812,N_19512);
and U22660 (N_22660,N_21763,N_21049);
xnor U22661 (N_22661,N_19764,N_21263);
nor U22662 (N_22662,N_19327,N_19400);
nor U22663 (N_22663,N_19202,N_20177);
or U22664 (N_22664,N_21758,N_19372);
xnor U22665 (N_22665,N_19771,N_21215);
nor U22666 (N_22666,N_21402,N_21408);
or U22667 (N_22667,N_21130,N_21099);
or U22668 (N_22668,N_19885,N_18869);
nand U22669 (N_22669,N_20855,N_19719);
nor U22670 (N_22670,N_20812,N_20289);
or U22671 (N_22671,N_19662,N_21172);
or U22672 (N_22672,N_21092,N_21750);
xor U22673 (N_22673,N_18961,N_19183);
and U22674 (N_22674,N_21270,N_19729);
nor U22675 (N_22675,N_21551,N_19703);
and U22676 (N_22676,N_19968,N_20481);
or U22677 (N_22677,N_19681,N_20886);
nand U22678 (N_22678,N_20158,N_21106);
and U22679 (N_22679,N_21838,N_19902);
nor U22680 (N_22680,N_21211,N_20310);
and U22681 (N_22681,N_19855,N_20837);
nand U22682 (N_22682,N_21165,N_21774);
and U22683 (N_22683,N_18890,N_20876);
or U22684 (N_22684,N_20030,N_21176);
nor U22685 (N_22685,N_21703,N_19309);
or U22686 (N_22686,N_21087,N_21656);
or U22687 (N_22687,N_19387,N_19560);
xnor U22688 (N_22688,N_21666,N_19421);
or U22689 (N_22689,N_19677,N_20401);
or U22690 (N_22690,N_20636,N_21742);
and U22691 (N_22691,N_20755,N_19103);
nor U22692 (N_22692,N_21474,N_21806);
nand U22693 (N_22693,N_20293,N_19405);
nor U22694 (N_22694,N_19292,N_18800);
and U22695 (N_22695,N_20618,N_21072);
nand U22696 (N_22696,N_20336,N_20688);
xor U22697 (N_22697,N_19702,N_19900);
nor U22698 (N_22698,N_21308,N_19019);
and U22699 (N_22699,N_19943,N_20074);
or U22700 (N_22700,N_19625,N_20370);
nor U22701 (N_22701,N_19234,N_19739);
nor U22702 (N_22702,N_19274,N_20044);
nor U22703 (N_22703,N_20977,N_21229);
nand U22704 (N_22704,N_21212,N_21803);
and U22705 (N_22705,N_20112,N_19223);
and U22706 (N_22706,N_21208,N_20852);
nand U22707 (N_22707,N_19107,N_19586);
nand U22708 (N_22708,N_18889,N_19842);
nand U22709 (N_22709,N_19368,N_21213);
or U22710 (N_22710,N_21623,N_18779);
nor U22711 (N_22711,N_20589,N_20161);
nand U22712 (N_22712,N_20268,N_20317);
and U22713 (N_22713,N_20364,N_20411);
or U22714 (N_22714,N_19092,N_21862);
nand U22715 (N_22715,N_20981,N_21853);
or U22716 (N_22716,N_21570,N_19006);
nand U22717 (N_22717,N_19974,N_19758);
or U22718 (N_22718,N_19407,N_19365);
nor U22719 (N_22719,N_18795,N_20569);
xor U22720 (N_22720,N_20002,N_20658);
and U22721 (N_22721,N_21086,N_20446);
nand U22722 (N_22722,N_20715,N_21016);
or U22723 (N_22723,N_18912,N_18894);
nand U22724 (N_22724,N_20247,N_21310);
or U22725 (N_22725,N_21329,N_19030);
and U22726 (N_22726,N_20664,N_21262);
nor U22727 (N_22727,N_19000,N_20735);
nor U22728 (N_22728,N_20961,N_20463);
xor U22729 (N_22729,N_19406,N_19585);
nor U22730 (N_22730,N_19931,N_18947);
or U22731 (N_22731,N_19022,N_19559);
nor U22732 (N_22732,N_19775,N_21662);
and U22733 (N_22733,N_21521,N_21471);
or U22734 (N_22734,N_21604,N_21074);
nor U22735 (N_22735,N_21144,N_20912);
nand U22736 (N_22736,N_20018,N_19317);
nor U22737 (N_22737,N_19084,N_21162);
or U22738 (N_22738,N_19659,N_20684);
xor U22739 (N_22739,N_20439,N_21121);
xnor U22740 (N_22740,N_21809,N_19198);
and U22741 (N_22741,N_20816,N_19345);
or U22742 (N_22742,N_20700,N_19652);
nor U22743 (N_22743,N_21081,N_20619);
and U22744 (N_22744,N_19881,N_21457);
nand U22745 (N_22745,N_19284,N_19026);
and U22746 (N_22746,N_21094,N_20400);
nor U22747 (N_22747,N_21873,N_18750);
nor U22748 (N_22748,N_18839,N_21648);
nor U22749 (N_22749,N_19653,N_21804);
and U22750 (N_22750,N_20311,N_20123);
nor U22751 (N_22751,N_20927,N_21500);
xor U22752 (N_22752,N_21552,N_20656);
nand U22753 (N_22753,N_20957,N_19657);
and U22754 (N_22754,N_19037,N_21487);
and U22755 (N_22755,N_20986,N_21403);
and U22756 (N_22756,N_20355,N_20025);
nand U22757 (N_22757,N_19875,N_20203);
or U22758 (N_22758,N_20340,N_21849);
and U22759 (N_22759,N_20037,N_20713);
nor U22760 (N_22760,N_20617,N_21015);
and U22761 (N_22761,N_21681,N_19483);
nor U22762 (N_22762,N_21567,N_21088);
nand U22763 (N_22763,N_21864,N_20227);
nor U22764 (N_22764,N_19250,N_20150);
xnor U22765 (N_22765,N_21557,N_20906);
nand U22766 (N_22766,N_20717,N_20571);
and U22767 (N_22767,N_19322,N_19063);
or U22768 (N_22768,N_21687,N_18864);
nor U22769 (N_22769,N_21705,N_19566);
xnor U22770 (N_22770,N_20167,N_19912);
nor U22771 (N_22771,N_20546,N_21317);
and U22772 (N_22772,N_20625,N_21832);
nor U22773 (N_22773,N_19964,N_21716);
nand U22774 (N_22774,N_20794,N_21255);
nand U22775 (N_22775,N_21063,N_19506);
and U22776 (N_22776,N_20901,N_19082);
nor U22777 (N_22777,N_20108,N_20849);
nand U22778 (N_22778,N_21794,N_19298);
xnor U22779 (N_22779,N_20758,N_20584);
nor U22780 (N_22780,N_20639,N_19649);
nand U22781 (N_22781,N_19171,N_19820);
or U22782 (N_22782,N_18930,N_19282);
or U22783 (N_22783,N_19366,N_21736);
nor U22784 (N_22784,N_21449,N_21415);
nand U22785 (N_22785,N_21246,N_21036);
or U22786 (N_22786,N_21628,N_18859);
and U22787 (N_22787,N_21405,N_21839);
xnor U22788 (N_22788,N_21254,N_21332);
xor U22789 (N_22789,N_20073,N_18952);
nand U22790 (N_22790,N_19529,N_20013);
nand U22791 (N_22791,N_18999,N_20962);
and U22792 (N_22792,N_19634,N_19098);
nor U22793 (N_22793,N_19106,N_21823);
nor U22794 (N_22794,N_20188,N_21530);
nand U22795 (N_22795,N_20373,N_21518);
nor U22796 (N_22796,N_20104,N_20499);
nand U22797 (N_22797,N_18790,N_21589);
or U22798 (N_22798,N_20866,N_19520);
and U22799 (N_22799,N_20205,N_19477);
nand U22800 (N_22800,N_20815,N_20098);
or U22801 (N_22801,N_18910,N_21135);
xor U22802 (N_22802,N_19343,N_21412);
and U22803 (N_22803,N_21692,N_18762);
and U22804 (N_22804,N_20674,N_20863);
nand U22805 (N_22805,N_20223,N_20577);
or U22806 (N_22806,N_20450,N_19930);
or U22807 (N_22807,N_21241,N_20208);
and U22808 (N_22808,N_19511,N_19928);
nor U22809 (N_22809,N_21326,N_20048);
xor U22810 (N_22810,N_20679,N_20266);
nor U22811 (N_22811,N_20207,N_20657);
xor U22812 (N_22812,N_20974,N_21783);
nor U22813 (N_22813,N_19540,N_19261);
nand U22814 (N_22814,N_20440,N_18819);
xnor U22815 (N_22815,N_18877,N_20841);
and U22816 (N_22816,N_21634,N_21489);
nand U22817 (N_22817,N_21050,N_20874);
and U22818 (N_22818,N_18968,N_18855);
xor U22819 (N_22819,N_21805,N_19819);
nor U22820 (N_22820,N_21465,N_19348);
xor U22821 (N_22821,N_21869,N_20544);
nand U22822 (N_22822,N_21218,N_20771);
nor U22823 (N_22823,N_19992,N_20604);
or U22824 (N_22824,N_19371,N_21068);
nand U22825 (N_22825,N_20689,N_20007);
nor U22826 (N_22826,N_19746,N_20923);
nor U22827 (N_22827,N_21011,N_19538);
nor U22828 (N_22828,N_18917,N_19381);
nor U22829 (N_22829,N_20412,N_20882);
or U22830 (N_22830,N_19279,N_20046);
nand U22831 (N_22831,N_18941,N_21017);
and U22832 (N_22832,N_19565,N_20231);
or U22833 (N_22833,N_20367,N_19260);
nor U22834 (N_22834,N_20635,N_21731);
xnor U22835 (N_22835,N_21280,N_20381);
and U22836 (N_22836,N_19950,N_18970);
and U22837 (N_22837,N_19880,N_21520);
or U22838 (N_22838,N_19424,N_20165);
nand U22839 (N_22839,N_20102,N_19823);
or U22840 (N_22840,N_19631,N_20718);
nor U22841 (N_22841,N_19256,N_18838);
and U22842 (N_22842,N_19894,N_20392);
or U22843 (N_22843,N_19737,N_20415);
nand U22844 (N_22844,N_19887,N_19138);
nor U22845 (N_22845,N_20997,N_18981);
or U22846 (N_22846,N_20178,N_21043);
or U22847 (N_22847,N_20447,N_20479);
or U22848 (N_22848,N_20219,N_21525);
or U22849 (N_22849,N_21146,N_19227);
nand U22850 (N_22850,N_21362,N_20989);
nor U22851 (N_22851,N_19888,N_19110);
and U22852 (N_22852,N_19850,N_21810);
nand U22853 (N_22853,N_19225,N_20836);
or U22854 (N_22854,N_19328,N_21269);
nor U22855 (N_22855,N_21762,N_21006);
and U22856 (N_22856,N_21060,N_19020);
nand U22857 (N_22857,N_21867,N_21486);
nor U22858 (N_22858,N_19735,N_21338);
nor U22859 (N_22859,N_19567,N_19382);
nor U22860 (N_22860,N_20896,N_21631);
nor U22861 (N_22861,N_21328,N_20061);
nand U22862 (N_22862,N_19913,N_19334);
nor U22863 (N_22863,N_21586,N_18832);
or U22864 (N_22864,N_20210,N_18937);
or U22865 (N_22865,N_19374,N_20126);
xor U22866 (N_22866,N_20461,N_19940);
nor U22867 (N_22867,N_20116,N_20386);
xnor U22868 (N_22868,N_19800,N_19532);
nand U22869 (N_22869,N_18771,N_21154);
nor U22870 (N_22870,N_20531,N_19457);
nor U22871 (N_22871,N_19926,N_21178);
nor U22872 (N_22872,N_21769,N_19217);
nor U22873 (N_22873,N_21373,N_20049);
nand U22874 (N_22874,N_20383,N_19938);
and U22875 (N_22875,N_19663,N_20438);
or U22876 (N_22876,N_20432,N_20902);
and U22877 (N_22877,N_19010,N_21495);
or U22878 (N_22878,N_19096,N_19906);
nand U22879 (N_22879,N_21502,N_21009);
or U22880 (N_22880,N_19821,N_19645);
or U22881 (N_22881,N_20344,N_20605);
nand U22882 (N_22882,N_19473,N_19029);
nand U22883 (N_22883,N_18807,N_19384);
xor U22884 (N_22884,N_21419,N_19561);
nor U22885 (N_22885,N_21363,N_21221);
xor U22886 (N_22886,N_20024,N_19358);
or U22887 (N_22887,N_19169,N_20120);
or U22888 (N_22888,N_21350,N_19535);
xnor U22889 (N_22889,N_20298,N_21309);
nor U22890 (N_22890,N_20527,N_19414);
nand U22891 (N_22891,N_19269,N_21259);
nand U22892 (N_22892,N_21756,N_19949);
nand U22893 (N_22893,N_21102,N_21174);
xnor U22894 (N_22894,N_18763,N_21621);
and U22895 (N_22895,N_20274,N_18754);
nor U22896 (N_22896,N_20610,N_21295);
and U22897 (N_22897,N_21724,N_20789);
or U22898 (N_22898,N_21299,N_20491);
and U22899 (N_22899,N_20253,N_19937);
and U22900 (N_22900,N_20258,N_19526);
nand U22901 (N_22901,N_21496,N_18834);
or U22902 (N_22902,N_19058,N_21075);
or U22903 (N_22903,N_20720,N_20591);
nor U22904 (N_22904,N_18966,N_20984);
or U22905 (N_22905,N_20382,N_19264);
or U22906 (N_22906,N_18862,N_21571);
nor U22907 (N_22907,N_20212,N_19591);
or U22908 (N_22908,N_21515,N_20221);
nor U22909 (N_22909,N_19354,N_21399);
nor U22910 (N_22910,N_18817,N_21166);
and U22911 (N_22911,N_19644,N_19979);
and U22912 (N_22912,N_19689,N_19798);
nor U22913 (N_22913,N_21605,N_19190);
nor U22914 (N_22914,N_21082,N_19826);
nand U22915 (N_22915,N_19972,N_20186);
nor U22916 (N_22916,N_20498,N_19860);
and U22917 (N_22917,N_21374,N_19021);
xor U22918 (N_22918,N_20056,N_19178);
and U22919 (N_22919,N_20800,N_20330);
nor U22920 (N_22920,N_21287,N_21633);
nor U22921 (N_22921,N_19852,N_19693);
nand U22922 (N_22922,N_21133,N_21207);
or U22923 (N_22923,N_21527,N_19033);
or U22924 (N_22924,N_19822,N_19080);
and U22925 (N_22925,N_19857,N_20409);
nor U22926 (N_22926,N_20777,N_20222);
nor U22927 (N_22927,N_21743,N_19621);
and U22928 (N_22928,N_21673,N_21452);
nand U22929 (N_22929,N_20817,N_18871);
and U22930 (N_22930,N_19590,N_21516);
and U22931 (N_22931,N_18943,N_18988);
and U22932 (N_22932,N_20345,N_19521);
or U22933 (N_22933,N_19497,N_19420);
nand U22934 (N_22934,N_21700,N_19831);
nand U22935 (N_22935,N_19130,N_18936);
nand U22936 (N_22936,N_19664,N_20050);
nand U22937 (N_22937,N_21796,N_21640);
or U22938 (N_22938,N_19754,N_19465);
nor U22939 (N_22939,N_20322,N_19433);
nor U22940 (N_22940,N_18777,N_19073);
or U22941 (N_22941,N_21404,N_20163);
nand U22942 (N_22942,N_20885,N_20925);
or U22943 (N_22943,N_21004,N_20979);
nor U22944 (N_22944,N_20512,N_19231);
and U22945 (N_22945,N_21776,N_19824);
nor U22946 (N_22946,N_21334,N_19373);
nand U22947 (N_22947,N_21505,N_19045);
nand U22948 (N_22948,N_21042,N_19196);
or U22949 (N_22949,N_18909,N_18903);
nand U22950 (N_22950,N_18991,N_20096);
nand U22951 (N_22951,N_18956,N_18818);
nor U22952 (N_22952,N_19493,N_20474);
xor U22953 (N_22953,N_21105,N_21114);
xor U22954 (N_22954,N_20225,N_20572);
and U22955 (N_22955,N_20821,N_20448);
nand U22956 (N_22956,N_20683,N_20170);
or U22957 (N_22957,N_20305,N_20189);
and U22958 (N_22958,N_21107,N_20759);
or U22959 (N_22959,N_19074,N_19650);
nor U22960 (N_22960,N_19478,N_21707);
or U22961 (N_22961,N_20858,N_19983);
xnor U22962 (N_22962,N_19487,N_19226);
nand U22963 (N_22963,N_18925,N_19195);
nor U22964 (N_22964,N_20012,N_18902);
and U22965 (N_22965,N_20839,N_21550);
or U22966 (N_22966,N_20739,N_20698);
or U22967 (N_22967,N_20093,N_21436);
nand U22968 (N_22968,N_19851,N_18976);
nor U22969 (N_22969,N_19054,N_20365);
nor U22970 (N_22970,N_20982,N_21163);
and U22971 (N_22971,N_21219,N_20005);
nor U22972 (N_22972,N_20348,N_20403);
nand U22973 (N_22973,N_20019,N_19732);
or U22974 (N_22974,N_20965,N_20480);
or U22975 (N_22975,N_19610,N_21720);
or U22976 (N_22976,N_19921,N_19429);
xnor U22977 (N_22977,N_18769,N_21501);
or U22978 (N_22978,N_21815,N_21696);
or U22979 (N_22979,N_20751,N_20848);
nor U22980 (N_22980,N_21612,N_21344);
nand U22981 (N_22981,N_18949,N_19355);
or U22982 (N_22982,N_21693,N_19609);
or U22983 (N_22983,N_21069,N_19997);
nor U22984 (N_22984,N_19265,N_20822);
nor U22985 (N_22985,N_19128,N_19179);
xnor U22986 (N_22986,N_21777,N_20653);
and U22987 (N_22987,N_19336,N_19514);
and U22988 (N_22988,N_21083,N_20375);
nand U22989 (N_22989,N_18955,N_19601);
nor U22990 (N_22990,N_18848,N_19841);
xnor U22991 (N_22991,N_19830,N_19882);
or U22992 (N_22992,N_20810,N_20372);
nand U22993 (N_22993,N_19268,N_19375);
and U22994 (N_22994,N_19867,N_21093);
nand U22995 (N_22995,N_21784,N_21080);
and U22996 (N_22996,N_20872,N_19635);
and U22997 (N_22997,N_21148,N_19050);
or U22998 (N_22998,N_19350,N_20732);
nor U22999 (N_22999,N_18939,N_21519);
nand U23000 (N_23000,N_21152,N_21240);
and U23001 (N_23001,N_19524,N_20883);
nand U23002 (N_23002,N_21782,N_20425);
xor U23003 (N_23003,N_21034,N_19028);
xnor U23004 (N_23004,N_21298,N_20261);
nand U23005 (N_23005,N_19109,N_19244);
or U23006 (N_23006,N_20462,N_19356);
nand U23007 (N_23007,N_19398,N_19573);
xor U23008 (N_23008,N_20229,N_20995);
and U23009 (N_23009,N_20832,N_21608);
nand U23010 (N_23010,N_20761,N_21432);
nor U23011 (N_23011,N_19438,N_19847);
and U23012 (N_23012,N_21103,N_19544);
nor U23013 (N_23013,N_21037,N_19464);
nor U23014 (N_23014,N_19165,N_20723);
nor U23015 (N_23015,N_21180,N_20441);
nand U23016 (N_23016,N_21356,N_20911);
nor U23017 (N_23017,N_18824,N_19214);
or U23018 (N_23018,N_21115,N_20347);
nand U23019 (N_23019,N_18802,N_20978);
or U23020 (N_23020,N_19853,N_19896);
and U23021 (N_23021,N_20059,N_19756);
or U23022 (N_23022,N_19001,N_20539);
or U23023 (N_23023,N_19959,N_21690);
and U23024 (N_23024,N_20265,N_21555);
nand U23025 (N_23025,N_20043,N_19844);
nand U23026 (N_23026,N_21753,N_20827);
nand U23027 (N_23027,N_21652,N_19944);
nor U23028 (N_23028,N_20754,N_19323);
nor U23029 (N_23029,N_20361,N_19680);
nor U23030 (N_23030,N_20711,N_21141);
and U23031 (N_23031,N_20956,N_21779);
nand U23032 (N_23032,N_21517,N_21671);
or U23033 (N_23033,N_21313,N_20780);
xor U23034 (N_23034,N_19571,N_21333);
or U23035 (N_23035,N_19720,N_19589);
nor U23036 (N_23036,N_19736,N_20680);
or U23037 (N_23037,N_21276,N_20805);
or U23038 (N_23038,N_19153,N_19210);
and U23039 (N_23039,N_21129,N_21772);
nor U23040 (N_23040,N_19132,N_21636);
and U23041 (N_23041,N_19236,N_19612);
nand U23042 (N_23042,N_18843,N_21627);
nor U23043 (N_23043,N_21565,N_19905);
nand U23044 (N_23044,N_19810,N_19083);
nor U23045 (N_23045,N_18812,N_19112);
xor U23046 (N_23046,N_21564,N_21159);
or U23047 (N_23047,N_20524,N_20749);
nand U23048 (N_23048,N_20041,N_19879);
xor U23049 (N_23049,N_19723,N_20652);
nand U23050 (N_23050,N_19273,N_21470);
or U23051 (N_23051,N_21575,N_20621);
and U23052 (N_23052,N_20454,N_18962);
nand U23053 (N_23053,N_19734,N_21437);
and U23054 (N_23054,N_20607,N_20477);
nand U23055 (N_23055,N_19395,N_21251);
nor U23056 (N_23056,N_18854,N_21532);
nor U23057 (N_23057,N_21646,N_21689);
nor U23058 (N_23058,N_21051,N_19466);
and U23059 (N_23059,N_20076,N_21569);
and U23060 (N_23060,N_20813,N_20753);
nand U23061 (N_23061,N_21253,N_21855);
nor U23062 (N_23062,N_21020,N_19043);
nor U23063 (N_23063,N_19147,N_18935);
or U23064 (N_23064,N_20948,N_21847);
and U23065 (N_23065,N_19197,N_20118);
nor U23066 (N_23066,N_18811,N_21822);
xnor U23067 (N_23067,N_20129,N_20421);
and U23068 (N_23068,N_19187,N_21727);
or U23069 (N_23069,N_20408,N_20823);
and U23070 (N_23070,N_21169,N_21265);
and U23071 (N_23071,N_19299,N_20084);
nor U23072 (N_23072,N_21236,N_21685);
nand U23073 (N_23073,N_20750,N_19957);
and U23074 (N_23074,N_21661,N_21136);
nor U23075 (N_23075,N_20940,N_19017);
nor U23076 (N_23076,N_19031,N_21307);
or U23077 (N_23077,N_21400,N_20142);
and U23078 (N_23078,N_19351,N_20502);
and U23079 (N_23079,N_20449,N_20269);
or U23080 (N_23080,N_19893,N_21235);
nor U23081 (N_23081,N_20125,N_21528);
xnor U23082 (N_23082,N_19079,N_19488);
nor U23083 (N_23083,N_19874,N_20501);
and U23084 (N_23084,N_21479,N_18874);
and U23085 (N_23085,N_20307,N_21209);
or U23086 (N_23086,N_19791,N_19951);
nand U23087 (N_23087,N_19357,N_19553);
xor U23088 (N_23088,N_20632,N_19733);
nand U23089 (N_23089,N_20548,N_20384);
nor U23090 (N_23090,N_19182,N_21300);
and U23091 (N_23091,N_21061,N_20179);
or U23092 (N_23092,N_18772,N_21147);
nand U23093 (N_23093,N_18901,N_20009);
or U23094 (N_23094,N_21858,N_21160);
or U23095 (N_23095,N_19953,N_18915);
nor U23096 (N_23096,N_19632,N_21651);
or U23097 (N_23097,N_18891,N_19123);
nand U23098 (N_23098,N_19716,N_20168);
and U23099 (N_23099,N_21161,N_21177);
or U23100 (N_23100,N_20139,N_19812);
and U23101 (N_23101,N_19229,N_19301);
and U23102 (N_23102,N_21000,N_21874);
or U23103 (N_23103,N_20328,N_19932);
nor U23104 (N_23104,N_19759,N_20040);
and U23105 (N_23105,N_18822,N_20820);
or U23106 (N_23106,N_21609,N_21728);
and U23107 (N_23107,N_18786,N_18766);
xnor U23108 (N_23108,N_19956,N_18828);
nand U23109 (N_23109,N_19525,N_21722);
nand U23110 (N_23110,N_18857,N_20295);
xnor U23111 (N_23111,N_18872,N_21434);
nor U23112 (N_23112,N_21584,N_20063);
xnor U23113 (N_23113,N_21677,N_19711);
or U23114 (N_23114,N_20620,N_21155);
nor U23115 (N_23115,N_19996,N_19890);
nand U23116 (N_23116,N_18826,N_21381);
or U23117 (N_23117,N_19787,N_20631);
nand U23118 (N_23118,N_19864,N_20374);
or U23119 (N_23119,N_19040,N_19148);
or U23120 (N_23120,N_19377,N_18844);
xor U23121 (N_23121,N_20235,N_19077);
or U23122 (N_23122,N_19908,N_20551);
nor U23123 (N_23123,N_21534,N_21747);
and U23124 (N_23124,N_20010,N_20728);
nor U23125 (N_23125,N_20281,N_19439);
xnor U23126 (N_23126,N_20614,N_18865);
and U23127 (N_23127,N_20628,N_20637);
nand U23128 (N_23128,N_21322,N_19251);
and U23129 (N_23129,N_19731,N_19364);
and U23130 (N_23130,N_20893,N_19212);
or U23131 (N_23131,N_18820,N_21430);
nand U23132 (N_23132,N_21359,N_18996);
and U23133 (N_23133,N_20731,N_20921);
nor U23134 (N_23134,N_20537,N_21820);
or U23135 (N_23135,N_19235,N_19789);
and U23136 (N_23136,N_19656,N_21347);
and U23137 (N_23137,N_21351,N_20873);
and U23138 (N_23138,N_20793,N_19815);
nor U23139 (N_23139,N_20457,N_19089);
nand U23140 (N_23140,N_20695,N_21833);
nor U23141 (N_23141,N_21170,N_20881);
or U23142 (N_23142,N_19638,N_18975);
nor U23143 (N_23143,N_21639,N_19136);
nor U23144 (N_23144,N_19597,N_20467);
nor U23145 (N_23145,N_20192,N_21600);
or U23146 (N_23146,N_20747,N_20694);
nor U23147 (N_23147,N_19485,N_19667);
nand U23148 (N_23148,N_19809,N_20545);
nor U23149 (N_23149,N_20707,N_19582);
and U23150 (N_23150,N_19331,N_20599);
nand U23151 (N_23151,N_20746,N_20493);
nand U23152 (N_23152,N_21697,N_21841);
nor U23153 (N_23153,N_19211,N_19713);
nand U23154 (N_23154,N_20148,N_19294);
nand U23155 (N_23155,N_20490,N_19603);
or U23156 (N_23156,N_19929,N_21248);
nand U23157 (N_23157,N_19062,N_19833);
nor U23158 (N_23158,N_19688,N_19773);
nor U23159 (N_23159,N_18831,N_20897);
nand U23160 (N_23160,N_18752,N_19388);
nand U23161 (N_23161,N_20600,N_19971);
and U23162 (N_23162,N_21469,N_21057);
nor U23163 (N_23163,N_20824,N_20422);
or U23164 (N_23164,N_18785,N_20790);
or U23165 (N_23165,N_19505,N_20920);
and U23166 (N_23166,N_20483,N_20299);
and U23167 (N_23167,N_19922,N_21282);
or U23168 (N_23168,N_19085,N_20353);
and U23169 (N_23169,N_18887,N_20834);
nor U23170 (N_23170,N_20303,N_21409);
nand U23171 (N_23171,N_21066,N_21484);
nand U23172 (N_23172,N_20505,N_19233);
and U23173 (N_23173,N_19482,N_19101);
nor U23174 (N_23174,N_20795,N_19779);
xnor U23175 (N_23175,N_20721,N_21137);
or U23176 (N_23176,N_18842,N_19973);
nor U23177 (N_23177,N_18954,N_20406);
nor U23178 (N_23178,N_21657,N_21744);
nand U23179 (N_23179,N_19143,N_19426);
or U23180 (N_23180,N_21524,N_20803);
or U23181 (N_23181,N_18963,N_21153);
nor U23182 (N_23182,N_21010,N_20141);
or U23183 (N_23183,N_21150,N_19618);
nor U23184 (N_23184,N_19480,N_19672);
nand U23185 (N_23185,N_21540,N_20606);
or U23186 (N_23186,N_20907,N_21507);
and U23187 (N_23187,N_20898,N_19172);
nor U23188 (N_23188,N_18920,N_19164);
nand U23189 (N_23189,N_18971,N_20094);
or U23190 (N_23190,N_21343,N_21714);
nor U23191 (N_23191,N_19342,N_21840);
nor U23192 (N_23192,N_20504,N_19135);
xor U23193 (N_23193,N_20830,N_19122);
xnor U23194 (N_23194,N_19642,N_20325);
and U23195 (N_23195,N_21179,N_21695);
nand U23196 (N_23196,N_18830,N_19117);
nor U23197 (N_23197,N_20100,N_19475);
and U23198 (N_23198,N_19536,N_19035);
and U23199 (N_23199,N_19678,N_20029);
xor U23200 (N_23200,N_19757,N_19319);
and U23201 (N_23201,N_20146,N_20124);
nor U23202 (N_23202,N_21143,N_20070);
and U23203 (N_23203,N_19280,N_21297);
xor U23204 (N_23204,N_21245,N_20991);
nor U23205 (N_23205,N_20338,N_20869);
nor U23206 (N_23206,N_21142,N_19133);
or U23207 (N_23207,N_21819,N_20080);
or U23208 (N_23208,N_18860,N_21440);
and U23209 (N_23209,N_21357,N_21607);
xnor U23210 (N_23210,N_19307,N_21008);
and U23211 (N_23211,N_19070,N_18856);
or U23212 (N_23212,N_19167,N_21089);
or U23213 (N_23213,N_20028,N_19090);
or U23214 (N_23214,N_20470,N_19088);
or U23215 (N_23215,N_21079,N_19448);
or U23216 (N_23216,N_21024,N_19607);
nand U23217 (N_23217,N_19919,N_20701);
nor U23218 (N_23218,N_21223,N_20588);
nor U23219 (N_23219,N_21045,N_20066);
xor U23220 (N_23220,N_20312,N_20774);
or U23221 (N_23221,N_19205,N_20489);
and U23222 (N_23222,N_20115,N_19843);
xor U23223 (N_23223,N_21073,N_18964);
nand U23224 (N_23224,N_18945,N_21369);
or U23225 (N_23225,N_21827,N_21239);
nand U23226 (N_23226,N_20175,N_20245);
nand U23227 (N_23227,N_20875,N_19636);
or U23228 (N_23228,N_19011,N_19963);
and U23229 (N_23229,N_19813,N_19624);
or U23230 (N_23230,N_20064,N_21740);
and U23231 (N_23231,N_20315,N_21598);
nand U23232 (N_23232,N_21522,N_20181);
and U23233 (N_23233,N_21019,N_21816);
nand U23234 (N_23234,N_19394,N_19976);
nor U23235 (N_23235,N_19543,N_20359);
or U23236 (N_23236,N_18953,N_21702);
nor U23237 (N_23237,N_19209,N_20938);
and U23238 (N_23238,N_21389,N_20511);
xor U23239 (N_23239,N_19241,N_19337);
or U23240 (N_23240,N_19156,N_19066);
xnor U23241 (N_23241,N_20513,N_19140);
and U23242 (N_23242,N_21388,N_21232);
nand U23243 (N_23243,N_19239,N_19403);
and U23244 (N_23244,N_20287,N_19362);
nor U23245 (N_23245,N_21546,N_20153);
and U23246 (N_23246,N_18896,N_20613);
xnor U23247 (N_23247,N_19834,N_20402);
or U23248 (N_23248,N_20593,N_20703);
nand U23249 (N_23249,N_19829,N_19836);
nand U23250 (N_23250,N_21427,N_20932);
nand U23251 (N_23251,N_21579,N_20380);
nor U23252 (N_23252,N_19314,N_18987);
nand U23253 (N_23253,N_21786,N_20054);
nand U23254 (N_23254,N_19494,N_20928);
and U23255 (N_23255,N_20987,N_20807);
nor U23256 (N_23256,N_19783,N_20236);
nand U23257 (N_23257,N_18760,N_19129);
or U23258 (N_23258,N_20263,N_21553);
nor U23259 (N_23259,N_19828,N_20291);
nor U23260 (N_23260,N_21012,N_20622);
nor U23261 (N_23261,N_21845,N_20047);
nand U23262 (N_23262,N_21444,N_21537);
nand U23263 (N_23263,N_19288,N_20568);
xor U23264 (N_23264,N_21325,N_20342);
nor U23265 (N_23265,N_19646,N_20052);
nor U23266 (N_23266,N_20270,N_19748);
or U23267 (N_23267,N_21047,N_19238);
xnor U23268 (N_23268,N_19304,N_20672);
or U23269 (N_23269,N_20878,N_19685);
nand U23270 (N_23270,N_21134,N_18997);
nand U23271 (N_23271,N_19046,N_19302);
xor U23272 (N_23272,N_19344,N_19174);
nand U23273 (N_23273,N_21201,N_20740);
nor U23274 (N_23274,N_19417,N_18900);
and U23275 (N_23275,N_19287,N_21587);
and U23276 (N_23276,N_21225,N_21711);
or U23277 (N_23277,N_21870,N_21775);
or U23278 (N_23278,N_20629,N_20586);
xor U23279 (N_23279,N_21603,N_21244);
or U23280 (N_23280,N_19470,N_19898);
nor U23281 (N_23281,N_18793,N_19859);
or U23282 (N_23282,N_21175,N_19698);
and U23283 (N_23283,N_21193,N_21678);
and U23284 (N_23284,N_19151,N_21198);
nand U23285 (N_23285,N_20420,N_21818);
nor U23286 (N_23286,N_19246,N_19039);
or U23287 (N_23287,N_21477,N_19091);
and U23288 (N_23288,N_20478,N_21583);
or U23289 (N_23289,N_21694,N_20671);
and U23290 (N_23290,N_19389,N_20114);
and U23291 (N_23291,N_19945,N_18809);
nand U23292 (N_23292,N_19697,N_19878);
and U23293 (N_23293,N_20857,N_18923);
nand U23294 (N_23294,N_20506,N_18841);
nor U23295 (N_23295,N_20542,N_19548);
nor U23296 (N_23296,N_19665,N_19580);
or U23297 (N_23297,N_21271,N_20602);
and U23298 (N_23298,N_20884,N_20909);
nand U23299 (N_23299,N_21355,N_20518);
and U23300 (N_23300,N_19428,N_18948);
or U23301 (N_23301,N_21158,N_19877);
xor U23302 (N_23302,N_19604,N_21766);
and U23303 (N_23303,N_19341,N_20806);
and U23304 (N_23304,N_21679,N_21795);
and U23305 (N_23305,N_18895,N_19619);
nor U23306 (N_23306,N_20556,N_20194);
and U23307 (N_23307,N_21752,N_20716);
and U23308 (N_23308,N_19911,N_21842);
and U23309 (N_23309,N_18933,N_19661);
and U23310 (N_23310,N_20547,N_20469);
or U23311 (N_23311,N_21423,N_21260);
or U23312 (N_23312,N_21610,N_20423);
nand U23313 (N_23313,N_21184,N_21658);
or U23314 (N_23314,N_20482,N_19295);
nor U23315 (N_23315,N_21578,N_20536);
and U23316 (N_23316,N_19048,N_21787);
and U23317 (N_23317,N_20130,N_21268);
and U23318 (N_23318,N_21442,N_21523);
or U23319 (N_23319,N_18815,N_21231);
nand U23320 (N_23320,N_20574,N_20971);
nand U23321 (N_23321,N_20500,N_19262);
nor U23322 (N_23322,N_20580,N_19041);
or U23323 (N_23323,N_19861,N_19835);
nor U23324 (N_23324,N_21104,N_19072);
or U23325 (N_23325,N_20596,N_19611);
nand U23326 (N_23326,N_20973,N_20496);
nor U23327 (N_23327,N_21058,N_18904);
nor U23328 (N_23328,N_19316,N_20465);
and U23329 (N_23329,N_19925,N_21084);
and U23330 (N_23330,N_20226,N_21151);
nand U23331 (N_23331,N_19053,N_21733);
or U23332 (N_23332,N_21632,N_20840);
nor U23333 (N_23333,N_21046,N_20072);
and U23334 (N_23334,N_20727,N_19704);
nand U23335 (N_23335,N_20941,N_19425);
or U23336 (N_23336,N_21616,N_19897);
and U23337 (N_23337,N_20559,N_21064);
or U23338 (N_23338,N_18792,N_20809);
or U23339 (N_23339,N_20460,N_19660);
or U23340 (N_23340,N_20387,N_19863);
nand U23341 (N_23341,N_21668,N_21345);
or U23342 (N_23342,N_19450,N_20516);
nor U23343 (N_23343,N_18791,N_19556);
nand U23344 (N_23344,N_21770,N_21461);
nor U23345 (N_23345,N_20078,N_20472);
nor U23346 (N_23346,N_18969,N_20241);
nor U23347 (N_23347,N_20939,N_21249);
and U23348 (N_23348,N_21445,N_19504);
nand U23349 (N_23349,N_20782,N_20926);
nor U23350 (N_23350,N_20252,N_19978);
nand U23351 (N_23351,N_20304,N_20134);
and U23352 (N_23352,N_19668,N_21637);
xor U23353 (N_23353,N_21194,N_20742);
or U23354 (N_23354,N_18861,N_21850);
nor U23355 (N_23355,N_20352,N_20829);
and U23356 (N_23356,N_18916,N_19042);
or U23357 (N_23357,N_20944,N_19437);
nor U23358 (N_23358,N_20346,N_20895);
and U23359 (N_23359,N_19289,N_19449);
nand U23360 (N_23360,N_21065,N_21238);
nor U23361 (N_23361,N_20889,N_20092);
nand U23362 (N_23362,N_20155,N_20038);
and U23363 (N_23363,N_19606,N_20418);
nor U23364 (N_23364,N_20643,N_21719);
and U23365 (N_23365,N_19184,N_21688);
nor U23366 (N_23366,N_19629,N_19730);
nand U23367 (N_23367,N_19320,N_19687);
or U23368 (N_23368,N_19415,N_21670);
nor U23369 (N_23369,N_20316,N_21413);
or U23370 (N_23370,N_20879,N_20535);
xnor U23371 (N_23371,N_19463,N_20509);
xor U23372 (N_23372,N_19367,N_19534);
nand U23373 (N_23373,N_21509,N_20597);
xnor U23374 (N_23374,N_20332,N_19145);
or U23375 (N_23375,N_18837,N_20292);
xnor U23376 (N_23376,N_21382,N_20937);
or U23377 (N_23377,N_21392,N_20741);
xnor U23378 (N_23378,N_20201,N_19312);
and U23379 (N_23379,N_20796,N_20650);
or U23380 (N_23380,N_20748,N_19181);
and U23381 (N_23381,N_21113,N_20942);
or U23382 (N_23382,N_19267,N_21531);
and U23383 (N_23383,N_20642,N_19023);
and U23384 (N_23384,N_19115,N_21543);
nand U23385 (N_23385,N_20143,N_21868);
nor U23386 (N_23386,N_20553,N_19232);
xnor U23387 (N_23387,N_20240,N_20950);
nand U23388 (N_23388,N_19263,N_21454);
or U23389 (N_23389,N_19166,N_20847);
nor U23390 (N_23390,N_20257,N_20853);
and U23391 (N_23391,N_21116,N_18770);
and U23392 (N_23392,N_21267,N_18823);
nor U23393 (N_23393,N_18825,N_19445);
and U23394 (N_23394,N_20180,N_19254);
or U23395 (N_23395,N_20930,N_21304);
nand U23396 (N_23396,N_20356,N_20541);
or U23397 (N_23397,N_19640,N_20647);
or U23398 (N_23398,N_19002,N_19958);
or U23399 (N_23399,N_19369,N_21378);
nor U23400 (N_23400,N_19207,N_20182);
and U23401 (N_23401,N_18870,N_19161);
xnor U23402 (N_23402,N_20565,N_20947);
nor U23403 (N_23403,N_20494,N_21667);
xor U23404 (N_23404,N_20331,N_21871);
and U23405 (N_23405,N_18767,N_19518);
or U23406 (N_23406,N_19728,N_19935);
xor U23407 (N_23407,N_21852,N_20808);
nand U23408 (N_23408,N_20197,N_21127);
xor U23409 (N_23409,N_21857,N_19452);
nand U23410 (N_23410,N_19218,N_20196);
xor U23411 (N_23411,N_21290,N_21472);
xnor U23412 (N_23412,N_20594,N_19479);
nand U23413 (N_23413,N_20554,N_19596);
or U23414 (N_23414,N_21726,N_20908);
and U23415 (N_23415,N_20868,N_20756);
nand U23416 (N_23416,N_19311,N_18907);
xnor U23417 (N_23417,N_20833,N_18794);
nor U23418 (N_23418,N_20121,N_20564);
or U23419 (N_23419,N_19213,N_19936);
or U23420 (N_23420,N_20001,N_21026);
and U23421 (N_23421,N_18892,N_18796);
xor U23422 (N_23422,N_21601,N_21602);
and U23423 (N_23423,N_21588,N_20861);
nand U23424 (N_23424,N_19383,N_19955);
and U23425 (N_23425,N_20844,N_20136);
and U23426 (N_23426,N_21311,N_20195);
nand U23427 (N_23427,N_21292,N_20378);
and U23428 (N_23428,N_21737,N_18774);
xnor U23429 (N_23429,N_19496,N_21096);
and U23430 (N_23430,N_21353,N_19969);
or U23431 (N_23431,N_19471,N_21395);
nand U23432 (N_23432,N_19712,N_19918);
or U23433 (N_23433,N_18816,N_20508);
nor U23434 (N_23434,N_20764,N_21319);
nor U23435 (N_23435,N_19623,N_21033);
and U23436 (N_23436,N_20433,N_21680);
and U23437 (N_23437,N_20667,N_21081);
and U23438 (N_23438,N_19682,N_18814);
or U23439 (N_23439,N_19794,N_21552);
nand U23440 (N_23440,N_19245,N_20256);
xor U23441 (N_23441,N_21551,N_20403);
and U23442 (N_23442,N_21697,N_21330);
nor U23443 (N_23443,N_18911,N_21475);
xnor U23444 (N_23444,N_19901,N_19293);
nand U23445 (N_23445,N_20482,N_20081);
nand U23446 (N_23446,N_21709,N_21129);
nand U23447 (N_23447,N_20891,N_21105);
nor U23448 (N_23448,N_20260,N_21472);
nor U23449 (N_23449,N_21804,N_20792);
or U23450 (N_23450,N_19806,N_21574);
nand U23451 (N_23451,N_20146,N_19354);
nand U23452 (N_23452,N_20299,N_20340);
and U23453 (N_23453,N_19668,N_20252);
or U23454 (N_23454,N_19129,N_21304);
and U23455 (N_23455,N_20993,N_19758);
and U23456 (N_23456,N_19286,N_20168);
or U23457 (N_23457,N_19733,N_20310);
nor U23458 (N_23458,N_21299,N_21151);
nor U23459 (N_23459,N_20188,N_21350);
and U23460 (N_23460,N_20210,N_21676);
nand U23461 (N_23461,N_21345,N_20367);
nor U23462 (N_23462,N_21782,N_21846);
and U23463 (N_23463,N_19523,N_19126);
nand U23464 (N_23464,N_19193,N_20724);
nor U23465 (N_23465,N_21223,N_19521);
nand U23466 (N_23466,N_20209,N_20511);
and U23467 (N_23467,N_18856,N_19911);
and U23468 (N_23468,N_19530,N_21738);
or U23469 (N_23469,N_21595,N_19406);
or U23470 (N_23470,N_21796,N_21022);
nor U23471 (N_23471,N_21380,N_20628);
nand U23472 (N_23472,N_20636,N_20146);
and U23473 (N_23473,N_20992,N_21040);
nor U23474 (N_23474,N_20739,N_21477);
xor U23475 (N_23475,N_21776,N_21054);
and U23476 (N_23476,N_21101,N_19166);
and U23477 (N_23477,N_21168,N_19848);
or U23478 (N_23478,N_20141,N_19062);
nand U23479 (N_23479,N_19223,N_21129);
or U23480 (N_23480,N_19589,N_20615);
xor U23481 (N_23481,N_19868,N_20855);
xnor U23482 (N_23482,N_19692,N_21509);
xnor U23483 (N_23483,N_21159,N_21300);
or U23484 (N_23484,N_21329,N_21494);
nand U23485 (N_23485,N_20749,N_21685);
and U23486 (N_23486,N_20965,N_20150);
nor U23487 (N_23487,N_19635,N_19467);
or U23488 (N_23488,N_20979,N_20493);
xnor U23489 (N_23489,N_20197,N_20433);
nor U23490 (N_23490,N_21367,N_20668);
nand U23491 (N_23491,N_19260,N_18767);
and U23492 (N_23492,N_21774,N_19654);
and U23493 (N_23493,N_20464,N_21565);
and U23494 (N_23494,N_21218,N_19919);
nand U23495 (N_23495,N_21627,N_19769);
nor U23496 (N_23496,N_19260,N_20028);
or U23497 (N_23497,N_21590,N_20609);
nand U23498 (N_23498,N_19136,N_19331);
and U23499 (N_23499,N_19967,N_18793);
or U23500 (N_23500,N_20632,N_21512);
and U23501 (N_23501,N_18811,N_21518);
nor U23502 (N_23502,N_20470,N_19751);
and U23503 (N_23503,N_20182,N_21665);
xor U23504 (N_23504,N_20189,N_21596);
nor U23505 (N_23505,N_20394,N_19528);
and U23506 (N_23506,N_19710,N_19860);
and U23507 (N_23507,N_21196,N_19352);
and U23508 (N_23508,N_20849,N_21566);
and U23509 (N_23509,N_20492,N_19887);
nor U23510 (N_23510,N_21290,N_18857);
or U23511 (N_23511,N_19383,N_20021);
nand U23512 (N_23512,N_21356,N_19569);
nand U23513 (N_23513,N_18806,N_19978);
and U23514 (N_23514,N_19014,N_19199);
nor U23515 (N_23515,N_21216,N_21520);
or U23516 (N_23516,N_19256,N_20487);
and U23517 (N_23517,N_20638,N_20947);
and U23518 (N_23518,N_20512,N_18896);
nand U23519 (N_23519,N_21485,N_20318);
and U23520 (N_23520,N_19271,N_18796);
xor U23521 (N_23521,N_20907,N_19424);
and U23522 (N_23522,N_18833,N_21274);
nor U23523 (N_23523,N_19037,N_21659);
and U23524 (N_23524,N_20692,N_19460);
nand U23525 (N_23525,N_18853,N_19142);
and U23526 (N_23526,N_21446,N_19713);
and U23527 (N_23527,N_19607,N_21152);
nand U23528 (N_23528,N_20495,N_20758);
and U23529 (N_23529,N_21027,N_21000);
nand U23530 (N_23530,N_21651,N_20376);
and U23531 (N_23531,N_19295,N_19468);
or U23532 (N_23532,N_18868,N_19038);
or U23533 (N_23533,N_18968,N_20719);
and U23534 (N_23534,N_20934,N_18875);
nor U23535 (N_23535,N_19355,N_21354);
xor U23536 (N_23536,N_21359,N_19256);
and U23537 (N_23537,N_19466,N_19512);
nor U23538 (N_23538,N_19485,N_21384);
and U23539 (N_23539,N_19721,N_20085);
xnor U23540 (N_23540,N_18835,N_21516);
and U23541 (N_23541,N_19463,N_21524);
nand U23542 (N_23542,N_19025,N_21582);
and U23543 (N_23543,N_21486,N_20509);
or U23544 (N_23544,N_19751,N_19367);
xor U23545 (N_23545,N_19150,N_21568);
and U23546 (N_23546,N_20832,N_20706);
and U23547 (N_23547,N_21021,N_19836);
or U23548 (N_23548,N_19462,N_21631);
and U23549 (N_23549,N_18750,N_20562);
nand U23550 (N_23550,N_21599,N_19928);
or U23551 (N_23551,N_20342,N_20815);
nand U23552 (N_23552,N_19049,N_19067);
nand U23553 (N_23553,N_18817,N_21469);
nor U23554 (N_23554,N_20912,N_19572);
nand U23555 (N_23555,N_20633,N_21616);
xnor U23556 (N_23556,N_19835,N_21557);
nand U23557 (N_23557,N_19593,N_20976);
and U23558 (N_23558,N_18969,N_21735);
xor U23559 (N_23559,N_19394,N_21737);
nor U23560 (N_23560,N_20380,N_19262);
nor U23561 (N_23561,N_21394,N_20072);
and U23562 (N_23562,N_19420,N_19603);
or U23563 (N_23563,N_19318,N_20259);
or U23564 (N_23564,N_19071,N_18950);
or U23565 (N_23565,N_19139,N_20935);
and U23566 (N_23566,N_21587,N_20007);
and U23567 (N_23567,N_19544,N_19253);
xnor U23568 (N_23568,N_20461,N_21794);
xor U23569 (N_23569,N_20709,N_18817);
and U23570 (N_23570,N_21386,N_21368);
nor U23571 (N_23571,N_19403,N_19593);
nor U23572 (N_23572,N_21512,N_21409);
nand U23573 (N_23573,N_20259,N_20113);
and U23574 (N_23574,N_21840,N_20802);
nand U23575 (N_23575,N_21210,N_19530);
or U23576 (N_23576,N_19811,N_20624);
or U23577 (N_23577,N_20487,N_19173);
or U23578 (N_23578,N_21439,N_19631);
or U23579 (N_23579,N_19958,N_19016);
or U23580 (N_23580,N_18753,N_19580);
or U23581 (N_23581,N_20367,N_20628);
or U23582 (N_23582,N_19792,N_20124);
nor U23583 (N_23583,N_20870,N_19077);
nand U23584 (N_23584,N_21300,N_19575);
nor U23585 (N_23585,N_20720,N_19378);
nand U23586 (N_23586,N_21398,N_19576);
and U23587 (N_23587,N_20835,N_18775);
nor U23588 (N_23588,N_19790,N_21068);
nand U23589 (N_23589,N_20248,N_19008);
nor U23590 (N_23590,N_21487,N_19619);
or U23591 (N_23591,N_20376,N_18895);
nand U23592 (N_23592,N_19466,N_20039);
or U23593 (N_23593,N_19767,N_19460);
xor U23594 (N_23594,N_19230,N_19302);
nor U23595 (N_23595,N_19483,N_20390);
nor U23596 (N_23596,N_21528,N_20546);
or U23597 (N_23597,N_21385,N_21111);
nand U23598 (N_23598,N_21771,N_18985);
nand U23599 (N_23599,N_18930,N_20478);
or U23600 (N_23600,N_19414,N_19747);
nor U23601 (N_23601,N_21088,N_19580);
nor U23602 (N_23602,N_19532,N_21490);
and U23603 (N_23603,N_19820,N_21109);
nand U23604 (N_23604,N_18913,N_21675);
or U23605 (N_23605,N_21824,N_20503);
nand U23606 (N_23606,N_19510,N_19451);
nand U23607 (N_23607,N_21289,N_20197);
and U23608 (N_23608,N_21544,N_19803);
nand U23609 (N_23609,N_21408,N_19293);
or U23610 (N_23610,N_19462,N_21421);
or U23611 (N_23611,N_20162,N_21403);
xor U23612 (N_23612,N_20081,N_19046);
or U23613 (N_23613,N_19287,N_19598);
or U23614 (N_23614,N_21674,N_21069);
and U23615 (N_23615,N_20166,N_21356);
xor U23616 (N_23616,N_21291,N_20958);
or U23617 (N_23617,N_21073,N_20559);
nor U23618 (N_23618,N_20501,N_20277);
nand U23619 (N_23619,N_20785,N_20770);
and U23620 (N_23620,N_21370,N_20772);
nand U23621 (N_23621,N_21782,N_20101);
nand U23622 (N_23622,N_18816,N_21744);
and U23623 (N_23623,N_21856,N_20320);
nor U23624 (N_23624,N_21631,N_20560);
or U23625 (N_23625,N_20867,N_21477);
nand U23626 (N_23626,N_20845,N_21868);
or U23627 (N_23627,N_21006,N_19144);
nor U23628 (N_23628,N_21271,N_20003);
nand U23629 (N_23629,N_20061,N_19022);
and U23630 (N_23630,N_18892,N_19321);
and U23631 (N_23631,N_20914,N_21712);
nor U23632 (N_23632,N_19844,N_19275);
and U23633 (N_23633,N_21334,N_19524);
nand U23634 (N_23634,N_21529,N_20337);
nor U23635 (N_23635,N_21048,N_20472);
xnor U23636 (N_23636,N_21538,N_21176);
nor U23637 (N_23637,N_18913,N_21084);
nand U23638 (N_23638,N_19851,N_18959);
and U23639 (N_23639,N_20928,N_20778);
or U23640 (N_23640,N_19760,N_21480);
nor U23641 (N_23641,N_19815,N_20918);
or U23642 (N_23642,N_21132,N_19960);
or U23643 (N_23643,N_18965,N_19061);
xor U23644 (N_23644,N_21434,N_20788);
nor U23645 (N_23645,N_19996,N_20283);
or U23646 (N_23646,N_20468,N_19269);
and U23647 (N_23647,N_20443,N_19696);
nand U23648 (N_23648,N_21048,N_18824);
nand U23649 (N_23649,N_19581,N_20746);
or U23650 (N_23650,N_21643,N_20444);
or U23651 (N_23651,N_20939,N_18981);
or U23652 (N_23652,N_19274,N_20725);
and U23653 (N_23653,N_19127,N_19886);
or U23654 (N_23654,N_20193,N_21003);
nand U23655 (N_23655,N_18872,N_20179);
nand U23656 (N_23656,N_19480,N_21674);
or U23657 (N_23657,N_20187,N_18982);
or U23658 (N_23658,N_20026,N_20595);
or U23659 (N_23659,N_21491,N_20662);
nand U23660 (N_23660,N_20334,N_21086);
nor U23661 (N_23661,N_20785,N_21453);
nand U23662 (N_23662,N_19247,N_20778);
nor U23663 (N_23663,N_20544,N_21619);
nand U23664 (N_23664,N_21833,N_20554);
and U23665 (N_23665,N_20691,N_19384);
nand U23666 (N_23666,N_20887,N_20251);
xnor U23667 (N_23667,N_21722,N_19603);
nor U23668 (N_23668,N_21160,N_19181);
and U23669 (N_23669,N_20231,N_19751);
nor U23670 (N_23670,N_21734,N_19980);
nor U23671 (N_23671,N_20256,N_21233);
nor U23672 (N_23672,N_20206,N_19647);
xnor U23673 (N_23673,N_21210,N_19650);
nor U23674 (N_23674,N_19745,N_19913);
and U23675 (N_23675,N_21388,N_21387);
xor U23676 (N_23676,N_18950,N_21587);
nand U23677 (N_23677,N_21738,N_20320);
nand U23678 (N_23678,N_21343,N_20521);
nor U23679 (N_23679,N_20957,N_19243);
nand U23680 (N_23680,N_20802,N_20278);
nor U23681 (N_23681,N_21514,N_21687);
and U23682 (N_23682,N_20433,N_20138);
and U23683 (N_23683,N_20129,N_19551);
and U23684 (N_23684,N_21660,N_19487);
or U23685 (N_23685,N_20137,N_21709);
xor U23686 (N_23686,N_19672,N_19065);
xor U23687 (N_23687,N_21579,N_20572);
or U23688 (N_23688,N_20289,N_21068);
nor U23689 (N_23689,N_20650,N_19635);
or U23690 (N_23690,N_19957,N_19541);
nand U23691 (N_23691,N_21769,N_19088);
or U23692 (N_23692,N_20378,N_21741);
nor U23693 (N_23693,N_19576,N_19694);
or U23694 (N_23694,N_19496,N_18848);
or U23695 (N_23695,N_21593,N_21624);
nor U23696 (N_23696,N_21531,N_19452);
or U23697 (N_23697,N_21610,N_21533);
nand U23698 (N_23698,N_19739,N_19489);
and U23699 (N_23699,N_20858,N_20683);
and U23700 (N_23700,N_19453,N_20220);
and U23701 (N_23701,N_20875,N_20076);
or U23702 (N_23702,N_18935,N_20415);
nor U23703 (N_23703,N_19838,N_18998);
and U23704 (N_23704,N_19698,N_21743);
or U23705 (N_23705,N_19248,N_18897);
or U23706 (N_23706,N_20010,N_20460);
or U23707 (N_23707,N_20332,N_19865);
and U23708 (N_23708,N_21573,N_21774);
and U23709 (N_23709,N_20057,N_20945);
nand U23710 (N_23710,N_19786,N_19421);
and U23711 (N_23711,N_21132,N_19378);
nor U23712 (N_23712,N_18784,N_21157);
xnor U23713 (N_23713,N_19493,N_21724);
and U23714 (N_23714,N_20306,N_20111);
xnor U23715 (N_23715,N_20720,N_21224);
or U23716 (N_23716,N_20608,N_18944);
and U23717 (N_23717,N_19537,N_19246);
xnor U23718 (N_23718,N_21693,N_20630);
nor U23719 (N_23719,N_19513,N_19705);
or U23720 (N_23720,N_19558,N_20849);
or U23721 (N_23721,N_19814,N_20045);
nand U23722 (N_23722,N_19186,N_20100);
nor U23723 (N_23723,N_19295,N_20825);
nand U23724 (N_23724,N_19085,N_20764);
and U23725 (N_23725,N_21761,N_20271);
xnor U23726 (N_23726,N_20157,N_18943);
nand U23727 (N_23727,N_19676,N_21384);
nor U23728 (N_23728,N_19452,N_18977);
or U23729 (N_23729,N_19050,N_21151);
or U23730 (N_23730,N_20304,N_19058);
or U23731 (N_23731,N_21324,N_19927);
nor U23732 (N_23732,N_19954,N_19023);
nand U23733 (N_23733,N_20067,N_20790);
xor U23734 (N_23734,N_19986,N_19399);
and U23735 (N_23735,N_18976,N_21617);
and U23736 (N_23736,N_21105,N_21708);
or U23737 (N_23737,N_19733,N_21337);
nor U23738 (N_23738,N_20706,N_21359);
nand U23739 (N_23739,N_20287,N_20321);
nand U23740 (N_23740,N_20214,N_19062);
xor U23741 (N_23741,N_20244,N_19517);
nand U23742 (N_23742,N_19515,N_20883);
nor U23743 (N_23743,N_19363,N_19300);
nor U23744 (N_23744,N_18887,N_21198);
nand U23745 (N_23745,N_20487,N_18847);
and U23746 (N_23746,N_21196,N_20849);
nor U23747 (N_23747,N_19656,N_19617);
nor U23748 (N_23748,N_21606,N_21256);
nor U23749 (N_23749,N_21831,N_19724);
or U23750 (N_23750,N_21254,N_20356);
xor U23751 (N_23751,N_21032,N_19045);
xor U23752 (N_23752,N_21771,N_20417);
and U23753 (N_23753,N_20047,N_18997);
xor U23754 (N_23754,N_20144,N_20889);
xnor U23755 (N_23755,N_20001,N_21598);
or U23756 (N_23756,N_20368,N_20851);
and U23757 (N_23757,N_20844,N_21109);
nand U23758 (N_23758,N_20212,N_21125);
nand U23759 (N_23759,N_20619,N_21617);
nor U23760 (N_23760,N_21440,N_20974);
or U23761 (N_23761,N_20496,N_20593);
nor U23762 (N_23762,N_19211,N_19353);
nand U23763 (N_23763,N_19803,N_21215);
nor U23764 (N_23764,N_18770,N_21790);
and U23765 (N_23765,N_20659,N_20292);
nand U23766 (N_23766,N_20802,N_21288);
xnor U23767 (N_23767,N_20356,N_20392);
and U23768 (N_23768,N_20902,N_21523);
or U23769 (N_23769,N_21326,N_20854);
or U23770 (N_23770,N_21702,N_21369);
nand U23771 (N_23771,N_19562,N_21712);
xor U23772 (N_23772,N_20023,N_21361);
and U23773 (N_23773,N_19646,N_18763);
and U23774 (N_23774,N_21098,N_21241);
nor U23775 (N_23775,N_21770,N_21381);
nand U23776 (N_23776,N_19216,N_20115);
and U23777 (N_23777,N_21132,N_19537);
and U23778 (N_23778,N_19963,N_20642);
nor U23779 (N_23779,N_19593,N_20141);
nand U23780 (N_23780,N_18765,N_20519);
nand U23781 (N_23781,N_18801,N_21660);
nand U23782 (N_23782,N_21008,N_21646);
or U23783 (N_23783,N_20352,N_18814);
nor U23784 (N_23784,N_19713,N_18864);
and U23785 (N_23785,N_19489,N_20165);
xor U23786 (N_23786,N_19540,N_19734);
or U23787 (N_23787,N_21781,N_21815);
or U23788 (N_23788,N_21069,N_19896);
or U23789 (N_23789,N_21001,N_19327);
or U23790 (N_23790,N_21436,N_21643);
and U23791 (N_23791,N_20253,N_19567);
nand U23792 (N_23792,N_20151,N_20556);
nand U23793 (N_23793,N_20615,N_20917);
and U23794 (N_23794,N_18869,N_20331);
and U23795 (N_23795,N_19332,N_21872);
nor U23796 (N_23796,N_21720,N_20186);
nand U23797 (N_23797,N_19491,N_20873);
xor U23798 (N_23798,N_21074,N_19363);
nand U23799 (N_23799,N_21415,N_19463);
or U23800 (N_23800,N_19866,N_20622);
or U23801 (N_23801,N_19693,N_20046);
nor U23802 (N_23802,N_20148,N_20713);
nand U23803 (N_23803,N_20491,N_20621);
or U23804 (N_23804,N_19776,N_21782);
and U23805 (N_23805,N_20594,N_20860);
and U23806 (N_23806,N_21137,N_19293);
nor U23807 (N_23807,N_21445,N_19805);
and U23808 (N_23808,N_19566,N_21330);
nor U23809 (N_23809,N_20003,N_21860);
or U23810 (N_23810,N_21038,N_20313);
and U23811 (N_23811,N_19695,N_19823);
and U23812 (N_23812,N_20060,N_19713);
nand U23813 (N_23813,N_20746,N_20229);
nor U23814 (N_23814,N_21432,N_18942);
or U23815 (N_23815,N_20064,N_19759);
and U23816 (N_23816,N_18857,N_19325);
or U23817 (N_23817,N_21241,N_21439);
nor U23818 (N_23818,N_21019,N_19666);
and U23819 (N_23819,N_20436,N_20990);
nand U23820 (N_23820,N_20962,N_20833);
xnor U23821 (N_23821,N_18887,N_20938);
nand U23822 (N_23822,N_21232,N_19867);
or U23823 (N_23823,N_18993,N_20521);
or U23824 (N_23824,N_20936,N_21104);
and U23825 (N_23825,N_21635,N_21741);
or U23826 (N_23826,N_21848,N_21338);
and U23827 (N_23827,N_21569,N_21431);
or U23828 (N_23828,N_19293,N_19988);
or U23829 (N_23829,N_20928,N_18929);
xor U23830 (N_23830,N_19166,N_20765);
nor U23831 (N_23831,N_20113,N_19961);
nand U23832 (N_23832,N_18988,N_18944);
or U23833 (N_23833,N_18941,N_19843);
and U23834 (N_23834,N_20901,N_21639);
nor U23835 (N_23835,N_18950,N_20250);
nor U23836 (N_23836,N_20355,N_21815);
nand U23837 (N_23837,N_20233,N_19583);
nand U23838 (N_23838,N_18852,N_18949);
xnor U23839 (N_23839,N_20670,N_21661);
and U23840 (N_23840,N_21408,N_20352);
or U23841 (N_23841,N_19632,N_19320);
nand U23842 (N_23842,N_20989,N_19493);
nor U23843 (N_23843,N_20135,N_21726);
and U23844 (N_23844,N_19882,N_18831);
or U23845 (N_23845,N_21633,N_21693);
nor U23846 (N_23846,N_19957,N_19261);
nand U23847 (N_23847,N_21670,N_19841);
or U23848 (N_23848,N_21492,N_21657);
xnor U23849 (N_23849,N_20702,N_19982);
and U23850 (N_23850,N_19320,N_19197);
nor U23851 (N_23851,N_21365,N_19319);
and U23852 (N_23852,N_19337,N_18938);
nor U23853 (N_23853,N_20419,N_20181);
nor U23854 (N_23854,N_19212,N_18916);
nor U23855 (N_23855,N_21596,N_21178);
xor U23856 (N_23856,N_18857,N_20585);
xor U23857 (N_23857,N_21869,N_20745);
nand U23858 (N_23858,N_18923,N_21216);
nand U23859 (N_23859,N_20148,N_21574);
nand U23860 (N_23860,N_18950,N_20891);
nor U23861 (N_23861,N_19691,N_19926);
xnor U23862 (N_23862,N_19246,N_20089);
nand U23863 (N_23863,N_20618,N_20187);
nand U23864 (N_23864,N_19127,N_20790);
and U23865 (N_23865,N_20885,N_19748);
or U23866 (N_23866,N_18779,N_19750);
or U23867 (N_23867,N_20273,N_21434);
nand U23868 (N_23868,N_21375,N_20018);
nand U23869 (N_23869,N_19092,N_18972);
nand U23870 (N_23870,N_20599,N_21840);
xor U23871 (N_23871,N_21478,N_19507);
nand U23872 (N_23872,N_19528,N_20841);
xor U23873 (N_23873,N_19322,N_21132);
and U23874 (N_23874,N_20471,N_19317);
or U23875 (N_23875,N_21075,N_20988);
nand U23876 (N_23876,N_20001,N_20648);
and U23877 (N_23877,N_19101,N_20675);
nor U23878 (N_23878,N_19067,N_21856);
and U23879 (N_23879,N_19257,N_20585);
nor U23880 (N_23880,N_21843,N_21811);
nand U23881 (N_23881,N_19129,N_21852);
or U23882 (N_23882,N_19023,N_19081);
nand U23883 (N_23883,N_19174,N_21649);
nand U23884 (N_23884,N_19089,N_20605);
or U23885 (N_23885,N_19806,N_20452);
or U23886 (N_23886,N_21724,N_19451);
or U23887 (N_23887,N_21551,N_20689);
and U23888 (N_23888,N_20169,N_20456);
and U23889 (N_23889,N_20547,N_20135);
and U23890 (N_23890,N_19912,N_20874);
or U23891 (N_23891,N_19469,N_19394);
nand U23892 (N_23892,N_19132,N_21318);
or U23893 (N_23893,N_18864,N_19730);
and U23894 (N_23894,N_21250,N_19145);
nand U23895 (N_23895,N_21765,N_19446);
nand U23896 (N_23896,N_20015,N_21377);
nand U23897 (N_23897,N_21733,N_19844);
xnor U23898 (N_23898,N_20603,N_20994);
nand U23899 (N_23899,N_21383,N_21100);
nand U23900 (N_23900,N_21563,N_20060);
nand U23901 (N_23901,N_20181,N_19499);
nand U23902 (N_23902,N_21688,N_20045);
nor U23903 (N_23903,N_20750,N_20300);
or U23904 (N_23904,N_19437,N_19122);
xor U23905 (N_23905,N_20281,N_19549);
or U23906 (N_23906,N_20655,N_18781);
or U23907 (N_23907,N_21381,N_21160);
nand U23908 (N_23908,N_20276,N_19009);
or U23909 (N_23909,N_20571,N_19065);
or U23910 (N_23910,N_20556,N_21102);
xnor U23911 (N_23911,N_19067,N_19042);
nor U23912 (N_23912,N_21689,N_18809);
or U23913 (N_23913,N_20393,N_21856);
or U23914 (N_23914,N_20361,N_19902);
nand U23915 (N_23915,N_20216,N_19936);
or U23916 (N_23916,N_19620,N_19453);
or U23917 (N_23917,N_20182,N_19128);
nand U23918 (N_23918,N_18806,N_19891);
nand U23919 (N_23919,N_19297,N_19470);
nand U23920 (N_23920,N_18776,N_20704);
nor U23921 (N_23921,N_20367,N_21199);
nor U23922 (N_23922,N_21343,N_18876);
or U23923 (N_23923,N_20014,N_21423);
xor U23924 (N_23924,N_20247,N_20202);
and U23925 (N_23925,N_19478,N_19747);
nand U23926 (N_23926,N_19643,N_21081);
and U23927 (N_23927,N_19503,N_21380);
xnor U23928 (N_23928,N_21691,N_19764);
or U23929 (N_23929,N_21162,N_18956);
or U23930 (N_23930,N_21495,N_21337);
or U23931 (N_23931,N_18751,N_19313);
nor U23932 (N_23932,N_21542,N_19769);
nand U23933 (N_23933,N_21450,N_20161);
nand U23934 (N_23934,N_20058,N_21486);
nor U23935 (N_23935,N_20669,N_19990);
nor U23936 (N_23936,N_19853,N_21688);
nand U23937 (N_23937,N_21544,N_20194);
or U23938 (N_23938,N_20663,N_21759);
and U23939 (N_23939,N_19665,N_18910);
nor U23940 (N_23940,N_20894,N_18886);
nor U23941 (N_23941,N_19760,N_18926);
and U23942 (N_23942,N_20415,N_21595);
nand U23943 (N_23943,N_20149,N_21366);
nor U23944 (N_23944,N_19088,N_19371);
and U23945 (N_23945,N_21128,N_21375);
nand U23946 (N_23946,N_19005,N_21740);
nand U23947 (N_23947,N_20970,N_21032);
or U23948 (N_23948,N_19350,N_20190);
and U23949 (N_23949,N_18934,N_21487);
nor U23950 (N_23950,N_19462,N_20188);
nor U23951 (N_23951,N_20641,N_19379);
and U23952 (N_23952,N_21174,N_19227);
nor U23953 (N_23953,N_20508,N_20176);
nor U23954 (N_23954,N_21242,N_19300);
or U23955 (N_23955,N_21375,N_18958);
nor U23956 (N_23956,N_21383,N_21812);
and U23957 (N_23957,N_21739,N_20225);
and U23958 (N_23958,N_19193,N_20773);
nand U23959 (N_23959,N_21334,N_18862);
or U23960 (N_23960,N_20150,N_20137);
or U23961 (N_23961,N_20374,N_19806);
and U23962 (N_23962,N_19370,N_20088);
and U23963 (N_23963,N_21868,N_21125);
nor U23964 (N_23964,N_20784,N_19332);
nand U23965 (N_23965,N_20108,N_19861);
or U23966 (N_23966,N_20712,N_21426);
or U23967 (N_23967,N_19586,N_19837);
and U23968 (N_23968,N_21605,N_21592);
and U23969 (N_23969,N_20832,N_20491);
or U23970 (N_23970,N_20185,N_20029);
or U23971 (N_23971,N_19959,N_21659);
nand U23972 (N_23972,N_19892,N_20049);
nor U23973 (N_23973,N_19501,N_19673);
or U23974 (N_23974,N_21378,N_19520);
and U23975 (N_23975,N_21228,N_20634);
xor U23976 (N_23976,N_19349,N_19189);
or U23977 (N_23977,N_19693,N_20173);
nand U23978 (N_23978,N_18974,N_20430);
or U23979 (N_23979,N_19586,N_20883);
and U23980 (N_23980,N_21474,N_21081);
or U23981 (N_23981,N_20114,N_19549);
and U23982 (N_23982,N_18868,N_20872);
nor U23983 (N_23983,N_19178,N_19410);
and U23984 (N_23984,N_21167,N_19108);
or U23985 (N_23985,N_21239,N_19722);
nor U23986 (N_23986,N_21829,N_19101);
or U23987 (N_23987,N_19712,N_20227);
or U23988 (N_23988,N_19923,N_21118);
nor U23989 (N_23989,N_19800,N_19132);
nor U23990 (N_23990,N_19841,N_19409);
nor U23991 (N_23991,N_21448,N_21166);
nor U23992 (N_23992,N_20545,N_19765);
nor U23993 (N_23993,N_19140,N_21775);
nand U23994 (N_23994,N_20255,N_20865);
nand U23995 (N_23995,N_19811,N_19901);
nor U23996 (N_23996,N_20896,N_21843);
or U23997 (N_23997,N_19383,N_18944);
nor U23998 (N_23998,N_19533,N_19993);
or U23999 (N_23999,N_20219,N_20346);
xnor U24000 (N_24000,N_20396,N_21226);
xnor U24001 (N_24001,N_21562,N_20801);
nand U24002 (N_24002,N_19645,N_20111);
nor U24003 (N_24003,N_19102,N_19380);
or U24004 (N_24004,N_19639,N_19048);
and U24005 (N_24005,N_21304,N_21028);
nand U24006 (N_24006,N_20109,N_20172);
nand U24007 (N_24007,N_19396,N_21083);
nor U24008 (N_24008,N_21711,N_20881);
or U24009 (N_24009,N_21322,N_20965);
nor U24010 (N_24010,N_18848,N_20510);
or U24011 (N_24011,N_21532,N_19872);
nand U24012 (N_24012,N_21408,N_19725);
nor U24013 (N_24013,N_20533,N_19626);
or U24014 (N_24014,N_21411,N_21598);
nor U24015 (N_24015,N_19489,N_20019);
nor U24016 (N_24016,N_20751,N_19223);
or U24017 (N_24017,N_20938,N_19176);
or U24018 (N_24018,N_19611,N_21831);
and U24019 (N_24019,N_18826,N_21597);
nand U24020 (N_24020,N_20397,N_21799);
nor U24021 (N_24021,N_20784,N_19417);
nor U24022 (N_24022,N_20358,N_19883);
and U24023 (N_24023,N_20433,N_21631);
nor U24024 (N_24024,N_20745,N_19383);
or U24025 (N_24025,N_20158,N_18929);
nand U24026 (N_24026,N_19565,N_20520);
nor U24027 (N_24027,N_20206,N_21144);
xnor U24028 (N_24028,N_20575,N_21448);
and U24029 (N_24029,N_21157,N_20245);
nand U24030 (N_24030,N_19601,N_19804);
or U24031 (N_24031,N_19546,N_19986);
or U24032 (N_24032,N_20865,N_21237);
and U24033 (N_24033,N_21827,N_20347);
xnor U24034 (N_24034,N_19936,N_19663);
nand U24035 (N_24035,N_20939,N_18969);
nand U24036 (N_24036,N_20757,N_19326);
and U24037 (N_24037,N_19408,N_20427);
nor U24038 (N_24038,N_20942,N_20814);
nor U24039 (N_24039,N_20495,N_21427);
xnor U24040 (N_24040,N_21701,N_20618);
or U24041 (N_24041,N_20562,N_21175);
nor U24042 (N_24042,N_20697,N_21150);
nor U24043 (N_24043,N_20391,N_21019);
nor U24044 (N_24044,N_21724,N_20852);
and U24045 (N_24045,N_19032,N_21761);
nor U24046 (N_24046,N_20912,N_19643);
xnor U24047 (N_24047,N_21011,N_19428);
nand U24048 (N_24048,N_19866,N_18934);
nand U24049 (N_24049,N_19802,N_21175);
xor U24050 (N_24050,N_20354,N_19244);
or U24051 (N_24051,N_21229,N_21646);
nor U24052 (N_24052,N_21442,N_20861);
or U24053 (N_24053,N_21710,N_21212);
or U24054 (N_24054,N_19294,N_19953);
and U24055 (N_24055,N_20950,N_20544);
or U24056 (N_24056,N_20718,N_21845);
nand U24057 (N_24057,N_21852,N_21129);
and U24058 (N_24058,N_20936,N_19216);
nand U24059 (N_24059,N_19002,N_21466);
nor U24060 (N_24060,N_21130,N_21652);
and U24061 (N_24061,N_18857,N_18782);
xor U24062 (N_24062,N_19604,N_19450);
or U24063 (N_24063,N_21434,N_20235);
nand U24064 (N_24064,N_20684,N_21342);
and U24065 (N_24065,N_19565,N_21553);
or U24066 (N_24066,N_20771,N_21299);
and U24067 (N_24067,N_21484,N_19733);
or U24068 (N_24068,N_19213,N_21019);
or U24069 (N_24069,N_20371,N_20059);
nand U24070 (N_24070,N_20887,N_21739);
nor U24071 (N_24071,N_20984,N_18930);
xor U24072 (N_24072,N_19876,N_21449);
nor U24073 (N_24073,N_21562,N_19999);
and U24074 (N_24074,N_20914,N_20604);
and U24075 (N_24075,N_21772,N_20083);
xor U24076 (N_24076,N_20352,N_19686);
nand U24077 (N_24077,N_19660,N_19500);
xnor U24078 (N_24078,N_19931,N_20846);
xnor U24079 (N_24079,N_21104,N_18946);
or U24080 (N_24080,N_20351,N_19088);
xor U24081 (N_24081,N_20271,N_18945);
and U24082 (N_24082,N_20109,N_18888);
xor U24083 (N_24083,N_19615,N_21559);
and U24084 (N_24084,N_21020,N_21449);
nor U24085 (N_24085,N_19512,N_20581);
nand U24086 (N_24086,N_20045,N_21558);
or U24087 (N_24087,N_19740,N_19237);
or U24088 (N_24088,N_21091,N_20058);
nand U24089 (N_24089,N_21796,N_19479);
nand U24090 (N_24090,N_20826,N_21793);
and U24091 (N_24091,N_21649,N_18822);
and U24092 (N_24092,N_21170,N_21177);
or U24093 (N_24093,N_21740,N_19552);
xor U24094 (N_24094,N_21673,N_20996);
nand U24095 (N_24095,N_19352,N_20447);
and U24096 (N_24096,N_19730,N_18898);
and U24097 (N_24097,N_21749,N_21357);
xnor U24098 (N_24098,N_18993,N_20977);
nand U24099 (N_24099,N_20709,N_20186);
nand U24100 (N_24100,N_20248,N_20923);
nor U24101 (N_24101,N_20464,N_20889);
xor U24102 (N_24102,N_20251,N_21091);
and U24103 (N_24103,N_21728,N_20428);
nand U24104 (N_24104,N_19893,N_20706);
and U24105 (N_24105,N_20726,N_20607);
nand U24106 (N_24106,N_18968,N_21434);
nand U24107 (N_24107,N_19483,N_19186);
nor U24108 (N_24108,N_19732,N_20104);
nand U24109 (N_24109,N_19623,N_18899);
and U24110 (N_24110,N_19268,N_19752);
or U24111 (N_24111,N_18904,N_18860);
nand U24112 (N_24112,N_20372,N_21305);
or U24113 (N_24113,N_20850,N_19778);
or U24114 (N_24114,N_20565,N_21533);
nor U24115 (N_24115,N_18810,N_20879);
nand U24116 (N_24116,N_19817,N_20746);
or U24117 (N_24117,N_20456,N_20010);
nor U24118 (N_24118,N_19752,N_21565);
or U24119 (N_24119,N_19197,N_19034);
nor U24120 (N_24120,N_19517,N_19501);
and U24121 (N_24121,N_21422,N_19380);
or U24122 (N_24122,N_19340,N_21135);
nor U24123 (N_24123,N_20276,N_21229);
or U24124 (N_24124,N_20136,N_21623);
or U24125 (N_24125,N_20498,N_18868);
or U24126 (N_24126,N_21824,N_19226);
xor U24127 (N_24127,N_19000,N_21781);
and U24128 (N_24128,N_21102,N_19759);
or U24129 (N_24129,N_20720,N_20166);
nand U24130 (N_24130,N_19978,N_19850);
nand U24131 (N_24131,N_18785,N_20803);
and U24132 (N_24132,N_21566,N_21580);
nor U24133 (N_24133,N_20758,N_19259);
and U24134 (N_24134,N_20618,N_19343);
or U24135 (N_24135,N_21660,N_20525);
nor U24136 (N_24136,N_21553,N_19081);
or U24137 (N_24137,N_19160,N_18831);
or U24138 (N_24138,N_18758,N_21359);
xor U24139 (N_24139,N_21377,N_20488);
nand U24140 (N_24140,N_19705,N_20318);
xor U24141 (N_24141,N_21671,N_20741);
nor U24142 (N_24142,N_21276,N_20019);
nand U24143 (N_24143,N_21341,N_20767);
xnor U24144 (N_24144,N_19063,N_19214);
and U24145 (N_24145,N_20850,N_21702);
xnor U24146 (N_24146,N_19947,N_20282);
and U24147 (N_24147,N_21262,N_20501);
or U24148 (N_24148,N_20599,N_19630);
and U24149 (N_24149,N_21593,N_20842);
nor U24150 (N_24150,N_20512,N_19443);
or U24151 (N_24151,N_19767,N_20694);
nor U24152 (N_24152,N_20600,N_20193);
nor U24153 (N_24153,N_18936,N_21001);
nand U24154 (N_24154,N_19739,N_21074);
nand U24155 (N_24155,N_20673,N_19652);
nor U24156 (N_24156,N_19197,N_19264);
nand U24157 (N_24157,N_21562,N_20926);
xnor U24158 (N_24158,N_19141,N_21531);
xnor U24159 (N_24159,N_21063,N_19766);
xor U24160 (N_24160,N_20606,N_21291);
nand U24161 (N_24161,N_20135,N_19211);
nand U24162 (N_24162,N_19384,N_21631);
and U24163 (N_24163,N_20937,N_19254);
xnor U24164 (N_24164,N_19967,N_19331);
nand U24165 (N_24165,N_20816,N_20136);
nor U24166 (N_24166,N_20121,N_21783);
and U24167 (N_24167,N_19968,N_19872);
nor U24168 (N_24168,N_18851,N_19560);
and U24169 (N_24169,N_21440,N_19543);
nor U24170 (N_24170,N_21806,N_20849);
or U24171 (N_24171,N_18763,N_19756);
nor U24172 (N_24172,N_19137,N_18977);
nor U24173 (N_24173,N_21269,N_19763);
xor U24174 (N_24174,N_21539,N_21532);
and U24175 (N_24175,N_19724,N_21338);
nor U24176 (N_24176,N_20887,N_21137);
and U24177 (N_24177,N_19932,N_21251);
or U24178 (N_24178,N_18823,N_21387);
xnor U24179 (N_24179,N_20940,N_20409);
nor U24180 (N_24180,N_20242,N_20903);
or U24181 (N_24181,N_21641,N_19889);
nor U24182 (N_24182,N_20325,N_21371);
nand U24183 (N_24183,N_20269,N_20372);
nand U24184 (N_24184,N_20724,N_20885);
or U24185 (N_24185,N_20893,N_19478);
or U24186 (N_24186,N_21506,N_18890);
and U24187 (N_24187,N_19218,N_20271);
nand U24188 (N_24188,N_20466,N_21114);
nand U24189 (N_24189,N_18840,N_19051);
or U24190 (N_24190,N_20601,N_21170);
and U24191 (N_24191,N_20176,N_19629);
nor U24192 (N_24192,N_20299,N_19053);
nor U24193 (N_24193,N_19644,N_19642);
nor U24194 (N_24194,N_19429,N_20167);
nor U24195 (N_24195,N_20439,N_21838);
and U24196 (N_24196,N_20176,N_19057);
nor U24197 (N_24197,N_21075,N_19740);
nand U24198 (N_24198,N_21371,N_21380);
nor U24199 (N_24199,N_20873,N_19328);
nor U24200 (N_24200,N_21379,N_21548);
nand U24201 (N_24201,N_19399,N_20024);
xor U24202 (N_24202,N_19454,N_18752);
and U24203 (N_24203,N_20790,N_20958);
nor U24204 (N_24204,N_19564,N_19902);
nand U24205 (N_24205,N_20797,N_20017);
or U24206 (N_24206,N_18976,N_19256);
nand U24207 (N_24207,N_19245,N_21557);
or U24208 (N_24208,N_19091,N_19774);
nand U24209 (N_24209,N_19422,N_20775);
nand U24210 (N_24210,N_21167,N_20426);
or U24211 (N_24211,N_19696,N_21078);
nor U24212 (N_24212,N_20249,N_21045);
and U24213 (N_24213,N_19720,N_20598);
nor U24214 (N_24214,N_20087,N_18905);
and U24215 (N_24215,N_18842,N_19344);
nor U24216 (N_24216,N_21657,N_21195);
nand U24217 (N_24217,N_19128,N_19368);
nor U24218 (N_24218,N_20768,N_20663);
nor U24219 (N_24219,N_19720,N_21672);
nor U24220 (N_24220,N_20895,N_21670);
and U24221 (N_24221,N_18944,N_18819);
nor U24222 (N_24222,N_21567,N_21091);
nand U24223 (N_24223,N_21252,N_19364);
nand U24224 (N_24224,N_19137,N_20831);
nand U24225 (N_24225,N_18750,N_18956);
or U24226 (N_24226,N_19714,N_20170);
nand U24227 (N_24227,N_21262,N_20605);
nand U24228 (N_24228,N_20044,N_19423);
or U24229 (N_24229,N_19733,N_19667);
nor U24230 (N_24230,N_18927,N_21171);
and U24231 (N_24231,N_20396,N_18811);
or U24232 (N_24232,N_19078,N_20178);
or U24233 (N_24233,N_19325,N_21739);
and U24234 (N_24234,N_19890,N_21468);
nor U24235 (N_24235,N_21717,N_21038);
and U24236 (N_24236,N_19898,N_20377);
nand U24237 (N_24237,N_19980,N_21586);
nand U24238 (N_24238,N_19197,N_21551);
nand U24239 (N_24239,N_19680,N_19383);
nand U24240 (N_24240,N_21355,N_20987);
and U24241 (N_24241,N_19510,N_20903);
and U24242 (N_24242,N_21216,N_21596);
nand U24243 (N_24243,N_20136,N_20754);
nor U24244 (N_24244,N_20101,N_21134);
xnor U24245 (N_24245,N_20792,N_19643);
or U24246 (N_24246,N_21042,N_20258);
nand U24247 (N_24247,N_18892,N_20537);
nor U24248 (N_24248,N_19766,N_20823);
xnor U24249 (N_24249,N_20354,N_21823);
xnor U24250 (N_24250,N_21761,N_20905);
nor U24251 (N_24251,N_21081,N_21197);
nand U24252 (N_24252,N_20920,N_19665);
nor U24253 (N_24253,N_21098,N_21340);
xor U24254 (N_24254,N_19680,N_20566);
or U24255 (N_24255,N_21833,N_20431);
nand U24256 (N_24256,N_20195,N_21505);
or U24257 (N_24257,N_19823,N_21731);
and U24258 (N_24258,N_21602,N_19133);
nor U24259 (N_24259,N_21143,N_21004);
xor U24260 (N_24260,N_21335,N_20587);
or U24261 (N_24261,N_21582,N_20121);
nor U24262 (N_24262,N_19366,N_18774);
and U24263 (N_24263,N_21304,N_20776);
or U24264 (N_24264,N_20659,N_21239);
and U24265 (N_24265,N_18936,N_20588);
nand U24266 (N_24266,N_18750,N_18786);
nor U24267 (N_24267,N_20865,N_20775);
nand U24268 (N_24268,N_19675,N_20659);
or U24269 (N_24269,N_21647,N_21517);
nand U24270 (N_24270,N_21838,N_20654);
or U24271 (N_24271,N_20058,N_19572);
nand U24272 (N_24272,N_21098,N_21257);
nor U24273 (N_24273,N_20815,N_21067);
or U24274 (N_24274,N_21604,N_21805);
and U24275 (N_24275,N_21787,N_19436);
or U24276 (N_24276,N_21177,N_21795);
or U24277 (N_24277,N_20208,N_20532);
nor U24278 (N_24278,N_21137,N_20051);
nor U24279 (N_24279,N_20068,N_19609);
nand U24280 (N_24280,N_18865,N_19289);
xor U24281 (N_24281,N_18879,N_19792);
or U24282 (N_24282,N_21586,N_21419);
or U24283 (N_24283,N_19754,N_19168);
nor U24284 (N_24284,N_20438,N_19274);
and U24285 (N_24285,N_19454,N_21695);
or U24286 (N_24286,N_19036,N_20969);
or U24287 (N_24287,N_20431,N_19299);
or U24288 (N_24288,N_21753,N_20099);
nand U24289 (N_24289,N_21555,N_19094);
and U24290 (N_24290,N_20511,N_21588);
nor U24291 (N_24291,N_19035,N_20409);
or U24292 (N_24292,N_20925,N_19896);
nor U24293 (N_24293,N_19914,N_19157);
and U24294 (N_24294,N_19010,N_18980);
nor U24295 (N_24295,N_19229,N_21700);
xnor U24296 (N_24296,N_21536,N_21047);
and U24297 (N_24297,N_19878,N_20194);
nand U24298 (N_24298,N_20553,N_21585);
nand U24299 (N_24299,N_19463,N_20207);
or U24300 (N_24300,N_21053,N_20511);
nor U24301 (N_24301,N_20831,N_21799);
nand U24302 (N_24302,N_20790,N_20883);
or U24303 (N_24303,N_19167,N_20170);
and U24304 (N_24304,N_20115,N_20939);
and U24305 (N_24305,N_19398,N_19727);
xor U24306 (N_24306,N_19752,N_19082);
xor U24307 (N_24307,N_19860,N_19845);
nand U24308 (N_24308,N_21767,N_19888);
and U24309 (N_24309,N_19207,N_20771);
and U24310 (N_24310,N_21155,N_19259);
xor U24311 (N_24311,N_19982,N_19306);
xnor U24312 (N_24312,N_18901,N_21533);
xnor U24313 (N_24313,N_21716,N_19269);
nand U24314 (N_24314,N_19290,N_21616);
or U24315 (N_24315,N_18892,N_19939);
and U24316 (N_24316,N_21815,N_21311);
nor U24317 (N_24317,N_21831,N_19900);
or U24318 (N_24318,N_18973,N_21794);
nor U24319 (N_24319,N_19575,N_20703);
xor U24320 (N_24320,N_21283,N_19360);
or U24321 (N_24321,N_21676,N_20824);
and U24322 (N_24322,N_21341,N_20604);
or U24323 (N_24323,N_19917,N_19107);
or U24324 (N_24324,N_20669,N_20606);
and U24325 (N_24325,N_19757,N_21630);
and U24326 (N_24326,N_18941,N_21701);
and U24327 (N_24327,N_19767,N_19694);
or U24328 (N_24328,N_21324,N_21546);
xor U24329 (N_24329,N_21235,N_21522);
nor U24330 (N_24330,N_20734,N_19933);
nand U24331 (N_24331,N_20889,N_19833);
xor U24332 (N_24332,N_19123,N_18854);
nand U24333 (N_24333,N_19386,N_18845);
and U24334 (N_24334,N_21359,N_18992);
and U24335 (N_24335,N_18765,N_19871);
and U24336 (N_24336,N_21486,N_21102);
xnor U24337 (N_24337,N_19340,N_21453);
nand U24338 (N_24338,N_19208,N_21045);
nand U24339 (N_24339,N_21491,N_18970);
nor U24340 (N_24340,N_20605,N_20366);
nor U24341 (N_24341,N_20435,N_20780);
nor U24342 (N_24342,N_20692,N_20121);
nand U24343 (N_24343,N_20631,N_19627);
and U24344 (N_24344,N_20986,N_20644);
or U24345 (N_24345,N_19751,N_19932);
nor U24346 (N_24346,N_20220,N_21394);
nor U24347 (N_24347,N_19872,N_19673);
and U24348 (N_24348,N_20252,N_19533);
or U24349 (N_24349,N_21347,N_20096);
nand U24350 (N_24350,N_19406,N_20285);
nand U24351 (N_24351,N_21721,N_20840);
nand U24352 (N_24352,N_21404,N_19662);
nand U24353 (N_24353,N_21304,N_21776);
nor U24354 (N_24354,N_21434,N_20685);
nand U24355 (N_24355,N_21577,N_21670);
or U24356 (N_24356,N_21279,N_21249);
and U24357 (N_24357,N_20340,N_19808);
nor U24358 (N_24358,N_21251,N_21650);
or U24359 (N_24359,N_21728,N_20213);
nor U24360 (N_24360,N_21276,N_20900);
and U24361 (N_24361,N_19757,N_21499);
and U24362 (N_24362,N_19628,N_19987);
or U24363 (N_24363,N_20969,N_20308);
or U24364 (N_24364,N_20268,N_19720);
nand U24365 (N_24365,N_18964,N_21576);
and U24366 (N_24366,N_20312,N_21248);
and U24367 (N_24367,N_21603,N_20727);
xor U24368 (N_24368,N_20615,N_21154);
nand U24369 (N_24369,N_20845,N_21608);
nor U24370 (N_24370,N_21714,N_20761);
or U24371 (N_24371,N_21482,N_21744);
or U24372 (N_24372,N_20264,N_21338);
nand U24373 (N_24373,N_20417,N_19203);
nand U24374 (N_24374,N_19829,N_19170);
or U24375 (N_24375,N_18822,N_20680);
nor U24376 (N_24376,N_19293,N_21010);
nand U24377 (N_24377,N_21767,N_19399);
nor U24378 (N_24378,N_20819,N_19137);
or U24379 (N_24379,N_21500,N_19564);
and U24380 (N_24380,N_21382,N_19371);
and U24381 (N_24381,N_19546,N_20774);
nand U24382 (N_24382,N_19019,N_21637);
xnor U24383 (N_24383,N_19874,N_21223);
and U24384 (N_24384,N_19545,N_20674);
nand U24385 (N_24385,N_21119,N_20916);
nor U24386 (N_24386,N_20302,N_21316);
nor U24387 (N_24387,N_20835,N_18834);
and U24388 (N_24388,N_21343,N_20378);
nor U24389 (N_24389,N_20774,N_21196);
and U24390 (N_24390,N_21459,N_21153);
and U24391 (N_24391,N_21095,N_19855);
and U24392 (N_24392,N_20058,N_18879);
nor U24393 (N_24393,N_18779,N_19027);
nand U24394 (N_24394,N_21848,N_20187);
and U24395 (N_24395,N_21746,N_20083);
or U24396 (N_24396,N_19498,N_20836);
nand U24397 (N_24397,N_20554,N_19807);
and U24398 (N_24398,N_21148,N_18816);
and U24399 (N_24399,N_20074,N_20407);
or U24400 (N_24400,N_21307,N_19490);
or U24401 (N_24401,N_20652,N_19129);
nand U24402 (N_24402,N_19895,N_21044);
nor U24403 (N_24403,N_18984,N_20777);
or U24404 (N_24404,N_21025,N_19451);
nand U24405 (N_24405,N_20620,N_21356);
nand U24406 (N_24406,N_18988,N_20392);
and U24407 (N_24407,N_19089,N_20215);
nand U24408 (N_24408,N_20398,N_20086);
nand U24409 (N_24409,N_19837,N_19372);
and U24410 (N_24410,N_20633,N_21278);
and U24411 (N_24411,N_19633,N_21483);
nand U24412 (N_24412,N_20438,N_21644);
xnor U24413 (N_24413,N_21335,N_20334);
nor U24414 (N_24414,N_19789,N_20243);
nor U24415 (N_24415,N_21436,N_21570);
or U24416 (N_24416,N_19895,N_19584);
nand U24417 (N_24417,N_19134,N_20118);
and U24418 (N_24418,N_19112,N_20352);
and U24419 (N_24419,N_21775,N_20469);
nor U24420 (N_24420,N_21496,N_20551);
or U24421 (N_24421,N_18901,N_19085);
nor U24422 (N_24422,N_21398,N_21685);
nand U24423 (N_24423,N_18900,N_18833);
nor U24424 (N_24424,N_21676,N_19481);
or U24425 (N_24425,N_20993,N_20470);
xor U24426 (N_24426,N_21150,N_20835);
or U24427 (N_24427,N_19626,N_20364);
nor U24428 (N_24428,N_21499,N_21529);
and U24429 (N_24429,N_21097,N_19314);
nand U24430 (N_24430,N_19956,N_21534);
nor U24431 (N_24431,N_19585,N_20832);
nor U24432 (N_24432,N_21855,N_19893);
nand U24433 (N_24433,N_19591,N_21802);
nand U24434 (N_24434,N_21307,N_21847);
nor U24435 (N_24435,N_20647,N_21356);
nor U24436 (N_24436,N_20399,N_20886);
nor U24437 (N_24437,N_19328,N_18855);
nand U24438 (N_24438,N_21281,N_21021);
nor U24439 (N_24439,N_19241,N_21830);
nand U24440 (N_24440,N_19068,N_19445);
or U24441 (N_24441,N_20028,N_19278);
nand U24442 (N_24442,N_20615,N_20989);
and U24443 (N_24443,N_20226,N_21308);
and U24444 (N_24444,N_18841,N_18987);
or U24445 (N_24445,N_20922,N_21676);
nor U24446 (N_24446,N_18949,N_20570);
nand U24447 (N_24447,N_19152,N_19958);
or U24448 (N_24448,N_20341,N_19182);
and U24449 (N_24449,N_21243,N_19239);
nand U24450 (N_24450,N_21456,N_20529);
nand U24451 (N_24451,N_19565,N_19839);
nand U24452 (N_24452,N_21113,N_19707);
and U24453 (N_24453,N_21232,N_21774);
xnor U24454 (N_24454,N_20421,N_21399);
xor U24455 (N_24455,N_21279,N_21671);
and U24456 (N_24456,N_19788,N_20836);
or U24457 (N_24457,N_21855,N_21761);
nor U24458 (N_24458,N_18793,N_19342);
and U24459 (N_24459,N_21262,N_20504);
nand U24460 (N_24460,N_19526,N_20774);
nor U24461 (N_24461,N_19424,N_20749);
xor U24462 (N_24462,N_21049,N_18865);
and U24463 (N_24463,N_18835,N_19647);
nor U24464 (N_24464,N_20511,N_21593);
nand U24465 (N_24465,N_20956,N_21780);
xor U24466 (N_24466,N_21040,N_21771);
or U24467 (N_24467,N_19148,N_20170);
or U24468 (N_24468,N_19471,N_19043);
and U24469 (N_24469,N_20543,N_21652);
nand U24470 (N_24470,N_20331,N_19059);
nor U24471 (N_24471,N_20013,N_20167);
nor U24472 (N_24472,N_19020,N_21421);
and U24473 (N_24473,N_19565,N_21851);
and U24474 (N_24474,N_19357,N_18838);
nand U24475 (N_24475,N_21707,N_19211);
nor U24476 (N_24476,N_21658,N_19461);
and U24477 (N_24477,N_21492,N_20200);
xor U24478 (N_24478,N_18910,N_20127);
and U24479 (N_24479,N_20997,N_18852);
nor U24480 (N_24480,N_21124,N_20928);
and U24481 (N_24481,N_19779,N_19850);
nor U24482 (N_24482,N_19731,N_21698);
nand U24483 (N_24483,N_21490,N_21652);
xnor U24484 (N_24484,N_19012,N_18932);
or U24485 (N_24485,N_18864,N_19406);
nor U24486 (N_24486,N_18760,N_18802);
nor U24487 (N_24487,N_20467,N_19494);
xnor U24488 (N_24488,N_20274,N_19567);
nand U24489 (N_24489,N_19983,N_21789);
and U24490 (N_24490,N_19719,N_21462);
nand U24491 (N_24491,N_21164,N_20693);
and U24492 (N_24492,N_19564,N_21373);
nand U24493 (N_24493,N_21611,N_19186);
nor U24494 (N_24494,N_21684,N_19523);
nor U24495 (N_24495,N_20324,N_19839);
nor U24496 (N_24496,N_20948,N_21707);
and U24497 (N_24497,N_20270,N_21010);
nand U24498 (N_24498,N_19976,N_21534);
nor U24499 (N_24499,N_19079,N_19546);
nor U24500 (N_24500,N_21353,N_21625);
nor U24501 (N_24501,N_19445,N_18929);
nor U24502 (N_24502,N_19271,N_20012);
nor U24503 (N_24503,N_21160,N_18924);
nor U24504 (N_24504,N_18949,N_20604);
nand U24505 (N_24505,N_19967,N_20971);
xor U24506 (N_24506,N_20279,N_19479);
or U24507 (N_24507,N_19094,N_21593);
or U24508 (N_24508,N_21389,N_21432);
nor U24509 (N_24509,N_21325,N_19715);
or U24510 (N_24510,N_20433,N_21446);
or U24511 (N_24511,N_20585,N_20663);
nand U24512 (N_24512,N_21713,N_19334);
nor U24513 (N_24513,N_21746,N_21212);
or U24514 (N_24514,N_20061,N_21145);
or U24515 (N_24515,N_21490,N_21018);
or U24516 (N_24516,N_19847,N_21711);
and U24517 (N_24517,N_21687,N_21766);
nor U24518 (N_24518,N_20290,N_20127);
nor U24519 (N_24519,N_19732,N_19135);
nand U24520 (N_24520,N_20565,N_21391);
xnor U24521 (N_24521,N_20304,N_18948);
nand U24522 (N_24522,N_18848,N_19788);
or U24523 (N_24523,N_21831,N_19809);
and U24524 (N_24524,N_20326,N_21060);
and U24525 (N_24525,N_20235,N_20379);
and U24526 (N_24526,N_19252,N_21235);
and U24527 (N_24527,N_19682,N_21535);
and U24528 (N_24528,N_20924,N_21318);
nor U24529 (N_24529,N_20811,N_19807);
xor U24530 (N_24530,N_19713,N_21581);
and U24531 (N_24531,N_21118,N_21860);
or U24532 (N_24532,N_20586,N_20487);
and U24533 (N_24533,N_19479,N_21728);
and U24534 (N_24534,N_21069,N_21531);
or U24535 (N_24535,N_20778,N_19795);
or U24536 (N_24536,N_19329,N_20301);
xor U24537 (N_24537,N_21182,N_21635);
or U24538 (N_24538,N_20851,N_20987);
nand U24539 (N_24539,N_20794,N_20269);
or U24540 (N_24540,N_19930,N_21654);
nand U24541 (N_24541,N_21629,N_19811);
and U24542 (N_24542,N_18938,N_21380);
and U24543 (N_24543,N_19358,N_19979);
nor U24544 (N_24544,N_20117,N_19049);
and U24545 (N_24545,N_18926,N_19697);
and U24546 (N_24546,N_19149,N_21378);
nor U24547 (N_24547,N_19302,N_21869);
nand U24548 (N_24548,N_20184,N_21441);
nand U24549 (N_24549,N_19665,N_19355);
nor U24550 (N_24550,N_20248,N_19777);
or U24551 (N_24551,N_19344,N_21828);
nand U24552 (N_24552,N_21598,N_21013);
nor U24553 (N_24553,N_21546,N_21206);
nand U24554 (N_24554,N_20236,N_20474);
and U24555 (N_24555,N_19644,N_20251);
nand U24556 (N_24556,N_20932,N_21360);
nor U24557 (N_24557,N_20426,N_20944);
and U24558 (N_24558,N_21604,N_19206);
nor U24559 (N_24559,N_21232,N_20167);
or U24560 (N_24560,N_20132,N_19154);
nor U24561 (N_24561,N_21176,N_19619);
xnor U24562 (N_24562,N_20679,N_20540);
nand U24563 (N_24563,N_20413,N_21204);
nand U24564 (N_24564,N_20369,N_21651);
nor U24565 (N_24565,N_20477,N_21391);
xnor U24566 (N_24566,N_20130,N_18917);
xnor U24567 (N_24567,N_19639,N_19251);
or U24568 (N_24568,N_18883,N_20575);
or U24569 (N_24569,N_19882,N_20127);
and U24570 (N_24570,N_19121,N_19992);
nor U24571 (N_24571,N_19080,N_19178);
xor U24572 (N_24572,N_19968,N_20623);
nor U24573 (N_24573,N_18984,N_20643);
or U24574 (N_24574,N_20459,N_19988);
or U24575 (N_24575,N_21568,N_20941);
nand U24576 (N_24576,N_20847,N_21710);
nand U24577 (N_24577,N_19205,N_19849);
nor U24578 (N_24578,N_19800,N_20100);
and U24579 (N_24579,N_21757,N_19231);
nand U24580 (N_24580,N_20441,N_20141);
nor U24581 (N_24581,N_21273,N_18952);
or U24582 (N_24582,N_20205,N_21709);
nor U24583 (N_24583,N_21072,N_21653);
nor U24584 (N_24584,N_21368,N_21269);
and U24585 (N_24585,N_21160,N_20339);
or U24586 (N_24586,N_20718,N_20429);
nand U24587 (N_24587,N_21170,N_21172);
nand U24588 (N_24588,N_19160,N_19886);
and U24589 (N_24589,N_19737,N_21731);
or U24590 (N_24590,N_21452,N_18941);
nand U24591 (N_24591,N_20802,N_19182);
and U24592 (N_24592,N_19299,N_19457);
nor U24593 (N_24593,N_19782,N_19658);
or U24594 (N_24594,N_19054,N_21753);
nand U24595 (N_24595,N_21540,N_21731);
nor U24596 (N_24596,N_20385,N_21750);
nand U24597 (N_24597,N_20258,N_19847);
nand U24598 (N_24598,N_19197,N_19486);
nor U24599 (N_24599,N_20764,N_21115);
nand U24600 (N_24600,N_21212,N_18980);
and U24601 (N_24601,N_19531,N_20480);
and U24602 (N_24602,N_19325,N_20756);
nor U24603 (N_24603,N_19315,N_19352);
and U24604 (N_24604,N_19210,N_20675);
nand U24605 (N_24605,N_20690,N_18905);
or U24606 (N_24606,N_20717,N_19947);
nor U24607 (N_24607,N_21066,N_20961);
or U24608 (N_24608,N_20096,N_19536);
nand U24609 (N_24609,N_19932,N_20672);
nand U24610 (N_24610,N_21839,N_20617);
nand U24611 (N_24611,N_21085,N_19018);
nand U24612 (N_24612,N_20835,N_18785);
and U24613 (N_24613,N_20605,N_20360);
xnor U24614 (N_24614,N_21071,N_19405);
nor U24615 (N_24615,N_19360,N_19797);
and U24616 (N_24616,N_18914,N_19548);
and U24617 (N_24617,N_20501,N_21255);
or U24618 (N_24618,N_21767,N_19218);
or U24619 (N_24619,N_21533,N_18868);
and U24620 (N_24620,N_21862,N_19139);
nor U24621 (N_24621,N_21834,N_20782);
xnor U24622 (N_24622,N_19252,N_19571);
nor U24623 (N_24623,N_19934,N_20220);
nor U24624 (N_24624,N_20832,N_19417);
and U24625 (N_24625,N_20436,N_19916);
nand U24626 (N_24626,N_20200,N_21526);
or U24627 (N_24627,N_19622,N_20185);
nor U24628 (N_24628,N_20144,N_20282);
nand U24629 (N_24629,N_20878,N_21455);
nor U24630 (N_24630,N_20028,N_21275);
nor U24631 (N_24631,N_21456,N_20726);
or U24632 (N_24632,N_21414,N_21621);
nand U24633 (N_24633,N_21039,N_21504);
nor U24634 (N_24634,N_19165,N_20891);
or U24635 (N_24635,N_21626,N_21671);
nand U24636 (N_24636,N_19391,N_21239);
and U24637 (N_24637,N_21538,N_19464);
xnor U24638 (N_24638,N_18925,N_20328);
nor U24639 (N_24639,N_21683,N_20759);
or U24640 (N_24640,N_21313,N_19903);
nand U24641 (N_24641,N_20910,N_19294);
xor U24642 (N_24642,N_21358,N_21228);
nand U24643 (N_24643,N_21717,N_21024);
or U24644 (N_24644,N_20477,N_21728);
nor U24645 (N_24645,N_21850,N_20605);
and U24646 (N_24646,N_19345,N_20879);
xor U24647 (N_24647,N_21305,N_21626);
nor U24648 (N_24648,N_21701,N_21734);
or U24649 (N_24649,N_19514,N_20664);
and U24650 (N_24650,N_20738,N_21401);
and U24651 (N_24651,N_21309,N_20318);
or U24652 (N_24652,N_20167,N_20871);
nor U24653 (N_24653,N_18832,N_19042);
nor U24654 (N_24654,N_21100,N_20127);
and U24655 (N_24655,N_19855,N_19310);
or U24656 (N_24656,N_20775,N_19799);
xnor U24657 (N_24657,N_21705,N_18763);
and U24658 (N_24658,N_19945,N_19496);
nor U24659 (N_24659,N_19075,N_20542);
or U24660 (N_24660,N_21497,N_19777);
and U24661 (N_24661,N_20554,N_19453);
or U24662 (N_24662,N_19935,N_20842);
nor U24663 (N_24663,N_20517,N_21223);
or U24664 (N_24664,N_21033,N_19524);
nand U24665 (N_24665,N_20335,N_19583);
nor U24666 (N_24666,N_21672,N_20093);
nor U24667 (N_24667,N_21519,N_20684);
or U24668 (N_24668,N_20740,N_20321);
and U24669 (N_24669,N_21695,N_21679);
and U24670 (N_24670,N_20550,N_19227);
and U24671 (N_24671,N_20997,N_20266);
xor U24672 (N_24672,N_20423,N_18853);
or U24673 (N_24673,N_21250,N_19920);
nand U24674 (N_24674,N_19250,N_21294);
nor U24675 (N_24675,N_19271,N_19623);
or U24676 (N_24676,N_20785,N_19292);
and U24677 (N_24677,N_19191,N_18993);
nor U24678 (N_24678,N_20818,N_19325);
xnor U24679 (N_24679,N_18872,N_20417);
and U24680 (N_24680,N_20778,N_19317);
nand U24681 (N_24681,N_19842,N_20827);
nand U24682 (N_24682,N_20414,N_20438);
or U24683 (N_24683,N_21029,N_20770);
nor U24684 (N_24684,N_20031,N_20369);
nand U24685 (N_24685,N_19100,N_19415);
or U24686 (N_24686,N_21003,N_20727);
or U24687 (N_24687,N_19446,N_19269);
or U24688 (N_24688,N_20733,N_20857);
nor U24689 (N_24689,N_21067,N_20369);
nor U24690 (N_24690,N_20133,N_20982);
xor U24691 (N_24691,N_20642,N_19142);
nor U24692 (N_24692,N_20763,N_18794);
and U24693 (N_24693,N_19132,N_19230);
nor U24694 (N_24694,N_21111,N_20601);
nand U24695 (N_24695,N_20313,N_21561);
xor U24696 (N_24696,N_21826,N_21616);
and U24697 (N_24697,N_20077,N_20085);
and U24698 (N_24698,N_21850,N_19310);
nand U24699 (N_24699,N_20216,N_21214);
and U24700 (N_24700,N_19062,N_20762);
nand U24701 (N_24701,N_19323,N_19045);
nor U24702 (N_24702,N_21546,N_19376);
nor U24703 (N_24703,N_20458,N_20767);
nand U24704 (N_24704,N_20231,N_19235);
nand U24705 (N_24705,N_19570,N_19518);
or U24706 (N_24706,N_20459,N_19000);
and U24707 (N_24707,N_21769,N_20864);
nand U24708 (N_24708,N_19610,N_19933);
nand U24709 (N_24709,N_19134,N_19468);
xnor U24710 (N_24710,N_21427,N_20646);
or U24711 (N_24711,N_19200,N_21662);
or U24712 (N_24712,N_21400,N_20155);
nand U24713 (N_24713,N_19481,N_21144);
nand U24714 (N_24714,N_21046,N_19613);
nor U24715 (N_24715,N_19419,N_20578);
and U24716 (N_24716,N_21028,N_21527);
or U24717 (N_24717,N_20816,N_19325);
xnor U24718 (N_24718,N_21790,N_19810);
nand U24719 (N_24719,N_20377,N_19533);
nand U24720 (N_24720,N_20336,N_21007);
nand U24721 (N_24721,N_20785,N_21189);
xnor U24722 (N_24722,N_21674,N_20135);
or U24723 (N_24723,N_18840,N_21499);
nand U24724 (N_24724,N_21530,N_21793);
nand U24725 (N_24725,N_21613,N_18927);
nand U24726 (N_24726,N_20559,N_21732);
or U24727 (N_24727,N_20751,N_21103);
and U24728 (N_24728,N_21329,N_19806);
nand U24729 (N_24729,N_21756,N_19739);
nor U24730 (N_24730,N_18779,N_19189);
xnor U24731 (N_24731,N_19590,N_19505);
and U24732 (N_24732,N_18968,N_18882);
and U24733 (N_24733,N_21041,N_20417);
nand U24734 (N_24734,N_19388,N_21753);
or U24735 (N_24735,N_20577,N_20624);
nor U24736 (N_24736,N_19728,N_21223);
xnor U24737 (N_24737,N_19720,N_20773);
nor U24738 (N_24738,N_19352,N_21490);
and U24739 (N_24739,N_21009,N_20805);
or U24740 (N_24740,N_19895,N_19363);
xor U24741 (N_24741,N_19373,N_20455);
or U24742 (N_24742,N_18818,N_20931);
nor U24743 (N_24743,N_19208,N_21609);
nor U24744 (N_24744,N_19330,N_19526);
xnor U24745 (N_24745,N_20631,N_18787);
nand U24746 (N_24746,N_21784,N_20330);
nand U24747 (N_24747,N_21108,N_19341);
nor U24748 (N_24748,N_19841,N_18883);
or U24749 (N_24749,N_21616,N_20356);
xor U24750 (N_24750,N_20228,N_21736);
or U24751 (N_24751,N_20568,N_20133);
nand U24752 (N_24752,N_18848,N_20851);
or U24753 (N_24753,N_21360,N_20533);
nor U24754 (N_24754,N_19526,N_21086);
or U24755 (N_24755,N_21492,N_20988);
and U24756 (N_24756,N_21639,N_19544);
nor U24757 (N_24757,N_20505,N_19345);
xor U24758 (N_24758,N_21426,N_20609);
and U24759 (N_24759,N_21116,N_19651);
and U24760 (N_24760,N_21827,N_19670);
or U24761 (N_24761,N_20398,N_19242);
or U24762 (N_24762,N_20831,N_21422);
nand U24763 (N_24763,N_20895,N_19193);
xnor U24764 (N_24764,N_19623,N_21673);
and U24765 (N_24765,N_19946,N_18967);
or U24766 (N_24766,N_21359,N_20689);
and U24767 (N_24767,N_18759,N_21463);
or U24768 (N_24768,N_21093,N_20541);
or U24769 (N_24769,N_20405,N_21699);
xor U24770 (N_24770,N_20699,N_21850);
nor U24771 (N_24771,N_20832,N_19817);
nor U24772 (N_24772,N_20247,N_18787);
xor U24773 (N_24773,N_19058,N_21506);
and U24774 (N_24774,N_20432,N_21055);
and U24775 (N_24775,N_19889,N_21847);
nand U24776 (N_24776,N_20202,N_21185);
and U24777 (N_24777,N_20213,N_21118);
nand U24778 (N_24778,N_21060,N_21699);
xnor U24779 (N_24779,N_20161,N_21370);
nor U24780 (N_24780,N_19092,N_21068);
xor U24781 (N_24781,N_19427,N_21698);
and U24782 (N_24782,N_19660,N_20140);
or U24783 (N_24783,N_18777,N_19862);
nand U24784 (N_24784,N_19982,N_20127);
nand U24785 (N_24785,N_19122,N_19858);
nand U24786 (N_24786,N_19989,N_18781);
or U24787 (N_24787,N_19530,N_21829);
or U24788 (N_24788,N_19412,N_19021);
nor U24789 (N_24789,N_19121,N_19442);
nor U24790 (N_24790,N_21567,N_20255);
and U24791 (N_24791,N_20623,N_20535);
and U24792 (N_24792,N_20020,N_19141);
or U24793 (N_24793,N_21441,N_19288);
nor U24794 (N_24794,N_21730,N_19334);
or U24795 (N_24795,N_21222,N_20525);
nand U24796 (N_24796,N_21344,N_19085);
nand U24797 (N_24797,N_20819,N_20412);
and U24798 (N_24798,N_21609,N_19424);
nor U24799 (N_24799,N_18857,N_20021);
or U24800 (N_24800,N_21509,N_20296);
or U24801 (N_24801,N_21063,N_20197);
xnor U24802 (N_24802,N_19744,N_19616);
nand U24803 (N_24803,N_21151,N_21129);
or U24804 (N_24804,N_21617,N_20864);
nand U24805 (N_24805,N_20657,N_19102);
or U24806 (N_24806,N_19460,N_20416);
or U24807 (N_24807,N_19551,N_19277);
or U24808 (N_24808,N_20277,N_19541);
nor U24809 (N_24809,N_20501,N_20946);
nor U24810 (N_24810,N_19241,N_19386);
nand U24811 (N_24811,N_21822,N_19901);
nand U24812 (N_24812,N_21410,N_19682);
nor U24813 (N_24813,N_21282,N_19920);
or U24814 (N_24814,N_18776,N_21674);
xor U24815 (N_24815,N_21265,N_19906);
nor U24816 (N_24816,N_19750,N_20527);
and U24817 (N_24817,N_20844,N_21289);
nand U24818 (N_24818,N_20473,N_21350);
nand U24819 (N_24819,N_21748,N_21235);
nor U24820 (N_24820,N_19177,N_18850);
xor U24821 (N_24821,N_20203,N_19752);
or U24822 (N_24822,N_19360,N_20174);
nand U24823 (N_24823,N_21843,N_21531);
xnor U24824 (N_24824,N_20724,N_21545);
nor U24825 (N_24825,N_21701,N_19902);
xor U24826 (N_24826,N_20233,N_20635);
nand U24827 (N_24827,N_20766,N_20391);
and U24828 (N_24828,N_20753,N_19266);
or U24829 (N_24829,N_21018,N_19079);
and U24830 (N_24830,N_20513,N_19689);
nor U24831 (N_24831,N_19562,N_20194);
nand U24832 (N_24832,N_19578,N_21263);
or U24833 (N_24833,N_19825,N_19119);
and U24834 (N_24834,N_19811,N_20866);
and U24835 (N_24835,N_21858,N_21491);
nor U24836 (N_24836,N_18823,N_20181);
nand U24837 (N_24837,N_18921,N_19124);
or U24838 (N_24838,N_19432,N_20036);
and U24839 (N_24839,N_20216,N_21513);
nor U24840 (N_24840,N_21183,N_18830);
nand U24841 (N_24841,N_19372,N_19653);
or U24842 (N_24842,N_20498,N_21045);
and U24843 (N_24843,N_20815,N_21577);
or U24844 (N_24844,N_19047,N_21406);
nand U24845 (N_24845,N_21452,N_18973);
nor U24846 (N_24846,N_20255,N_19785);
and U24847 (N_24847,N_19170,N_21180);
xor U24848 (N_24848,N_19754,N_19719);
nor U24849 (N_24849,N_20109,N_21602);
nand U24850 (N_24850,N_21682,N_20581);
or U24851 (N_24851,N_21404,N_20251);
nor U24852 (N_24852,N_20863,N_21366);
and U24853 (N_24853,N_19143,N_19106);
or U24854 (N_24854,N_20040,N_20552);
xnor U24855 (N_24855,N_19236,N_20740);
nand U24856 (N_24856,N_21256,N_19764);
and U24857 (N_24857,N_21541,N_21438);
nand U24858 (N_24858,N_20779,N_20469);
nor U24859 (N_24859,N_20663,N_21527);
and U24860 (N_24860,N_19928,N_18781);
nor U24861 (N_24861,N_20573,N_20093);
and U24862 (N_24862,N_19976,N_21127);
nor U24863 (N_24863,N_19966,N_20424);
and U24864 (N_24864,N_21854,N_20995);
or U24865 (N_24865,N_20725,N_19708);
and U24866 (N_24866,N_20046,N_21390);
xor U24867 (N_24867,N_21770,N_19474);
or U24868 (N_24868,N_21259,N_19922);
or U24869 (N_24869,N_21776,N_18852);
xnor U24870 (N_24870,N_21633,N_21058);
or U24871 (N_24871,N_21532,N_18831);
nand U24872 (N_24872,N_18961,N_21861);
or U24873 (N_24873,N_20866,N_21450);
nor U24874 (N_24874,N_20741,N_20577);
or U24875 (N_24875,N_19837,N_19593);
or U24876 (N_24876,N_21725,N_20174);
or U24877 (N_24877,N_20961,N_20686);
nand U24878 (N_24878,N_20069,N_20625);
nand U24879 (N_24879,N_19769,N_19065);
xor U24880 (N_24880,N_19384,N_21356);
nand U24881 (N_24881,N_20917,N_20872);
nor U24882 (N_24882,N_21749,N_21808);
nand U24883 (N_24883,N_19621,N_21717);
and U24884 (N_24884,N_19529,N_21369);
and U24885 (N_24885,N_21178,N_19365);
nor U24886 (N_24886,N_20023,N_20645);
nor U24887 (N_24887,N_19734,N_19894);
nor U24888 (N_24888,N_20396,N_21541);
nand U24889 (N_24889,N_20265,N_18898);
xnor U24890 (N_24890,N_19239,N_19583);
nor U24891 (N_24891,N_21028,N_21770);
nand U24892 (N_24892,N_20645,N_19393);
nand U24893 (N_24893,N_19683,N_21007);
nand U24894 (N_24894,N_21114,N_18908);
or U24895 (N_24895,N_21226,N_18843);
and U24896 (N_24896,N_20149,N_18813);
and U24897 (N_24897,N_20932,N_21156);
or U24898 (N_24898,N_20248,N_21489);
or U24899 (N_24899,N_19619,N_21284);
nand U24900 (N_24900,N_19909,N_19262);
and U24901 (N_24901,N_19123,N_19245);
or U24902 (N_24902,N_18805,N_18750);
and U24903 (N_24903,N_18964,N_19137);
and U24904 (N_24904,N_20186,N_20655);
or U24905 (N_24905,N_20933,N_19348);
nor U24906 (N_24906,N_21824,N_20626);
or U24907 (N_24907,N_21017,N_20741);
or U24908 (N_24908,N_20328,N_21047);
nor U24909 (N_24909,N_21198,N_21219);
xnor U24910 (N_24910,N_20553,N_21660);
nor U24911 (N_24911,N_19827,N_18990);
nor U24912 (N_24912,N_19532,N_21150);
nand U24913 (N_24913,N_19257,N_20330);
nor U24914 (N_24914,N_20726,N_21408);
or U24915 (N_24915,N_21784,N_20849);
nand U24916 (N_24916,N_19884,N_20701);
nor U24917 (N_24917,N_19661,N_20523);
or U24918 (N_24918,N_19138,N_20742);
and U24919 (N_24919,N_20409,N_19033);
xor U24920 (N_24920,N_21807,N_19134);
or U24921 (N_24921,N_19773,N_20669);
or U24922 (N_24922,N_19249,N_18833);
and U24923 (N_24923,N_21187,N_19148);
or U24924 (N_24924,N_20979,N_19540);
and U24925 (N_24925,N_21566,N_21117);
or U24926 (N_24926,N_19609,N_21674);
and U24927 (N_24927,N_20447,N_18905);
or U24928 (N_24928,N_21116,N_18881);
nor U24929 (N_24929,N_18841,N_20255);
nand U24930 (N_24930,N_19017,N_19851);
nand U24931 (N_24931,N_21831,N_18846);
or U24932 (N_24932,N_18834,N_19528);
or U24933 (N_24933,N_21645,N_19466);
xor U24934 (N_24934,N_19044,N_20037);
and U24935 (N_24935,N_20563,N_20426);
or U24936 (N_24936,N_21614,N_21101);
nor U24937 (N_24937,N_21358,N_19277);
nand U24938 (N_24938,N_21460,N_21805);
nand U24939 (N_24939,N_20957,N_20098);
nand U24940 (N_24940,N_19366,N_21587);
nand U24941 (N_24941,N_20079,N_19781);
and U24942 (N_24942,N_20421,N_21587);
nand U24943 (N_24943,N_19068,N_21565);
or U24944 (N_24944,N_21592,N_20133);
nand U24945 (N_24945,N_20426,N_21699);
and U24946 (N_24946,N_18870,N_19136);
and U24947 (N_24947,N_21422,N_19574);
or U24948 (N_24948,N_19251,N_19616);
nand U24949 (N_24949,N_19787,N_19143);
nor U24950 (N_24950,N_20442,N_19001);
nand U24951 (N_24951,N_21111,N_18803);
and U24952 (N_24952,N_21123,N_20036);
nand U24953 (N_24953,N_19185,N_18849);
nor U24954 (N_24954,N_18864,N_19247);
nor U24955 (N_24955,N_20206,N_21532);
and U24956 (N_24956,N_19398,N_21434);
and U24957 (N_24957,N_20908,N_19623);
or U24958 (N_24958,N_19674,N_20322);
or U24959 (N_24959,N_21241,N_21791);
nor U24960 (N_24960,N_20227,N_20890);
nor U24961 (N_24961,N_21602,N_21203);
nor U24962 (N_24962,N_20704,N_19819);
nor U24963 (N_24963,N_21747,N_19593);
and U24964 (N_24964,N_20729,N_20852);
xor U24965 (N_24965,N_21842,N_21747);
nor U24966 (N_24966,N_21164,N_21100);
nand U24967 (N_24967,N_18897,N_21550);
or U24968 (N_24968,N_20240,N_19329);
nand U24969 (N_24969,N_19530,N_21038);
nor U24970 (N_24970,N_20449,N_20162);
and U24971 (N_24971,N_20407,N_19459);
or U24972 (N_24972,N_19142,N_21173);
or U24973 (N_24973,N_19462,N_21355);
or U24974 (N_24974,N_19139,N_21514);
and U24975 (N_24975,N_21434,N_21575);
or U24976 (N_24976,N_20389,N_18986);
or U24977 (N_24977,N_18884,N_21841);
nor U24978 (N_24978,N_20521,N_19972);
nand U24979 (N_24979,N_19236,N_19836);
nand U24980 (N_24980,N_20287,N_21393);
nor U24981 (N_24981,N_21117,N_18868);
or U24982 (N_24982,N_19012,N_20493);
and U24983 (N_24983,N_19062,N_18966);
xor U24984 (N_24984,N_21410,N_20966);
nand U24985 (N_24985,N_21104,N_21682);
and U24986 (N_24986,N_19355,N_19253);
or U24987 (N_24987,N_19979,N_21585);
or U24988 (N_24988,N_21048,N_19566);
and U24989 (N_24989,N_18755,N_20758);
nor U24990 (N_24990,N_19956,N_21137);
nand U24991 (N_24991,N_21328,N_20259);
nor U24992 (N_24992,N_21151,N_21828);
and U24993 (N_24993,N_20878,N_21180);
nor U24994 (N_24994,N_19500,N_21191);
nor U24995 (N_24995,N_21224,N_21824);
and U24996 (N_24996,N_19681,N_19555);
nand U24997 (N_24997,N_21738,N_18901);
and U24998 (N_24998,N_21517,N_20514);
nor U24999 (N_24999,N_19812,N_19383);
or UO_0 (O_0,N_23760,N_24805);
nor UO_1 (O_1,N_24714,N_22481);
or UO_2 (O_2,N_24122,N_24645);
or UO_3 (O_3,N_23154,N_23955);
and UO_4 (O_4,N_24051,N_24960);
nand UO_5 (O_5,N_22107,N_22797);
and UO_6 (O_6,N_24050,N_21964);
nor UO_7 (O_7,N_23579,N_22817);
xnor UO_8 (O_8,N_23457,N_24628);
nand UO_9 (O_9,N_24647,N_24396);
and UO_10 (O_10,N_23329,N_22049);
and UO_11 (O_11,N_22093,N_24015);
or UO_12 (O_12,N_22763,N_23821);
xnor UO_13 (O_13,N_22581,N_24848);
nor UO_14 (O_14,N_21918,N_24035);
nor UO_15 (O_15,N_22517,N_22976);
nand UO_16 (O_16,N_23657,N_24638);
nor UO_17 (O_17,N_24988,N_24721);
or UO_18 (O_18,N_24253,N_23722);
nor UO_19 (O_19,N_24288,N_23950);
xor UO_20 (O_20,N_22782,N_23290);
nor UO_21 (O_21,N_24662,N_22619);
nor UO_22 (O_22,N_22360,N_22243);
and UO_23 (O_23,N_23803,N_24926);
xnor UO_24 (O_24,N_24843,N_23951);
nand UO_25 (O_25,N_23309,N_24224);
nor UO_26 (O_26,N_23819,N_24434);
xor UO_27 (O_27,N_23436,N_24249);
or UO_28 (O_28,N_24517,N_22105);
or UO_29 (O_29,N_23670,N_23197);
nor UO_30 (O_30,N_22706,N_24295);
and UO_31 (O_31,N_23785,N_22847);
nand UO_32 (O_32,N_22810,N_23652);
or UO_33 (O_33,N_23391,N_24333);
and UO_34 (O_34,N_24591,N_24451);
or UO_35 (O_35,N_24460,N_22666);
nand UO_36 (O_36,N_23081,N_22341);
and UO_37 (O_37,N_24423,N_24703);
or UO_38 (O_38,N_23285,N_24707);
or UO_39 (O_39,N_24470,N_22074);
nand UO_40 (O_40,N_24189,N_22024);
and UO_41 (O_41,N_23859,N_23039);
nand UO_42 (O_42,N_24832,N_22048);
and UO_43 (O_43,N_22438,N_24398);
nor UO_44 (O_44,N_22597,N_22409);
and UO_45 (O_45,N_22121,N_22855);
nand UO_46 (O_46,N_23627,N_23608);
nand UO_47 (O_47,N_23614,N_23183);
xor UO_48 (O_48,N_22940,N_22367);
nand UO_49 (O_49,N_23289,N_23891);
or UO_50 (O_50,N_24261,N_24323);
nor UO_51 (O_51,N_21919,N_23105);
and UO_52 (O_52,N_24768,N_22411);
nor UO_53 (O_53,N_24632,N_24860);
and UO_54 (O_54,N_24927,N_23902);
nand UO_55 (O_55,N_23501,N_23866);
nand UO_56 (O_56,N_23581,N_24479);
or UO_57 (O_57,N_22334,N_23211);
and UO_58 (O_58,N_23116,N_23621);
or UO_59 (O_59,N_23447,N_24990);
nand UO_60 (O_60,N_24448,N_22203);
or UO_61 (O_61,N_23299,N_23212);
or UO_62 (O_62,N_22931,N_22480);
nand UO_63 (O_63,N_21953,N_23326);
or UO_64 (O_64,N_23537,N_22189);
or UO_65 (O_65,N_23966,N_24369);
or UO_66 (O_66,N_22960,N_22679);
nand UO_67 (O_67,N_23536,N_24871);
nand UO_68 (O_68,N_23871,N_24840);
nand UO_69 (O_69,N_24153,N_22368);
and UO_70 (O_70,N_24180,N_22654);
and UO_71 (O_71,N_23339,N_24314);
or UO_72 (O_72,N_23179,N_23741);
or UO_73 (O_73,N_22485,N_22874);
nand UO_74 (O_74,N_24294,N_23086);
nor UO_75 (O_75,N_22917,N_22443);
and UO_76 (O_76,N_22171,N_22195);
or UO_77 (O_77,N_23172,N_22290);
and UO_78 (O_78,N_23907,N_22859);
or UO_79 (O_79,N_24718,N_22769);
or UO_80 (O_80,N_23952,N_23522);
nor UO_81 (O_81,N_24354,N_22008);
nand UO_82 (O_82,N_23142,N_23108);
nor UO_83 (O_83,N_22349,N_23720);
and UO_84 (O_84,N_24363,N_22780);
and UO_85 (O_85,N_23698,N_23558);
xnor UO_86 (O_86,N_24762,N_22030);
or UO_87 (O_87,N_24538,N_23982);
nor UO_88 (O_88,N_22956,N_24390);
nor UO_89 (O_89,N_24586,N_23257);
and UO_90 (O_90,N_24709,N_22773);
nor UO_91 (O_91,N_24164,N_23707);
or UO_92 (O_92,N_22651,N_22882);
and UO_93 (O_93,N_24684,N_23607);
and UO_94 (O_94,N_21915,N_22986);
or UO_95 (O_95,N_23931,N_24306);
or UO_96 (O_96,N_24968,N_22110);
nand UO_97 (O_97,N_23682,N_23458);
nor UO_98 (O_98,N_24534,N_23502);
xor UO_99 (O_99,N_23188,N_22149);
or UO_100 (O_100,N_24811,N_22629);
nor UO_101 (O_101,N_22725,N_24523);
or UO_102 (O_102,N_24338,N_24063);
and UO_103 (O_103,N_24610,N_24175);
nand UO_104 (O_104,N_23876,N_23481);
nor UO_105 (O_105,N_23918,N_22310);
and UO_106 (O_106,N_23420,N_23487);
and UO_107 (O_107,N_24242,N_23750);
and UO_108 (O_108,N_22661,N_23667);
or UO_109 (O_109,N_23439,N_24230);
or UO_110 (O_110,N_22636,N_22196);
nand UO_111 (O_111,N_21947,N_22785);
and UO_112 (O_112,N_24627,N_22467);
and UO_113 (O_113,N_23157,N_21949);
nor UO_114 (O_114,N_22138,N_23362);
nand UO_115 (O_115,N_24930,N_23830);
nand UO_116 (O_116,N_22113,N_23195);
or UO_117 (O_117,N_22742,N_24594);
and UO_118 (O_118,N_24207,N_21928);
or UO_119 (O_119,N_24644,N_22760);
xor UO_120 (O_120,N_22887,N_23280);
nor UO_121 (O_121,N_23994,N_23926);
nor UO_122 (O_122,N_24076,N_22757);
nor UO_123 (O_123,N_23307,N_23820);
nor UO_124 (O_124,N_23292,N_24849);
or UO_125 (O_125,N_23019,N_22789);
nor UO_126 (O_126,N_22621,N_24255);
or UO_127 (O_127,N_24459,N_21893);
xnor UO_128 (O_128,N_24218,N_22090);
nand UO_129 (O_129,N_24982,N_22431);
xnor UO_130 (O_130,N_23184,N_24400);
nand UO_131 (O_131,N_22820,N_22217);
and UO_132 (O_132,N_23654,N_22015);
nor UO_133 (O_133,N_23409,N_22415);
or UO_134 (O_134,N_24842,N_23113);
nand UO_135 (O_135,N_23156,N_23322);
nand UO_136 (O_136,N_22447,N_24521);
xor UO_137 (O_137,N_23602,N_23605);
nor UO_138 (O_138,N_24496,N_24943);
xnor UO_139 (O_139,N_24222,N_24085);
and UO_140 (O_140,N_23533,N_23041);
and UO_141 (O_141,N_23323,N_24098);
and UO_142 (O_142,N_24743,N_23161);
nand UO_143 (O_143,N_22944,N_24075);
xor UO_144 (O_144,N_22028,N_24724);
nor UO_145 (O_145,N_23435,N_23864);
or UO_146 (O_146,N_23867,N_24600);
and UO_147 (O_147,N_22212,N_23890);
or UO_148 (O_148,N_23240,N_22292);
or UO_149 (O_149,N_22169,N_22697);
nor UO_150 (O_150,N_23745,N_23571);
nor UO_151 (O_151,N_23650,N_22045);
nor UO_152 (O_152,N_22372,N_24522);
or UO_153 (O_153,N_23776,N_23526);
or UO_154 (O_154,N_22703,N_22159);
xnor UO_155 (O_155,N_22058,N_21940);
nand UO_156 (O_156,N_24786,N_24206);
nor UO_157 (O_157,N_24000,N_24851);
nand UO_158 (O_158,N_22178,N_22907);
or UO_159 (O_159,N_23151,N_24009);
nor UO_160 (O_160,N_22059,N_21938);
nor UO_161 (O_161,N_22949,N_23958);
nor UO_162 (O_162,N_22357,N_24066);
and UO_163 (O_163,N_24007,N_22803);
and UO_164 (O_164,N_22036,N_22700);
nor UO_165 (O_165,N_23730,N_24228);
or UO_166 (O_166,N_24838,N_24212);
xor UO_167 (O_167,N_23794,N_23315);
nand UO_168 (O_168,N_22454,N_23740);
nand UO_169 (O_169,N_24512,N_22380);
and UO_170 (O_170,N_23628,N_22614);
nand UO_171 (O_171,N_24781,N_22516);
or UO_172 (O_172,N_22115,N_23408);
or UO_173 (O_173,N_22604,N_24486);
nor UO_174 (O_174,N_24734,N_22375);
nor UO_175 (O_175,N_24145,N_21891);
or UO_176 (O_176,N_21966,N_24996);
nor UO_177 (O_177,N_24682,N_23972);
and UO_178 (O_178,N_23219,N_23368);
or UO_179 (O_179,N_22741,N_24944);
or UO_180 (O_180,N_23646,N_24862);
nand UO_181 (O_181,N_22131,N_24174);
nand UO_182 (O_182,N_24331,N_23726);
and UO_183 (O_183,N_24214,N_24623);
and UO_184 (O_184,N_23059,N_24322);
or UO_185 (O_185,N_23564,N_24308);
or UO_186 (O_186,N_24760,N_23078);
or UO_187 (O_187,N_23947,N_21988);
and UO_188 (O_188,N_24090,N_24317);
nand UO_189 (O_189,N_24771,N_22507);
nand UO_190 (O_190,N_22278,N_24678);
xor UO_191 (O_191,N_24258,N_23150);
and UO_192 (O_192,N_24956,N_23512);
and UO_193 (O_193,N_23016,N_22012);
nand UO_194 (O_194,N_23675,N_22823);
nor UO_195 (O_195,N_24116,N_24565);
and UO_196 (O_196,N_22937,N_24782);
nor UO_197 (O_197,N_23499,N_24531);
nor UO_198 (O_198,N_21897,N_22222);
nor UO_199 (O_199,N_24213,N_22816);
or UO_200 (O_200,N_23459,N_22762);
and UO_201 (O_201,N_24827,N_24658);
nor UO_202 (O_202,N_23206,N_22497);
and UO_203 (O_203,N_23045,N_24710);
nor UO_204 (O_204,N_22205,N_23539);
or UO_205 (O_205,N_24118,N_24494);
nand UO_206 (O_206,N_24328,N_24487);
xor UO_207 (O_207,N_23773,N_23495);
xor UO_208 (O_208,N_23400,N_23699);
nor UO_209 (O_209,N_24360,N_23026);
nand UO_210 (O_210,N_24110,N_22892);
and UO_211 (O_211,N_24028,N_22401);
nand UO_212 (O_212,N_22470,N_24023);
nor UO_213 (O_213,N_24598,N_23412);
or UO_214 (O_214,N_22704,N_22201);
xor UO_215 (O_215,N_22686,N_23460);
and UO_216 (O_216,N_22183,N_22003);
or UO_217 (O_217,N_22851,N_22649);
xor UO_218 (O_218,N_23567,N_23523);
nand UO_219 (O_219,N_21934,N_23983);
nand UO_220 (O_220,N_24621,N_23208);
nor UO_221 (O_221,N_24095,N_22391);
or UO_222 (O_222,N_21914,N_22064);
or UO_223 (O_223,N_22968,N_23075);
nand UO_224 (O_224,N_23549,N_23014);
nand UO_225 (O_225,N_22740,N_23110);
or UO_226 (O_226,N_23297,N_23111);
nand UO_227 (O_227,N_24711,N_23656);
nand UO_228 (O_228,N_22256,N_24029);
nand UO_229 (O_229,N_22002,N_22077);
or UO_230 (O_230,N_24651,N_23347);
xor UO_231 (O_231,N_22079,N_24749);
nor UO_232 (O_232,N_23247,N_22471);
and UO_233 (O_233,N_22580,N_22673);
nor UO_234 (O_234,N_24587,N_24217);
nand UO_235 (O_235,N_22425,N_22439);
xnor UO_236 (O_236,N_23937,N_23274);
nor UO_237 (O_237,N_23239,N_24379);
nor UO_238 (O_238,N_24411,N_22839);
or UO_239 (O_239,N_23189,N_23968);
or UO_240 (O_240,N_24895,N_22548);
and UO_241 (O_241,N_24361,N_22726);
and UO_242 (O_242,N_22728,N_22599);
nand UO_243 (O_243,N_22687,N_22230);
nand UO_244 (O_244,N_24093,N_22618);
nand UO_245 (O_245,N_24819,N_22366);
xor UO_246 (O_246,N_22933,N_24747);
and UO_247 (O_247,N_24624,N_22116);
nand UO_248 (O_248,N_24466,N_24143);
nand UO_249 (O_249,N_24399,N_24863);
or UO_250 (O_250,N_23777,N_22111);
xnor UO_251 (O_251,N_24829,N_22043);
or UO_252 (O_252,N_23747,N_22530);
xnor UO_253 (O_253,N_22297,N_24391);
and UO_254 (O_254,N_22206,N_23671);
nand UO_255 (O_255,N_23023,N_23079);
xor UO_256 (O_256,N_24527,N_23648);
xor UO_257 (O_257,N_22386,N_23603);
xnor UO_258 (O_258,N_22020,N_24185);
or UO_259 (O_259,N_23573,N_23258);
nand UO_260 (O_260,N_23162,N_23528);
nand UO_261 (O_261,N_22466,N_24570);
nor UO_262 (O_262,N_24103,N_22369);
or UO_263 (O_263,N_23152,N_22495);
or UO_264 (O_264,N_24650,N_24204);
nor UO_265 (O_265,N_23957,N_21921);
xor UO_266 (O_266,N_23749,N_24952);
or UO_267 (O_267,N_22458,N_23869);
and UO_268 (O_268,N_23087,N_22493);
or UO_269 (O_269,N_23538,N_24022);
and UO_270 (O_270,N_23281,N_23555);
nor UO_271 (O_271,N_24488,N_23886);
and UO_272 (O_272,N_24528,N_24789);
nand UO_273 (O_273,N_24089,N_24526);
or UO_274 (O_274,N_23963,N_23916);
or UO_275 (O_275,N_24705,N_22583);
nor UO_276 (O_276,N_22050,N_22716);
nand UO_277 (O_277,N_22707,N_23361);
xnor UO_278 (O_278,N_22743,N_22009);
or UO_279 (O_279,N_24584,N_23532);
or UO_280 (O_280,N_24904,N_24043);
xnor UO_281 (O_281,N_23974,N_24237);
or UO_282 (O_282,N_24962,N_23592);
and UO_283 (O_283,N_22691,N_23805);
nand UO_284 (O_284,N_23180,N_23898);
or UO_285 (O_285,N_23370,N_23328);
or UO_286 (O_286,N_23076,N_23012);
nor UO_287 (O_287,N_23787,N_22306);
and UO_288 (O_288,N_24349,N_23742);
and UO_289 (O_289,N_23992,N_22300);
or UO_290 (O_290,N_23417,N_23753);
nor UO_291 (O_291,N_22041,N_22199);
nand UO_292 (O_292,N_23256,N_24184);
or UO_293 (O_293,N_23810,N_22615);
nand UO_294 (O_294,N_24004,N_22815);
nor UO_295 (O_295,N_22753,N_23831);
and UO_296 (O_296,N_22525,N_24319);
or UO_297 (O_297,N_24558,N_24515);
or UO_298 (O_298,N_24774,N_23278);
or UO_299 (O_299,N_24967,N_23205);
and UO_300 (O_300,N_24113,N_22296);
nand UO_301 (O_301,N_21905,N_23393);
nand UO_302 (O_302,N_23949,N_22643);
nand UO_303 (O_303,N_22157,N_21941);
and UO_304 (O_304,N_24683,N_24005);
or UO_305 (O_305,N_23757,N_22927);
or UO_306 (O_306,N_24088,N_24065);
nand UO_307 (O_307,N_23715,N_24903);
nor UO_308 (O_308,N_23480,N_24304);
or UO_309 (O_309,N_23641,N_24769);
or UO_310 (O_310,N_23882,N_23633);
xnor UO_311 (O_311,N_24611,N_22318);
nor UO_312 (O_312,N_22544,N_24188);
or UO_313 (O_313,N_22570,N_23270);
xor UO_314 (O_314,N_22492,N_23367);
or UO_315 (O_315,N_22498,N_22903);
or UO_316 (O_316,N_23071,N_23330);
and UO_317 (O_317,N_23756,N_23489);
nor UO_318 (O_318,N_22957,N_24156);
nor UO_319 (O_319,N_23381,N_22881);
nor UO_320 (O_320,N_24563,N_24439);
nand UO_321 (O_321,N_23248,N_22130);
xnor UO_322 (O_322,N_24757,N_22972);
nor UO_323 (O_323,N_22648,N_22824);
xnor UO_324 (O_324,N_23478,N_23732);
or UO_325 (O_325,N_22985,N_22249);
or UO_326 (O_326,N_24588,N_22518);
xnor UO_327 (O_327,N_23193,N_22453);
or UO_328 (O_328,N_23975,N_23689);
nand UO_329 (O_329,N_23979,N_23948);
or UO_330 (O_330,N_24947,N_24582);
nand UO_331 (O_331,N_22229,N_22238);
nand UO_332 (O_332,N_24663,N_24745);
nand UO_333 (O_333,N_23121,N_23739);
and UO_334 (O_334,N_21971,N_24209);
nand UO_335 (O_335,N_24480,N_23575);
nor UO_336 (O_336,N_22579,N_22564);
xor UO_337 (O_337,N_23848,N_23123);
nand UO_338 (O_338,N_24514,N_23973);
nand UO_339 (O_339,N_23283,N_22371);
xor UO_340 (O_340,N_22647,N_23097);
nor UO_341 (O_341,N_22552,N_23768);
or UO_342 (O_342,N_24231,N_23941);
or UO_343 (O_343,N_22098,N_23818);
nand UO_344 (O_344,N_23935,N_23473);
nand UO_345 (O_345,N_22920,N_24267);
xor UO_346 (O_346,N_24060,N_22496);
nor UO_347 (O_347,N_24321,N_24637);
nand UO_348 (O_348,N_23342,N_24833);
nand UO_349 (O_349,N_22450,N_24419);
nand UO_350 (O_350,N_24585,N_23915);
nor UO_351 (O_351,N_22734,N_24081);
nand UO_352 (O_352,N_22016,N_24173);
and UO_353 (O_353,N_23235,N_22560);
nand UO_354 (O_354,N_24036,N_22692);
xnor UO_355 (O_355,N_22455,N_24096);
xnor UO_356 (O_356,N_22218,N_23229);
nor UO_357 (O_357,N_22756,N_23040);
and UO_358 (O_358,N_24355,N_22818);
and UO_359 (O_359,N_22754,N_24350);
nor UO_360 (O_360,N_23182,N_24019);
and UO_361 (O_361,N_23231,N_21959);
nand UO_362 (O_362,N_23680,N_23314);
nand UO_363 (O_363,N_24746,N_22658);
or UO_364 (O_364,N_22213,N_24375);
nand UO_365 (O_365,N_22919,N_21911);
or UO_366 (O_366,N_22587,N_24537);
nor UO_367 (O_367,N_22922,N_22977);
nor UO_368 (O_368,N_23761,N_22276);
xor UO_369 (O_369,N_24821,N_22633);
xor UO_370 (O_370,N_23634,N_24491);
nor UO_371 (O_371,N_23424,N_22025);
xor UO_372 (O_372,N_23717,N_24476);
nand UO_373 (O_373,N_24282,N_22299);
nor UO_374 (O_374,N_24497,N_22317);
and UO_375 (O_375,N_22699,N_24449);
nor UO_376 (O_376,N_22640,N_24802);
or UO_377 (O_377,N_23548,N_22677);
and UO_378 (O_378,N_23909,N_23175);
or UO_379 (O_379,N_24373,N_24420);
nor UO_380 (O_380,N_22711,N_21944);
nand UO_381 (O_381,N_23692,N_23686);
and UO_382 (O_382,N_22154,N_24775);
xnor UO_383 (O_383,N_24311,N_23286);
nor UO_384 (O_384,N_24418,N_23415);
nor UO_385 (O_385,N_23816,N_24884);
nand UO_386 (O_386,N_22427,N_22500);
or UO_387 (O_387,N_23827,N_22293);
or UO_388 (O_388,N_24999,N_22112);
or UO_389 (O_389,N_21948,N_23335);
or UO_390 (O_390,N_22071,N_24545);
nand UO_391 (O_391,N_22421,N_24928);
nor UO_392 (O_392,N_24720,N_23067);
nor UO_393 (O_393,N_23174,N_22186);
nand UO_394 (O_394,N_24911,N_22392);
and UO_395 (O_395,N_23333,N_23010);
and UO_396 (O_396,N_21989,N_21977);
or UO_397 (O_397,N_23492,N_23124);
and UO_398 (O_398,N_23325,N_22835);
or UO_399 (O_399,N_23243,N_22814);
and UO_400 (O_400,N_23246,N_24935);
nor UO_401 (O_401,N_24755,N_24371);
and UO_402 (O_402,N_23792,N_23535);
or UO_403 (O_403,N_24790,N_24607);
nand UO_404 (O_404,N_22047,N_24190);
and UO_405 (O_405,N_22849,N_22646);
nor UO_406 (O_406,N_23065,N_22227);
and UO_407 (O_407,N_22524,N_22204);
or UO_408 (O_408,N_22543,N_22042);
nand UO_409 (O_409,N_22906,N_22842);
nor UO_410 (O_410,N_23001,N_22489);
and UO_411 (O_411,N_23542,N_22232);
or UO_412 (O_412,N_21954,N_23047);
nand UO_413 (O_413,N_23098,N_24123);
and UO_414 (O_414,N_24200,N_24640);
and UO_415 (O_415,N_23629,N_23238);
or UO_416 (O_416,N_22277,N_22275);
and UO_417 (O_417,N_24454,N_22331);
nor UO_418 (O_418,N_22553,N_24394);
xnor UO_419 (O_419,N_23861,N_24908);
nor UO_420 (O_420,N_22744,N_24704);
nor UO_421 (O_421,N_23900,N_22608);
nor UO_422 (O_422,N_24412,N_24408);
nand UO_423 (O_423,N_22035,N_23386);
nand UO_424 (O_424,N_23378,N_24455);
nand UO_425 (O_425,N_23106,N_24378);
and UO_426 (O_426,N_24803,N_23999);
nor UO_427 (O_427,N_23568,N_22767);
nand UO_428 (O_428,N_24725,N_23933);
nand UO_429 (O_429,N_23808,N_22139);
nand UO_430 (O_430,N_24872,N_21906);
or UO_431 (O_431,N_23022,N_24529);
xnor UO_432 (O_432,N_23505,N_23399);
nand UO_433 (O_433,N_23406,N_24402);
nand UO_434 (O_434,N_22029,N_23889);
nor UO_435 (O_435,N_23600,N_22774);
or UO_436 (O_436,N_22622,N_23660);
and UO_437 (O_437,N_23702,N_22219);
or UO_438 (O_438,N_22582,N_24111);
nor UO_439 (O_439,N_24955,N_23485);
nor UO_440 (O_440,N_24826,N_23031);
and UO_441 (O_441,N_22979,N_22787);
nor UO_442 (O_442,N_24335,N_24524);
or UO_443 (O_443,N_23976,N_22689);
or UO_444 (O_444,N_23637,N_22394);
or UO_445 (O_445,N_24182,N_23829);
xnor UO_446 (O_446,N_24272,N_23885);
nor UO_447 (O_447,N_24263,N_24388);
and UO_448 (O_448,N_22819,N_23241);
or UO_449 (O_449,N_22348,N_22118);
or UO_450 (O_450,N_22312,N_23425);
and UO_451 (O_451,N_22676,N_22837);
and UO_452 (O_452,N_24866,N_24203);
nor UO_453 (O_453,N_22559,N_21894);
and UO_454 (O_454,N_22076,N_22260);
and UO_455 (O_455,N_23261,N_24717);
xnor UO_456 (O_456,N_23880,N_23448);
nor UO_457 (O_457,N_23883,N_23877);
nor UO_458 (O_458,N_23028,N_22990);
and UO_459 (O_459,N_22721,N_23594);
or UO_460 (O_460,N_22092,N_22684);
nor UO_461 (O_461,N_22938,N_23669);
or UO_462 (O_462,N_23013,N_22239);
nor UO_463 (O_463,N_23164,N_22182);
and UO_464 (O_464,N_22941,N_23562);
nor UO_465 (O_465,N_21956,N_22433);
nand UO_466 (O_466,N_22273,N_22326);
nand UO_467 (O_467,N_23483,N_24450);
xor UO_468 (O_468,N_22574,N_23438);
or UO_469 (O_469,N_22342,N_22430);
and UO_470 (O_470,N_22281,N_23431);
xor UO_471 (O_471,N_22536,N_23856);
nand UO_472 (O_472,N_23132,N_23475);
nor UO_473 (O_473,N_22996,N_24221);
and UO_474 (O_474,N_23057,N_22729);
nor UO_475 (O_475,N_24162,N_22935);
and UO_476 (O_476,N_24334,N_22175);
and UO_477 (O_477,N_23996,N_22595);
and UO_478 (O_478,N_22084,N_22683);
and UO_479 (O_479,N_22511,N_23080);
nor UO_480 (O_480,N_23355,N_24949);
or UO_481 (O_481,N_21903,N_22936);
nand UO_482 (O_482,N_24347,N_22625);
nor UO_483 (O_483,N_22613,N_23721);
nand UO_484 (O_484,N_24899,N_24812);
and UO_485 (O_485,N_22448,N_22840);
xnor UO_486 (O_486,N_22894,N_24958);
nand UO_487 (O_487,N_24176,N_22969);
xor UO_488 (O_488,N_24381,N_22735);
or UO_489 (O_489,N_23198,N_24235);
or UO_490 (O_490,N_22542,N_23863);
or UO_491 (O_491,N_22843,N_24887);
and UO_492 (O_492,N_22800,N_23337);
or UO_493 (O_493,N_24765,N_24744);
nand UO_494 (O_494,N_23601,N_24767);
nand UO_495 (O_495,N_23940,N_23868);
and UO_496 (O_496,N_22325,N_24299);
nor UO_497 (O_497,N_22083,N_23100);
nor UO_498 (O_498,N_22539,N_22033);
or UO_499 (O_499,N_22813,N_24027);
xnor UO_500 (O_500,N_22771,N_24691);
nor UO_501 (O_501,N_22503,N_24841);
or UO_502 (O_502,N_24079,N_21998);
xor UO_503 (O_503,N_23168,N_22383);
and UO_504 (O_504,N_22961,N_21942);
nor UO_505 (O_505,N_23396,N_21933);
or UO_506 (O_506,N_22054,N_22514);
nand UO_507 (O_507,N_22039,N_22953);
nand UO_508 (O_508,N_22627,N_24722);
and UO_509 (O_509,N_24868,N_24216);
nor UO_510 (O_510,N_23236,N_22280);
nand UO_511 (O_511,N_23755,N_24026);
nand UO_512 (O_512,N_22825,N_24877);
or UO_513 (O_513,N_22340,N_21986);
or UO_514 (O_514,N_24792,N_22695);
nand UO_515 (O_515,N_23569,N_24977);
or UO_516 (O_516,N_24974,N_23137);
and UO_517 (O_517,N_23096,N_22174);
nand UO_518 (O_518,N_23030,N_23520);
nand UO_519 (O_519,N_22305,N_22730);
nor UO_520 (O_520,N_23350,N_23872);
or UO_521 (O_521,N_23479,N_23120);
nor UO_522 (O_522,N_24754,N_23550);
or UO_523 (O_523,N_23965,N_23843);
nand UO_524 (O_524,N_22445,N_24502);
nand UO_525 (O_525,N_23062,N_22473);
and UO_526 (O_526,N_24791,N_22484);
and UO_527 (O_527,N_22124,N_23178);
or UO_528 (O_528,N_24431,N_24766);
or UO_529 (O_529,N_22713,N_24706);
and UO_530 (O_530,N_24874,N_22790);
or UO_531 (O_531,N_22404,N_23956);
nor UO_532 (O_532,N_22868,N_23407);
and UO_533 (O_533,N_23514,N_24161);
xor UO_534 (O_534,N_22491,N_23524);
and UO_535 (O_535,N_24395,N_22052);
nor UO_536 (O_536,N_23403,N_22314);
nor UO_537 (O_537,N_23273,N_24969);
nand UO_538 (O_538,N_24748,N_22739);
and UO_539 (O_539,N_24629,N_23875);
and UO_540 (O_540,N_24062,N_24112);
or UO_541 (O_541,N_24902,N_22457);
nor UO_542 (O_542,N_23049,N_22531);
or UO_543 (O_543,N_22027,N_24069);
nor UO_544 (O_544,N_21961,N_23678);
nor UO_545 (O_545,N_24397,N_21975);
nor UO_546 (O_546,N_23262,N_22623);
and UO_547 (O_547,N_22173,N_22632);
or UO_548 (O_548,N_23332,N_22541);
and UO_549 (O_549,N_21885,N_22593);
and UO_550 (O_550,N_22179,N_22418);
nand UO_551 (O_551,N_23673,N_22974);
xnor UO_552 (O_552,N_24474,N_24254);
nand UO_553 (O_553,N_22307,N_22528);
or UO_554 (O_554,N_23507,N_22952);
or UO_555 (O_555,N_23841,N_23027);
or UO_556 (O_556,N_22563,N_23371);
nor UO_557 (O_557,N_23985,N_23226);
or UO_558 (O_558,N_24879,N_23083);
or UO_559 (O_559,N_23181,N_24845);
nand UO_560 (O_560,N_22225,N_24787);
nor UO_561 (O_561,N_23731,N_22829);
and UO_562 (O_562,N_24433,N_24875);
xor UO_563 (O_563,N_22575,N_23155);
and UO_564 (O_564,N_24693,N_24152);
and UO_565 (O_565,N_23260,N_23357);
nor UO_566 (O_566,N_23077,N_24702);
or UO_567 (O_567,N_24380,N_24495);
and UO_568 (O_568,N_24816,N_22022);
nand UO_569 (O_569,N_24873,N_24286);
nor UO_570 (O_570,N_22529,N_23824);
nor UO_571 (O_571,N_23529,N_22114);
nand UO_572 (O_572,N_22339,N_22142);
nand UO_573 (O_573,N_22123,N_23623);
and UO_574 (O_574,N_22459,N_22185);
xor UO_575 (O_575,N_24278,N_23844);
and UO_576 (O_576,N_24010,N_22807);
nand UO_577 (O_577,N_24125,N_23611);
nor UO_578 (O_578,N_24386,N_23897);
xnor UO_579 (O_579,N_24681,N_22765);
or UO_580 (O_580,N_22051,N_24339);
or UO_581 (O_581,N_23585,N_22791);
or UO_582 (O_582,N_21904,N_24508);
xor UO_583 (O_583,N_24820,N_24126);
nor UO_584 (O_584,N_23645,N_22216);
or UO_585 (O_585,N_24823,N_23990);
nand UO_586 (O_586,N_24452,N_22021);
nand UO_587 (O_587,N_24130,N_22750);
and UO_588 (O_588,N_21950,N_24266);
nor UO_589 (O_589,N_22845,N_22639);
or UO_590 (O_590,N_23349,N_22365);
nor UO_591 (O_591,N_23874,N_23711);
nand UO_592 (O_592,N_24303,N_23578);
and UO_593 (O_593,N_23397,N_23302);
xnor UO_594 (O_594,N_24250,N_24121);
xnor UO_595 (O_595,N_22209,N_22795);
or UO_596 (O_596,N_24318,N_24625);
xor UO_597 (O_597,N_24679,N_22226);
nor UO_598 (O_598,N_24507,N_24251);
nand UO_599 (O_599,N_24392,N_22220);
or UO_600 (O_600,N_23177,N_24094);
or UO_601 (O_601,N_22980,N_22928);
nand UO_602 (O_602,N_24822,N_23713);
or UO_603 (O_603,N_24012,N_23008);
and UO_604 (O_604,N_23519,N_24830);
and UO_605 (O_605,N_23163,N_23833);
or UO_606 (O_606,N_24492,N_23791);
nand UO_607 (O_607,N_22959,N_24183);
nand UO_608 (O_608,N_23218,N_22151);
nor UO_609 (O_609,N_24660,N_21952);
nor UO_610 (O_610,N_22971,N_23490);
or UO_611 (O_611,N_23849,N_24580);
nor UO_612 (O_612,N_24659,N_24426);
or UO_613 (O_613,N_22521,N_22158);
xor UO_614 (O_614,N_24808,N_22452);
or UO_615 (O_615,N_23630,N_22916);
nor UO_616 (O_616,N_24421,N_24234);
or UO_617 (O_617,N_23410,N_24793);
and UO_618 (O_618,N_23005,N_24038);
nor UO_619 (O_619,N_22821,N_23939);
nand UO_620 (O_620,N_22826,N_23455);
and UO_621 (O_621,N_23638,N_22268);
or UO_622 (O_622,N_23194,N_24835);
or UO_623 (O_623,N_24154,N_23434);
nor UO_624 (O_624,N_22811,N_22954);
nor UO_625 (O_625,N_24031,N_23468);
nor UO_626 (O_626,N_23170,N_24602);
and UO_627 (O_627,N_23806,N_22248);
nor UO_628 (O_628,N_23221,N_23998);
or UO_629 (O_629,N_23383,N_22382);
nor UO_630 (O_630,N_24888,N_22432);
nor UO_631 (O_631,N_22656,N_23069);
or UO_632 (O_632,N_23129,N_23659);
nand UO_633 (O_633,N_24441,N_24108);
or UO_634 (O_634,N_22251,N_24763);
or UO_635 (O_635,N_22652,N_22476);
or UO_636 (O_636,N_23305,N_22017);
nor UO_637 (O_637,N_24959,N_23472);
nand UO_638 (O_638,N_24554,N_22019);
and UO_639 (O_639,N_22384,N_23836);
or UO_640 (O_640,N_23015,N_22330);
or UO_641 (O_641,N_24546,N_22089);
and UO_642 (O_642,N_23946,N_24933);
or UO_643 (O_643,N_22958,N_22598);
and UO_644 (O_644,N_22407,N_23217);
and UO_645 (O_645,N_22663,N_23066);
or UO_646 (O_646,N_21912,N_23056);
or UO_647 (O_647,N_23574,N_22428);
or UO_648 (O_648,N_23103,N_24648);
nand UO_649 (O_649,N_22257,N_24006);
nand UO_650 (O_650,N_23786,N_23597);
nand UO_651 (O_651,N_23595,N_23167);
and UO_652 (O_652,N_23825,N_24536);
nor UO_653 (O_653,N_22809,N_24264);
nor UO_654 (O_654,N_22465,N_23636);
or UO_655 (O_655,N_23296,N_24676);
nand UO_656 (O_656,N_22208,N_23759);
nor UO_657 (O_657,N_23694,N_23727);
and UO_658 (O_658,N_22680,N_24603);
nand UO_659 (O_659,N_24401,N_23488);
or UO_660 (O_660,N_24867,N_22252);
nor UO_661 (O_661,N_23687,N_22638);
nand UO_662 (O_662,N_23826,N_22833);
nand UO_663 (O_663,N_24337,N_24422);
nand UO_664 (O_664,N_22932,N_22429);
and UO_665 (O_665,N_24751,N_23576);
or UO_666 (O_666,N_24064,N_24828);
and UO_667 (O_667,N_22072,N_22828);
or UO_668 (O_668,N_23341,N_24670);
nand UO_669 (O_669,N_21968,N_24285);
nor UO_670 (O_670,N_22682,N_22295);
nand UO_671 (O_671,N_24886,N_23919);
nor UO_672 (O_672,N_22589,N_23530);
and UO_673 (O_673,N_23847,N_23304);
nor UO_674 (O_674,N_24970,N_23873);
and UO_675 (O_675,N_23316,N_24385);
nand UO_676 (O_676,N_23099,N_24614);
and UO_677 (O_677,N_24296,N_21987);
nand UO_678 (O_678,N_23580,N_23604);
and UO_679 (O_679,N_23427,N_24896);
xnor UO_680 (O_680,N_24464,N_24442);
xnor UO_681 (O_681,N_23553,N_24359);
xor UO_682 (O_682,N_22806,N_24002);
nor UO_683 (O_683,N_22435,N_22712);
nand UO_684 (O_684,N_22235,N_24465);
xnor UO_685 (O_685,N_22412,N_22827);
nor UO_686 (O_686,N_24134,N_22207);
xnor UO_687 (O_687,N_24336,N_23515);
or UO_688 (O_688,N_23186,N_21967);
nand UO_689 (O_689,N_23746,N_24986);
and UO_690 (O_690,N_22477,N_23073);
and UO_691 (O_691,N_22904,N_24456);
and UO_692 (O_692,N_23840,N_22104);
and UO_693 (O_693,N_24329,N_24635);
nor UO_694 (O_694,N_23224,N_24906);
and UO_695 (O_695,N_22499,N_22523);
or UO_696 (O_696,N_23101,N_22873);
nand UO_697 (O_697,N_24518,N_23879);
nor UO_698 (O_698,N_23035,N_23469);
nand UO_699 (O_699,N_23476,N_24300);
or UO_700 (O_700,N_24983,N_23954);
nand UO_701 (O_701,N_21908,N_23068);
and UO_702 (O_702,N_24309,N_24172);
nand UO_703 (O_703,N_21896,N_22202);
nor UO_704 (O_704,N_24992,N_23672);
and UO_705 (O_705,N_22267,N_23610);
and UO_706 (O_706,N_24194,N_23359);
and UO_707 (O_707,N_24074,N_23936);
nand UO_708 (O_708,N_23894,N_22328);
nor UO_709 (O_709,N_23213,N_22605);
nand UO_710 (O_710,N_22596,N_24890);
nand UO_711 (O_711,N_22805,N_22984);
or UO_712 (O_712,N_24953,N_22350);
xor UO_713 (O_713,N_22592,N_22872);
xor UO_714 (O_714,N_24310,N_23815);
or UO_715 (O_715,N_22344,N_23599);
or UO_716 (O_716,N_24241,N_24128);
or UO_717 (O_717,N_24776,N_23665);
nand UO_718 (O_718,N_24785,N_24428);
and UO_719 (O_719,N_21985,N_21974);
and UO_720 (O_720,N_24796,N_22351);
nor UO_721 (O_721,N_22167,N_23709);
nor UO_722 (O_722,N_23398,N_24655);
or UO_723 (O_723,N_24211,N_24461);
or UO_724 (O_724,N_23102,N_23615);
and UO_725 (O_725,N_23249,N_23588);
nor UO_726 (O_726,N_23679,N_22588);
nand UO_727 (O_727,N_24965,N_22934);
nand UO_728 (O_728,N_23042,N_24493);
or UO_729 (O_729,N_23038,N_22436);
or UO_730 (O_730,N_24738,N_22891);
or UO_731 (O_731,N_22718,N_24801);
nor UO_732 (O_732,N_22889,N_23450);
and UO_733 (O_733,N_23744,N_23771);
or UO_734 (O_734,N_24239,N_23209);
and UO_735 (O_735,N_24572,N_23570);
nor UO_736 (O_736,N_24916,N_24171);
nand UO_737 (O_737,N_24736,N_23503);
or UO_738 (O_738,N_24469,N_22254);
nor UO_739 (O_739,N_24675,N_23461);
nor UO_740 (O_740,N_23018,N_24236);
xnor UO_741 (O_741,N_23969,N_22166);
nor UO_742 (O_742,N_22385,N_22616);
nor UO_743 (O_743,N_23887,N_24976);
nor UO_744 (O_744,N_23823,N_23513);
or UO_745 (O_745,N_24430,N_24934);
nor UO_746 (O_746,N_23159,N_21997);
or UO_747 (O_747,N_21929,N_23632);
and UO_748 (O_748,N_24199,N_22558);
nand UO_749 (O_749,N_23545,N_23910);
and UO_750 (O_750,N_24044,N_24936);
and UO_751 (O_751,N_23321,N_23674);
nand UO_752 (O_752,N_23372,N_23232);
nand UO_753 (O_753,N_21955,N_22620);
nand UO_754 (O_754,N_23782,N_23596);
and UO_755 (O_755,N_24246,N_24574);
nor UO_756 (O_756,N_23318,N_23266);
or UO_757 (O_757,N_24210,N_24853);
or UO_758 (O_758,N_24674,N_24556);
and UO_759 (O_759,N_24332,N_22352);
nand UO_760 (O_760,N_24876,N_22150);
nand UO_761 (O_761,N_23007,N_22399);
or UO_762 (O_762,N_23697,N_24937);
and UO_763 (O_763,N_24087,N_23960);
and UO_764 (O_764,N_23681,N_23547);
nand UO_765 (O_765,N_23938,N_23423);
and UO_766 (O_766,N_24458,N_24383);
nor UO_767 (O_767,N_23703,N_24274);
or UO_768 (O_768,N_24136,N_24078);
or UO_769 (O_769,N_24201,N_22527);
xnor UO_770 (O_770,N_24345,N_22668);
and UO_771 (O_771,N_23945,N_23310);
or UO_772 (O_772,N_24750,N_24040);
or UO_773 (O_773,N_24124,N_24208);
or UO_774 (O_774,N_24995,N_22119);
nand UO_775 (O_775,N_22160,N_24283);
nand UO_776 (O_776,N_22946,N_24665);
nand UO_777 (O_777,N_22451,N_22948);
nand UO_778 (O_778,N_23613,N_23906);
nand UO_779 (O_779,N_22128,N_22942);
and UO_780 (O_780,N_24961,N_22981);
xor UO_781 (O_781,N_24325,N_23878);
nand UO_782 (O_782,N_24865,N_24667);
nor UO_783 (O_783,N_23118,N_24045);
nor UO_784 (O_784,N_24018,N_24901);
nor UO_785 (O_785,N_23923,N_23250);
or UO_786 (O_786,N_24579,N_23796);
xor UO_787 (O_787,N_21927,N_24672);
nor UO_788 (O_788,N_23140,N_22337);
xor UO_789 (O_789,N_23508,N_24315);
and UO_790 (O_790,N_24568,N_22417);
nand UO_791 (O_791,N_23058,N_23214);
nand UO_792 (O_792,N_24815,N_22788);
nor UO_793 (O_793,N_24351,N_22863);
xnor UO_794 (O_794,N_23725,N_23800);
nand UO_795 (O_795,N_22146,N_24138);
nor UO_796 (O_796,N_23858,N_22390);
or UO_797 (O_797,N_23405,N_22321);
and UO_798 (O_798,N_23752,N_22719);
nor UO_799 (O_799,N_22947,N_24856);
or UO_800 (O_800,N_22200,N_22912);
nor UO_801 (O_801,N_23351,N_24578);
or UO_802 (O_802,N_21925,N_22600);
nor UO_803 (O_803,N_22549,N_23336);
or UO_804 (O_804,N_24140,N_23500);
nor UO_805 (O_805,N_23509,N_22475);
or UO_806 (O_806,N_22534,N_22566);
xor UO_807 (O_807,N_23587,N_22120);
nand UO_808 (O_808,N_24197,N_22420);
nand UO_809 (O_809,N_22554,N_22617);
nor UO_810 (O_810,N_23775,N_24055);
nor UO_811 (O_811,N_23735,N_22738);
and UO_812 (O_812,N_24445,N_21890);
nand UO_813 (O_813,N_22876,N_23700);
nand UO_814 (O_814,N_22410,N_23774);
nor UO_815 (O_815,N_23147,N_23072);
nand UO_816 (O_816,N_22561,N_24477);
nor UO_817 (O_817,N_24740,N_23668);
or UO_818 (O_818,N_23090,N_23977);
nor UO_819 (O_819,N_24167,N_24993);
nand UO_820 (O_820,N_24233,N_24855);
xnor UO_821 (O_821,N_23556,N_23811);
nand UO_822 (O_822,N_22783,N_23340);
nor UO_823 (O_823,N_24498,N_22586);
or UO_824 (O_824,N_24429,N_22053);
or UO_825 (O_825,N_22786,N_24731);
and UO_826 (O_826,N_22522,N_22885);
and UO_827 (O_827,N_21980,N_24284);
and UO_828 (O_828,N_22644,N_22665);
nand UO_829 (O_829,N_22004,N_24557);
nor UO_830 (O_830,N_22091,N_22097);
nor UO_831 (O_831,N_22127,N_24804);
and UO_832 (O_832,N_22362,N_22709);
or UO_833 (O_833,N_24192,N_23413);
and UO_834 (O_834,N_22603,N_23839);
nor UO_835 (O_835,N_24642,N_22264);
and UO_836 (O_836,N_22988,N_23997);
xnor UO_837 (O_837,N_23653,N_22346);
nor UO_838 (O_838,N_24686,N_21926);
nor UO_839 (O_839,N_24389,N_23643);
nor UO_840 (O_840,N_24067,N_23451);
and UO_841 (O_841,N_21909,N_23264);
or UO_842 (O_842,N_22951,N_22088);
nand UO_843 (O_843,N_22993,N_24071);
nor UO_844 (O_844,N_22537,N_23622);
nand UO_845 (O_845,N_22509,N_22908);
nor UO_846 (O_846,N_23589,N_24613);
or UO_847 (O_847,N_24914,N_22573);
nand UO_848 (O_848,N_22520,N_23590);
nand UO_849 (O_849,N_24483,N_24169);
or UO_850 (O_850,N_22370,N_22291);
nand UO_851 (O_851,N_23275,N_24478);
nand UO_852 (O_852,N_24699,N_23401);
nor UO_853 (O_853,N_22073,N_22336);
nor UO_854 (O_854,N_23743,N_24275);
nand UO_855 (O_855,N_22838,N_22555);
nand UO_856 (O_856,N_24257,N_24646);
xor UO_857 (O_857,N_22246,N_21995);
or UO_858 (O_858,N_22856,N_22846);
nand UO_859 (O_859,N_24034,N_23854);
xnor UO_860 (O_860,N_23685,N_23557);
nor UO_861 (O_861,N_24215,N_23287);
or UO_862 (O_862,N_24202,N_24880);
nor UO_863 (O_863,N_23388,N_22504);
nand UO_864 (O_864,N_23207,N_23442);
nor UO_865 (O_865,N_24846,N_23430);
xnor UO_866 (O_866,N_22354,N_22376);
and UO_867 (O_867,N_23925,N_23060);
or UO_868 (O_868,N_24547,N_22822);
nand UO_869 (O_869,N_22488,N_24119);
nand UO_870 (O_870,N_23011,N_23911);
or UO_871 (O_871,N_23429,N_22287);
or UO_872 (O_872,N_23271,N_22999);
nand UO_873 (O_873,N_24265,N_24915);
xnor UO_874 (O_874,N_23191,N_22764);
or UO_875 (O_875,N_23444,N_24139);
nor UO_876 (O_876,N_21951,N_23724);
or UO_877 (O_877,N_23577,N_24271);
nand UO_878 (O_878,N_21876,N_22446);
and UO_879 (O_879,N_24021,N_22197);
and UO_880 (O_880,N_24057,N_24656);
or UO_881 (O_881,N_21875,N_22347);
nor UO_882 (O_882,N_23932,N_22271);
and UO_883 (O_883,N_22101,N_22562);
xor UO_884 (O_884,N_24994,N_24513);
xor UO_885 (O_885,N_24752,N_23778);
nor UO_886 (O_886,N_22710,N_23642);
or UO_887 (O_887,N_24252,N_22215);
nand UO_888 (O_888,N_22177,N_24160);
or UO_889 (O_889,N_23363,N_21913);
nand UO_890 (O_890,N_22965,N_22374);
nand UO_891 (O_891,N_24077,N_22324);
and UO_892 (O_892,N_22886,N_24368);
nand UO_893 (O_893,N_24797,N_24084);
nand UO_894 (O_894,N_22395,N_23922);
nand UO_895 (O_895,N_24297,N_23649);
or UO_896 (O_896,N_22266,N_24909);
nor UO_897 (O_897,N_23964,N_22705);
and UO_898 (O_898,N_22675,N_23141);
and UO_899 (O_899,N_22242,N_22361);
or UO_900 (O_900,N_22645,N_24327);
nor UO_901 (O_901,N_21878,N_22624);
and UO_902 (O_902,N_22026,N_22141);
nor UO_903 (O_903,N_23390,N_23003);
nor UO_904 (O_904,N_24925,N_22396);
nor UO_905 (O_905,N_23764,N_22316);
nand UO_906 (O_906,N_24435,N_22975);
xor UO_907 (O_907,N_21923,N_24227);
and UO_908 (O_908,N_24831,N_22356);
or UO_909 (O_909,N_23255,N_23995);
or UO_910 (O_910,N_24891,N_23445);
and UO_911 (O_911,N_22224,N_24519);
and UO_912 (O_912,N_22610,N_21976);
nor UO_913 (O_913,N_22781,N_22441);
and UO_914 (O_914,N_22888,N_22836);
nor UO_915 (O_915,N_23009,N_22770);
and UO_916 (O_916,N_22322,N_23356);
nor UO_917 (O_917,N_24599,N_23467);
or UO_918 (O_918,N_21935,N_23021);
and UO_919 (O_919,N_22100,N_21993);
nor UO_920 (O_920,N_23619,N_24417);
nand UO_921 (O_921,N_22701,N_23432);
or UO_922 (O_922,N_24612,N_22233);
nor UO_923 (O_923,N_24484,N_22865);
nand UO_924 (O_924,N_24326,N_24181);
or UO_925 (O_925,N_24109,N_23115);
or UO_926 (O_926,N_24824,N_22001);
nor UO_927 (O_927,N_22655,N_21910);
xor UO_928 (O_928,N_21917,N_24618);
nand UO_929 (O_929,N_22152,N_24370);
or UO_930 (O_930,N_23301,N_24276);
nand UO_931 (O_931,N_22899,N_24179);
xnor UO_932 (O_932,N_22727,N_24511);
and UO_933 (O_933,N_23127,N_23384);
and UO_934 (O_934,N_23220,N_23303);
nor UO_935 (O_935,N_23924,N_22335);
xnor UO_936 (O_936,N_22013,N_23862);
nor UO_937 (O_937,N_22148,N_21884);
or UO_938 (O_938,N_24885,N_22038);
nor UO_939 (O_939,N_24059,N_22506);
nor UO_940 (O_940,N_23712,N_24577);
and UO_941 (O_941,N_24616,N_23655);
or UO_942 (O_942,N_24932,N_23082);
nor UO_943 (O_943,N_21879,N_24193);
or UO_944 (O_944,N_21887,N_23358);
nor UO_945 (O_945,N_22547,N_23860);
nand UO_946 (O_946,N_24409,N_22018);
nor UO_947 (O_947,N_24680,N_22298);
or UO_948 (O_948,N_24198,N_24780);
or UO_949 (O_949,N_22221,N_23640);
or UO_950 (O_950,N_24567,N_23884);
or UO_951 (O_951,N_24592,N_22259);
nor UO_952 (O_952,N_24773,N_23993);
nand UO_953 (O_953,N_24506,N_22117);
and UO_954 (O_954,N_22389,N_24798);
nor UO_955 (O_955,N_23706,N_24273);
and UO_956 (O_956,N_21946,N_22681);
or UO_957 (O_957,N_23055,N_24905);
or UO_958 (O_958,N_22995,N_23494);
or UO_959 (O_959,N_23484,N_22103);
nor UO_960 (O_960,N_24741,N_23166);
and UO_961 (O_961,N_21979,N_22844);
nor UO_962 (O_962,N_22405,N_22802);
nand UO_963 (O_963,N_24427,N_24413);
nand UO_964 (O_964,N_23223,N_24912);
xnor UO_965 (O_965,N_23584,N_24003);
and UO_966 (O_966,N_24313,N_22456);
or UO_967 (O_967,N_22363,N_24229);
or UO_968 (O_968,N_24945,N_23971);
xnor UO_969 (O_969,N_22749,N_23043);
or UO_970 (O_970,N_24761,N_23606);
and UO_971 (O_971,N_22776,N_22060);
or UO_972 (O_972,N_22910,N_21991);
or UO_973 (O_973,N_23560,N_23644);
and UO_974 (O_974,N_22078,N_22099);
or UO_975 (O_975,N_24024,N_22069);
xor UO_976 (O_976,N_23000,N_24520);
and UO_977 (O_977,N_23165,N_23563);
and UO_978 (O_978,N_23306,N_23767);
and UO_979 (O_979,N_22538,N_23091);
or UO_980 (O_980,N_21990,N_24245);
or UO_981 (O_981,N_24166,N_23895);
nor UO_982 (O_982,N_24649,N_23169);
or UO_983 (O_983,N_24425,N_24951);
nor UO_984 (O_984,N_24834,N_22926);
xor UO_985 (O_985,N_21916,N_23705);
nand UO_986 (O_986,N_22955,N_23242);
nand UO_987 (O_987,N_22569,N_22642);
or UO_988 (O_988,N_24468,N_23498);
or UO_989 (O_989,N_23404,N_22463);
nor UO_990 (O_990,N_23376,N_22875);
or UO_991 (O_991,N_23109,N_22106);
nand UO_992 (O_992,N_24357,N_24571);
and UO_993 (O_993,N_24922,N_22585);
nor UO_994 (O_994,N_22796,N_22129);
nand UO_995 (O_995,N_23136,N_21936);
nand UO_996 (O_996,N_22338,N_22397);
nand UO_997 (O_997,N_23527,N_23210);
nor UO_998 (O_998,N_22180,N_22478);
xnor UO_999 (O_999,N_23268,N_23691);
or UO_1000 (O_1000,N_23454,N_22736);
nor UO_1001 (O_1001,N_22210,N_24605);
and UO_1002 (O_1002,N_23801,N_23870);
or UO_1003 (O_1003,N_24052,N_22461);
nand UO_1004 (O_1004,N_23544,N_23092);
and UO_1005 (O_1005,N_22877,N_22464);
or UO_1006 (O_1006,N_22244,N_22801);
or UO_1007 (O_1007,N_23493,N_22419);
nand UO_1008 (O_1008,N_23662,N_22572);
nor UO_1009 (O_1009,N_22966,N_24053);
or UO_1010 (O_1010,N_23719,N_22532);
xnor UO_1011 (O_1011,N_24946,N_24844);
and UO_1012 (O_1012,N_22468,N_23267);
or UO_1013 (O_1013,N_24287,N_23809);
nand UO_1014 (O_1014,N_24131,N_23710);
xor UO_1015 (O_1015,N_23565,N_22857);
nor UO_1016 (O_1016,N_24716,N_23837);
nand UO_1017 (O_1017,N_23265,N_22678);
or UO_1018 (O_1018,N_23176,N_23626);
xnor UO_1019 (O_1019,N_24290,N_22963);
or UO_1020 (O_1020,N_22294,N_23050);
xnor UO_1021 (O_1021,N_22556,N_24482);
or UO_1022 (O_1022,N_23551,N_23300);
xnor UO_1023 (O_1023,N_23276,N_24692);
and UO_1024 (O_1024,N_24432,N_24320);
and UO_1025 (O_1025,N_22777,N_23620);
or UO_1026 (O_1026,N_24219,N_23293);
or UO_1027 (O_1027,N_23385,N_24046);
nand UO_1028 (O_1028,N_21939,N_22010);
or UO_1029 (O_1029,N_24525,N_23437);
nor UO_1030 (O_1030,N_24772,N_24120);
nor UO_1031 (O_1031,N_24115,N_22037);
nand UO_1032 (O_1032,N_23253,N_22191);
xnor UO_1033 (O_1033,N_24117,N_24609);
and UO_1034 (O_1034,N_22890,N_24620);
xor UO_1035 (O_1035,N_22308,N_22469);
and UO_1036 (O_1036,N_22327,N_22095);
xor UO_1037 (O_1037,N_23904,N_24177);
or UO_1038 (O_1038,N_24907,N_22653);
nor UO_1039 (O_1039,N_23842,N_23259);
or UO_1040 (O_1040,N_23618,N_21883);
nor UO_1041 (O_1041,N_22402,N_24291);
nand UO_1042 (O_1042,N_24240,N_22332);
and UO_1043 (O_1043,N_22240,N_23228);
nor UO_1044 (O_1044,N_24950,N_24719);
nand UO_1045 (O_1045,N_23187,N_22799);
xor UO_1046 (O_1046,N_23006,N_24377);
and UO_1047 (O_1047,N_23192,N_23324);
nand UO_1048 (O_1048,N_22755,N_23908);
or UO_1049 (O_1049,N_22082,N_23497);
and UO_1050 (O_1050,N_22594,N_24552);
or UO_1051 (O_1051,N_22670,N_22992);
or UO_1052 (O_1052,N_23534,N_24366);
xnor UO_1053 (O_1053,N_24636,N_24957);
or UO_1054 (O_1054,N_22241,N_22031);
xnor UO_1055 (O_1055,N_23762,N_22373);
nor UO_1056 (O_1056,N_22994,N_22272);
nand UO_1057 (O_1057,N_23269,N_22449);
nor UO_1058 (O_1058,N_24105,N_22081);
nand UO_1059 (O_1059,N_24293,N_24393);
or UO_1060 (O_1060,N_24539,N_22861);
nor UO_1061 (O_1061,N_24346,N_22970);
nor UO_1062 (O_1062,N_24799,N_24305);
nand UO_1063 (O_1063,N_23200,N_24342);
nand UO_1064 (O_1064,N_22126,N_24516);
and UO_1065 (O_1065,N_22408,N_23052);
nor UO_1066 (O_1066,N_24324,N_22501);
or UO_1067 (O_1067,N_22062,N_24817);
or UO_1068 (O_1068,N_23227,N_22913);
nand UO_1069 (O_1069,N_23986,N_23375);
nand UO_1070 (O_1070,N_22144,N_22400);
nand UO_1071 (O_1071,N_23617,N_24301);
and UO_1072 (O_1072,N_23591,N_24129);
or UO_1073 (O_1073,N_23048,N_23252);
nand UO_1074 (O_1074,N_24367,N_22535);
nor UO_1075 (O_1075,N_22163,N_24989);
nor UO_1076 (O_1076,N_23203,N_23651);
nor UO_1077 (O_1077,N_24715,N_24777);
or UO_1078 (O_1078,N_23374,N_22657);
nor UO_1079 (O_1079,N_24196,N_22245);
nand UO_1080 (O_1080,N_24727,N_23978);
nand UO_1081 (O_1081,N_23145,N_24042);
nand UO_1082 (O_1082,N_23272,N_22571);
and UO_1083 (O_1083,N_23134,N_24165);
or UO_1084 (O_1084,N_22909,N_24080);
nand UO_1085 (O_1085,N_23582,N_22192);
and UO_1086 (O_1086,N_24742,N_22717);
and UO_1087 (O_1087,N_24878,N_23799);
nor UO_1088 (O_1088,N_23748,N_23846);
and UO_1089 (O_1089,N_22688,N_22329);
nor UO_1090 (O_1090,N_24666,N_22831);
nand UO_1091 (O_1091,N_22378,N_22398);
and UO_1092 (O_1092,N_23037,N_23354);
and UO_1093 (O_1093,N_22747,N_22893);
xnor UO_1094 (O_1094,N_22698,N_24689);
or UO_1095 (O_1095,N_23173,N_21962);
nand UO_1096 (O_1096,N_23353,N_24759);
nand UO_1097 (O_1097,N_22567,N_24356);
nand UO_1098 (O_1098,N_24730,N_24155);
nor UO_1099 (O_1099,N_23284,N_24382);
nand UO_1100 (O_1100,N_24280,N_23004);
or UO_1101 (O_1101,N_23462,N_22565);
nor UO_1102 (O_1102,N_21978,N_23893);
nor UO_1103 (O_1103,N_24025,N_23433);
and UO_1104 (O_1104,N_23788,N_23084);
and UO_1105 (O_1105,N_23331,N_24712);
or UO_1106 (O_1106,N_23814,N_24307);
nand UO_1107 (O_1107,N_23784,N_22945);
or UO_1108 (O_1108,N_23112,N_22724);
or UO_1109 (O_1109,N_24133,N_22285);
and UO_1110 (O_1110,N_21888,N_22591);
nand UO_1111 (O_1111,N_24376,N_22046);
and UO_1112 (O_1112,N_21996,N_24407);
nor UO_1113 (O_1113,N_23032,N_22364);
and UO_1114 (O_1114,N_23913,N_23237);
nand UO_1115 (O_1115,N_24583,N_24447);
nand UO_1116 (O_1116,N_21945,N_23263);
nand UO_1117 (O_1117,N_24852,N_24362);
or UO_1118 (O_1118,N_21882,N_22284);
nand UO_1119 (O_1119,N_23128,N_23346);
nor UO_1120 (O_1120,N_22898,N_22145);
nor UO_1121 (O_1121,N_22462,N_24729);
nand UO_1122 (O_1122,N_22584,N_24106);
and UO_1123 (O_1123,N_23516,N_24569);
nor UO_1124 (O_1124,N_24654,N_23419);
and UO_1125 (O_1125,N_24446,N_22490);
nor UO_1126 (O_1126,N_22546,N_23348);
nand UO_1127 (O_1127,N_23987,N_22474);
nand UO_1128 (O_1128,N_22274,N_21958);
nor UO_1129 (O_1129,N_22472,N_23024);
or UO_1130 (O_1130,N_22626,N_24615);
xnor UO_1131 (O_1131,N_23482,N_23769);
nor UO_1132 (O_1132,N_23892,N_23813);
nor UO_1133 (O_1133,N_24509,N_23201);
and UO_1134 (O_1134,N_24643,N_23029);
nor UO_1135 (O_1135,N_23244,N_24581);
nand UO_1136 (O_1136,N_24187,N_22007);
xor UO_1137 (O_1137,N_24114,N_21994);
or UO_1138 (O_1138,N_23117,N_23046);
xnor UO_1139 (O_1139,N_24737,N_22135);
or UO_1140 (O_1140,N_23984,N_24340);
nor UO_1141 (O_1141,N_23317,N_24931);
or UO_1142 (O_1142,N_24941,N_24020);
or UO_1143 (O_1143,N_24471,N_22737);
nor UO_1144 (O_1144,N_22611,N_22997);
nand UO_1145 (O_1145,N_24810,N_22289);
and UO_1146 (O_1146,N_24358,N_22792);
and UO_1147 (O_1147,N_24921,N_22540);
and UO_1148 (O_1148,N_24882,N_23093);
and UO_1149 (O_1149,N_24341,N_23541);
nor UO_1150 (O_1150,N_22672,N_22253);
nand UO_1151 (O_1151,N_22702,N_24713);
or UO_1152 (O_1152,N_24462,N_22696);
nand UO_1153 (O_1153,N_23598,N_24641);
and UO_1154 (O_1154,N_24269,N_23828);
nand UO_1155 (O_1155,N_24778,N_22869);
nand UO_1156 (O_1156,N_22258,N_23639);
or UO_1157 (O_1157,N_23135,N_24898);
xor UO_1158 (O_1158,N_24047,N_21889);
nor UO_1159 (O_1159,N_24149,N_22133);
or UO_1160 (O_1160,N_24424,N_23313);
xnor UO_1161 (O_1161,N_24086,N_23779);
xnor UO_1162 (O_1162,N_23930,N_23291);
xor UO_1163 (O_1163,N_24260,N_23254);
xor UO_1164 (O_1164,N_23807,N_22723);
xor UO_1165 (O_1165,N_24150,N_24859);
and UO_1166 (O_1166,N_23822,N_24041);
nor UO_1167 (O_1167,N_22998,N_23510);
nand UO_1168 (O_1168,N_21992,N_24617);
or UO_1169 (O_1169,N_23295,N_23572);
nor UO_1170 (O_1170,N_22607,N_24857);
nand UO_1171 (O_1171,N_24929,N_23051);
nor UO_1172 (O_1172,N_23766,N_24549);
or UO_1173 (O_1173,N_22576,N_23696);
nor UO_1174 (O_1174,N_24622,N_22355);
and UO_1175 (O_1175,N_22650,N_24779);
or UO_1176 (O_1176,N_24850,N_23934);
nand UO_1177 (O_1177,N_22983,N_22406);
and UO_1178 (O_1178,N_23126,N_22793);
nand UO_1179 (O_1179,N_24924,N_24353);
nand UO_1180 (O_1180,N_24626,N_24544);
nor UO_1181 (O_1181,N_23802,N_24701);
and UO_1182 (O_1182,N_22165,N_23471);
nand UO_1183 (O_1183,N_24532,N_22108);
and UO_1184 (O_1184,N_21907,N_22250);
nor UO_1185 (O_1185,N_24978,N_23942);
nand UO_1186 (O_1186,N_22858,N_24072);
nor UO_1187 (O_1187,N_22779,N_22333);
nand UO_1188 (O_1188,N_23927,N_22261);
nand UO_1189 (O_1189,N_22502,N_22057);
or UO_1190 (O_1190,N_24292,N_22211);
and UO_1191 (O_1191,N_23944,N_24918);
nor UO_1192 (O_1192,N_24948,N_22122);
and UO_1193 (O_1193,N_24281,N_23449);
or UO_1194 (O_1194,N_24312,N_21920);
nor UO_1195 (O_1195,N_22732,N_24013);
and UO_1196 (O_1196,N_23338,N_22895);
nor UO_1197 (O_1197,N_24595,N_24697);
and UO_1198 (O_1198,N_24406,N_22748);
xnor UO_1199 (O_1199,N_24404,N_21931);
and UO_1200 (O_1200,N_24606,N_24223);
nor UO_1201 (O_1201,N_22143,N_21892);
nand UO_1202 (O_1202,N_24981,N_23074);
nor UO_1203 (O_1203,N_22923,N_24559);
or UO_1204 (O_1204,N_22198,N_23804);
or UO_1205 (O_1205,N_22323,N_24892);
and UO_1206 (O_1206,N_22512,N_22733);
or UO_1207 (O_1207,N_23754,N_24861);
nand UO_1208 (O_1208,N_24695,N_23496);
xor UO_1209 (O_1209,N_23453,N_24017);
xor UO_1210 (O_1210,N_22479,N_24688);
nor UO_1211 (O_1211,N_23474,N_23033);
and UO_1212 (O_1212,N_23095,N_24437);
nor UO_1213 (O_1213,N_24963,N_24576);
nor UO_1214 (O_1214,N_21880,N_22282);
nand UO_1215 (O_1215,N_23929,N_22830);
and UO_1216 (O_1216,N_24814,N_23988);
and UO_1217 (O_1217,N_24783,N_23728);
nand UO_1218 (O_1218,N_22181,N_22853);
xor UO_1219 (O_1219,N_22660,N_24316);
and UO_1220 (O_1220,N_24102,N_22915);
and UO_1221 (O_1221,N_23465,N_24543);
nand UO_1222 (O_1222,N_22102,N_22884);
or UO_1223 (O_1223,N_24440,N_22080);
xor UO_1224 (O_1224,N_24485,N_24504);
and UO_1225 (O_1225,N_24107,N_24923);
nand UO_1226 (O_1226,N_21943,N_24739);
nor UO_1227 (O_1227,N_23282,N_22896);
or UO_1228 (O_1228,N_22722,N_24186);
or UO_1229 (O_1229,N_23693,N_23751);
nor UO_1230 (O_1230,N_24302,N_22637);
nor UO_1231 (O_1231,N_23658,N_24813);
nor UO_1232 (O_1232,N_23817,N_24997);
nor UO_1233 (O_1233,N_23504,N_24530);
and UO_1234 (O_1234,N_21881,N_24608);
or UO_1235 (O_1235,N_22358,N_24270);
or UO_1236 (O_1236,N_24467,N_22125);
nor UO_1237 (O_1237,N_24436,N_23763);
or UO_1238 (O_1238,N_23583,N_23216);
nand UO_1239 (O_1239,N_23245,N_22577);
and UO_1240 (O_1240,N_24919,N_23635);
or UO_1241 (O_1241,N_23912,N_24913);
nand UO_1242 (O_1242,N_22487,N_22557);
xor UO_1243 (O_1243,N_24864,N_22659);
nand UO_1244 (O_1244,N_24756,N_21999);
nand UO_1245 (O_1245,N_24343,N_24148);
or UO_1246 (O_1246,N_23114,N_24975);
or UO_1247 (O_1247,N_21973,N_23845);
and UO_1248 (O_1248,N_24696,N_22414);
and UO_1249 (O_1249,N_24444,N_24938);
xnor UO_1250 (O_1250,N_23531,N_23392);
or UO_1251 (O_1251,N_22635,N_22866);
nand UO_1252 (O_1252,N_23320,N_24728);
and UO_1253 (O_1253,N_23812,N_24475);
nand UO_1254 (O_1254,N_22444,N_24039);
or UO_1255 (O_1255,N_23380,N_22302);
xor UO_1256 (O_1256,N_24973,N_22834);
nand UO_1257 (O_1257,N_23838,N_23790);
nand UO_1258 (O_1258,N_21898,N_21963);
nand UO_1259 (O_1259,N_23464,N_23738);
and UO_1260 (O_1260,N_22510,N_24238);
or UO_1261 (O_1261,N_23158,N_22905);
and UO_1262 (O_1262,N_24061,N_23373);
and UO_1263 (O_1263,N_22345,N_22545);
and UO_1264 (O_1264,N_24794,N_22132);
nand UO_1265 (O_1265,N_23119,N_24092);
or UO_1266 (O_1266,N_24137,N_22270);
or UO_1267 (O_1267,N_22301,N_23855);
and UO_1268 (O_1268,N_24942,N_23967);
nand UO_1269 (O_1269,N_24920,N_24037);
and UO_1270 (O_1270,N_22359,N_21899);
xor UO_1271 (O_1271,N_24416,N_22393);
nor UO_1272 (O_1272,N_22590,N_23943);
nor UO_1273 (O_1273,N_22867,N_24881);
xor UO_1274 (O_1274,N_22379,N_23143);
or UO_1275 (O_1275,N_24147,N_22343);
xor UO_1276 (O_1276,N_24839,N_22303);
xor UO_1277 (O_1277,N_22533,N_22136);
nand UO_1278 (O_1278,N_22087,N_23025);
and UO_1279 (O_1279,N_23729,N_24244);
nand UO_1280 (O_1280,N_24940,N_24414);
and UO_1281 (O_1281,N_23131,N_22187);
and UO_1282 (O_1282,N_23561,N_24553);
and UO_1283 (O_1283,N_22231,N_23718);
and UO_1284 (O_1284,N_22902,N_23308);
nor UO_1285 (O_1285,N_23770,N_24146);
nor UO_1286 (O_1286,N_22320,N_24157);
nand UO_1287 (O_1287,N_24700,N_22883);
xor UO_1288 (O_1288,N_22794,N_22304);
or UO_1289 (O_1289,N_21981,N_22924);
or UO_1290 (O_1290,N_22841,N_24897);
nand UO_1291 (O_1291,N_23714,N_22731);
nand UO_1292 (O_1292,N_22228,N_22860);
and UO_1293 (O_1293,N_24535,N_22901);
or UO_1294 (O_1294,N_22628,N_23379);
or UO_1295 (O_1295,N_23981,N_24964);
or UO_1296 (O_1296,N_23344,N_23104);
nand UO_1297 (O_1297,N_22319,N_24631);
and UO_1298 (O_1298,N_22879,N_24708);
and UO_1299 (O_1299,N_23517,N_24966);
nand UO_1300 (O_1300,N_24634,N_23609);
or UO_1301 (O_1301,N_24352,N_24795);
and UO_1302 (O_1302,N_23962,N_24410);
nand UO_1303 (O_1303,N_21972,N_24259);
and UO_1304 (O_1304,N_24016,N_22040);
nor UO_1305 (O_1305,N_24364,N_23624);
and UO_1306 (O_1306,N_23540,N_24365);
and UO_1307 (O_1307,N_24344,N_21982);
nand UO_1308 (O_1308,N_24807,N_23463);
or UO_1309 (O_1309,N_22184,N_23616);
nand UO_1310 (O_1310,N_22377,N_23160);
and UO_1311 (O_1311,N_22061,N_24220);
or UO_1312 (O_1312,N_21932,N_24499);
nor UO_1313 (O_1313,N_23017,N_23896);
and UO_1314 (O_1314,N_23723,N_22075);
nand UO_1315 (O_1315,N_24225,N_22426);
and UO_1316 (O_1316,N_24438,N_23733);
or UO_1317 (O_1317,N_23586,N_24178);
xnor UO_1318 (O_1318,N_23204,N_23511);
nor UO_1319 (O_1319,N_22508,N_22641);
nor UO_1320 (O_1320,N_23366,N_24677);
nand UO_1321 (O_1321,N_23708,N_24443);
nor UO_1322 (O_1322,N_22550,N_23146);
nor UO_1323 (O_1323,N_21901,N_22434);
and UO_1324 (O_1324,N_24917,N_22388);
nor UO_1325 (O_1325,N_23153,N_24758);
nand UO_1326 (O_1326,N_24032,N_23426);
or UO_1327 (O_1327,N_22852,N_23980);
or UO_1328 (O_1328,N_24127,N_23970);
and UO_1329 (O_1329,N_22939,N_24405);
nand UO_1330 (O_1330,N_23612,N_22921);
or UO_1331 (O_1331,N_22808,N_22153);
nand UO_1332 (O_1332,N_22416,N_24083);
or UO_1333 (O_1333,N_23036,N_22067);
nand UO_1334 (O_1334,N_22671,N_24510);
xor UO_1335 (O_1335,N_23345,N_24573);
nand UO_1336 (O_1336,N_23677,N_22758);
nand UO_1337 (O_1337,N_24894,N_23428);
nor UO_1338 (O_1338,N_24753,N_23054);
or UO_1339 (O_1339,N_22424,N_22486);
nand UO_1340 (O_1340,N_22745,N_22194);
and UO_1341 (O_1341,N_22631,N_23466);
nand UO_1342 (O_1342,N_22551,N_22634);
or UO_1343 (O_1343,N_22190,N_23991);
nor UO_1344 (O_1344,N_23414,N_23961);
and UO_1345 (O_1345,N_23716,N_23085);
nor UO_1346 (O_1346,N_24971,N_24048);
or UO_1347 (O_1347,N_24593,N_24158);
nand UO_1348 (O_1348,N_24939,N_23298);
or UO_1349 (O_1349,N_22288,N_24500);
nand UO_1350 (O_1350,N_24068,N_23422);
or UO_1351 (O_1351,N_24277,N_24889);
and UO_1352 (O_1352,N_23684,N_23061);
and UO_1353 (O_1353,N_23857,N_23365);
nor UO_1354 (O_1354,N_23676,N_23666);
nor UO_1355 (O_1355,N_24262,N_23850);
or UO_1356 (O_1356,N_24030,N_24910);
and UO_1357 (O_1357,N_21895,N_23044);
nand UO_1358 (O_1358,N_22140,N_24575);
or UO_1359 (O_1359,N_24991,N_24735);
nand UO_1360 (O_1360,N_22759,N_23319);
and UO_1361 (O_1361,N_22247,N_23149);
xor UO_1362 (O_1362,N_23185,N_24540);
nand UO_1363 (O_1363,N_23486,N_22989);
xor UO_1364 (O_1364,N_22056,N_23914);
or UO_1365 (O_1365,N_24168,N_23138);
and UO_1366 (O_1366,N_24690,N_24163);
nand UO_1367 (O_1367,N_24191,N_23905);
nor UO_1368 (O_1368,N_22714,N_22880);
or UO_1369 (O_1369,N_24550,N_22483);
xnor UO_1370 (O_1370,N_22715,N_21965);
nor UO_1371 (O_1371,N_24985,N_23387);
nor UO_1372 (O_1372,N_22170,N_22752);
nand UO_1373 (O_1373,N_24800,N_24668);
or UO_1374 (O_1374,N_24247,N_22011);
nor UO_1375 (O_1375,N_22612,N_22720);
nor UO_1376 (O_1376,N_22034,N_23020);
nand UO_1377 (O_1377,N_23139,N_22066);
or UO_1378 (O_1378,N_22000,N_22578);
or UO_1379 (O_1379,N_24900,N_24694);
and UO_1380 (O_1380,N_24195,N_24893);
nand UO_1381 (O_1381,N_23377,N_22134);
or UO_1382 (O_1382,N_24818,N_23543);
or UO_1383 (O_1383,N_23795,N_24248);
nand UO_1384 (O_1384,N_23959,N_22848);
nand UO_1385 (O_1385,N_24298,N_22987);
or UO_1386 (O_1386,N_22494,N_24457);
nor UO_1387 (O_1387,N_22313,N_24566);
and UO_1388 (O_1388,N_24954,N_22223);
or UO_1389 (O_1389,N_23566,N_22943);
and UO_1390 (O_1390,N_22086,N_23920);
nand UO_1391 (O_1391,N_23133,N_23402);
nand UO_1392 (O_1392,N_23352,N_23953);
nor UO_1393 (O_1393,N_22515,N_24669);
or UO_1394 (O_1394,N_22897,N_24732);
or UO_1395 (O_1395,N_24330,N_24159);
and UO_1396 (O_1396,N_22162,N_23470);
nand UO_1397 (O_1397,N_23789,N_24984);
nand UO_1398 (O_1398,N_23190,N_23122);
nor UO_1399 (O_1399,N_24073,N_22669);
nand UO_1400 (O_1400,N_22286,N_23928);
nor UO_1401 (O_1401,N_23446,N_22798);
xor UO_1402 (O_1402,N_24883,N_24100);
or UO_1403 (O_1403,N_24001,N_22746);
and UO_1404 (O_1404,N_23772,N_24170);
nor UO_1405 (O_1405,N_22991,N_23663);
nor UO_1406 (O_1406,N_23418,N_21960);
and UO_1407 (O_1407,N_24664,N_22315);
or UO_1408 (O_1408,N_24415,N_22381);
nor UO_1409 (O_1409,N_23089,N_22085);
and UO_1410 (O_1410,N_22068,N_22156);
and UO_1411 (O_1411,N_22964,N_23593);
xnor UO_1412 (O_1412,N_24542,N_23202);
nor UO_1413 (O_1413,N_22096,N_24633);
and UO_1414 (O_1414,N_24403,N_23736);
or UO_1415 (O_1415,N_24014,N_23421);
or UO_1416 (O_1416,N_24243,N_23737);
nand UO_1417 (O_1417,N_24639,N_24555);
xor UO_1418 (O_1418,N_23088,N_23865);
nand UO_1419 (O_1419,N_23279,N_23233);
and UO_1420 (O_1420,N_22854,N_22505);
or UO_1421 (O_1421,N_23064,N_24987);
nor UO_1422 (O_1422,N_23734,N_22667);
or UO_1423 (O_1423,N_22900,N_22413);
or UO_1424 (O_1424,N_22006,N_23899);
nand UO_1425 (O_1425,N_23171,N_23411);
xor UO_1426 (O_1426,N_24481,N_24082);
nand UO_1427 (O_1427,N_23225,N_22109);
xor UO_1428 (O_1428,N_23793,N_23695);
and UO_1429 (O_1429,N_23834,N_24733);
and UO_1430 (O_1430,N_22768,N_22911);
nor UO_1431 (O_1431,N_21937,N_22914);
xor UO_1432 (O_1432,N_24661,N_24726);
xor UO_1433 (O_1433,N_22237,N_22214);
and UO_1434 (O_1434,N_23683,N_23144);
and UO_1435 (O_1435,N_22353,N_23661);
and UO_1436 (O_1436,N_22662,N_22032);
or UO_1437 (O_1437,N_23783,N_24049);
nand UO_1438 (O_1438,N_24054,N_24256);
and UO_1439 (O_1439,N_22437,N_24268);
xnor UO_1440 (O_1440,N_24453,N_24011);
and UO_1441 (O_1441,N_22176,N_24348);
nand UO_1442 (O_1442,N_23781,N_23288);
and UO_1443 (O_1443,N_22460,N_23546);
or UO_1444 (O_1444,N_24723,N_23107);
xnor UO_1445 (O_1445,N_23704,N_24541);
and UO_1446 (O_1446,N_22234,N_22482);
and UO_1447 (O_1447,N_24836,N_23901);
nor UO_1448 (O_1448,N_24788,N_24151);
and UO_1449 (O_1449,N_23452,N_23125);
nand UO_1450 (O_1450,N_24854,N_22387);
and UO_1451 (O_1451,N_24099,N_22161);
nand UO_1452 (O_1452,N_22147,N_22918);
xnor UO_1453 (O_1453,N_23852,N_23765);
nor UO_1454 (O_1454,N_24847,N_22440);
nor UO_1455 (O_1455,N_23343,N_21969);
and UO_1456 (O_1456,N_22442,N_22602);
nor UO_1457 (O_1457,N_22044,N_24979);
xor UO_1458 (O_1458,N_24764,N_22236);
nor UO_1459 (O_1459,N_24564,N_24806);
or UO_1460 (O_1460,N_24590,N_23688);
xnor UO_1461 (O_1461,N_24132,N_21957);
and UO_1462 (O_1462,N_23389,N_21984);
nand UO_1463 (O_1463,N_21877,N_23395);
nor UO_1464 (O_1464,N_24008,N_22967);
nor UO_1465 (O_1465,N_24673,N_24869);
nor UO_1466 (O_1466,N_24289,N_22526);
nand UO_1467 (O_1467,N_23441,N_22871);
nor UO_1468 (O_1468,N_22606,N_22005);
nor UO_1469 (O_1469,N_24687,N_24619);
nand UO_1470 (O_1470,N_22137,N_24372);
nand UO_1471 (O_1471,N_24551,N_23063);
and UO_1472 (O_1472,N_24630,N_22812);
nand UO_1473 (O_1473,N_22070,N_22690);
nand UO_1474 (O_1474,N_22693,N_22878);
and UO_1475 (O_1475,N_22188,N_24671);
nor UO_1476 (O_1476,N_24472,N_24463);
and UO_1477 (O_1477,N_24232,N_24505);
nand UO_1478 (O_1478,N_22262,N_23832);
and UO_1479 (O_1479,N_24597,N_24653);
and UO_1480 (O_1480,N_24784,N_23456);
nor UO_1481 (O_1481,N_22832,N_24533);
nand UO_1482 (O_1482,N_23835,N_22982);
or UO_1483 (O_1483,N_23222,N_22269);
or UO_1484 (O_1484,N_24601,N_24503);
nand UO_1485 (O_1485,N_23053,N_23888);
or UO_1486 (O_1486,N_23002,N_23251);
and UO_1487 (O_1487,N_23034,N_23327);
nand UO_1488 (O_1488,N_22751,N_22761);
nor UO_1489 (O_1489,N_23881,N_22664);
and UO_1490 (O_1490,N_22265,N_23631);
and UO_1491 (O_1491,N_22601,N_22609);
or UO_1492 (O_1492,N_23690,N_22950);
xnor UO_1493 (O_1493,N_23989,N_24473);
nand UO_1494 (O_1494,N_21902,N_24490);
nor UO_1495 (O_1495,N_22925,N_22164);
or UO_1496 (O_1496,N_24226,N_23647);
nor UO_1497 (O_1497,N_22094,N_22685);
and UO_1498 (O_1498,N_23443,N_23394);
or UO_1499 (O_1499,N_24589,N_22423);
nor UO_1500 (O_1500,N_22279,N_22962);
and UO_1501 (O_1501,N_21922,N_24070);
nor UO_1502 (O_1502,N_22772,N_23312);
and UO_1503 (O_1503,N_22978,N_23798);
nor UO_1504 (O_1504,N_22930,N_23758);
nor UO_1505 (O_1505,N_23199,N_23311);
nand UO_1506 (O_1506,N_23917,N_22055);
nand UO_1507 (O_1507,N_23521,N_24144);
xor UO_1508 (O_1508,N_23701,N_24596);
nand UO_1509 (O_1509,N_23525,N_24972);
nand UO_1510 (O_1510,N_23334,N_24058);
nor UO_1511 (O_1511,N_23294,N_24657);
nand UO_1512 (O_1512,N_23230,N_22309);
nor UO_1513 (O_1513,N_21924,N_22784);
and UO_1514 (O_1514,N_23277,N_24998);
nand UO_1515 (O_1515,N_24101,N_24652);
or UO_1516 (O_1516,N_23664,N_23416);
nand UO_1517 (O_1517,N_23070,N_24384);
or UO_1518 (O_1518,N_24562,N_21886);
nor UO_1519 (O_1519,N_22708,N_24770);
and UO_1520 (O_1520,N_23518,N_22862);
or UO_1521 (O_1521,N_24033,N_22850);
nand UO_1522 (O_1522,N_24091,N_22263);
or UO_1523 (O_1523,N_24825,N_22155);
nand UO_1524 (O_1524,N_24698,N_23130);
nor UO_1525 (O_1525,N_23797,N_24205);
or UO_1526 (O_1526,N_24548,N_24142);
nand UO_1527 (O_1527,N_23094,N_24141);
or UO_1528 (O_1528,N_24489,N_24685);
nor UO_1529 (O_1529,N_23554,N_22775);
or UO_1530 (O_1530,N_22870,N_24501);
or UO_1531 (O_1531,N_21970,N_24560);
and UO_1532 (O_1532,N_22630,N_23853);
nor UO_1533 (O_1533,N_23215,N_22513);
and UO_1534 (O_1534,N_24104,N_24387);
nand UO_1535 (O_1535,N_24980,N_22864);
or UO_1536 (O_1536,N_22014,N_24374);
nand UO_1537 (O_1537,N_21983,N_23196);
or UO_1538 (O_1538,N_24056,N_23360);
xnor UO_1539 (O_1539,N_22973,N_22311);
nand UO_1540 (O_1540,N_22403,N_24097);
nand UO_1541 (O_1541,N_22065,N_21930);
nand UO_1542 (O_1542,N_22568,N_23506);
nor UO_1543 (O_1543,N_22255,N_23851);
and UO_1544 (O_1544,N_22172,N_23364);
nor UO_1545 (O_1545,N_23477,N_23903);
and UO_1546 (O_1546,N_24870,N_22778);
nor UO_1547 (O_1547,N_22283,N_24135);
and UO_1548 (O_1548,N_22766,N_22519);
nor UO_1549 (O_1549,N_24604,N_22804);
nor UO_1550 (O_1550,N_24809,N_22674);
xor UO_1551 (O_1551,N_23491,N_23369);
nor UO_1552 (O_1552,N_24279,N_22929);
and UO_1553 (O_1553,N_23148,N_23382);
xor UO_1554 (O_1554,N_23780,N_23552);
or UO_1555 (O_1555,N_23234,N_22063);
nand UO_1556 (O_1556,N_22694,N_24858);
nand UO_1557 (O_1557,N_24837,N_23625);
nand UO_1558 (O_1558,N_23921,N_23559);
nand UO_1559 (O_1559,N_24561,N_22422);
or UO_1560 (O_1560,N_21900,N_22023);
or UO_1561 (O_1561,N_22193,N_23440);
and UO_1562 (O_1562,N_22168,N_24656);
and UO_1563 (O_1563,N_23322,N_24706);
nor UO_1564 (O_1564,N_22580,N_22719);
nor UO_1565 (O_1565,N_24603,N_22276);
nand UO_1566 (O_1566,N_22446,N_24971);
nand UO_1567 (O_1567,N_23776,N_22044);
nor UO_1568 (O_1568,N_22837,N_23578);
nand UO_1569 (O_1569,N_22792,N_23947);
and UO_1570 (O_1570,N_23278,N_23831);
or UO_1571 (O_1571,N_24728,N_24349);
nor UO_1572 (O_1572,N_22739,N_24399);
nand UO_1573 (O_1573,N_23457,N_22267);
xnor UO_1574 (O_1574,N_24586,N_24407);
or UO_1575 (O_1575,N_22426,N_23413);
nand UO_1576 (O_1576,N_24248,N_23253);
and UO_1577 (O_1577,N_24434,N_22696);
or UO_1578 (O_1578,N_23970,N_23759);
nand UO_1579 (O_1579,N_23572,N_23732);
nor UO_1580 (O_1580,N_22169,N_22966);
nor UO_1581 (O_1581,N_24099,N_24029);
xor UO_1582 (O_1582,N_22767,N_23700);
or UO_1583 (O_1583,N_22311,N_24276);
xor UO_1584 (O_1584,N_24419,N_22461);
nand UO_1585 (O_1585,N_23225,N_24510);
nand UO_1586 (O_1586,N_24876,N_22121);
nor UO_1587 (O_1587,N_22083,N_22454);
or UO_1588 (O_1588,N_24003,N_23767);
nand UO_1589 (O_1589,N_23215,N_23232);
and UO_1590 (O_1590,N_23140,N_22582);
nor UO_1591 (O_1591,N_23898,N_24199);
xor UO_1592 (O_1592,N_23644,N_22904);
or UO_1593 (O_1593,N_22865,N_24410);
and UO_1594 (O_1594,N_24706,N_23515);
or UO_1595 (O_1595,N_22633,N_24592);
or UO_1596 (O_1596,N_22380,N_23536);
nor UO_1597 (O_1597,N_24042,N_22922);
nand UO_1598 (O_1598,N_23297,N_24704);
nor UO_1599 (O_1599,N_23903,N_23892);
and UO_1600 (O_1600,N_23468,N_23909);
or UO_1601 (O_1601,N_22578,N_22527);
or UO_1602 (O_1602,N_23238,N_24878);
and UO_1603 (O_1603,N_21951,N_22826);
and UO_1604 (O_1604,N_22554,N_24137);
or UO_1605 (O_1605,N_24612,N_24543);
nor UO_1606 (O_1606,N_23153,N_22321);
or UO_1607 (O_1607,N_24548,N_24970);
or UO_1608 (O_1608,N_23677,N_24506);
and UO_1609 (O_1609,N_22773,N_24555);
nor UO_1610 (O_1610,N_24193,N_22781);
or UO_1611 (O_1611,N_24096,N_24765);
nand UO_1612 (O_1612,N_21969,N_24540);
and UO_1613 (O_1613,N_23332,N_23469);
nor UO_1614 (O_1614,N_23254,N_22242);
nand UO_1615 (O_1615,N_24388,N_22196);
or UO_1616 (O_1616,N_22158,N_24409);
or UO_1617 (O_1617,N_22993,N_23579);
nand UO_1618 (O_1618,N_22701,N_23315);
or UO_1619 (O_1619,N_22217,N_22676);
nor UO_1620 (O_1620,N_23733,N_22925);
xnor UO_1621 (O_1621,N_23613,N_21896);
and UO_1622 (O_1622,N_22852,N_24713);
or UO_1623 (O_1623,N_24165,N_24634);
or UO_1624 (O_1624,N_22050,N_23472);
and UO_1625 (O_1625,N_23560,N_22182);
nor UO_1626 (O_1626,N_24855,N_23341);
nand UO_1627 (O_1627,N_23722,N_22623);
or UO_1628 (O_1628,N_24303,N_24762);
nor UO_1629 (O_1629,N_23614,N_24912);
xor UO_1630 (O_1630,N_23343,N_24998);
and UO_1631 (O_1631,N_23523,N_22136);
or UO_1632 (O_1632,N_22430,N_22698);
nand UO_1633 (O_1633,N_24948,N_23981);
nor UO_1634 (O_1634,N_24704,N_24619);
nor UO_1635 (O_1635,N_23755,N_24141);
and UO_1636 (O_1636,N_22401,N_24901);
or UO_1637 (O_1637,N_22079,N_22537);
nor UO_1638 (O_1638,N_24002,N_24867);
nand UO_1639 (O_1639,N_22644,N_23631);
nand UO_1640 (O_1640,N_24704,N_24715);
or UO_1641 (O_1641,N_23603,N_24545);
or UO_1642 (O_1642,N_23750,N_24222);
nand UO_1643 (O_1643,N_24356,N_22401);
and UO_1644 (O_1644,N_22954,N_23348);
xnor UO_1645 (O_1645,N_23814,N_24472);
and UO_1646 (O_1646,N_24681,N_24459);
xor UO_1647 (O_1647,N_21991,N_24287);
nand UO_1648 (O_1648,N_24363,N_23815);
nor UO_1649 (O_1649,N_24360,N_22559);
nand UO_1650 (O_1650,N_24514,N_24579);
nor UO_1651 (O_1651,N_23005,N_23822);
nor UO_1652 (O_1652,N_23097,N_24396);
and UO_1653 (O_1653,N_22328,N_24419);
nor UO_1654 (O_1654,N_24597,N_24056);
nand UO_1655 (O_1655,N_24596,N_22885);
or UO_1656 (O_1656,N_24780,N_23747);
nand UO_1657 (O_1657,N_23749,N_22063);
nor UO_1658 (O_1658,N_22971,N_23384);
nor UO_1659 (O_1659,N_22899,N_23901);
xor UO_1660 (O_1660,N_22126,N_22353);
nor UO_1661 (O_1661,N_23709,N_23295);
xnor UO_1662 (O_1662,N_24167,N_24624);
nand UO_1663 (O_1663,N_23932,N_22408);
or UO_1664 (O_1664,N_23421,N_24748);
nand UO_1665 (O_1665,N_23397,N_22727);
and UO_1666 (O_1666,N_22768,N_23260);
nand UO_1667 (O_1667,N_21935,N_24659);
and UO_1668 (O_1668,N_21941,N_24395);
nand UO_1669 (O_1669,N_24628,N_24981);
or UO_1670 (O_1670,N_23110,N_23713);
nor UO_1671 (O_1671,N_24319,N_22459);
nand UO_1672 (O_1672,N_24538,N_24338);
nor UO_1673 (O_1673,N_22038,N_23823);
or UO_1674 (O_1674,N_22548,N_23178);
or UO_1675 (O_1675,N_23717,N_22741);
nand UO_1676 (O_1676,N_23249,N_22176);
nor UO_1677 (O_1677,N_22577,N_24906);
or UO_1678 (O_1678,N_24444,N_24266);
nand UO_1679 (O_1679,N_23250,N_21946);
nor UO_1680 (O_1680,N_24883,N_22229);
or UO_1681 (O_1681,N_22515,N_24680);
nand UO_1682 (O_1682,N_24894,N_24501);
or UO_1683 (O_1683,N_23943,N_22393);
or UO_1684 (O_1684,N_22233,N_22142);
nor UO_1685 (O_1685,N_23115,N_24378);
nor UO_1686 (O_1686,N_24735,N_24016);
nand UO_1687 (O_1687,N_22831,N_22173);
nor UO_1688 (O_1688,N_24592,N_24970);
nor UO_1689 (O_1689,N_21946,N_22817);
and UO_1690 (O_1690,N_22223,N_22093);
nand UO_1691 (O_1691,N_22093,N_22655);
or UO_1692 (O_1692,N_23544,N_22769);
and UO_1693 (O_1693,N_23138,N_23156);
nand UO_1694 (O_1694,N_23202,N_22401);
or UO_1695 (O_1695,N_24942,N_23393);
nand UO_1696 (O_1696,N_23905,N_24251);
or UO_1697 (O_1697,N_22371,N_22451);
nor UO_1698 (O_1698,N_22867,N_24924);
and UO_1699 (O_1699,N_24787,N_24858);
nand UO_1700 (O_1700,N_23982,N_22684);
or UO_1701 (O_1701,N_23905,N_24936);
and UO_1702 (O_1702,N_24346,N_24481);
and UO_1703 (O_1703,N_22495,N_21946);
or UO_1704 (O_1704,N_24128,N_24683);
nand UO_1705 (O_1705,N_24283,N_24239);
and UO_1706 (O_1706,N_22276,N_22854);
and UO_1707 (O_1707,N_23975,N_22148);
nor UO_1708 (O_1708,N_22159,N_24803);
nor UO_1709 (O_1709,N_22645,N_22876);
or UO_1710 (O_1710,N_22791,N_24960);
or UO_1711 (O_1711,N_22304,N_24293);
or UO_1712 (O_1712,N_24586,N_24339);
nand UO_1713 (O_1713,N_22183,N_22420);
nand UO_1714 (O_1714,N_23278,N_23999);
nor UO_1715 (O_1715,N_24332,N_24616);
and UO_1716 (O_1716,N_24436,N_24973);
nor UO_1717 (O_1717,N_24472,N_24247);
xnor UO_1718 (O_1718,N_23913,N_24195);
nand UO_1719 (O_1719,N_22427,N_23841);
nor UO_1720 (O_1720,N_24427,N_22811);
and UO_1721 (O_1721,N_23814,N_23891);
or UO_1722 (O_1722,N_22308,N_24527);
or UO_1723 (O_1723,N_23230,N_24115);
or UO_1724 (O_1724,N_24647,N_24094);
nor UO_1725 (O_1725,N_24371,N_23612);
nor UO_1726 (O_1726,N_22084,N_23131);
or UO_1727 (O_1727,N_24179,N_22597);
or UO_1728 (O_1728,N_24697,N_22384);
nand UO_1729 (O_1729,N_24658,N_24623);
and UO_1730 (O_1730,N_21980,N_23396);
and UO_1731 (O_1731,N_22889,N_21978);
xnor UO_1732 (O_1732,N_23458,N_24352);
xor UO_1733 (O_1733,N_23363,N_24214);
nor UO_1734 (O_1734,N_23125,N_24592);
nor UO_1735 (O_1735,N_24263,N_24479);
xor UO_1736 (O_1736,N_22980,N_24549);
and UO_1737 (O_1737,N_23444,N_22479);
xor UO_1738 (O_1738,N_23519,N_23556);
nor UO_1739 (O_1739,N_23670,N_24811);
nand UO_1740 (O_1740,N_23873,N_22689);
and UO_1741 (O_1741,N_23511,N_23944);
and UO_1742 (O_1742,N_21925,N_24798);
or UO_1743 (O_1743,N_22834,N_23817);
nand UO_1744 (O_1744,N_24398,N_24595);
nor UO_1745 (O_1745,N_22411,N_24145);
nor UO_1746 (O_1746,N_23342,N_24078);
xor UO_1747 (O_1747,N_23708,N_24496);
nor UO_1748 (O_1748,N_22592,N_24498);
nand UO_1749 (O_1749,N_22775,N_23911);
or UO_1750 (O_1750,N_23138,N_23487);
xor UO_1751 (O_1751,N_23989,N_23787);
nor UO_1752 (O_1752,N_24037,N_24181);
and UO_1753 (O_1753,N_22831,N_23016);
nand UO_1754 (O_1754,N_22545,N_23327);
nor UO_1755 (O_1755,N_24474,N_24599);
nor UO_1756 (O_1756,N_22697,N_23182);
or UO_1757 (O_1757,N_23286,N_22676);
nand UO_1758 (O_1758,N_24477,N_24424);
nor UO_1759 (O_1759,N_22341,N_24827);
nor UO_1760 (O_1760,N_24301,N_24473);
or UO_1761 (O_1761,N_22468,N_24145);
nor UO_1762 (O_1762,N_24924,N_22017);
nor UO_1763 (O_1763,N_22475,N_23661);
and UO_1764 (O_1764,N_24880,N_24359);
nor UO_1765 (O_1765,N_22646,N_23386);
nand UO_1766 (O_1766,N_21954,N_22942);
or UO_1767 (O_1767,N_22793,N_24338);
and UO_1768 (O_1768,N_23467,N_24468);
and UO_1769 (O_1769,N_22078,N_24249);
nor UO_1770 (O_1770,N_23875,N_23390);
or UO_1771 (O_1771,N_22097,N_24863);
or UO_1772 (O_1772,N_24996,N_23153);
and UO_1773 (O_1773,N_22627,N_23082);
or UO_1774 (O_1774,N_24879,N_22866);
nand UO_1775 (O_1775,N_24510,N_22579);
nor UO_1776 (O_1776,N_23458,N_24710);
or UO_1777 (O_1777,N_24346,N_22035);
nand UO_1778 (O_1778,N_23691,N_23501);
or UO_1779 (O_1779,N_22100,N_23545);
or UO_1780 (O_1780,N_24260,N_24628);
nor UO_1781 (O_1781,N_23027,N_22708);
or UO_1782 (O_1782,N_24151,N_24146);
xor UO_1783 (O_1783,N_24477,N_22823);
and UO_1784 (O_1784,N_24346,N_24448);
nor UO_1785 (O_1785,N_24089,N_24719);
and UO_1786 (O_1786,N_22220,N_24728);
nand UO_1787 (O_1787,N_24864,N_23963);
nand UO_1788 (O_1788,N_23876,N_22531);
xor UO_1789 (O_1789,N_23459,N_24880);
xor UO_1790 (O_1790,N_22319,N_24878);
and UO_1791 (O_1791,N_22291,N_24684);
nor UO_1792 (O_1792,N_23414,N_24340);
or UO_1793 (O_1793,N_22746,N_23803);
nor UO_1794 (O_1794,N_24345,N_24932);
or UO_1795 (O_1795,N_21964,N_24674);
xor UO_1796 (O_1796,N_23034,N_23144);
or UO_1797 (O_1797,N_24703,N_22946);
or UO_1798 (O_1798,N_23476,N_24784);
nand UO_1799 (O_1799,N_22221,N_23838);
or UO_1800 (O_1800,N_23971,N_23425);
nor UO_1801 (O_1801,N_21954,N_24914);
or UO_1802 (O_1802,N_23110,N_23104);
nor UO_1803 (O_1803,N_23810,N_24097);
nor UO_1804 (O_1804,N_24525,N_24751);
or UO_1805 (O_1805,N_24766,N_23373);
and UO_1806 (O_1806,N_24724,N_23805);
or UO_1807 (O_1807,N_23643,N_23332);
or UO_1808 (O_1808,N_24639,N_24542);
nand UO_1809 (O_1809,N_22064,N_23658);
nor UO_1810 (O_1810,N_22409,N_22959);
or UO_1811 (O_1811,N_22931,N_23123);
and UO_1812 (O_1812,N_22845,N_22505);
nor UO_1813 (O_1813,N_24201,N_22348);
nand UO_1814 (O_1814,N_23322,N_24658);
nor UO_1815 (O_1815,N_23616,N_23146);
nor UO_1816 (O_1816,N_24142,N_22832);
and UO_1817 (O_1817,N_22325,N_24234);
nor UO_1818 (O_1818,N_22928,N_23379);
nor UO_1819 (O_1819,N_23259,N_23356);
and UO_1820 (O_1820,N_23080,N_22691);
or UO_1821 (O_1821,N_22702,N_24270);
nand UO_1822 (O_1822,N_23014,N_23828);
xor UO_1823 (O_1823,N_23373,N_23655);
nand UO_1824 (O_1824,N_22545,N_24776);
nor UO_1825 (O_1825,N_23565,N_22621);
nor UO_1826 (O_1826,N_23414,N_24788);
or UO_1827 (O_1827,N_23701,N_22342);
nand UO_1828 (O_1828,N_23444,N_23578);
and UO_1829 (O_1829,N_24381,N_24941);
nand UO_1830 (O_1830,N_23911,N_23320);
and UO_1831 (O_1831,N_23379,N_22554);
or UO_1832 (O_1832,N_22889,N_22626);
xor UO_1833 (O_1833,N_23935,N_24722);
nand UO_1834 (O_1834,N_22160,N_22284);
nand UO_1835 (O_1835,N_22994,N_21941);
and UO_1836 (O_1836,N_22618,N_22042);
and UO_1837 (O_1837,N_23801,N_24603);
or UO_1838 (O_1838,N_24204,N_23723);
nor UO_1839 (O_1839,N_22470,N_22390);
nor UO_1840 (O_1840,N_23772,N_22665);
nor UO_1841 (O_1841,N_21968,N_24604);
and UO_1842 (O_1842,N_22510,N_23761);
nand UO_1843 (O_1843,N_24984,N_23220);
nor UO_1844 (O_1844,N_23318,N_22670);
and UO_1845 (O_1845,N_23509,N_23882);
xnor UO_1846 (O_1846,N_22068,N_24700);
and UO_1847 (O_1847,N_22427,N_24601);
and UO_1848 (O_1848,N_21896,N_23209);
or UO_1849 (O_1849,N_24651,N_23341);
or UO_1850 (O_1850,N_24281,N_24140);
xnor UO_1851 (O_1851,N_22151,N_24585);
nor UO_1852 (O_1852,N_23328,N_23582);
nand UO_1853 (O_1853,N_24927,N_22545);
xnor UO_1854 (O_1854,N_24404,N_23792);
xnor UO_1855 (O_1855,N_22675,N_24569);
nor UO_1856 (O_1856,N_22912,N_24143);
or UO_1857 (O_1857,N_22770,N_22385);
nor UO_1858 (O_1858,N_23154,N_24649);
nor UO_1859 (O_1859,N_24207,N_22994);
or UO_1860 (O_1860,N_24454,N_22604);
xnor UO_1861 (O_1861,N_23336,N_22288);
and UO_1862 (O_1862,N_22182,N_23843);
nand UO_1863 (O_1863,N_23525,N_24869);
or UO_1864 (O_1864,N_24511,N_22690);
nand UO_1865 (O_1865,N_23236,N_23909);
nand UO_1866 (O_1866,N_23285,N_23931);
nor UO_1867 (O_1867,N_24828,N_24914);
and UO_1868 (O_1868,N_24465,N_23689);
nand UO_1869 (O_1869,N_23311,N_23872);
and UO_1870 (O_1870,N_24740,N_22488);
nor UO_1871 (O_1871,N_23633,N_22584);
nor UO_1872 (O_1872,N_22001,N_23445);
xnor UO_1873 (O_1873,N_23016,N_23592);
xor UO_1874 (O_1874,N_24589,N_24876);
and UO_1875 (O_1875,N_22940,N_22623);
nor UO_1876 (O_1876,N_24985,N_24394);
nand UO_1877 (O_1877,N_23001,N_23148);
or UO_1878 (O_1878,N_22627,N_22079);
and UO_1879 (O_1879,N_23113,N_21923);
and UO_1880 (O_1880,N_22414,N_24277);
xnor UO_1881 (O_1881,N_22195,N_24871);
xor UO_1882 (O_1882,N_22154,N_24688);
nand UO_1883 (O_1883,N_23751,N_23210);
or UO_1884 (O_1884,N_24468,N_24061);
nor UO_1885 (O_1885,N_24507,N_23851);
and UO_1886 (O_1886,N_22692,N_23208);
xnor UO_1887 (O_1887,N_22250,N_22663);
nand UO_1888 (O_1888,N_23169,N_23562);
and UO_1889 (O_1889,N_24601,N_22565);
and UO_1890 (O_1890,N_23507,N_23194);
and UO_1891 (O_1891,N_22017,N_24008);
nand UO_1892 (O_1892,N_21987,N_23632);
and UO_1893 (O_1893,N_23376,N_23653);
xnor UO_1894 (O_1894,N_22912,N_23360);
and UO_1895 (O_1895,N_24642,N_24686);
and UO_1896 (O_1896,N_22185,N_24511);
nor UO_1897 (O_1897,N_23008,N_21995);
nor UO_1898 (O_1898,N_23003,N_23098);
or UO_1899 (O_1899,N_23234,N_22833);
nor UO_1900 (O_1900,N_23675,N_23193);
or UO_1901 (O_1901,N_22562,N_22679);
nor UO_1902 (O_1902,N_23837,N_23298);
and UO_1903 (O_1903,N_23740,N_22871);
nor UO_1904 (O_1904,N_22819,N_24066);
nand UO_1905 (O_1905,N_23798,N_23771);
and UO_1906 (O_1906,N_23274,N_22920);
nand UO_1907 (O_1907,N_24288,N_22482);
and UO_1908 (O_1908,N_22657,N_22138);
nor UO_1909 (O_1909,N_22967,N_23690);
or UO_1910 (O_1910,N_23456,N_23013);
or UO_1911 (O_1911,N_24979,N_22707);
or UO_1912 (O_1912,N_23776,N_22545);
nand UO_1913 (O_1913,N_22962,N_22742);
and UO_1914 (O_1914,N_23981,N_22048);
and UO_1915 (O_1915,N_21966,N_24735);
and UO_1916 (O_1916,N_24698,N_22544);
nor UO_1917 (O_1917,N_23766,N_24477);
or UO_1918 (O_1918,N_23863,N_24115);
nand UO_1919 (O_1919,N_22781,N_22387);
and UO_1920 (O_1920,N_24451,N_21941);
nand UO_1921 (O_1921,N_24177,N_22599);
or UO_1922 (O_1922,N_22943,N_24323);
or UO_1923 (O_1923,N_23341,N_22635);
or UO_1924 (O_1924,N_23951,N_23106);
nand UO_1925 (O_1925,N_24678,N_22339);
xnor UO_1926 (O_1926,N_22771,N_23114);
and UO_1927 (O_1927,N_24638,N_23581);
or UO_1928 (O_1928,N_22874,N_22306);
nand UO_1929 (O_1929,N_24576,N_24749);
and UO_1930 (O_1930,N_24033,N_23079);
and UO_1931 (O_1931,N_23293,N_24446);
nor UO_1932 (O_1932,N_21984,N_21986);
and UO_1933 (O_1933,N_22670,N_23256);
nor UO_1934 (O_1934,N_24539,N_22212);
and UO_1935 (O_1935,N_24179,N_23774);
or UO_1936 (O_1936,N_22373,N_23160);
xor UO_1937 (O_1937,N_22195,N_24268);
nor UO_1938 (O_1938,N_24320,N_23724);
and UO_1939 (O_1939,N_23065,N_23461);
nor UO_1940 (O_1940,N_24204,N_23706);
xnor UO_1941 (O_1941,N_23308,N_22564);
nand UO_1942 (O_1942,N_24178,N_23256);
or UO_1943 (O_1943,N_24914,N_24664);
nand UO_1944 (O_1944,N_24753,N_24535);
xor UO_1945 (O_1945,N_23480,N_24606);
xnor UO_1946 (O_1946,N_21921,N_22671);
nand UO_1947 (O_1947,N_24308,N_24119);
and UO_1948 (O_1948,N_23631,N_22741);
and UO_1949 (O_1949,N_24935,N_24380);
nand UO_1950 (O_1950,N_22229,N_23392);
nand UO_1951 (O_1951,N_22166,N_23425);
nor UO_1952 (O_1952,N_23284,N_22873);
nor UO_1953 (O_1953,N_24349,N_24897);
and UO_1954 (O_1954,N_24556,N_23360);
and UO_1955 (O_1955,N_22775,N_24598);
nand UO_1956 (O_1956,N_24938,N_22845);
xnor UO_1957 (O_1957,N_22430,N_23278);
nand UO_1958 (O_1958,N_24736,N_24922);
or UO_1959 (O_1959,N_24527,N_24043);
or UO_1960 (O_1960,N_23561,N_22267);
nor UO_1961 (O_1961,N_22649,N_22174);
xnor UO_1962 (O_1962,N_23691,N_24438);
and UO_1963 (O_1963,N_23280,N_23076);
nor UO_1964 (O_1964,N_24266,N_22184);
nand UO_1965 (O_1965,N_24612,N_23280);
or UO_1966 (O_1966,N_23900,N_23786);
nand UO_1967 (O_1967,N_23657,N_23160);
or UO_1968 (O_1968,N_24632,N_24346);
or UO_1969 (O_1969,N_24518,N_24003);
nor UO_1970 (O_1970,N_22140,N_23779);
or UO_1971 (O_1971,N_22380,N_22984);
or UO_1972 (O_1972,N_24559,N_24339);
or UO_1973 (O_1973,N_22807,N_22116);
or UO_1974 (O_1974,N_22853,N_23970);
nor UO_1975 (O_1975,N_22615,N_23077);
or UO_1976 (O_1976,N_23865,N_22835);
nor UO_1977 (O_1977,N_24899,N_24214);
nor UO_1978 (O_1978,N_24921,N_23950);
nor UO_1979 (O_1979,N_24560,N_23989);
xor UO_1980 (O_1980,N_24565,N_24408);
nand UO_1981 (O_1981,N_23066,N_23090);
nor UO_1982 (O_1982,N_23886,N_24941);
nor UO_1983 (O_1983,N_24859,N_24149);
or UO_1984 (O_1984,N_23502,N_23140);
nand UO_1985 (O_1985,N_22232,N_23582);
nand UO_1986 (O_1986,N_22909,N_23233);
and UO_1987 (O_1987,N_22275,N_22167);
nand UO_1988 (O_1988,N_23797,N_21960);
or UO_1989 (O_1989,N_24026,N_22439);
or UO_1990 (O_1990,N_23433,N_23319);
or UO_1991 (O_1991,N_22994,N_23702);
nor UO_1992 (O_1992,N_24007,N_23531);
nor UO_1993 (O_1993,N_21918,N_23704);
and UO_1994 (O_1994,N_24376,N_24538);
or UO_1995 (O_1995,N_24244,N_22495);
nor UO_1996 (O_1996,N_22675,N_22144);
and UO_1997 (O_1997,N_23639,N_22307);
nor UO_1998 (O_1998,N_24561,N_24669);
nor UO_1999 (O_1999,N_24802,N_24509);
nand UO_2000 (O_2000,N_22798,N_22885);
or UO_2001 (O_2001,N_23206,N_24556);
xor UO_2002 (O_2002,N_24737,N_24137);
nor UO_2003 (O_2003,N_23426,N_22554);
and UO_2004 (O_2004,N_22259,N_22943);
nand UO_2005 (O_2005,N_24206,N_24997);
nand UO_2006 (O_2006,N_22091,N_24021);
or UO_2007 (O_2007,N_22057,N_22183);
nand UO_2008 (O_2008,N_24576,N_23817);
xnor UO_2009 (O_2009,N_22395,N_23875);
and UO_2010 (O_2010,N_24297,N_24001);
and UO_2011 (O_2011,N_23562,N_22970);
or UO_2012 (O_2012,N_22055,N_22871);
nor UO_2013 (O_2013,N_23741,N_22220);
nand UO_2014 (O_2014,N_23327,N_23750);
or UO_2015 (O_2015,N_24763,N_24764);
nand UO_2016 (O_2016,N_23479,N_22351);
nand UO_2017 (O_2017,N_22500,N_24230);
xnor UO_2018 (O_2018,N_22915,N_24032);
nand UO_2019 (O_2019,N_23762,N_22767);
xor UO_2020 (O_2020,N_23854,N_22279);
and UO_2021 (O_2021,N_23461,N_22475);
xnor UO_2022 (O_2022,N_22135,N_24890);
nand UO_2023 (O_2023,N_23149,N_24659);
nor UO_2024 (O_2024,N_24929,N_23294);
nor UO_2025 (O_2025,N_23807,N_24326);
xor UO_2026 (O_2026,N_23172,N_24292);
nor UO_2027 (O_2027,N_24838,N_24178);
and UO_2028 (O_2028,N_23044,N_21890);
nor UO_2029 (O_2029,N_22496,N_22833);
or UO_2030 (O_2030,N_22821,N_23255);
or UO_2031 (O_2031,N_23531,N_23439);
nor UO_2032 (O_2032,N_22947,N_22896);
xor UO_2033 (O_2033,N_23218,N_24186);
and UO_2034 (O_2034,N_22674,N_22738);
and UO_2035 (O_2035,N_24279,N_24421);
and UO_2036 (O_2036,N_22727,N_21984);
nor UO_2037 (O_2037,N_24824,N_22145);
or UO_2038 (O_2038,N_24999,N_21981);
or UO_2039 (O_2039,N_23934,N_24017);
nand UO_2040 (O_2040,N_23868,N_22747);
nand UO_2041 (O_2041,N_24061,N_24409);
or UO_2042 (O_2042,N_22991,N_22877);
and UO_2043 (O_2043,N_23969,N_22510);
nor UO_2044 (O_2044,N_22650,N_23208);
nor UO_2045 (O_2045,N_23873,N_23904);
nor UO_2046 (O_2046,N_22054,N_24713);
nor UO_2047 (O_2047,N_22442,N_24114);
or UO_2048 (O_2048,N_23543,N_23992);
nor UO_2049 (O_2049,N_23924,N_22330);
nand UO_2050 (O_2050,N_24154,N_24441);
nand UO_2051 (O_2051,N_24112,N_22071);
or UO_2052 (O_2052,N_24788,N_23455);
or UO_2053 (O_2053,N_24402,N_24203);
and UO_2054 (O_2054,N_23507,N_22138);
nor UO_2055 (O_2055,N_23258,N_22887);
and UO_2056 (O_2056,N_23834,N_22976);
nor UO_2057 (O_2057,N_24811,N_23386);
nand UO_2058 (O_2058,N_24042,N_24662);
nand UO_2059 (O_2059,N_23347,N_23800);
or UO_2060 (O_2060,N_24240,N_22929);
or UO_2061 (O_2061,N_22024,N_24970);
and UO_2062 (O_2062,N_24396,N_23291);
nor UO_2063 (O_2063,N_24294,N_23668);
nor UO_2064 (O_2064,N_21927,N_23496);
nor UO_2065 (O_2065,N_24351,N_23148);
and UO_2066 (O_2066,N_22045,N_22839);
and UO_2067 (O_2067,N_24260,N_23750);
nor UO_2068 (O_2068,N_24421,N_23159);
nand UO_2069 (O_2069,N_22488,N_22665);
or UO_2070 (O_2070,N_24187,N_22655);
or UO_2071 (O_2071,N_23846,N_24464);
nand UO_2072 (O_2072,N_23374,N_23825);
or UO_2073 (O_2073,N_22341,N_22614);
nand UO_2074 (O_2074,N_23475,N_23460);
and UO_2075 (O_2075,N_23266,N_23041);
nor UO_2076 (O_2076,N_24150,N_23905);
nor UO_2077 (O_2077,N_24602,N_24458);
and UO_2078 (O_2078,N_22781,N_23720);
nor UO_2079 (O_2079,N_24041,N_24871);
or UO_2080 (O_2080,N_23437,N_24808);
nand UO_2081 (O_2081,N_23107,N_24889);
or UO_2082 (O_2082,N_22702,N_23730);
xor UO_2083 (O_2083,N_23724,N_22146);
and UO_2084 (O_2084,N_23293,N_24312);
nand UO_2085 (O_2085,N_23929,N_24012);
and UO_2086 (O_2086,N_22396,N_23895);
xnor UO_2087 (O_2087,N_23666,N_24836);
and UO_2088 (O_2088,N_24584,N_23620);
and UO_2089 (O_2089,N_24905,N_23225);
and UO_2090 (O_2090,N_24712,N_22786);
nor UO_2091 (O_2091,N_24434,N_23339);
nand UO_2092 (O_2092,N_22582,N_23038);
nor UO_2093 (O_2093,N_23091,N_23559);
nor UO_2094 (O_2094,N_23072,N_22494);
or UO_2095 (O_2095,N_23688,N_24650);
xnor UO_2096 (O_2096,N_22047,N_23059);
and UO_2097 (O_2097,N_22503,N_23281);
or UO_2098 (O_2098,N_22295,N_22236);
nand UO_2099 (O_2099,N_23954,N_22934);
and UO_2100 (O_2100,N_23831,N_24100);
and UO_2101 (O_2101,N_23698,N_24611);
nor UO_2102 (O_2102,N_23691,N_23972);
xor UO_2103 (O_2103,N_23264,N_24352);
nand UO_2104 (O_2104,N_23965,N_22444);
or UO_2105 (O_2105,N_22635,N_24566);
nand UO_2106 (O_2106,N_24882,N_22939);
nor UO_2107 (O_2107,N_24286,N_21965);
or UO_2108 (O_2108,N_24254,N_21923);
xnor UO_2109 (O_2109,N_22829,N_22714);
xor UO_2110 (O_2110,N_24016,N_24325);
xor UO_2111 (O_2111,N_23816,N_23653);
nor UO_2112 (O_2112,N_23484,N_23189);
xor UO_2113 (O_2113,N_23880,N_21878);
nand UO_2114 (O_2114,N_24059,N_23382);
and UO_2115 (O_2115,N_23141,N_24161);
or UO_2116 (O_2116,N_24395,N_23858);
nand UO_2117 (O_2117,N_23091,N_22113);
and UO_2118 (O_2118,N_23666,N_24145);
and UO_2119 (O_2119,N_24650,N_22357);
nand UO_2120 (O_2120,N_22845,N_23995);
nor UO_2121 (O_2121,N_23654,N_24843);
nor UO_2122 (O_2122,N_24572,N_24001);
nand UO_2123 (O_2123,N_24326,N_21989);
or UO_2124 (O_2124,N_22345,N_22712);
or UO_2125 (O_2125,N_23106,N_24112);
or UO_2126 (O_2126,N_24395,N_22385);
or UO_2127 (O_2127,N_23650,N_22778);
or UO_2128 (O_2128,N_23038,N_24453);
nor UO_2129 (O_2129,N_22581,N_22305);
or UO_2130 (O_2130,N_23193,N_23908);
nand UO_2131 (O_2131,N_22507,N_24350);
or UO_2132 (O_2132,N_24325,N_22740);
or UO_2133 (O_2133,N_23550,N_23459);
nor UO_2134 (O_2134,N_22814,N_24918);
nor UO_2135 (O_2135,N_24388,N_24222);
and UO_2136 (O_2136,N_22721,N_22827);
or UO_2137 (O_2137,N_22867,N_22673);
nand UO_2138 (O_2138,N_22580,N_22584);
xor UO_2139 (O_2139,N_22497,N_24549);
xnor UO_2140 (O_2140,N_23642,N_22188);
nor UO_2141 (O_2141,N_22827,N_23946);
nand UO_2142 (O_2142,N_24039,N_21891);
nor UO_2143 (O_2143,N_24335,N_24459);
and UO_2144 (O_2144,N_23170,N_22965);
nand UO_2145 (O_2145,N_22135,N_23561);
or UO_2146 (O_2146,N_24154,N_24552);
nand UO_2147 (O_2147,N_22452,N_23524);
or UO_2148 (O_2148,N_22043,N_23902);
or UO_2149 (O_2149,N_22628,N_23685);
nor UO_2150 (O_2150,N_22825,N_22729);
nand UO_2151 (O_2151,N_24560,N_24675);
nand UO_2152 (O_2152,N_21898,N_22089);
nor UO_2153 (O_2153,N_23709,N_24949);
nor UO_2154 (O_2154,N_24096,N_22501);
nand UO_2155 (O_2155,N_24523,N_23376);
nor UO_2156 (O_2156,N_23810,N_22912);
or UO_2157 (O_2157,N_22917,N_24569);
and UO_2158 (O_2158,N_22796,N_24947);
nand UO_2159 (O_2159,N_23619,N_24289);
nor UO_2160 (O_2160,N_22615,N_24679);
nor UO_2161 (O_2161,N_24887,N_21903);
and UO_2162 (O_2162,N_21988,N_23198);
nand UO_2163 (O_2163,N_23836,N_22353);
nand UO_2164 (O_2164,N_23587,N_23153);
or UO_2165 (O_2165,N_23882,N_22943);
nor UO_2166 (O_2166,N_23804,N_21878);
xor UO_2167 (O_2167,N_22928,N_24262);
and UO_2168 (O_2168,N_24752,N_24015);
xnor UO_2169 (O_2169,N_24929,N_22743);
nor UO_2170 (O_2170,N_23250,N_23960);
xnor UO_2171 (O_2171,N_22996,N_24032);
and UO_2172 (O_2172,N_21904,N_23132);
and UO_2173 (O_2173,N_22657,N_23716);
nor UO_2174 (O_2174,N_23278,N_23455);
and UO_2175 (O_2175,N_23152,N_24094);
and UO_2176 (O_2176,N_23425,N_24645);
nor UO_2177 (O_2177,N_24862,N_23142);
or UO_2178 (O_2178,N_22613,N_23683);
and UO_2179 (O_2179,N_22007,N_24769);
or UO_2180 (O_2180,N_23509,N_24233);
nor UO_2181 (O_2181,N_23572,N_23287);
nor UO_2182 (O_2182,N_24342,N_23335);
or UO_2183 (O_2183,N_24475,N_22670);
xnor UO_2184 (O_2184,N_24270,N_23827);
nand UO_2185 (O_2185,N_23832,N_24954);
nor UO_2186 (O_2186,N_23887,N_22594);
nor UO_2187 (O_2187,N_23971,N_23289);
or UO_2188 (O_2188,N_23028,N_22365);
nor UO_2189 (O_2189,N_22104,N_23896);
nand UO_2190 (O_2190,N_24368,N_22252);
nor UO_2191 (O_2191,N_22372,N_23252);
and UO_2192 (O_2192,N_22171,N_22435);
or UO_2193 (O_2193,N_23775,N_23958);
nor UO_2194 (O_2194,N_23896,N_22092);
or UO_2195 (O_2195,N_22400,N_22124);
or UO_2196 (O_2196,N_24015,N_22967);
or UO_2197 (O_2197,N_22177,N_24616);
nor UO_2198 (O_2198,N_21951,N_24357);
or UO_2199 (O_2199,N_24649,N_24332);
nand UO_2200 (O_2200,N_24019,N_21982);
xnor UO_2201 (O_2201,N_24258,N_22182);
or UO_2202 (O_2202,N_22975,N_23255);
and UO_2203 (O_2203,N_23494,N_24067);
nor UO_2204 (O_2204,N_24264,N_22657);
or UO_2205 (O_2205,N_21958,N_24173);
and UO_2206 (O_2206,N_24034,N_24734);
and UO_2207 (O_2207,N_23485,N_23458);
nor UO_2208 (O_2208,N_24656,N_22385);
nand UO_2209 (O_2209,N_23309,N_22441);
nor UO_2210 (O_2210,N_22596,N_23350);
nand UO_2211 (O_2211,N_23975,N_23550);
or UO_2212 (O_2212,N_22493,N_23046);
nand UO_2213 (O_2213,N_23582,N_22160);
or UO_2214 (O_2214,N_24736,N_24299);
xor UO_2215 (O_2215,N_21903,N_21977);
xnor UO_2216 (O_2216,N_24943,N_22343);
nand UO_2217 (O_2217,N_23018,N_23148);
and UO_2218 (O_2218,N_24145,N_24176);
or UO_2219 (O_2219,N_24436,N_24926);
and UO_2220 (O_2220,N_24932,N_22747);
and UO_2221 (O_2221,N_23450,N_23556);
and UO_2222 (O_2222,N_24002,N_22761);
and UO_2223 (O_2223,N_24344,N_23789);
nor UO_2224 (O_2224,N_22658,N_23304);
and UO_2225 (O_2225,N_23230,N_22362);
and UO_2226 (O_2226,N_23983,N_22686);
and UO_2227 (O_2227,N_22152,N_22891);
nand UO_2228 (O_2228,N_23671,N_24835);
nand UO_2229 (O_2229,N_22357,N_24691);
xor UO_2230 (O_2230,N_24758,N_23703);
nor UO_2231 (O_2231,N_21965,N_23963);
nor UO_2232 (O_2232,N_24012,N_22674);
xnor UO_2233 (O_2233,N_24239,N_22676);
nand UO_2234 (O_2234,N_23357,N_24378);
or UO_2235 (O_2235,N_22508,N_22126);
nor UO_2236 (O_2236,N_21915,N_24321);
or UO_2237 (O_2237,N_21967,N_24702);
or UO_2238 (O_2238,N_23442,N_24870);
and UO_2239 (O_2239,N_23417,N_21931);
and UO_2240 (O_2240,N_23950,N_24275);
and UO_2241 (O_2241,N_24381,N_23604);
nor UO_2242 (O_2242,N_22617,N_22789);
and UO_2243 (O_2243,N_24007,N_23543);
and UO_2244 (O_2244,N_22426,N_24650);
nor UO_2245 (O_2245,N_22141,N_22196);
nor UO_2246 (O_2246,N_24027,N_24104);
nand UO_2247 (O_2247,N_22701,N_24935);
nand UO_2248 (O_2248,N_22582,N_22478);
nor UO_2249 (O_2249,N_23867,N_23402);
nand UO_2250 (O_2250,N_23196,N_22947);
or UO_2251 (O_2251,N_22505,N_22575);
nand UO_2252 (O_2252,N_24970,N_23863);
or UO_2253 (O_2253,N_24826,N_22012);
or UO_2254 (O_2254,N_22025,N_22140);
and UO_2255 (O_2255,N_24825,N_24333);
nand UO_2256 (O_2256,N_23536,N_23623);
and UO_2257 (O_2257,N_22950,N_22560);
nand UO_2258 (O_2258,N_24084,N_24452);
nor UO_2259 (O_2259,N_24764,N_22223);
and UO_2260 (O_2260,N_22543,N_23112);
or UO_2261 (O_2261,N_23022,N_24918);
nand UO_2262 (O_2262,N_23362,N_23953);
or UO_2263 (O_2263,N_23115,N_24499);
nand UO_2264 (O_2264,N_22759,N_23260);
nor UO_2265 (O_2265,N_21917,N_22828);
nand UO_2266 (O_2266,N_24696,N_23007);
and UO_2267 (O_2267,N_22359,N_23639);
nor UO_2268 (O_2268,N_23186,N_24187);
and UO_2269 (O_2269,N_22762,N_23998);
or UO_2270 (O_2270,N_24222,N_24248);
nor UO_2271 (O_2271,N_24441,N_24814);
nor UO_2272 (O_2272,N_23929,N_24134);
nand UO_2273 (O_2273,N_23788,N_24377);
and UO_2274 (O_2274,N_23413,N_22203);
or UO_2275 (O_2275,N_22852,N_22872);
or UO_2276 (O_2276,N_22267,N_24077);
or UO_2277 (O_2277,N_23753,N_23113);
nor UO_2278 (O_2278,N_22295,N_22511);
and UO_2279 (O_2279,N_23669,N_21912);
nor UO_2280 (O_2280,N_22919,N_23317);
nor UO_2281 (O_2281,N_23003,N_22740);
or UO_2282 (O_2282,N_24021,N_24758);
or UO_2283 (O_2283,N_24408,N_23220);
or UO_2284 (O_2284,N_23470,N_23692);
or UO_2285 (O_2285,N_24660,N_23611);
and UO_2286 (O_2286,N_22573,N_22445);
or UO_2287 (O_2287,N_23894,N_22958);
nor UO_2288 (O_2288,N_23724,N_23775);
nor UO_2289 (O_2289,N_24252,N_23018);
nor UO_2290 (O_2290,N_23877,N_22639);
or UO_2291 (O_2291,N_23570,N_23114);
and UO_2292 (O_2292,N_22703,N_24163);
or UO_2293 (O_2293,N_22086,N_24554);
nor UO_2294 (O_2294,N_24689,N_24238);
xnor UO_2295 (O_2295,N_24470,N_23622);
nand UO_2296 (O_2296,N_23037,N_22916);
or UO_2297 (O_2297,N_23989,N_24969);
and UO_2298 (O_2298,N_23862,N_22945);
or UO_2299 (O_2299,N_23999,N_24958);
nor UO_2300 (O_2300,N_23538,N_24906);
and UO_2301 (O_2301,N_23566,N_22710);
and UO_2302 (O_2302,N_21889,N_23900);
nor UO_2303 (O_2303,N_22799,N_24315);
nor UO_2304 (O_2304,N_22601,N_24475);
and UO_2305 (O_2305,N_23725,N_23074);
nand UO_2306 (O_2306,N_23904,N_23076);
nor UO_2307 (O_2307,N_22366,N_23984);
and UO_2308 (O_2308,N_24794,N_24982);
nor UO_2309 (O_2309,N_23595,N_23793);
or UO_2310 (O_2310,N_21952,N_23941);
xor UO_2311 (O_2311,N_22216,N_24397);
or UO_2312 (O_2312,N_24221,N_24735);
or UO_2313 (O_2313,N_22649,N_22816);
and UO_2314 (O_2314,N_24879,N_23831);
or UO_2315 (O_2315,N_24969,N_22090);
nand UO_2316 (O_2316,N_24498,N_24217);
and UO_2317 (O_2317,N_22298,N_22140);
and UO_2318 (O_2318,N_23292,N_22085);
and UO_2319 (O_2319,N_22637,N_23080);
and UO_2320 (O_2320,N_23534,N_23107);
and UO_2321 (O_2321,N_23382,N_24409);
and UO_2322 (O_2322,N_22723,N_24675);
nor UO_2323 (O_2323,N_22990,N_23621);
nor UO_2324 (O_2324,N_21876,N_22899);
or UO_2325 (O_2325,N_22564,N_24190);
nand UO_2326 (O_2326,N_24901,N_22466);
and UO_2327 (O_2327,N_22196,N_22848);
nor UO_2328 (O_2328,N_23739,N_22070);
nand UO_2329 (O_2329,N_23194,N_23249);
and UO_2330 (O_2330,N_21966,N_23654);
or UO_2331 (O_2331,N_24740,N_23537);
or UO_2332 (O_2332,N_23128,N_22852);
nand UO_2333 (O_2333,N_23234,N_22690);
nand UO_2334 (O_2334,N_23096,N_23854);
or UO_2335 (O_2335,N_24415,N_23390);
nor UO_2336 (O_2336,N_23044,N_23050);
or UO_2337 (O_2337,N_23358,N_24808);
nor UO_2338 (O_2338,N_23718,N_23212);
or UO_2339 (O_2339,N_23520,N_23074);
nand UO_2340 (O_2340,N_22695,N_24284);
or UO_2341 (O_2341,N_24717,N_24672);
nor UO_2342 (O_2342,N_21988,N_23763);
or UO_2343 (O_2343,N_24635,N_22105);
nor UO_2344 (O_2344,N_24489,N_23931);
or UO_2345 (O_2345,N_23776,N_23563);
nand UO_2346 (O_2346,N_24622,N_22932);
or UO_2347 (O_2347,N_23203,N_24290);
and UO_2348 (O_2348,N_22227,N_21892);
nand UO_2349 (O_2349,N_23534,N_22519);
nor UO_2350 (O_2350,N_23366,N_22450);
and UO_2351 (O_2351,N_23361,N_23735);
xnor UO_2352 (O_2352,N_24302,N_22108);
or UO_2353 (O_2353,N_23627,N_23646);
xor UO_2354 (O_2354,N_24752,N_23575);
nand UO_2355 (O_2355,N_22885,N_22423);
nor UO_2356 (O_2356,N_24232,N_22246);
nand UO_2357 (O_2357,N_22867,N_22681);
nor UO_2358 (O_2358,N_24456,N_22806);
and UO_2359 (O_2359,N_24448,N_23478);
nor UO_2360 (O_2360,N_21933,N_23179);
or UO_2361 (O_2361,N_23596,N_24510);
nand UO_2362 (O_2362,N_22427,N_22347);
nor UO_2363 (O_2363,N_22607,N_24509);
or UO_2364 (O_2364,N_22014,N_23641);
or UO_2365 (O_2365,N_22118,N_22748);
or UO_2366 (O_2366,N_22868,N_23854);
or UO_2367 (O_2367,N_23952,N_23637);
or UO_2368 (O_2368,N_22767,N_22620);
nand UO_2369 (O_2369,N_22557,N_23388);
or UO_2370 (O_2370,N_24004,N_23593);
or UO_2371 (O_2371,N_22745,N_24143);
nand UO_2372 (O_2372,N_23885,N_24366);
nand UO_2373 (O_2373,N_23588,N_24587);
or UO_2374 (O_2374,N_23948,N_21951);
xnor UO_2375 (O_2375,N_22003,N_23708);
or UO_2376 (O_2376,N_24623,N_21900);
nand UO_2377 (O_2377,N_23307,N_24096);
and UO_2378 (O_2378,N_23872,N_23281);
nand UO_2379 (O_2379,N_22592,N_22959);
nor UO_2380 (O_2380,N_22537,N_24105);
nor UO_2381 (O_2381,N_22917,N_22184);
or UO_2382 (O_2382,N_22898,N_23307);
and UO_2383 (O_2383,N_23461,N_23420);
nor UO_2384 (O_2384,N_23042,N_22745);
nor UO_2385 (O_2385,N_22480,N_22531);
and UO_2386 (O_2386,N_22375,N_23476);
xor UO_2387 (O_2387,N_22203,N_24208);
xor UO_2388 (O_2388,N_24276,N_22344);
nor UO_2389 (O_2389,N_22752,N_24817);
nand UO_2390 (O_2390,N_22324,N_22578);
nand UO_2391 (O_2391,N_22792,N_22470);
or UO_2392 (O_2392,N_23464,N_22802);
nand UO_2393 (O_2393,N_22236,N_23541);
and UO_2394 (O_2394,N_23093,N_24440);
nand UO_2395 (O_2395,N_22997,N_22895);
nor UO_2396 (O_2396,N_22124,N_23321);
xor UO_2397 (O_2397,N_21917,N_22327);
xor UO_2398 (O_2398,N_24080,N_22099);
nor UO_2399 (O_2399,N_22994,N_24685);
and UO_2400 (O_2400,N_22460,N_24588);
or UO_2401 (O_2401,N_24262,N_24095);
nor UO_2402 (O_2402,N_23414,N_24587);
or UO_2403 (O_2403,N_24679,N_24828);
nand UO_2404 (O_2404,N_21947,N_24821);
nand UO_2405 (O_2405,N_24023,N_24545);
nand UO_2406 (O_2406,N_22526,N_23427);
and UO_2407 (O_2407,N_23526,N_21991);
nand UO_2408 (O_2408,N_22411,N_22102);
nand UO_2409 (O_2409,N_24482,N_24847);
nor UO_2410 (O_2410,N_24502,N_24279);
nor UO_2411 (O_2411,N_23638,N_23853);
xnor UO_2412 (O_2412,N_23600,N_23644);
or UO_2413 (O_2413,N_24967,N_24854);
or UO_2414 (O_2414,N_24229,N_23331);
nor UO_2415 (O_2415,N_23374,N_23238);
xor UO_2416 (O_2416,N_23874,N_23056);
nor UO_2417 (O_2417,N_24408,N_24288);
nand UO_2418 (O_2418,N_24806,N_24553);
or UO_2419 (O_2419,N_23911,N_22586);
and UO_2420 (O_2420,N_23401,N_23939);
or UO_2421 (O_2421,N_24971,N_22630);
nor UO_2422 (O_2422,N_24899,N_22979);
nor UO_2423 (O_2423,N_22354,N_23284);
nor UO_2424 (O_2424,N_23331,N_24554);
and UO_2425 (O_2425,N_22432,N_22073);
nor UO_2426 (O_2426,N_23740,N_21934);
xor UO_2427 (O_2427,N_22773,N_23633);
nand UO_2428 (O_2428,N_22229,N_22162);
nor UO_2429 (O_2429,N_22213,N_23235);
nand UO_2430 (O_2430,N_23895,N_22802);
nand UO_2431 (O_2431,N_22743,N_23708);
and UO_2432 (O_2432,N_22738,N_24702);
and UO_2433 (O_2433,N_23728,N_24278);
nor UO_2434 (O_2434,N_24955,N_24948);
or UO_2435 (O_2435,N_22877,N_22898);
and UO_2436 (O_2436,N_23683,N_22695);
and UO_2437 (O_2437,N_24893,N_22095);
nand UO_2438 (O_2438,N_22303,N_22198);
xor UO_2439 (O_2439,N_22471,N_24023);
or UO_2440 (O_2440,N_24199,N_23844);
nand UO_2441 (O_2441,N_24688,N_23068);
or UO_2442 (O_2442,N_22903,N_23390);
xor UO_2443 (O_2443,N_24780,N_22857);
or UO_2444 (O_2444,N_23859,N_23697);
nand UO_2445 (O_2445,N_24534,N_22854);
and UO_2446 (O_2446,N_23015,N_22687);
nor UO_2447 (O_2447,N_22934,N_24703);
nor UO_2448 (O_2448,N_23187,N_24965);
or UO_2449 (O_2449,N_23462,N_22489);
nor UO_2450 (O_2450,N_23815,N_24922);
or UO_2451 (O_2451,N_24137,N_22615);
nand UO_2452 (O_2452,N_22723,N_24738);
nor UO_2453 (O_2453,N_22107,N_24977);
or UO_2454 (O_2454,N_23114,N_24922);
or UO_2455 (O_2455,N_23903,N_24653);
xor UO_2456 (O_2456,N_23106,N_23059);
or UO_2457 (O_2457,N_24629,N_22015);
and UO_2458 (O_2458,N_24662,N_23534);
and UO_2459 (O_2459,N_24535,N_22723);
nand UO_2460 (O_2460,N_24301,N_23322);
nand UO_2461 (O_2461,N_22271,N_23548);
xnor UO_2462 (O_2462,N_24294,N_24529);
xnor UO_2463 (O_2463,N_22171,N_22892);
nand UO_2464 (O_2464,N_24926,N_24536);
nor UO_2465 (O_2465,N_23566,N_23938);
and UO_2466 (O_2466,N_23588,N_22981);
nor UO_2467 (O_2467,N_22283,N_22252);
xnor UO_2468 (O_2468,N_21986,N_24675);
nand UO_2469 (O_2469,N_24967,N_21898);
and UO_2470 (O_2470,N_23535,N_24383);
and UO_2471 (O_2471,N_22200,N_24493);
and UO_2472 (O_2472,N_23426,N_22528);
and UO_2473 (O_2473,N_24760,N_24021);
nand UO_2474 (O_2474,N_24787,N_23768);
nand UO_2475 (O_2475,N_22674,N_23276);
nor UO_2476 (O_2476,N_21907,N_23486);
or UO_2477 (O_2477,N_22443,N_24382);
or UO_2478 (O_2478,N_23441,N_23934);
or UO_2479 (O_2479,N_24169,N_23673);
xor UO_2480 (O_2480,N_21990,N_23130);
and UO_2481 (O_2481,N_22318,N_23178);
nor UO_2482 (O_2482,N_24738,N_22999);
and UO_2483 (O_2483,N_22745,N_22901);
or UO_2484 (O_2484,N_23926,N_24784);
nor UO_2485 (O_2485,N_24857,N_23600);
and UO_2486 (O_2486,N_23900,N_22455);
or UO_2487 (O_2487,N_22253,N_23868);
or UO_2488 (O_2488,N_23463,N_22719);
nand UO_2489 (O_2489,N_22676,N_24775);
nand UO_2490 (O_2490,N_24047,N_23931);
and UO_2491 (O_2491,N_24596,N_22977);
nand UO_2492 (O_2492,N_22369,N_24829);
or UO_2493 (O_2493,N_23039,N_24737);
nor UO_2494 (O_2494,N_23157,N_23769);
and UO_2495 (O_2495,N_23819,N_22326);
xnor UO_2496 (O_2496,N_23019,N_24718);
and UO_2497 (O_2497,N_24223,N_23699);
or UO_2498 (O_2498,N_22747,N_24915);
nand UO_2499 (O_2499,N_22279,N_23612);
or UO_2500 (O_2500,N_22084,N_22921);
xnor UO_2501 (O_2501,N_23608,N_23713);
or UO_2502 (O_2502,N_23402,N_24242);
and UO_2503 (O_2503,N_23500,N_22406);
nand UO_2504 (O_2504,N_23355,N_23249);
or UO_2505 (O_2505,N_23990,N_24855);
nor UO_2506 (O_2506,N_23839,N_22642);
or UO_2507 (O_2507,N_23236,N_24450);
or UO_2508 (O_2508,N_23384,N_24773);
nor UO_2509 (O_2509,N_23559,N_22456);
nand UO_2510 (O_2510,N_23984,N_22308);
or UO_2511 (O_2511,N_24545,N_22475);
or UO_2512 (O_2512,N_22616,N_21881);
nor UO_2513 (O_2513,N_23987,N_22133);
and UO_2514 (O_2514,N_23142,N_22533);
nor UO_2515 (O_2515,N_23836,N_23950);
nand UO_2516 (O_2516,N_23664,N_23053);
or UO_2517 (O_2517,N_22236,N_22766);
or UO_2518 (O_2518,N_24915,N_24755);
nor UO_2519 (O_2519,N_22275,N_24643);
or UO_2520 (O_2520,N_22606,N_23461);
or UO_2521 (O_2521,N_24928,N_23602);
and UO_2522 (O_2522,N_24121,N_23788);
nand UO_2523 (O_2523,N_24318,N_22260);
or UO_2524 (O_2524,N_24079,N_23541);
and UO_2525 (O_2525,N_23088,N_24900);
nor UO_2526 (O_2526,N_22470,N_23344);
and UO_2527 (O_2527,N_24085,N_23773);
nor UO_2528 (O_2528,N_24427,N_23621);
or UO_2529 (O_2529,N_23878,N_23521);
or UO_2530 (O_2530,N_22987,N_22044);
xnor UO_2531 (O_2531,N_22567,N_23150);
xnor UO_2532 (O_2532,N_24780,N_22341);
or UO_2533 (O_2533,N_24937,N_23955);
nand UO_2534 (O_2534,N_23202,N_24941);
nor UO_2535 (O_2535,N_22970,N_22174);
nor UO_2536 (O_2536,N_22304,N_24382);
nor UO_2537 (O_2537,N_22641,N_24639);
and UO_2538 (O_2538,N_24141,N_24912);
or UO_2539 (O_2539,N_23839,N_22926);
xor UO_2540 (O_2540,N_23260,N_22320);
nor UO_2541 (O_2541,N_23972,N_22651);
nor UO_2542 (O_2542,N_24709,N_23383);
nor UO_2543 (O_2543,N_24839,N_24217);
nor UO_2544 (O_2544,N_24160,N_22799);
nor UO_2545 (O_2545,N_24711,N_22538);
or UO_2546 (O_2546,N_23494,N_22342);
nor UO_2547 (O_2547,N_24701,N_23015);
nor UO_2548 (O_2548,N_24140,N_23558);
nand UO_2549 (O_2549,N_23352,N_24325);
xnor UO_2550 (O_2550,N_24258,N_23017);
nor UO_2551 (O_2551,N_22630,N_21901);
nand UO_2552 (O_2552,N_23690,N_24852);
or UO_2553 (O_2553,N_23232,N_24267);
nand UO_2554 (O_2554,N_24094,N_24941);
and UO_2555 (O_2555,N_22991,N_23386);
nor UO_2556 (O_2556,N_24711,N_24886);
nor UO_2557 (O_2557,N_23049,N_22510);
nand UO_2558 (O_2558,N_23931,N_23241);
nand UO_2559 (O_2559,N_22368,N_23948);
nor UO_2560 (O_2560,N_24600,N_23513);
xor UO_2561 (O_2561,N_23645,N_24470);
nand UO_2562 (O_2562,N_24314,N_22063);
and UO_2563 (O_2563,N_22730,N_22012);
or UO_2564 (O_2564,N_24730,N_23775);
or UO_2565 (O_2565,N_24297,N_24426);
nand UO_2566 (O_2566,N_23422,N_22489);
nand UO_2567 (O_2567,N_22507,N_22964);
and UO_2568 (O_2568,N_22815,N_24760);
and UO_2569 (O_2569,N_21910,N_23209);
xnor UO_2570 (O_2570,N_24479,N_23498);
nor UO_2571 (O_2571,N_23904,N_24540);
or UO_2572 (O_2572,N_22747,N_22204);
xor UO_2573 (O_2573,N_24389,N_22601);
or UO_2574 (O_2574,N_23526,N_24476);
nand UO_2575 (O_2575,N_21916,N_22716);
and UO_2576 (O_2576,N_22142,N_23023);
nor UO_2577 (O_2577,N_24900,N_23534);
nand UO_2578 (O_2578,N_23915,N_24954);
nand UO_2579 (O_2579,N_22718,N_24522);
or UO_2580 (O_2580,N_24272,N_23408);
nor UO_2581 (O_2581,N_22657,N_24735);
and UO_2582 (O_2582,N_24539,N_24895);
nor UO_2583 (O_2583,N_22974,N_24373);
and UO_2584 (O_2584,N_22069,N_23526);
nand UO_2585 (O_2585,N_22163,N_23478);
nor UO_2586 (O_2586,N_24636,N_22736);
nand UO_2587 (O_2587,N_22143,N_22938);
xor UO_2588 (O_2588,N_23202,N_23628);
nand UO_2589 (O_2589,N_24796,N_24662);
nor UO_2590 (O_2590,N_23997,N_21926);
and UO_2591 (O_2591,N_23948,N_24875);
nor UO_2592 (O_2592,N_21953,N_23348);
nor UO_2593 (O_2593,N_24545,N_24865);
or UO_2594 (O_2594,N_23138,N_22987);
and UO_2595 (O_2595,N_24951,N_22655);
and UO_2596 (O_2596,N_21881,N_24184);
xnor UO_2597 (O_2597,N_23112,N_24083);
or UO_2598 (O_2598,N_22547,N_23198);
or UO_2599 (O_2599,N_24482,N_22805);
nor UO_2600 (O_2600,N_24583,N_22187);
or UO_2601 (O_2601,N_24235,N_24862);
nor UO_2602 (O_2602,N_23350,N_23603);
nor UO_2603 (O_2603,N_22836,N_24385);
nand UO_2604 (O_2604,N_22246,N_24096);
or UO_2605 (O_2605,N_22083,N_23288);
or UO_2606 (O_2606,N_22181,N_22383);
and UO_2607 (O_2607,N_22738,N_24822);
or UO_2608 (O_2608,N_22419,N_22292);
nor UO_2609 (O_2609,N_24876,N_24563);
nor UO_2610 (O_2610,N_23031,N_24031);
or UO_2611 (O_2611,N_24009,N_24725);
and UO_2612 (O_2612,N_23141,N_22828);
and UO_2613 (O_2613,N_21910,N_22974);
nor UO_2614 (O_2614,N_24290,N_22992);
or UO_2615 (O_2615,N_22213,N_22763);
nand UO_2616 (O_2616,N_22351,N_22034);
or UO_2617 (O_2617,N_24921,N_24911);
nor UO_2618 (O_2618,N_23242,N_24488);
or UO_2619 (O_2619,N_23128,N_22097);
or UO_2620 (O_2620,N_22764,N_23454);
and UO_2621 (O_2621,N_23177,N_22127);
nand UO_2622 (O_2622,N_22321,N_23093);
nand UO_2623 (O_2623,N_22874,N_22550);
nor UO_2624 (O_2624,N_23307,N_24884);
nand UO_2625 (O_2625,N_22773,N_23550);
or UO_2626 (O_2626,N_24598,N_22464);
nand UO_2627 (O_2627,N_22768,N_24579);
xor UO_2628 (O_2628,N_24186,N_23658);
or UO_2629 (O_2629,N_24171,N_24768);
nand UO_2630 (O_2630,N_22139,N_23527);
and UO_2631 (O_2631,N_23189,N_24552);
or UO_2632 (O_2632,N_24731,N_24693);
and UO_2633 (O_2633,N_24137,N_24643);
nor UO_2634 (O_2634,N_24692,N_23656);
or UO_2635 (O_2635,N_24157,N_24959);
and UO_2636 (O_2636,N_23166,N_22949);
and UO_2637 (O_2637,N_24416,N_23020);
or UO_2638 (O_2638,N_22463,N_24243);
nand UO_2639 (O_2639,N_22770,N_22252);
and UO_2640 (O_2640,N_22096,N_24393);
nor UO_2641 (O_2641,N_24029,N_24135);
or UO_2642 (O_2642,N_24308,N_24355);
nor UO_2643 (O_2643,N_23512,N_22264);
nand UO_2644 (O_2644,N_24447,N_22361);
nand UO_2645 (O_2645,N_23017,N_23248);
nand UO_2646 (O_2646,N_23168,N_22747);
and UO_2647 (O_2647,N_24467,N_23635);
nand UO_2648 (O_2648,N_21962,N_22927);
nand UO_2649 (O_2649,N_23636,N_24945);
or UO_2650 (O_2650,N_23939,N_22908);
xor UO_2651 (O_2651,N_23279,N_22251);
nor UO_2652 (O_2652,N_24070,N_22401);
nor UO_2653 (O_2653,N_22992,N_23450);
xnor UO_2654 (O_2654,N_23998,N_24492);
or UO_2655 (O_2655,N_21899,N_24552);
or UO_2656 (O_2656,N_22646,N_22690);
nand UO_2657 (O_2657,N_24111,N_22359);
nor UO_2658 (O_2658,N_23892,N_22144);
nor UO_2659 (O_2659,N_22198,N_23354);
nand UO_2660 (O_2660,N_24238,N_22341);
nand UO_2661 (O_2661,N_22744,N_23241);
nor UO_2662 (O_2662,N_24201,N_22983);
or UO_2663 (O_2663,N_21960,N_24992);
or UO_2664 (O_2664,N_23566,N_22504);
nand UO_2665 (O_2665,N_22602,N_24538);
or UO_2666 (O_2666,N_24842,N_22314);
nor UO_2667 (O_2667,N_22679,N_24859);
xnor UO_2668 (O_2668,N_23126,N_23190);
or UO_2669 (O_2669,N_22042,N_24911);
or UO_2670 (O_2670,N_23169,N_23832);
nand UO_2671 (O_2671,N_22029,N_22088);
nand UO_2672 (O_2672,N_23415,N_23236);
and UO_2673 (O_2673,N_23163,N_24145);
xor UO_2674 (O_2674,N_23639,N_22651);
nand UO_2675 (O_2675,N_22276,N_24825);
or UO_2676 (O_2676,N_24957,N_24275);
and UO_2677 (O_2677,N_22416,N_22663);
and UO_2678 (O_2678,N_23875,N_23658);
nor UO_2679 (O_2679,N_24727,N_23127);
nand UO_2680 (O_2680,N_24745,N_23163);
and UO_2681 (O_2681,N_22266,N_24971);
nand UO_2682 (O_2682,N_24263,N_23608);
xor UO_2683 (O_2683,N_22001,N_24563);
and UO_2684 (O_2684,N_23181,N_22380);
nor UO_2685 (O_2685,N_23667,N_23173);
and UO_2686 (O_2686,N_22467,N_24157);
nand UO_2687 (O_2687,N_23272,N_24354);
nor UO_2688 (O_2688,N_23634,N_21962);
xor UO_2689 (O_2689,N_24100,N_21894);
or UO_2690 (O_2690,N_23813,N_23602);
xor UO_2691 (O_2691,N_22047,N_23972);
and UO_2692 (O_2692,N_24301,N_22223);
xnor UO_2693 (O_2693,N_23682,N_24167);
or UO_2694 (O_2694,N_22882,N_23048);
and UO_2695 (O_2695,N_23662,N_24675);
and UO_2696 (O_2696,N_22246,N_21884);
or UO_2697 (O_2697,N_22332,N_22492);
nor UO_2698 (O_2698,N_24339,N_21975);
nor UO_2699 (O_2699,N_24459,N_21889);
xor UO_2700 (O_2700,N_23694,N_24699);
nor UO_2701 (O_2701,N_21962,N_21912);
xnor UO_2702 (O_2702,N_23837,N_23553);
nor UO_2703 (O_2703,N_22120,N_22755);
or UO_2704 (O_2704,N_22590,N_23077);
nand UO_2705 (O_2705,N_24530,N_22777);
and UO_2706 (O_2706,N_24246,N_24857);
nor UO_2707 (O_2707,N_22713,N_22198);
nand UO_2708 (O_2708,N_24460,N_24916);
nor UO_2709 (O_2709,N_24525,N_23831);
or UO_2710 (O_2710,N_23369,N_23372);
nand UO_2711 (O_2711,N_23640,N_23765);
or UO_2712 (O_2712,N_22325,N_22309);
and UO_2713 (O_2713,N_23502,N_22919);
nor UO_2714 (O_2714,N_23912,N_22185);
nand UO_2715 (O_2715,N_24410,N_23890);
nand UO_2716 (O_2716,N_24932,N_23001);
and UO_2717 (O_2717,N_24085,N_22824);
or UO_2718 (O_2718,N_23454,N_24801);
and UO_2719 (O_2719,N_24747,N_24836);
and UO_2720 (O_2720,N_23608,N_23838);
or UO_2721 (O_2721,N_23114,N_22555);
nor UO_2722 (O_2722,N_22224,N_24649);
nor UO_2723 (O_2723,N_22750,N_22143);
nor UO_2724 (O_2724,N_22095,N_24536);
and UO_2725 (O_2725,N_22567,N_24275);
and UO_2726 (O_2726,N_23640,N_22804);
xnor UO_2727 (O_2727,N_22806,N_24232);
and UO_2728 (O_2728,N_23477,N_22156);
nor UO_2729 (O_2729,N_22544,N_24745);
or UO_2730 (O_2730,N_24732,N_22443);
or UO_2731 (O_2731,N_23608,N_22017);
and UO_2732 (O_2732,N_24235,N_24860);
or UO_2733 (O_2733,N_22926,N_24527);
or UO_2734 (O_2734,N_24410,N_22192);
xor UO_2735 (O_2735,N_21934,N_24592);
nor UO_2736 (O_2736,N_24564,N_24129);
nand UO_2737 (O_2737,N_24539,N_23727);
or UO_2738 (O_2738,N_23977,N_23309);
nor UO_2739 (O_2739,N_24158,N_24582);
nand UO_2740 (O_2740,N_23403,N_24655);
nand UO_2741 (O_2741,N_22773,N_24633);
nand UO_2742 (O_2742,N_23882,N_23403);
and UO_2743 (O_2743,N_23015,N_23139);
nand UO_2744 (O_2744,N_24421,N_23248);
nor UO_2745 (O_2745,N_23234,N_24069);
xor UO_2746 (O_2746,N_23028,N_24872);
or UO_2747 (O_2747,N_23999,N_23117);
and UO_2748 (O_2748,N_23006,N_24812);
nor UO_2749 (O_2749,N_21934,N_23258);
nor UO_2750 (O_2750,N_23324,N_22245);
xnor UO_2751 (O_2751,N_23555,N_22515);
or UO_2752 (O_2752,N_22869,N_23564);
and UO_2753 (O_2753,N_23848,N_24633);
nor UO_2754 (O_2754,N_22029,N_22853);
nand UO_2755 (O_2755,N_22637,N_23514);
nand UO_2756 (O_2756,N_22405,N_22762);
xnor UO_2757 (O_2757,N_22068,N_22295);
or UO_2758 (O_2758,N_22118,N_23841);
nand UO_2759 (O_2759,N_22942,N_23443);
xnor UO_2760 (O_2760,N_24384,N_23416);
or UO_2761 (O_2761,N_22151,N_22114);
nor UO_2762 (O_2762,N_24480,N_24944);
and UO_2763 (O_2763,N_23647,N_23609);
or UO_2764 (O_2764,N_24019,N_24888);
nand UO_2765 (O_2765,N_23195,N_24423);
nand UO_2766 (O_2766,N_22913,N_23724);
or UO_2767 (O_2767,N_23942,N_23866);
nor UO_2768 (O_2768,N_22415,N_24974);
and UO_2769 (O_2769,N_24914,N_22514);
and UO_2770 (O_2770,N_23938,N_22815);
nor UO_2771 (O_2771,N_23671,N_22910);
or UO_2772 (O_2772,N_24622,N_22922);
nor UO_2773 (O_2773,N_23460,N_24900);
nand UO_2774 (O_2774,N_22406,N_24056);
nand UO_2775 (O_2775,N_21931,N_24466);
nand UO_2776 (O_2776,N_23096,N_23627);
and UO_2777 (O_2777,N_22780,N_23695);
nor UO_2778 (O_2778,N_23994,N_24459);
or UO_2779 (O_2779,N_21876,N_24648);
and UO_2780 (O_2780,N_23201,N_24037);
and UO_2781 (O_2781,N_24243,N_23618);
nand UO_2782 (O_2782,N_22199,N_24489);
xnor UO_2783 (O_2783,N_23529,N_23889);
nor UO_2784 (O_2784,N_24829,N_23460);
or UO_2785 (O_2785,N_21889,N_22125);
nand UO_2786 (O_2786,N_23419,N_24618);
nor UO_2787 (O_2787,N_23177,N_24380);
and UO_2788 (O_2788,N_22758,N_22340);
xor UO_2789 (O_2789,N_24370,N_24093);
xor UO_2790 (O_2790,N_24942,N_22542);
and UO_2791 (O_2791,N_22594,N_23216);
or UO_2792 (O_2792,N_23318,N_22253);
xor UO_2793 (O_2793,N_22040,N_24763);
or UO_2794 (O_2794,N_23862,N_22947);
nand UO_2795 (O_2795,N_23645,N_22143);
or UO_2796 (O_2796,N_23837,N_23525);
xnor UO_2797 (O_2797,N_23171,N_21996);
or UO_2798 (O_2798,N_24891,N_22971);
and UO_2799 (O_2799,N_22970,N_22654);
nor UO_2800 (O_2800,N_23834,N_22937);
xnor UO_2801 (O_2801,N_22758,N_22081);
or UO_2802 (O_2802,N_23866,N_23148);
and UO_2803 (O_2803,N_22210,N_23584);
xor UO_2804 (O_2804,N_24490,N_23593);
nand UO_2805 (O_2805,N_24548,N_23488);
and UO_2806 (O_2806,N_22795,N_24949);
or UO_2807 (O_2807,N_23379,N_23928);
and UO_2808 (O_2808,N_23571,N_23710);
or UO_2809 (O_2809,N_24218,N_23867);
and UO_2810 (O_2810,N_24262,N_24816);
and UO_2811 (O_2811,N_22600,N_23236);
nand UO_2812 (O_2812,N_22414,N_24786);
and UO_2813 (O_2813,N_22101,N_22666);
nor UO_2814 (O_2814,N_23303,N_23886);
and UO_2815 (O_2815,N_24958,N_24456);
and UO_2816 (O_2816,N_23101,N_22197);
xnor UO_2817 (O_2817,N_23734,N_24758);
and UO_2818 (O_2818,N_22686,N_24265);
nor UO_2819 (O_2819,N_22859,N_22003);
nand UO_2820 (O_2820,N_23167,N_22202);
xor UO_2821 (O_2821,N_22704,N_23314);
nand UO_2822 (O_2822,N_22738,N_22404);
or UO_2823 (O_2823,N_22985,N_22010);
or UO_2824 (O_2824,N_22322,N_21901);
and UO_2825 (O_2825,N_22406,N_24656);
or UO_2826 (O_2826,N_23479,N_24474);
nand UO_2827 (O_2827,N_23058,N_24167);
nand UO_2828 (O_2828,N_24181,N_22532);
and UO_2829 (O_2829,N_22278,N_22298);
and UO_2830 (O_2830,N_23542,N_23220);
and UO_2831 (O_2831,N_22570,N_22838);
and UO_2832 (O_2832,N_24293,N_22374);
nor UO_2833 (O_2833,N_21876,N_22501);
and UO_2834 (O_2834,N_21887,N_23403);
or UO_2835 (O_2835,N_24414,N_24142);
or UO_2836 (O_2836,N_23675,N_22959);
nand UO_2837 (O_2837,N_23327,N_23870);
nand UO_2838 (O_2838,N_24826,N_24641);
nor UO_2839 (O_2839,N_23142,N_23238);
or UO_2840 (O_2840,N_23130,N_23299);
and UO_2841 (O_2841,N_24376,N_23211);
or UO_2842 (O_2842,N_22800,N_23217);
nor UO_2843 (O_2843,N_24688,N_22852);
and UO_2844 (O_2844,N_23660,N_22531);
or UO_2845 (O_2845,N_22864,N_24982);
nor UO_2846 (O_2846,N_23815,N_23493);
and UO_2847 (O_2847,N_23359,N_22433);
or UO_2848 (O_2848,N_24132,N_22375);
and UO_2849 (O_2849,N_23063,N_23952);
or UO_2850 (O_2850,N_22611,N_24139);
xor UO_2851 (O_2851,N_24580,N_24268);
nand UO_2852 (O_2852,N_24936,N_23048);
and UO_2853 (O_2853,N_22377,N_23679);
nand UO_2854 (O_2854,N_22444,N_24155);
nand UO_2855 (O_2855,N_23194,N_23592);
nand UO_2856 (O_2856,N_21936,N_24910);
and UO_2857 (O_2857,N_24846,N_23009);
or UO_2858 (O_2858,N_23340,N_24079);
or UO_2859 (O_2859,N_23549,N_23447);
nand UO_2860 (O_2860,N_22916,N_23178);
nand UO_2861 (O_2861,N_23506,N_24427);
nand UO_2862 (O_2862,N_23117,N_24847);
and UO_2863 (O_2863,N_22027,N_22053);
nand UO_2864 (O_2864,N_24079,N_22045);
or UO_2865 (O_2865,N_22745,N_24133);
nor UO_2866 (O_2866,N_23154,N_24837);
or UO_2867 (O_2867,N_22859,N_22004);
or UO_2868 (O_2868,N_24324,N_24055);
nand UO_2869 (O_2869,N_22123,N_23464);
xor UO_2870 (O_2870,N_24402,N_23164);
and UO_2871 (O_2871,N_24262,N_22906);
or UO_2872 (O_2872,N_23406,N_22076);
and UO_2873 (O_2873,N_22769,N_22687);
nor UO_2874 (O_2874,N_24097,N_22262);
or UO_2875 (O_2875,N_23507,N_22495);
or UO_2876 (O_2876,N_21917,N_24251);
and UO_2877 (O_2877,N_23306,N_24890);
nor UO_2878 (O_2878,N_23908,N_24940);
and UO_2879 (O_2879,N_23869,N_24446);
or UO_2880 (O_2880,N_22498,N_23160);
nor UO_2881 (O_2881,N_22304,N_22524);
and UO_2882 (O_2882,N_22915,N_22391);
and UO_2883 (O_2883,N_23060,N_23481);
nor UO_2884 (O_2884,N_22509,N_24928);
and UO_2885 (O_2885,N_24366,N_22475);
nand UO_2886 (O_2886,N_23773,N_23415);
nor UO_2887 (O_2887,N_23609,N_24871);
nor UO_2888 (O_2888,N_23352,N_23326);
xnor UO_2889 (O_2889,N_22288,N_23774);
and UO_2890 (O_2890,N_24308,N_22244);
nor UO_2891 (O_2891,N_23753,N_24961);
or UO_2892 (O_2892,N_22226,N_23505);
or UO_2893 (O_2893,N_24436,N_22064);
and UO_2894 (O_2894,N_24354,N_23138);
nor UO_2895 (O_2895,N_23399,N_22205);
nor UO_2896 (O_2896,N_22860,N_22018);
nor UO_2897 (O_2897,N_23928,N_24867);
nor UO_2898 (O_2898,N_24336,N_23014);
nor UO_2899 (O_2899,N_22799,N_24188);
and UO_2900 (O_2900,N_23191,N_24240);
and UO_2901 (O_2901,N_23955,N_22875);
nand UO_2902 (O_2902,N_24802,N_24423);
and UO_2903 (O_2903,N_22625,N_21976);
and UO_2904 (O_2904,N_24501,N_24181);
and UO_2905 (O_2905,N_24734,N_24299);
nor UO_2906 (O_2906,N_22132,N_23360);
or UO_2907 (O_2907,N_23932,N_23669);
nand UO_2908 (O_2908,N_24807,N_22662);
and UO_2909 (O_2909,N_24390,N_22308);
or UO_2910 (O_2910,N_24622,N_23931);
or UO_2911 (O_2911,N_23371,N_22939);
or UO_2912 (O_2912,N_24439,N_23229);
nand UO_2913 (O_2913,N_22729,N_23644);
nor UO_2914 (O_2914,N_23342,N_22640);
nor UO_2915 (O_2915,N_22453,N_22682);
and UO_2916 (O_2916,N_23720,N_24728);
and UO_2917 (O_2917,N_24497,N_24226);
nor UO_2918 (O_2918,N_22365,N_24926);
and UO_2919 (O_2919,N_23940,N_24657);
nor UO_2920 (O_2920,N_23756,N_23452);
and UO_2921 (O_2921,N_24361,N_23714);
xnor UO_2922 (O_2922,N_23843,N_24425);
or UO_2923 (O_2923,N_24110,N_24678);
or UO_2924 (O_2924,N_23552,N_22805);
or UO_2925 (O_2925,N_24929,N_23168);
xor UO_2926 (O_2926,N_24955,N_22358);
or UO_2927 (O_2927,N_24365,N_22590);
nand UO_2928 (O_2928,N_24475,N_23212);
nand UO_2929 (O_2929,N_22783,N_24671);
or UO_2930 (O_2930,N_22538,N_23422);
nand UO_2931 (O_2931,N_21975,N_23133);
nand UO_2932 (O_2932,N_22653,N_22943);
nor UO_2933 (O_2933,N_22256,N_23037);
nand UO_2934 (O_2934,N_23564,N_22527);
nor UO_2935 (O_2935,N_23576,N_21894);
nand UO_2936 (O_2936,N_22660,N_24742);
nor UO_2937 (O_2937,N_24767,N_21948);
or UO_2938 (O_2938,N_23091,N_24581);
nand UO_2939 (O_2939,N_24769,N_23490);
nor UO_2940 (O_2940,N_22978,N_21991);
nor UO_2941 (O_2941,N_22313,N_23539);
nand UO_2942 (O_2942,N_24816,N_24735);
nand UO_2943 (O_2943,N_23880,N_22013);
or UO_2944 (O_2944,N_24876,N_22293);
and UO_2945 (O_2945,N_22404,N_22774);
xor UO_2946 (O_2946,N_22542,N_24724);
and UO_2947 (O_2947,N_24213,N_24981);
nor UO_2948 (O_2948,N_22068,N_24471);
nand UO_2949 (O_2949,N_24731,N_22534);
or UO_2950 (O_2950,N_24657,N_22534);
nor UO_2951 (O_2951,N_23152,N_24070);
or UO_2952 (O_2952,N_24325,N_22969);
or UO_2953 (O_2953,N_23902,N_24577);
nand UO_2954 (O_2954,N_23271,N_22803);
nand UO_2955 (O_2955,N_24873,N_22904);
and UO_2956 (O_2956,N_23695,N_23991);
nand UO_2957 (O_2957,N_23865,N_24532);
or UO_2958 (O_2958,N_22714,N_24139);
or UO_2959 (O_2959,N_24560,N_23081);
or UO_2960 (O_2960,N_22925,N_23894);
nor UO_2961 (O_2961,N_22502,N_22333);
and UO_2962 (O_2962,N_21912,N_23467);
nand UO_2963 (O_2963,N_23609,N_24556);
nor UO_2964 (O_2964,N_23207,N_23901);
nor UO_2965 (O_2965,N_24652,N_22924);
and UO_2966 (O_2966,N_23541,N_22400);
nor UO_2967 (O_2967,N_23931,N_23299);
nand UO_2968 (O_2968,N_21962,N_22550);
xor UO_2969 (O_2969,N_22290,N_24160);
and UO_2970 (O_2970,N_23631,N_23653);
and UO_2971 (O_2971,N_24304,N_23520);
or UO_2972 (O_2972,N_24892,N_21955);
nand UO_2973 (O_2973,N_24463,N_21933);
nor UO_2974 (O_2974,N_24248,N_23946);
and UO_2975 (O_2975,N_24259,N_23090);
nand UO_2976 (O_2976,N_24942,N_23629);
or UO_2977 (O_2977,N_24968,N_23687);
and UO_2978 (O_2978,N_22610,N_22473);
or UO_2979 (O_2979,N_22541,N_24447);
nand UO_2980 (O_2980,N_24936,N_22646);
nor UO_2981 (O_2981,N_23602,N_23608);
nor UO_2982 (O_2982,N_23412,N_22719);
or UO_2983 (O_2983,N_24135,N_22299);
or UO_2984 (O_2984,N_22430,N_23049);
nor UO_2985 (O_2985,N_22982,N_23845);
and UO_2986 (O_2986,N_22249,N_22742);
and UO_2987 (O_2987,N_22588,N_24385);
xnor UO_2988 (O_2988,N_21880,N_22734);
nor UO_2989 (O_2989,N_23966,N_24667);
nand UO_2990 (O_2990,N_22333,N_22230);
nand UO_2991 (O_2991,N_22619,N_22939);
or UO_2992 (O_2992,N_24047,N_22359);
nor UO_2993 (O_2993,N_22537,N_23609);
nor UO_2994 (O_2994,N_22768,N_24790);
or UO_2995 (O_2995,N_22570,N_24694);
and UO_2996 (O_2996,N_22122,N_24351);
nor UO_2997 (O_2997,N_23370,N_24372);
and UO_2998 (O_2998,N_22359,N_23332);
and UO_2999 (O_2999,N_24698,N_23811);
endmodule