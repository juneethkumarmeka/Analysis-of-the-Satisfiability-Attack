module basic_1500_15000_2000_60_levels_5xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_1331,In_560);
nand U1 (N_1,In_1468,In_874);
and U2 (N_2,In_162,In_700);
and U3 (N_3,In_173,In_1172);
or U4 (N_4,In_774,In_835);
and U5 (N_5,In_1350,In_40);
nand U6 (N_6,In_260,In_799);
and U7 (N_7,In_812,In_531);
and U8 (N_8,In_653,In_1335);
or U9 (N_9,In_636,In_332);
and U10 (N_10,In_570,In_1240);
nand U11 (N_11,In_1090,In_809);
and U12 (N_12,In_578,In_575);
xnor U13 (N_13,In_280,In_879);
nand U14 (N_14,In_655,In_859);
nor U15 (N_15,In_1360,In_480);
and U16 (N_16,In_1388,In_20);
xnor U17 (N_17,In_338,In_768);
and U18 (N_18,In_1216,In_1481);
nand U19 (N_19,In_400,In_72);
or U20 (N_20,In_42,In_968);
or U21 (N_21,In_1249,In_194);
or U22 (N_22,In_600,In_702);
and U23 (N_23,In_329,In_439);
nand U24 (N_24,In_287,In_839);
nor U25 (N_25,In_16,In_448);
nand U26 (N_26,In_89,In_668);
or U27 (N_27,In_1494,In_84);
and U28 (N_28,In_1395,In_221);
nor U29 (N_29,In_973,In_142);
nor U30 (N_30,In_550,In_340);
nor U31 (N_31,In_723,In_1265);
nor U32 (N_32,In_820,In_766);
nor U33 (N_33,In_1327,In_241);
and U34 (N_34,In_395,In_709);
nand U35 (N_35,In_326,In_1186);
nor U36 (N_36,In_518,In_313);
and U37 (N_37,In_1378,In_713);
nor U38 (N_38,In_154,In_236);
nand U39 (N_39,In_145,In_232);
nand U40 (N_40,In_424,In_905);
nand U41 (N_41,In_1351,In_1349);
xor U42 (N_42,In_180,In_1269);
nand U43 (N_43,In_673,In_649);
nand U44 (N_44,In_936,In_698);
nor U45 (N_45,In_1021,In_354);
nor U46 (N_46,In_1165,In_867);
nor U47 (N_47,In_735,In_422);
nand U48 (N_48,In_239,In_383);
or U49 (N_49,In_1044,In_117);
xor U50 (N_50,In_265,In_467);
xor U51 (N_51,In_1211,In_1347);
or U52 (N_52,In_171,In_1342);
and U53 (N_53,In_1278,In_670);
nand U54 (N_54,In_681,In_1092);
and U55 (N_55,In_24,In_127);
xor U56 (N_56,In_858,In_1079);
nand U57 (N_57,In_219,In_6);
and U58 (N_58,In_780,In_710);
nand U59 (N_59,In_302,In_815);
or U60 (N_60,In_1073,In_1287);
and U61 (N_61,In_996,In_1045);
and U62 (N_62,In_598,In_1141);
nand U63 (N_63,In_1416,In_394);
and U64 (N_64,In_626,In_955);
or U65 (N_65,In_1406,In_293);
nor U66 (N_66,In_1352,In_992);
and U67 (N_67,In_793,In_421);
nand U68 (N_68,In_2,In_1422);
or U69 (N_69,In_1066,In_1322);
xor U70 (N_70,In_167,In_149);
xnor U71 (N_71,In_1376,In_747);
and U72 (N_72,In_634,In_44);
nor U73 (N_73,In_1285,In_1194);
or U74 (N_74,In_1267,In_10);
or U75 (N_75,In_1030,In_1438);
nand U76 (N_76,In_1482,In_1131);
nand U77 (N_77,In_915,In_25);
or U78 (N_78,In_1324,In_918);
and U79 (N_79,In_984,In_1384);
nand U80 (N_80,In_386,In_1332);
and U81 (N_81,In_899,In_1158);
nor U82 (N_82,In_868,In_1389);
nand U83 (N_83,In_1370,In_853);
nand U84 (N_84,In_621,In_1022);
nor U85 (N_85,In_1358,In_869);
and U86 (N_86,In_91,In_1355);
or U87 (N_87,In_113,In_695);
nor U88 (N_88,In_1181,In_997);
nand U89 (N_89,In_453,In_1371);
nand U90 (N_90,In_1225,In_790);
xnor U91 (N_91,In_1493,In_1444);
and U92 (N_92,In_295,In_1190);
nand U93 (N_93,In_1036,In_216);
or U94 (N_94,In_530,In_100);
and U95 (N_95,In_322,In_160);
or U96 (N_96,In_958,In_398);
and U97 (N_97,In_1268,In_848);
nand U98 (N_98,In_498,In_916);
nor U99 (N_99,In_660,In_851);
xnor U100 (N_100,In_586,In_1374);
nor U101 (N_101,In_910,In_515);
or U102 (N_102,In_588,In_526);
nand U103 (N_103,In_310,In_1424);
xnor U104 (N_104,In_164,In_240);
or U105 (N_105,In_805,In_615);
or U106 (N_106,In_985,In_837);
or U107 (N_107,In_8,In_94);
or U108 (N_108,In_405,In_499);
and U109 (N_109,In_646,In_64);
nand U110 (N_110,In_1011,In_857);
or U111 (N_111,In_696,In_546);
nand U112 (N_112,In_654,In_1043);
nor U113 (N_113,In_836,In_1382);
nor U114 (N_114,In_23,In_407);
and U115 (N_115,In_103,In_979);
or U116 (N_116,In_462,In_388);
or U117 (N_117,In_500,In_775);
xor U118 (N_118,In_244,In_903);
or U119 (N_119,In_311,In_408);
nor U120 (N_120,In_174,In_1058);
nor U121 (N_121,In_1139,In_28);
nand U122 (N_122,In_687,In_108);
and U123 (N_123,In_1298,In_427);
or U124 (N_124,In_343,In_344);
or U125 (N_125,In_157,In_524);
xor U126 (N_126,In_1257,In_949);
nor U127 (N_127,In_1193,In_933);
and U128 (N_128,In_1230,In_1333);
or U129 (N_129,In_352,In_350);
or U130 (N_130,In_946,In_252);
or U131 (N_131,In_1323,In_596);
or U132 (N_132,In_1032,In_935);
xor U133 (N_133,In_1297,In_1274);
or U134 (N_134,In_489,In_337);
nor U135 (N_135,In_1235,In_704);
nor U136 (N_136,In_827,In_1238);
nand U137 (N_137,In_952,In_1487);
or U138 (N_138,In_685,In_963);
or U139 (N_139,In_986,In_1288);
or U140 (N_140,In_1227,In_902);
nor U141 (N_141,In_889,In_671);
or U142 (N_142,In_819,In_658);
nand U143 (N_143,In_732,In_1033);
nand U144 (N_144,In_107,In_34);
and U145 (N_145,In_1078,In_1334);
or U146 (N_146,In_866,In_118);
nand U147 (N_147,In_576,In_291);
or U148 (N_148,In_1229,In_301);
nand U149 (N_149,In_177,In_1310);
and U150 (N_150,In_559,In_82);
nand U151 (N_151,In_1222,In_940);
xnor U152 (N_152,In_186,In_442);
nor U153 (N_153,In_122,In_151);
nor U154 (N_154,In_503,In_1166);
nor U155 (N_155,In_268,In_966);
nand U156 (N_156,In_729,In_604);
nor U157 (N_157,In_939,In_1242);
nand U158 (N_158,In_921,In_415);
and U159 (N_159,In_1375,In_1280);
and U160 (N_160,In_169,In_431);
xnor U161 (N_161,In_248,In_676);
and U162 (N_162,In_189,In_1050);
nand U163 (N_163,In_445,In_1425);
and U164 (N_164,In_1113,In_476);
and U165 (N_165,In_571,In_823);
nor U166 (N_166,In_464,In_657);
nor U167 (N_167,In_843,In_458);
and U168 (N_168,In_981,In_254);
and U169 (N_169,In_587,In_229);
and U170 (N_170,In_284,In_41);
or U171 (N_171,In_1233,In_1248);
or U172 (N_172,In_624,In_614);
and U173 (N_173,In_1049,In_788);
or U174 (N_174,In_1137,In_1122);
nand U175 (N_175,In_1452,In_1127);
or U176 (N_176,In_286,In_1364);
and U177 (N_177,In_1489,In_1266);
xnor U178 (N_178,In_1289,In_250);
nand U179 (N_179,In_1053,In_926);
nor U180 (N_180,In_1423,In_893);
nand U181 (N_181,In_369,In_97);
nand U182 (N_182,In_510,In_1448);
or U183 (N_183,In_787,In_817);
nor U184 (N_184,In_368,In_1029);
nor U185 (N_185,In_1302,In_930);
and U186 (N_186,In_1463,In_730);
nor U187 (N_187,In_1219,In_237);
and U188 (N_188,In_502,In_1234);
nor U189 (N_189,In_758,In_150);
nand U190 (N_190,In_594,In_1074);
or U191 (N_191,In_456,In_1420);
nor U192 (N_192,In_1136,In_1415);
and U193 (N_193,In_374,In_243);
nand U194 (N_194,In_1069,In_1001);
nand U195 (N_195,In_102,In_539);
or U196 (N_196,In_290,In_1407);
nor U197 (N_197,In_1381,In_473);
xnor U198 (N_198,In_1457,In_607);
xnor U199 (N_199,In_534,In_617);
nand U200 (N_200,In_296,In_205);
nand U201 (N_201,In_1112,In_226);
nand U202 (N_202,In_1404,In_862);
nand U203 (N_203,In_1167,In_277);
or U204 (N_204,In_1123,In_1120);
and U205 (N_205,In_308,In_803);
nand U206 (N_206,In_516,In_715);
or U207 (N_207,In_1142,In_60);
nor U208 (N_208,In_175,In_1373);
and U209 (N_209,In_602,In_611);
nand U210 (N_210,In_477,In_533);
xnor U211 (N_211,In_392,In_1411);
and U212 (N_212,In_155,In_378);
nor U213 (N_213,In_767,In_1035);
or U214 (N_214,In_773,In_912);
nand U215 (N_215,In_1236,In_1202);
or U216 (N_216,In_964,In_807);
and U217 (N_217,In_152,In_1402);
nor U218 (N_218,In_1296,In_897);
or U219 (N_219,In_1383,In_542);
and U220 (N_220,In_1379,In_852);
and U221 (N_221,In_1070,In_1409);
nor U222 (N_222,In_17,In_1117);
or U223 (N_223,In_629,In_1465);
xor U224 (N_224,In_358,In_1390);
nand U225 (N_225,In_1188,In_599);
or U226 (N_226,In_1345,In_255);
and U227 (N_227,In_230,In_1002);
or U228 (N_228,In_782,In_1319);
nand U229 (N_229,In_70,In_204);
nor U230 (N_230,In_892,In_1151);
nor U231 (N_231,In_1086,In_138);
or U232 (N_232,In_491,In_842);
or U233 (N_233,In_849,In_71);
or U234 (N_234,In_1130,In_1312);
and U235 (N_235,In_66,In_80);
nor U236 (N_236,In_661,In_708);
and U237 (N_237,In_390,In_1232);
or U238 (N_238,In_207,In_891);
xor U239 (N_239,In_1072,In_1040);
nor U240 (N_240,In_251,In_1241);
nor U241 (N_241,In_1100,In_375);
or U242 (N_242,In_29,In_620);
and U243 (N_243,In_703,In_1000);
and U244 (N_244,In_1476,In_1432);
or U245 (N_245,In_1254,In_1125);
nor U246 (N_246,In_304,In_1221);
or U247 (N_247,In_522,In_783);
nor U248 (N_248,In_796,In_146);
nand U249 (N_249,In_62,In_562);
and U250 (N_250,In_908,In_556);
nor U251 (N_251,In_523,In_1330);
xor U252 (N_252,In_124,In_76);
or U253 (N_253,N_54,In_1293);
or U254 (N_254,In_397,In_345);
or U255 (N_255,In_1150,In_971);
nand U256 (N_256,In_1198,In_436);
nand U257 (N_257,In_856,N_23);
nand U258 (N_258,In_472,In_1212);
or U259 (N_259,In_437,In_956);
nor U260 (N_260,N_36,In_1006);
nor U261 (N_261,In_403,In_1307);
or U262 (N_262,In_307,In_443);
or U263 (N_263,In_123,In_667);
nor U264 (N_264,In_465,N_182);
nor U265 (N_265,In_4,In_420);
or U266 (N_266,In_957,In_924);
or U267 (N_267,In_37,In_1206);
or U268 (N_268,In_417,In_1168);
nand U269 (N_269,In_1026,In_1);
nor U270 (N_270,In_960,N_166);
nor U271 (N_271,In_1051,In_929);
or U272 (N_272,In_188,In_1397);
or U273 (N_273,In_266,In_200);
nand U274 (N_274,In_133,In_520);
and U275 (N_275,In_1133,In_132);
nand U276 (N_276,In_1204,In_1408);
or U277 (N_277,In_585,In_922);
nor U278 (N_278,In_633,In_1365);
nand U279 (N_279,In_228,In_1308);
nor U280 (N_280,N_160,In_1325);
nor U281 (N_281,In_1437,In_147);
or U282 (N_282,N_41,In_791);
nor U283 (N_283,In_253,In_1152);
nand U284 (N_284,N_219,In_755);
and U285 (N_285,In_1318,In_1111);
nor U286 (N_286,In_569,N_65);
or U287 (N_287,In_557,In_300);
xnor U288 (N_288,N_45,In_770);
and U289 (N_289,In_724,In_449);
or U290 (N_290,In_1174,N_105);
or U291 (N_291,In_651,In_365);
xor U292 (N_292,N_55,In_69);
xor U293 (N_293,In_469,In_235);
and U294 (N_294,In_1108,In_878);
nor U295 (N_295,N_172,In_1007);
nor U296 (N_296,N_79,In_830);
nor U297 (N_297,In_595,In_810);
nand U298 (N_298,In_1191,In_894);
nand U299 (N_299,In_1094,In_941);
or U300 (N_300,In_1281,In_135);
and U301 (N_301,In_1396,In_1237);
nor U302 (N_302,In_931,In_829);
and U303 (N_303,In_276,N_49);
nand U304 (N_304,In_1446,In_890);
or U305 (N_305,In_1417,N_210);
nand U306 (N_306,In_551,N_44);
or U307 (N_307,In_187,In_744);
nor U308 (N_308,In_165,In_932);
nand U309 (N_309,In_275,N_66);
nand U310 (N_310,In_504,In_1075);
or U311 (N_311,In_195,In_541);
nor U312 (N_312,N_16,N_78);
and U313 (N_313,In_1129,In_764);
xnor U314 (N_314,In_691,In_233);
and U315 (N_315,In_666,In_261);
nand U316 (N_316,In_278,In_1275);
nand U317 (N_317,In_911,In_426);
and U318 (N_318,In_1300,In_238);
or U319 (N_319,In_56,N_25);
and U320 (N_320,N_188,In_292);
or U321 (N_321,In_712,In_728);
and U322 (N_322,N_42,In_825);
and U323 (N_323,In_1459,In_743);
xor U324 (N_324,N_163,N_33);
nor U325 (N_325,N_142,In_1445);
nor U326 (N_326,N_175,In_1246);
and U327 (N_327,In_1273,N_7);
nor U328 (N_328,In_792,N_52);
nor U329 (N_329,N_27,In_1231);
and U330 (N_330,In_1441,In_26);
nand U331 (N_331,In_1144,N_71);
and U332 (N_332,In_754,In_273);
nand U333 (N_333,In_218,In_227);
xnor U334 (N_334,In_1362,In_170);
or U335 (N_335,In_1189,N_88);
nor U336 (N_336,In_760,N_164);
and U337 (N_337,In_683,In_855);
nand U338 (N_338,N_205,In_444);
nand U339 (N_339,In_880,In_1039);
and U340 (N_340,In_1017,In_1412);
nor U341 (N_341,In_1037,N_97);
nor U342 (N_342,In_1024,N_204);
nor U343 (N_343,In_934,In_330);
nand U344 (N_344,In_90,In_1385);
nand U345 (N_345,In_474,In_1203);
or U346 (N_346,In_1290,N_68);
nand U347 (N_347,In_1138,N_83);
nor U348 (N_348,N_48,In_1245);
and U349 (N_349,In_801,In_1048);
or U350 (N_350,In_609,N_109);
nor U351 (N_351,In_877,In_1009);
nand U352 (N_352,In_1054,In_1015);
nand U353 (N_353,N_184,N_46);
or U354 (N_354,In_1259,In_36);
xnor U355 (N_355,N_237,In_1251);
nand U356 (N_356,In_1292,In_505);
nand U357 (N_357,In_898,In_267);
or U358 (N_358,In_537,In_434);
and U359 (N_359,N_183,In_1449);
and U360 (N_360,In_1343,N_148);
nor U361 (N_361,N_144,In_980);
or U362 (N_362,In_1279,N_108);
nand U363 (N_363,In_674,In_15);
xnor U364 (N_364,In_828,N_195);
nand U365 (N_365,N_70,In_1064);
nor U366 (N_366,In_1479,N_216);
nand U367 (N_367,In_1426,In_1196);
or U368 (N_368,In_1065,In_1013);
and U369 (N_369,In_65,In_1436);
or U370 (N_370,N_8,In_938);
nand U371 (N_371,N_117,In_1096);
or U372 (N_372,In_172,In_1215);
nand U373 (N_373,In_579,In_1456);
xnor U374 (N_374,In_716,In_638);
and U375 (N_375,In_1276,In_711);
or U376 (N_376,In_9,N_203);
nand U377 (N_377,In_347,N_98);
and U378 (N_378,In_561,In_206);
or U379 (N_379,N_74,In_475);
xor U380 (N_380,N_107,In_57);
nand U381 (N_381,In_989,In_1173);
nor U382 (N_382,N_229,In_54);
and U383 (N_383,N_80,In_92);
nand U384 (N_384,In_425,In_509);
or U385 (N_385,N_30,In_494);
xnor U386 (N_386,N_22,In_613);
and U387 (N_387,In_264,In_572);
nor U388 (N_388,In_360,N_171);
and U389 (N_389,N_181,In_1076);
nand U390 (N_390,In_789,N_103);
or U391 (N_391,In_274,N_90);
or U392 (N_392,In_131,In_1004);
nor U393 (N_393,In_88,In_497);
or U394 (N_394,In_1414,N_151);
and U395 (N_395,In_895,N_146);
nand U396 (N_396,In_1271,In_625);
nand U397 (N_397,In_1313,N_165);
and U398 (N_398,In_410,In_970);
and U399 (N_399,In_699,In_1357);
or U400 (N_400,N_227,In_1068);
or U401 (N_401,N_21,In_1473);
and U402 (N_402,In_978,In_725);
nand U403 (N_403,In_454,N_153);
nand U404 (N_404,In_1220,N_10);
or U405 (N_405,In_887,N_11);
and U406 (N_406,In_1088,In_129);
nand U407 (N_407,In_12,In_413);
xor U408 (N_408,In_840,In_457);
or U409 (N_409,In_1480,In_1027);
nor U410 (N_410,In_1099,In_1466);
nor U411 (N_411,In_1386,In_762);
or U412 (N_412,In_1458,N_194);
xnor U413 (N_413,In_1484,N_245);
and U414 (N_414,In_331,In_406);
and U415 (N_415,In_944,In_5);
xor U416 (N_416,In_813,In_1453);
or U417 (N_417,In_463,In_1294);
or U418 (N_418,In_377,N_162);
or U419 (N_419,In_38,In_959);
nand U420 (N_420,N_116,In_920);
or U421 (N_421,In_256,In_50);
and U422 (N_422,N_87,In_656);
nand U423 (N_423,In_1055,In_1316);
and U424 (N_424,N_24,In_865);
xor U425 (N_425,In_748,In_679);
nand U426 (N_426,In_734,In_327);
or U427 (N_427,In_27,N_155);
nor U428 (N_428,N_191,In_109);
nor U429 (N_429,In_106,In_800);
xor U430 (N_430,In_833,In_67);
nand U431 (N_431,In_318,In_583);
and U432 (N_432,In_1368,In_348);
or U433 (N_433,In_919,In_485);
xor U434 (N_434,In_137,N_99);
nand U435 (N_435,In_130,In_564);
and U436 (N_436,In_1105,In_976);
or U437 (N_437,In_423,In_391);
xnor U438 (N_438,In_808,In_223);
or U439 (N_439,In_689,In_972);
or U440 (N_440,In_873,In_482);
nor U441 (N_441,In_763,N_125);
nor U442 (N_442,In_79,N_234);
or U443 (N_443,In_416,N_129);
nand U444 (N_444,In_860,In_148);
nand U445 (N_445,In_51,In_1083);
nor U446 (N_446,In_876,In_370);
nand U447 (N_447,In_336,N_138);
or U448 (N_448,In_328,In_1183);
or U449 (N_449,In_35,In_795);
and U450 (N_450,In_1447,In_119);
and U451 (N_451,N_134,N_197);
nand U452 (N_452,N_147,In_1057);
nand U453 (N_453,In_584,In_451);
nand U454 (N_454,In_1205,In_418);
and U455 (N_455,In_419,In_589);
nand U456 (N_456,In_30,In_496);
and U457 (N_457,In_279,N_231);
and U458 (N_458,In_652,In_298);
nand U459 (N_459,In_1367,In_22);
or U460 (N_460,In_371,N_5);
or U461 (N_461,In_727,In_937);
or U462 (N_462,In_495,In_197);
and U463 (N_463,In_144,In_776);
or U464 (N_464,In_577,In_785);
or U465 (N_465,N_212,N_111);
and U466 (N_466,In_74,In_156);
nand U467 (N_467,N_156,In_19);
or U468 (N_468,In_1299,N_150);
or U469 (N_469,N_15,In_178);
and U470 (N_470,In_158,In_756);
nor U471 (N_471,In_640,N_113);
nor U472 (N_472,N_149,In_357);
xnor U473 (N_473,In_389,In_622);
and U474 (N_474,In_281,In_612);
nand U475 (N_475,N_127,In_565);
and U476 (N_476,In_1433,In_590);
nand U477 (N_477,In_925,In_376);
nor U478 (N_478,In_96,In_411);
xnor U479 (N_479,In_545,In_886);
and U480 (N_480,In_1471,In_382);
or U481 (N_481,In_1428,In_1431);
xor U482 (N_482,N_235,In_619);
nand U483 (N_483,In_1361,In_818);
and U484 (N_484,In_1060,In_693);
nand U485 (N_485,In_751,In_1495);
or U486 (N_486,In_717,In_182);
nand U487 (N_487,In_128,In_294);
nand U488 (N_488,In_1171,In_98);
or U489 (N_489,N_200,In_1084);
nand U490 (N_490,In_974,N_115);
xnor U491 (N_491,In_798,In_948);
or U492 (N_492,In_1391,In_447);
xnor U493 (N_493,In_120,In_1244);
nand U494 (N_494,N_50,In_535);
and U495 (N_495,In_645,N_139);
or U496 (N_496,In_269,In_47);
and U497 (N_497,In_1107,In_1008);
xnor U498 (N_498,N_0,In_196);
nand U499 (N_499,In_581,In_271);
nor U500 (N_500,N_121,N_95);
nor U501 (N_501,N_384,N_288);
xor U502 (N_502,In_141,N_60);
xnor U503 (N_503,N_269,N_380);
or U504 (N_504,In_1419,N_441);
nand U505 (N_505,In_1209,N_220);
nand U506 (N_506,In_1126,In_111);
or U507 (N_507,N_370,In_884);
and U508 (N_508,In_1145,N_301);
nor U509 (N_509,In_87,In_1135);
and U510 (N_510,N_345,In_272);
nor U511 (N_511,N_201,N_81);
xor U512 (N_512,N_333,N_17);
or U513 (N_513,In_33,In_1175);
xnor U514 (N_514,In_648,In_213);
or U515 (N_515,In_847,N_438);
or U516 (N_516,In_478,N_140);
nand U517 (N_517,In_597,In_479);
and U518 (N_518,N_402,N_187);
and U519 (N_519,N_314,In_1208);
nand U520 (N_520,In_675,In_731);
and U521 (N_521,In_387,N_316);
nor U522 (N_522,N_85,In_692);
and U523 (N_523,In_459,In_826);
or U524 (N_524,In_962,N_86);
and U525 (N_525,N_317,N_102);
nor U526 (N_526,In_58,N_76);
or U527 (N_527,N_465,N_418);
and U528 (N_528,N_386,N_429);
nor U529 (N_529,In_324,N_124);
or U530 (N_530,N_471,N_255);
nor U531 (N_531,In_18,In_192);
and U532 (N_532,In_380,N_295);
nand U533 (N_533,N_328,N_456);
xor U534 (N_534,N_393,In_1038);
and U535 (N_535,N_332,N_446);
nor U536 (N_536,In_1369,In_319);
nor U537 (N_537,N_62,In_1109);
or U538 (N_538,In_567,N_217);
xor U539 (N_539,In_824,N_266);
nor U540 (N_540,N_338,In_306);
or U541 (N_541,In_470,In_738);
xnor U542 (N_542,In_1272,In_714);
nand U543 (N_543,N_489,In_512);
and U544 (N_544,N_59,In_1046);
nand U545 (N_545,In_555,In_1477);
or U546 (N_546,In_1082,N_308);
nor U547 (N_547,N_413,In_525);
or U548 (N_548,N_267,In_1461);
nor U549 (N_549,N_126,In_901);
or U550 (N_550,In_297,In_379);
and U551 (N_551,N_92,In_608);
and U552 (N_552,In_245,In_104);
nand U553 (N_553,N_335,In_1067);
nor U554 (N_554,N_450,N_303);
nor U555 (N_555,N_89,N_239);
nor U556 (N_556,In_740,N_334);
and U557 (N_557,In_481,N_327);
nor U558 (N_558,N_364,In_642);
nor U559 (N_559,In_993,In_593);
and U560 (N_560,In_707,N_331);
and U561 (N_561,N_279,N_104);
nand U562 (N_562,In_746,In_1329);
or U563 (N_563,In_529,In_52);
or U564 (N_564,In_461,In_341);
or U565 (N_565,N_35,N_118);
and U566 (N_566,N_388,In_988);
xor U567 (N_567,In_493,In_1405);
xor U568 (N_568,In_220,In_202);
and U569 (N_569,N_120,In_896);
and U570 (N_570,In_1363,In_259);
nor U571 (N_571,N_100,N_356);
and U572 (N_572,N_241,N_312);
nand U573 (N_573,N_484,In_201);
nand U574 (N_574,In_110,N_344);
and U575 (N_575,In_802,In_519);
and U576 (N_576,N_223,In_351);
or U577 (N_577,N_270,In_558);
nand U578 (N_578,In_367,N_401);
or U579 (N_579,In_166,In_161);
nand U580 (N_580,In_1148,In_1091);
nor U581 (N_581,In_1258,N_466);
nor U582 (N_582,In_1474,In_1217);
and U583 (N_583,N_12,N_361);
or U584 (N_584,N_490,In_1486);
nor U585 (N_585,N_474,In_1421);
nand U586 (N_586,N_369,In_1399);
nand U587 (N_587,In_566,N_381);
or U588 (N_588,N_34,N_271);
or U589 (N_589,N_274,In_452);
nor U590 (N_590,In_136,In_1087);
nand U591 (N_591,In_488,N_460);
nor U592 (N_592,N_143,In_1499);
or U593 (N_593,In_409,In_969);
nor U594 (N_594,In_433,In_907);
or U595 (N_595,N_13,In_1354);
nand U596 (N_596,In_1020,N_64);
nor U597 (N_597,N_298,In_871);
xnor U598 (N_598,In_961,N_193);
nand U599 (N_599,In_31,N_315);
nand U600 (N_600,In_393,N_63);
nand U601 (N_601,N_321,In_1115);
or U602 (N_602,N_20,In_289);
nand U603 (N_603,In_844,N_273);
nand U604 (N_604,In_349,In_455);
nand U605 (N_605,In_1147,In_270);
nand U606 (N_606,In_1023,N_259);
nand U607 (N_607,N_367,In_115);
nand U608 (N_608,N_340,In_603);
nor U609 (N_609,In_994,In_544);
nor U610 (N_610,In_3,In_55);
nor U611 (N_611,N_481,In_1387);
and U612 (N_612,N_1,In_521);
nand U613 (N_613,In_726,N_427);
and U614 (N_614,N_351,In_888);
and U615 (N_615,In_325,N_268);
or U616 (N_616,N_224,In_1326);
or U617 (N_617,In_761,In_1178);
nor U618 (N_618,N_487,In_943);
nand U619 (N_619,In_501,N_174);
nand U620 (N_620,N_199,N_93);
xor U621 (N_621,N_320,In_511);
and U622 (N_622,N_323,N_448);
nand U623 (N_623,In_249,In_582);
xor U624 (N_624,N_464,In_385);
nor U625 (N_625,N_215,N_178);
nand U626 (N_626,N_96,In_428);
nor U627 (N_627,In_1018,N_496);
xor U628 (N_628,N_82,In_225);
and U629 (N_629,In_323,In_282);
nor U630 (N_630,N_348,In_1306);
and U631 (N_631,In_845,In_362);
nand U632 (N_632,In_1062,N_31);
nor U633 (N_633,In_1451,N_264);
or U634 (N_634,In_1394,N_75);
and U635 (N_635,In_1121,In_384);
and U636 (N_636,N_373,In_563);
nor U637 (N_637,In_1180,In_1012);
nand U638 (N_638,N_73,N_284);
nand U639 (N_639,In_1098,In_1016);
and U640 (N_640,In_592,N_412);
nand U641 (N_641,In_1256,N_176);
nor U642 (N_642,In_315,In_682);
nand U643 (N_643,In_1140,N_475);
or U644 (N_644,In_1470,In_299);
and U645 (N_645,In_353,In_312);
and U646 (N_646,In_784,In_1469);
and U647 (N_647,N_265,In_81);
or U648 (N_648,N_252,In_1185);
xor U649 (N_649,In_1089,In_1176);
and U650 (N_650,N_425,N_453);
nor U651 (N_651,In_536,N_179);
nor U652 (N_652,In_637,N_389);
xnor U653 (N_653,N_387,N_84);
nand U654 (N_654,In_441,N_294);
and U655 (N_655,In_1377,N_233);
nor U656 (N_656,In_528,In_492);
nand U657 (N_657,In_806,In_722);
nor U658 (N_658,In_314,In_1028);
nand U659 (N_659,In_635,In_1252);
or U660 (N_660,In_663,N_420);
xor U661 (N_661,N_479,N_488);
and U662 (N_662,In_1025,In_779);
nand U663 (N_663,N_275,In_547);
and U664 (N_664,In_1286,In_257);
nand U665 (N_665,In_1478,In_900);
and U666 (N_666,N_206,In_552);
or U667 (N_667,In_1475,N_325);
nand U668 (N_668,In_678,N_372);
and U669 (N_669,N_18,N_359);
nor U670 (N_670,In_1164,In_736);
nand U671 (N_671,In_85,In_1488);
or U672 (N_672,In_258,In_632);
nor U673 (N_673,N_157,In_450);
or U674 (N_674,N_404,In_1253);
nand U675 (N_675,In_1162,In_412);
nor U676 (N_676,In_1118,In_333);
nor U677 (N_677,In_1134,In_672);
nor U678 (N_678,N_434,In_1311);
and U679 (N_679,N_394,In_1262);
or U680 (N_680,N_411,In_95);
or U681 (N_681,In_605,In_303);
or U682 (N_682,In_372,N_180);
nand U683 (N_683,In_1034,In_466);
xnor U684 (N_684,In_1344,In_686);
nand U685 (N_685,In_850,N_408);
or U686 (N_686,N_222,In_1019);
nor U687 (N_687,In_184,In_1491);
xnor U688 (N_688,In_288,In_1101);
nand U689 (N_689,In_1169,N_136);
nor U690 (N_690,In_863,In_1283);
nand U691 (N_691,N_106,In_193);
nand U692 (N_692,In_1031,N_132);
xnor U693 (N_693,N_468,In_39);
or U694 (N_694,In_11,N_141);
or U695 (N_695,In_139,In_1392);
nand U696 (N_696,In_1192,In_749);
and U697 (N_697,In_1346,N_458);
and U698 (N_698,N_167,N_198);
nor U699 (N_699,N_58,N_170);
nand U700 (N_700,In_183,In_861);
and U701 (N_701,N_414,In_1496);
or U702 (N_702,In_641,N_349);
or U703 (N_703,N_486,N_431);
and U704 (N_704,In_432,N_305);
nand U705 (N_705,In_1149,In_1041);
nand U706 (N_706,In_404,In_665);
nor U707 (N_707,In_399,In_53);
nor U708 (N_708,N_405,N_360);
nor U709 (N_709,In_1356,N_3);
nor U710 (N_710,In_942,In_804);
nand U711 (N_711,N_190,In_644);
or U712 (N_712,N_213,N_318);
nand U713 (N_713,In_601,N_218);
nor U714 (N_714,In_772,N_276);
nand U715 (N_715,N_72,In_1282);
nand U716 (N_716,In_1103,In_591);
nor U717 (N_717,In_334,In_373);
xor U718 (N_718,In_1443,N_110);
or U719 (N_719,In_954,N_395);
and U720 (N_720,In_983,N_322);
or U721 (N_721,In_647,In_757);
xnor U722 (N_722,In_1061,In_1197);
nand U723 (N_723,In_116,In_1321);
and U724 (N_724,N_355,In_1124);
nand U725 (N_725,In_543,N_463);
nand U726 (N_726,N_306,In_540);
nor U727 (N_727,N_406,In_834);
nand U728 (N_728,In_342,N_29);
and U729 (N_729,In_1097,N_366);
or U730 (N_730,In_1182,N_480);
or U731 (N_731,N_2,In_1010);
or U732 (N_732,In_208,In_1153);
nand U733 (N_733,In_705,In_263);
xor U734 (N_734,In_982,In_1304);
and U735 (N_735,In_1309,In_309);
and U736 (N_736,N_311,N_272);
xnor U737 (N_737,N_302,In_1314);
or U738 (N_738,In_1250,N_499);
nand U739 (N_739,In_1261,N_391);
or U740 (N_740,In_1485,In_7);
nor U741 (N_741,N_447,N_119);
and U742 (N_742,N_422,In_1187);
or U743 (N_743,N_374,N_177);
or U744 (N_744,N_262,In_1201);
or U745 (N_745,N_77,In_203);
and U746 (N_746,In_1157,N_4);
or U747 (N_747,In_1260,In_1059);
nand U748 (N_748,In_1155,In_630);
xor U749 (N_749,N_358,In_93);
or U750 (N_750,N_592,In_631);
nor U751 (N_751,In_568,In_1214);
or U752 (N_752,N_561,In_1372);
and U753 (N_753,In_1228,N_697);
and U754 (N_754,N_432,N_527);
xnor U755 (N_755,In_1341,In_998);
or U756 (N_756,N_663,N_504);
nand U757 (N_757,In_1490,In_364);
nor U758 (N_758,N_291,N_399);
xor U759 (N_759,In_487,In_402);
nand U760 (N_760,N_604,N_628);
nand U761 (N_761,In_777,N_688);
nor U762 (N_762,N_297,N_469);
or U763 (N_763,N_657,In_429);
nand U764 (N_764,N_722,N_661);
nand U765 (N_765,N_507,N_495);
nand U766 (N_766,In_483,In_1210);
xnor U767 (N_767,N_741,N_249);
and U768 (N_768,N_512,In_181);
or U769 (N_769,N_717,In_231);
nand U770 (N_770,In_553,In_864);
or U771 (N_771,In_490,N_354);
nand U772 (N_772,In_914,In_967);
or U773 (N_773,N_591,In_1450);
nand U774 (N_774,N_703,In_143);
xnor U775 (N_775,N_670,In_759);
or U776 (N_776,N_283,N_528);
or U777 (N_777,In_1440,N_440);
xor U778 (N_778,N_6,In_821);
nand U779 (N_779,N_551,In_870);
nor U780 (N_780,N_701,In_1497);
nand U781 (N_781,N_559,N_290);
xor U782 (N_782,In_574,N_173);
xor U783 (N_783,In_1223,N_698);
and U784 (N_784,In_77,N_720);
and U785 (N_785,N_589,In_1492);
and U786 (N_786,In_750,In_1247);
nor U787 (N_787,In_643,N_627);
nor U788 (N_788,In_841,In_1156);
nand U789 (N_789,In_1200,N_545);
nand U790 (N_790,N_564,In_1184);
and U791 (N_791,N_652,N_641);
nand U792 (N_792,N_673,N_400);
nor U793 (N_793,N_565,N_671);
and U794 (N_794,In_191,In_317);
nand U795 (N_795,N_577,In_1454);
or U796 (N_796,N_472,In_1301);
xor U797 (N_797,In_513,N_228);
and U798 (N_798,In_659,In_61);
xnor U799 (N_799,In_59,In_1305);
nand U800 (N_800,In_883,In_73);
and U801 (N_801,N_533,In_1413);
nand U802 (N_802,In_335,In_548);
nand U803 (N_803,N_686,N_694);
or U804 (N_804,In_1339,In_1366);
and U805 (N_805,N_513,N_609);
nand U806 (N_806,In_739,N_56);
nand U807 (N_807,In_742,N_397);
or U808 (N_808,In_786,N_729);
or U809 (N_809,N_28,N_730);
nor U810 (N_810,N_256,N_597);
xnor U811 (N_811,N_368,N_749);
nand U812 (N_812,N_517,N_159);
nor U813 (N_813,N_467,N_588);
nand U814 (N_814,N_497,N_436);
and U815 (N_815,In_1093,In_606);
nor U816 (N_816,In_706,N_626);
nor U817 (N_817,N_616,N_506);
or U818 (N_818,In_975,In_906);
and U819 (N_819,In_1340,In_210);
and U820 (N_820,In_1434,N_539);
nand U821 (N_821,In_1427,In_176);
and U822 (N_822,In_1102,In_1442);
or U823 (N_823,N_500,N_693);
nand U824 (N_824,N_32,In_741);
xnor U825 (N_825,In_140,In_1455);
nor U826 (N_826,N_649,N_313);
nor U827 (N_827,In_46,N_674);
nor U828 (N_828,In_1077,In_126);
and U829 (N_829,In_923,N_114);
nor U830 (N_830,N_529,N_696);
xor U831 (N_831,N_683,N_581);
and U832 (N_832,N_740,N_721);
nor U833 (N_833,N_637,N_624);
nor U834 (N_834,In_814,In_381);
or U835 (N_835,N_130,In_1328);
or U836 (N_836,N_664,In_697);
nand U837 (N_837,N_731,N_417);
or U838 (N_838,N_576,N_678);
nand U839 (N_839,In_1317,In_684);
nor U840 (N_840,N_599,N_398);
nor U841 (N_841,N_346,N_336);
xnor U842 (N_842,N_716,N_424);
and U843 (N_843,N_656,In_913);
nand U844 (N_844,N_737,N_392);
or U845 (N_845,N_154,N_736);
nor U846 (N_846,N_482,In_1114);
or U847 (N_847,N_746,N_342);
xor U848 (N_848,N_553,N_337);
or U849 (N_849,N_611,In_1239);
or U850 (N_850,In_769,N_725);
or U851 (N_851,In_1439,N_14);
xor U852 (N_852,N_378,N_37);
nor U853 (N_853,N_462,In_1063);
and U854 (N_854,N_537,N_726);
or U855 (N_855,In_1003,N_169);
nand U856 (N_856,N_633,N_362);
nor U857 (N_857,N_685,N_590);
and U858 (N_858,N_610,N_459);
nor U859 (N_859,N_550,In_1400);
nand U860 (N_860,N_202,In_435);
and U861 (N_861,N_257,N_133);
nor U862 (N_862,In_977,In_1320);
and U863 (N_863,In_854,N_690);
nor U864 (N_864,N_379,N_211);
nor U865 (N_865,In_1080,N_442);
nand U866 (N_866,N_713,N_575);
nor U867 (N_867,In_965,N_518);
nand U868 (N_868,N_363,N_629);
nor U869 (N_869,N_509,In_953);
nand U870 (N_870,N_145,N_692);
and U871 (N_871,N_710,In_669);
or U872 (N_872,In_359,N_744);
and U873 (N_873,N_745,In_794);
nand U874 (N_874,In_1464,In_1460);
or U875 (N_875,N_236,In_1085);
nand U876 (N_876,In_872,In_339);
or U877 (N_877,N_415,N_455);
nor U878 (N_878,In_1146,In_765);
and U879 (N_879,N_723,N_625);
nand U880 (N_880,N_280,N_541);
nor U881 (N_881,N_530,N_523);
nor U882 (N_882,N_734,In_832);
nand U883 (N_883,N_546,N_571);
nor U884 (N_884,N_665,N_324);
or U885 (N_885,N_407,N_714);
nand U886 (N_886,In_1467,N_522);
xnor U887 (N_887,N_232,N_570);
xnor U888 (N_888,N_43,N_650);
nor U889 (N_889,In_320,N_587);
nand U890 (N_890,N_708,In_1398);
xnor U891 (N_891,In_438,In_401);
or U892 (N_892,N_260,N_491);
or U893 (N_893,N_137,In_650);
xor U894 (N_894,N_385,N_501);
or U895 (N_895,N_739,N_573);
nand U896 (N_896,N_350,In_68);
or U897 (N_897,In_517,N_377);
nor U898 (N_898,N_214,N_630);
or U899 (N_899,In_1195,N_292);
or U900 (N_900,N_326,N_615);
xnor U901 (N_901,In_1179,In_1071);
and U902 (N_902,N_544,In_507);
nor U903 (N_903,N_572,In_396);
and U904 (N_904,N_67,In_951);
or U905 (N_905,In_1116,In_680);
or U906 (N_906,In_885,In_214);
or U907 (N_907,In_430,N_357);
nand U908 (N_908,In_242,In_121);
nor U909 (N_909,N_525,In_1143);
and U910 (N_910,In_316,N_423);
nor U911 (N_911,N_602,N_555);
nand U912 (N_912,In_882,N_365);
and U913 (N_913,In_366,In_1315);
or U914 (N_914,In_14,In_664);
or U915 (N_915,N_226,In_1483);
nor U916 (N_916,In_190,N_648);
xnor U917 (N_917,In_346,In_246);
or U918 (N_918,In_486,N_607);
and U919 (N_919,N_569,In_999);
or U920 (N_920,N_261,N_208);
and U921 (N_921,N_632,In_508);
and U922 (N_922,In_1243,N_38);
nor U923 (N_923,N_242,N_672);
nand U924 (N_924,N_667,In_1226);
nor U925 (N_925,In_13,N_691);
nor U926 (N_926,In_1270,In_1295);
nand U927 (N_927,N_562,N_421);
nand U928 (N_928,N_700,In_610);
or U929 (N_929,In_616,N_281);
or U930 (N_930,In_1095,In_112);
and U931 (N_931,N_521,N_563);
nand U932 (N_932,In_1338,N_352);
or U933 (N_933,N_396,In_105);
and U934 (N_934,N_742,In_720);
xnor U935 (N_935,N_556,In_101);
or U936 (N_936,In_1429,N_383);
or U937 (N_937,N_339,In_1410);
nor U938 (N_938,N_614,In_446);
and U939 (N_939,N_514,N_477);
or U940 (N_940,N_454,N_549);
nand U941 (N_941,N_601,N_285);
or U942 (N_942,N_376,In_1255);
or U943 (N_943,In_990,N_595);
nor U944 (N_944,N_707,N_687);
and U945 (N_945,In_1159,N_743);
nor U946 (N_946,In_514,N_654);
nor U947 (N_947,N_185,N_186);
and U948 (N_948,In_1264,In_32);
or U949 (N_949,In_224,N_619);
nor U950 (N_950,N_738,In_991);
or U951 (N_951,N_547,N_286);
and U952 (N_952,In_639,N_263);
nor U953 (N_953,In_1170,In_875);
nor U954 (N_954,N_461,N_457);
or U955 (N_955,In_846,In_719);
or U956 (N_956,In_1177,In_745);
xnor U957 (N_957,In_1081,In_1056);
xor U958 (N_958,In_355,N_9);
nor U959 (N_959,N_519,N_594);
or U960 (N_960,In_532,N_244);
nor U961 (N_961,N_330,In_928);
and U962 (N_962,In_1336,N_445);
nand U963 (N_963,In_1128,N_483);
and U964 (N_964,In_917,N_341);
or U965 (N_965,In_211,N_307);
nand U966 (N_966,N_711,In_1119);
and U967 (N_967,In_1005,N_300);
or U968 (N_968,N_733,In_527);
or U969 (N_969,In_1163,N_304);
or U970 (N_970,In_285,N_532);
nor U971 (N_971,N_596,In_1435);
and U972 (N_972,N_593,N_583);
xor U973 (N_973,N_508,N_51);
xnor U974 (N_974,N_449,In_471);
and U975 (N_975,In_209,In_1047);
nor U976 (N_976,N_554,In_945);
nor U977 (N_977,In_904,N_681);
nor U978 (N_978,N_524,In_1224);
or U979 (N_979,In_1042,In_1277);
nor U980 (N_980,In_752,N_196);
nand U981 (N_981,N_47,In_733);
and U982 (N_982,N_503,N_439);
nand U983 (N_983,N_498,In_321);
nor U984 (N_984,In_0,N_123);
or U985 (N_985,N_510,N_293);
nor U986 (N_986,In_114,In_484);
nor U987 (N_987,N_579,In_1218);
nor U988 (N_988,N_666,N_643);
nand U989 (N_989,N_329,N_419);
nand U990 (N_990,N_732,In_134);
nor U991 (N_991,N_437,In_573);
xnor U992 (N_992,In_538,N_580);
xor U993 (N_993,In_822,In_222);
nor U994 (N_994,In_212,N_409);
nor U995 (N_995,N_152,In_1263);
or U996 (N_996,N_682,N_516);
nor U997 (N_997,N_675,N_705);
and U998 (N_998,In_1498,N_646);
or U999 (N_999,In_627,N_189);
or U1000 (N_1000,In_987,N_299);
or U1001 (N_1001,N_968,In_1161);
and U1002 (N_1002,In_460,In_48);
and U1003 (N_1003,N_820,In_1462);
and U1004 (N_1004,N_854,In_21);
or U1005 (N_1005,N_724,N_786);
and U1006 (N_1006,N_862,N_403);
nand U1007 (N_1007,N_988,N_526);
nor U1008 (N_1008,N_578,N_895);
and U1009 (N_1009,N_603,N_112);
nor U1010 (N_1010,N_251,N_128);
or U1011 (N_1011,In_838,N_855);
or U1012 (N_1012,N_882,N_828);
nor U1013 (N_1013,In_662,N_924);
nand U1014 (N_1014,In_1348,N_531);
xor U1015 (N_1015,N_435,N_976);
nand U1016 (N_1016,N_574,N_779);
nand U1017 (N_1017,N_826,N_221);
and U1018 (N_1018,N_444,N_872);
and U1019 (N_1019,N_788,N_347);
nor U1020 (N_1020,N_844,N_240);
nor U1021 (N_1021,N_473,N_931);
or U1022 (N_1022,N_927,N_906);
or U1023 (N_1023,N_827,In_125);
and U1024 (N_1024,N_763,In_690);
and U1025 (N_1025,N_877,N_645);
or U1026 (N_1026,N_542,N_890);
and U1027 (N_1027,N_225,N_796);
nor U1028 (N_1028,N_959,N_606);
or U1029 (N_1029,In_83,N_760);
nor U1030 (N_1030,N_131,N_905);
nand U1031 (N_1031,In_1303,In_356);
nand U1032 (N_1032,In_947,N_909);
and U1033 (N_1033,N_792,N_842);
nand U1034 (N_1034,N_880,N_973);
or U1035 (N_1035,N_859,N_998);
and U1036 (N_1036,N_797,N_793);
nand U1037 (N_1037,N_791,N_704);
and U1038 (N_1038,N_861,N_825);
nor U1039 (N_1039,N_543,N_91);
xor U1040 (N_1040,N_642,N_932);
and U1041 (N_1041,N_727,N_248);
and U1042 (N_1042,N_892,N_798);
nand U1043 (N_1043,In_549,In_440);
nor U1044 (N_1044,N_761,N_787);
and U1045 (N_1045,N_289,N_161);
xor U1046 (N_1046,N_718,In_1154);
or U1047 (N_1047,N_598,N_878);
or U1048 (N_1048,N_958,N_969);
nor U1049 (N_1049,N_608,N_916);
nand U1050 (N_1050,N_794,N_94);
or U1051 (N_1051,N_712,N_702);
or U1052 (N_1052,N_122,N_904);
xnor U1053 (N_1053,N_709,N_908);
nor U1054 (N_1054,N_258,N_492);
or U1055 (N_1055,N_869,N_635);
and U1056 (N_1056,N_853,N_639);
or U1057 (N_1057,N_505,In_153);
nand U1058 (N_1058,N_850,N_662);
or U1059 (N_1059,N_963,N_789);
and U1060 (N_1060,N_799,N_804);
and U1061 (N_1061,N_911,N_954);
nand U1062 (N_1062,N_852,N_600);
and U1063 (N_1063,N_951,N_808);
and U1064 (N_1064,N_978,In_781);
or U1065 (N_1065,N_885,N_975);
nor U1066 (N_1066,N_669,N_679);
nand U1067 (N_1067,N_699,N_61);
or U1068 (N_1068,In_950,N_989);
xnor U1069 (N_1069,N_319,In_199);
nand U1070 (N_1070,N_902,In_63);
nor U1071 (N_1071,N_899,N_896);
nor U1072 (N_1072,N_620,N_928);
or U1073 (N_1073,N_668,N_846);
nand U1074 (N_1074,N_640,N_772);
or U1075 (N_1075,In_1418,N_695);
and U1076 (N_1076,In_43,N_751);
or U1077 (N_1077,N_728,N_747);
nand U1078 (N_1078,N_919,N_209);
and U1079 (N_1079,N_69,N_863);
and U1080 (N_1080,N_343,N_990);
nand U1081 (N_1081,N_375,In_506);
nor U1082 (N_1082,In_623,N_821);
or U1083 (N_1083,N_972,In_737);
or U1084 (N_1084,N_898,In_618);
and U1085 (N_1085,N_382,N_631);
xnor U1086 (N_1086,N_900,In_701);
or U1087 (N_1087,N_971,N_762);
or U1088 (N_1088,N_961,N_893);
or U1089 (N_1089,N_764,N_824);
nand U1090 (N_1090,N_586,N_992);
and U1091 (N_1091,N_889,In_1132);
xor U1092 (N_1092,N_478,N_247);
nor U1093 (N_1093,In_688,N_887);
and U1094 (N_1094,N_848,N_950);
xnor U1095 (N_1095,N_884,N_921);
or U1096 (N_1096,N_838,N_910);
and U1097 (N_1097,N_433,N_948);
nand U1098 (N_1098,N_867,N_230);
nand U1099 (N_1099,N_253,In_185);
nand U1100 (N_1100,N_659,N_40);
and U1101 (N_1101,N_955,N_502);
xnor U1102 (N_1102,N_612,N_868);
nor U1103 (N_1103,N_644,In_305);
nand U1104 (N_1104,N_567,N_939);
and U1105 (N_1105,N_735,In_628);
nand U1106 (N_1106,In_1160,N_775);
and U1107 (N_1107,N_582,N_979);
and U1108 (N_1108,N_912,N_829);
nor U1109 (N_1109,In_1106,N_997);
or U1110 (N_1110,N_984,N_936);
nor U1111 (N_1111,N_560,N_934);
or U1112 (N_1112,N_585,N_830);
nand U1113 (N_1113,N_782,N_897);
xnor U1114 (N_1114,N_901,N_676);
and U1115 (N_1115,N_822,N_557);
nand U1116 (N_1116,N_801,N_282);
nor U1117 (N_1117,N_778,N_53);
nand U1118 (N_1118,In_86,In_580);
or U1119 (N_1119,In_831,N_832);
nand U1120 (N_1120,N_774,N_653);
and U1121 (N_1121,N_278,N_858);
nor U1122 (N_1122,N_677,N_839);
nor U1123 (N_1123,N_660,N_296);
and U1124 (N_1124,N_617,In_995);
or U1125 (N_1125,In_778,N_658);
nand U1126 (N_1126,N_991,In_1110);
nand U1127 (N_1127,N_19,N_962);
nor U1128 (N_1128,N_765,N_783);
or U1129 (N_1129,N_849,In_1104);
xor U1130 (N_1130,N_920,N_956);
nor U1131 (N_1131,N_811,In_1430);
nand U1132 (N_1132,N_622,N_277);
nand U1133 (N_1133,In_234,In_771);
nor U1134 (N_1134,N_894,N_903);
or U1135 (N_1135,In_1393,N_953);
or U1136 (N_1136,N_970,N_795);
or U1137 (N_1137,N_800,In_1213);
and U1138 (N_1138,N_207,N_876);
or U1139 (N_1139,N_840,In_1403);
nand U1140 (N_1140,N_999,N_888);
and U1141 (N_1141,In_1014,N_922);
or U1142 (N_1142,N_818,N_485);
xor U1143 (N_1143,N_836,N_470);
or U1144 (N_1144,N_773,In_1207);
nor U1145 (N_1145,N_715,N_535);
and U1146 (N_1146,N_974,N_390);
nand U1147 (N_1147,N_250,In_217);
nor U1148 (N_1148,In_811,N_443);
nor U1149 (N_1149,N_719,N_875);
and U1150 (N_1150,N_881,N_947);
nor U1151 (N_1151,In_1291,In_179);
or U1152 (N_1152,N_638,N_845);
or U1153 (N_1153,N_841,N_879);
nand U1154 (N_1154,N_520,N_371);
nor U1155 (N_1155,N_870,N_952);
nor U1156 (N_1156,N_949,N_945);
xnor U1157 (N_1157,N_39,In_1052);
xor U1158 (N_1158,N_605,N_940);
and U1159 (N_1159,N_918,N_655);
nor U1160 (N_1160,N_917,N_759);
nor U1161 (N_1161,N_771,In_49);
and U1162 (N_1162,N_925,N_552);
nand U1163 (N_1163,N_777,N_192);
and U1164 (N_1164,N_993,N_613);
or U1165 (N_1165,In_909,In_1284);
and U1166 (N_1166,N_101,N_865);
and U1167 (N_1167,In_75,N_494);
and U1168 (N_1168,N_946,N_915);
nor U1169 (N_1169,N_996,N_254);
nand U1170 (N_1170,N_965,In_78);
xor U1171 (N_1171,In_1401,N_944);
or U1172 (N_1172,In_168,N_860);
xor U1173 (N_1173,N_287,In_554);
nand U1174 (N_1174,N_618,N_689);
and U1175 (N_1175,N_835,N_812);
or U1176 (N_1176,N_158,N_977);
nand U1177 (N_1177,N_807,N_769);
and U1178 (N_1178,In_816,N_982);
nand U1179 (N_1179,N_753,N_623);
xor U1180 (N_1180,N_857,N_748);
or U1181 (N_1181,N_802,N_935);
xnor U1182 (N_1182,In_99,N_987);
nand U1183 (N_1183,N_540,N_416);
and U1184 (N_1184,In_694,N_980);
nor U1185 (N_1185,N_883,N_636);
and U1186 (N_1186,N_871,N_785);
nor U1187 (N_1187,N_943,In_718);
nor U1188 (N_1188,In_262,N_452);
nor U1189 (N_1189,N_756,N_534);
xnor U1190 (N_1190,N_823,N_810);
and U1191 (N_1191,In_159,N_983);
or U1192 (N_1192,N_309,In_881);
or U1193 (N_1193,In_677,N_851);
nand U1194 (N_1194,N_752,N_26);
nand U1195 (N_1195,N_476,N_930);
nor U1196 (N_1196,N_914,N_938);
or U1197 (N_1197,In_468,N_837);
nand U1198 (N_1198,N_843,N_428);
nor U1199 (N_1199,N_493,N_757);
and U1200 (N_1200,N_647,N_886);
nor U1201 (N_1201,N_515,N_754);
nor U1202 (N_1202,N_929,In_1359);
or U1203 (N_1203,In_721,N_933);
or U1204 (N_1204,N_706,N_538);
nand U1205 (N_1205,N_937,N_856);
and U1206 (N_1206,N_942,N_926);
nand U1207 (N_1207,N_548,N_750);
and U1208 (N_1208,N_430,N_790);
or U1209 (N_1209,N_168,N_680);
and U1210 (N_1210,N_767,N_986);
nand U1211 (N_1211,N_864,N_994);
nor U1212 (N_1212,In_215,N_833);
nand U1213 (N_1213,In_1380,In_198);
and U1214 (N_1214,N_813,N_353);
or U1215 (N_1215,N_451,N_770);
xor U1216 (N_1216,N_831,N_805);
nand U1217 (N_1217,N_923,N_967);
xor U1218 (N_1218,N_766,N_913);
or U1219 (N_1219,In_753,N_310);
nor U1220 (N_1220,In_163,N_758);
and U1221 (N_1221,In_1353,N_941);
nand U1222 (N_1222,N_243,N_964);
or U1223 (N_1223,N_960,N_781);
or U1224 (N_1224,N_985,N_651);
and U1225 (N_1225,N_684,N_847);
xnor U1226 (N_1226,In_1472,N_957);
nor U1227 (N_1227,In_1199,N_566);
nand U1228 (N_1228,N_806,N_816);
xor U1229 (N_1229,In_45,N_776);
nand U1230 (N_1230,N_891,N_768);
and U1231 (N_1231,N_238,N_834);
and U1232 (N_1232,N_780,N_784);
or U1233 (N_1233,N_246,N_634);
nand U1234 (N_1234,N_817,N_815);
or U1235 (N_1235,N_511,In_247);
nor U1236 (N_1236,N_809,N_621);
or U1237 (N_1237,In_927,In_363);
and U1238 (N_1238,N_907,N_568);
nor U1239 (N_1239,N_410,N_966);
or U1240 (N_1240,N_755,N_866);
nor U1241 (N_1241,In_283,In_361);
nand U1242 (N_1242,N_803,N_981);
nand U1243 (N_1243,In_797,N_814);
xor U1244 (N_1244,N_874,N_873);
nor U1245 (N_1245,N_819,In_414);
and U1246 (N_1246,N_536,N_57);
nand U1247 (N_1247,N_135,N_426);
nand U1248 (N_1248,In_1337,N_995);
and U1249 (N_1249,N_584,N_558);
and U1250 (N_1250,N_1026,N_1109);
nor U1251 (N_1251,N_1065,N_1012);
and U1252 (N_1252,N_1149,N_1217);
and U1253 (N_1253,N_1180,N_1073);
nand U1254 (N_1254,N_1183,N_1014);
nor U1255 (N_1255,N_1061,N_1132);
and U1256 (N_1256,N_1146,N_1164);
nor U1257 (N_1257,N_1140,N_1001);
or U1258 (N_1258,N_1209,N_1128);
nor U1259 (N_1259,N_1249,N_1176);
or U1260 (N_1260,N_1143,N_1122);
and U1261 (N_1261,N_1063,N_1011);
nand U1262 (N_1262,N_1033,N_1238);
or U1263 (N_1263,N_1064,N_1053);
and U1264 (N_1264,N_1071,N_1177);
nand U1265 (N_1265,N_1067,N_1150);
nand U1266 (N_1266,N_1188,N_1197);
and U1267 (N_1267,N_1145,N_1165);
and U1268 (N_1268,N_1050,N_1038);
nor U1269 (N_1269,N_1178,N_1156);
and U1270 (N_1270,N_1153,N_1151);
or U1271 (N_1271,N_1204,N_1055);
or U1272 (N_1272,N_1019,N_1057);
nand U1273 (N_1273,N_1195,N_1084);
nor U1274 (N_1274,N_1208,N_1003);
nand U1275 (N_1275,N_1102,N_1191);
nand U1276 (N_1276,N_1111,N_1192);
nand U1277 (N_1277,N_1189,N_1173);
nand U1278 (N_1278,N_1056,N_1096);
and U1279 (N_1279,N_1058,N_1235);
or U1280 (N_1280,N_1239,N_1248);
or U1281 (N_1281,N_1004,N_1022);
and U1282 (N_1282,N_1231,N_1039);
nor U1283 (N_1283,N_1009,N_1021);
or U1284 (N_1284,N_1069,N_1095);
and U1285 (N_1285,N_1129,N_1030);
nand U1286 (N_1286,N_1170,N_1085);
xnor U1287 (N_1287,N_1115,N_1166);
and U1288 (N_1288,N_1097,N_1052);
and U1289 (N_1289,N_1007,N_1114);
nand U1290 (N_1290,N_1182,N_1081);
and U1291 (N_1291,N_1229,N_1136);
and U1292 (N_1292,N_1112,N_1040);
and U1293 (N_1293,N_1142,N_1131);
nor U1294 (N_1294,N_1123,N_1193);
and U1295 (N_1295,N_1005,N_1155);
and U1296 (N_1296,N_1218,N_1206);
and U1297 (N_1297,N_1046,N_1186);
or U1298 (N_1298,N_1137,N_1162);
nor U1299 (N_1299,N_1087,N_1032);
or U1300 (N_1300,N_1010,N_1232);
and U1301 (N_1301,N_1121,N_1219);
and U1302 (N_1302,N_1041,N_1037);
nand U1303 (N_1303,N_1138,N_1211);
or U1304 (N_1304,N_1075,N_1023);
or U1305 (N_1305,N_1077,N_1029);
nor U1306 (N_1306,N_1194,N_1015);
or U1307 (N_1307,N_1089,N_1220);
or U1308 (N_1308,N_1134,N_1017);
nand U1309 (N_1309,N_1043,N_1099);
nand U1310 (N_1310,N_1190,N_1158);
nand U1311 (N_1311,N_1243,N_1044);
nand U1312 (N_1312,N_1078,N_1117);
or U1313 (N_1313,N_1094,N_1100);
nor U1314 (N_1314,N_1199,N_1124);
nand U1315 (N_1315,N_1000,N_1020);
xor U1316 (N_1316,N_1181,N_1148);
nand U1317 (N_1317,N_1163,N_1223);
and U1318 (N_1318,N_1125,N_1161);
nand U1319 (N_1319,N_1226,N_1072);
nand U1320 (N_1320,N_1068,N_1215);
or U1321 (N_1321,N_1224,N_1247);
nor U1322 (N_1322,N_1228,N_1090);
nand U1323 (N_1323,N_1059,N_1086);
nand U1324 (N_1324,N_1093,N_1016);
nand U1325 (N_1325,N_1244,N_1113);
xnor U1326 (N_1326,N_1152,N_1042);
nand U1327 (N_1327,N_1002,N_1144);
nor U1328 (N_1328,N_1105,N_1074);
or U1329 (N_1329,N_1047,N_1227);
and U1330 (N_1330,N_1175,N_1207);
and U1331 (N_1331,N_1066,N_1008);
xnor U1332 (N_1332,N_1205,N_1234);
nor U1333 (N_1333,N_1240,N_1101);
nand U1334 (N_1334,N_1187,N_1060);
or U1335 (N_1335,N_1006,N_1076);
nor U1336 (N_1336,N_1103,N_1118);
or U1337 (N_1337,N_1168,N_1045);
nor U1338 (N_1338,N_1082,N_1147);
nand U1339 (N_1339,N_1200,N_1230);
and U1340 (N_1340,N_1167,N_1212);
nand U1341 (N_1341,N_1083,N_1013);
nor U1342 (N_1342,N_1172,N_1237);
nand U1343 (N_1343,N_1119,N_1036);
nor U1344 (N_1344,N_1091,N_1120);
and U1345 (N_1345,N_1171,N_1031);
and U1346 (N_1346,N_1127,N_1018);
and U1347 (N_1347,N_1196,N_1027);
nand U1348 (N_1348,N_1092,N_1159);
or U1349 (N_1349,N_1203,N_1174);
xor U1350 (N_1350,N_1169,N_1035);
xnor U1351 (N_1351,N_1139,N_1216);
nor U1352 (N_1352,N_1201,N_1116);
nand U1353 (N_1353,N_1051,N_1202);
and U1354 (N_1354,N_1241,N_1225);
xor U1355 (N_1355,N_1107,N_1079);
or U1356 (N_1356,N_1049,N_1160);
nor U1357 (N_1357,N_1236,N_1080);
nand U1358 (N_1358,N_1135,N_1104);
or U1359 (N_1359,N_1246,N_1157);
and U1360 (N_1360,N_1184,N_1214);
or U1361 (N_1361,N_1070,N_1126);
or U1362 (N_1362,N_1025,N_1048);
nand U1363 (N_1363,N_1054,N_1210);
nor U1364 (N_1364,N_1179,N_1233);
xor U1365 (N_1365,N_1106,N_1130);
nand U1366 (N_1366,N_1185,N_1108);
and U1367 (N_1367,N_1141,N_1154);
and U1368 (N_1368,N_1133,N_1221);
nand U1369 (N_1369,N_1245,N_1222);
nor U1370 (N_1370,N_1242,N_1034);
or U1371 (N_1371,N_1088,N_1213);
nor U1372 (N_1372,N_1024,N_1110);
or U1373 (N_1373,N_1028,N_1198);
nor U1374 (N_1374,N_1062,N_1098);
nor U1375 (N_1375,N_1095,N_1010);
xor U1376 (N_1376,N_1010,N_1184);
and U1377 (N_1377,N_1022,N_1086);
or U1378 (N_1378,N_1027,N_1057);
nor U1379 (N_1379,N_1177,N_1120);
and U1380 (N_1380,N_1116,N_1047);
xnor U1381 (N_1381,N_1191,N_1237);
and U1382 (N_1382,N_1154,N_1248);
xor U1383 (N_1383,N_1104,N_1181);
or U1384 (N_1384,N_1050,N_1222);
nand U1385 (N_1385,N_1051,N_1022);
and U1386 (N_1386,N_1222,N_1172);
and U1387 (N_1387,N_1125,N_1133);
xnor U1388 (N_1388,N_1181,N_1112);
or U1389 (N_1389,N_1165,N_1060);
and U1390 (N_1390,N_1170,N_1191);
or U1391 (N_1391,N_1138,N_1022);
or U1392 (N_1392,N_1161,N_1097);
or U1393 (N_1393,N_1160,N_1131);
nor U1394 (N_1394,N_1199,N_1021);
nor U1395 (N_1395,N_1124,N_1033);
nand U1396 (N_1396,N_1088,N_1198);
nor U1397 (N_1397,N_1100,N_1159);
or U1398 (N_1398,N_1239,N_1225);
or U1399 (N_1399,N_1154,N_1114);
or U1400 (N_1400,N_1196,N_1185);
nand U1401 (N_1401,N_1013,N_1227);
xnor U1402 (N_1402,N_1088,N_1142);
and U1403 (N_1403,N_1156,N_1025);
and U1404 (N_1404,N_1137,N_1063);
or U1405 (N_1405,N_1014,N_1240);
or U1406 (N_1406,N_1204,N_1031);
nand U1407 (N_1407,N_1146,N_1076);
or U1408 (N_1408,N_1091,N_1080);
or U1409 (N_1409,N_1035,N_1207);
and U1410 (N_1410,N_1115,N_1110);
or U1411 (N_1411,N_1156,N_1126);
or U1412 (N_1412,N_1185,N_1144);
nor U1413 (N_1413,N_1249,N_1180);
and U1414 (N_1414,N_1099,N_1239);
or U1415 (N_1415,N_1170,N_1096);
nor U1416 (N_1416,N_1152,N_1012);
nor U1417 (N_1417,N_1040,N_1004);
nand U1418 (N_1418,N_1221,N_1066);
nand U1419 (N_1419,N_1059,N_1103);
and U1420 (N_1420,N_1018,N_1240);
and U1421 (N_1421,N_1060,N_1115);
nor U1422 (N_1422,N_1105,N_1111);
nand U1423 (N_1423,N_1036,N_1173);
nand U1424 (N_1424,N_1211,N_1219);
or U1425 (N_1425,N_1139,N_1001);
nor U1426 (N_1426,N_1188,N_1124);
nor U1427 (N_1427,N_1119,N_1068);
nor U1428 (N_1428,N_1062,N_1093);
and U1429 (N_1429,N_1039,N_1093);
nor U1430 (N_1430,N_1061,N_1129);
and U1431 (N_1431,N_1223,N_1046);
nor U1432 (N_1432,N_1040,N_1237);
and U1433 (N_1433,N_1128,N_1240);
or U1434 (N_1434,N_1114,N_1081);
nor U1435 (N_1435,N_1035,N_1188);
or U1436 (N_1436,N_1191,N_1217);
nand U1437 (N_1437,N_1072,N_1086);
nand U1438 (N_1438,N_1166,N_1061);
and U1439 (N_1439,N_1203,N_1161);
xor U1440 (N_1440,N_1198,N_1027);
and U1441 (N_1441,N_1134,N_1141);
and U1442 (N_1442,N_1069,N_1207);
nand U1443 (N_1443,N_1155,N_1206);
and U1444 (N_1444,N_1203,N_1019);
and U1445 (N_1445,N_1239,N_1176);
or U1446 (N_1446,N_1200,N_1227);
or U1447 (N_1447,N_1181,N_1228);
or U1448 (N_1448,N_1044,N_1094);
nor U1449 (N_1449,N_1017,N_1185);
nand U1450 (N_1450,N_1102,N_1103);
nand U1451 (N_1451,N_1113,N_1199);
xor U1452 (N_1452,N_1042,N_1003);
or U1453 (N_1453,N_1024,N_1091);
nand U1454 (N_1454,N_1106,N_1125);
and U1455 (N_1455,N_1059,N_1032);
nand U1456 (N_1456,N_1053,N_1080);
nor U1457 (N_1457,N_1022,N_1095);
nor U1458 (N_1458,N_1100,N_1107);
or U1459 (N_1459,N_1082,N_1157);
or U1460 (N_1460,N_1164,N_1032);
and U1461 (N_1461,N_1068,N_1151);
and U1462 (N_1462,N_1113,N_1003);
or U1463 (N_1463,N_1144,N_1188);
nor U1464 (N_1464,N_1003,N_1111);
and U1465 (N_1465,N_1071,N_1170);
nand U1466 (N_1466,N_1134,N_1129);
nand U1467 (N_1467,N_1108,N_1040);
or U1468 (N_1468,N_1005,N_1129);
or U1469 (N_1469,N_1017,N_1033);
or U1470 (N_1470,N_1072,N_1187);
and U1471 (N_1471,N_1134,N_1164);
or U1472 (N_1472,N_1163,N_1083);
or U1473 (N_1473,N_1128,N_1046);
or U1474 (N_1474,N_1119,N_1104);
or U1475 (N_1475,N_1226,N_1215);
nor U1476 (N_1476,N_1220,N_1158);
or U1477 (N_1477,N_1130,N_1009);
nor U1478 (N_1478,N_1105,N_1053);
and U1479 (N_1479,N_1245,N_1233);
and U1480 (N_1480,N_1151,N_1054);
nor U1481 (N_1481,N_1020,N_1206);
nor U1482 (N_1482,N_1188,N_1097);
nor U1483 (N_1483,N_1194,N_1029);
or U1484 (N_1484,N_1106,N_1219);
and U1485 (N_1485,N_1049,N_1128);
xor U1486 (N_1486,N_1139,N_1042);
nor U1487 (N_1487,N_1191,N_1099);
nand U1488 (N_1488,N_1095,N_1063);
nor U1489 (N_1489,N_1201,N_1018);
and U1490 (N_1490,N_1191,N_1028);
or U1491 (N_1491,N_1070,N_1010);
nor U1492 (N_1492,N_1185,N_1190);
nor U1493 (N_1493,N_1138,N_1228);
nor U1494 (N_1494,N_1211,N_1155);
nor U1495 (N_1495,N_1043,N_1223);
and U1496 (N_1496,N_1222,N_1234);
and U1497 (N_1497,N_1049,N_1179);
and U1498 (N_1498,N_1176,N_1070);
nand U1499 (N_1499,N_1209,N_1161);
and U1500 (N_1500,N_1445,N_1457);
nand U1501 (N_1501,N_1470,N_1343);
nand U1502 (N_1502,N_1352,N_1392);
or U1503 (N_1503,N_1363,N_1347);
or U1504 (N_1504,N_1288,N_1495);
or U1505 (N_1505,N_1431,N_1446);
nand U1506 (N_1506,N_1432,N_1357);
or U1507 (N_1507,N_1306,N_1256);
nor U1508 (N_1508,N_1451,N_1327);
or U1509 (N_1509,N_1421,N_1391);
or U1510 (N_1510,N_1349,N_1354);
nand U1511 (N_1511,N_1268,N_1289);
xnor U1512 (N_1512,N_1266,N_1386);
or U1513 (N_1513,N_1498,N_1373);
nand U1514 (N_1514,N_1441,N_1379);
and U1515 (N_1515,N_1486,N_1479);
nor U1516 (N_1516,N_1448,N_1286);
nor U1517 (N_1517,N_1272,N_1338);
and U1518 (N_1518,N_1359,N_1316);
nand U1519 (N_1519,N_1489,N_1455);
nand U1520 (N_1520,N_1290,N_1324);
nand U1521 (N_1521,N_1459,N_1399);
and U1522 (N_1522,N_1488,N_1303);
and U1523 (N_1523,N_1331,N_1253);
xnor U1524 (N_1524,N_1396,N_1468);
nor U1525 (N_1525,N_1458,N_1333);
nor U1526 (N_1526,N_1430,N_1395);
xor U1527 (N_1527,N_1323,N_1465);
or U1528 (N_1528,N_1274,N_1315);
and U1529 (N_1529,N_1460,N_1319);
nand U1530 (N_1530,N_1302,N_1414);
nor U1531 (N_1531,N_1282,N_1318);
nor U1532 (N_1532,N_1275,N_1404);
and U1533 (N_1533,N_1280,N_1464);
nor U1534 (N_1534,N_1314,N_1341);
and U1535 (N_1535,N_1297,N_1440);
nand U1536 (N_1536,N_1376,N_1371);
and U1537 (N_1537,N_1361,N_1393);
xnor U1538 (N_1538,N_1418,N_1409);
xor U1539 (N_1539,N_1471,N_1362);
nand U1540 (N_1540,N_1330,N_1267);
and U1541 (N_1541,N_1408,N_1473);
nor U1542 (N_1542,N_1405,N_1255);
nand U1543 (N_1543,N_1287,N_1372);
or U1544 (N_1544,N_1251,N_1291);
or U1545 (N_1545,N_1353,N_1420);
nor U1546 (N_1546,N_1485,N_1276);
and U1547 (N_1547,N_1322,N_1284);
or U1548 (N_1548,N_1309,N_1452);
nor U1549 (N_1549,N_1425,N_1262);
or U1550 (N_1550,N_1348,N_1499);
nand U1551 (N_1551,N_1346,N_1412);
nand U1552 (N_1552,N_1497,N_1356);
and U1553 (N_1553,N_1403,N_1340);
nand U1554 (N_1554,N_1450,N_1400);
xnor U1555 (N_1555,N_1461,N_1258);
nor U1556 (N_1556,N_1261,N_1295);
and U1557 (N_1557,N_1493,N_1381);
nand U1558 (N_1558,N_1370,N_1467);
nor U1559 (N_1559,N_1398,N_1438);
or U1560 (N_1560,N_1285,N_1326);
nor U1561 (N_1561,N_1328,N_1380);
or U1562 (N_1562,N_1427,N_1476);
nand U1563 (N_1563,N_1320,N_1475);
or U1564 (N_1564,N_1435,N_1423);
and U1565 (N_1565,N_1394,N_1298);
nand U1566 (N_1566,N_1442,N_1250);
nor U1567 (N_1567,N_1387,N_1336);
nor U1568 (N_1568,N_1345,N_1337);
nor U1569 (N_1569,N_1310,N_1439);
and U1570 (N_1570,N_1252,N_1269);
or U1571 (N_1571,N_1351,N_1263);
or U1572 (N_1572,N_1454,N_1296);
or U1573 (N_1573,N_1254,N_1355);
and U1574 (N_1574,N_1389,N_1417);
nand U1575 (N_1575,N_1325,N_1321);
nor U1576 (N_1576,N_1483,N_1301);
and U1577 (N_1577,N_1474,N_1367);
nand U1578 (N_1578,N_1294,N_1329);
xor U1579 (N_1579,N_1419,N_1490);
and U1580 (N_1580,N_1368,N_1384);
and U1581 (N_1581,N_1273,N_1463);
nor U1582 (N_1582,N_1334,N_1410);
xor U1583 (N_1583,N_1304,N_1312);
and U1584 (N_1584,N_1364,N_1481);
nand U1585 (N_1585,N_1437,N_1335);
or U1586 (N_1586,N_1277,N_1426);
xor U1587 (N_1587,N_1478,N_1480);
nand U1588 (N_1588,N_1482,N_1271);
nor U1589 (N_1589,N_1388,N_1494);
xnor U1590 (N_1590,N_1411,N_1443);
xnor U1591 (N_1591,N_1358,N_1434);
or U1592 (N_1592,N_1265,N_1449);
or U1593 (N_1593,N_1402,N_1378);
nand U1594 (N_1594,N_1390,N_1270);
and U1595 (N_1595,N_1484,N_1444);
xnor U1596 (N_1596,N_1424,N_1292);
and U1597 (N_1597,N_1456,N_1436);
or U1598 (N_1598,N_1416,N_1365);
xor U1599 (N_1599,N_1278,N_1307);
or U1600 (N_1600,N_1466,N_1491);
and U1601 (N_1601,N_1281,N_1453);
nor U1602 (N_1602,N_1308,N_1350);
and U1603 (N_1603,N_1311,N_1413);
or U1604 (N_1604,N_1305,N_1283);
nor U1605 (N_1605,N_1487,N_1422);
nor U1606 (N_1606,N_1382,N_1299);
nor U1607 (N_1607,N_1257,N_1279);
nor U1608 (N_1608,N_1383,N_1293);
nand U1609 (N_1609,N_1375,N_1433);
nand U1610 (N_1610,N_1344,N_1415);
and U1611 (N_1611,N_1332,N_1264);
nand U1612 (N_1612,N_1492,N_1406);
nand U1613 (N_1613,N_1401,N_1313);
nand U1614 (N_1614,N_1360,N_1259);
nor U1615 (N_1615,N_1342,N_1462);
or U1616 (N_1616,N_1429,N_1339);
nor U1617 (N_1617,N_1369,N_1300);
or U1618 (N_1618,N_1374,N_1397);
or U1619 (N_1619,N_1447,N_1385);
and U1620 (N_1620,N_1260,N_1428);
nand U1621 (N_1621,N_1469,N_1407);
nand U1622 (N_1622,N_1496,N_1477);
nor U1623 (N_1623,N_1472,N_1377);
or U1624 (N_1624,N_1317,N_1366);
nand U1625 (N_1625,N_1310,N_1411);
nor U1626 (N_1626,N_1255,N_1300);
xor U1627 (N_1627,N_1273,N_1468);
nand U1628 (N_1628,N_1404,N_1371);
nand U1629 (N_1629,N_1362,N_1492);
nor U1630 (N_1630,N_1313,N_1460);
and U1631 (N_1631,N_1369,N_1381);
or U1632 (N_1632,N_1371,N_1309);
and U1633 (N_1633,N_1355,N_1465);
and U1634 (N_1634,N_1414,N_1492);
nor U1635 (N_1635,N_1295,N_1307);
nand U1636 (N_1636,N_1373,N_1260);
nor U1637 (N_1637,N_1441,N_1473);
and U1638 (N_1638,N_1257,N_1250);
and U1639 (N_1639,N_1406,N_1366);
and U1640 (N_1640,N_1401,N_1361);
or U1641 (N_1641,N_1488,N_1339);
nor U1642 (N_1642,N_1429,N_1461);
and U1643 (N_1643,N_1475,N_1416);
and U1644 (N_1644,N_1317,N_1293);
or U1645 (N_1645,N_1406,N_1323);
and U1646 (N_1646,N_1367,N_1380);
or U1647 (N_1647,N_1451,N_1309);
or U1648 (N_1648,N_1393,N_1457);
nor U1649 (N_1649,N_1403,N_1290);
nor U1650 (N_1650,N_1337,N_1406);
or U1651 (N_1651,N_1423,N_1279);
or U1652 (N_1652,N_1405,N_1441);
nor U1653 (N_1653,N_1456,N_1429);
nand U1654 (N_1654,N_1454,N_1466);
nor U1655 (N_1655,N_1298,N_1280);
nor U1656 (N_1656,N_1381,N_1426);
or U1657 (N_1657,N_1309,N_1261);
nor U1658 (N_1658,N_1487,N_1263);
or U1659 (N_1659,N_1315,N_1461);
nor U1660 (N_1660,N_1335,N_1304);
or U1661 (N_1661,N_1452,N_1427);
xnor U1662 (N_1662,N_1269,N_1345);
nor U1663 (N_1663,N_1400,N_1300);
nor U1664 (N_1664,N_1453,N_1327);
nor U1665 (N_1665,N_1376,N_1305);
xor U1666 (N_1666,N_1485,N_1345);
nand U1667 (N_1667,N_1350,N_1466);
nor U1668 (N_1668,N_1270,N_1289);
nor U1669 (N_1669,N_1285,N_1423);
or U1670 (N_1670,N_1381,N_1326);
nand U1671 (N_1671,N_1368,N_1379);
nand U1672 (N_1672,N_1291,N_1354);
and U1673 (N_1673,N_1382,N_1492);
and U1674 (N_1674,N_1276,N_1284);
nor U1675 (N_1675,N_1490,N_1293);
nor U1676 (N_1676,N_1410,N_1428);
and U1677 (N_1677,N_1434,N_1284);
nor U1678 (N_1678,N_1394,N_1446);
nor U1679 (N_1679,N_1315,N_1452);
xor U1680 (N_1680,N_1307,N_1436);
nor U1681 (N_1681,N_1438,N_1335);
nor U1682 (N_1682,N_1471,N_1480);
or U1683 (N_1683,N_1274,N_1298);
and U1684 (N_1684,N_1455,N_1369);
nor U1685 (N_1685,N_1269,N_1497);
nand U1686 (N_1686,N_1417,N_1331);
nand U1687 (N_1687,N_1458,N_1387);
or U1688 (N_1688,N_1382,N_1311);
or U1689 (N_1689,N_1319,N_1450);
or U1690 (N_1690,N_1416,N_1284);
nand U1691 (N_1691,N_1476,N_1292);
xor U1692 (N_1692,N_1269,N_1348);
nand U1693 (N_1693,N_1332,N_1423);
nand U1694 (N_1694,N_1376,N_1446);
nand U1695 (N_1695,N_1287,N_1409);
nor U1696 (N_1696,N_1463,N_1346);
nor U1697 (N_1697,N_1433,N_1385);
nand U1698 (N_1698,N_1368,N_1491);
and U1699 (N_1699,N_1284,N_1372);
nand U1700 (N_1700,N_1482,N_1371);
or U1701 (N_1701,N_1261,N_1329);
and U1702 (N_1702,N_1308,N_1288);
and U1703 (N_1703,N_1260,N_1415);
xnor U1704 (N_1704,N_1276,N_1316);
nor U1705 (N_1705,N_1409,N_1254);
and U1706 (N_1706,N_1408,N_1468);
and U1707 (N_1707,N_1462,N_1281);
nand U1708 (N_1708,N_1405,N_1338);
nand U1709 (N_1709,N_1334,N_1492);
or U1710 (N_1710,N_1320,N_1264);
or U1711 (N_1711,N_1425,N_1446);
or U1712 (N_1712,N_1396,N_1282);
nand U1713 (N_1713,N_1324,N_1414);
nand U1714 (N_1714,N_1385,N_1273);
xnor U1715 (N_1715,N_1484,N_1490);
and U1716 (N_1716,N_1433,N_1259);
and U1717 (N_1717,N_1349,N_1496);
nor U1718 (N_1718,N_1488,N_1263);
and U1719 (N_1719,N_1485,N_1480);
nand U1720 (N_1720,N_1412,N_1265);
or U1721 (N_1721,N_1380,N_1320);
nor U1722 (N_1722,N_1472,N_1314);
nand U1723 (N_1723,N_1421,N_1278);
nor U1724 (N_1724,N_1377,N_1285);
nand U1725 (N_1725,N_1261,N_1346);
and U1726 (N_1726,N_1294,N_1333);
or U1727 (N_1727,N_1482,N_1324);
and U1728 (N_1728,N_1253,N_1329);
nand U1729 (N_1729,N_1451,N_1303);
and U1730 (N_1730,N_1352,N_1496);
and U1731 (N_1731,N_1307,N_1410);
nor U1732 (N_1732,N_1293,N_1272);
and U1733 (N_1733,N_1280,N_1431);
nand U1734 (N_1734,N_1347,N_1281);
nor U1735 (N_1735,N_1475,N_1267);
or U1736 (N_1736,N_1414,N_1280);
xor U1737 (N_1737,N_1345,N_1431);
nand U1738 (N_1738,N_1470,N_1352);
nor U1739 (N_1739,N_1429,N_1491);
nand U1740 (N_1740,N_1299,N_1435);
nand U1741 (N_1741,N_1446,N_1359);
and U1742 (N_1742,N_1347,N_1321);
nor U1743 (N_1743,N_1252,N_1460);
nor U1744 (N_1744,N_1452,N_1479);
or U1745 (N_1745,N_1302,N_1373);
nand U1746 (N_1746,N_1398,N_1377);
xor U1747 (N_1747,N_1343,N_1369);
and U1748 (N_1748,N_1456,N_1336);
nand U1749 (N_1749,N_1423,N_1434);
nor U1750 (N_1750,N_1660,N_1630);
and U1751 (N_1751,N_1704,N_1604);
or U1752 (N_1752,N_1529,N_1712);
or U1753 (N_1753,N_1510,N_1585);
nand U1754 (N_1754,N_1749,N_1505);
or U1755 (N_1755,N_1594,N_1747);
or U1756 (N_1756,N_1745,N_1540);
nor U1757 (N_1757,N_1654,N_1705);
nand U1758 (N_1758,N_1658,N_1526);
nor U1759 (N_1759,N_1680,N_1545);
nand U1760 (N_1760,N_1564,N_1702);
nor U1761 (N_1761,N_1703,N_1619);
and U1762 (N_1762,N_1563,N_1713);
nand U1763 (N_1763,N_1531,N_1632);
or U1764 (N_1764,N_1512,N_1681);
nor U1765 (N_1765,N_1655,N_1506);
nand U1766 (N_1766,N_1559,N_1589);
nand U1767 (N_1767,N_1501,N_1537);
nor U1768 (N_1768,N_1666,N_1700);
and U1769 (N_1769,N_1565,N_1732);
nor U1770 (N_1770,N_1688,N_1514);
or U1771 (N_1771,N_1687,N_1611);
or U1772 (N_1772,N_1715,N_1689);
nand U1773 (N_1773,N_1581,N_1708);
xor U1774 (N_1774,N_1595,N_1603);
nor U1775 (N_1775,N_1651,N_1530);
nor U1776 (N_1776,N_1624,N_1523);
and U1777 (N_1777,N_1590,N_1612);
or U1778 (N_1778,N_1676,N_1601);
and U1779 (N_1779,N_1527,N_1509);
or U1780 (N_1780,N_1742,N_1574);
and U1781 (N_1781,N_1562,N_1728);
or U1782 (N_1782,N_1692,N_1580);
and U1783 (N_1783,N_1733,N_1606);
xnor U1784 (N_1784,N_1672,N_1519);
nor U1785 (N_1785,N_1738,N_1570);
nand U1786 (N_1786,N_1522,N_1552);
nand U1787 (N_1787,N_1507,N_1588);
nand U1788 (N_1788,N_1635,N_1697);
and U1789 (N_1789,N_1536,N_1516);
or U1790 (N_1790,N_1546,N_1723);
nand U1791 (N_1791,N_1698,N_1549);
nor U1792 (N_1792,N_1679,N_1504);
nor U1793 (N_1793,N_1620,N_1548);
nand U1794 (N_1794,N_1664,N_1542);
and U1795 (N_1795,N_1541,N_1613);
and U1796 (N_1796,N_1616,N_1724);
or U1797 (N_1797,N_1568,N_1710);
or U1798 (N_1798,N_1627,N_1716);
xor U1799 (N_1799,N_1577,N_1650);
nand U1800 (N_1800,N_1561,N_1633);
nor U1801 (N_1801,N_1520,N_1736);
or U1802 (N_1802,N_1730,N_1513);
and U1803 (N_1803,N_1569,N_1727);
and U1804 (N_1804,N_1586,N_1711);
and U1805 (N_1805,N_1631,N_1684);
or U1806 (N_1806,N_1642,N_1503);
nor U1807 (N_1807,N_1634,N_1709);
nor U1808 (N_1808,N_1535,N_1538);
or U1809 (N_1809,N_1582,N_1722);
or U1810 (N_1810,N_1502,N_1525);
nand U1811 (N_1811,N_1739,N_1553);
or U1812 (N_1812,N_1572,N_1593);
nand U1813 (N_1813,N_1640,N_1534);
and U1814 (N_1814,N_1626,N_1682);
or U1815 (N_1815,N_1659,N_1748);
and U1816 (N_1816,N_1584,N_1638);
nand U1817 (N_1817,N_1677,N_1648);
nor U1818 (N_1818,N_1695,N_1521);
nand U1819 (N_1819,N_1614,N_1735);
xnor U1820 (N_1820,N_1579,N_1557);
nand U1821 (N_1821,N_1696,N_1701);
and U1822 (N_1822,N_1587,N_1720);
nor U1823 (N_1823,N_1737,N_1678);
xnor U1824 (N_1824,N_1741,N_1707);
nand U1825 (N_1825,N_1556,N_1734);
and U1826 (N_1826,N_1656,N_1667);
or U1827 (N_1827,N_1669,N_1524);
and U1828 (N_1828,N_1691,N_1625);
or U1829 (N_1829,N_1591,N_1743);
nor U1830 (N_1830,N_1628,N_1517);
nand U1831 (N_1831,N_1636,N_1539);
nor U1832 (N_1832,N_1641,N_1718);
nor U1833 (N_1833,N_1533,N_1726);
or U1834 (N_1834,N_1685,N_1602);
and U1835 (N_1835,N_1573,N_1609);
nor U1836 (N_1836,N_1637,N_1621);
and U1837 (N_1837,N_1551,N_1744);
xor U1838 (N_1838,N_1583,N_1615);
or U1839 (N_1839,N_1694,N_1663);
and U1840 (N_1840,N_1729,N_1508);
nor U1841 (N_1841,N_1693,N_1605);
and U1842 (N_1842,N_1511,N_1717);
nand U1843 (N_1843,N_1600,N_1518);
nand U1844 (N_1844,N_1560,N_1647);
and U1845 (N_1845,N_1653,N_1674);
and U1846 (N_1846,N_1622,N_1657);
xnor U1847 (N_1847,N_1532,N_1592);
and U1848 (N_1848,N_1629,N_1596);
nor U1849 (N_1849,N_1670,N_1683);
nand U1850 (N_1850,N_1607,N_1699);
and U1851 (N_1851,N_1686,N_1618);
nand U1852 (N_1852,N_1721,N_1675);
and U1853 (N_1853,N_1610,N_1746);
or U1854 (N_1854,N_1500,N_1643);
nor U1855 (N_1855,N_1608,N_1567);
and U1856 (N_1856,N_1644,N_1578);
nand U1857 (N_1857,N_1673,N_1719);
nand U1858 (N_1858,N_1575,N_1555);
nand U1859 (N_1859,N_1665,N_1571);
or U1860 (N_1860,N_1671,N_1597);
and U1861 (N_1861,N_1662,N_1547);
or U1862 (N_1862,N_1661,N_1740);
nor U1863 (N_1863,N_1543,N_1550);
or U1864 (N_1864,N_1646,N_1652);
nor U1865 (N_1865,N_1617,N_1599);
or U1866 (N_1866,N_1566,N_1725);
nor U1867 (N_1867,N_1544,N_1649);
and U1868 (N_1868,N_1731,N_1576);
xor U1869 (N_1869,N_1668,N_1645);
and U1870 (N_1870,N_1598,N_1558);
nand U1871 (N_1871,N_1515,N_1554);
or U1872 (N_1872,N_1706,N_1690);
nand U1873 (N_1873,N_1639,N_1714);
and U1874 (N_1874,N_1623,N_1528);
and U1875 (N_1875,N_1626,N_1558);
nand U1876 (N_1876,N_1537,N_1615);
nand U1877 (N_1877,N_1513,N_1554);
or U1878 (N_1878,N_1505,N_1529);
and U1879 (N_1879,N_1632,N_1532);
or U1880 (N_1880,N_1714,N_1707);
nand U1881 (N_1881,N_1536,N_1690);
nor U1882 (N_1882,N_1744,N_1516);
nor U1883 (N_1883,N_1589,N_1672);
nand U1884 (N_1884,N_1626,N_1671);
or U1885 (N_1885,N_1622,N_1570);
nand U1886 (N_1886,N_1614,N_1717);
nor U1887 (N_1887,N_1660,N_1677);
nand U1888 (N_1888,N_1733,N_1507);
xnor U1889 (N_1889,N_1618,N_1685);
and U1890 (N_1890,N_1508,N_1515);
nor U1891 (N_1891,N_1644,N_1559);
xnor U1892 (N_1892,N_1533,N_1672);
and U1893 (N_1893,N_1541,N_1744);
nor U1894 (N_1894,N_1566,N_1504);
and U1895 (N_1895,N_1749,N_1685);
and U1896 (N_1896,N_1615,N_1675);
nand U1897 (N_1897,N_1551,N_1579);
nand U1898 (N_1898,N_1720,N_1586);
or U1899 (N_1899,N_1693,N_1540);
nor U1900 (N_1900,N_1592,N_1619);
or U1901 (N_1901,N_1591,N_1649);
or U1902 (N_1902,N_1605,N_1644);
or U1903 (N_1903,N_1741,N_1530);
or U1904 (N_1904,N_1642,N_1725);
and U1905 (N_1905,N_1697,N_1597);
nand U1906 (N_1906,N_1590,N_1504);
nor U1907 (N_1907,N_1614,N_1541);
and U1908 (N_1908,N_1560,N_1681);
or U1909 (N_1909,N_1733,N_1598);
nand U1910 (N_1910,N_1510,N_1652);
nand U1911 (N_1911,N_1633,N_1749);
nand U1912 (N_1912,N_1714,N_1648);
nand U1913 (N_1913,N_1728,N_1677);
and U1914 (N_1914,N_1526,N_1673);
and U1915 (N_1915,N_1637,N_1642);
nand U1916 (N_1916,N_1584,N_1532);
nor U1917 (N_1917,N_1731,N_1659);
nand U1918 (N_1918,N_1708,N_1695);
nor U1919 (N_1919,N_1566,N_1505);
and U1920 (N_1920,N_1700,N_1590);
or U1921 (N_1921,N_1506,N_1613);
nand U1922 (N_1922,N_1589,N_1590);
xor U1923 (N_1923,N_1556,N_1559);
xor U1924 (N_1924,N_1542,N_1594);
or U1925 (N_1925,N_1690,N_1623);
nand U1926 (N_1926,N_1680,N_1745);
nand U1927 (N_1927,N_1600,N_1650);
and U1928 (N_1928,N_1625,N_1556);
and U1929 (N_1929,N_1724,N_1579);
xor U1930 (N_1930,N_1717,N_1638);
nand U1931 (N_1931,N_1609,N_1586);
and U1932 (N_1932,N_1702,N_1737);
nor U1933 (N_1933,N_1631,N_1663);
nor U1934 (N_1934,N_1635,N_1609);
nor U1935 (N_1935,N_1682,N_1649);
and U1936 (N_1936,N_1646,N_1541);
nand U1937 (N_1937,N_1591,N_1512);
and U1938 (N_1938,N_1648,N_1526);
xor U1939 (N_1939,N_1536,N_1611);
nor U1940 (N_1940,N_1644,N_1510);
or U1941 (N_1941,N_1728,N_1602);
or U1942 (N_1942,N_1721,N_1509);
nor U1943 (N_1943,N_1530,N_1574);
xor U1944 (N_1944,N_1689,N_1706);
nor U1945 (N_1945,N_1611,N_1612);
or U1946 (N_1946,N_1715,N_1684);
and U1947 (N_1947,N_1655,N_1712);
nor U1948 (N_1948,N_1559,N_1540);
xor U1949 (N_1949,N_1694,N_1664);
nand U1950 (N_1950,N_1632,N_1735);
nand U1951 (N_1951,N_1521,N_1558);
nor U1952 (N_1952,N_1635,N_1501);
nor U1953 (N_1953,N_1679,N_1691);
xor U1954 (N_1954,N_1715,N_1548);
or U1955 (N_1955,N_1719,N_1743);
and U1956 (N_1956,N_1618,N_1593);
nand U1957 (N_1957,N_1670,N_1666);
or U1958 (N_1958,N_1701,N_1604);
and U1959 (N_1959,N_1620,N_1729);
nor U1960 (N_1960,N_1543,N_1738);
nor U1961 (N_1961,N_1633,N_1584);
nor U1962 (N_1962,N_1696,N_1730);
nand U1963 (N_1963,N_1656,N_1570);
and U1964 (N_1964,N_1687,N_1522);
and U1965 (N_1965,N_1629,N_1594);
or U1966 (N_1966,N_1607,N_1731);
and U1967 (N_1967,N_1520,N_1597);
or U1968 (N_1968,N_1561,N_1669);
nand U1969 (N_1969,N_1749,N_1644);
nor U1970 (N_1970,N_1731,N_1735);
or U1971 (N_1971,N_1694,N_1523);
nand U1972 (N_1972,N_1611,N_1680);
nand U1973 (N_1973,N_1590,N_1721);
nand U1974 (N_1974,N_1589,N_1655);
nor U1975 (N_1975,N_1745,N_1660);
nand U1976 (N_1976,N_1694,N_1646);
and U1977 (N_1977,N_1546,N_1628);
or U1978 (N_1978,N_1715,N_1545);
and U1979 (N_1979,N_1733,N_1506);
or U1980 (N_1980,N_1646,N_1673);
xnor U1981 (N_1981,N_1598,N_1678);
nor U1982 (N_1982,N_1696,N_1540);
or U1983 (N_1983,N_1549,N_1586);
xor U1984 (N_1984,N_1590,N_1564);
nand U1985 (N_1985,N_1577,N_1581);
nor U1986 (N_1986,N_1686,N_1537);
nand U1987 (N_1987,N_1715,N_1553);
or U1988 (N_1988,N_1586,N_1747);
or U1989 (N_1989,N_1568,N_1507);
and U1990 (N_1990,N_1747,N_1580);
xnor U1991 (N_1991,N_1581,N_1628);
or U1992 (N_1992,N_1660,N_1563);
nor U1993 (N_1993,N_1732,N_1684);
and U1994 (N_1994,N_1733,N_1693);
or U1995 (N_1995,N_1632,N_1554);
nand U1996 (N_1996,N_1565,N_1637);
or U1997 (N_1997,N_1502,N_1659);
nor U1998 (N_1998,N_1677,N_1511);
nand U1999 (N_1999,N_1515,N_1711);
nor U2000 (N_2000,N_1821,N_1799);
or U2001 (N_2001,N_1981,N_1861);
or U2002 (N_2002,N_1776,N_1947);
or U2003 (N_2003,N_1915,N_1779);
nand U2004 (N_2004,N_1899,N_1844);
nand U2005 (N_2005,N_1818,N_1983);
or U2006 (N_2006,N_1880,N_1771);
or U2007 (N_2007,N_1960,N_1887);
nand U2008 (N_2008,N_1843,N_1751);
nor U2009 (N_2009,N_1874,N_1951);
nand U2010 (N_2010,N_1988,N_1793);
nor U2011 (N_2011,N_1854,N_1858);
and U2012 (N_2012,N_1830,N_1949);
and U2013 (N_2013,N_1929,N_1872);
nor U2014 (N_2014,N_1803,N_1897);
nand U2015 (N_2015,N_1800,N_1927);
nor U2016 (N_2016,N_1797,N_1795);
nand U2017 (N_2017,N_1754,N_1848);
and U2018 (N_2018,N_1817,N_1807);
nand U2019 (N_2019,N_1783,N_1878);
and U2020 (N_2020,N_1856,N_1928);
nand U2021 (N_2021,N_1908,N_1785);
nand U2022 (N_2022,N_1999,N_1823);
or U2023 (N_2023,N_1790,N_1774);
or U2024 (N_2024,N_1812,N_1913);
and U2025 (N_2025,N_1882,N_1796);
nand U2026 (N_2026,N_1995,N_1936);
and U2027 (N_2027,N_1922,N_1868);
xnor U2028 (N_2028,N_1946,N_1903);
or U2029 (N_2029,N_1784,N_1879);
nor U2030 (N_2030,N_1850,N_1905);
nand U2031 (N_2031,N_1883,N_1820);
xnor U2032 (N_2032,N_1923,N_1958);
or U2033 (N_2033,N_1842,N_1808);
xor U2034 (N_2034,N_1849,N_1998);
or U2035 (N_2035,N_1930,N_1968);
or U2036 (N_2036,N_1901,N_1953);
and U2037 (N_2037,N_1889,N_1787);
nor U2038 (N_2038,N_1891,N_1833);
and U2039 (N_2039,N_1926,N_1943);
or U2040 (N_2040,N_1839,N_1909);
and U2041 (N_2041,N_1965,N_1869);
or U2042 (N_2042,N_1758,N_1841);
nand U2043 (N_2043,N_1788,N_1757);
xor U2044 (N_2044,N_1977,N_1910);
or U2045 (N_2045,N_1851,N_1822);
xor U2046 (N_2046,N_1945,N_1881);
nand U2047 (N_2047,N_1764,N_1917);
and U2048 (N_2048,N_1873,N_1840);
nand U2049 (N_2049,N_1786,N_1907);
and U2050 (N_2050,N_1763,N_1975);
nand U2051 (N_2051,N_1978,N_1811);
nand U2052 (N_2052,N_1974,N_1939);
and U2053 (N_2053,N_1898,N_1932);
nor U2054 (N_2054,N_1914,N_1919);
and U2055 (N_2055,N_1967,N_1772);
and U2056 (N_2056,N_1831,N_1985);
xor U2057 (N_2057,N_1924,N_1934);
nor U2058 (N_2058,N_1806,N_1896);
and U2059 (N_2059,N_1954,N_1775);
or U2060 (N_2060,N_1885,N_1753);
nor U2061 (N_2061,N_1778,N_1816);
and U2062 (N_2062,N_1752,N_1791);
nor U2063 (N_2063,N_1768,N_1870);
or U2064 (N_2064,N_1987,N_1838);
and U2065 (N_2065,N_1759,N_1931);
or U2066 (N_2066,N_1859,N_1895);
or U2067 (N_2067,N_1962,N_1765);
or U2068 (N_2068,N_1888,N_1846);
nor U2069 (N_2069,N_1819,N_1837);
nor U2070 (N_2070,N_1828,N_1971);
xnor U2071 (N_2071,N_1857,N_1862);
nor U2072 (N_2072,N_1762,N_1760);
nor U2073 (N_2073,N_1836,N_1884);
nor U2074 (N_2074,N_1886,N_1855);
nor U2075 (N_2075,N_1921,N_1911);
nor U2076 (N_2076,N_1990,N_1991);
and U2077 (N_2077,N_1918,N_1860);
and U2078 (N_2078,N_1773,N_1809);
nand U2079 (N_2079,N_1876,N_1890);
nand U2080 (N_2080,N_1813,N_1864);
and U2081 (N_2081,N_1847,N_1994);
nor U2082 (N_2082,N_1997,N_1794);
or U2083 (N_2083,N_1940,N_1979);
nor U2084 (N_2084,N_1866,N_1970);
xor U2085 (N_2085,N_1877,N_1916);
nor U2086 (N_2086,N_1982,N_1989);
and U2087 (N_2087,N_1777,N_1938);
or U2088 (N_2088,N_1755,N_1829);
or U2089 (N_2089,N_1972,N_1766);
xor U2090 (N_2090,N_1825,N_1845);
nor U2091 (N_2091,N_1832,N_1941);
or U2092 (N_2092,N_1875,N_1781);
nand U2093 (N_2093,N_1902,N_1935);
and U2094 (N_2094,N_1944,N_1792);
nor U2095 (N_2095,N_1814,N_1892);
nand U2096 (N_2096,N_1770,N_1893);
nand U2097 (N_2097,N_1801,N_1992);
or U2098 (N_2098,N_1925,N_1980);
and U2099 (N_2099,N_1802,N_1853);
and U2100 (N_2100,N_1789,N_1761);
nand U2101 (N_2101,N_1769,N_1782);
xnor U2102 (N_2102,N_1948,N_1933);
nand U2103 (N_2103,N_1986,N_1993);
nor U2104 (N_2104,N_1942,N_1984);
xor U2105 (N_2105,N_1950,N_1867);
nor U2106 (N_2106,N_1804,N_1956);
or U2107 (N_2107,N_1805,N_1952);
or U2108 (N_2108,N_1996,N_1969);
xnor U2109 (N_2109,N_1973,N_1920);
xor U2110 (N_2110,N_1912,N_1815);
nand U2111 (N_2111,N_1767,N_1959);
xor U2112 (N_2112,N_1894,N_1756);
nor U2113 (N_2113,N_1750,N_1871);
nor U2114 (N_2114,N_1835,N_1826);
or U2115 (N_2115,N_1906,N_1852);
nor U2116 (N_2116,N_1780,N_1966);
nand U2117 (N_2117,N_1810,N_1937);
nor U2118 (N_2118,N_1955,N_1904);
and U2119 (N_2119,N_1865,N_1834);
nor U2120 (N_2120,N_1957,N_1827);
and U2121 (N_2121,N_1964,N_1976);
nor U2122 (N_2122,N_1963,N_1863);
nand U2123 (N_2123,N_1824,N_1798);
nor U2124 (N_2124,N_1961,N_1900);
nor U2125 (N_2125,N_1954,N_1944);
xnor U2126 (N_2126,N_1811,N_1868);
nand U2127 (N_2127,N_1774,N_1843);
nor U2128 (N_2128,N_1956,N_1986);
nor U2129 (N_2129,N_1872,N_1955);
nand U2130 (N_2130,N_1869,N_1810);
nor U2131 (N_2131,N_1819,N_1991);
nor U2132 (N_2132,N_1820,N_1962);
and U2133 (N_2133,N_1985,N_1816);
nor U2134 (N_2134,N_1807,N_1899);
nand U2135 (N_2135,N_1882,N_1982);
or U2136 (N_2136,N_1969,N_1977);
nand U2137 (N_2137,N_1848,N_1925);
and U2138 (N_2138,N_1864,N_1934);
nand U2139 (N_2139,N_1898,N_1993);
nand U2140 (N_2140,N_1907,N_1770);
and U2141 (N_2141,N_1867,N_1783);
nand U2142 (N_2142,N_1993,N_1875);
xor U2143 (N_2143,N_1919,N_1830);
and U2144 (N_2144,N_1993,N_1870);
nand U2145 (N_2145,N_1830,N_1907);
nor U2146 (N_2146,N_1810,N_1947);
nand U2147 (N_2147,N_1805,N_1964);
nor U2148 (N_2148,N_1925,N_1755);
nor U2149 (N_2149,N_1785,N_1993);
nor U2150 (N_2150,N_1924,N_1995);
xnor U2151 (N_2151,N_1891,N_1923);
and U2152 (N_2152,N_1928,N_1838);
xnor U2153 (N_2153,N_1955,N_1780);
or U2154 (N_2154,N_1925,N_1805);
nand U2155 (N_2155,N_1832,N_1778);
nor U2156 (N_2156,N_1945,N_1994);
nor U2157 (N_2157,N_1821,N_1901);
or U2158 (N_2158,N_1925,N_1989);
or U2159 (N_2159,N_1920,N_1860);
nand U2160 (N_2160,N_1875,N_1980);
nor U2161 (N_2161,N_1888,N_1857);
or U2162 (N_2162,N_1751,N_1955);
xor U2163 (N_2163,N_1852,N_1830);
and U2164 (N_2164,N_1769,N_1965);
and U2165 (N_2165,N_1751,N_1898);
or U2166 (N_2166,N_1801,N_1809);
and U2167 (N_2167,N_1823,N_1810);
nand U2168 (N_2168,N_1907,N_1920);
xor U2169 (N_2169,N_1782,N_1881);
nand U2170 (N_2170,N_1863,N_1976);
nor U2171 (N_2171,N_1901,N_1800);
and U2172 (N_2172,N_1941,N_1787);
nor U2173 (N_2173,N_1861,N_1896);
and U2174 (N_2174,N_1959,N_1970);
nand U2175 (N_2175,N_1810,N_1955);
or U2176 (N_2176,N_1980,N_1909);
nand U2177 (N_2177,N_1750,N_1764);
nor U2178 (N_2178,N_1859,N_1838);
or U2179 (N_2179,N_1772,N_1836);
nor U2180 (N_2180,N_1788,N_1948);
or U2181 (N_2181,N_1843,N_1764);
nor U2182 (N_2182,N_1820,N_1818);
nand U2183 (N_2183,N_1858,N_1828);
or U2184 (N_2184,N_1898,N_1927);
nand U2185 (N_2185,N_1964,N_1819);
or U2186 (N_2186,N_1797,N_1984);
nand U2187 (N_2187,N_1962,N_1848);
nand U2188 (N_2188,N_1829,N_1977);
nand U2189 (N_2189,N_1915,N_1967);
and U2190 (N_2190,N_1780,N_1947);
nand U2191 (N_2191,N_1917,N_1961);
or U2192 (N_2192,N_1987,N_1793);
nand U2193 (N_2193,N_1971,N_1836);
and U2194 (N_2194,N_1904,N_1917);
and U2195 (N_2195,N_1798,N_1750);
xnor U2196 (N_2196,N_1761,N_1930);
nand U2197 (N_2197,N_1955,N_1948);
nor U2198 (N_2198,N_1848,N_1966);
or U2199 (N_2199,N_1774,N_1927);
or U2200 (N_2200,N_1927,N_1847);
nand U2201 (N_2201,N_1948,N_1899);
nand U2202 (N_2202,N_1811,N_1786);
and U2203 (N_2203,N_1909,N_1827);
xnor U2204 (N_2204,N_1946,N_1886);
xor U2205 (N_2205,N_1923,N_1942);
xnor U2206 (N_2206,N_1794,N_1836);
or U2207 (N_2207,N_1977,N_1896);
nor U2208 (N_2208,N_1850,N_1788);
and U2209 (N_2209,N_1864,N_1765);
xor U2210 (N_2210,N_1878,N_1942);
nor U2211 (N_2211,N_1879,N_1844);
nand U2212 (N_2212,N_1963,N_1986);
nand U2213 (N_2213,N_1991,N_1768);
nand U2214 (N_2214,N_1938,N_1794);
nand U2215 (N_2215,N_1908,N_1827);
or U2216 (N_2216,N_1849,N_1985);
nor U2217 (N_2217,N_1766,N_1848);
and U2218 (N_2218,N_1938,N_1940);
and U2219 (N_2219,N_1917,N_1945);
and U2220 (N_2220,N_1825,N_1808);
xnor U2221 (N_2221,N_1846,N_1980);
xor U2222 (N_2222,N_1966,N_1807);
or U2223 (N_2223,N_1995,N_1879);
nor U2224 (N_2224,N_1995,N_1935);
and U2225 (N_2225,N_1964,N_1983);
and U2226 (N_2226,N_1824,N_1765);
xor U2227 (N_2227,N_1969,N_1939);
or U2228 (N_2228,N_1895,N_1972);
and U2229 (N_2229,N_1978,N_1812);
nand U2230 (N_2230,N_1943,N_1930);
and U2231 (N_2231,N_1922,N_1950);
nand U2232 (N_2232,N_1929,N_1867);
nor U2233 (N_2233,N_1933,N_1905);
nor U2234 (N_2234,N_1950,N_1854);
or U2235 (N_2235,N_1897,N_1995);
and U2236 (N_2236,N_1885,N_1902);
nor U2237 (N_2237,N_1888,N_1825);
nor U2238 (N_2238,N_1795,N_1982);
and U2239 (N_2239,N_1934,N_1999);
nand U2240 (N_2240,N_1945,N_1933);
and U2241 (N_2241,N_1906,N_1841);
nor U2242 (N_2242,N_1953,N_1972);
xnor U2243 (N_2243,N_1910,N_1846);
and U2244 (N_2244,N_1883,N_1828);
or U2245 (N_2245,N_1988,N_1765);
nand U2246 (N_2246,N_1770,N_1884);
and U2247 (N_2247,N_1911,N_1750);
and U2248 (N_2248,N_1885,N_1992);
or U2249 (N_2249,N_1988,N_1822);
or U2250 (N_2250,N_2152,N_2073);
nand U2251 (N_2251,N_2081,N_2174);
nor U2252 (N_2252,N_2013,N_2211);
nor U2253 (N_2253,N_2091,N_2237);
nor U2254 (N_2254,N_2228,N_2162);
and U2255 (N_2255,N_2136,N_2017);
and U2256 (N_2256,N_2012,N_2109);
or U2257 (N_2257,N_2210,N_2236);
or U2258 (N_2258,N_2242,N_2238);
nand U2259 (N_2259,N_2239,N_2010);
nor U2260 (N_2260,N_2104,N_2035);
and U2261 (N_2261,N_2085,N_2209);
nor U2262 (N_2262,N_2173,N_2131);
and U2263 (N_2263,N_2002,N_2096);
and U2264 (N_2264,N_2037,N_2023);
or U2265 (N_2265,N_2086,N_2044);
xor U2266 (N_2266,N_2189,N_2093);
nor U2267 (N_2267,N_2186,N_2125);
or U2268 (N_2268,N_2166,N_2171);
xnor U2269 (N_2269,N_2099,N_2215);
and U2270 (N_2270,N_2089,N_2062);
nor U2271 (N_2271,N_2103,N_2151);
nor U2272 (N_2272,N_2119,N_2076);
nor U2273 (N_2273,N_2144,N_2146);
nor U2274 (N_2274,N_2030,N_2059);
or U2275 (N_2275,N_2056,N_2153);
nor U2276 (N_2276,N_2090,N_2080);
nor U2277 (N_2277,N_2155,N_2219);
nand U2278 (N_2278,N_2129,N_2118);
and U2279 (N_2279,N_2208,N_2034);
or U2280 (N_2280,N_2001,N_2018);
nand U2281 (N_2281,N_2248,N_2177);
and U2282 (N_2282,N_2126,N_2184);
nor U2283 (N_2283,N_2112,N_2038);
or U2284 (N_2284,N_2054,N_2050);
or U2285 (N_2285,N_2247,N_2102);
or U2286 (N_2286,N_2212,N_2113);
nand U2287 (N_2287,N_2156,N_2074);
or U2288 (N_2288,N_2019,N_2180);
or U2289 (N_2289,N_2154,N_2198);
or U2290 (N_2290,N_2231,N_2217);
nand U2291 (N_2291,N_2032,N_2027);
nand U2292 (N_2292,N_2048,N_2135);
and U2293 (N_2293,N_2088,N_2222);
nor U2294 (N_2294,N_2123,N_2213);
and U2295 (N_2295,N_2058,N_2133);
or U2296 (N_2296,N_2064,N_2087);
nand U2297 (N_2297,N_2061,N_2092);
nand U2298 (N_2298,N_2235,N_2043);
or U2299 (N_2299,N_2097,N_2006);
or U2300 (N_2300,N_2063,N_2070);
xor U2301 (N_2301,N_2114,N_2117);
or U2302 (N_2302,N_2022,N_2132);
nand U2303 (N_2303,N_2069,N_2004);
nand U2304 (N_2304,N_2115,N_2082);
xnor U2305 (N_2305,N_2026,N_2221);
nand U2306 (N_2306,N_2077,N_2163);
nand U2307 (N_2307,N_2137,N_2127);
nor U2308 (N_2308,N_2128,N_2033);
and U2309 (N_2309,N_2003,N_2158);
and U2310 (N_2310,N_2078,N_2047);
xnor U2311 (N_2311,N_2145,N_2108);
xnor U2312 (N_2312,N_2110,N_2071);
and U2313 (N_2313,N_2233,N_2200);
or U2314 (N_2314,N_2224,N_2192);
nor U2315 (N_2315,N_2182,N_2005);
and U2316 (N_2316,N_2230,N_2055);
or U2317 (N_2317,N_2201,N_2101);
and U2318 (N_2318,N_2220,N_2130);
nor U2319 (N_2319,N_2160,N_2246);
xor U2320 (N_2320,N_2095,N_2020);
or U2321 (N_2321,N_2169,N_2147);
nand U2322 (N_2322,N_2046,N_2111);
nor U2323 (N_2323,N_2040,N_2203);
nor U2324 (N_2324,N_2134,N_2140);
nor U2325 (N_2325,N_2249,N_2143);
nand U2326 (N_2326,N_2083,N_2161);
or U2327 (N_2327,N_2051,N_2036);
or U2328 (N_2328,N_2185,N_2214);
nor U2329 (N_2329,N_2165,N_2207);
nor U2330 (N_2330,N_2011,N_2183);
nand U2331 (N_2331,N_2194,N_2164);
nand U2332 (N_2332,N_2138,N_2039);
nand U2333 (N_2333,N_2124,N_2049);
and U2334 (N_2334,N_2148,N_2052);
nor U2335 (N_2335,N_2016,N_2045);
xnor U2336 (N_2336,N_2014,N_2168);
xnor U2337 (N_2337,N_2170,N_2084);
xor U2338 (N_2338,N_2150,N_2245);
and U2339 (N_2339,N_2065,N_2015);
and U2340 (N_2340,N_2100,N_2167);
or U2341 (N_2341,N_2141,N_2218);
and U2342 (N_2342,N_2009,N_2157);
nand U2343 (N_2343,N_2031,N_2240);
xnor U2344 (N_2344,N_2204,N_2116);
nor U2345 (N_2345,N_2067,N_2243);
and U2346 (N_2346,N_2206,N_2178);
nor U2347 (N_2347,N_2190,N_2007);
or U2348 (N_2348,N_2199,N_2205);
and U2349 (N_2349,N_2191,N_2008);
nand U2350 (N_2350,N_2120,N_2028);
or U2351 (N_2351,N_2042,N_2176);
and U2352 (N_2352,N_2029,N_2232);
and U2353 (N_2353,N_2227,N_2041);
nand U2354 (N_2354,N_2244,N_2021);
nor U2355 (N_2355,N_2106,N_2060);
nor U2356 (N_2356,N_2195,N_2181);
and U2357 (N_2357,N_2197,N_2229);
nand U2358 (N_2358,N_2053,N_2068);
nand U2359 (N_2359,N_2188,N_2098);
or U2360 (N_2360,N_2225,N_2066);
xor U2361 (N_2361,N_2179,N_2142);
or U2362 (N_2362,N_2079,N_2025);
xor U2363 (N_2363,N_2187,N_2094);
nand U2364 (N_2364,N_2216,N_2196);
or U2365 (N_2365,N_2202,N_2226);
or U2366 (N_2366,N_2000,N_2159);
or U2367 (N_2367,N_2075,N_2241);
nand U2368 (N_2368,N_2149,N_2234);
nor U2369 (N_2369,N_2105,N_2107);
and U2370 (N_2370,N_2172,N_2072);
and U2371 (N_2371,N_2139,N_2223);
nor U2372 (N_2372,N_2122,N_2175);
or U2373 (N_2373,N_2057,N_2024);
xor U2374 (N_2374,N_2121,N_2193);
or U2375 (N_2375,N_2091,N_2187);
nor U2376 (N_2376,N_2025,N_2059);
and U2377 (N_2377,N_2155,N_2019);
nor U2378 (N_2378,N_2101,N_2089);
or U2379 (N_2379,N_2039,N_2071);
or U2380 (N_2380,N_2238,N_2209);
or U2381 (N_2381,N_2030,N_2097);
or U2382 (N_2382,N_2093,N_2117);
nor U2383 (N_2383,N_2215,N_2092);
and U2384 (N_2384,N_2197,N_2073);
nand U2385 (N_2385,N_2077,N_2168);
or U2386 (N_2386,N_2026,N_2147);
xnor U2387 (N_2387,N_2132,N_2155);
nand U2388 (N_2388,N_2012,N_2054);
nor U2389 (N_2389,N_2232,N_2151);
nor U2390 (N_2390,N_2230,N_2022);
or U2391 (N_2391,N_2111,N_2229);
nand U2392 (N_2392,N_2118,N_2237);
nand U2393 (N_2393,N_2057,N_2135);
and U2394 (N_2394,N_2181,N_2084);
nand U2395 (N_2395,N_2022,N_2069);
xnor U2396 (N_2396,N_2115,N_2182);
and U2397 (N_2397,N_2094,N_2227);
and U2398 (N_2398,N_2047,N_2110);
and U2399 (N_2399,N_2111,N_2233);
or U2400 (N_2400,N_2210,N_2161);
and U2401 (N_2401,N_2246,N_2167);
and U2402 (N_2402,N_2146,N_2081);
or U2403 (N_2403,N_2133,N_2165);
xor U2404 (N_2404,N_2239,N_2220);
xnor U2405 (N_2405,N_2125,N_2054);
and U2406 (N_2406,N_2173,N_2089);
nand U2407 (N_2407,N_2144,N_2249);
xor U2408 (N_2408,N_2192,N_2155);
nand U2409 (N_2409,N_2093,N_2107);
or U2410 (N_2410,N_2026,N_2241);
and U2411 (N_2411,N_2038,N_2113);
nor U2412 (N_2412,N_2242,N_2207);
and U2413 (N_2413,N_2124,N_2178);
and U2414 (N_2414,N_2099,N_2041);
and U2415 (N_2415,N_2112,N_2066);
and U2416 (N_2416,N_2168,N_2248);
nand U2417 (N_2417,N_2229,N_2004);
nand U2418 (N_2418,N_2077,N_2060);
nor U2419 (N_2419,N_2001,N_2098);
and U2420 (N_2420,N_2236,N_2049);
xor U2421 (N_2421,N_2213,N_2085);
nand U2422 (N_2422,N_2167,N_2127);
or U2423 (N_2423,N_2099,N_2167);
nor U2424 (N_2424,N_2226,N_2170);
or U2425 (N_2425,N_2064,N_2048);
nand U2426 (N_2426,N_2020,N_2072);
and U2427 (N_2427,N_2223,N_2236);
and U2428 (N_2428,N_2041,N_2178);
or U2429 (N_2429,N_2142,N_2177);
or U2430 (N_2430,N_2119,N_2224);
nand U2431 (N_2431,N_2022,N_2249);
xor U2432 (N_2432,N_2133,N_2203);
xnor U2433 (N_2433,N_2097,N_2159);
and U2434 (N_2434,N_2079,N_2089);
and U2435 (N_2435,N_2236,N_2077);
nor U2436 (N_2436,N_2150,N_2120);
nand U2437 (N_2437,N_2113,N_2201);
nor U2438 (N_2438,N_2138,N_2163);
or U2439 (N_2439,N_2075,N_2214);
and U2440 (N_2440,N_2080,N_2107);
nand U2441 (N_2441,N_2240,N_2204);
xor U2442 (N_2442,N_2068,N_2088);
or U2443 (N_2443,N_2105,N_2097);
and U2444 (N_2444,N_2223,N_2237);
and U2445 (N_2445,N_2086,N_2195);
xor U2446 (N_2446,N_2133,N_2102);
nor U2447 (N_2447,N_2009,N_2228);
nand U2448 (N_2448,N_2178,N_2031);
nor U2449 (N_2449,N_2146,N_2060);
or U2450 (N_2450,N_2227,N_2065);
or U2451 (N_2451,N_2033,N_2182);
nor U2452 (N_2452,N_2116,N_2054);
nand U2453 (N_2453,N_2041,N_2225);
or U2454 (N_2454,N_2211,N_2097);
nor U2455 (N_2455,N_2160,N_2121);
xor U2456 (N_2456,N_2110,N_2134);
and U2457 (N_2457,N_2143,N_2090);
or U2458 (N_2458,N_2242,N_2206);
or U2459 (N_2459,N_2044,N_2093);
or U2460 (N_2460,N_2051,N_2187);
nor U2461 (N_2461,N_2073,N_2133);
and U2462 (N_2462,N_2030,N_2094);
nor U2463 (N_2463,N_2246,N_2060);
nand U2464 (N_2464,N_2106,N_2215);
nor U2465 (N_2465,N_2238,N_2026);
and U2466 (N_2466,N_2209,N_2001);
and U2467 (N_2467,N_2020,N_2200);
nand U2468 (N_2468,N_2189,N_2128);
nand U2469 (N_2469,N_2224,N_2189);
nand U2470 (N_2470,N_2188,N_2215);
xor U2471 (N_2471,N_2087,N_2201);
and U2472 (N_2472,N_2075,N_2246);
and U2473 (N_2473,N_2244,N_2243);
and U2474 (N_2474,N_2002,N_2008);
nor U2475 (N_2475,N_2130,N_2215);
or U2476 (N_2476,N_2126,N_2105);
and U2477 (N_2477,N_2042,N_2223);
nor U2478 (N_2478,N_2145,N_2189);
nand U2479 (N_2479,N_2148,N_2127);
xor U2480 (N_2480,N_2157,N_2004);
or U2481 (N_2481,N_2148,N_2211);
or U2482 (N_2482,N_2051,N_2094);
xor U2483 (N_2483,N_2195,N_2025);
nand U2484 (N_2484,N_2157,N_2023);
or U2485 (N_2485,N_2248,N_2167);
nor U2486 (N_2486,N_2154,N_2211);
nor U2487 (N_2487,N_2143,N_2165);
nand U2488 (N_2488,N_2092,N_2076);
and U2489 (N_2489,N_2131,N_2062);
nor U2490 (N_2490,N_2061,N_2057);
xor U2491 (N_2491,N_2011,N_2211);
nor U2492 (N_2492,N_2098,N_2215);
nor U2493 (N_2493,N_2167,N_2188);
and U2494 (N_2494,N_2225,N_2199);
or U2495 (N_2495,N_2054,N_2238);
or U2496 (N_2496,N_2225,N_2111);
or U2497 (N_2497,N_2080,N_2196);
nor U2498 (N_2498,N_2237,N_2039);
or U2499 (N_2499,N_2172,N_2156);
xnor U2500 (N_2500,N_2472,N_2311);
or U2501 (N_2501,N_2275,N_2367);
nand U2502 (N_2502,N_2491,N_2328);
nand U2503 (N_2503,N_2404,N_2264);
nand U2504 (N_2504,N_2457,N_2292);
and U2505 (N_2505,N_2305,N_2389);
and U2506 (N_2506,N_2450,N_2485);
and U2507 (N_2507,N_2296,N_2459);
or U2508 (N_2508,N_2256,N_2252);
nor U2509 (N_2509,N_2384,N_2463);
or U2510 (N_2510,N_2373,N_2496);
or U2511 (N_2511,N_2345,N_2475);
nand U2512 (N_2512,N_2458,N_2383);
or U2513 (N_2513,N_2417,N_2385);
nor U2514 (N_2514,N_2461,N_2453);
xor U2515 (N_2515,N_2494,N_2375);
and U2516 (N_2516,N_2312,N_2327);
and U2517 (N_2517,N_2456,N_2486);
nand U2518 (N_2518,N_2452,N_2393);
and U2519 (N_2519,N_2271,N_2396);
nor U2520 (N_2520,N_2445,N_2407);
xnor U2521 (N_2521,N_2350,N_2257);
nand U2522 (N_2522,N_2465,N_2480);
nand U2523 (N_2523,N_2451,N_2278);
and U2524 (N_2524,N_2388,N_2268);
nand U2525 (N_2525,N_2467,N_2354);
nor U2526 (N_2526,N_2267,N_2443);
or U2527 (N_2527,N_2430,N_2444);
nand U2528 (N_2528,N_2338,N_2374);
nand U2529 (N_2529,N_2322,N_2454);
or U2530 (N_2530,N_2497,N_2253);
nand U2531 (N_2531,N_2413,N_2394);
nor U2532 (N_2532,N_2474,N_2390);
and U2533 (N_2533,N_2318,N_2325);
and U2534 (N_2534,N_2351,N_2326);
nor U2535 (N_2535,N_2381,N_2462);
or U2536 (N_2536,N_2477,N_2418);
xnor U2537 (N_2537,N_2449,N_2287);
or U2538 (N_2538,N_2265,N_2419);
or U2539 (N_2539,N_2498,N_2464);
or U2540 (N_2540,N_2358,N_2258);
or U2541 (N_2541,N_2291,N_2364);
and U2542 (N_2542,N_2282,N_2307);
nand U2543 (N_2543,N_2435,N_2378);
nand U2544 (N_2544,N_2355,N_2340);
nand U2545 (N_2545,N_2481,N_2290);
and U2546 (N_2546,N_2269,N_2308);
and U2547 (N_2547,N_2370,N_2335);
nand U2548 (N_2548,N_2427,N_2360);
nor U2549 (N_2549,N_2425,N_2423);
and U2550 (N_2550,N_2493,N_2377);
xor U2551 (N_2551,N_2402,N_2330);
or U2552 (N_2552,N_2342,N_2420);
or U2553 (N_2553,N_2470,N_2428);
or U2554 (N_2554,N_2403,N_2429);
nand U2555 (N_2555,N_2436,N_2277);
and U2556 (N_2556,N_2380,N_2460);
or U2557 (N_2557,N_2295,N_2487);
nor U2558 (N_2558,N_2424,N_2365);
nor U2559 (N_2559,N_2489,N_2441);
nor U2560 (N_2560,N_2431,N_2434);
nand U2561 (N_2561,N_2426,N_2309);
nand U2562 (N_2562,N_2280,N_2484);
and U2563 (N_2563,N_2276,N_2310);
nand U2564 (N_2564,N_2259,N_2398);
nand U2565 (N_2565,N_2333,N_2408);
xnor U2566 (N_2566,N_2397,N_2255);
nor U2567 (N_2567,N_2285,N_2409);
nand U2568 (N_2568,N_2324,N_2303);
and U2569 (N_2569,N_2414,N_2415);
nand U2570 (N_2570,N_2349,N_2306);
or U2571 (N_2571,N_2416,N_2321);
nand U2572 (N_2572,N_2437,N_2371);
xor U2573 (N_2573,N_2284,N_2438);
nor U2574 (N_2574,N_2392,N_2395);
nor U2575 (N_2575,N_2356,N_2298);
nor U2576 (N_2576,N_2283,N_2313);
or U2577 (N_2577,N_2254,N_2293);
nand U2578 (N_2578,N_2379,N_2359);
nor U2579 (N_2579,N_2368,N_2301);
or U2580 (N_2580,N_2270,N_2251);
xor U2581 (N_2581,N_2369,N_2250);
xor U2582 (N_2582,N_2446,N_2422);
xor U2583 (N_2583,N_2387,N_2319);
xnor U2584 (N_2584,N_2421,N_2316);
or U2585 (N_2585,N_2412,N_2299);
and U2586 (N_2586,N_2286,N_2279);
xnor U2587 (N_2587,N_2410,N_2447);
and U2588 (N_2588,N_2372,N_2439);
nor U2589 (N_2589,N_2432,N_2346);
and U2590 (N_2590,N_2281,N_2341);
nand U2591 (N_2591,N_2411,N_2482);
and U2592 (N_2592,N_2288,N_2334);
and U2593 (N_2593,N_2323,N_2440);
nand U2594 (N_2594,N_2260,N_2405);
nor U2595 (N_2595,N_2337,N_2391);
and U2596 (N_2596,N_2483,N_2336);
or U2597 (N_2597,N_2320,N_2304);
and U2598 (N_2598,N_2348,N_2471);
and U2599 (N_2599,N_2294,N_2315);
nor U2600 (N_2600,N_2400,N_2478);
nor U2601 (N_2601,N_2363,N_2386);
nor U2602 (N_2602,N_2332,N_2466);
xnor U2603 (N_2603,N_2317,N_2455);
and U2604 (N_2604,N_2476,N_2469);
or U2605 (N_2605,N_2399,N_2473);
or U2606 (N_2606,N_2366,N_2344);
nand U2607 (N_2607,N_2261,N_2263);
or U2608 (N_2608,N_2361,N_2274);
or U2609 (N_2609,N_2401,N_2266);
or U2610 (N_2610,N_2488,N_2499);
and U2611 (N_2611,N_2448,N_2289);
and U2612 (N_2612,N_2329,N_2357);
nand U2613 (N_2613,N_2376,N_2262);
and U2614 (N_2614,N_2442,N_2406);
and U2615 (N_2615,N_2492,N_2352);
xor U2616 (N_2616,N_2314,N_2297);
xnor U2617 (N_2617,N_2468,N_2353);
and U2618 (N_2618,N_2302,N_2300);
nor U2619 (N_2619,N_2433,N_2479);
and U2620 (N_2620,N_2490,N_2495);
and U2621 (N_2621,N_2331,N_2339);
and U2622 (N_2622,N_2362,N_2343);
and U2623 (N_2623,N_2382,N_2272);
and U2624 (N_2624,N_2273,N_2347);
nor U2625 (N_2625,N_2361,N_2334);
or U2626 (N_2626,N_2297,N_2402);
or U2627 (N_2627,N_2272,N_2330);
nor U2628 (N_2628,N_2314,N_2483);
and U2629 (N_2629,N_2364,N_2326);
nand U2630 (N_2630,N_2343,N_2452);
or U2631 (N_2631,N_2456,N_2492);
and U2632 (N_2632,N_2356,N_2325);
nor U2633 (N_2633,N_2473,N_2481);
xnor U2634 (N_2634,N_2451,N_2474);
nor U2635 (N_2635,N_2418,N_2293);
nand U2636 (N_2636,N_2274,N_2260);
nor U2637 (N_2637,N_2393,N_2353);
nor U2638 (N_2638,N_2259,N_2418);
nor U2639 (N_2639,N_2465,N_2261);
nand U2640 (N_2640,N_2389,N_2332);
or U2641 (N_2641,N_2494,N_2276);
or U2642 (N_2642,N_2363,N_2429);
or U2643 (N_2643,N_2281,N_2327);
or U2644 (N_2644,N_2479,N_2476);
nand U2645 (N_2645,N_2377,N_2253);
and U2646 (N_2646,N_2325,N_2352);
nand U2647 (N_2647,N_2297,N_2281);
nor U2648 (N_2648,N_2350,N_2456);
xnor U2649 (N_2649,N_2299,N_2341);
xor U2650 (N_2650,N_2319,N_2405);
or U2651 (N_2651,N_2466,N_2302);
nor U2652 (N_2652,N_2382,N_2285);
and U2653 (N_2653,N_2364,N_2419);
xor U2654 (N_2654,N_2400,N_2454);
and U2655 (N_2655,N_2282,N_2333);
or U2656 (N_2656,N_2301,N_2466);
nor U2657 (N_2657,N_2422,N_2313);
nand U2658 (N_2658,N_2471,N_2488);
nor U2659 (N_2659,N_2488,N_2411);
nor U2660 (N_2660,N_2381,N_2299);
nand U2661 (N_2661,N_2478,N_2374);
and U2662 (N_2662,N_2343,N_2498);
or U2663 (N_2663,N_2321,N_2477);
nor U2664 (N_2664,N_2250,N_2396);
and U2665 (N_2665,N_2346,N_2469);
or U2666 (N_2666,N_2257,N_2343);
nor U2667 (N_2667,N_2425,N_2488);
or U2668 (N_2668,N_2322,N_2330);
nor U2669 (N_2669,N_2456,N_2301);
nor U2670 (N_2670,N_2405,N_2442);
and U2671 (N_2671,N_2379,N_2290);
nor U2672 (N_2672,N_2496,N_2342);
and U2673 (N_2673,N_2486,N_2368);
nand U2674 (N_2674,N_2398,N_2270);
or U2675 (N_2675,N_2478,N_2277);
nand U2676 (N_2676,N_2430,N_2438);
nor U2677 (N_2677,N_2367,N_2482);
nor U2678 (N_2678,N_2403,N_2260);
or U2679 (N_2679,N_2332,N_2290);
nor U2680 (N_2680,N_2264,N_2256);
or U2681 (N_2681,N_2270,N_2289);
nor U2682 (N_2682,N_2339,N_2381);
nor U2683 (N_2683,N_2272,N_2314);
nand U2684 (N_2684,N_2259,N_2281);
nor U2685 (N_2685,N_2325,N_2254);
xor U2686 (N_2686,N_2308,N_2280);
or U2687 (N_2687,N_2345,N_2287);
or U2688 (N_2688,N_2310,N_2326);
or U2689 (N_2689,N_2499,N_2259);
xnor U2690 (N_2690,N_2456,N_2337);
or U2691 (N_2691,N_2294,N_2379);
nand U2692 (N_2692,N_2408,N_2270);
nor U2693 (N_2693,N_2256,N_2364);
and U2694 (N_2694,N_2281,N_2353);
nor U2695 (N_2695,N_2369,N_2370);
xor U2696 (N_2696,N_2366,N_2393);
and U2697 (N_2697,N_2415,N_2321);
and U2698 (N_2698,N_2255,N_2360);
xor U2699 (N_2699,N_2480,N_2430);
or U2700 (N_2700,N_2441,N_2432);
and U2701 (N_2701,N_2289,N_2345);
and U2702 (N_2702,N_2494,N_2481);
nor U2703 (N_2703,N_2394,N_2306);
nor U2704 (N_2704,N_2303,N_2481);
nand U2705 (N_2705,N_2285,N_2256);
or U2706 (N_2706,N_2350,N_2273);
nand U2707 (N_2707,N_2458,N_2286);
or U2708 (N_2708,N_2332,N_2451);
nor U2709 (N_2709,N_2446,N_2431);
nor U2710 (N_2710,N_2422,N_2271);
nor U2711 (N_2711,N_2468,N_2314);
nor U2712 (N_2712,N_2473,N_2293);
xnor U2713 (N_2713,N_2388,N_2291);
nand U2714 (N_2714,N_2421,N_2434);
nand U2715 (N_2715,N_2372,N_2273);
and U2716 (N_2716,N_2412,N_2418);
or U2717 (N_2717,N_2334,N_2392);
nand U2718 (N_2718,N_2376,N_2450);
or U2719 (N_2719,N_2419,N_2460);
nor U2720 (N_2720,N_2435,N_2262);
nand U2721 (N_2721,N_2480,N_2289);
nor U2722 (N_2722,N_2310,N_2268);
or U2723 (N_2723,N_2440,N_2489);
nand U2724 (N_2724,N_2459,N_2455);
nand U2725 (N_2725,N_2261,N_2324);
xnor U2726 (N_2726,N_2283,N_2344);
or U2727 (N_2727,N_2459,N_2354);
or U2728 (N_2728,N_2281,N_2398);
nor U2729 (N_2729,N_2270,N_2414);
nand U2730 (N_2730,N_2339,N_2484);
and U2731 (N_2731,N_2283,N_2342);
and U2732 (N_2732,N_2450,N_2325);
and U2733 (N_2733,N_2267,N_2263);
or U2734 (N_2734,N_2390,N_2431);
and U2735 (N_2735,N_2264,N_2421);
nand U2736 (N_2736,N_2288,N_2402);
and U2737 (N_2737,N_2393,N_2438);
or U2738 (N_2738,N_2351,N_2406);
and U2739 (N_2739,N_2333,N_2393);
nand U2740 (N_2740,N_2358,N_2484);
and U2741 (N_2741,N_2400,N_2489);
nor U2742 (N_2742,N_2472,N_2439);
and U2743 (N_2743,N_2298,N_2339);
nor U2744 (N_2744,N_2498,N_2295);
nor U2745 (N_2745,N_2372,N_2298);
nor U2746 (N_2746,N_2395,N_2334);
or U2747 (N_2747,N_2363,N_2456);
nand U2748 (N_2748,N_2379,N_2430);
or U2749 (N_2749,N_2253,N_2273);
nand U2750 (N_2750,N_2721,N_2702);
xnor U2751 (N_2751,N_2588,N_2616);
nand U2752 (N_2752,N_2723,N_2509);
and U2753 (N_2753,N_2724,N_2615);
and U2754 (N_2754,N_2583,N_2548);
nor U2755 (N_2755,N_2729,N_2526);
nor U2756 (N_2756,N_2672,N_2574);
nor U2757 (N_2757,N_2551,N_2715);
and U2758 (N_2758,N_2695,N_2680);
and U2759 (N_2759,N_2567,N_2537);
nand U2760 (N_2760,N_2611,N_2656);
nor U2761 (N_2761,N_2601,N_2618);
nor U2762 (N_2762,N_2722,N_2595);
and U2763 (N_2763,N_2538,N_2740);
xor U2764 (N_2764,N_2657,N_2590);
nor U2765 (N_2765,N_2637,N_2536);
xnor U2766 (N_2766,N_2597,N_2596);
nor U2767 (N_2767,N_2599,N_2564);
nor U2768 (N_2768,N_2562,N_2727);
and U2769 (N_2769,N_2553,N_2534);
nor U2770 (N_2770,N_2510,N_2710);
nor U2771 (N_2771,N_2593,N_2560);
and U2772 (N_2772,N_2716,N_2687);
xnor U2773 (N_2773,N_2576,N_2508);
nor U2774 (N_2774,N_2500,N_2513);
nand U2775 (N_2775,N_2625,N_2559);
nand U2776 (N_2776,N_2706,N_2745);
and U2777 (N_2777,N_2717,N_2686);
nand U2778 (N_2778,N_2524,N_2688);
nor U2779 (N_2779,N_2623,N_2598);
nor U2780 (N_2780,N_2654,N_2644);
nor U2781 (N_2781,N_2643,N_2628);
xor U2782 (N_2782,N_2572,N_2698);
or U2783 (N_2783,N_2659,N_2569);
nand U2784 (N_2784,N_2684,N_2676);
nand U2785 (N_2785,N_2501,N_2591);
or U2786 (N_2786,N_2606,N_2674);
or U2787 (N_2787,N_2507,N_2622);
and U2788 (N_2788,N_2518,N_2638);
nor U2789 (N_2789,N_2681,N_2587);
nand U2790 (N_2790,N_2580,N_2520);
and U2791 (N_2791,N_2707,N_2734);
and U2792 (N_2792,N_2713,N_2645);
nor U2793 (N_2793,N_2529,N_2581);
or U2794 (N_2794,N_2696,N_2749);
nand U2795 (N_2795,N_2530,N_2515);
nor U2796 (N_2796,N_2624,N_2699);
nand U2797 (N_2797,N_2570,N_2585);
or U2798 (N_2798,N_2555,N_2741);
or U2799 (N_2799,N_2661,N_2641);
or U2800 (N_2800,N_2631,N_2691);
nand U2801 (N_2801,N_2739,N_2711);
nor U2802 (N_2802,N_2636,N_2610);
nor U2803 (N_2803,N_2511,N_2655);
nand U2804 (N_2804,N_2709,N_2700);
nor U2805 (N_2805,N_2516,N_2635);
nor U2806 (N_2806,N_2626,N_2602);
xor U2807 (N_2807,N_2658,N_2621);
nand U2808 (N_2808,N_2682,N_2603);
or U2809 (N_2809,N_2693,N_2646);
and U2810 (N_2810,N_2665,N_2629);
nand U2811 (N_2811,N_2728,N_2650);
and U2812 (N_2812,N_2521,N_2666);
nand U2813 (N_2813,N_2527,N_2748);
and U2814 (N_2814,N_2642,N_2539);
nor U2815 (N_2815,N_2719,N_2725);
nand U2816 (N_2816,N_2514,N_2565);
and U2817 (N_2817,N_2605,N_2664);
nand U2818 (N_2818,N_2578,N_2546);
nand U2819 (N_2819,N_2523,N_2726);
nand U2820 (N_2820,N_2543,N_2549);
nor U2821 (N_2821,N_2633,N_2732);
nor U2822 (N_2822,N_2502,N_2525);
nor U2823 (N_2823,N_2685,N_2697);
nand U2824 (N_2824,N_2568,N_2608);
nor U2825 (N_2825,N_2573,N_2705);
or U2826 (N_2826,N_2594,N_2584);
xor U2827 (N_2827,N_2662,N_2663);
nor U2828 (N_2828,N_2531,N_2577);
or U2829 (N_2829,N_2694,N_2604);
nor U2830 (N_2830,N_2586,N_2634);
or U2831 (N_2831,N_2517,N_2667);
nand U2832 (N_2832,N_2701,N_2651);
and U2833 (N_2833,N_2600,N_2630);
nor U2834 (N_2834,N_2545,N_2718);
or U2835 (N_2835,N_2566,N_2532);
or U2836 (N_2836,N_2708,N_2668);
or U2837 (N_2837,N_2746,N_2535);
nand U2838 (N_2838,N_2689,N_2678);
and U2839 (N_2839,N_2519,N_2714);
or U2840 (N_2840,N_2743,N_2649);
and U2841 (N_2841,N_2677,N_2670);
nand U2842 (N_2842,N_2554,N_2541);
nand U2843 (N_2843,N_2561,N_2544);
nor U2844 (N_2844,N_2614,N_2582);
and U2845 (N_2845,N_2730,N_2557);
and U2846 (N_2846,N_2575,N_2742);
xor U2847 (N_2847,N_2669,N_2550);
nor U2848 (N_2848,N_2613,N_2653);
and U2849 (N_2849,N_2528,N_2503);
nand U2850 (N_2850,N_2505,N_2736);
nor U2851 (N_2851,N_2617,N_2571);
and U2852 (N_2852,N_2720,N_2673);
nor U2853 (N_2853,N_2556,N_2640);
nor U2854 (N_2854,N_2737,N_2639);
or U2855 (N_2855,N_2683,N_2632);
and U2856 (N_2856,N_2533,N_2506);
and U2857 (N_2857,N_2619,N_2675);
nor U2858 (N_2858,N_2660,N_2542);
or U2859 (N_2859,N_2522,N_2609);
nor U2860 (N_2860,N_2731,N_2671);
nand U2861 (N_2861,N_2704,N_2703);
nor U2862 (N_2862,N_2744,N_2627);
nor U2863 (N_2863,N_2563,N_2733);
xor U2864 (N_2864,N_2679,N_2552);
or U2865 (N_2865,N_2547,N_2512);
nor U2866 (N_2866,N_2692,N_2647);
xor U2867 (N_2867,N_2712,N_2747);
or U2868 (N_2868,N_2589,N_2690);
nor U2869 (N_2869,N_2592,N_2620);
nor U2870 (N_2870,N_2735,N_2558);
nor U2871 (N_2871,N_2540,N_2504);
nand U2872 (N_2872,N_2652,N_2738);
and U2873 (N_2873,N_2648,N_2579);
or U2874 (N_2874,N_2612,N_2607);
or U2875 (N_2875,N_2722,N_2737);
and U2876 (N_2876,N_2617,N_2621);
nand U2877 (N_2877,N_2593,N_2645);
nor U2878 (N_2878,N_2505,N_2592);
and U2879 (N_2879,N_2637,N_2741);
and U2880 (N_2880,N_2504,N_2635);
and U2881 (N_2881,N_2668,N_2621);
or U2882 (N_2882,N_2556,N_2550);
or U2883 (N_2883,N_2505,N_2588);
and U2884 (N_2884,N_2729,N_2734);
xor U2885 (N_2885,N_2710,N_2667);
or U2886 (N_2886,N_2555,N_2739);
or U2887 (N_2887,N_2560,N_2548);
or U2888 (N_2888,N_2697,N_2739);
nand U2889 (N_2889,N_2621,N_2727);
nand U2890 (N_2890,N_2586,N_2576);
and U2891 (N_2891,N_2513,N_2612);
nand U2892 (N_2892,N_2539,N_2689);
nor U2893 (N_2893,N_2643,N_2679);
and U2894 (N_2894,N_2672,N_2584);
and U2895 (N_2895,N_2658,N_2719);
nor U2896 (N_2896,N_2682,N_2680);
xor U2897 (N_2897,N_2533,N_2593);
and U2898 (N_2898,N_2520,N_2533);
nor U2899 (N_2899,N_2581,N_2559);
nand U2900 (N_2900,N_2544,N_2567);
and U2901 (N_2901,N_2559,N_2538);
and U2902 (N_2902,N_2565,N_2673);
or U2903 (N_2903,N_2519,N_2663);
xnor U2904 (N_2904,N_2634,N_2744);
and U2905 (N_2905,N_2505,N_2644);
or U2906 (N_2906,N_2622,N_2602);
xnor U2907 (N_2907,N_2605,N_2745);
or U2908 (N_2908,N_2706,N_2505);
xnor U2909 (N_2909,N_2671,N_2574);
nor U2910 (N_2910,N_2543,N_2627);
xnor U2911 (N_2911,N_2500,N_2613);
nand U2912 (N_2912,N_2698,N_2719);
or U2913 (N_2913,N_2540,N_2517);
and U2914 (N_2914,N_2654,N_2609);
nand U2915 (N_2915,N_2557,N_2537);
nand U2916 (N_2916,N_2506,N_2548);
or U2917 (N_2917,N_2662,N_2597);
nor U2918 (N_2918,N_2504,N_2719);
nand U2919 (N_2919,N_2730,N_2540);
nor U2920 (N_2920,N_2663,N_2547);
or U2921 (N_2921,N_2581,N_2653);
and U2922 (N_2922,N_2560,N_2654);
nor U2923 (N_2923,N_2672,N_2623);
nor U2924 (N_2924,N_2685,N_2601);
and U2925 (N_2925,N_2709,N_2503);
or U2926 (N_2926,N_2742,N_2548);
and U2927 (N_2927,N_2713,N_2530);
nor U2928 (N_2928,N_2645,N_2559);
nor U2929 (N_2929,N_2641,N_2555);
or U2930 (N_2930,N_2737,N_2723);
or U2931 (N_2931,N_2748,N_2568);
xor U2932 (N_2932,N_2523,N_2709);
nor U2933 (N_2933,N_2743,N_2682);
nand U2934 (N_2934,N_2717,N_2705);
and U2935 (N_2935,N_2520,N_2501);
and U2936 (N_2936,N_2705,N_2720);
nor U2937 (N_2937,N_2720,N_2566);
and U2938 (N_2938,N_2556,N_2690);
xor U2939 (N_2939,N_2581,N_2734);
nand U2940 (N_2940,N_2545,N_2603);
nand U2941 (N_2941,N_2705,N_2667);
or U2942 (N_2942,N_2638,N_2643);
nand U2943 (N_2943,N_2688,N_2729);
and U2944 (N_2944,N_2545,N_2536);
or U2945 (N_2945,N_2733,N_2684);
and U2946 (N_2946,N_2503,N_2737);
nand U2947 (N_2947,N_2628,N_2721);
nor U2948 (N_2948,N_2657,N_2503);
nor U2949 (N_2949,N_2540,N_2630);
xor U2950 (N_2950,N_2670,N_2695);
nand U2951 (N_2951,N_2655,N_2521);
nor U2952 (N_2952,N_2727,N_2505);
xnor U2953 (N_2953,N_2692,N_2737);
xnor U2954 (N_2954,N_2621,N_2584);
nand U2955 (N_2955,N_2586,N_2533);
or U2956 (N_2956,N_2669,N_2542);
nand U2957 (N_2957,N_2676,N_2723);
nand U2958 (N_2958,N_2692,N_2564);
and U2959 (N_2959,N_2554,N_2642);
xnor U2960 (N_2960,N_2678,N_2577);
nand U2961 (N_2961,N_2682,N_2602);
xnor U2962 (N_2962,N_2641,N_2671);
nand U2963 (N_2963,N_2674,N_2530);
nor U2964 (N_2964,N_2731,N_2601);
xor U2965 (N_2965,N_2613,N_2718);
xor U2966 (N_2966,N_2510,N_2719);
and U2967 (N_2967,N_2546,N_2506);
and U2968 (N_2968,N_2535,N_2648);
nand U2969 (N_2969,N_2563,N_2555);
nor U2970 (N_2970,N_2724,N_2602);
nand U2971 (N_2971,N_2560,N_2636);
nor U2972 (N_2972,N_2571,N_2650);
xor U2973 (N_2973,N_2508,N_2533);
nor U2974 (N_2974,N_2596,N_2686);
and U2975 (N_2975,N_2552,N_2577);
nor U2976 (N_2976,N_2573,N_2711);
nor U2977 (N_2977,N_2613,N_2738);
and U2978 (N_2978,N_2659,N_2704);
nor U2979 (N_2979,N_2668,N_2670);
nor U2980 (N_2980,N_2502,N_2594);
xor U2981 (N_2981,N_2527,N_2714);
nor U2982 (N_2982,N_2644,N_2727);
xor U2983 (N_2983,N_2692,N_2741);
and U2984 (N_2984,N_2686,N_2742);
and U2985 (N_2985,N_2545,N_2512);
nand U2986 (N_2986,N_2626,N_2650);
nand U2987 (N_2987,N_2531,N_2683);
nor U2988 (N_2988,N_2514,N_2613);
or U2989 (N_2989,N_2564,N_2674);
nand U2990 (N_2990,N_2586,N_2555);
xnor U2991 (N_2991,N_2677,N_2703);
and U2992 (N_2992,N_2667,N_2746);
nor U2993 (N_2993,N_2681,N_2607);
and U2994 (N_2994,N_2657,N_2560);
nor U2995 (N_2995,N_2703,N_2501);
or U2996 (N_2996,N_2565,N_2738);
nor U2997 (N_2997,N_2661,N_2509);
and U2998 (N_2998,N_2671,N_2664);
and U2999 (N_2999,N_2587,N_2646);
and U3000 (N_3000,N_2927,N_2984);
nor U3001 (N_3001,N_2810,N_2892);
xor U3002 (N_3002,N_2960,N_2854);
nand U3003 (N_3003,N_2944,N_2820);
and U3004 (N_3004,N_2968,N_2890);
nand U3005 (N_3005,N_2797,N_2809);
or U3006 (N_3006,N_2818,N_2817);
xnor U3007 (N_3007,N_2763,N_2812);
xnor U3008 (N_3008,N_2974,N_2774);
nor U3009 (N_3009,N_2853,N_2872);
and U3010 (N_3010,N_2967,N_2806);
nor U3011 (N_3011,N_2827,N_2884);
or U3012 (N_3012,N_2837,N_2869);
nand U3013 (N_3013,N_2859,N_2989);
xnor U3014 (N_3014,N_2966,N_2938);
or U3015 (N_3015,N_2945,N_2929);
or U3016 (N_3016,N_2877,N_2808);
or U3017 (N_3017,N_2782,N_2897);
nor U3018 (N_3018,N_2755,N_2780);
nand U3019 (N_3019,N_2828,N_2993);
nor U3020 (N_3020,N_2758,N_2952);
nand U3021 (N_3021,N_2958,N_2916);
and U3022 (N_3022,N_2752,N_2814);
nor U3023 (N_3023,N_2979,N_2992);
nor U3024 (N_3024,N_2868,N_2756);
nor U3025 (N_3025,N_2874,N_2923);
or U3026 (N_3026,N_2829,N_2832);
nor U3027 (N_3027,N_2863,N_2922);
or U3028 (N_3028,N_2838,N_2981);
xor U3029 (N_3029,N_2994,N_2911);
nor U3030 (N_3030,N_2821,N_2865);
nand U3031 (N_3031,N_2835,N_2954);
or U3032 (N_3032,N_2751,N_2856);
nand U3033 (N_3033,N_2824,N_2924);
nor U3034 (N_3034,N_2764,N_2775);
nor U3035 (N_3035,N_2771,N_2910);
or U3036 (N_3036,N_2932,N_2840);
nand U3037 (N_3037,N_2912,N_2772);
and U3038 (N_3038,N_2867,N_2915);
nor U3039 (N_3039,N_2947,N_2861);
nor U3040 (N_3040,N_2843,N_2901);
nand U3041 (N_3041,N_2970,N_2870);
xnor U3042 (N_3042,N_2760,N_2893);
and U3043 (N_3043,N_2790,N_2822);
or U3044 (N_3044,N_2811,N_2896);
or U3045 (N_3045,N_2961,N_2955);
xnor U3046 (N_3046,N_2900,N_2753);
nor U3047 (N_3047,N_2798,N_2878);
nor U3048 (N_3048,N_2852,N_2873);
nand U3049 (N_3049,N_2953,N_2830);
nor U3050 (N_3050,N_2899,N_2881);
xor U3051 (N_3051,N_2841,N_2788);
xor U3052 (N_3052,N_2847,N_2860);
xor U3053 (N_3053,N_2792,N_2985);
xnor U3054 (N_3054,N_2972,N_2980);
nor U3055 (N_3055,N_2937,N_2768);
and U3056 (N_3056,N_2754,N_2846);
nand U3057 (N_3057,N_2796,N_2987);
and U3058 (N_3058,N_2826,N_2762);
nor U3059 (N_3059,N_2907,N_2908);
nand U3060 (N_3060,N_2882,N_2895);
nand U3061 (N_3061,N_2759,N_2894);
xnor U3062 (N_3062,N_2969,N_2998);
nor U3063 (N_3063,N_2943,N_2804);
nor U3064 (N_3064,N_2813,N_2793);
or U3065 (N_3065,N_2799,N_2802);
nor U3066 (N_3066,N_2983,N_2842);
nor U3067 (N_3067,N_2951,N_2905);
nand U3068 (N_3068,N_2904,N_2925);
nor U3069 (N_3069,N_2935,N_2785);
and U3070 (N_3070,N_2988,N_2779);
nand U3071 (N_3071,N_2833,N_2851);
nor U3072 (N_3072,N_2930,N_2995);
and U3073 (N_3073,N_2794,N_2964);
and U3074 (N_3074,N_2934,N_2781);
xnor U3075 (N_3075,N_2773,N_2864);
xor U3076 (N_3076,N_2991,N_2948);
and U3077 (N_3077,N_2917,N_2848);
nand U3078 (N_3078,N_2928,N_2902);
or U3079 (N_3079,N_2950,N_2766);
nor U3080 (N_3080,N_2918,N_2919);
and U3081 (N_3081,N_2839,N_2757);
nor U3082 (N_3082,N_2996,N_2957);
and U3083 (N_3083,N_2777,N_2844);
nor U3084 (N_3084,N_2823,N_2949);
xor U3085 (N_3085,N_2886,N_2769);
or U3086 (N_3086,N_2962,N_2906);
and U3087 (N_3087,N_2803,N_2933);
or U3088 (N_3088,N_2982,N_2845);
xnor U3089 (N_3089,N_2920,N_2926);
nor U3090 (N_3090,N_2836,N_2765);
nand U3091 (N_3091,N_2921,N_2939);
xnor U3092 (N_3092,N_2850,N_2789);
and U3093 (N_3093,N_2816,N_2963);
and U3094 (N_3094,N_2795,N_2914);
or U3095 (N_3095,N_2857,N_2891);
nand U3096 (N_3096,N_2815,N_2800);
nor U3097 (N_3097,N_2977,N_2778);
or U3098 (N_3098,N_2879,N_2990);
or U3099 (N_3099,N_2876,N_2889);
and U3100 (N_3100,N_2942,N_2787);
and U3101 (N_3101,N_2913,N_2941);
nand U3102 (N_3102,N_2909,N_2767);
nor U3103 (N_3103,N_2971,N_2883);
or U3104 (N_3104,N_2940,N_2761);
or U3105 (N_3105,N_2871,N_2965);
or U3106 (N_3106,N_2825,N_2776);
and U3107 (N_3107,N_2855,N_2819);
nor U3108 (N_3108,N_2887,N_2783);
nor U3109 (N_3109,N_2750,N_2976);
or U3110 (N_3110,N_2898,N_2862);
or U3111 (N_3111,N_2956,N_2959);
or U3112 (N_3112,N_2849,N_2999);
nand U3113 (N_3113,N_2936,N_2770);
xnor U3114 (N_3114,N_2888,N_2831);
or U3115 (N_3115,N_2931,N_2973);
and U3116 (N_3116,N_2885,N_2866);
or U3117 (N_3117,N_2807,N_2801);
nand U3118 (N_3118,N_2858,N_2903);
nor U3119 (N_3119,N_2986,N_2805);
nand U3120 (N_3120,N_2784,N_2834);
xnor U3121 (N_3121,N_2880,N_2791);
nand U3122 (N_3122,N_2975,N_2946);
xor U3123 (N_3123,N_2997,N_2875);
nand U3124 (N_3124,N_2978,N_2786);
xnor U3125 (N_3125,N_2783,N_2959);
or U3126 (N_3126,N_2783,N_2814);
xnor U3127 (N_3127,N_2794,N_2895);
xnor U3128 (N_3128,N_2862,N_2826);
or U3129 (N_3129,N_2910,N_2824);
and U3130 (N_3130,N_2974,N_2793);
xor U3131 (N_3131,N_2848,N_2981);
and U3132 (N_3132,N_2768,N_2962);
and U3133 (N_3133,N_2773,N_2777);
or U3134 (N_3134,N_2839,N_2890);
or U3135 (N_3135,N_2969,N_2787);
or U3136 (N_3136,N_2955,N_2886);
nand U3137 (N_3137,N_2814,N_2966);
nor U3138 (N_3138,N_2785,N_2978);
or U3139 (N_3139,N_2986,N_2985);
and U3140 (N_3140,N_2934,N_2802);
and U3141 (N_3141,N_2953,N_2752);
and U3142 (N_3142,N_2952,N_2924);
nor U3143 (N_3143,N_2839,N_2969);
or U3144 (N_3144,N_2945,N_2865);
nand U3145 (N_3145,N_2990,N_2954);
or U3146 (N_3146,N_2925,N_2946);
or U3147 (N_3147,N_2869,N_2885);
or U3148 (N_3148,N_2975,N_2879);
xnor U3149 (N_3149,N_2899,N_2975);
nand U3150 (N_3150,N_2777,N_2930);
nor U3151 (N_3151,N_2932,N_2938);
or U3152 (N_3152,N_2897,N_2760);
xor U3153 (N_3153,N_2864,N_2948);
or U3154 (N_3154,N_2839,N_2782);
or U3155 (N_3155,N_2840,N_2805);
and U3156 (N_3156,N_2953,N_2766);
nor U3157 (N_3157,N_2870,N_2890);
nor U3158 (N_3158,N_2875,N_2991);
nand U3159 (N_3159,N_2800,N_2920);
and U3160 (N_3160,N_2875,N_2864);
or U3161 (N_3161,N_2914,N_2988);
or U3162 (N_3162,N_2774,N_2945);
or U3163 (N_3163,N_2845,N_2803);
nor U3164 (N_3164,N_2772,N_2894);
nand U3165 (N_3165,N_2754,N_2892);
xor U3166 (N_3166,N_2879,N_2938);
nor U3167 (N_3167,N_2760,N_2966);
and U3168 (N_3168,N_2862,N_2982);
nor U3169 (N_3169,N_2918,N_2890);
and U3170 (N_3170,N_2903,N_2845);
or U3171 (N_3171,N_2902,N_2932);
and U3172 (N_3172,N_2837,N_2865);
nand U3173 (N_3173,N_2956,N_2931);
nand U3174 (N_3174,N_2835,N_2897);
or U3175 (N_3175,N_2975,N_2969);
xnor U3176 (N_3176,N_2759,N_2974);
xor U3177 (N_3177,N_2955,N_2795);
and U3178 (N_3178,N_2828,N_2894);
xnor U3179 (N_3179,N_2942,N_2848);
nor U3180 (N_3180,N_2848,N_2975);
xnor U3181 (N_3181,N_2817,N_2836);
xnor U3182 (N_3182,N_2910,N_2758);
nand U3183 (N_3183,N_2997,N_2984);
nor U3184 (N_3184,N_2890,N_2953);
and U3185 (N_3185,N_2771,N_2828);
nor U3186 (N_3186,N_2791,N_2919);
or U3187 (N_3187,N_2763,N_2984);
nor U3188 (N_3188,N_2793,N_2841);
nor U3189 (N_3189,N_2971,N_2830);
or U3190 (N_3190,N_2759,N_2779);
nor U3191 (N_3191,N_2945,N_2952);
or U3192 (N_3192,N_2811,N_2889);
and U3193 (N_3193,N_2772,N_2917);
or U3194 (N_3194,N_2981,N_2975);
and U3195 (N_3195,N_2978,N_2964);
and U3196 (N_3196,N_2795,N_2822);
or U3197 (N_3197,N_2994,N_2956);
nor U3198 (N_3198,N_2999,N_2960);
and U3199 (N_3199,N_2869,N_2998);
nand U3200 (N_3200,N_2942,N_2979);
nor U3201 (N_3201,N_2772,N_2852);
nor U3202 (N_3202,N_2891,N_2997);
or U3203 (N_3203,N_2949,N_2835);
or U3204 (N_3204,N_2983,N_2774);
or U3205 (N_3205,N_2818,N_2811);
and U3206 (N_3206,N_2862,N_2859);
or U3207 (N_3207,N_2990,N_2937);
or U3208 (N_3208,N_2902,N_2806);
nand U3209 (N_3209,N_2903,N_2963);
or U3210 (N_3210,N_2869,N_2907);
nand U3211 (N_3211,N_2754,N_2938);
nand U3212 (N_3212,N_2829,N_2918);
nor U3213 (N_3213,N_2817,N_2763);
nor U3214 (N_3214,N_2884,N_2879);
nor U3215 (N_3215,N_2948,N_2994);
nor U3216 (N_3216,N_2793,N_2773);
or U3217 (N_3217,N_2833,N_2857);
xor U3218 (N_3218,N_2791,N_2939);
or U3219 (N_3219,N_2961,N_2864);
nor U3220 (N_3220,N_2910,N_2906);
nand U3221 (N_3221,N_2805,N_2785);
nand U3222 (N_3222,N_2792,N_2797);
or U3223 (N_3223,N_2813,N_2949);
nand U3224 (N_3224,N_2891,N_2965);
or U3225 (N_3225,N_2936,N_2933);
nand U3226 (N_3226,N_2904,N_2905);
or U3227 (N_3227,N_2954,N_2866);
nand U3228 (N_3228,N_2996,N_2866);
nand U3229 (N_3229,N_2756,N_2810);
xor U3230 (N_3230,N_2788,N_2854);
nand U3231 (N_3231,N_2750,N_2890);
nor U3232 (N_3232,N_2895,N_2859);
and U3233 (N_3233,N_2767,N_2790);
nand U3234 (N_3234,N_2903,N_2750);
nor U3235 (N_3235,N_2857,N_2979);
or U3236 (N_3236,N_2863,N_2969);
nor U3237 (N_3237,N_2954,N_2883);
nand U3238 (N_3238,N_2786,N_2754);
and U3239 (N_3239,N_2860,N_2859);
nor U3240 (N_3240,N_2807,N_2995);
nand U3241 (N_3241,N_2936,N_2772);
nor U3242 (N_3242,N_2762,N_2874);
nand U3243 (N_3243,N_2913,N_2932);
nor U3244 (N_3244,N_2805,N_2855);
and U3245 (N_3245,N_2988,N_2896);
nand U3246 (N_3246,N_2941,N_2865);
nand U3247 (N_3247,N_2822,N_2888);
nand U3248 (N_3248,N_2797,N_2961);
and U3249 (N_3249,N_2833,N_2894);
and U3250 (N_3250,N_3095,N_3047);
nand U3251 (N_3251,N_3166,N_3038);
and U3252 (N_3252,N_3097,N_3058);
or U3253 (N_3253,N_3176,N_3165);
nand U3254 (N_3254,N_3052,N_3148);
nor U3255 (N_3255,N_3001,N_3159);
and U3256 (N_3256,N_3205,N_3168);
and U3257 (N_3257,N_3073,N_3172);
and U3258 (N_3258,N_3040,N_3241);
or U3259 (N_3259,N_3138,N_3034);
nor U3260 (N_3260,N_3015,N_3014);
and U3261 (N_3261,N_3157,N_3077);
nor U3262 (N_3262,N_3169,N_3065);
nand U3263 (N_3263,N_3163,N_3170);
nor U3264 (N_3264,N_3107,N_3217);
nor U3265 (N_3265,N_3190,N_3211);
xnor U3266 (N_3266,N_3142,N_3013);
nor U3267 (N_3267,N_3234,N_3067);
nand U3268 (N_3268,N_3048,N_3027);
or U3269 (N_3269,N_3066,N_3146);
nand U3270 (N_3270,N_3192,N_3150);
xor U3271 (N_3271,N_3120,N_3186);
nor U3272 (N_3272,N_3009,N_3042);
nand U3273 (N_3273,N_3237,N_3227);
nand U3274 (N_3274,N_3083,N_3208);
nor U3275 (N_3275,N_3119,N_3080);
and U3276 (N_3276,N_3152,N_3000);
nand U3277 (N_3277,N_3210,N_3092);
or U3278 (N_3278,N_3082,N_3122);
or U3279 (N_3279,N_3200,N_3236);
or U3280 (N_3280,N_3071,N_3232);
xor U3281 (N_3281,N_3091,N_3156);
and U3282 (N_3282,N_3002,N_3088);
nor U3283 (N_3283,N_3145,N_3089);
nor U3284 (N_3284,N_3063,N_3188);
nor U3285 (N_3285,N_3182,N_3036);
nor U3286 (N_3286,N_3181,N_3112);
or U3287 (N_3287,N_3102,N_3174);
xor U3288 (N_3288,N_3243,N_3116);
nand U3289 (N_3289,N_3031,N_3184);
nor U3290 (N_3290,N_3106,N_3161);
or U3291 (N_3291,N_3032,N_3151);
xor U3292 (N_3292,N_3085,N_3129);
xnor U3293 (N_3293,N_3059,N_3053);
and U3294 (N_3294,N_3203,N_3007);
or U3295 (N_3295,N_3149,N_3127);
and U3296 (N_3296,N_3055,N_3228);
nor U3297 (N_3297,N_3075,N_3191);
and U3298 (N_3298,N_3219,N_3074);
xor U3299 (N_3299,N_3030,N_3160);
and U3300 (N_3300,N_3134,N_3117);
or U3301 (N_3301,N_3179,N_3024);
nand U3302 (N_3302,N_3239,N_3054);
and U3303 (N_3303,N_3212,N_3143);
or U3304 (N_3304,N_3155,N_3115);
nand U3305 (N_3305,N_3056,N_3235);
nor U3306 (N_3306,N_3213,N_3123);
or U3307 (N_3307,N_3189,N_3049);
and U3308 (N_3308,N_3060,N_3139);
or U3309 (N_3309,N_3197,N_3064);
nor U3310 (N_3310,N_3051,N_3206);
and U3311 (N_3311,N_3187,N_3005);
or U3312 (N_3312,N_3025,N_3231);
nor U3313 (N_3313,N_3238,N_3140);
nand U3314 (N_3314,N_3041,N_3098);
or U3315 (N_3315,N_3185,N_3247);
or U3316 (N_3316,N_3183,N_3039);
or U3317 (N_3317,N_3158,N_3099);
nor U3318 (N_3318,N_3124,N_3068);
nor U3319 (N_3319,N_3101,N_3126);
or U3320 (N_3320,N_3010,N_3028);
and U3321 (N_3321,N_3195,N_3125);
or U3322 (N_3322,N_3130,N_3220);
or U3323 (N_3323,N_3100,N_3128);
or U3324 (N_3324,N_3105,N_3114);
nor U3325 (N_3325,N_3233,N_3164);
nor U3326 (N_3326,N_3118,N_3147);
and U3327 (N_3327,N_3173,N_3214);
and U3328 (N_3328,N_3222,N_3196);
and U3329 (N_3329,N_3070,N_3198);
or U3330 (N_3330,N_3135,N_3094);
nor U3331 (N_3331,N_3076,N_3061);
xnor U3332 (N_3332,N_3072,N_3090);
nor U3333 (N_3333,N_3225,N_3035);
nor U3334 (N_3334,N_3242,N_3137);
and U3335 (N_3335,N_3177,N_3045);
and U3336 (N_3336,N_3141,N_3218);
or U3337 (N_3337,N_3215,N_3103);
nand U3338 (N_3338,N_3171,N_3050);
nor U3339 (N_3339,N_3162,N_3021);
nand U3340 (N_3340,N_3023,N_3110);
or U3341 (N_3341,N_3223,N_3104);
and U3342 (N_3342,N_3136,N_3019);
and U3343 (N_3343,N_3093,N_3224);
and U3344 (N_3344,N_3230,N_3006);
or U3345 (N_3345,N_3193,N_3046);
xor U3346 (N_3346,N_3249,N_3244);
and U3347 (N_3347,N_3062,N_3026);
nor U3348 (N_3348,N_3167,N_3180);
or U3349 (N_3349,N_3087,N_3086);
or U3350 (N_3350,N_3069,N_3044);
or U3351 (N_3351,N_3144,N_3022);
and U3352 (N_3352,N_3109,N_3154);
nand U3353 (N_3353,N_3018,N_3121);
xor U3354 (N_3354,N_3079,N_3003);
nor U3355 (N_3355,N_3016,N_3043);
nor U3356 (N_3356,N_3078,N_3108);
or U3357 (N_3357,N_3096,N_3229);
or U3358 (N_3358,N_3153,N_3057);
and U3359 (N_3359,N_3199,N_3081);
and U3360 (N_3360,N_3240,N_3111);
and U3361 (N_3361,N_3029,N_3216);
and U3362 (N_3362,N_3246,N_3209);
nor U3363 (N_3363,N_3113,N_3033);
nor U3364 (N_3364,N_3037,N_3194);
xor U3365 (N_3365,N_3202,N_3011);
and U3366 (N_3366,N_3084,N_3226);
and U3367 (N_3367,N_3175,N_3008);
or U3368 (N_3368,N_3132,N_3201);
nand U3369 (N_3369,N_3012,N_3178);
nand U3370 (N_3370,N_3245,N_3017);
or U3371 (N_3371,N_3207,N_3004);
nor U3372 (N_3372,N_3248,N_3221);
xnor U3373 (N_3373,N_3020,N_3204);
or U3374 (N_3374,N_3131,N_3133);
nand U3375 (N_3375,N_3077,N_3117);
or U3376 (N_3376,N_3066,N_3015);
nor U3377 (N_3377,N_3141,N_3237);
and U3378 (N_3378,N_3161,N_3007);
or U3379 (N_3379,N_3216,N_3103);
nor U3380 (N_3380,N_3200,N_3192);
or U3381 (N_3381,N_3193,N_3215);
nor U3382 (N_3382,N_3135,N_3175);
nor U3383 (N_3383,N_3042,N_3180);
and U3384 (N_3384,N_3185,N_3042);
nand U3385 (N_3385,N_3146,N_3236);
and U3386 (N_3386,N_3200,N_3021);
or U3387 (N_3387,N_3230,N_3183);
or U3388 (N_3388,N_3197,N_3001);
xnor U3389 (N_3389,N_3102,N_3189);
nor U3390 (N_3390,N_3145,N_3162);
or U3391 (N_3391,N_3225,N_3184);
and U3392 (N_3392,N_3143,N_3246);
or U3393 (N_3393,N_3031,N_3053);
or U3394 (N_3394,N_3154,N_3203);
nor U3395 (N_3395,N_3084,N_3056);
and U3396 (N_3396,N_3065,N_3044);
xor U3397 (N_3397,N_3122,N_3019);
and U3398 (N_3398,N_3145,N_3033);
xnor U3399 (N_3399,N_3063,N_3122);
nand U3400 (N_3400,N_3158,N_3074);
and U3401 (N_3401,N_3094,N_3132);
nand U3402 (N_3402,N_3034,N_3240);
nand U3403 (N_3403,N_3168,N_3093);
or U3404 (N_3404,N_3110,N_3098);
or U3405 (N_3405,N_3248,N_3183);
and U3406 (N_3406,N_3144,N_3090);
xnor U3407 (N_3407,N_3238,N_3063);
and U3408 (N_3408,N_3026,N_3154);
or U3409 (N_3409,N_3048,N_3136);
and U3410 (N_3410,N_3230,N_3137);
and U3411 (N_3411,N_3070,N_3029);
nand U3412 (N_3412,N_3086,N_3059);
nand U3413 (N_3413,N_3033,N_3107);
nor U3414 (N_3414,N_3074,N_3189);
nand U3415 (N_3415,N_3195,N_3210);
nand U3416 (N_3416,N_3136,N_3169);
or U3417 (N_3417,N_3130,N_3132);
nor U3418 (N_3418,N_3172,N_3146);
and U3419 (N_3419,N_3015,N_3064);
nor U3420 (N_3420,N_3102,N_3052);
or U3421 (N_3421,N_3118,N_3212);
and U3422 (N_3422,N_3135,N_3186);
nand U3423 (N_3423,N_3177,N_3235);
or U3424 (N_3424,N_3096,N_3243);
xor U3425 (N_3425,N_3052,N_3031);
xor U3426 (N_3426,N_3184,N_3016);
and U3427 (N_3427,N_3209,N_3225);
or U3428 (N_3428,N_3186,N_3039);
xnor U3429 (N_3429,N_3179,N_3197);
nand U3430 (N_3430,N_3195,N_3106);
nor U3431 (N_3431,N_3187,N_3021);
nand U3432 (N_3432,N_3187,N_3049);
and U3433 (N_3433,N_3084,N_3247);
and U3434 (N_3434,N_3015,N_3186);
or U3435 (N_3435,N_3178,N_3156);
or U3436 (N_3436,N_3096,N_3058);
or U3437 (N_3437,N_3080,N_3185);
or U3438 (N_3438,N_3221,N_3211);
or U3439 (N_3439,N_3193,N_3174);
or U3440 (N_3440,N_3008,N_3137);
nand U3441 (N_3441,N_3166,N_3181);
xnor U3442 (N_3442,N_3209,N_3223);
or U3443 (N_3443,N_3216,N_3162);
and U3444 (N_3444,N_3088,N_3097);
or U3445 (N_3445,N_3213,N_3118);
nand U3446 (N_3446,N_3156,N_3176);
nand U3447 (N_3447,N_3074,N_3177);
or U3448 (N_3448,N_3060,N_3126);
and U3449 (N_3449,N_3121,N_3242);
nand U3450 (N_3450,N_3132,N_3023);
or U3451 (N_3451,N_3033,N_3129);
nand U3452 (N_3452,N_3248,N_3161);
or U3453 (N_3453,N_3035,N_3126);
nand U3454 (N_3454,N_3135,N_3034);
xor U3455 (N_3455,N_3028,N_3006);
nor U3456 (N_3456,N_3086,N_3100);
or U3457 (N_3457,N_3245,N_3244);
and U3458 (N_3458,N_3148,N_3145);
and U3459 (N_3459,N_3247,N_3016);
nor U3460 (N_3460,N_3034,N_3069);
nor U3461 (N_3461,N_3041,N_3034);
nand U3462 (N_3462,N_3131,N_3109);
and U3463 (N_3463,N_3135,N_3209);
or U3464 (N_3464,N_3195,N_3134);
and U3465 (N_3465,N_3119,N_3214);
or U3466 (N_3466,N_3050,N_3076);
or U3467 (N_3467,N_3055,N_3131);
and U3468 (N_3468,N_3016,N_3092);
nor U3469 (N_3469,N_3156,N_3145);
nand U3470 (N_3470,N_3173,N_3239);
nor U3471 (N_3471,N_3190,N_3195);
or U3472 (N_3472,N_3035,N_3037);
or U3473 (N_3473,N_3188,N_3154);
nor U3474 (N_3474,N_3162,N_3207);
nand U3475 (N_3475,N_3101,N_3062);
nand U3476 (N_3476,N_3172,N_3018);
xnor U3477 (N_3477,N_3082,N_3069);
nor U3478 (N_3478,N_3012,N_3087);
and U3479 (N_3479,N_3030,N_3204);
xor U3480 (N_3480,N_3186,N_3220);
and U3481 (N_3481,N_3149,N_3247);
nand U3482 (N_3482,N_3013,N_3247);
and U3483 (N_3483,N_3194,N_3126);
and U3484 (N_3484,N_3222,N_3081);
xnor U3485 (N_3485,N_3043,N_3186);
and U3486 (N_3486,N_3049,N_3142);
nor U3487 (N_3487,N_3075,N_3105);
nand U3488 (N_3488,N_3111,N_3083);
and U3489 (N_3489,N_3140,N_3209);
nor U3490 (N_3490,N_3003,N_3016);
and U3491 (N_3491,N_3043,N_3182);
nor U3492 (N_3492,N_3036,N_3224);
xor U3493 (N_3493,N_3211,N_3068);
xnor U3494 (N_3494,N_3203,N_3186);
and U3495 (N_3495,N_3005,N_3214);
and U3496 (N_3496,N_3074,N_3152);
nand U3497 (N_3497,N_3193,N_3138);
nand U3498 (N_3498,N_3199,N_3119);
nor U3499 (N_3499,N_3240,N_3044);
nor U3500 (N_3500,N_3350,N_3363);
nor U3501 (N_3501,N_3274,N_3337);
or U3502 (N_3502,N_3425,N_3342);
or U3503 (N_3503,N_3491,N_3432);
nor U3504 (N_3504,N_3398,N_3410);
nor U3505 (N_3505,N_3348,N_3376);
or U3506 (N_3506,N_3275,N_3367);
nand U3507 (N_3507,N_3377,N_3346);
or U3508 (N_3508,N_3356,N_3314);
nor U3509 (N_3509,N_3412,N_3389);
or U3510 (N_3510,N_3490,N_3263);
or U3511 (N_3511,N_3401,N_3400);
and U3512 (N_3512,N_3324,N_3315);
nor U3513 (N_3513,N_3321,N_3374);
nand U3514 (N_3514,N_3347,N_3396);
nor U3515 (N_3515,N_3497,N_3351);
or U3516 (N_3516,N_3279,N_3434);
or U3517 (N_3517,N_3406,N_3345);
and U3518 (N_3518,N_3286,N_3302);
nand U3519 (N_3519,N_3454,N_3301);
nor U3520 (N_3520,N_3478,N_3357);
nand U3521 (N_3521,N_3253,N_3372);
nor U3522 (N_3522,N_3289,N_3424);
or U3523 (N_3523,N_3267,N_3467);
nor U3524 (N_3524,N_3387,N_3362);
nand U3525 (N_3525,N_3499,N_3404);
and U3526 (N_3526,N_3353,N_3473);
or U3527 (N_3527,N_3438,N_3441);
nor U3528 (N_3528,N_3493,N_3299);
nand U3529 (N_3529,N_3278,N_3392);
or U3530 (N_3530,N_3468,N_3307);
xnor U3531 (N_3531,N_3369,N_3272);
nor U3532 (N_3532,N_3329,N_3413);
and U3533 (N_3533,N_3257,N_3365);
nor U3534 (N_3534,N_3487,N_3332);
nand U3535 (N_3535,N_3291,N_3323);
and U3536 (N_3536,N_3316,N_3339);
and U3537 (N_3537,N_3284,N_3384);
xor U3538 (N_3538,N_3481,N_3447);
nor U3539 (N_3539,N_3443,N_3453);
nand U3540 (N_3540,N_3411,N_3422);
or U3541 (N_3541,N_3444,N_3264);
and U3542 (N_3542,N_3488,N_3474);
nand U3543 (N_3543,N_3255,N_3446);
or U3544 (N_3544,N_3417,N_3309);
nand U3545 (N_3545,N_3330,N_3418);
nor U3546 (N_3546,N_3416,N_3254);
nor U3547 (N_3547,N_3431,N_3471);
and U3548 (N_3548,N_3451,N_3340);
nand U3549 (N_3549,N_3496,N_3300);
and U3550 (N_3550,N_3318,N_3368);
nor U3551 (N_3551,N_3360,N_3378);
nand U3552 (N_3552,N_3495,N_3338);
or U3553 (N_3553,N_3386,N_3359);
or U3554 (N_3554,N_3297,N_3426);
nand U3555 (N_3555,N_3343,N_3269);
nand U3556 (N_3556,N_3482,N_3409);
xnor U3557 (N_3557,N_3405,N_3383);
nor U3558 (N_3558,N_3415,N_3427);
nand U3559 (N_3559,N_3327,N_3288);
nor U3560 (N_3560,N_3258,N_3421);
and U3561 (N_3561,N_3399,N_3322);
nand U3562 (N_3562,N_3290,N_3485);
or U3563 (N_3563,N_3388,N_3437);
nand U3564 (N_3564,N_3465,N_3260);
and U3565 (N_3565,N_3268,N_3334);
and U3566 (N_3566,N_3270,N_3449);
nor U3567 (N_3567,N_3335,N_3381);
and U3568 (N_3568,N_3464,N_3402);
xor U3569 (N_3569,N_3331,N_3414);
nand U3570 (N_3570,N_3475,N_3479);
or U3571 (N_3571,N_3470,N_3296);
nand U3572 (N_3572,N_3480,N_3472);
nor U3573 (N_3573,N_3294,N_3458);
and U3574 (N_3574,N_3484,N_3283);
or U3575 (N_3575,N_3379,N_3361);
or U3576 (N_3576,N_3375,N_3498);
nand U3577 (N_3577,N_3256,N_3463);
xor U3578 (N_3578,N_3304,N_3469);
or U3579 (N_3579,N_3380,N_3419);
or U3580 (N_3580,N_3273,N_3276);
nand U3581 (N_3581,N_3312,N_3349);
or U3582 (N_3582,N_3298,N_3287);
nor U3583 (N_3583,N_3476,N_3460);
or U3584 (N_3584,N_3433,N_3407);
nand U3585 (N_3585,N_3391,N_3371);
nand U3586 (N_3586,N_3259,N_3428);
nand U3587 (N_3587,N_3262,N_3429);
and U3588 (N_3588,N_3445,N_3341);
and U3589 (N_3589,N_3494,N_3320);
nand U3590 (N_3590,N_3352,N_3281);
nor U3591 (N_3591,N_3282,N_3489);
or U3592 (N_3592,N_3293,N_3306);
or U3593 (N_3593,N_3395,N_3370);
nand U3594 (N_3594,N_3382,N_3450);
nand U3595 (N_3595,N_3285,N_3265);
xor U3596 (N_3596,N_3251,N_3313);
xnor U3597 (N_3597,N_3492,N_3461);
xnor U3598 (N_3598,N_3252,N_3403);
nand U3599 (N_3599,N_3394,N_3477);
xnor U3600 (N_3600,N_3336,N_3483);
and U3601 (N_3601,N_3326,N_3390);
nand U3602 (N_3602,N_3430,N_3397);
and U3603 (N_3603,N_3442,N_3385);
nand U3604 (N_3604,N_3455,N_3261);
xor U3605 (N_3605,N_3408,N_3393);
or U3606 (N_3606,N_3452,N_3355);
nand U3607 (N_3607,N_3319,N_3311);
nor U3608 (N_3608,N_3358,N_3325);
and U3609 (N_3609,N_3308,N_3456);
nor U3610 (N_3610,N_3328,N_3364);
nand U3611 (N_3611,N_3266,N_3459);
nor U3612 (N_3612,N_3317,N_3486);
and U3613 (N_3613,N_3292,N_3344);
nor U3614 (N_3614,N_3280,N_3466);
nor U3615 (N_3615,N_3277,N_3310);
xor U3616 (N_3616,N_3295,N_3271);
nand U3617 (N_3617,N_3435,N_3439);
nand U3618 (N_3618,N_3333,N_3303);
and U3619 (N_3619,N_3440,N_3420);
and U3620 (N_3620,N_3373,N_3354);
nor U3621 (N_3621,N_3366,N_3457);
or U3622 (N_3622,N_3250,N_3423);
and U3623 (N_3623,N_3436,N_3462);
nor U3624 (N_3624,N_3448,N_3305);
and U3625 (N_3625,N_3289,N_3436);
or U3626 (N_3626,N_3397,N_3265);
nor U3627 (N_3627,N_3278,N_3272);
or U3628 (N_3628,N_3498,N_3441);
nor U3629 (N_3629,N_3466,N_3284);
or U3630 (N_3630,N_3299,N_3288);
or U3631 (N_3631,N_3492,N_3296);
nand U3632 (N_3632,N_3261,N_3395);
nor U3633 (N_3633,N_3399,N_3496);
nand U3634 (N_3634,N_3417,N_3366);
nor U3635 (N_3635,N_3403,N_3273);
xnor U3636 (N_3636,N_3418,N_3423);
or U3637 (N_3637,N_3449,N_3327);
xor U3638 (N_3638,N_3257,N_3324);
nor U3639 (N_3639,N_3256,N_3389);
nor U3640 (N_3640,N_3411,N_3339);
and U3641 (N_3641,N_3476,N_3334);
or U3642 (N_3642,N_3448,N_3352);
nand U3643 (N_3643,N_3387,N_3304);
nand U3644 (N_3644,N_3304,N_3289);
nand U3645 (N_3645,N_3476,N_3342);
nand U3646 (N_3646,N_3475,N_3269);
xor U3647 (N_3647,N_3286,N_3421);
or U3648 (N_3648,N_3326,N_3452);
nand U3649 (N_3649,N_3394,N_3457);
or U3650 (N_3650,N_3347,N_3384);
nand U3651 (N_3651,N_3478,N_3333);
xor U3652 (N_3652,N_3442,N_3485);
and U3653 (N_3653,N_3321,N_3467);
xnor U3654 (N_3654,N_3308,N_3337);
nor U3655 (N_3655,N_3444,N_3265);
and U3656 (N_3656,N_3476,N_3401);
or U3657 (N_3657,N_3375,N_3389);
nand U3658 (N_3658,N_3282,N_3342);
nand U3659 (N_3659,N_3434,N_3462);
and U3660 (N_3660,N_3415,N_3265);
nor U3661 (N_3661,N_3344,N_3426);
or U3662 (N_3662,N_3455,N_3276);
nand U3663 (N_3663,N_3460,N_3269);
or U3664 (N_3664,N_3264,N_3416);
xor U3665 (N_3665,N_3359,N_3451);
nor U3666 (N_3666,N_3308,N_3463);
or U3667 (N_3667,N_3474,N_3485);
nand U3668 (N_3668,N_3290,N_3266);
nand U3669 (N_3669,N_3432,N_3307);
nor U3670 (N_3670,N_3371,N_3311);
nor U3671 (N_3671,N_3361,N_3382);
or U3672 (N_3672,N_3396,N_3315);
nor U3673 (N_3673,N_3384,N_3265);
nor U3674 (N_3674,N_3398,N_3421);
and U3675 (N_3675,N_3492,N_3361);
nor U3676 (N_3676,N_3327,N_3303);
nor U3677 (N_3677,N_3489,N_3468);
nor U3678 (N_3678,N_3361,N_3272);
or U3679 (N_3679,N_3348,N_3264);
or U3680 (N_3680,N_3455,N_3312);
or U3681 (N_3681,N_3461,N_3256);
nor U3682 (N_3682,N_3391,N_3473);
or U3683 (N_3683,N_3403,N_3290);
or U3684 (N_3684,N_3274,N_3410);
and U3685 (N_3685,N_3442,N_3488);
nand U3686 (N_3686,N_3328,N_3348);
and U3687 (N_3687,N_3403,N_3496);
xor U3688 (N_3688,N_3323,N_3466);
and U3689 (N_3689,N_3322,N_3496);
or U3690 (N_3690,N_3419,N_3466);
nor U3691 (N_3691,N_3406,N_3277);
or U3692 (N_3692,N_3437,N_3334);
xnor U3693 (N_3693,N_3254,N_3392);
and U3694 (N_3694,N_3424,N_3257);
nand U3695 (N_3695,N_3317,N_3480);
or U3696 (N_3696,N_3337,N_3384);
nor U3697 (N_3697,N_3328,N_3347);
nor U3698 (N_3698,N_3342,N_3484);
and U3699 (N_3699,N_3323,N_3328);
and U3700 (N_3700,N_3290,N_3305);
nor U3701 (N_3701,N_3457,N_3305);
and U3702 (N_3702,N_3295,N_3476);
nor U3703 (N_3703,N_3255,N_3490);
nor U3704 (N_3704,N_3320,N_3425);
xor U3705 (N_3705,N_3303,N_3253);
and U3706 (N_3706,N_3478,N_3411);
or U3707 (N_3707,N_3368,N_3299);
nor U3708 (N_3708,N_3317,N_3469);
and U3709 (N_3709,N_3295,N_3333);
nand U3710 (N_3710,N_3335,N_3372);
and U3711 (N_3711,N_3498,N_3309);
nand U3712 (N_3712,N_3491,N_3286);
nor U3713 (N_3713,N_3329,N_3266);
xor U3714 (N_3714,N_3347,N_3403);
or U3715 (N_3715,N_3408,N_3378);
nor U3716 (N_3716,N_3431,N_3477);
or U3717 (N_3717,N_3403,N_3357);
nand U3718 (N_3718,N_3460,N_3265);
or U3719 (N_3719,N_3334,N_3370);
or U3720 (N_3720,N_3460,N_3259);
nor U3721 (N_3721,N_3322,N_3457);
and U3722 (N_3722,N_3472,N_3399);
and U3723 (N_3723,N_3470,N_3370);
nor U3724 (N_3724,N_3294,N_3330);
and U3725 (N_3725,N_3448,N_3361);
nand U3726 (N_3726,N_3465,N_3480);
and U3727 (N_3727,N_3488,N_3392);
xor U3728 (N_3728,N_3351,N_3429);
or U3729 (N_3729,N_3282,N_3362);
and U3730 (N_3730,N_3367,N_3464);
nand U3731 (N_3731,N_3468,N_3339);
nor U3732 (N_3732,N_3281,N_3348);
nand U3733 (N_3733,N_3462,N_3457);
or U3734 (N_3734,N_3305,N_3475);
nor U3735 (N_3735,N_3414,N_3360);
nor U3736 (N_3736,N_3476,N_3481);
xor U3737 (N_3737,N_3458,N_3422);
and U3738 (N_3738,N_3283,N_3360);
nand U3739 (N_3739,N_3306,N_3405);
or U3740 (N_3740,N_3353,N_3270);
xnor U3741 (N_3741,N_3257,N_3396);
or U3742 (N_3742,N_3325,N_3313);
and U3743 (N_3743,N_3446,N_3266);
nor U3744 (N_3744,N_3478,N_3448);
nand U3745 (N_3745,N_3373,N_3497);
nand U3746 (N_3746,N_3292,N_3381);
xor U3747 (N_3747,N_3313,N_3378);
nand U3748 (N_3748,N_3497,N_3355);
xnor U3749 (N_3749,N_3305,N_3430);
and U3750 (N_3750,N_3657,N_3627);
nand U3751 (N_3751,N_3505,N_3547);
and U3752 (N_3752,N_3518,N_3563);
and U3753 (N_3753,N_3595,N_3671);
or U3754 (N_3754,N_3559,N_3571);
nand U3755 (N_3755,N_3646,N_3531);
nand U3756 (N_3756,N_3726,N_3558);
xnor U3757 (N_3757,N_3743,N_3517);
and U3758 (N_3758,N_3672,N_3556);
nand U3759 (N_3759,N_3693,N_3707);
xor U3760 (N_3760,N_3695,N_3676);
nor U3761 (N_3761,N_3539,N_3670);
nor U3762 (N_3762,N_3679,N_3544);
xnor U3763 (N_3763,N_3614,N_3585);
and U3764 (N_3764,N_3618,N_3749);
and U3765 (N_3765,N_3526,N_3554);
nand U3766 (N_3766,N_3713,N_3669);
nand U3767 (N_3767,N_3717,N_3740);
or U3768 (N_3768,N_3573,N_3660);
and U3769 (N_3769,N_3723,N_3674);
and U3770 (N_3770,N_3626,N_3581);
or U3771 (N_3771,N_3711,N_3644);
nand U3772 (N_3772,N_3694,N_3523);
nor U3773 (N_3773,N_3634,N_3649);
nand U3774 (N_3774,N_3586,N_3729);
or U3775 (N_3775,N_3620,N_3654);
or U3776 (N_3776,N_3622,N_3632);
or U3777 (N_3777,N_3642,N_3511);
and U3778 (N_3778,N_3550,N_3655);
xnor U3779 (N_3779,N_3639,N_3576);
and U3780 (N_3780,N_3537,N_3746);
or U3781 (N_3781,N_3663,N_3500);
and U3782 (N_3782,N_3716,N_3587);
or U3783 (N_3783,N_3513,N_3661);
nor U3784 (N_3784,N_3527,N_3534);
or U3785 (N_3785,N_3609,N_3745);
and U3786 (N_3786,N_3744,N_3536);
nand U3787 (N_3787,N_3675,N_3580);
or U3788 (N_3788,N_3708,N_3548);
and U3789 (N_3789,N_3608,N_3700);
and U3790 (N_3790,N_3619,N_3565);
nor U3791 (N_3791,N_3724,N_3666);
nand U3792 (N_3792,N_3545,N_3611);
or U3793 (N_3793,N_3612,N_3709);
and U3794 (N_3794,N_3507,N_3502);
nor U3795 (N_3795,N_3570,N_3630);
or U3796 (N_3796,N_3682,N_3692);
nand U3797 (N_3797,N_3561,N_3728);
nand U3798 (N_3798,N_3635,N_3647);
or U3799 (N_3799,N_3651,N_3699);
and U3800 (N_3800,N_3582,N_3520);
and U3801 (N_3801,N_3673,N_3541);
and U3802 (N_3802,N_3702,N_3731);
nor U3803 (N_3803,N_3638,N_3564);
and U3804 (N_3804,N_3680,N_3653);
and U3805 (N_3805,N_3562,N_3577);
or U3806 (N_3806,N_3516,N_3735);
and U3807 (N_3807,N_3528,N_3597);
and U3808 (N_3808,N_3667,N_3602);
or U3809 (N_3809,N_3583,N_3538);
or U3810 (N_3810,N_3610,N_3519);
xnor U3811 (N_3811,N_3560,N_3738);
or U3812 (N_3812,N_3697,N_3688);
and U3813 (N_3813,N_3549,N_3687);
xor U3814 (N_3814,N_3515,N_3631);
and U3815 (N_3815,N_3637,N_3529);
and U3816 (N_3816,N_3720,N_3621);
or U3817 (N_3817,N_3650,N_3551);
or U3818 (N_3818,N_3590,N_3579);
nor U3819 (N_3819,N_3705,N_3625);
or U3820 (N_3820,N_3569,N_3691);
nand U3821 (N_3821,N_3601,N_3512);
nand U3822 (N_3822,N_3659,N_3623);
nand U3823 (N_3823,N_3574,N_3546);
or U3824 (N_3824,N_3533,N_3522);
nand U3825 (N_3825,N_3572,N_3690);
nand U3826 (N_3826,N_3521,N_3555);
nor U3827 (N_3827,N_3501,N_3696);
and U3828 (N_3828,N_3600,N_3591);
and U3829 (N_3829,N_3605,N_3575);
xor U3830 (N_3830,N_3589,N_3506);
xor U3831 (N_3831,N_3662,N_3596);
nand U3832 (N_3832,N_3739,N_3540);
nand U3833 (N_3833,N_3509,N_3730);
nor U3834 (N_3834,N_3742,N_3629);
nand U3835 (N_3835,N_3734,N_3725);
nor U3836 (N_3836,N_3567,N_3508);
nand U3837 (N_3837,N_3736,N_3503);
xnor U3838 (N_3838,N_3727,N_3604);
and U3839 (N_3839,N_3584,N_3525);
and U3840 (N_3840,N_3636,N_3656);
nand U3841 (N_3841,N_3748,N_3645);
nor U3842 (N_3842,N_3652,N_3504);
nor U3843 (N_3843,N_3624,N_3588);
nand U3844 (N_3844,N_3747,N_3594);
or U3845 (N_3845,N_3568,N_3703);
xnor U3846 (N_3846,N_3607,N_3566);
or U3847 (N_3847,N_3681,N_3686);
nand U3848 (N_3848,N_3712,N_3603);
nor U3849 (N_3849,N_3633,N_3543);
or U3850 (N_3850,N_3641,N_3606);
nor U3851 (N_3851,N_3704,N_3643);
nor U3852 (N_3852,N_3698,N_3710);
nand U3853 (N_3853,N_3532,N_3578);
xnor U3854 (N_3854,N_3557,N_3732);
or U3855 (N_3855,N_3721,N_3719);
or U3856 (N_3856,N_3689,N_3542);
or U3857 (N_3857,N_3640,N_3598);
and U3858 (N_3858,N_3514,N_3685);
or U3859 (N_3859,N_3648,N_3741);
nand U3860 (N_3860,N_3510,N_3718);
nor U3861 (N_3861,N_3722,N_3733);
nor U3862 (N_3862,N_3678,N_3714);
nor U3863 (N_3863,N_3553,N_3616);
or U3864 (N_3864,N_3737,N_3628);
and U3865 (N_3865,N_3613,N_3658);
and U3866 (N_3866,N_3706,N_3701);
nand U3867 (N_3867,N_3552,N_3683);
and U3868 (N_3868,N_3599,N_3617);
or U3869 (N_3869,N_3665,N_3592);
nand U3870 (N_3870,N_3615,N_3684);
and U3871 (N_3871,N_3524,N_3664);
and U3872 (N_3872,N_3593,N_3530);
nand U3873 (N_3873,N_3715,N_3668);
nor U3874 (N_3874,N_3535,N_3677);
and U3875 (N_3875,N_3731,N_3587);
or U3876 (N_3876,N_3666,N_3742);
nand U3877 (N_3877,N_3625,N_3691);
nor U3878 (N_3878,N_3739,N_3657);
nand U3879 (N_3879,N_3600,N_3648);
or U3880 (N_3880,N_3685,N_3591);
and U3881 (N_3881,N_3525,N_3589);
xnor U3882 (N_3882,N_3542,N_3622);
and U3883 (N_3883,N_3696,N_3536);
xor U3884 (N_3884,N_3563,N_3583);
xor U3885 (N_3885,N_3695,N_3570);
nor U3886 (N_3886,N_3722,N_3734);
nand U3887 (N_3887,N_3561,N_3537);
nor U3888 (N_3888,N_3549,N_3606);
nor U3889 (N_3889,N_3684,N_3680);
and U3890 (N_3890,N_3566,N_3678);
xnor U3891 (N_3891,N_3677,N_3526);
xor U3892 (N_3892,N_3689,N_3643);
nor U3893 (N_3893,N_3638,N_3566);
nor U3894 (N_3894,N_3501,N_3630);
nor U3895 (N_3895,N_3643,N_3573);
and U3896 (N_3896,N_3500,N_3586);
xor U3897 (N_3897,N_3664,N_3544);
nor U3898 (N_3898,N_3642,N_3549);
nand U3899 (N_3899,N_3616,N_3632);
and U3900 (N_3900,N_3524,N_3739);
and U3901 (N_3901,N_3743,N_3515);
nor U3902 (N_3902,N_3710,N_3552);
or U3903 (N_3903,N_3674,N_3560);
or U3904 (N_3904,N_3524,N_3532);
or U3905 (N_3905,N_3621,N_3567);
or U3906 (N_3906,N_3696,N_3585);
and U3907 (N_3907,N_3695,N_3515);
or U3908 (N_3908,N_3568,N_3740);
nor U3909 (N_3909,N_3539,N_3740);
and U3910 (N_3910,N_3630,N_3669);
nand U3911 (N_3911,N_3661,N_3512);
nor U3912 (N_3912,N_3739,N_3710);
and U3913 (N_3913,N_3654,N_3562);
nor U3914 (N_3914,N_3549,N_3670);
and U3915 (N_3915,N_3740,N_3593);
or U3916 (N_3916,N_3568,N_3533);
or U3917 (N_3917,N_3528,N_3527);
or U3918 (N_3918,N_3644,N_3582);
or U3919 (N_3919,N_3632,N_3709);
nor U3920 (N_3920,N_3733,N_3649);
nor U3921 (N_3921,N_3664,N_3678);
nand U3922 (N_3922,N_3532,N_3508);
nand U3923 (N_3923,N_3690,N_3700);
xnor U3924 (N_3924,N_3631,N_3605);
nand U3925 (N_3925,N_3636,N_3681);
xnor U3926 (N_3926,N_3511,N_3684);
and U3927 (N_3927,N_3611,N_3721);
nand U3928 (N_3928,N_3544,N_3563);
and U3929 (N_3929,N_3602,N_3592);
and U3930 (N_3930,N_3538,N_3617);
or U3931 (N_3931,N_3596,N_3688);
nand U3932 (N_3932,N_3705,N_3620);
xnor U3933 (N_3933,N_3631,N_3555);
or U3934 (N_3934,N_3709,N_3719);
nor U3935 (N_3935,N_3522,N_3600);
and U3936 (N_3936,N_3508,N_3642);
and U3937 (N_3937,N_3633,N_3610);
or U3938 (N_3938,N_3598,N_3557);
and U3939 (N_3939,N_3542,N_3621);
or U3940 (N_3940,N_3704,N_3541);
or U3941 (N_3941,N_3524,N_3571);
and U3942 (N_3942,N_3620,N_3746);
xnor U3943 (N_3943,N_3717,N_3735);
or U3944 (N_3944,N_3615,N_3629);
and U3945 (N_3945,N_3713,N_3652);
and U3946 (N_3946,N_3560,N_3589);
or U3947 (N_3947,N_3728,N_3512);
nand U3948 (N_3948,N_3658,N_3501);
and U3949 (N_3949,N_3696,N_3620);
nand U3950 (N_3950,N_3540,N_3501);
nand U3951 (N_3951,N_3627,N_3650);
or U3952 (N_3952,N_3668,N_3552);
or U3953 (N_3953,N_3510,N_3663);
or U3954 (N_3954,N_3611,N_3653);
and U3955 (N_3955,N_3628,N_3548);
and U3956 (N_3956,N_3717,N_3744);
and U3957 (N_3957,N_3646,N_3737);
or U3958 (N_3958,N_3538,N_3736);
nor U3959 (N_3959,N_3500,N_3553);
and U3960 (N_3960,N_3553,N_3514);
nand U3961 (N_3961,N_3676,N_3539);
nand U3962 (N_3962,N_3590,N_3580);
nand U3963 (N_3963,N_3549,N_3716);
or U3964 (N_3964,N_3562,N_3710);
or U3965 (N_3965,N_3719,N_3645);
and U3966 (N_3966,N_3625,N_3500);
and U3967 (N_3967,N_3642,N_3577);
nor U3968 (N_3968,N_3629,N_3607);
and U3969 (N_3969,N_3697,N_3709);
or U3970 (N_3970,N_3684,N_3516);
or U3971 (N_3971,N_3628,N_3646);
nor U3972 (N_3972,N_3667,N_3569);
or U3973 (N_3973,N_3646,N_3537);
nor U3974 (N_3974,N_3589,N_3556);
and U3975 (N_3975,N_3556,N_3615);
nand U3976 (N_3976,N_3611,N_3575);
and U3977 (N_3977,N_3553,N_3594);
nand U3978 (N_3978,N_3720,N_3538);
and U3979 (N_3979,N_3709,N_3684);
and U3980 (N_3980,N_3629,N_3635);
or U3981 (N_3981,N_3525,N_3542);
nor U3982 (N_3982,N_3548,N_3596);
and U3983 (N_3983,N_3622,N_3512);
nor U3984 (N_3984,N_3512,N_3638);
or U3985 (N_3985,N_3668,N_3532);
nor U3986 (N_3986,N_3555,N_3635);
nor U3987 (N_3987,N_3680,N_3504);
nand U3988 (N_3988,N_3584,N_3685);
nand U3989 (N_3989,N_3730,N_3627);
nor U3990 (N_3990,N_3562,N_3568);
or U3991 (N_3991,N_3705,N_3523);
and U3992 (N_3992,N_3579,N_3553);
or U3993 (N_3993,N_3675,N_3613);
xor U3994 (N_3994,N_3693,N_3573);
and U3995 (N_3995,N_3702,N_3696);
nand U3996 (N_3996,N_3544,N_3613);
xnor U3997 (N_3997,N_3574,N_3567);
or U3998 (N_3998,N_3583,N_3595);
or U3999 (N_3999,N_3624,N_3712);
nand U4000 (N_4000,N_3910,N_3893);
and U4001 (N_4001,N_3760,N_3797);
xor U4002 (N_4002,N_3874,N_3912);
nand U4003 (N_4003,N_3911,N_3775);
or U4004 (N_4004,N_3882,N_3751);
or U4005 (N_4005,N_3790,N_3856);
or U4006 (N_4006,N_3791,N_3991);
nor U4007 (N_4007,N_3984,N_3754);
or U4008 (N_4008,N_3805,N_3941);
or U4009 (N_4009,N_3782,N_3927);
nor U4010 (N_4010,N_3809,N_3871);
xnor U4011 (N_4011,N_3982,N_3973);
nand U4012 (N_4012,N_3811,N_3855);
or U4013 (N_4013,N_3944,N_3960);
or U4014 (N_4014,N_3956,N_3950);
nor U4015 (N_4015,N_3847,N_3819);
and U4016 (N_4016,N_3995,N_3878);
or U4017 (N_4017,N_3920,N_3965);
nand U4018 (N_4018,N_3824,N_3986);
or U4019 (N_4019,N_3774,N_3947);
nand U4020 (N_4020,N_3903,N_3955);
and U4021 (N_4021,N_3755,N_3859);
nor U4022 (N_4022,N_3877,N_3786);
nand U4023 (N_4023,N_3817,N_3904);
nand U4024 (N_4024,N_3821,N_3867);
nand U4025 (N_4025,N_3770,N_3784);
xnor U4026 (N_4026,N_3943,N_3834);
or U4027 (N_4027,N_3979,N_3967);
or U4028 (N_4028,N_3829,N_3895);
nand U4029 (N_4029,N_3917,N_3822);
or U4030 (N_4030,N_3861,N_3849);
or U4031 (N_4031,N_3933,N_3778);
nand U4032 (N_4032,N_3814,N_3899);
nor U4033 (N_4033,N_3988,N_3891);
or U4034 (N_4034,N_3881,N_3905);
nor U4035 (N_4035,N_3923,N_3862);
xor U4036 (N_4036,N_3919,N_3883);
or U4037 (N_4037,N_3966,N_3866);
nand U4038 (N_4038,N_3793,N_3981);
nor U4039 (N_4039,N_3900,N_3975);
and U4040 (N_4040,N_3873,N_3785);
xor U4041 (N_4041,N_3974,N_3752);
or U4042 (N_4042,N_3964,N_3922);
nand U4043 (N_4043,N_3761,N_3827);
nand U4044 (N_4044,N_3940,N_3845);
or U4045 (N_4045,N_3875,N_3779);
or U4046 (N_4046,N_3803,N_3997);
or U4047 (N_4047,N_3870,N_3958);
and U4048 (N_4048,N_3976,N_3896);
nand U4049 (N_4049,N_3839,N_3840);
nor U4050 (N_4050,N_3852,N_3915);
nand U4051 (N_4051,N_3837,N_3977);
nor U4052 (N_4052,N_3906,N_3796);
and U4053 (N_4053,N_3804,N_3853);
nor U4054 (N_4054,N_3913,N_3812);
or U4055 (N_4055,N_3970,N_3934);
and U4056 (N_4056,N_3802,N_3808);
and U4057 (N_4057,N_3777,N_3789);
nand U4058 (N_4058,N_3836,N_3929);
or U4059 (N_4059,N_3924,N_3825);
or U4060 (N_4060,N_3949,N_3901);
and U4061 (N_4061,N_3945,N_3928);
xor U4062 (N_4062,N_3869,N_3816);
nand U4063 (N_4063,N_3807,N_3897);
or U4064 (N_4064,N_3783,N_3936);
and U4065 (N_4065,N_3946,N_3983);
nand U4066 (N_4066,N_3892,N_3963);
nand U4067 (N_4067,N_3762,N_3801);
xor U4068 (N_4068,N_3880,N_3833);
or U4069 (N_4069,N_3888,N_3794);
or U4070 (N_4070,N_3787,N_3843);
nand U4071 (N_4071,N_3926,N_3772);
or U4072 (N_4072,N_3872,N_3930);
and U4073 (N_4073,N_3889,N_3876);
nor U4074 (N_4074,N_3818,N_3885);
or U4075 (N_4075,N_3962,N_3854);
or U4076 (N_4076,N_3771,N_3992);
and U4077 (N_4077,N_3769,N_3850);
or U4078 (N_4078,N_3815,N_3894);
and U4079 (N_4079,N_3792,N_3863);
nor U4080 (N_4080,N_3914,N_3971);
and U4081 (N_4081,N_3952,N_3980);
and U4082 (N_4082,N_3753,N_3806);
xnor U4083 (N_4083,N_3957,N_3954);
nand U4084 (N_4084,N_3961,N_3830);
or U4085 (N_4085,N_3842,N_3820);
nor U4086 (N_4086,N_3908,N_3826);
nor U4087 (N_4087,N_3886,N_3994);
nor U4088 (N_4088,N_3953,N_3884);
nor U4089 (N_4089,N_3993,N_3758);
and U4090 (N_4090,N_3773,N_3989);
xor U4091 (N_4091,N_3844,N_3799);
or U4092 (N_4092,N_3925,N_3764);
nand U4093 (N_4093,N_3767,N_3813);
and U4094 (N_4094,N_3838,N_3841);
nand U4095 (N_4095,N_3931,N_3985);
nand U4096 (N_4096,N_3781,N_3951);
nor U4097 (N_4097,N_3831,N_3902);
xor U4098 (N_4098,N_3865,N_3959);
and U4099 (N_4099,N_3823,N_3935);
nand U4100 (N_4100,N_3757,N_3969);
nor U4101 (N_4101,N_3750,N_3909);
or U4102 (N_4102,N_3851,N_3978);
and U4103 (N_4103,N_3763,N_3998);
nor U4104 (N_4104,N_3828,N_3756);
nor U4105 (N_4105,N_3898,N_3968);
nand U4106 (N_4106,N_3759,N_3810);
and U4107 (N_4107,N_3937,N_3798);
xnor U4108 (N_4108,N_3846,N_3864);
nand U4109 (N_4109,N_3848,N_3832);
nor U4110 (N_4110,N_3942,N_3860);
nor U4111 (N_4111,N_3918,N_3921);
nor U4112 (N_4112,N_3990,N_3948);
and U4113 (N_4113,N_3795,N_3765);
nor U4114 (N_4114,N_3788,N_3932);
nand U4115 (N_4115,N_3887,N_3890);
and U4116 (N_4116,N_3916,N_3996);
and U4117 (N_4117,N_3858,N_3776);
nand U4118 (N_4118,N_3879,N_3766);
or U4119 (N_4119,N_3939,N_3800);
or U4120 (N_4120,N_3857,N_3907);
nor U4121 (N_4121,N_3780,N_3938);
nand U4122 (N_4122,N_3768,N_3999);
nand U4123 (N_4123,N_3868,N_3835);
xor U4124 (N_4124,N_3987,N_3972);
xor U4125 (N_4125,N_3830,N_3960);
nand U4126 (N_4126,N_3815,N_3938);
nor U4127 (N_4127,N_3803,N_3919);
nand U4128 (N_4128,N_3961,N_3757);
nor U4129 (N_4129,N_3821,N_3873);
and U4130 (N_4130,N_3931,N_3973);
and U4131 (N_4131,N_3992,N_3851);
nand U4132 (N_4132,N_3894,N_3823);
nand U4133 (N_4133,N_3862,N_3981);
xnor U4134 (N_4134,N_3866,N_3784);
xor U4135 (N_4135,N_3942,N_3972);
and U4136 (N_4136,N_3843,N_3980);
and U4137 (N_4137,N_3963,N_3825);
or U4138 (N_4138,N_3956,N_3786);
or U4139 (N_4139,N_3771,N_3975);
xnor U4140 (N_4140,N_3896,N_3955);
and U4141 (N_4141,N_3938,N_3980);
nor U4142 (N_4142,N_3820,N_3966);
or U4143 (N_4143,N_3755,N_3918);
xor U4144 (N_4144,N_3806,N_3971);
or U4145 (N_4145,N_3991,N_3763);
xnor U4146 (N_4146,N_3960,N_3753);
and U4147 (N_4147,N_3834,N_3803);
xor U4148 (N_4148,N_3865,N_3784);
and U4149 (N_4149,N_3778,N_3755);
or U4150 (N_4150,N_3893,N_3813);
nand U4151 (N_4151,N_3993,N_3940);
nor U4152 (N_4152,N_3909,N_3973);
nor U4153 (N_4153,N_3999,N_3761);
nor U4154 (N_4154,N_3875,N_3765);
and U4155 (N_4155,N_3853,N_3966);
and U4156 (N_4156,N_3844,N_3855);
or U4157 (N_4157,N_3836,N_3858);
nor U4158 (N_4158,N_3966,N_3828);
and U4159 (N_4159,N_3751,N_3989);
or U4160 (N_4160,N_3875,N_3993);
or U4161 (N_4161,N_3754,N_3839);
and U4162 (N_4162,N_3946,N_3801);
nor U4163 (N_4163,N_3815,N_3872);
nor U4164 (N_4164,N_3911,N_3870);
or U4165 (N_4165,N_3814,N_3849);
or U4166 (N_4166,N_3874,N_3872);
and U4167 (N_4167,N_3944,N_3753);
and U4168 (N_4168,N_3936,N_3874);
nand U4169 (N_4169,N_3815,N_3838);
nand U4170 (N_4170,N_3786,N_3837);
nand U4171 (N_4171,N_3924,N_3901);
nand U4172 (N_4172,N_3941,N_3834);
nor U4173 (N_4173,N_3756,N_3948);
nand U4174 (N_4174,N_3855,N_3820);
xnor U4175 (N_4175,N_3750,N_3985);
nand U4176 (N_4176,N_3987,N_3868);
and U4177 (N_4177,N_3888,N_3835);
or U4178 (N_4178,N_3986,N_3786);
xnor U4179 (N_4179,N_3849,N_3993);
nand U4180 (N_4180,N_3921,N_3776);
or U4181 (N_4181,N_3973,N_3824);
nor U4182 (N_4182,N_3971,N_3821);
nor U4183 (N_4183,N_3943,N_3763);
or U4184 (N_4184,N_3773,N_3811);
xnor U4185 (N_4185,N_3917,N_3860);
and U4186 (N_4186,N_3992,N_3831);
nand U4187 (N_4187,N_3769,N_3952);
nor U4188 (N_4188,N_3997,N_3831);
nor U4189 (N_4189,N_3877,N_3913);
xor U4190 (N_4190,N_3932,N_3899);
and U4191 (N_4191,N_3853,N_3975);
nor U4192 (N_4192,N_3768,N_3952);
xor U4193 (N_4193,N_3783,N_3985);
nand U4194 (N_4194,N_3867,N_3876);
nand U4195 (N_4195,N_3792,N_3820);
nand U4196 (N_4196,N_3852,N_3963);
nand U4197 (N_4197,N_3806,N_3769);
xor U4198 (N_4198,N_3801,N_3885);
xor U4199 (N_4199,N_3751,N_3982);
nor U4200 (N_4200,N_3814,N_3957);
nand U4201 (N_4201,N_3893,N_3901);
or U4202 (N_4202,N_3921,N_3941);
nand U4203 (N_4203,N_3906,N_3838);
xnor U4204 (N_4204,N_3827,N_3982);
nor U4205 (N_4205,N_3908,N_3754);
xor U4206 (N_4206,N_3998,N_3973);
and U4207 (N_4207,N_3976,N_3975);
nor U4208 (N_4208,N_3917,N_3955);
and U4209 (N_4209,N_3750,N_3912);
nand U4210 (N_4210,N_3758,N_3864);
nor U4211 (N_4211,N_3842,N_3944);
or U4212 (N_4212,N_3965,N_3933);
nand U4213 (N_4213,N_3753,N_3810);
nor U4214 (N_4214,N_3880,N_3894);
nor U4215 (N_4215,N_3758,N_3861);
or U4216 (N_4216,N_3778,N_3979);
xor U4217 (N_4217,N_3753,N_3852);
or U4218 (N_4218,N_3871,N_3990);
nand U4219 (N_4219,N_3965,N_3855);
nand U4220 (N_4220,N_3828,N_3944);
xor U4221 (N_4221,N_3820,N_3939);
xor U4222 (N_4222,N_3807,N_3981);
and U4223 (N_4223,N_3989,N_3898);
or U4224 (N_4224,N_3770,N_3941);
nand U4225 (N_4225,N_3989,N_3972);
or U4226 (N_4226,N_3879,N_3963);
or U4227 (N_4227,N_3996,N_3913);
and U4228 (N_4228,N_3777,N_3821);
nor U4229 (N_4229,N_3937,N_3993);
nor U4230 (N_4230,N_3853,N_3867);
nor U4231 (N_4231,N_3927,N_3985);
nor U4232 (N_4232,N_3900,N_3907);
and U4233 (N_4233,N_3751,N_3785);
and U4234 (N_4234,N_3891,N_3908);
and U4235 (N_4235,N_3920,N_3917);
nor U4236 (N_4236,N_3886,N_3764);
and U4237 (N_4237,N_3982,N_3829);
and U4238 (N_4238,N_3960,N_3865);
xor U4239 (N_4239,N_3831,N_3908);
nand U4240 (N_4240,N_3882,N_3780);
or U4241 (N_4241,N_3917,N_3806);
nand U4242 (N_4242,N_3759,N_3859);
nor U4243 (N_4243,N_3994,N_3988);
nand U4244 (N_4244,N_3889,N_3772);
and U4245 (N_4245,N_3946,N_3923);
nor U4246 (N_4246,N_3797,N_3830);
and U4247 (N_4247,N_3953,N_3782);
nand U4248 (N_4248,N_3919,N_3782);
nand U4249 (N_4249,N_3961,N_3984);
nor U4250 (N_4250,N_4113,N_4181);
nand U4251 (N_4251,N_4235,N_4156);
nand U4252 (N_4252,N_4141,N_4026);
or U4253 (N_4253,N_4098,N_4065);
and U4254 (N_4254,N_4241,N_4204);
and U4255 (N_4255,N_4202,N_4240);
and U4256 (N_4256,N_4226,N_4243);
nor U4257 (N_4257,N_4110,N_4080);
and U4258 (N_4258,N_4022,N_4219);
xnor U4259 (N_4259,N_4200,N_4155);
nor U4260 (N_4260,N_4099,N_4063);
and U4261 (N_4261,N_4059,N_4143);
nor U4262 (N_4262,N_4034,N_4210);
or U4263 (N_4263,N_4031,N_4159);
nand U4264 (N_4264,N_4029,N_4108);
and U4265 (N_4265,N_4225,N_4051);
xnor U4266 (N_4266,N_4006,N_4162);
nand U4267 (N_4267,N_4238,N_4077);
nand U4268 (N_4268,N_4095,N_4030);
nor U4269 (N_4269,N_4092,N_4045);
or U4270 (N_4270,N_4193,N_4014);
and U4271 (N_4271,N_4061,N_4198);
and U4272 (N_4272,N_4067,N_4245);
xor U4273 (N_4273,N_4154,N_4121);
nand U4274 (N_4274,N_4220,N_4038);
nor U4275 (N_4275,N_4044,N_4184);
or U4276 (N_4276,N_4056,N_4140);
or U4277 (N_4277,N_4179,N_4124);
nor U4278 (N_4278,N_4027,N_4107);
nor U4279 (N_4279,N_4066,N_4015);
nor U4280 (N_4280,N_4187,N_4132);
nor U4281 (N_4281,N_4151,N_4138);
and U4282 (N_4282,N_4091,N_4103);
or U4283 (N_4283,N_4105,N_4192);
nand U4284 (N_4284,N_4131,N_4052);
nor U4285 (N_4285,N_4212,N_4033);
or U4286 (N_4286,N_4088,N_4017);
nand U4287 (N_4287,N_4137,N_4116);
or U4288 (N_4288,N_4188,N_4048);
or U4289 (N_4289,N_4023,N_4157);
nand U4290 (N_4290,N_4201,N_4093);
nor U4291 (N_4291,N_4036,N_4199);
nand U4292 (N_4292,N_4130,N_4094);
and U4293 (N_4293,N_4150,N_4003);
and U4294 (N_4294,N_4142,N_4076);
nand U4295 (N_4295,N_4019,N_4050);
xnor U4296 (N_4296,N_4008,N_4125);
nand U4297 (N_4297,N_4222,N_4106);
nor U4298 (N_4298,N_4046,N_4249);
nand U4299 (N_4299,N_4166,N_4054);
nand U4300 (N_4300,N_4191,N_4170);
or U4301 (N_4301,N_4083,N_4216);
or U4302 (N_4302,N_4004,N_4037);
xor U4303 (N_4303,N_4104,N_4160);
xor U4304 (N_4304,N_4163,N_4224);
nand U4305 (N_4305,N_4028,N_4135);
nor U4306 (N_4306,N_4239,N_4119);
or U4307 (N_4307,N_4176,N_4000);
nor U4308 (N_4308,N_4042,N_4011);
or U4309 (N_4309,N_4089,N_4002);
or U4310 (N_4310,N_4177,N_4069);
and U4311 (N_4311,N_4190,N_4009);
nor U4312 (N_4312,N_4208,N_4161);
nand U4313 (N_4313,N_4115,N_4024);
and U4314 (N_4314,N_4174,N_4172);
nor U4315 (N_4315,N_4248,N_4025);
and U4316 (N_4316,N_4246,N_4182);
xnor U4317 (N_4317,N_4072,N_4085);
nand U4318 (N_4318,N_4207,N_4203);
nand U4319 (N_4319,N_4185,N_4068);
nand U4320 (N_4320,N_4144,N_4139);
or U4321 (N_4321,N_4096,N_4134);
nor U4322 (N_4322,N_4232,N_4169);
and U4323 (N_4323,N_4165,N_4057);
nor U4324 (N_4324,N_4167,N_4087);
nor U4325 (N_4325,N_4237,N_4097);
and U4326 (N_4326,N_4064,N_4229);
or U4327 (N_4327,N_4230,N_4129);
or U4328 (N_4328,N_4039,N_4171);
nand U4329 (N_4329,N_4244,N_4149);
or U4330 (N_4330,N_4058,N_4062);
or U4331 (N_4331,N_4242,N_4227);
nor U4332 (N_4332,N_4111,N_4117);
and U4333 (N_4333,N_4120,N_4205);
nand U4334 (N_4334,N_4211,N_4118);
nor U4335 (N_4335,N_4081,N_4209);
or U4336 (N_4336,N_4128,N_4152);
nand U4337 (N_4337,N_4221,N_4016);
or U4338 (N_4338,N_4082,N_4147);
and U4339 (N_4339,N_4197,N_4136);
nand U4340 (N_4340,N_4041,N_4100);
and U4341 (N_4341,N_4175,N_4234);
or U4342 (N_4342,N_4070,N_4043);
or U4343 (N_4343,N_4173,N_4231);
nor U4344 (N_4344,N_4112,N_4178);
or U4345 (N_4345,N_4233,N_4153);
xor U4346 (N_4346,N_4049,N_4223);
or U4347 (N_4347,N_4047,N_4164);
nand U4348 (N_4348,N_4005,N_4228);
nand U4349 (N_4349,N_4180,N_4020);
or U4350 (N_4350,N_4146,N_4102);
and U4351 (N_4351,N_4018,N_4010);
or U4352 (N_4352,N_4194,N_4122);
and U4353 (N_4353,N_4218,N_4021);
and U4354 (N_4354,N_4079,N_4148);
nand U4355 (N_4355,N_4001,N_4126);
nand U4356 (N_4356,N_4032,N_4007);
nand U4357 (N_4357,N_4078,N_4123);
and U4358 (N_4358,N_4145,N_4012);
and U4359 (N_4359,N_4168,N_4215);
nand U4360 (N_4360,N_4086,N_4040);
and U4361 (N_4361,N_4127,N_4158);
nor U4362 (N_4362,N_4053,N_4109);
and U4363 (N_4363,N_4213,N_4206);
nand U4364 (N_4364,N_4060,N_4084);
nor U4365 (N_4365,N_4195,N_4133);
xor U4366 (N_4366,N_4196,N_4214);
nand U4367 (N_4367,N_4183,N_4090);
or U4368 (N_4368,N_4035,N_4073);
nor U4369 (N_4369,N_4186,N_4074);
nand U4370 (N_4370,N_4247,N_4071);
xor U4371 (N_4371,N_4114,N_4075);
nand U4372 (N_4372,N_4217,N_4013);
nand U4373 (N_4373,N_4101,N_4189);
xor U4374 (N_4374,N_4055,N_4236);
nor U4375 (N_4375,N_4098,N_4188);
nand U4376 (N_4376,N_4046,N_4081);
nand U4377 (N_4377,N_4111,N_4071);
nor U4378 (N_4378,N_4190,N_4013);
and U4379 (N_4379,N_4063,N_4015);
nor U4380 (N_4380,N_4080,N_4042);
nand U4381 (N_4381,N_4060,N_4142);
nand U4382 (N_4382,N_4189,N_4034);
and U4383 (N_4383,N_4009,N_4183);
nor U4384 (N_4384,N_4133,N_4030);
nand U4385 (N_4385,N_4064,N_4041);
nand U4386 (N_4386,N_4210,N_4123);
nor U4387 (N_4387,N_4151,N_4244);
nor U4388 (N_4388,N_4094,N_4087);
and U4389 (N_4389,N_4132,N_4108);
nor U4390 (N_4390,N_4182,N_4003);
nand U4391 (N_4391,N_4168,N_4038);
or U4392 (N_4392,N_4238,N_4112);
and U4393 (N_4393,N_4017,N_4191);
nor U4394 (N_4394,N_4230,N_4080);
or U4395 (N_4395,N_4035,N_4085);
and U4396 (N_4396,N_4088,N_4111);
and U4397 (N_4397,N_4051,N_4221);
or U4398 (N_4398,N_4213,N_4019);
or U4399 (N_4399,N_4210,N_4009);
nor U4400 (N_4400,N_4054,N_4209);
nor U4401 (N_4401,N_4161,N_4103);
nand U4402 (N_4402,N_4074,N_4009);
or U4403 (N_4403,N_4222,N_4066);
or U4404 (N_4404,N_4015,N_4211);
nand U4405 (N_4405,N_4131,N_4222);
and U4406 (N_4406,N_4180,N_4231);
and U4407 (N_4407,N_4056,N_4108);
nand U4408 (N_4408,N_4225,N_4135);
nor U4409 (N_4409,N_4027,N_4039);
nand U4410 (N_4410,N_4212,N_4125);
nor U4411 (N_4411,N_4235,N_4117);
nor U4412 (N_4412,N_4192,N_4063);
and U4413 (N_4413,N_4209,N_4053);
xnor U4414 (N_4414,N_4203,N_4086);
nand U4415 (N_4415,N_4015,N_4093);
and U4416 (N_4416,N_4012,N_4229);
and U4417 (N_4417,N_4205,N_4186);
nand U4418 (N_4418,N_4224,N_4126);
nor U4419 (N_4419,N_4074,N_4235);
and U4420 (N_4420,N_4249,N_4094);
or U4421 (N_4421,N_4235,N_4085);
or U4422 (N_4422,N_4209,N_4004);
nand U4423 (N_4423,N_4207,N_4103);
nor U4424 (N_4424,N_4249,N_4025);
or U4425 (N_4425,N_4167,N_4008);
nand U4426 (N_4426,N_4006,N_4067);
nand U4427 (N_4427,N_4149,N_4051);
xnor U4428 (N_4428,N_4219,N_4125);
nor U4429 (N_4429,N_4147,N_4166);
or U4430 (N_4430,N_4132,N_4061);
nor U4431 (N_4431,N_4033,N_4168);
nor U4432 (N_4432,N_4207,N_4123);
nand U4433 (N_4433,N_4031,N_4122);
nand U4434 (N_4434,N_4230,N_4185);
nor U4435 (N_4435,N_4098,N_4228);
and U4436 (N_4436,N_4246,N_4088);
and U4437 (N_4437,N_4035,N_4054);
and U4438 (N_4438,N_4207,N_4014);
nor U4439 (N_4439,N_4095,N_4235);
nand U4440 (N_4440,N_4043,N_4090);
or U4441 (N_4441,N_4238,N_4176);
or U4442 (N_4442,N_4137,N_4035);
xnor U4443 (N_4443,N_4033,N_4222);
nor U4444 (N_4444,N_4004,N_4232);
nor U4445 (N_4445,N_4095,N_4067);
nor U4446 (N_4446,N_4059,N_4193);
or U4447 (N_4447,N_4154,N_4206);
and U4448 (N_4448,N_4049,N_4242);
and U4449 (N_4449,N_4112,N_4120);
or U4450 (N_4450,N_4156,N_4028);
or U4451 (N_4451,N_4133,N_4209);
or U4452 (N_4452,N_4088,N_4044);
and U4453 (N_4453,N_4151,N_4115);
and U4454 (N_4454,N_4199,N_4029);
nor U4455 (N_4455,N_4072,N_4024);
or U4456 (N_4456,N_4082,N_4244);
or U4457 (N_4457,N_4186,N_4208);
and U4458 (N_4458,N_4009,N_4245);
nor U4459 (N_4459,N_4166,N_4039);
and U4460 (N_4460,N_4205,N_4231);
nor U4461 (N_4461,N_4097,N_4123);
nor U4462 (N_4462,N_4143,N_4174);
nor U4463 (N_4463,N_4183,N_4226);
nand U4464 (N_4464,N_4058,N_4225);
xor U4465 (N_4465,N_4119,N_4156);
nor U4466 (N_4466,N_4123,N_4224);
nand U4467 (N_4467,N_4169,N_4131);
nand U4468 (N_4468,N_4115,N_4219);
and U4469 (N_4469,N_4086,N_4171);
nor U4470 (N_4470,N_4090,N_4078);
nor U4471 (N_4471,N_4152,N_4136);
nand U4472 (N_4472,N_4245,N_4021);
nand U4473 (N_4473,N_4050,N_4214);
nand U4474 (N_4474,N_4176,N_4146);
and U4475 (N_4475,N_4074,N_4140);
or U4476 (N_4476,N_4049,N_4210);
or U4477 (N_4477,N_4207,N_4130);
xor U4478 (N_4478,N_4157,N_4046);
or U4479 (N_4479,N_4190,N_4035);
nand U4480 (N_4480,N_4005,N_4126);
nand U4481 (N_4481,N_4125,N_4032);
or U4482 (N_4482,N_4239,N_4201);
nor U4483 (N_4483,N_4239,N_4085);
or U4484 (N_4484,N_4150,N_4037);
or U4485 (N_4485,N_4244,N_4010);
xor U4486 (N_4486,N_4092,N_4021);
and U4487 (N_4487,N_4049,N_4067);
and U4488 (N_4488,N_4235,N_4037);
and U4489 (N_4489,N_4054,N_4079);
nand U4490 (N_4490,N_4128,N_4221);
nand U4491 (N_4491,N_4066,N_4074);
or U4492 (N_4492,N_4151,N_4032);
nor U4493 (N_4493,N_4113,N_4236);
or U4494 (N_4494,N_4249,N_4221);
nor U4495 (N_4495,N_4126,N_4223);
nand U4496 (N_4496,N_4056,N_4020);
nor U4497 (N_4497,N_4126,N_4085);
and U4498 (N_4498,N_4151,N_4106);
nand U4499 (N_4499,N_4248,N_4084);
nand U4500 (N_4500,N_4307,N_4397);
or U4501 (N_4501,N_4445,N_4409);
nand U4502 (N_4502,N_4317,N_4320);
and U4503 (N_4503,N_4416,N_4434);
and U4504 (N_4504,N_4310,N_4346);
or U4505 (N_4505,N_4414,N_4447);
nand U4506 (N_4506,N_4327,N_4436);
nand U4507 (N_4507,N_4478,N_4396);
nor U4508 (N_4508,N_4257,N_4267);
nor U4509 (N_4509,N_4472,N_4432);
and U4510 (N_4510,N_4334,N_4493);
xnor U4511 (N_4511,N_4328,N_4381);
and U4512 (N_4512,N_4356,N_4344);
and U4513 (N_4513,N_4252,N_4302);
xnor U4514 (N_4514,N_4378,N_4486);
nor U4515 (N_4515,N_4446,N_4311);
xnor U4516 (N_4516,N_4336,N_4287);
xnor U4517 (N_4517,N_4412,N_4401);
or U4518 (N_4518,N_4359,N_4376);
and U4519 (N_4519,N_4384,N_4382);
nand U4520 (N_4520,N_4392,N_4497);
nand U4521 (N_4521,N_4452,N_4329);
and U4522 (N_4522,N_4324,N_4372);
nor U4523 (N_4523,N_4464,N_4460);
nor U4524 (N_4524,N_4348,N_4449);
nand U4525 (N_4525,N_4333,N_4321);
or U4526 (N_4526,N_4484,N_4264);
nor U4527 (N_4527,N_4278,N_4270);
or U4528 (N_4528,N_4255,N_4400);
nand U4529 (N_4529,N_4425,N_4439);
nor U4530 (N_4530,N_4456,N_4413);
nand U4531 (N_4531,N_4479,N_4387);
or U4532 (N_4532,N_4319,N_4315);
nand U4533 (N_4533,N_4351,N_4426);
nor U4534 (N_4534,N_4306,N_4294);
and U4535 (N_4535,N_4305,N_4268);
and U4536 (N_4536,N_4411,N_4337);
xor U4537 (N_4537,N_4471,N_4386);
and U4538 (N_4538,N_4263,N_4345);
nor U4539 (N_4539,N_4448,N_4379);
and U4540 (N_4540,N_4298,N_4314);
xnor U4541 (N_4541,N_4440,N_4459);
nand U4542 (N_4542,N_4364,N_4262);
nand U4543 (N_4543,N_4404,N_4395);
or U4544 (N_4544,N_4466,N_4318);
or U4545 (N_4545,N_4304,N_4398);
and U4546 (N_4546,N_4366,N_4251);
nand U4547 (N_4547,N_4418,N_4431);
nand U4548 (N_4548,N_4303,N_4408);
nand U4549 (N_4549,N_4476,N_4335);
nor U4550 (N_4550,N_4343,N_4483);
nor U4551 (N_4551,N_4290,N_4367);
nand U4552 (N_4552,N_4261,N_4347);
nand U4553 (N_4553,N_4377,N_4374);
or U4554 (N_4554,N_4259,N_4429);
nand U4555 (N_4555,N_4361,N_4465);
and U4556 (N_4556,N_4383,N_4313);
nor U4557 (N_4557,N_4371,N_4453);
nand U4558 (N_4558,N_4326,N_4406);
nor U4559 (N_4559,N_4402,N_4286);
nand U4560 (N_4560,N_4292,N_4389);
and U4561 (N_4561,N_4457,N_4424);
xnor U4562 (N_4562,N_4492,N_4342);
or U4563 (N_4563,N_4325,N_4297);
xnor U4564 (N_4564,N_4481,N_4323);
nor U4565 (N_4565,N_4475,N_4291);
nand U4566 (N_4566,N_4385,N_4300);
nor U4567 (N_4567,N_4288,N_4419);
or U4568 (N_4568,N_4322,N_4357);
and U4569 (N_4569,N_4258,N_4433);
xnor U4570 (N_4570,N_4265,N_4423);
nor U4571 (N_4571,N_4410,N_4394);
nor U4572 (N_4572,N_4271,N_4461);
nand U4573 (N_4573,N_4266,N_4399);
and U4574 (N_4574,N_4390,N_4365);
nand U4575 (N_4575,N_4430,N_4282);
nand U4576 (N_4576,N_4468,N_4438);
nand U4577 (N_4577,N_4280,N_4256);
xnor U4578 (N_4578,N_4380,N_4340);
nor U4579 (N_4579,N_4393,N_4269);
xnor U4580 (N_4580,N_4276,N_4455);
and U4581 (N_4581,N_4308,N_4443);
and U4582 (N_4582,N_4281,N_4353);
or U4583 (N_4583,N_4358,N_4369);
nand U4584 (N_4584,N_4474,N_4415);
or U4585 (N_4585,N_4316,N_4437);
and U4586 (N_4586,N_4373,N_4285);
or U4587 (N_4587,N_4331,N_4469);
xor U4588 (N_4588,N_4442,N_4350);
and U4589 (N_4589,N_4428,N_4421);
nand U4590 (N_4590,N_4289,N_4405);
nand U4591 (N_4591,N_4274,N_4296);
nand U4592 (N_4592,N_4458,N_4467);
and U4593 (N_4593,N_4253,N_4477);
nand U4594 (N_4594,N_4470,N_4283);
nor U4595 (N_4595,N_4463,N_4250);
and U4596 (N_4596,N_4489,N_4352);
nor U4597 (N_4597,N_4272,N_4368);
nor U4598 (N_4598,N_4349,N_4427);
nor U4599 (N_4599,N_4494,N_4355);
nand U4600 (N_4600,N_4444,N_4480);
and U4601 (N_4601,N_4388,N_4339);
or U4602 (N_4602,N_4312,N_4473);
nand U4603 (N_4603,N_4435,N_4417);
nand U4604 (N_4604,N_4488,N_4284);
nor U4605 (N_4605,N_4391,N_4277);
xor U4606 (N_4606,N_4341,N_4332);
nor U4607 (N_4607,N_4330,N_4254);
xnor U4608 (N_4608,N_4370,N_4495);
and U4609 (N_4609,N_4462,N_4275);
nor U4610 (N_4610,N_4420,N_4485);
nor U4611 (N_4611,N_4362,N_4375);
or U4612 (N_4612,N_4422,N_4273);
nor U4613 (N_4613,N_4454,N_4450);
nand U4614 (N_4614,N_4451,N_4403);
nor U4615 (N_4615,N_4299,N_4279);
and U4616 (N_4616,N_4360,N_4482);
or U4617 (N_4617,N_4301,N_4441);
and U4618 (N_4618,N_4309,N_4487);
and U4619 (N_4619,N_4407,N_4490);
nor U4620 (N_4620,N_4295,N_4363);
nor U4621 (N_4621,N_4293,N_4496);
and U4622 (N_4622,N_4491,N_4354);
and U4623 (N_4623,N_4499,N_4260);
and U4624 (N_4624,N_4338,N_4498);
or U4625 (N_4625,N_4432,N_4474);
and U4626 (N_4626,N_4369,N_4273);
and U4627 (N_4627,N_4457,N_4401);
nand U4628 (N_4628,N_4367,N_4287);
nor U4629 (N_4629,N_4368,N_4451);
and U4630 (N_4630,N_4326,N_4477);
nor U4631 (N_4631,N_4419,N_4311);
or U4632 (N_4632,N_4260,N_4365);
or U4633 (N_4633,N_4254,N_4350);
and U4634 (N_4634,N_4286,N_4476);
and U4635 (N_4635,N_4497,N_4408);
nand U4636 (N_4636,N_4440,N_4328);
and U4637 (N_4637,N_4383,N_4331);
nor U4638 (N_4638,N_4482,N_4487);
nor U4639 (N_4639,N_4474,N_4280);
nand U4640 (N_4640,N_4425,N_4302);
nor U4641 (N_4641,N_4336,N_4412);
and U4642 (N_4642,N_4493,N_4329);
xnor U4643 (N_4643,N_4498,N_4276);
nor U4644 (N_4644,N_4322,N_4378);
nand U4645 (N_4645,N_4435,N_4460);
xnor U4646 (N_4646,N_4305,N_4396);
nor U4647 (N_4647,N_4479,N_4469);
and U4648 (N_4648,N_4482,N_4441);
and U4649 (N_4649,N_4281,N_4463);
nand U4650 (N_4650,N_4351,N_4427);
xor U4651 (N_4651,N_4466,N_4281);
nor U4652 (N_4652,N_4254,N_4300);
and U4653 (N_4653,N_4383,N_4256);
or U4654 (N_4654,N_4477,N_4415);
nand U4655 (N_4655,N_4350,N_4483);
or U4656 (N_4656,N_4263,N_4367);
nand U4657 (N_4657,N_4408,N_4444);
nor U4658 (N_4658,N_4412,N_4382);
or U4659 (N_4659,N_4392,N_4269);
or U4660 (N_4660,N_4303,N_4320);
nor U4661 (N_4661,N_4434,N_4422);
xor U4662 (N_4662,N_4253,N_4360);
and U4663 (N_4663,N_4337,N_4371);
and U4664 (N_4664,N_4428,N_4474);
and U4665 (N_4665,N_4258,N_4499);
nor U4666 (N_4666,N_4486,N_4254);
nor U4667 (N_4667,N_4260,N_4342);
nand U4668 (N_4668,N_4455,N_4296);
nand U4669 (N_4669,N_4432,N_4250);
nand U4670 (N_4670,N_4475,N_4324);
and U4671 (N_4671,N_4424,N_4274);
and U4672 (N_4672,N_4337,N_4329);
and U4673 (N_4673,N_4273,N_4353);
nand U4674 (N_4674,N_4444,N_4397);
or U4675 (N_4675,N_4341,N_4292);
or U4676 (N_4676,N_4367,N_4449);
and U4677 (N_4677,N_4433,N_4463);
or U4678 (N_4678,N_4388,N_4295);
nor U4679 (N_4679,N_4284,N_4259);
nor U4680 (N_4680,N_4324,N_4456);
and U4681 (N_4681,N_4324,N_4289);
xor U4682 (N_4682,N_4376,N_4442);
nand U4683 (N_4683,N_4254,N_4371);
or U4684 (N_4684,N_4326,N_4265);
or U4685 (N_4685,N_4325,N_4468);
or U4686 (N_4686,N_4490,N_4480);
nand U4687 (N_4687,N_4466,N_4296);
nand U4688 (N_4688,N_4275,N_4402);
xor U4689 (N_4689,N_4424,N_4268);
or U4690 (N_4690,N_4284,N_4480);
or U4691 (N_4691,N_4332,N_4264);
nor U4692 (N_4692,N_4480,N_4492);
or U4693 (N_4693,N_4460,N_4451);
nor U4694 (N_4694,N_4274,N_4293);
nor U4695 (N_4695,N_4359,N_4264);
nand U4696 (N_4696,N_4373,N_4440);
or U4697 (N_4697,N_4493,N_4326);
nand U4698 (N_4698,N_4382,N_4338);
or U4699 (N_4699,N_4495,N_4417);
nor U4700 (N_4700,N_4272,N_4461);
nor U4701 (N_4701,N_4322,N_4269);
nor U4702 (N_4702,N_4353,N_4473);
xnor U4703 (N_4703,N_4360,N_4271);
and U4704 (N_4704,N_4322,N_4448);
or U4705 (N_4705,N_4271,N_4476);
or U4706 (N_4706,N_4332,N_4345);
and U4707 (N_4707,N_4411,N_4361);
or U4708 (N_4708,N_4266,N_4350);
or U4709 (N_4709,N_4350,N_4434);
nand U4710 (N_4710,N_4271,N_4269);
and U4711 (N_4711,N_4271,N_4327);
and U4712 (N_4712,N_4416,N_4381);
nand U4713 (N_4713,N_4432,N_4351);
nor U4714 (N_4714,N_4308,N_4340);
or U4715 (N_4715,N_4273,N_4346);
or U4716 (N_4716,N_4352,N_4342);
or U4717 (N_4717,N_4457,N_4285);
and U4718 (N_4718,N_4445,N_4316);
nand U4719 (N_4719,N_4431,N_4426);
nand U4720 (N_4720,N_4343,N_4254);
nand U4721 (N_4721,N_4479,N_4498);
xnor U4722 (N_4722,N_4404,N_4430);
or U4723 (N_4723,N_4437,N_4347);
and U4724 (N_4724,N_4420,N_4268);
xor U4725 (N_4725,N_4492,N_4362);
nand U4726 (N_4726,N_4294,N_4290);
xnor U4727 (N_4727,N_4407,N_4260);
nor U4728 (N_4728,N_4441,N_4255);
xnor U4729 (N_4729,N_4356,N_4269);
and U4730 (N_4730,N_4412,N_4483);
or U4731 (N_4731,N_4303,N_4333);
nor U4732 (N_4732,N_4266,N_4432);
or U4733 (N_4733,N_4399,N_4442);
and U4734 (N_4734,N_4377,N_4385);
nand U4735 (N_4735,N_4303,N_4250);
or U4736 (N_4736,N_4338,N_4332);
nor U4737 (N_4737,N_4283,N_4327);
nor U4738 (N_4738,N_4298,N_4261);
nor U4739 (N_4739,N_4389,N_4454);
and U4740 (N_4740,N_4413,N_4384);
and U4741 (N_4741,N_4439,N_4437);
and U4742 (N_4742,N_4271,N_4257);
or U4743 (N_4743,N_4310,N_4459);
nor U4744 (N_4744,N_4398,N_4413);
xnor U4745 (N_4745,N_4469,N_4492);
nand U4746 (N_4746,N_4390,N_4358);
and U4747 (N_4747,N_4416,N_4432);
and U4748 (N_4748,N_4313,N_4386);
nand U4749 (N_4749,N_4452,N_4346);
nor U4750 (N_4750,N_4639,N_4704);
or U4751 (N_4751,N_4724,N_4619);
nand U4752 (N_4752,N_4741,N_4609);
nor U4753 (N_4753,N_4713,N_4682);
or U4754 (N_4754,N_4522,N_4694);
or U4755 (N_4755,N_4562,N_4614);
or U4756 (N_4756,N_4660,N_4630);
nand U4757 (N_4757,N_4645,N_4581);
nor U4758 (N_4758,N_4740,N_4621);
nand U4759 (N_4759,N_4595,N_4561);
nand U4760 (N_4760,N_4612,N_4699);
and U4761 (N_4761,N_4593,N_4571);
nor U4762 (N_4762,N_4610,N_4698);
and U4763 (N_4763,N_4644,N_4517);
or U4764 (N_4764,N_4541,N_4733);
nand U4765 (N_4765,N_4594,N_4606);
and U4766 (N_4766,N_4695,N_4501);
or U4767 (N_4767,N_4693,N_4678);
nand U4768 (N_4768,N_4686,N_4749);
nand U4769 (N_4769,N_4565,N_4563);
nor U4770 (N_4770,N_4586,N_4676);
xor U4771 (N_4771,N_4528,N_4726);
or U4772 (N_4772,N_4714,N_4620);
nand U4773 (N_4773,N_4521,N_4711);
and U4774 (N_4774,N_4533,N_4661);
nor U4775 (N_4775,N_4587,N_4531);
nand U4776 (N_4776,N_4516,N_4723);
nor U4777 (N_4777,N_4654,N_4671);
xnor U4778 (N_4778,N_4657,N_4721);
or U4779 (N_4779,N_4702,N_4582);
or U4780 (N_4780,N_4601,N_4722);
or U4781 (N_4781,N_4575,N_4731);
or U4782 (N_4782,N_4667,N_4748);
nor U4783 (N_4783,N_4534,N_4712);
nor U4784 (N_4784,N_4705,N_4738);
nor U4785 (N_4785,N_4685,N_4503);
or U4786 (N_4786,N_4656,N_4641);
nor U4787 (N_4787,N_4681,N_4546);
nor U4788 (N_4788,N_4734,N_4577);
and U4789 (N_4789,N_4513,N_4732);
nand U4790 (N_4790,N_4636,N_4629);
and U4791 (N_4791,N_4613,N_4692);
xnor U4792 (N_4792,N_4701,N_4728);
and U4793 (N_4793,N_4596,N_4638);
nor U4794 (N_4794,N_4715,N_4616);
xnor U4795 (N_4795,N_4523,N_4525);
nor U4796 (N_4796,N_4649,N_4703);
or U4797 (N_4797,N_4570,N_4555);
nand U4798 (N_4798,N_4739,N_4542);
nand U4799 (N_4799,N_4536,N_4623);
and U4800 (N_4800,N_4684,N_4735);
nor U4801 (N_4801,N_4524,N_4604);
nor U4802 (N_4802,N_4535,N_4743);
nor U4803 (N_4803,N_4668,N_4742);
and U4804 (N_4804,N_4519,N_4674);
and U4805 (N_4805,N_4583,N_4666);
nor U4806 (N_4806,N_4591,N_4709);
and U4807 (N_4807,N_4512,N_4554);
nor U4808 (N_4808,N_4632,N_4653);
xor U4809 (N_4809,N_4574,N_4627);
or U4810 (N_4810,N_4689,N_4706);
nand U4811 (N_4811,N_4505,N_4500);
nand U4812 (N_4812,N_4727,N_4566);
or U4813 (N_4813,N_4502,N_4576);
nand U4814 (N_4814,N_4592,N_4568);
nand U4815 (N_4815,N_4691,N_4696);
or U4816 (N_4816,N_4643,N_4560);
nor U4817 (N_4817,N_4650,N_4746);
and U4818 (N_4818,N_4527,N_4507);
nor U4819 (N_4819,N_4737,N_4633);
nand U4820 (N_4820,N_4646,N_4687);
xor U4821 (N_4821,N_4585,N_4579);
and U4822 (N_4822,N_4677,N_4615);
or U4823 (N_4823,N_4659,N_4572);
xnor U4824 (N_4824,N_4551,N_4611);
nand U4825 (N_4825,N_4506,N_4607);
nor U4826 (N_4826,N_4569,N_4597);
and U4827 (N_4827,N_4635,N_4665);
nand U4828 (N_4828,N_4647,N_4549);
xor U4829 (N_4829,N_4548,N_4637);
or U4830 (N_4830,N_4539,N_4608);
nor U4831 (N_4831,N_4518,N_4618);
and U4832 (N_4832,N_4651,N_4617);
nand U4833 (N_4833,N_4543,N_4710);
and U4834 (N_4834,N_4510,N_4526);
nand U4835 (N_4835,N_4573,N_4547);
and U4836 (N_4836,N_4508,N_4688);
nand U4837 (N_4837,N_4662,N_4590);
or U4838 (N_4838,N_4605,N_4509);
nor U4839 (N_4839,N_4550,N_4652);
nand U4840 (N_4840,N_4603,N_4716);
and U4841 (N_4841,N_4642,N_4669);
nand U4842 (N_4842,N_4558,N_4744);
and U4843 (N_4843,N_4504,N_4663);
nor U4844 (N_4844,N_4624,N_4602);
nand U4845 (N_4845,N_4537,N_4552);
or U4846 (N_4846,N_4600,N_4584);
or U4847 (N_4847,N_4529,N_4559);
or U4848 (N_4848,N_4736,N_4514);
and U4849 (N_4849,N_4628,N_4673);
or U4850 (N_4850,N_4680,N_4707);
nand U4851 (N_4851,N_4717,N_4683);
nor U4852 (N_4852,N_4718,N_4670);
or U4853 (N_4853,N_4530,N_4690);
nor U4854 (N_4854,N_4700,N_4567);
and U4855 (N_4855,N_4511,N_4599);
nor U4856 (N_4856,N_4729,N_4538);
or U4857 (N_4857,N_4578,N_4580);
or U4858 (N_4858,N_4545,N_4520);
and U4859 (N_4859,N_4658,N_4598);
nand U4860 (N_4860,N_4564,N_4664);
nor U4861 (N_4861,N_4544,N_4626);
nand U4862 (N_4862,N_4745,N_4720);
nand U4863 (N_4863,N_4589,N_4747);
xor U4864 (N_4864,N_4515,N_4625);
and U4865 (N_4865,N_4588,N_4675);
nand U4866 (N_4866,N_4634,N_4725);
and U4867 (N_4867,N_4622,N_4532);
nand U4868 (N_4868,N_4655,N_4672);
or U4869 (N_4869,N_4648,N_4631);
nand U4870 (N_4870,N_4556,N_4719);
nand U4871 (N_4871,N_4697,N_4540);
nand U4872 (N_4872,N_4557,N_4679);
nand U4873 (N_4873,N_4640,N_4553);
nor U4874 (N_4874,N_4730,N_4708);
nand U4875 (N_4875,N_4569,N_4578);
nor U4876 (N_4876,N_4635,N_4574);
nand U4877 (N_4877,N_4615,N_4667);
nor U4878 (N_4878,N_4733,N_4634);
or U4879 (N_4879,N_4517,N_4594);
xor U4880 (N_4880,N_4680,N_4682);
nor U4881 (N_4881,N_4684,N_4683);
or U4882 (N_4882,N_4667,N_4588);
xnor U4883 (N_4883,N_4674,N_4734);
nand U4884 (N_4884,N_4593,N_4681);
xnor U4885 (N_4885,N_4712,N_4688);
nor U4886 (N_4886,N_4597,N_4524);
nand U4887 (N_4887,N_4698,N_4595);
or U4888 (N_4888,N_4504,N_4678);
nor U4889 (N_4889,N_4645,N_4579);
nand U4890 (N_4890,N_4519,N_4533);
nand U4891 (N_4891,N_4646,N_4568);
nand U4892 (N_4892,N_4642,N_4564);
nand U4893 (N_4893,N_4656,N_4747);
nor U4894 (N_4894,N_4555,N_4674);
or U4895 (N_4895,N_4541,N_4736);
nor U4896 (N_4896,N_4692,N_4534);
nand U4897 (N_4897,N_4686,N_4651);
and U4898 (N_4898,N_4670,N_4688);
xor U4899 (N_4899,N_4561,N_4632);
xnor U4900 (N_4900,N_4532,N_4587);
and U4901 (N_4901,N_4539,N_4586);
xor U4902 (N_4902,N_4741,N_4696);
and U4903 (N_4903,N_4654,N_4501);
nand U4904 (N_4904,N_4648,N_4558);
and U4905 (N_4905,N_4592,N_4711);
or U4906 (N_4906,N_4595,N_4515);
and U4907 (N_4907,N_4607,N_4531);
nand U4908 (N_4908,N_4551,N_4653);
or U4909 (N_4909,N_4658,N_4657);
nor U4910 (N_4910,N_4639,N_4687);
nand U4911 (N_4911,N_4694,N_4639);
or U4912 (N_4912,N_4702,N_4732);
nand U4913 (N_4913,N_4717,N_4523);
and U4914 (N_4914,N_4576,N_4643);
or U4915 (N_4915,N_4670,N_4619);
nor U4916 (N_4916,N_4602,N_4526);
nand U4917 (N_4917,N_4549,N_4739);
nand U4918 (N_4918,N_4571,N_4629);
and U4919 (N_4919,N_4741,N_4538);
nor U4920 (N_4920,N_4689,N_4569);
or U4921 (N_4921,N_4620,N_4694);
nor U4922 (N_4922,N_4547,N_4733);
nor U4923 (N_4923,N_4734,N_4604);
or U4924 (N_4924,N_4532,N_4507);
nor U4925 (N_4925,N_4549,N_4558);
xor U4926 (N_4926,N_4721,N_4726);
nand U4927 (N_4927,N_4688,N_4536);
nand U4928 (N_4928,N_4695,N_4597);
and U4929 (N_4929,N_4542,N_4575);
nand U4930 (N_4930,N_4549,N_4500);
and U4931 (N_4931,N_4531,N_4563);
and U4932 (N_4932,N_4727,N_4595);
or U4933 (N_4933,N_4686,N_4728);
and U4934 (N_4934,N_4576,N_4709);
xor U4935 (N_4935,N_4673,N_4634);
or U4936 (N_4936,N_4653,N_4673);
nand U4937 (N_4937,N_4578,N_4643);
nand U4938 (N_4938,N_4558,N_4603);
or U4939 (N_4939,N_4571,N_4505);
xor U4940 (N_4940,N_4690,N_4502);
nand U4941 (N_4941,N_4647,N_4603);
xor U4942 (N_4942,N_4541,N_4596);
nor U4943 (N_4943,N_4604,N_4624);
or U4944 (N_4944,N_4721,N_4598);
nor U4945 (N_4945,N_4541,N_4584);
nor U4946 (N_4946,N_4696,N_4736);
and U4947 (N_4947,N_4616,N_4710);
or U4948 (N_4948,N_4747,N_4553);
and U4949 (N_4949,N_4581,N_4546);
xnor U4950 (N_4950,N_4585,N_4588);
nand U4951 (N_4951,N_4574,N_4584);
nor U4952 (N_4952,N_4704,N_4543);
nand U4953 (N_4953,N_4600,N_4627);
nor U4954 (N_4954,N_4575,N_4532);
or U4955 (N_4955,N_4560,N_4506);
and U4956 (N_4956,N_4728,N_4682);
nand U4957 (N_4957,N_4513,N_4736);
xnor U4958 (N_4958,N_4676,N_4660);
or U4959 (N_4959,N_4649,N_4605);
and U4960 (N_4960,N_4677,N_4508);
and U4961 (N_4961,N_4612,N_4506);
or U4962 (N_4962,N_4513,N_4728);
and U4963 (N_4963,N_4722,N_4598);
nor U4964 (N_4964,N_4588,N_4549);
or U4965 (N_4965,N_4539,N_4615);
or U4966 (N_4966,N_4566,N_4542);
and U4967 (N_4967,N_4731,N_4649);
xor U4968 (N_4968,N_4702,N_4655);
and U4969 (N_4969,N_4689,N_4710);
nand U4970 (N_4970,N_4728,N_4678);
nor U4971 (N_4971,N_4550,N_4619);
nand U4972 (N_4972,N_4591,N_4569);
or U4973 (N_4973,N_4630,N_4739);
nand U4974 (N_4974,N_4629,N_4604);
nor U4975 (N_4975,N_4680,N_4573);
nor U4976 (N_4976,N_4686,N_4537);
or U4977 (N_4977,N_4642,N_4615);
or U4978 (N_4978,N_4636,N_4744);
nand U4979 (N_4979,N_4565,N_4645);
nor U4980 (N_4980,N_4620,N_4622);
nor U4981 (N_4981,N_4708,N_4726);
or U4982 (N_4982,N_4518,N_4531);
and U4983 (N_4983,N_4682,N_4502);
or U4984 (N_4984,N_4586,N_4704);
and U4985 (N_4985,N_4511,N_4630);
or U4986 (N_4986,N_4547,N_4503);
xor U4987 (N_4987,N_4546,N_4672);
and U4988 (N_4988,N_4635,N_4568);
and U4989 (N_4989,N_4640,N_4702);
nor U4990 (N_4990,N_4619,N_4707);
nand U4991 (N_4991,N_4579,N_4729);
nand U4992 (N_4992,N_4614,N_4558);
or U4993 (N_4993,N_4578,N_4612);
nor U4994 (N_4994,N_4662,N_4640);
nor U4995 (N_4995,N_4654,N_4560);
and U4996 (N_4996,N_4672,N_4519);
nor U4997 (N_4997,N_4516,N_4586);
nand U4998 (N_4998,N_4633,N_4717);
nand U4999 (N_4999,N_4704,N_4684);
nor U5000 (N_5000,N_4968,N_4786);
nor U5001 (N_5001,N_4815,N_4939);
nand U5002 (N_5002,N_4856,N_4936);
or U5003 (N_5003,N_4987,N_4915);
or U5004 (N_5004,N_4942,N_4959);
and U5005 (N_5005,N_4895,N_4905);
nand U5006 (N_5006,N_4873,N_4876);
or U5007 (N_5007,N_4930,N_4805);
or U5008 (N_5008,N_4871,N_4765);
and U5009 (N_5009,N_4864,N_4977);
nand U5010 (N_5010,N_4878,N_4853);
xnor U5011 (N_5011,N_4940,N_4751);
and U5012 (N_5012,N_4798,N_4830);
or U5013 (N_5013,N_4803,N_4778);
or U5014 (N_5014,N_4902,N_4833);
and U5015 (N_5015,N_4956,N_4842);
nor U5016 (N_5016,N_4789,N_4850);
and U5017 (N_5017,N_4886,N_4870);
or U5018 (N_5018,N_4756,N_4843);
and U5019 (N_5019,N_4967,N_4800);
or U5020 (N_5020,N_4837,N_4901);
nor U5021 (N_5021,N_4891,N_4937);
nand U5022 (N_5022,N_4954,N_4929);
nand U5023 (N_5023,N_4770,N_4923);
nand U5024 (N_5024,N_4863,N_4974);
or U5025 (N_5025,N_4917,N_4866);
xnor U5026 (N_5026,N_4875,N_4962);
or U5027 (N_5027,N_4797,N_4861);
nor U5028 (N_5028,N_4801,N_4963);
or U5029 (N_5029,N_4951,N_4918);
nand U5030 (N_5030,N_4986,N_4855);
and U5031 (N_5031,N_4818,N_4958);
or U5032 (N_5032,N_4980,N_4758);
and U5033 (N_5033,N_4872,N_4966);
or U5034 (N_5034,N_4907,N_4900);
nor U5035 (N_5035,N_4828,N_4976);
nand U5036 (N_5036,N_4788,N_4916);
nor U5037 (N_5037,N_4931,N_4983);
and U5038 (N_5038,N_4944,N_4793);
nor U5039 (N_5039,N_4946,N_4911);
nand U5040 (N_5040,N_4825,N_4846);
or U5041 (N_5041,N_4972,N_4919);
and U5042 (N_5042,N_4964,N_4928);
and U5043 (N_5043,N_4898,N_4945);
nor U5044 (N_5044,N_4988,N_4948);
or U5045 (N_5045,N_4883,N_4978);
nand U5046 (N_5046,N_4808,N_4790);
nor U5047 (N_5047,N_4985,N_4762);
and U5048 (N_5048,N_4764,N_4840);
nand U5049 (N_5049,N_4781,N_4971);
or U5050 (N_5050,N_4995,N_4975);
and U5051 (N_5051,N_4777,N_4841);
nand U5052 (N_5052,N_4812,N_4903);
nor U5053 (N_5053,N_4949,N_4816);
and U5054 (N_5054,N_4953,N_4994);
and U5055 (N_5055,N_4992,N_4938);
nor U5056 (N_5056,N_4854,N_4965);
xnor U5057 (N_5057,N_4769,N_4784);
or U5058 (N_5058,N_4943,N_4998);
nor U5059 (N_5059,N_4970,N_4759);
and U5060 (N_5060,N_4822,N_4757);
nor U5061 (N_5061,N_4997,N_4750);
and U5062 (N_5062,N_4912,N_4982);
or U5063 (N_5063,N_4981,N_4922);
nor U5064 (N_5064,N_4804,N_4783);
nand U5065 (N_5065,N_4823,N_4831);
or U5066 (N_5066,N_4859,N_4862);
xor U5067 (N_5067,N_4924,N_4882);
or U5068 (N_5068,N_4814,N_4774);
or U5069 (N_5069,N_4791,N_4827);
and U5070 (N_5070,N_4835,N_4889);
or U5071 (N_5071,N_4897,N_4752);
or U5072 (N_5072,N_4910,N_4755);
and U5073 (N_5073,N_4754,N_4847);
and U5074 (N_5074,N_4996,N_4807);
xnor U5075 (N_5075,N_4799,N_4858);
nand U5076 (N_5076,N_4780,N_4773);
nand U5077 (N_5077,N_4969,N_4874);
and U5078 (N_5078,N_4810,N_4979);
and U5079 (N_5079,N_4955,N_4787);
or U5080 (N_5080,N_4796,N_4957);
nand U5081 (N_5081,N_4834,N_4921);
xnor U5082 (N_5082,N_4826,N_4961);
xor U5083 (N_5083,N_4806,N_4884);
nor U5084 (N_5084,N_4999,N_4868);
nor U5085 (N_5085,N_4887,N_4989);
nor U5086 (N_5086,N_4893,N_4768);
nor U5087 (N_5087,N_4851,N_4824);
and U5088 (N_5088,N_4888,N_4771);
and U5089 (N_5089,N_4792,N_4811);
nor U5090 (N_5090,N_4894,N_4821);
and U5091 (N_5091,N_4817,N_4760);
or U5092 (N_5092,N_4899,N_4785);
or U5093 (N_5093,N_4795,N_4775);
nor U5094 (N_5094,N_4913,N_4947);
or U5095 (N_5095,N_4926,N_4932);
or U5096 (N_5096,N_4766,N_4819);
xor U5097 (N_5097,N_4952,N_4925);
xnor U5098 (N_5098,N_4839,N_4935);
nor U5099 (N_5099,N_4906,N_4767);
or U5100 (N_5100,N_4753,N_4860);
nand U5101 (N_5101,N_4761,N_4869);
nor U5102 (N_5102,N_4927,N_4794);
xnor U5103 (N_5103,N_4877,N_4896);
nand U5104 (N_5104,N_4904,N_4867);
nor U5105 (N_5105,N_4908,N_4829);
nor U5106 (N_5106,N_4885,N_4802);
nor U5107 (N_5107,N_4838,N_4832);
and U5108 (N_5108,N_4984,N_4934);
and U5109 (N_5109,N_4836,N_4772);
and U5110 (N_5110,N_4892,N_4865);
or U5111 (N_5111,N_4845,N_4782);
nand U5112 (N_5112,N_4857,N_4881);
or U5113 (N_5113,N_4991,N_4993);
and U5114 (N_5114,N_4909,N_4920);
and U5115 (N_5115,N_4941,N_4933);
nand U5116 (N_5116,N_4914,N_4779);
and U5117 (N_5117,N_4813,N_4776);
nand U5118 (N_5118,N_4990,N_4879);
or U5119 (N_5119,N_4848,N_4849);
nor U5120 (N_5120,N_4950,N_4890);
or U5121 (N_5121,N_4763,N_4880);
xor U5122 (N_5122,N_4820,N_4852);
nand U5123 (N_5123,N_4960,N_4809);
nor U5124 (N_5124,N_4973,N_4844);
xor U5125 (N_5125,N_4964,N_4949);
and U5126 (N_5126,N_4911,N_4872);
nor U5127 (N_5127,N_4811,N_4835);
nand U5128 (N_5128,N_4962,N_4770);
or U5129 (N_5129,N_4855,N_4774);
and U5130 (N_5130,N_4810,N_4956);
xnor U5131 (N_5131,N_4821,N_4965);
nand U5132 (N_5132,N_4961,N_4827);
nand U5133 (N_5133,N_4803,N_4843);
xor U5134 (N_5134,N_4873,N_4923);
and U5135 (N_5135,N_4913,N_4776);
nand U5136 (N_5136,N_4934,N_4948);
xnor U5137 (N_5137,N_4836,N_4834);
and U5138 (N_5138,N_4807,N_4969);
or U5139 (N_5139,N_4970,N_4979);
nor U5140 (N_5140,N_4867,N_4812);
and U5141 (N_5141,N_4918,N_4899);
nor U5142 (N_5142,N_4834,N_4787);
and U5143 (N_5143,N_4856,N_4976);
nor U5144 (N_5144,N_4994,N_4819);
or U5145 (N_5145,N_4810,N_4771);
nor U5146 (N_5146,N_4848,N_4840);
or U5147 (N_5147,N_4776,N_4832);
nor U5148 (N_5148,N_4773,N_4817);
xor U5149 (N_5149,N_4873,N_4981);
nand U5150 (N_5150,N_4965,N_4865);
nor U5151 (N_5151,N_4754,N_4892);
or U5152 (N_5152,N_4995,N_4876);
nor U5153 (N_5153,N_4798,N_4881);
and U5154 (N_5154,N_4877,N_4954);
nor U5155 (N_5155,N_4968,N_4909);
or U5156 (N_5156,N_4808,N_4861);
xor U5157 (N_5157,N_4900,N_4761);
nor U5158 (N_5158,N_4995,N_4751);
and U5159 (N_5159,N_4870,N_4803);
nand U5160 (N_5160,N_4956,N_4780);
nor U5161 (N_5161,N_4898,N_4885);
nand U5162 (N_5162,N_4991,N_4952);
xor U5163 (N_5163,N_4751,N_4882);
nand U5164 (N_5164,N_4955,N_4841);
and U5165 (N_5165,N_4813,N_4847);
nand U5166 (N_5166,N_4848,N_4828);
and U5167 (N_5167,N_4978,N_4783);
or U5168 (N_5168,N_4753,N_4931);
nor U5169 (N_5169,N_4833,N_4779);
nand U5170 (N_5170,N_4986,N_4954);
or U5171 (N_5171,N_4899,N_4846);
nand U5172 (N_5172,N_4789,N_4794);
or U5173 (N_5173,N_4949,N_4934);
nor U5174 (N_5174,N_4921,N_4933);
nor U5175 (N_5175,N_4936,N_4916);
or U5176 (N_5176,N_4964,N_4858);
nor U5177 (N_5177,N_4810,N_4934);
nand U5178 (N_5178,N_4903,N_4940);
nor U5179 (N_5179,N_4803,N_4836);
or U5180 (N_5180,N_4765,N_4847);
nand U5181 (N_5181,N_4880,N_4817);
nor U5182 (N_5182,N_4839,N_4761);
or U5183 (N_5183,N_4970,N_4961);
nor U5184 (N_5184,N_4993,N_4870);
and U5185 (N_5185,N_4771,N_4908);
nor U5186 (N_5186,N_4994,N_4956);
and U5187 (N_5187,N_4877,N_4936);
and U5188 (N_5188,N_4955,N_4930);
or U5189 (N_5189,N_4805,N_4994);
or U5190 (N_5190,N_4885,N_4962);
nand U5191 (N_5191,N_4944,N_4791);
and U5192 (N_5192,N_4772,N_4944);
nor U5193 (N_5193,N_4866,N_4893);
or U5194 (N_5194,N_4817,N_4992);
xor U5195 (N_5195,N_4839,N_4868);
nand U5196 (N_5196,N_4897,N_4905);
xor U5197 (N_5197,N_4808,N_4974);
nand U5198 (N_5198,N_4844,N_4903);
nand U5199 (N_5199,N_4810,N_4790);
nand U5200 (N_5200,N_4872,N_4915);
nor U5201 (N_5201,N_4924,N_4783);
nand U5202 (N_5202,N_4985,N_4915);
nor U5203 (N_5203,N_4945,N_4750);
or U5204 (N_5204,N_4946,N_4904);
nand U5205 (N_5205,N_4884,N_4803);
nor U5206 (N_5206,N_4823,N_4915);
or U5207 (N_5207,N_4878,N_4941);
nor U5208 (N_5208,N_4953,N_4855);
and U5209 (N_5209,N_4756,N_4832);
nor U5210 (N_5210,N_4789,N_4802);
xor U5211 (N_5211,N_4898,N_4878);
or U5212 (N_5212,N_4760,N_4967);
or U5213 (N_5213,N_4794,N_4969);
nor U5214 (N_5214,N_4982,N_4779);
or U5215 (N_5215,N_4779,N_4867);
xnor U5216 (N_5216,N_4902,N_4874);
or U5217 (N_5217,N_4873,N_4934);
xnor U5218 (N_5218,N_4942,N_4966);
nand U5219 (N_5219,N_4870,N_4750);
nor U5220 (N_5220,N_4877,N_4853);
nor U5221 (N_5221,N_4889,N_4918);
xor U5222 (N_5222,N_4966,N_4772);
nor U5223 (N_5223,N_4866,N_4814);
or U5224 (N_5224,N_4857,N_4959);
and U5225 (N_5225,N_4797,N_4758);
nand U5226 (N_5226,N_4949,N_4930);
nor U5227 (N_5227,N_4946,N_4780);
or U5228 (N_5228,N_4870,N_4987);
and U5229 (N_5229,N_4958,N_4845);
nor U5230 (N_5230,N_4971,N_4790);
xor U5231 (N_5231,N_4987,N_4883);
nand U5232 (N_5232,N_4954,N_4997);
or U5233 (N_5233,N_4857,N_4873);
nand U5234 (N_5234,N_4767,N_4924);
and U5235 (N_5235,N_4794,N_4865);
or U5236 (N_5236,N_4894,N_4805);
nand U5237 (N_5237,N_4937,N_4893);
nor U5238 (N_5238,N_4912,N_4756);
and U5239 (N_5239,N_4868,N_4895);
and U5240 (N_5240,N_4936,N_4774);
or U5241 (N_5241,N_4885,N_4881);
nand U5242 (N_5242,N_4810,N_4762);
or U5243 (N_5243,N_4757,N_4967);
nand U5244 (N_5244,N_4836,N_4992);
nand U5245 (N_5245,N_4866,N_4997);
and U5246 (N_5246,N_4778,N_4918);
nand U5247 (N_5247,N_4902,N_4883);
nor U5248 (N_5248,N_4951,N_4787);
nand U5249 (N_5249,N_4821,N_4950);
nor U5250 (N_5250,N_5242,N_5083);
nand U5251 (N_5251,N_5012,N_5247);
nand U5252 (N_5252,N_5137,N_5026);
nor U5253 (N_5253,N_5199,N_5087);
nand U5254 (N_5254,N_5148,N_5196);
and U5255 (N_5255,N_5176,N_5145);
nor U5256 (N_5256,N_5002,N_5102);
nand U5257 (N_5257,N_5014,N_5107);
nand U5258 (N_5258,N_5179,N_5141);
or U5259 (N_5259,N_5213,N_5139);
or U5260 (N_5260,N_5001,N_5010);
nand U5261 (N_5261,N_5067,N_5146);
xor U5262 (N_5262,N_5025,N_5097);
xnor U5263 (N_5263,N_5206,N_5129);
nand U5264 (N_5264,N_5197,N_5017);
nand U5265 (N_5265,N_5086,N_5153);
and U5266 (N_5266,N_5043,N_5122);
and U5267 (N_5267,N_5200,N_5155);
and U5268 (N_5268,N_5249,N_5223);
and U5269 (N_5269,N_5121,N_5116);
xor U5270 (N_5270,N_5073,N_5236);
nand U5271 (N_5271,N_5229,N_5050);
nand U5272 (N_5272,N_5100,N_5019);
or U5273 (N_5273,N_5047,N_5165);
or U5274 (N_5274,N_5127,N_5149);
or U5275 (N_5275,N_5048,N_5088);
nor U5276 (N_5276,N_5118,N_5140);
or U5277 (N_5277,N_5066,N_5074);
and U5278 (N_5278,N_5228,N_5160);
nor U5279 (N_5279,N_5104,N_5241);
and U5280 (N_5280,N_5054,N_5233);
nand U5281 (N_5281,N_5248,N_5150);
or U5282 (N_5282,N_5089,N_5082);
nand U5283 (N_5283,N_5027,N_5077);
xor U5284 (N_5284,N_5167,N_5243);
nand U5285 (N_5285,N_5235,N_5037);
and U5286 (N_5286,N_5214,N_5175);
nor U5287 (N_5287,N_5022,N_5065);
and U5288 (N_5288,N_5057,N_5166);
nand U5289 (N_5289,N_5171,N_5080);
nor U5290 (N_5290,N_5071,N_5177);
and U5291 (N_5291,N_5240,N_5103);
and U5292 (N_5292,N_5041,N_5046);
nand U5293 (N_5293,N_5062,N_5231);
nand U5294 (N_5294,N_5000,N_5207);
or U5295 (N_5295,N_5098,N_5044);
nand U5296 (N_5296,N_5009,N_5090);
nand U5297 (N_5297,N_5099,N_5034);
or U5298 (N_5298,N_5081,N_5115);
nor U5299 (N_5299,N_5004,N_5070);
and U5300 (N_5300,N_5016,N_5186);
nand U5301 (N_5301,N_5030,N_5072);
nor U5302 (N_5302,N_5052,N_5126);
and U5303 (N_5303,N_5079,N_5021);
nand U5304 (N_5304,N_5128,N_5239);
nand U5305 (N_5305,N_5147,N_5205);
nor U5306 (N_5306,N_5219,N_5131);
nor U5307 (N_5307,N_5192,N_5244);
and U5308 (N_5308,N_5018,N_5212);
nor U5309 (N_5309,N_5174,N_5216);
and U5310 (N_5310,N_5156,N_5020);
xnor U5311 (N_5311,N_5185,N_5078);
nand U5312 (N_5312,N_5005,N_5181);
or U5313 (N_5313,N_5180,N_5028);
nor U5314 (N_5314,N_5188,N_5217);
or U5315 (N_5315,N_5084,N_5218);
nand U5316 (N_5316,N_5003,N_5198);
nor U5317 (N_5317,N_5093,N_5201);
nor U5318 (N_5318,N_5096,N_5133);
and U5319 (N_5319,N_5068,N_5006);
or U5320 (N_5320,N_5036,N_5125);
nand U5321 (N_5321,N_5164,N_5045);
and U5322 (N_5322,N_5193,N_5151);
nor U5323 (N_5323,N_5210,N_5245);
nand U5324 (N_5324,N_5130,N_5161);
nand U5325 (N_5325,N_5120,N_5094);
or U5326 (N_5326,N_5154,N_5226);
or U5327 (N_5327,N_5106,N_5169);
and U5328 (N_5328,N_5013,N_5222);
or U5329 (N_5329,N_5195,N_5060);
nor U5330 (N_5330,N_5039,N_5112);
nand U5331 (N_5331,N_5110,N_5234);
nor U5332 (N_5332,N_5113,N_5051);
xor U5333 (N_5333,N_5095,N_5038);
nand U5334 (N_5334,N_5191,N_5172);
nor U5335 (N_5335,N_5237,N_5015);
or U5336 (N_5336,N_5055,N_5049);
or U5337 (N_5337,N_5033,N_5170);
and U5338 (N_5338,N_5183,N_5064);
nor U5339 (N_5339,N_5029,N_5238);
nand U5340 (N_5340,N_5076,N_5187);
or U5341 (N_5341,N_5159,N_5117);
nand U5342 (N_5342,N_5230,N_5123);
nand U5343 (N_5343,N_5132,N_5053);
nor U5344 (N_5344,N_5042,N_5152);
and U5345 (N_5345,N_5109,N_5190);
and U5346 (N_5346,N_5246,N_5056);
xor U5347 (N_5347,N_5158,N_5202);
nor U5348 (N_5348,N_5135,N_5142);
and U5349 (N_5349,N_5227,N_5136);
and U5350 (N_5350,N_5144,N_5111);
or U5351 (N_5351,N_5085,N_5203);
xor U5352 (N_5352,N_5220,N_5189);
nand U5353 (N_5353,N_5208,N_5225);
or U5354 (N_5354,N_5091,N_5092);
or U5355 (N_5355,N_5173,N_5163);
xor U5356 (N_5356,N_5209,N_5023);
nand U5357 (N_5357,N_5162,N_5105);
xnor U5358 (N_5358,N_5178,N_5011);
and U5359 (N_5359,N_5024,N_5182);
nor U5360 (N_5360,N_5134,N_5204);
xor U5361 (N_5361,N_5143,N_5008);
and U5362 (N_5362,N_5032,N_5138);
nand U5363 (N_5363,N_5101,N_5232);
and U5364 (N_5364,N_5215,N_5194);
nor U5365 (N_5365,N_5211,N_5124);
or U5366 (N_5366,N_5108,N_5035);
nor U5367 (N_5367,N_5119,N_5221);
or U5368 (N_5368,N_5061,N_5069);
and U5369 (N_5369,N_5114,N_5063);
nor U5370 (N_5370,N_5040,N_5059);
nand U5371 (N_5371,N_5168,N_5157);
nand U5372 (N_5372,N_5184,N_5224);
or U5373 (N_5373,N_5075,N_5007);
nor U5374 (N_5374,N_5031,N_5058);
or U5375 (N_5375,N_5044,N_5220);
nand U5376 (N_5376,N_5018,N_5175);
xor U5377 (N_5377,N_5211,N_5076);
xor U5378 (N_5378,N_5195,N_5132);
nor U5379 (N_5379,N_5061,N_5148);
and U5380 (N_5380,N_5193,N_5090);
or U5381 (N_5381,N_5202,N_5151);
nand U5382 (N_5382,N_5074,N_5029);
and U5383 (N_5383,N_5229,N_5179);
nor U5384 (N_5384,N_5037,N_5133);
nand U5385 (N_5385,N_5039,N_5119);
xor U5386 (N_5386,N_5118,N_5012);
or U5387 (N_5387,N_5071,N_5173);
nor U5388 (N_5388,N_5115,N_5143);
and U5389 (N_5389,N_5080,N_5031);
and U5390 (N_5390,N_5101,N_5235);
nor U5391 (N_5391,N_5130,N_5177);
nand U5392 (N_5392,N_5003,N_5168);
and U5393 (N_5393,N_5038,N_5099);
nor U5394 (N_5394,N_5238,N_5230);
and U5395 (N_5395,N_5039,N_5051);
xor U5396 (N_5396,N_5015,N_5177);
or U5397 (N_5397,N_5228,N_5067);
xnor U5398 (N_5398,N_5187,N_5015);
nand U5399 (N_5399,N_5204,N_5016);
and U5400 (N_5400,N_5156,N_5150);
nor U5401 (N_5401,N_5146,N_5228);
and U5402 (N_5402,N_5202,N_5065);
or U5403 (N_5403,N_5150,N_5247);
nor U5404 (N_5404,N_5133,N_5197);
xor U5405 (N_5405,N_5066,N_5235);
nand U5406 (N_5406,N_5122,N_5201);
and U5407 (N_5407,N_5209,N_5217);
or U5408 (N_5408,N_5058,N_5070);
nand U5409 (N_5409,N_5185,N_5028);
xor U5410 (N_5410,N_5230,N_5218);
and U5411 (N_5411,N_5196,N_5015);
xor U5412 (N_5412,N_5154,N_5013);
nor U5413 (N_5413,N_5190,N_5072);
nor U5414 (N_5414,N_5074,N_5062);
nor U5415 (N_5415,N_5035,N_5185);
or U5416 (N_5416,N_5082,N_5087);
nand U5417 (N_5417,N_5206,N_5211);
nor U5418 (N_5418,N_5233,N_5101);
and U5419 (N_5419,N_5075,N_5194);
nand U5420 (N_5420,N_5057,N_5034);
and U5421 (N_5421,N_5118,N_5029);
nand U5422 (N_5422,N_5142,N_5177);
nor U5423 (N_5423,N_5099,N_5220);
nand U5424 (N_5424,N_5221,N_5030);
or U5425 (N_5425,N_5122,N_5249);
xnor U5426 (N_5426,N_5153,N_5213);
and U5427 (N_5427,N_5224,N_5066);
nand U5428 (N_5428,N_5194,N_5096);
and U5429 (N_5429,N_5071,N_5124);
nand U5430 (N_5430,N_5088,N_5169);
nor U5431 (N_5431,N_5084,N_5134);
nand U5432 (N_5432,N_5114,N_5026);
nor U5433 (N_5433,N_5031,N_5093);
or U5434 (N_5434,N_5084,N_5002);
nand U5435 (N_5435,N_5213,N_5009);
or U5436 (N_5436,N_5228,N_5225);
or U5437 (N_5437,N_5053,N_5193);
nor U5438 (N_5438,N_5114,N_5220);
nand U5439 (N_5439,N_5023,N_5188);
nor U5440 (N_5440,N_5158,N_5052);
or U5441 (N_5441,N_5190,N_5060);
nor U5442 (N_5442,N_5004,N_5022);
nor U5443 (N_5443,N_5054,N_5026);
and U5444 (N_5444,N_5117,N_5221);
nand U5445 (N_5445,N_5230,N_5228);
or U5446 (N_5446,N_5114,N_5076);
or U5447 (N_5447,N_5015,N_5046);
or U5448 (N_5448,N_5147,N_5021);
nand U5449 (N_5449,N_5141,N_5056);
and U5450 (N_5450,N_5180,N_5002);
nor U5451 (N_5451,N_5229,N_5088);
or U5452 (N_5452,N_5067,N_5240);
nor U5453 (N_5453,N_5242,N_5080);
nor U5454 (N_5454,N_5114,N_5109);
xnor U5455 (N_5455,N_5033,N_5184);
or U5456 (N_5456,N_5090,N_5080);
or U5457 (N_5457,N_5042,N_5097);
xor U5458 (N_5458,N_5114,N_5187);
and U5459 (N_5459,N_5119,N_5205);
nor U5460 (N_5460,N_5010,N_5096);
nand U5461 (N_5461,N_5036,N_5038);
or U5462 (N_5462,N_5224,N_5206);
or U5463 (N_5463,N_5002,N_5052);
and U5464 (N_5464,N_5153,N_5081);
xnor U5465 (N_5465,N_5183,N_5195);
nor U5466 (N_5466,N_5222,N_5061);
nor U5467 (N_5467,N_5191,N_5023);
or U5468 (N_5468,N_5079,N_5164);
or U5469 (N_5469,N_5248,N_5109);
and U5470 (N_5470,N_5202,N_5078);
xnor U5471 (N_5471,N_5121,N_5053);
and U5472 (N_5472,N_5094,N_5025);
or U5473 (N_5473,N_5177,N_5145);
nand U5474 (N_5474,N_5201,N_5131);
or U5475 (N_5475,N_5003,N_5055);
and U5476 (N_5476,N_5195,N_5202);
and U5477 (N_5477,N_5219,N_5007);
and U5478 (N_5478,N_5185,N_5060);
and U5479 (N_5479,N_5160,N_5081);
nor U5480 (N_5480,N_5209,N_5222);
or U5481 (N_5481,N_5029,N_5135);
nor U5482 (N_5482,N_5110,N_5161);
or U5483 (N_5483,N_5212,N_5232);
or U5484 (N_5484,N_5224,N_5021);
or U5485 (N_5485,N_5019,N_5039);
or U5486 (N_5486,N_5166,N_5061);
nand U5487 (N_5487,N_5022,N_5106);
nor U5488 (N_5488,N_5214,N_5228);
nor U5489 (N_5489,N_5202,N_5168);
nand U5490 (N_5490,N_5085,N_5139);
or U5491 (N_5491,N_5234,N_5231);
and U5492 (N_5492,N_5121,N_5154);
nor U5493 (N_5493,N_5104,N_5146);
and U5494 (N_5494,N_5206,N_5135);
or U5495 (N_5495,N_5236,N_5149);
or U5496 (N_5496,N_5204,N_5193);
xor U5497 (N_5497,N_5249,N_5211);
nor U5498 (N_5498,N_5209,N_5035);
nand U5499 (N_5499,N_5174,N_5166);
nand U5500 (N_5500,N_5423,N_5326);
nand U5501 (N_5501,N_5364,N_5468);
nand U5502 (N_5502,N_5320,N_5370);
or U5503 (N_5503,N_5285,N_5410);
nor U5504 (N_5504,N_5475,N_5389);
nand U5505 (N_5505,N_5385,N_5388);
nor U5506 (N_5506,N_5278,N_5470);
nand U5507 (N_5507,N_5454,N_5315);
or U5508 (N_5508,N_5374,N_5260);
or U5509 (N_5509,N_5467,N_5484);
nor U5510 (N_5510,N_5395,N_5466);
nor U5511 (N_5511,N_5310,N_5299);
and U5512 (N_5512,N_5400,N_5489);
nor U5513 (N_5513,N_5426,N_5443);
and U5514 (N_5514,N_5486,N_5456);
or U5515 (N_5515,N_5396,N_5402);
or U5516 (N_5516,N_5414,N_5305);
or U5517 (N_5517,N_5386,N_5405);
or U5518 (N_5518,N_5322,N_5340);
nor U5519 (N_5519,N_5350,N_5252);
and U5520 (N_5520,N_5265,N_5452);
nor U5521 (N_5521,N_5391,N_5499);
nand U5522 (N_5522,N_5341,N_5330);
and U5523 (N_5523,N_5494,N_5301);
and U5524 (N_5524,N_5349,N_5453);
or U5525 (N_5525,N_5383,N_5417);
and U5526 (N_5526,N_5290,N_5259);
nor U5527 (N_5527,N_5471,N_5424);
nand U5528 (N_5528,N_5266,N_5380);
and U5529 (N_5529,N_5331,N_5309);
nor U5530 (N_5530,N_5358,N_5427);
and U5531 (N_5531,N_5455,N_5273);
nand U5532 (N_5532,N_5447,N_5367);
and U5533 (N_5533,N_5438,N_5378);
or U5534 (N_5534,N_5277,N_5377);
and U5535 (N_5535,N_5345,N_5360);
and U5536 (N_5536,N_5495,N_5291);
or U5537 (N_5537,N_5477,N_5419);
or U5538 (N_5538,N_5304,N_5382);
and U5539 (N_5539,N_5463,N_5297);
and U5540 (N_5540,N_5462,N_5413);
nand U5541 (N_5541,N_5319,N_5444);
nand U5542 (N_5542,N_5250,N_5284);
and U5543 (N_5543,N_5296,N_5357);
or U5544 (N_5544,N_5436,N_5256);
or U5545 (N_5545,N_5254,N_5399);
nor U5546 (N_5546,N_5381,N_5437);
nor U5547 (N_5547,N_5448,N_5488);
nand U5548 (N_5548,N_5253,N_5434);
nor U5549 (N_5549,N_5482,N_5406);
nor U5550 (N_5550,N_5450,N_5282);
and U5551 (N_5551,N_5420,N_5473);
or U5552 (N_5552,N_5474,N_5298);
and U5553 (N_5553,N_5283,N_5441);
nand U5554 (N_5554,N_5268,N_5408);
or U5555 (N_5555,N_5401,N_5311);
nor U5556 (N_5556,N_5257,N_5416);
nand U5557 (N_5557,N_5303,N_5449);
nand U5558 (N_5558,N_5313,N_5440);
and U5559 (N_5559,N_5365,N_5348);
xnor U5560 (N_5560,N_5371,N_5464);
nor U5561 (N_5561,N_5457,N_5289);
or U5562 (N_5562,N_5336,N_5317);
nand U5563 (N_5563,N_5433,N_5276);
xnor U5564 (N_5564,N_5342,N_5407);
xor U5565 (N_5565,N_5366,N_5429);
and U5566 (N_5566,N_5460,N_5267);
nand U5567 (N_5567,N_5498,N_5262);
xnor U5568 (N_5568,N_5432,N_5258);
nor U5569 (N_5569,N_5411,N_5431);
nor U5570 (N_5570,N_5343,N_5430);
nand U5571 (N_5571,N_5355,N_5392);
and U5572 (N_5572,N_5487,N_5333);
nand U5573 (N_5573,N_5393,N_5275);
xnor U5574 (N_5574,N_5479,N_5269);
xor U5575 (N_5575,N_5483,N_5264);
nor U5576 (N_5576,N_5497,N_5492);
and U5577 (N_5577,N_5325,N_5481);
nor U5578 (N_5578,N_5485,N_5314);
xor U5579 (N_5579,N_5270,N_5476);
nand U5580 (N_5580,N_5422,N_5318);
xnor U5581 (N_5581,N_5316,N_5327);
xor U5582 (N_5582,N_5403,N_5261);
and U5583 (N_5583,N_5306,N_5324);
or U5584 (N_5584,N_5287,N_5375);
and U5585 (N_5585,N_5361,N_5472);
xnor U5586 (N_5586,N_5335,N_5329);
nor U5587 (N_5587,N_5496,N_5384);
nand U5588 (N_5588,N_5478,N_5480);
nand U5589 (N_5589,N_5451,N_5465);
nor U5590 (N_5590,N_5363,N_5308);
nor U5591 (N_5591,N_5369,N_5294);
nor U5592 (N_5592,N_5387,N_5442);
or U5593 (N_5593,N_5286,N_5404);
nand U5594 (N_5594,N_5373,N_5354);
nor U5595 (N_5595,N_5418,N_5271);
xor U5596 (N_5596,N_5409,N_5255);
nor U5597 (N_5597,N_5293,N_5272);
or U5598 (N_5598,N_5288,N_5439);
nor U5599 (N_5599,N_5362,N_5263);
nor U5600 (N_5600,N_5328,N_5353);
and U5601 (N_5601,N_5300,N_5459);
nand U5602 (N_5602,N_5412,N_5394);
and U5603 (N_5603,N_5415,N_5428);
nand U5604 (N_5604,N_5425,N_5446);
nor U5605 (N_5605,N_5398,N_5344);
or U5606 (N_5606,N_5351,N_5279);
or U5607 (N_5607,N_5356,N_5491);
and U5608 (N_5608,N_5334,N_5359);
or U5609 (N_5609,N_5376,N_5461);
nor U5610 (N_5610,N_5280,N_5390);
xnor U5611 (N_5611,N_5352,N_5493);
nor U5612 (N_5612,N_5397,N_5368);
nor U5613 (N_5613,N_5321,N_5302);
nor U5614 (N_5614,N_5251,N_5372);
nor U5615 (N_5615,N_5292,N_5346);
nor U5616 (N_5616,N_5347,N_5337);
or U5617 (N_5617,N_5458,N_5490);
nor U5618 (N_5618,N_5295,N_5274);
xor U5619 (N_5619,N_5379,N_5338);
or U5620 (N_5620,N_5281,N_5339);
and U5621 (N_5621,N_5469,N_5332);
nand U5622 (N_5622,N_5435,N_5307);
nand U5623 (N_5623,N_5323,N_5445);
or U5624 (N_5624,N_5421,N_5312);
and U5625 (N_5625,N_5418,N_5331);
or U5626 (N_5626,N_5379,N_5386);
nor U5627 (N_5627,N_5467,N_5375);
or U5628 (N_5628,N_5359,N_5278);
or U5629 (N_5629,N_5413,N_5315);
or U5630 (N_5630,N_5398,N_5326);
or U5631 (N_5631,N_5358,N_5477);
nand U5632 (N_5632,N_5465,N_5495);
or U5633 (N_5633,N_5299,N_5374);
or U5634 (N_5634,N_5305,N_5372);
xnor U5635 (N_5635,N_5344,N_5397);
nor U5636 (N_5636,N_5491,N_5477);
and U5637 (N_5637,N_5396,N_5388);
nor U5638 (N_5638,N_5410,N_5250);
and U5639 (N_5639,N_5324,N_5393);
nor U5640 (N_5640,N_5343,N_5464);
nor U5641 (N_5641,N_5452,N_5456);
xnor U5642 (N_5642,N_5468,N_5378);
or U5643 (N_5643,N_5279,N_5367);
and U5644 (N_5644,N_5458,N_5347);
and U5645 (N_5645,N_5328,N_5449);
nand U5646 (N_5646,N_5302,N_5348);
or U5647 (N_5647,N_5467,N_5380);
nand U5648 (N_5648,N_5292,N_5469);
nor U5649 (N_5649,N_5326,N_5309);
xnor U5650 (N_5650,N_5259,N_5292);
nand U5651 (N_5651,N_5499,N_5358);
and U5652 (N_5652,N_5468,N_5393);
xor U5653 (N_5653,N_5485,N_5289);
nor U5654 (N_5654,N_5490,N_5485);
nor U5655 (N_5655,N_5486,N_5311);
or U5656 (N_5656,N_5414,N_5344);
xnor U5657 (N_5657,N_5271,N_5499);
nand U5658 (N_5658,N_5361,N_5486);
nand U5659 (N_5659,N_5419,N_5460);
nor U5660 (N_5660,N_5386,N_5253);
and U5661 (N_5661,N_5483,N_5443);
or U5662 (N_5662,N_5313,N_5339);
nand U5663 (N_5663,N_5345,N_5359);
nor U5664 (N_5664,N_5425,N_5390);
nand U5665 (N_5665,N_5336,N_5462);
or U5666 (N_5666,N_5447,N_5384);
and U5667 (N_5667,N_5388,N_5399);
nand U5668 (N_5668,N_5348,N_5374);
xor U5669 (N_5669,N_5365,N_5323);
xor U5670 (N_5670,N_5270,N_5406);
and U5671 (N_5671,N_5447,N_5425);
nor U5672 (N_5672,N_5422,N_5392);
and U5673 (N_5673,N_5322,N_5401);
nor U5674 (N_5674,N_5358,N_5322);
nor U5675 (N_5675,N_5435,N_5316);
nand U5676 (N_5676,N_5290,N_5365);
nand U5677 (N_5677,N_5283,N_5415);
nor U5678 (N_5678,N_5491,N_5346);
or U5679 (N_5679,N_5298,N_5396);
nand U5680 (N_5680,N_5321,N_5351);
nand U5681 (N_5681,N_5407,N_5480);
nand U5682 (N_5682,N_5460,N_5385);
nor U5683 (N_5683,N_5268,N_5421);
nor U5684 (N_5684,N_5459,N_5283);
nand U5685 (N_5685,N_5388,N_5336);
or U5686 (N_5686,N_5314,N_5379);
or U5687 (N_5687,N_5443,N_5463);
and U5688 (N_5688,N_5318,N_5254);
and U5689 (N_5689,N_5341,N_5489);
or U5690 (N_5690,N_5479,N_5364);
or U5691 (N_5691,N_5261,N_5321);
and U5692 (N_5692,N_5444,N_5264);
nor U5693 (N_5693,N_5252,N_5294);
or U5694 (N_5694,N_5294,N_5305);
or U5695 (N_5695,N_5384,N_5289);
or U5696 (N_5696,N_5277,N_5468);
nor U5697 (N_5697,N_5299,N_5366);
and U5698 (N_5698,N_5322,N_5385);
xor U5699 (N_5699,N_5364,N_5481);
nand U5700 (N_5700,N_5438,N_5386);
xnor U5701 (N_5701,N_5299,N_5499);
nor U5702 (N_5702,N_5251,N_5405);
or U5703 (N_5703,N_5294,N_5384);
nand U5704 (N_5704,N_5340,N_5328);
and U5705 (N_5705,N_5409,N_5374);
nor U5706 (N_5706,N_5392,N_5382);
nand U5707 (N_5707,N_5425,N_5256);
or U5708 (N_5708,N_5451,N_5453);
and U5709 (N_5709,N_5349,N_5328);
nand U5710 (N_5710,N_5481,N_5362);
nor U5711 (N_5711,N_5434,N_5307);
xnor U5712 (N_5712,N_5260,N_5271);
nand U5713 (N_5713,N_5458,N_5296);
or U5714 (N_5714,N_5419,N_5485);
or U5715 (N_5715,N_5375,N_5334);
nor U5716 (N_5716,N_5382,N_5367);
nand U5717 (N_5717,N_5377,N_5496);
nor U5718 (N_5718,N_5350,N_5311);
nand U5719 (N_5719,N_5272,N_5280);
xor U5720 (N_5720,N_5422,N_5489);
nor U5721 (N_5721,N_5455,N_5381);
nor U5722 (N_5722,N_5408,N_5285);
nor U5723 (N_5723,N_5359,N_5481);
nor U5724 (N_5724,N_5276,N_5393);
or U5725 (N_5725,N_5405,N_5479);
and U5726 (N_5726,N_5420,N_5276);
xnor U5727 (N_5727,N_5408,N_5394);
nand U5728 (N_5728,N_5259,N_5430);
nand U5729 (N_5729,N_5251,N_5375);
nor U5730 (N_5730,N_5364,N_5476);
nor U5731 (N_5731,N_5332,N_5344);
or U5732 (N_5732,N_5365,N_5317);
and U5733 (N_5733,N_5266,N_5316);
or U5734 (N_5734,N_5264,N_5318);
or U5735 (N_5735,N_5426,N_5449);
nand U5736 (N_5736,N_5386,N_5402);
or U5737 (N_5737,N_5417,N_5318);
and U5738 (N_5738,N_5308,N_5270);
nand U5739 (N_5739,N_5367,N_5354);
nor U5740 (N_5740,N_5314,N_5347);
xnor U5741 (N_5741,N_5365,N_5492);
nor U5742 (N_5742,N_5254,N_5404);
and U5743 (N_5743,N_5313,N_5408);
and U5744 (N_5744,N_5263,N_5392);
and U5745 (N_5745,N_5343,N_5257);
and U5746 (N_5746,N_5374,N_5279);
and U5747 (N_5747,N_5474,N_5273);
nor U5748 (N_5748,N_5475,N_5478);
nand U5749 (N_5749,N_5464,N_5266);
nor U5750 (N_5750,N_5545,N_5579);
nor U5751 (N_5751,N_5609,N_5543);
and U5752 (N_5752,N_5687,N_5550);
nand U5753 (N_5753,N_5696,N_5570);
nor U5754 (N_5754,N_5699,N_5680);
or U5755 (N_5755,N_5631,N_5530);
or U5756 (N_5756,N_5589,N_5618);
xnor U5757 (N_5757,N_5688,N_5627);
or U5758 (N_5758,N_5724,N_5639);
xor U5759 (N_5759,N_5528,N_5636);
or U5760 (N_5760,N_5526,N_5571);
nor U5761 (N_5761,N_5626,N_5660);
nand U5762 (N_5762,N_5506,N_5541);
xor U5763 (N_5763,N_5606,N_5709);
nand U5764 (N_5764,N_5652,N_5648);
or U5765 (N_5765,N_5519,N_5700);
nand U5766 (N_5766,N_5683,N_5516);
nor U5767 (N_5767,N_5518,N_5615);
and U5768 (N_5768,N_5720,N_5600);
nor U5769 (N_5769,N_5504,N_5632);
xor U5770 (N_5770,N_5686,N_5726);
and U5771 (N_5771,N_5583,N_5548);
and U5772 (N_5772,N_5634,N_5551);
or U5773 (N_5773,N_5509,N_5697);
or U5774 (N_5774,N_5559,N_5532);
or U5775 (N_5775,N_5647,N_5712);
and U5776 (N_5776,N_5710,N_5565);
or U5777 (N_5777,N_5538,N_5722);
and U5778 (N_5778,N_5597,N_5581);
or U5779 (N_5779,N_5733,N_5553);
or U5780 (N_5780,N_5662,N_5734);
and U5781 (N_5781,N_5555,N_5719);
nor U5782 (N_5782,N_5529,N_5507);
xnor U5783 (N_5783,N_5574,N_5547);
and U5784 (N_5784,N_5539,N_5706);
nand U5785 (N_5785,N_5681,N_5654);
nand U5786 (N_5786,N_5739,N_5513);
nor U5787 (N_5787,N_5588,N_5624);
or U5788 (N_5788,N_5748,N_5743);
and U5789 (N_5789,N_5694,N_5669);
and U5790 (N_5790,N_5691,N_5534);
nand U5791 (N_5791,N_5612,N_5501);
nand U5792 (N_5792,N_5586,N_5523);
nand U5793 (N_5793,N_5619,N_5564);
or U5794 (N_5794,N_5640,N_5704);
nor U5795 (N_5795,N_5718,N_5716);
or U5796 (N_5796,N_5708,N_5590);
and U5797 (N_5797,N_5741,N_5695);
and U5798 (N_5798,N_5749,N_5602);
and U5799 (N_5799,N_5663,N_5725);
or U5800 (N_5800,N_5653,N_5601);
nand U5801 (N_5801,N_5614,N_5670);
and U5802 (N_5802,N_5575,N_5587);
nor U5803 (N_5803,N_5536,N_5745);
or U5804 (N_5804,N_5641,N_5690);
nand U5805 (N_5805,N_5629,N_5702);
and U5806 (N_5806,N_5671,N_5540);
nor U5807 (N_5807,N_5525,N_5533);
nor U5808 (N_5808,N_5664,N_5630);
and U5809 (N_5809,N_5512,N_5567);
nand U5810 (N_5810,N_5578,N_5657);
or U5811 (N_5811,N_5582,N_5521);
or U5812 (N_5812,N_5591,N_5502);
and U5813 (N_5813,N_5542,N_5638);
or U5814 (N_5814,N_5572,N_5556);
nor U5815 (N_5815,N_5617,N_5595);
xnor U5816 (N_5816,N_5729,N_5684);
nor U5817 (N_5817,N_5593,N_5746);
nand U5818 (N_5818,N_5736,N_5577);
and U5819 (N_5819,N_5531,N_5679);
xor U5820 (N_5820,N_5744,N_5517);
or U5821 (N_5821,N_5611,N_5580);
nor U5822 (N_5822,N_5678,N_5658);
and U5823 (N_5823,N_5633,N_5735);
and U5824 (N_5824,N_5717,N_5723);
nor U5825 (N_5825,N_5625,N_5562);
and U5826 (N_5826,N_5705,N_5747);
nor U5827 (N_5827,N_5527,N_5650);
and U5828 (N_5828,N_5546,N_5620);
and U5829 (N_5829,N_5651,N_5558);
or U5830 (N_5830,N_5584,N_5605);
xor U5831 (N_5831,N_5596,N_5511);
or U5832 (N_5832,N_5676,N_5500);
and U5833 (N_5833,N_5552,N_5675);
nor U5834 (N_5834,N_5645,N_5635);
or U5835 (N_5835,N_5715,N_5714);
nor U5836 (N_5836,N_5674,N_5514);
or U5837 (N_5837,N_5549,N_5535);
nor U5838 (N_5838,N_5673,N_5659);
nor U5839 (N_5839,N_5701,N_5592);
or U5840 (N_5840,N_5731,N_5707);
and U5841 (N_5841,N_5505,N_5668);
or U5842 (N_5842,N_5522,N_5703);
nor U5843 (N_5843,N_5740,N_5585);
and U5844 (N_5844,N_5537,N_5561);
and U5845 (N_5845,N_5646,N_5616);
xor U5846 (N_5846,N_5693,N_5576);
nand U5847 (N_5847,N_5742,N_5728);
xor U5848 (N_5848,N_5613,N_5682);
and U5849 (N_5849,N_5510,N_5692);
nand U5850 (N_5850,N_5503,N_5594);
nand U5851 (N_5851,N_5544,N_5563);
and U5852 (N_5852,N_5608,N_5711);
and U5853 (N_5853,N_5643,N_5677);
or U5854 (N_5854,N_5738,N_5656);
or U5855 (N_5855,N_5721,N_5623);
and U5856 (N_5856,N_5573,N_5554);
and U5857 (N_5857,N_5732,N_5628);
and U5858 (N_5858,N_5621,N_5566);
or U5859 (N_5859,N_5644,N_5698);
and U5860 (N_5860,N_5637,N_5667);
xnor U5861 (N_5861,N_5730,N_5713);
nor U5862 (N_5862,N_5622,N_5560);
and U5863 (N_5863,N_5515,N_5665);
nor U5864 (N_5864,N_5568,N_5599);
nor U5865 (N_5865,N_5642,N_5569);
nor U5866 (N_5866,N_5557,N_5737);
nor U5867 (N_5867,N_5604,N_5661);
and U5868 (N_5868,N_5508,N_5685);
xor U5869 (N_5869,N_5598,N_5649);
nand U5870 (N_5870,N_5727,N_5666);
and U5871 (N_5871,N_5689,N_5520);
nor U5872 (N_5872,N_5672,N_5603);
or U5873 (N_5873,N_5524,N_5610);
or U5874 (N_5874,N_5607,N_5655);
or U5875 (N_5875,N_5714,N_5681);
and U5876 (N_5876,N_5599,N_5724);
and U5877 (N_5877,N_5671,N_5578);
nor U5878 (N_5878,N_5535,N_5552);
xor U5879 (N_5879,N_5533,N_5586);
or U5880 (N_5880,N_5568,N_5602);
or U5881 (N_5881,N_5725,N_5561);
xor U5882 (N_5882,N_5507,N_5552);
and U5883 (N_5883,N_5551,N_5638);
or U5884 (N_5884,N_5525,N_5596);
or U5885 (N_5885,N_5612,N_5623);
nand U5886 (N_5886,N_5607,N_5678);
nor U5887 (N_5887,N_5721,N_5625);
and U5888 (N_5888,N_5736,N_5573);
or U5889 (N_5889,N_5710,N_5576);
and U5890 (N_5890,N_5747,N_5732);
xnor U5891 (N_5891,N_5726,N_5502);
nor U5892 (N_5892,N_5504,N_5685);
nand U5893 (N_5893,N_5651,N_5517);
nand U5894 (N_5894,N_5651,N_5569);
nor U5895 (N_5895,N_5520,N_5748);
and U5896 (N_5896,N_5704,N_5645);
or U5897 (N_5897,N_5562,N_5633);
nor U5898 (N_5898,N_5672,N_5635);
and U5899 (N_5899,N_5533,N_5502);
xor U5900 (N_5900,N_5535,N_5619);
xnor U5901 (N_5901,N_5715,N_5591);
xor U5902 (N_5902,N_5543,N_5679);
or U5903 (N_5903,N_5666,N_5733);
and U5904 (N_5904,N_5521,N_5650);
or U5905 (N_5905,N_5567,N_5576);
and U5906 (N_5906,N_5520,N_5641);
and U5907 (N_5907,N_5620,N_5681);
or U5908 (N_5908,N_5558,N_5596);
nand U5909 (N_5909,N_5633,N_5563);
and U5910 (N_5910,N_5580,N_5541);
nor U5911 (N_5911,N_5734,N_5578);
nand U5912 (N_5912,N_5511,N_5609);
and U5913 (N_5913,N_5599,N_5709);
or U5914 (N_5914,N_5637,N_5540);
and U5915 (N_5915,N_5635,N_5684);
nor U5916 (N_5916,N_5603,N_5706);
nand U5917 (N_5917,N_5580,N_5683);
nor U5918 (N_5918,N_5712,N_5542);
nor U5919 (N_5919,N_5706,N_5740);
and U5920 (N_5920,N_5524,N_5528);
nor U5921 (N_5921,N_5512,N_5566);
or U5922 (N_5922,N_5613,N_5508);
nand U5923 (N_5923,N_5654,N_5700);
or U5924 (N_5924,N_5632,N_5720);
and U5925 (N_5925,N_5746,N_5634);
and U5926 (N_5926,N_5705,N_5669);
or U5927 (N_5927,N_5636,N_5534);
or U5928 (N_5928,N_5682,N_5635);
nor U5929 (N_5929,N_5675,N_5694);
and U5930 (N_5930,N_5536,N_5672);
or U5931 (N_5931,N_5596,N_5672);
or U5932 (N_5932,N_5534,N_5701);
nand U5933 (N_5933,N_5507,N_5524);
nand U5934 (N_5934,N_5732,N_5715);
or U5935 (N_5935,N_5667,N_5592);
and U5936 (N_5936,N_5583,N_5749);
nor U5937 (N_5937,N_5610,N_5690);
and U5938 (N_5938,N_5557,N_5551);
nor U5939 (N_5939,N_5517,N_5585);
nor U5940 (N_5940,N_5697,N_5711);
nor U5941 (N_5941,N_5565,N_5677);
xor U5942 (N_5942,N_5607,N_5533);
nand U5943 (N_5943,N_5667,N_5653);
or U5944 (N_5944,N_5541,N_5715);
or U5945 (N_5945,N_5536,N_5619);
and U5946 (N_5946,N_5743,N_5728);
and U5947 (N_5947,N_5702,N_5691);
or U5948 (N_5948,N_5516,N_5641);
nor U5949 (N_5949,N_5642,N_5664);
nor U5950 (N_5950,N_5623,N_5722);
and U5951 (N_5951,N_5636,N_5578);
nor U5952 (N_5952,N_5509,N_5546);
and U5953 (N_5953,N_5749,N_5658);
and U5954 (N_5954,N_5606,N_5718);
nand U5955 (N_5955,N_5585,N_5569);
nor U5956 (N_5956,N_5585,N_5686);
xnor U5957 (N_5957,N_5670,N_5618);
nor U5958 (N_5958,N_5586,N_5747);
or U5959 (N_5959,N_5573,N_5684);
xor U5960 (N_5960,N_5745,N_5686);
nand U5961 (N_5961,N_5584,N_5723);
nand U5962 (N_5962,N_5553,N_5547);
nand U5963 (N_5963,N_5728,N_5615);
nor U5964 (N_5964,N_5550,N_5652);
nor U5965 (N_5965,N_5713,N_5566);
nand U5966 (N_5966,N_5740,N_5618);
nand U5967 (N_5967,N_5520,N_5506);
nor U5968 (N_5968,N_5738,N_5735);
or U5969 (N_5969,N_5580,N_5722);
nor U5970 (N_5970,N_5508,N_5610);
or U5971 (N_5971,N_5580,N_5641);
and U5972 (N_5972,N_5505,N_5635);
nor U5973 (N_5973,N_5511,N_5718);
nand U5974 (N_5974,N_5506,N_5747);
or U5975 (N_5975,N_5573,N_5633);
or U5976 (N_5976,N_5573,N_5604);
nor U5977 (N_5977,N_5666,N_5651);
and U5978 (N_5978,N_5716,N_5507);
and U5979 (N_5979,N_5570,N_5564);
nand U5980 (N_5980,N_5612,N_5689);
or U5981 (N_5981,N_5719,N_5616);
nand U5982 (N_5982,N_5718,N_5507);
or U5983 (N_5983,N_5644,N_5581);
or U5984 (N_5984,N_5696,N_5731);
xnor U5985 (N_5985,N_5537,N_5623);
nor U5986 (N_5986,N_5625,N_5595);
nor U5987 (N_5987,N_5650,N_5670);
nor U5988 (N_5988,N_5747,N_5535);
and U5989 (N_5989,N_5726,N_5745);
xnor U5990 (N_5990,N_5730,N_5597);
nor U5991 (N_5991,N_5671,N_5678);
nor U5992 (N_5992,N_5570,N_5671);
nor U5993 (N_5993,N_5533,N_5567);
and U5994 (N_5994,N_5612,N_5603);
and U5995 (N_5995,N_5714,N_5710);
nand U5996 (N_5996,N_5533,N_5645);
nor U5997 (N_5997,N_5739,N_5516);
nand U5998 (N_5998,N_5596,N_5535);
xnor U5999 (N_5999,N_5680,N_5641);
nor U6000 (N_6000,N_5874,N_5913);
nor U6001 (N_6001,N_5832,N_5759);
and U6002 (N_6002,N_5948,N_5906);
or U6003 (N_6003,N_5815,N_5856);
and U6004 (N_6004,N_5890,N_5829);
and U6005 (N_6005,N_5784,N_5871);
or U6006 (N_6006,N_5845,N_5897);
or U6007 (N_6007,N_5786,N_5805);
and U6008 (N_6008,N_5953,N_5993);
xor U6009 (N_6009,N_5813,N_5797);
nand U6010 (N_6010,N_5831,N_5773);
nand U6011 (N_6011,N_5854,N_5892);
or U6012 (N_6012,N_5932,N_5981);
nand U6013 (N_6013,N_5764,N_5825);
and U6014 (N_6014,N_5954,N_5842);
or U6015 (N_6015,N_5859,N_5885);
nor U6016 (N_6016,N_5792,N_5976);
and U6017 (N_6017,N_5837,N_5939);
xor U6018 (N_6018,N_5836,N_5819);
xor U6019 (N_6019,N_5884,N_5956);
nand U6020 (N_6020,N_5811,N_5970);
and U6021 (N_6021,N_5794,N_5909);
or U6022 (N_6022,N_5750,N_5962);
nor U6023 (N_6023,N_5883,N_5992);
nor U6024 (N_6024,N_5843,N_5888);
nor U6025 (N_6025,N_5968,N_5991);
nand U6026 (N_6026,N_5933,N_5778);
and U6027 (N_6027,N_5938,N_5793);
xnor U6028 (N_6028,N_5789,N_5935);
and U6029 (N_6029,N_5766,N_5802);
nand U6030 (N_6030,N_5851,N_5965);
or U6031 (N_6031,N_5997,N_5882);
nand U6032 (N_6032,N_5881,N_5924);
nand U6033 (N_6033,N_5830,N_5969);
or U6034 (N_6034,N_5958,N_5860);
nor U6035 (N_6035,N_5966,N_5983);
nand U6036 (N_6036,N_5850,N_5790);
nand U6037 (N_6037,N_5855,N_5864);
nor U6038 (N_6038,N_5812,N_5910);
or U6039 (N_6039,N_5902,N_5770);
nor U6040 (N_6040,N_5899,N_5785);
xnor U6041 (N_6041,N_5868,N_5788);
nand U6042 (N_6042,N_5796,N_5753);
or U6043 (N_6043,N_5972,N_5936);
nor U6044 (N_6044,N_5781,N_5940);
or U6045 (N_6045,N_5853,N_5896);
or U6046 (N_6046,N_5922,N_5907);
or U6047 (N_6047,N_5877,N_5857);
and U6048 (N_6048,N_5893,N_5765);
or U6049 (N_6049,N_5973,N_5799);
nand U6050 (N_6050,N_5791,N_5921);
or U6051 (N_6051,N_5937,N_5756);
nand U6052 (N_6052,N_5801,N_5926);
nor U6053 (N_6053,N_5846,N_5995);
and U6054 (N_6054,N_5930,N_5951);
and U6055 (N_6055,N_5880,N_5964);
or U6056 (N_6056,N_5798,N_5984);
or U6057 (N_6057,N_5752,N_5823);
and U6058 (N_6058,N_5985,N_5818);
nor U6059 (N_6059,N_5863,N_5878);
nor U6060 (N_6060,N_5961,N_5783);
or U6061 (N_6061,N_5866,N_5996);
nor U6062 (N_6062,N_5959,N_5755);
nand U6063 (N_6063,N_5895,N_5879);
nand U6064 (N_6064,N_5894,N_5901);
and U6065 (N_6065,N_5840,N_5852);
xnor U6066 (N_6066,N_5967,N_5810);
or U6067 (N_6067,N_5987,N_5861);
nand U6068 (N_6068,N_5768,N_5862);
nor U6069 (N_6069,N_5787,N_5848);
nor U6070 (N_6070,N_5949,N_5898);
nand U6071 (N_6071,N_5931,N_5767);
nand U6072 (N_6072,N_5841,N_5941);
nand U6073 (N_6073,N_5919,N_5838);
nand U6074 (N_6074,N_5751,N_5988);
nand U6075 (N_6075,N_5809,N_5963);
nor U6076 (N_6076,N_5977,N_5771);
or U6077 (N_6077,N_5979,N_5975);
and U6078 (N_6078,N_5822,N_5908);
nor U6079 (N_6079,N_5986,N_5833);
nor U6080 (N_6080,N_5934,N_5777);
nand U6081 (N_6081,N_5955,N_5779);
nand U6082 (N_6082,N_5980,N_5903);
and U6083 (N_6083,N_5916,N_5914);
and U6084 (N_6084,N_5918,N_5917);
nor U6085 (N_6085,N_5816,N_5990);
nand U6086 (N_6086,N_5761,N_5891);
and U6087 (N_6087,N_5754,N_5904);
nor U6088 (N_6088,N_5849,N_5824);
and U6089 (N_6089,N_5873,N_5870);
and U6090 (N_6090,N_5839,N_5978);
or U6091 (N_6091,N_5814,N_5782);
nor U6092 (N_6092,N_5780,N_5875);
and U6093 (N_6093,N_5820,N_5945);
and U6094 (N_6094,N_5950,N_5947);
and U6095 (N_6095,N_5911,N_5808);
and U6096 (N_6096,N_5960,N_5905);
or U6097 (N_6097,N_5806,N_5974);
nor U6098 (N_6098,N_5869,N_5929);
or U6099 (N_6099,N_5925,N_5758);
nand U6100 (N_6100,N_5760,N_5847);
nand U6101 (N_6101,N_5774,N_5889);
and U6102 (N_6102,N_5776,N_5769);
nand U6103 (N_6103,N_5827,N_5920);
nand U6104 (N_6104,N_5867,N_5800);
nand U6105 (N_6105,N_5872,N_5757);
nand U6106 (N_6106,N_5982,N_5817);
and U6107 (N_6107,N_5858,N_5775);
nor U6108 (N_6108,N_5828,N_5928);
nand U6109 (N_6109,N_5989,N_5923);
or U6110 (N_6110,N_5772,N_5887);
or U6111 (N_6111,N_5942,N_5795);
and U6112 (N_6112,N_5971,N_5886);
nand U6113 (N_6113,N_5900,N_5912);
or U6114 (N_6114,N_5927,N_5803);
nor U6115 (N_6115,N_5844,N_5821);
and U6116 (N_6116,N_5943,N_5946);
and U6117 (N_6117,N_5826,N_5952);
or U6118 (N_6118,N_5994,N_5807);
nand U6119 (N_6119,N_5804,N_5944);
nor U6120 (N_6120,N_5957,N_5999);
nand U6121 (N_6121,N_5835,N_5834);
or U6122 (N_6122,N_5762,N_5763);
or U6123 (N_6123,N_5998,N_5876);
xnor U6124 (N_6124,N_5865,N_5915);
or U6125 (N_6125,N_5972,N_5929);
and U6126 (N_6126,N_5819,N_5788);
or U6127 (N_6127,N_5786,N_5980);
or U6128 (N_6128,N_5862,N_5940);
nand U6129 (N_6129,N_5973,N_5985);
nand U6130 (N_6130,N_5950,N_5920);
and U6131 (N_6131,N_5860,N_5939);
and U6132 (N_6132,N_5957,N_5985);
or U6133 (N_6133,N_5870,N_5840);
nand U6134 (N_6134,N_5939,N_5817);
and U6135 (N_6135,N_5999,N_5922);
or U6136 (N_6136,N_5849,N_5791);
nand U6137 (N_6137,N_5816,N_5963);
or U6138 (N_6138,N_5827,N_5876);
and U6139 (N_6139,N_5781,N_5796);
and U6140 (N_6140,N_5770,N_5810);
nand U6141 (N_6141,N_5761,N_5790);
nor U6142 (N_6142,N_5978,N_5932);
or U6143 (N_6143,N_5799,N_5994);
or U6144 (N_6144,N_5814,N_5942);
nand U6145 (N_6145,N_5851,N_5932);
or U6146 (N_6146,N_5927,N_5994);
nor U6147 (N_6147,N_5892,N_5903);
and U6148 (N_6148,N_5845,N_5941);
nor U6149 (N_6149,N_5879,N_5780);
nor U6150 (N_6150,N_5944,N_5978);
nor U6151 (N_6151,N_5940,N_5999);
and U6152 (N_6152,N_5906,N_5783);
and U6153 (N_6153,N_5848,N_5830);
nor U6154 (N_6154,N_5886,N_5852);
or U6155 (N_6155,N_5870,N_5805);
and U6156 (N_6156,N_5864,N_5852);
nand U6157 (N_6157,N_5910,N_5864);
nor U6158 (N_6158,N_5924,N_5905);
xnor U6159 (N_6159,N_5917,N_5772);
nor U6160 (N_6160,N_5788,N_5901);
nand U6161 (N_6161,N_5878,N_5956);
nor U6162 (N_6162,N_5934,N_5884);
nand U6163 (N_6163,N_5862,N_5847);
nand U6164 (N_6164,N_5980,N_5765);
and U6165 (N_6165,N_5836,N_5809);
xnor U6166 (N_6166,N_5804,N_5855);
nor U6167 (N_6167,N_5852,N_5761);
or U6168 (N_6168,N_5761,N_5859);
and U6169 (N_6169,N_5919,N_5912);
xnor U6170 (N_6170,N_5944,N_5989);
and U6171 (N_6171,N_5987,N_5767);
nand U6172 (N_6172,N_5968,N_5845);
nor U6173 (N_6173,N_5986,N_5911);
nor U6174 (N_6174,N_5951,N_5858);
or U6175 (N_6175,N_5759,N_5914);
nand U6176 (N_6176,N_5978,N_5976);
nand U6177 (N_6177,N_5933,N_5985);
and U6178 (N_6178,N_5838,N_5800);
nor U6179 (N_6179,N_5820,N_5943);
xor U6180 (N_6180,N_5843,N_5821);
nor U6181 (N_6181,N_5849,N_5872);
and U6182 (N_6182,N_5932,N_5760);
nor U6183 (N_6183,N_5842,N_5770);
and U6184 (N_6184,N_5920,N_5842);
nor U6185 (N_6185,N_5874,N_5778);
nor U6186 (N_6186,N_5886,N_5843);
or U6187 (N_6187,N_5925,N_5808);
and U6188 (N_6188,N_5822,N_5890);
and U6189 (N_6189,N_5768,N_5765);
and U6190 (N_6190,N_5790,N_5889);
nand U6191 (N_6191,N_5883,N_5977);
nor U6192 (N_6192,N_5822,N_5762);
or U6193 (N_6193,N_5879,N_5919);
or U6194 (N_6194,N_5775,N_5853);
nor U6195 (N_6195,N_5990,N_5928);
nor U6196 (N_6196,N_5955,N_5885);
nand U6197 (N_6197,N_5961,N_5946);
nand U6198 (N_6198,N_5972,N_5949);
or U6199 (N_6199,N_5960,N_5809);
nand U6200 (N_6200,N_5871,N_5981);
xnor U6201 (N_6201,N_5914,N_5795);
nor U6202 (N_6202,N_5757,N_5933);
nor U6203 (N_6203,N_5963,N_5924);
and U6204 (N_6204,N_5863,N_5964);
or U6205 (N_6205,N_5937,N_5966);
nor U6206 (N_6206,N_5881,N_5942);
nor U6207 (N_6207,N_5937,N_5926);
or U6208 (N_6208,N_5881,N_5776);
nor U6209 (N_6209,N_5942,N_5869);
or U6210 (N_6210,N_5813,N_5817);
nand U6211 (N_6211,N_5936,N_5990);
or U6212 (N_6212,N_5776,N_5972);
or U6213 (N_6213,N_5981,N_5794);
nor U6214 (N_6214,N_5836,N_5772);
nor U6215 (N_6215,N_5770,N_5903);
and U6216 (N_6216,N_5903,N_5936);
and U6217 (N_6217,N_5889,N_5893);
nor U6218 (N_6218,N_5842,N_5898);
nand U6219 (N_6219,N_5865,N_5987);
nand U6220 (N_6220,N_5922,N_5926);
nand U6221 (N_6221,N_5783,N_5925);
nand U6222 (N_6222,N_5799,N_5767);
and U6223 (N_6223,N_5984,N_5856);
nor U6224 (N_6224,N_5990,N_5981);
nand U6225 (N_6225,N_5785,N_5828);
or U6226 (N_6226,N_5869,N_5819);
nor U6227 (N_6227,N_5923,N_5766);
or U6228 (N_6228,N_5961,N_5774);
and U6229 (N_6229,N_5910,N_5935);
nor U6230 (N_6230,N_5772,N_5919);
nor U6231 (N_6231,N_5788,N_5896);
or U6232 (N_6232,N_5881,N_5926);
nand U6233 (N_6233,N_5955,N_5833);
and U6234 (N_6234,N_5984,N_5819);
nand U6235 (N_6235,N_5895,N_5923);
or U6236 (N_6236,N_5820,N_5853);
nand U6237 (N_6237,N_5904,N_5948);
xnor U6238 (N_6238,N_5890,N_5786);
nand U6239 (N_6239,N_5840,N_5882);
or U6240 (N_6240,N_5902,N_5823);
or U6241 (N_6241,N_5786,N_5944);
or U6242 (N_6242,N_5779,N_5891);
xnor U6243 (N_6243,N_5869,N_5844);
or U6244 (N_6244,N_5785,N_5879);
xnor U6245 (N_6245,N_5935,N_5927);
and U6246 (N_6246,N_5963,N_5755);
and U6247 (N_6247,N_5882,N_5754);
nor U6248 (N_6248,N_5926,N_5823);
or U6249 (N_6249,N_5932,N_5768);
nor U6250 (N_6250,N_6170,N_6150);
or U6251 (N_6251,N_6229,N_6165);
nand U6252 (N_6252,N_6242,N_6207);
or U6253 (N_6253,N_6070,N_6206);
nor U6254 (N_6254,N_6054,N_6064);
and U6255 (N_6255,N_6081,N_6208);
nand U6256 (N_6256,N_6084,N_6043);
nor U6257 (N_6257,N_6130,N_6205);
xor U6258 (N_6258,N_6066,N_6236);
nor U6259 (N_6259,N_6180,N_6055);
and U6260 (N_6260,N_6083,N_6216);
nand U6261 (N_6261,N_6020,N_6171);
or U6262 (N_6262,N_6169,N_6082);
or U6263 (N_6263,N_6154,N_6100);
nor U6264 (N_6264,N_6226,N_6010);
nand U6265 (N_6265,N_6155,N_6214);
nor U6266 (N_6266,N_6179,N_6118);
xnor U6267 (N_6267,N_6167,N_6005);
nor U6268 (N_6268,N_6058,N_6056);
or U6269 (N_6269,N_6107,N_6031);
or U6270 (N_6270,N_6124,N_6077);
and U6271 (N_6271,N_6157,N_6106);
nor U6272 (N_6272,N_6116,N_6046);
or U6273 (N_6273,N_6172,N_6194);
and U6274 (N_6274,N_6186,N_6249);
or U6275 (N_6275,N_6018,N_6240);
and U6276 (N_6276,N_6022,N_6193);
and U6277 (N_6277,N_6101,N_6023);
nor U6278 (N_6278,N_6080,N_6147);
and U6279 (N_6279,N_6132,N_6160);
nand U6280 (N_6280,N_6007,N_6033);
xor U6281 (N_6281,N_6145,N_6152);
nand U6282 (N_6282,N_6238,N_6036);
and U6283 (N_6283,N_6227,N_6091);
and U6284 (N_6284,N_6026,N_6168);
or U6285 (N_6285,N_6140,N_6177);
nand U6286 (N_6286,N_6039,N_6174);
xor U6287 (N_6287,N_6059,N_6137);
nand U6288 (N_6288,N_6089,N_6149);
and U6289 (N_6289,N_6196,N_6215);
or U6290 (N_6290,N_6004,N_6209);
xnor U6291 (N_6291,N_6025,N_6104);
or U6292 (N_6292,N_6146,N_6225);
nand U6293 (N_6293,N_6060,N_6203);
or U6294 (N_6294,N_6097,N_6049);
xnor U6295 (N_6295,N_6123,N_6078);
or U6296 (N_6296,N_6135,N_6173);
nand U6297 (N_6297,N_6204,N_6142);
or U6298 (N_6298,N_6245,N_6069);
or U6299 (N_6299,N_6028,N_6122);
nor U6300 (N_6300,N_6011,N_6000);
nor U6301 (N_6301,N_6079,N_6239);
nand U6302 (N_6302,N_6200,N_6029);
nand U6303 (N_6303,N_6187,N_6199);
and U6304 (N_6304,N_6190,N_6048);
or U6305 (N_6305,N_6153,N_6198);
xor U6306 (N_6306,N_6213,N_6073);
or U6307 (N_6307,N_6212,N_6136);
and U6308 (N_6308,N_6067,N_6144);
xor U6309 (N_6309,N_6158,N_6139);
or U6310 (N_6310,N_6098,N_6013);
nor U6311 (N_6311,N_6143,N_6201);
xnor U6312 (N_6312,N_6243,N_6181);
nand U6313 (N_6313,N_6197,N_6040);
and U6314 (N_6314,N_6138,N_6034);
or U6315 (N_6315,N_6113,N_6159);
nor U6316 (N_6316,N_6027,N_6095);
or U6317 (N_6317,N_6014,N_6217);
xnor U6318 (N_6318,N_6108,N_6006);
or U6319 (N_6319,N_6156,N_6244);
or U6320 (N_6320,N_6133,N_6176);
nand U6321 (N_6321,N_6182,N_6037);
nor U6322 (N_6322,N_6087,N_6072);
nor U6323 (N_6323,N_6131,N_6047);
or U6324 (N_6324,N_6052,N_6125);
and U6325 (N_6325,N_6185,N_6085);
or U6326 (N_6326,N_6162,N_6109);
nand U6327 (N_6327,N_6178,N_6112);
and U6328 (N_6328,N_6166,N_6231);
or U6329 (N_6329,N_6088,N_6202);
or U6330 (N_6330,N_6230,N_6045);
nor U6331 (N_6331,N_6105,N_6099);
or U6332 (N_6332,N_6161,N_6117);
and U6333 (N_6333,N_6235,N_6019);
or U6334 (N_6334,N_6042,N_6032);
and U6335 (N_6335,N_6062,N_6110);
and U6336 (N_6336,N_6188,N_6090);
nor U6337 (N_6337,N_6128,N_6017);
xnor U6338 (N_6338,N_6184,N_6102);
nand U6339 (N_6339,N_6057,N_6003);
nor U6340 (N_6340,N_6232,N_6223);
nor U6341 (N_6341,N_6041,N_6195);
nor U6342 (N_6342,N_6068,N_6044);
or U6343 (N_6343,N_6119,N_6224);
or U6344 (N_6344,N_6183,N_6129);
nor U6345 (N_6345,N_6115,N_6220);
or U6346 (N_6346,N_6141,N_6086);
or U6347 (N_6347,N_6071,N_6015);
nand U6348 (N_6348,N_6222,N_6246);
or U6349 (N_6349,N_6234,N_6211);
xor U6350 (N_6350,N_6189,N_6247);
nand U6351 (N_6351,N_6148,N_6038);
and U6352 (N_6352,N_6075,N_6035);
xor U6353 (N_6353,N_6093,N_6051);
nand U6354 (N_6354,N_6241,N_6103);
or U6355 (N_6355,N_6065,N_6218);
nand U6356 (N_6356,N_6175,N_6008);
or U6357 (N_6357,N_6050,N_6191);
or U6358 (N_6358,N_6016,N_6111);
nor U6359 (N_6359,N_6092,N_6021);
and U6360 (N_6360,N_6120,N_6076);
or U6361 (N_6361,N_6061,N_6074);
and U6362 (N_6362,N_6063,N_6163);
nand U6363 (N_6363,N_6053,N_6024);
nor U6364 (N_6364,N_6121,N_6210);
xnor U6365 (N_6365,N_6237,N_6192);
nor U6366 (N_6366,N_6009,N_6164);
or U6367 (N_6367,N_6114,N_6096);
nand U6368 (N_6368,N_6219,N_6094);
xnor U6369 (N_6369,N_6001,N_6248);
nand U6370 (N_6370,N_6221,N_6126);
nand U6371 (N_6371,N_6134,N_6127);
nand U6372 (N_6372,N_6012,N_6030);
nor U6373 (N_6373,N_6151,N_6002);
and U6374 (N_6374,N_6233,N_6228);
xnor U6375 (N_6375,N_6242,N_6239);
nand U6376 (N_6376,N_6104,N_6205);
nand U6377 (N_6377,N_6001,N_6029);
or U6378 (N_6378,N_6017,N_6137);
nand U6379 (N_6379,N_6137,N_6211);
nand U6380 (N_6380,N_6131,N_6097);
nand U6381 (N_6381,N_6170,N_6249);
nand U6382 (N_6382,N_6015,N_6248);
nor U6383 (N_6383,N_6164,N_6231);
or U6384 (N_6384,N_6093,N_6230);
and U6385 (N_6385,N_6077,N_6173);
and U6386 (N_6386,N_6129,N_6058);
and U6387 (N_6387,N_6170,N_6066);
or U6388 (N_6388,N_6084,N_6152);
nand U6389 (N_6389,N_6129,N_6003);
and U6390 (N_6390,N_6013,N_6169);
nor U6391 (N_6391,N_6203,N_6047);
and U6392 (N_6392,N_6104,N_6182);
or U6393 (N_6393,N_6005,N_6019);
nor U6394 (N_6394,N_6100,N_6041);
or U6395 (N_6395,N_6005,N_6194);
and U6396 (N_6396,N_6104,N_6136);
xnor U6397 (N_6397,N_6157,N_6025);
nand U6398 (N_6398,N_6041,N_6018);
or U6399 (N_6399,N_6009,N_6209);
or U6400 (N_6400,N_6044,N_6158);
or U6401 (N_6401,N_6133,N_6185);
or U6402 (N_6402,N_6055,N_6186);
or U6403 (N_6403,N_6118,N_6046);
xnor U6404 (N_6404,N_6169,N_6223);
nor U6405 (N_6405,N_6201,N_6160);
nand U6406 (N_6406,N_6047,N_6132);
nand U6407 (N_6407,N_6172,N_6189);
or U6408 (N_6408,N_6202,N_6118);
or U6409 (N_6409,N_6194,N_6102);
or U6410 (N_6410,N_6139,N_6227);
or U6411 (N_6411,N_6201,N_6172);
or U6412 (N_6412,N_6229,N_6021);
nor U6413 (N_6413,N_6166,N_6236);
nor U6414 (N_6414,N_6005,N_6190);
and U6415 (N_6415,N_6082,N_6022);
or U6416 (N_6416,N_6219,N_6093);
or U6417 (N_6417,N_6244,N_6041);
and U6418 (N_6418,N_6108,N_6174);
nand U6419 (N_6419,N_6015,N_6136);
and U6420 (N_6420,N_6029,N_6096);
and U6421 (N_6421,N_6181,N_6031);
nor U6422 (N_6422,N_6138,N_6230);
nor U6423 (N_6423,N_6086,N_6238);
nor U6424 (N_6424,N_6158,N_6197);
nand U6425 (N_6425,N_6183,N_6207);
nand U6426 (N_6426,N_6139,N_6054);
nand U6427 (N_6427,N_6207,N_6149);
and U6428 (N_6428,N_6160,N_6234);
nor U6429 (N_6429,N_6011,N_6062);
or U6430 (N_6430,N_6137,N_6098);
and U6431 (N_6431,N_6215,N_6130);
nor U6432 (N_6432,N_6079,N_6123);
nand U6433 (N_6433,N_6015,N_6201);
and U6434 (N_6434,N_6203,N_6131);
xor U6435 (N_6435,N_6036,N_6151);
or U6436 (N_6436,N_6042,N_6193);
nand U6437 (N_6437,N_6046,N_6146);
nor U6438 (N_6438,N_6064,N_6105);
or U6439 (N_6439,N_6038,N_6157);
nand U6440 (N_6440,N_6134,N_6090);
nand U6441 (N_6441,N_6234,N_6057);
nor U6442 (N_6442,N_6017,N_6088);
or U6443 (N_6443,N_6090,N_6192);
and U6444 (N_6444,N_6226,N_6126);
and U6445 (N_6445,N_6030,N_6170);
and U6446 (N_6446,N_6090,N_6011);
or U6447 (N_6447,N_6230,N_6132);
and U6448 (N_6448,N_6130,N_6185);
nor U6449 (N_6449,N_6038,N_6085);
nor U6450 (N_6450,N_6150,N_6101);
and U6451 (N_6451,N_6083,N_6221);
and U6452 (N_6452,N_6043,N_6172);
and U6453 (N_6453,N_6241,N_6197);
or U6454 (N_6454,N_6103,N_6179);
and U6455 (N_6455,N_6105,N_6167);
nand U6456 (N_6456,N_6207,N_6059);
or U6457 (N_6457,N_6190,N_6230);
xnor U6458 (N_6458,N_6210,N_6195);
or U6459 (N_6459,N_6021,N_6152);
nor U6460 (N_6460,N_6240,N_6141);
or U6461 (N_6461,N_6010,N_6180);
and U6462 (N_6462,N_6086,N_6101);
nand U6463 (N_6463,N_6062,N_6186);
or U6464 (N_6464,N_6030,N_6033);
and U6465 (N_6465,N_6147,N_6214);
and U6466 (N_6466,N_6095,N_6022);
nand U6467 (N_6467,N_6104,N_6084);
and U6468 (N_6468,N_6126,N_6087);
or U6469 (N_6469,N_6174,N_6215);
and U6470 (N_6470,N_6090,N_6142);
and U6471 (N_6471,N_6096,N_6147);
nor U6472 (N_6472,N_6202,N_6054);
and U6473 (N_6473,N_6148,N_6119);
nor U6474 (N_6474,N_6147,N_6024);
nor U6475 (N_6475,N_6032,N_6202);
and U6476 (N_6476,N_6223,N_6180);
nand U6477 (N_6477,N_6188,N_6185);
nor U6478 (N_6478,N_6181,N_6224);
nor U6479 (N_6479,N_6023,N_6246);
nand U6480 (N_6480,N_6160,N_6218);
or U6481 (N_6481,N_6027,N_6091);
nor U6482 (N_6482,N_6017,N_6049);
nand U6483 (N_6483,N_6131,N_6234);
xor U6484 (N_6484,N_6188,N_6144);
and U6485 (N_6485,N_6161,N_6114);
and U6486 (N_6486,N_6019,N_6056);
and U6487 (N_6487,N_6190,N_6000);
and U6488 (N_6488,N_6019,N_6144);
nand U6489 (N_6489,N_6198,N_6051);
xor U6490 (N_6490,N_6050,N_6005);
nor U6491 (N_6491,N_6231,N_6165);
and U6492 (N_6492,N_6239,N_6194);
nor U6493 (N_6493,N_6207,N_6063);
nand U6494 (N_6494,N_6238,N_6088);
or U6495 (N_6495,N_6016,N_6181);
and U6496 (N_6496,N_6108,N_6236);
xor U6497 (N_6497,N_6217,N_6037);
and U6498 (N_6498,N_6031,N_6218);
and U6499 (N_6499,N_6038,N_6245);
nand U6500 (N_6500,N_6389,N_6281);
nand U6501 (N_6501,N_6266,N_6378);
or U6502 (N_6502,N_6347,N_6338);
and U6503 (N_6503,N_6467,N_6363);
or U6504 (N_6504,N_6299,N_6447);
or U6505 (N_6505,N_6353,N_6448);
nand U6506 (N_6506,N_6316,N_6414);
nand U6507 (N_6507,N_6396,N_6436);
nor U6508 (N_6508,N_6428,N_6304);
and U6509 (N_6509,N_6290,N_6451);
and U6510 (N_6510,N_6477,N_6251);
nor U6511 (N_6511,N_6429,N_6466);
nor U6512 (N_6512,N_6276,N_6493);
nand U6513 (N_6513,N_6464,N_6397);
and U6514 (N_6514,N_6339,N_6291);
nand U6515 (N_6515,N_6384,N_6376);
nand U6516 (N_6516,N_6398,N_6342);
nand U6517 (N_6517,N_6293,N_6416);
nor U6518 (N_6518,N_6431,N_6337);
nand U6519 (N_6519,N_6418,N_6457);
nand U6520 (N_6520,N_6278,N_6300);
xor U6521 (N_6521,N_6285,N_6286);
and U6522 (N_6522,N_6483,N_6375);
and U6523 (N_6523,N_6322,N_6474);
nand U6524 (N_6524,N_6459,N_6253);
xor U6525 (N_6525,N_6379,N_6391);
or U6526 (N_6526,N_6308,N_6479);
and U6527 (N_6527,N_6445,N_6453);
xor U6528 (N_6528,N_6380,N_6471);
and U6529 (N_6529,N_6425,N_6364);
nor U6530 (N_6530,N_6463,N_6263);
nand U6531 (N_6531,N_6257,N_6478);
nor U6532 (N_6532,N_6410,N_6468);
and U6533 (N_6533,N_6438,N_6486);
or U6534 (N_6534,N_6327,N_6336);
nand U6535 (N_6535,N_6345,N_6250);
nand U6536 (N_6536,N_6313,N_6310);
or U6537 (N_6537,N_6390,N_6427);
or U6538 (N_6538,N_6444,N_6275);
nand U6539 (N_6539,N_6287,N_6309);
nor U6540 (N_6540,N_6489,N_6279);
or U6541 (N_6541,N_6295,N_6356);
nor U6542 (N_6542,N_6482,N_6476);
or U6543 (N_6543,N_6294,N_6374);
nor U6544 (N_6544,N_6443,N_6352);
nor U6545 (N_6545,N_6383,N_6446);
and U6546 (N_6546,N_6320,N_6402);
nor U6547 (N_6547,N_6417,N_6487);
and U6548 (N_6548,N_6317,N_6498);
nor U6549 (N_6549,N_6344,N_6490);
nor U6550 (N_6550,N_6454,N_6298);
nor U6551 (N_6551,N_6387,N_6452);
and U6552 (N_6552,N_6284,N_6289);
nor U6553 (N_6553,N_6472,N_6343);
nand U6554 (N_6554,N_6430,N_6456);
nand U6555 (N_6555,N_6368,N_6455);
and U6556 (N_6556,N_6485,N_6305);
or U6557 (N_6557,N_6423,N_6371);
nand U6558 (N_6558,N_6432,N_6357);
or U6559 (N_6559,N_6499,N_6328);
nor U6560 (N_6560,N_6302,N_6481);
xor U6561 (N_6561,N_6470,N_6497);
or U6562 (N_6562,N_6435,N_6326);
and U6563 (N_6563,N_6355,N_6319);
or U6564 (N_6564,N_6484,N_6400);
or U6565 (N_6565,N_6268,N_6492);
nor U6566 (N_6566,N_6488,N_6480);
nand U6567 (N_6567,N_6282,N_6329);
nand U6568 (N_6568,N_6462,N_6333);
nor U6569 (N_6569,N_6382,N_6312);
xnor U6570 (N_6570,N_6404,N_6261);
and U6571 (N_6571,N_6296,N_6341);
nor U6572 (N_6572,N_6349,N_6385);
nor U6573 (N_6573,N_6424,N_6366);
nor U6574 (N_6574,N_6254,N_6473);
nand U6575 (N_6575,N_6461,N_6450);
or U6576 (N_6576,N_6421,N_6439);
nor U6577 (N_6577,N_6274,N_6272);
and U6578 (N_6578,N_6370,N_6394);
or U6579 (N_6579,N_6465,N_6264);
xor U6580 (N_6580,N_6469,N_6408);
nor U6581 (N_6581,N_6406,N_6340);
nand U6582 (N_6582,N_6354,N_6323);
nor U6583 (N_6583,N_6360,N_6388);
nand U6584 (N_6584,N_6433,N_6365);
and U6585 (N_6585,N_6399,N_6386);
or U6586 (N_6586,N_6265,N_6409);
and U6587 (N_6587,N_6273,N_6334);
nor U6588 (N_6588,N_6392,N_6412);
nand U6589 (N_6589,N_6332,N_6362);
nor U6590 (N_6590,N_6351,N_6437);
nand U6591 (N_6591,N_6315,N_6395);
nor U6592 (N_6592,N_6411,N_6367);
nor U6593 (N_6593,N_6258,N_6441);
nor U6594 (N_6594,N_6311,N_6372);
nand U6595 (N_6595,N_6458,N_6495);
nand U6596 (N_6596,N_6301,N_6460);
and U6597 (N_6597,N_6449,N_6321);
nand U6598 (N_6598,N_6259,N_6252);
or U6599 (N_6599,N_6381,N_6434);
nand U6600 (N_6600,N_6361,N_6292);
nor U6601 (N_6601,N_6277,N_6420);
nand U6602 (N_6602,N_6325,N_6359);
nand U6603 (N_6603,N_6422,N_6283);
nand U6604 (N_6604,N_6335,N_6330);
or U6605 (N_6605,N_6297,N_6314);
nand U6606 (N_6606,N_6271,N_6324);
and U6607 (N_6607,N_6426,N_6288);
nand U6608 (N_6608,N_6331,N_6307);
or U6609 (N_6609,N_6496,N_6306);
or U6610 (N_6610,N_6413,N_6270);
nand U6611 (N_6611,N_6318,N_6267);
nor U6612 (N_6612,N_6256,N_6358);
nand U6613 (N_6613,N_6269,N_6303);
and U6614 (N_6614,N_6401,N_6442);
nand U6615 (N_6615,N_6494,N_6346);
nor U6616 (N_6616,N_6415,N_6440);
or U6617 (N_6617,N_6260,N_6475);
and U6618 (N_6618,N_6369,N_6280);
nand U6619 (N_6619,N_6373,N_6348);
xnor U6620 (N_6620,N_6262,N_6491);
nand U6621 (N_6621,N_6403,N_6377);
and U6622 (N_6622,N_6255,N_6405);
nor U6623 (N_6623,N_6350,N_6407);
and U6624 (N_6624,N_6419,N_6393);
and U6625 (N_6625,N_6276,N_6478);
nand U6626 (N_6626,N_6416,N_6440);
xor U6627 (N_6627,N_6371,N_6271);
xnor U6628 (N_6628,N_6425,N_6399);
xor U6629 (N_6629,N_6441,N_6444);
nor U6630 (N_6630,N_6457,N_6264);
nand U6631 (N_6631,N_6467,N_6354);
nor U6632 (N_6632,N_6295,N_6299);
or U6633 (N_6633,N_6372,N_6446);
xor U6634 (N_6634,N_6467,N_6476);
or U6635 (N_6635,N_6334,N_6371);
and U6636 (N_6636,N_6461,N_6466);
nor U6637 (N_6637,N_6481,N_6456);
nand U6638 (N_6638,N_6277,N_6292);
and U6639 (N_6639,N_6254,N_6339);
or U6640 (N_6640,N_6397,N_6385);
nand U6641 (N_6641,N_6397,N_6440);
and U6642 (N_6642,N_6307,N_6398);
xnor U6643 (N_6643,N_6376,N_6331);
and U6644 (N_6644,N_6437,N_6277);
or U6645 (N_6645,N_6340,N_6324);
and U6646 (N_6646,N_6476,N_6497);
nor U6647 (N_6647,N_6326,N_6316);
nand U6648 (N_6648,N_6378,N_6416);
and U6649 (N_6649,N_6411,N_6350);
nor U6650 (N_6650,N_6370,N_6269);
or U6651 (N_6651,N_6440,N_6403);
or U6652 (N_6652,N_6445,N_6293);
nor U6653 (N_6653,N_6433,N_6458);
and U6654 (N_6654,N_6299,N_6354);
and U6655 (N_6655,N_6490,N_6370);
and U6656 (N_6656,N_6349,N_6258);
nor U6657 (N_6657,N_6400,N_6260);
nand U6658 (N_6658,N_6421,N_6448);
and U6659 (N_6659,N_6302,N_6334);
or U6660 (N_6660,N_6487,N_6486);
and U6661 (N_6661,N_6494,N_6456);
nor U6662 (N_6662,N_6458,N_6320);
nand U6663 (N_6663,N_6271,N_6252);
nand U6664 (N_6664,N_6405,N_6366);
nor U6665 (N_6665,N_6433,N_6417);
and U6666 (N_6666,N_6366,N_6280);
nand U6667 (N_6667,N_6435,N_6493);
and U6668 (N_6668,N_6499,N_6428);
nor U6669 (N_6669,N_6279,N_6408);
and U6670 (N_6670,N_6391,N_6400);
or U6671 (N_6671,N_6384,N_6438);
nor U6672 (N_6672,N_6435,N_6496);
and U6673 (N_6673,N_6340,N_6292);
nor U6674 (N_6674,N_6304,N_6447);
nor U6675 (N_6675,N_6366,N_6413);
xor U6676 (N_6676,N_6289,N_6396);
and U6677 (N_6677,N_6272,N_6407);
xnor U6678 (N_6678,N_6362,N_6497);
nor U6679 (N_6679,N_6420,N_6290);
nand U6680 (N_6680,N_6411,N_6296);
nand U6681 (N_6681,N_6268,N_6309);
or U6682 (N_6682,N_6395,N_6417);
or U6683 (N_6683,N_6317,N_6475);
nor U6684 (N_6684,N_6441,N_6356);
or U6685 (N_6685,N_6348,N_6266);
nor U6686 (N_6686,N_6493,N_6497);
nor U6687 (N_6687,N_6264,N_6450);
xor U6688 (N_6688,N_6423,N_6333);
nand U6689 (N_6689,N_6351,N_6353);
or U6690 (N_6690,N_6405,N_6327);
nor U6691 (N_6691,N_6475,N_6306);
or U6692 (N_6692,N_6305,N_6306);
or U6693 (N_6693,N_6364,N_6277);
nor U6694 (N_6694,N_6454,N_6384);
or U6695 (N_6695,N_6280,N_6454);
nand U6696 (N_6696,N_6473,N_6284);
xor U6697 (N_6697,N_6263,N_6441);
and U6698 (N_6698,N_6327,N_6348);
nor U6699 (N_6699,N_6274,N_6306);
nor U6700 (N_6700,N_6290,N_6473);
nor U6701 (N_6701,N_6313,N_6448);
nor U6702 (N_6702,N_6414,N_6425);
nor U6703 (N_6703,N_6365,N_6311);
and U6704 (N_6704,N_6474,N_6424);
nor U6705 (N_6705,N_6420,N_6332);
nor U6706 (N_6706,N_6359,N_6391);
and U6707 (N_6707,N_6453,N_6308);
and U6708 (N_6708,N_6424,N_6440);
nand U6709 (N_6709,N_6297,N_6357);
nand U6710 (N_6710,N_6426,N_6375);
nor U6711 (N_6711,N_6379,N_6322);
xor U6712 (N_6712,N_6293,N_6263);
nand U6713 (N_6713,N_6430,N_6262);
nand U6714 (N_6714,N_6345,N_6468);
or U6715 (N_6715,N_6398,N_6252);
and U6716 (N_6716,N_6412,N_6416);
nor U6717 (N_6717,N_6296,N_6388);
nor U6718 (N_6718,N_6432,N_6358);
and U6719 (N_6719,N_6487,N_6400);
or U6720 (N_6720,N_6343,N_6401);
and U6721 (N_6721,N_6433,N_6288);
or U6722 (N_6722,N_6420,N_6463);
nand U6723 (N_6723,N_6305,N_6373);
nor U6724 (N_6724,N_6259,N_6271);
or U6725 (N_6725,N_6420,N_6498);
and U6726 (N_6726,N_6305,N_6328);
xnor U6727 (N_6727,N_6258,N_6428);
xor U6728 (N_6728,N_6456,N_6419);
or U6729 (N_6729,N_6282,N_6420);
and U6730 (N_6730,N_6389,N_6354);
xnor U6731 (N_6731,N_6416,N_6377);
xnor U6732 (N_6732,N_6448,N_6369);
and U6733 (N_6733,N_6351,N_6254);
and U6734 (N_6734,N_6360,N_6325);
and U6735 (N_6735,N_6381,N_6424);
nand U6736 (N_6736,N_6338,N_6384);
and U6737 (N_6737,N_6310,N_6345);
or U6738 (N_6738,N_6484,N_6410);
or U6739 (N_6739,N_6484,N_6397);
nand U6740 (N_6740,N_6311,N_6303);
nor U6741 (N_6741,N_6391,N_6422);
or U6742 (N_6742,N_6250,N_6429);
and U6743 (N_6743,N_6377,N_6286);
nand U6744 (N_6744,N_6457,N_6314);
nor U6745 (N_6745,N_6452,N_6451);
nand U6746 (N_6746,N_6418,N_6367);
or U6747 (N_6747,N_6391,N_6442);
nand U6748 (N_6748,N_6315,N_6342);
nand U6749 (N_6749,N_6285,N_6352);
or U6750 (N_6750,N_6672,N_6644);
and U6751 (N_6751,N_6581,N_6535);
nand U6752 (N_6752,N_6541,N_6542);
or U6753 (N_6753,N_6520,N_6736);
nand U6754 (N_6754,N_6621,N_6539);
nor U6755 (N_6755,N_6508,N_6507);
nor U6756 (N_6756,N_6579,N_6622);
nand U6757 (N_6757,N_6688,N_6724);
nor U6758 (N_6758,N_6668,N_6698);
and U6759 (N_6759,N_6589,N_6592);
and U6760 (N_6760,N_6675,N_6658);
nand U6761 (N_6761,N_6591,N_6551);
and U6762 (N_6762,N_6700,N_6739);
or U6763 (N_6763,N_6637,N_6561);
and U6764 (N_6764,N_6533,N_6543);
nand U6765 (N_6765,N_6529,N_6638);
nand U6766 (N_6766,N_6524,N_6619);
and U6767 (N_6767,N_6699,N_6580);
nor U6768 (N_6768,N_6671,N_6726);
and U6769 (N_6769,N_6646,N_6634);
and U6770 (N_6770,N_6596,N_6563);
and U6771 (N_6771,N_6704,N_6722);
xor U6772 (N_6772,N_6576,N_6661);
nand U6773 (N_6773,N_6626,N_6728);
and U6774 (N_6774,N_6662,N_6749);
xor U6775 (N_6775,N_6657,N_6606);
nand U6776 (N_6776,N_6603,N_6540);
nand U6777 (N_6777,N_6557,N_6531);
or U6778 (N_6778,N_6614,N_6690);
or U6779 (N_6779,N_6652,N_6546);
and U6780 (N_6780,N_6665,N_6547);
or U6781 (N_6781,N_6718,N_6641);
and U6782 (N_6782,N_6509,N_6569);
nor U6783 (N_6783,N_6677,N_6744);
xor U6784 (N_6784,N_6611,N_6574);
and U6785 (N_6785,N_6567,N_6600);
xnor U6786 (N_6786,N_6708,N_6727);
nor U6787 (N_6787,N_6512,N_6729);
or U6788 (N_6788,N_6740,N_6588);
nand U6789 (N_6789,N_6682,N_6716);
and U6790 (N_6790,N_6676,N_6679);
nand U6791 (N_6791,N_6544,N_6640);
and U6792 (N_6792,N_6526,N_6738);
and U6793 (N_6793,N_6659,N_6721);
nand U6794 (N_6794,N_6678,N_6697);
or U6795 (N_6795,N_6733,N_6734);
and U6796 (N_6796,N_6552,N_6564);
xor U6797 (N_6797,N_6627,N_6607);
nor U6798 (N_6798,N_6536,N_6655);
or U6799 (N_6799,N_6735,N_6712);
or U6800 (N_6800,N_6654,N_6573);
and U6801 (N_6801,N_6534,N_6667);
nor U6802 (N_6802,N_6685,N_6616);
nor U6803 (N_6803,N_6532,N_6683);
or U6804 (N_6804,N_6741,N_6503);
nor U6805 (N_6805,N_6710,N_6742);
nand U6806 (N_6806,N_6550,N_6702);
nor U6807 (N_6807,N_6624,N_6516);
and U6808 (N_6808,N_6554,N_6720);
or U6809 (N_6809,N_6649,N_6639);
and U6810 (N_6810,N_6594,N_6748);
nor U6811 (N_6811,N_6731,N_6703);
and U6812 (N_6812,N_6701,N_6537);
or U6813 (N_6813,N_6525,N_6610);
nand U6814 (N_6814,N_6743,N_6605);
nand U6815 (N_6815,N_6681,N_6625);
or U6816 (N_6816,N_6745,N_6713);
and U6817 (N_6817,N_6632,N_6715);
nor U6818 (N_6818,N_6617,N_6686);
nor U6819 (N_6819,N_6695,N_6631);
nand U6820 (N_6820,N_6527,N_6669);
nor U6821 (N_6821,N_6714,N_6555);
nand U6822 (N_6822,N_6664,N_6586);
and U6823 (N_6823,N_6500,N_6696);
xnor U6824 (N_6824,N_6663,N_6612);
or U6825 (N_6825,N_6666,N_6636);
nand U6826 (N_6826,N_6523,N_6577);
or U6827 (N_6827,N_6511,N_6583);
nor U6828 (N_6828,N_6684,N_6566);
nor U6829 (N_6829,N_6746,N_6515);
and U6830 (N_6830,N_6689,N_6693);
nor U6831 (N_6831,N_6687,N_6732);
nor U6832 (N_6832,N_6623,N_6629);
nand U6833 (N_6833,N_6502,N_6670);
nor U6834 (N_6834,N_6575,N_6584);
nand U6835 (N_6835,N_6694,N_6602);
nand U6836 (N_6836,N_6618,N_6571);
nor U6837 (N_6837,N_6530,N_6707);
and U6838 (N_6838,N_6706,N_6660);
and U6839 (N_6839,N_6674,N_6599);
nor U6840 (N_6840,N_6598,N_6538);
or U6841 (N_6841,N_6730,N_6514);
nor U6842 (N_6842,N_6609,N_6518);
nor U6843 (N_6843,N_6521,N_6717);
or U6844 (N_6844,N_6528,N_6590);
or U6845 (N_6845,N_6651,N_6513);
nor U6846 (N_6846,N_6711,N_6556);
nor U6847 (N_6847,N_6608,N_6656);
and U6848 (N_6848,N_6680,N_6747);
and U6849 (N_6849,N_6553,N_6595);
or U6850 (N_6850,N_6620,N_6559);
nand U6851 (N_6851,N_6692,N_6635);
nand U6852 (N_6852,N_6506,N_6504);
or U6853 (N_6853,N_6737,N_6725);
nand U6854 (N_6854,N_6723,N_6615);
nor U6855 (N_6855,N_6549,N_6572);
or U6856 (N_6856,N_6601,N_6593);
nand U6857 (N_6857,N_6645,N_6501);
or U6858 (N_6858,N_6709,N_6522);
nor U6859 (N_6859,N_6650,N_6673);
and U6860 (N_6860,N_6633,N_6691);
and U6861 (N_6861,N_6505,N_6587);
or U6862 (N_6862,N_6582,N_6604);
nand U6863 (N_6863,N_6578,N_6705);
and U6864 (N_6864,N_6519,N_6643);
and U6865 (N_6865,N_6653,N_6510);
and U6866 (N_6866,N_6642,N_6585);
or U6867 (N_6867,N_6548,N_6719);
and U6868 (N_6868,N_6613,N_6630);
or U6869 (N_6869,N_6560,N_6545);
xnor U6870 (N_6870,N_6558,N_6648);
and U6871 (N_6871,N_6570,N_6568);
and U6872 (N_6872,N_6517,N_6597);
or U6873 (N_6873,N_6628,N_6562);
and U6874 (N_6874,N_6565,N_6647);
nand U6875 (N_6875,N_6696,N_6580);
or U6876 (N_6876,N_6537,N_6529);
and U6877 (N_6877,N_6603,N_6549);
and U6878 (N_6878,N_6567,N_6546);
nand U6879 (N_6879,N_6589,N_6596);
nor U6880 (N_6880,N_6615,N_6613);
xor U6881 (N_6881,N_6620,N_6626);
xnor U6882 (N_6882,N_6626,N_6553);
and U6883 (N_6883,N_6611,N_6650);
or U6884 (N_6884,N_6664,N_6680);
and U6885 (N_6885,N_6581,N_6716);
nand U6886 (N_6886,N_6571,N_6744);
or U6887 (N_6887,N_6646,N_6676);
xor U6888 (N_6888,N_6621,N_6695);
nand U6889 (N_6889,N_6680,N_6612);
or U6890 (N_6890,N_6654,N_6558);
nand U6891 (N_6891,N_6601,N_6645);
nand U6892 (N_6892,N_6749,N_6657);
or U6893 (N_6893,N_6705,N_6534);
or U6894 (N_6894,N_6692,N_6654);
xor U6895 (N_6895,N_6710,N_6638);
or U6896 (N_6896,N_6729,N_6748);
and U6897 (N_6897,N_6529,N_6561);
xnor U6898 (N_6898,N_6509,N_6602);
or U6899 (N_6899,N_6742,N_6616);
or U6900 (N_6900,N_6664,N_6693);
and U6901 (N_6901,N_6531,N_6653);
nor U6902 (N_6902,N_6559,N_6502);
and U6903 (N_6903,N_6580,N_6575);
nand U6904 (N_6904,N_6500,N_6656);
nand U6905 (N_6905,N_6501,N_6629);
or U6906 (N_6906,N_6532,N_6555);
nor U6907 (N_6907,N_6512,N_6588);
or U6908 (N_6908,N_6599,N_6513);
nor U6909 (N_6909,N_6532,N_6678);
nor U6910 (N_6910,N_6521,N_6591);
nor U6911 (N_6911,N_6643,N_6646);
and U6912 (N_6912,N_6738,N_6706);
nand U6913 (N_6913,N_6517,N_6669);
nand U6914 (N_6914,N_6598,N_6607);
and U6915 (N_6915,N_6554,N_6517);
nand U6916 (N_6916,N_6683,N_6717);
and U6917 (N_6917,N_6589,N_6558);
nand U6918 (N_6918,N_6679,N_6655);
and U6919 (N_6919,N_6590,N_6554);
nor U6920 (N_6920,N_6565,N_6526);
xnor U6921 (N_6921,N_6656,N_6623);
and U6922 (N_6922,N_6628,N_6690);
and U6923 (N_6923,N_6749,N_6534);
nor U6924 (N_6924,N_6539,N_6506);
and U6925 (N_6925,N_6639,N_6577);
nor U6926 (N_6926,N_6592,N_6707);
or U6927 (N_6927,N_6710,N_6561);
nand U6928 (N_6928,N_6718,N_6539);
or U6929 (N_6929,N_6601,N_6643);
nand U6930 (N_6930,N_6704,N_6604);
or U6931 (N_6931,N_6662,N_6626);
nand U6932 (N_6932,N_6718,N_6609);
or U6933 (N_6933,N_6589,N_6542);
or U6934 (N_6934,N_6739,N_6540);
nand U6935 (N_6935,N_6599,N_6711);
or U6936 (N_6936,N_6732,N_6648);
nor U6937 (N_6937,N_6658,N_6670);
and U6938 (N_6938,N_6520,N_6711);
nand U6939 (N_6939,N_6582,N_6673);
and U6940 (N_6940,N_6680,N_6595);
nand U6941 (N_6941,N_6611,N_6506);
or U6942 (N_6942,N_6669,N_6602);
and U6943 (N_6943,N_6628,N_6595);
nor U6944 (N_6944,N_6562,N_6659);
nor U6945 (N_6945,N_6619,N_6696);
and U6946 (N_6946,N_6677,N_6719);
and U6947 (N_6947,N_6631,N_6641);
nor U6948 (N_6948,N_6541,N_6679);
nand U6949 (N_6949,N_6517,N_6729);
nor U6950 (N_6950,N_6673,N_6656);
and U6951 (N_6951,N_6568,N_6502);
or U6952 (N_6952,N_6702,N_6703);
or U6953 (N_6953,N_6718,N_6527);
xnor U6954 (N_6954,N_6731,N_6609);
or U6955 (N_6955,N_6565,N_6531);
nand U6956 (N_6956,N_6596,N_6597);
nor U6957 (N_6957,N_6576,N_6685);
and U6958 (N_6958,N_6688,N_6609);
or U6959 (N_6959,N_6638,N_6644);
and U6960 (N_6960,N_6670,N_6542);
nand U6961 (N_6961,N_6589,N_6556);
nor U6962 (N_6962,N_6635,N_6701);
and U6963 (N_6963,N_6552,N_6588);
xnor U6964 (N_6964,N_6528,N_6668);
nor U6965 (N_6965,N_6614,N_6699);
nand U6966 (N_6966,N_6512,N_6566);
and U6967 (N_6967,N_6552,N_6629);
nor U6968 (N_6968,N_6746,N_6675);
nor U6969 (N_6969,N_6569,N_6562);
or U6970 (N_6970,N_6704,N_6747);
nand U6971 (N_6971,N_6706,N_6740);
nor U6972 (N_6972,N_6640,N_6666);
nand U6973 (N_6973,N_6737,N_6541);
nand U6974 (N_6974,N_6505,N_6719);
or U6975 (N_6975,N_6644,N_6622);
nand U6976 (N_6976,N_6638,N_6715);
nand U6977 (N_6977,N_6582,N_6556);
xor U6978 (N_6978,N_6608,N_6567);
nand U6979 (N_6979,N_6677,N_6742);
nor U6980 (N_6980,N_6723,N_6611);
nand U6981 (N_6981,N_6608,N_6638);
nor U6982 (N_6982,N_6705,N_6653);
or U6983 (N_6983,N_6623,N_6633);
or U6984 (N_6984,N_6536,N_6706);
nand U6985 (N_6985,N_6575,N_6654);
nor U6986 (N_6986,N_6615,N_6638);
xor U6987 (N_6987,N_6588,N_6548);
and U6988 (N_6988,N_6570,N_6749);
xor U6989 (N_6989,N_6669,N_6715);
nor U6990 (N_6990,N_6555,N_6596);
or U6991 (N_6991,N_6721,N_6703);
or U6992 (N_6992,N_6740,N_6663);
and U6993 (N_6993,N_6661,N_6744);
nor U6994 (N_6994,N_6652,N_6585);
nor U6995 (N_6995,N_6717,N_6701);
or U6996 (N_6996,N_6512,N_6524);
nand U6997 (N_6997,N_6580,N_6569);
and U6998 (N_6998,N_6712,N_6505);
nor U6999 (N_6999,N_6519,N_6711);
and U7000 (N_7000,N_6759,N_6973);
and U7001 (N_7001,N_6876,N_6839);
and U7002 (N_7002,N_6821,N_6782);
and U7003 (N_7003,N_6988,N_6844);
xnor U7004 (N_7004,N_6853,N_6858);
and U7005 (N_7005,N_6984,N_6945);
xnor U7006 (N_7006,N_6770,N_6921);
and U7007 (N_7007,N_6942,N_6867);
xnor U7008 (N_7008,N_6775,N_6927);
nand U7009 (N_7009,N_6972,N_6818);
or U7010 (N_7010,N_6791,N_6767);
xor U7011 (N_7011,N_6847,N_6930);
xor U7012 (N_7012,N_6790,N_6856);
nor U7013 (N_7013,N_6769,N_6850);
or U7014 (N_7014,N_6914,N_6889);
and U7015 (N_7015,N_6750,N_6865);
and U7016 (N_7016,N_6830,N_6892);
and U7017 (N_7017,N_6875,N_6819);
or U7018 (N_7018,N_6840,N_6776);
or U7019 (N_7019,N_6869,N_6887);
or U7020 (N_7020,N_6779,N_6969);
xor U7021 (N_7021,N_6934,N_6998);
nor U7022 (N_7022,N_6783,N_6754);
xnor U7023 (N_7023,N_6809,N_6826);
nand U7024 (N_7024,N_6918,N_6986);
or U7025 (N_7025,N_6857,N_6981);
nand U7026 (N_7026,N_6859,N_6813);
xor U7027 (N_7027,N_6837,N_6824);
nor U7028 (N_7028,N_6982,N_6841);
and U7029 (N_7029,N_6868,N_6863);
and U7030 (N_7030,N_6956,N_6796);
nand U7031 (N_7031,N_6985,N_6810);
or U7032 (N_7032,N_6937,N_6975);
nor U7033 (N_7033,N_6756,N_6989);
nor U7034 (N_7034,N_6885,N_6992);
or U7035 (N_7035,N_6772,N_6835);
nand U7036 (N_7036,N_6913,N_6827);
or U7037 (N_7037,N_6999,N_6955);
or U7038 (N_7038,N_6890,N_6933);
and U7039 (N_7039,N_6952,N_6752);
or U7040 (N_7040,N_6792,N_6820);
nand U7041 (N_7041,N_6947,N_6838);
or U7042 (N_7042,N_6939,N_6798);
or U7043 (N_7043,N_6753,N_6911);
nor U7044 (N_7044,N_6823,N_6870);
or U7045 (N_7045,N_6996,N_6771);
or U7046 (N_7046,N_6967,N_6803);
nor U7047 (N_7047,N_6825,N_6938);
and U7048 (N_7048,N_6904,N_6966);
or U7049 (N_7049,N_6874,N_6815);
nand U7050 (N_7050,N_6860,N_6788);
nor U7051 (N_7051,N_6961,N_6912);
and U7052 (N_7052,N_6768,N_6916);
nor U7053 (N_7053,N_6968,N_6855);
nand U7054 (N_7054,N_6964,N_6854);
nor U7055 (N_7055,N_6900,N_6959);
or U7056 (N_7056,N_6757,N_6828);
nand U7057 (N_7057,N_6931,N_6953);
and U7058 (N_7058,N_6977,N_6751);
nor U7059 (N_7059,N_6777,N_6995);
nand U7060 (N_7060,N_6929,N_6878);
and U7061 (N_7061,N_6990,N_6943);
xor U7062 (N_7062,N_6979,N_6843);
xor U7063 (N_7063,N_6994,N_6795);
nand U7064 (N_7064,N_6877,N_6910);
nor U7065 (N_7065,N_6925,N_6766);
nand U7066 (N_7066,N_6905,N_6897);
or U7067 (N_7067,N_6954,N_6948);
and U7068 (N_7068,N_6906,N_6893);
nand U7069 (N_7069,N_6836,N_6957);
or U7070 (N_7070,N_6755,N_6882);
nor U7071 (N_7071,N_6781,N_6902);
nand U7072 (N_7072,N_6950,N_6935);
xor U7073 (N_7073,N_6780,N_6864);
and U7074 (N_7074,N_6845,N_6812);
nor U7075 (N_7075,N_6808,N_6800);
or U7076 (N_7076,N_6763,N_6817);
nand U7077 (N_7077,N_6849,N_6926);
and U7078 (N_7078,N_6949,N_6794);
and U7079 (N_7079,N_6806,N_6822);
nor U7080 (N_7080,N_6928,N_6899);
nand U7081 (N_7081,N_6903,N_6846);
nand U7082 (N_7082,N_6799,N_6778);
nor U7083 (N_7083,N_6980,N_6872);
nor U7084 (N_7084,N_6787,N_6842);
and U7085 (N_7085,N_6797,N_6915);
nand U7086 (N_7086,N_6758,N_6886);
nor U7087 (N_7087,N_6962,N_6978);
nand U7088 (N_7088,N_6786,N_6879);
and U7089 (N_7089,N_6805,N_6881);
xor U7090 (N_7090,N_6833,N_6991);
nand U7091 (N_7091,N_6866,N_6765);
and U7092 (N_7092,N_6764,N_6873);
nor U7093 (N_7093,N_6936,N_6832);
and U7094 (N_7094,N_6785,N_6804);
nor U7095 (N_7095,N_6920,N_6909);
nor U7096 (N_7096,N_6784,N_6871);
nor U7097 (N_7097,N_6919,N_6940);
xor U7098 (N_7098,N_6829,N_6970);
and U7099 (N_7099,N_6831,N_6880);
and U7100 (N_7100,N_6971,N_6908);
or U7101 (N_7101,N_6773,N_6997);
nor U7102 (N_7102,N_6802,N_6983);
or U7103 (N_7103,N_6974,N_6901);
nor U7104 (N_7104,N_6894,N_6896);
nor U7105 (N_7105,N_6944,N_6774);
or U7106 (N_7106,N_6898,N_6958);
nand U7107 (N_7107,N_6917,N_6891);
or U7108 (N_7108,N_6965,N_6976);
nor U7109 (N_7109,N_6834,N_6862);
and U7110 (N_7110,N_6814,N_6762);
nand U7111 (N_7111,N_6941,N_6816);
and U7112 (N_7112,N_6922,N_6895);
and U7113 (N_7113,N_6960,N_6761);
or U7114 (N_7114,N_6848,N_6924);
and U7115 (N_7115,N_6907,N_6852);
nor U7116 (N_7116,N_6888,N_6789);
nand U7117 (N_7117,N_6861,N_6884);
nand U7118 (N_7118,N_6807,N_6811);
or U7119 (N_7119,N_6987,N_6851);
and U7120 (N_7120,N_6801,N_6946);
or U7121 (N_7121,N_6760,N_6993);
nor U7122 (N_7122,N_6793,N_6963);
and U7123 (N_7123,N_6932,N_6951);
nor U7124 (N_7124,N_6923,N_6883);
nor U7125 (N_7125,N_6773,N_6899);
nor U7126 (N_7126,N_6792,N_6817);
and U7127 (N_7127,N_6770,N_6974);
nor U7128 (N_7128,N_6981,N_6901);
and U7129 (N_7129,N_6889,N_6993);
or U7130 (N_7130,N_6881,N_6761);
nand U7131 (N_7131,N_6922,N_6850);
and U7132 (N_7132,N_6879,N_6852);
or U7133 (N_7133,N_6991,N_6802);
or U7134 (N_7134,N_6781,N_6773);
or U7135 (N_7135,N_6776,N_6870);
nor U7136 (N_7136,N_6943,N_6958);
or U7137 (N_7137,N_6944,N_6865);
nand U7138 (N_7138,N_6971,N_6790);
nor U7139 (N_7139,N_6853,N_6899);
xnor U7140 (N_7140,N_6842,N_6917);
and U7141 (N_7141,N_6949,N_6913);
or U7142 (N_7142,N_6903,N_6793);
nand U7143 (N_7143,N_6788,N_6974);
xnor U7144 (N_7144,N_6821,N_6778);
nand U7145 (N_7145,N_6753,N_6774);
nor U7146 (N_7146,N_6951,N_6770);
or U7147 (N_7147,N_6948,N_6820);
nor U7148 (N_7148,N_6806,N_6883);
or U7149 (N_7149,N_6967,N_6788);
xor U7150 (N_7150,N_6875,N_6973);
nand U7151 (N_7151,N_6926,N_6897);
nand U7152 (N_7152,N_6770,N_6820);
and U7153 (N_7153,N_6978,N_6793);
nor U7154 (N_7154,N_6987,N_6926);
and U7155 (N_7155,N_6916,N_6781);
nor U7156 (N_7156,N_6907,N_6789);
or U7157 (N_7157,N_6827,N_6889);
and U7158 (N_7158,N_6948,N_6780);
nand U7159 (N_7159,N_6774,N_6958);
nand U7160 (N_7160,N_6762,N_6992);
xor U7161 (N_7161,N_6857,N_6962);
nor U7162 (N_7162,N_6987,N_6783);
nor U7163 (N_7163,N_6757,N_6829);
and U7164 (N_7164,N_6798,N_6879);
nor U7165 (N_7165,N_6876,N_6866);
xnor U7166 (N_7166,N_6835,N_6839);
and U7167 (N_7167,N_6771,N_6848);
nand U7168 (N_7168,N_6752,N_6972);
or U7169 (N_7169,N_6839,N_6943);
and U7170 (N_7170,N_6980,N_6894);
nand U7171 (N_7171,N_6829,N_6858);
or U7172 (N_7172,N_6923,N_6823);
nor U7173 (N_7173,N_6918,N_6985);
or U7174 (N_7174,N_6770,N_6878);
or U7175 (N_7175,N_6755,N_6963);
nor U7176 (N_7176,N_6761,N_6906);
nor U7177 (N_7177,N_6811,N_6839);
or U7178 (N_7178,N_6858,N_6776);
nand U7179 (N_7179,N_6785,N_6921);
nor U7180 (N_7180,N_6882,N_6981);
nand U7181 (N_7181,N_6850,N_6876);
and U7182 (N_7182,N_6916,N_6934);
or U7183 (N_7183,N_6924,N_6820);
or U7184 (N_7184,N_6782,N_6987);
xor U7185 (N_7185,N_6946,N_6953);
and U7186 (N_7186,N_6757,N_6755);
or U7187 (N_7187,N_6787,N_6853);
xnor U7188 (N_7188,N_6766,N_6887);
or U7189 (N_7189,N_6800,N_6870);
nand U7190 (N_7190,N_6862,N_6884);
nor U7191 (N_7191,N_6816,N_6878);
nand U7192 (N_7192,N_6830,N_6867);
nand U7193 (N_7193,N_6880,N_6901);
and U7194 (N_7194,N_6795,N_6875);
and U7195 (N_7195,N_6783,N_6763);
nand U7196 (N_7196,N_6815,N_6860);
xor U7197 (N_7197,N_6981,N_6928);
nand U7198 (N_7198,N_6954,N_6852);
or U7199 (N_7199,N_6873,N_6826);
nand U7200 (N_7200,N_6944,N_6858);
nand U7201 (N_7201,N_6796,N_6761);
and U7202 (N_7202,N_6798,N_6961);
nor U7203 (N_7203,N_6918,N_6882);
and U7204 (N_7204,N_6836,N_6896);
nor U7205 (N_7205,N_6820,N_6920);
nand U7206 (N_7206,N_6853,N_6876);
nor U7207 (N_7207,N_6790,N_6879);
or U7208 (N_7208,N_6970,N_6923);
and U7209 (N_7209,N_6825,N_6773);
nand U7210 (N_7210,N_6785,N_6813);
and U7211 (N_7211,N_6854,N_6856);
nand U7212 (N_7212,N_6869,N_6943);
nor U7213 (N_7213,N_6780,N_6930);
nand U7214 (N_7214,N_6897,N_6767);
nor U7215 (N_7215,N_6818,N_6933);
nor U7216 (N_7216,N_6835,N_6922);
nor U7217 (N_7217,N_6845,N_6985);
nand U7218 (N_7218,N_6991,N_6905);
nor U7219 (N_7219,N_6979,N_6888);
xnor U7220 (N_7220,N_6996,N_6830);
or U7221 (N_7221,N_6831,N_6797);
nor U7222 (N_7222,N_6881,N_6948);
nand U7223 (N_7223,N_6753,N_6873);
nor U7224 (N_7224,N_6944,N_6942);
or U7225 (N_7225,N_6989,N_6769);
nor U7226 (N_7226,N_6779,N_6820);
or U7227 (N_7227,N_6879,N_6956);
xnor U7228 (N_7228,N_6928,N_6919);
and U7229 (N_7229,N_6791,N_6986);
nor U7230 (N_7230,N_6882,N_6891);
nor U7231 (N_7231,N_6803,N_6842);
nand U7232 (N_7232,N_6955,N_6929);
xnor U7233 (N_7233,N_6852,N_6838);
nand U7234 (N_7234,N_6993,N_6884);
nand U7235 (N_7235,N_6876,N_6933);
xor U7236 (N_7236,N_6888,N_6942);
nor U7237 (N_7237,N_6851,N_6841);
nand U7238 (N_7238,N_6802,N_6833);
nor U7239 (N_7239,N_6836,N_6820);
xor U7240 (N_7240,N_6944,N_6872);
xnor U7241 (N_7241,N_6879,N_6855);
and U7242 (N_7242,N_6965,N_6822);
or U7243 (N_7243,N_6992,N_6930);
xnor U7244 (N_7244,N_6874,N_6955);
nand U7245 (N_7245,N_6787,N_6902);
and U7246 (N_7246,N_6812,N_6999);
xnor U7247 (N_7247,N_6959,N_6828);
nor U7248 (N_7248,N_6949,N_6943);
nor U7249 (N_7249,N_6957,N_6826);
or U7250 (N_7250,N_7021,N_7114);
and U7251 (N_7251,N_7006,N_7004);
and U7252 (N_7252,N_7226,N_7040);
nor U7253 (N_7253,N_7228,N_7137);
nor U7254 (N_7254,N_7094,N_7118);
xor U7255 (N_7255,N_7144,N_7057);
nor U7256 (N_7256,N_7190,N_7056);
nor U7257 (N_7257,N_7107,N_7022);
and U7258 (N_7258,N_7038,N_7090);
xnor U7259 (N_7259,N_7216,N_7229);
nor U7260 (N_7260,N_7187,N_7073);
nand U7261 (N_7261,N_7115,N_7189);
and U7262 (N_7262,N_7150,N_7134);
or U7263 (N_7263,N_7001,N_7178);
nand U7264 (N_7264,N_7171,N_7025);
nand U7265 (N_7265,N_7087,N_7033);
nand U7266 (N_7266,N_7145,N_7047);
xnor U7267 (N_7267,N_7129,N_7132);
nand U7268 (N_7268,N_7084,N_7170);
and U7269 (N_7269,N_7097,N_7247);
and U7270 (N_7270,N_7059,N_7031);
or U7271 (N_7271,N_7089,N_7002);
and U7272 (N_7272,N_7063,N_7160);
nor U7273 (N_7273,N_7196,N_7074);
nand U7274 (N_7274,N_7220,N_7029);
xor U7275 (N_7275,N_7245,N_7199);
or U7276 (N_7276,N_7109,N_7015);
and U7277 (N_7277,N_7076,N_7218);
or U7278 (N_7278,N_7058,N_7205);
xor U7279 (N_7279,N_7206,N_7140);
and U7280 (N_7280,N_7186,N_7207);
or U7281 (N_7281,N_7127,N_7039);
and U7282 (N_7282,N_7148,N_7195);
nand U7283 (N_7283,N_7158,N_7176);
or U7284 (N_7284,N_7019,N_7035);
nand U7285 (N_7285,N_7085,N_7236);
nand U7286 (N_7286,N_7146,N_7156);
nand U7287 (N_7287,N_7111,N_7182);
nor U7288 (N_7288,N_7154,N_7070);
nor U7289 (N_7289,N_7221,N_7248);
or U7290 (N_7290,N_7163,N_7212);
nor U7291 (N_7291,N_7012,N_7069);
xor U7292 (N_7292,N_7183,N_7034);
or U7293 (N_7293,N_7143,N_7238);
nand U7294 (N_7294,N_7102,N_7222);
or U7295 (N_7295,N_7082,N_7005);
or U7296 (N_7296,N_7065,N_7214);
or U7297 (N_7297,N_7213,N_7008);
nor U7298 (N_7298,N_7028,N_7131);
and U7299 (N_7299,N_7055,N_7128);
nor U7300 (N_7300,N_7123,N_7242);
nand U7301 (N_7301,N_7067,N_7110);
nor U7302 (N_7302,N_7061,N_7233);
nor U7303 (N_7303,N_7036,N_7192);
or U7304 (N_7304,N_7016,N_7180);
nand U7305 (N_7305,N_7017,N_7091);
and U7306 (N_7306,N_7217,N_7112);
nand U7307 (N_7307,N_7049,N_7026);
and U7308 (N_7308,N_7209,N_7201);
nand U7309 (N_7309,N_7007,N_7133);
nor U7310 (N_7310,N_7193,N_7227);
or U7311 (N_7311,N_7009,N_7077);
or U7312 (N_7312,N_7052,N_7232);
nand U7313 (N_7313,N_7105,N_7080);
nand U7314 (N_7314,N_7153,N_7211);
nand U7315 (N_7315,N_7152,N_7174);
nand U7316 (N_7316,N_7185,N_7135);
nand U7317 (N_7317,N_7215,N_7043);
and U7318 (N_7318,N_7239,N_7202);
and U7319 (N_7319,N_7064,N_7027);
nand U7320 (N_7320,N_7151,N_7106);
or U7321 (N_7321,N_7249,N_7120);
nor U7322 (N_7322,N_7068,N_7023);
xnor U7323 (N_7323,N_7054,N_7060);
xnor U7324 (N_7324,N_7194,N_7030);
nor U7325 (N_7325,N_7096,N_7093);
nor U7326 (N_7326,N_7075,N_7121);
and U7327 (N_7327,N_7136,N_7173);
nor U7328 (N_7328,N_7237,N_7010);
and U7329 (N_7329,N_7081,N_7161);
or U7330 (N_7330,N_7032,N_7088);
and U7331 (N_7331,N_7020,N_7051);
xnor U7332 (N_7332,N_7204,N_7125);
and U7333 (N_7333,N_7165,N_7072);
or U7334 (N_7334,N_7142,N_7188);
xor U7335 (N_7335,N_7168,N_7104);
nor U7336 (N_7336,N_7157,N_7095);
nand U7337 (N_7337,N_7053,N_7224);
and U7338 (N_7338,N_7079,N_7141);
nand U7339 (N_7339,N_7138,N_7169);
or U7340 (N_7340,N_7045,N_7042);
xor U7341 (N_7341,N_7092,N_7162);
nor U7342 (N_7342,N_7197,N_7086);
and U7343 (N_7343,N_7122,N_7159);
nor U7344 (N_7344,N_7208,N_7100);
nand U7345 (N_7345,N_7003,N_7062);
nand U7346 (N_7346,N_7116,N_7099);
or U7347 (N_7347,N_7241,N_7014);
nor U7348 (N_7348,N_7243,N_7164);
and U7349 (N_7349,N_7223,N_7000);
or U7350 (N_7350,N_7044,N_7130);
nor U7351 (N_7351,N_7066,N_7246);
or U7352 (N_7352,N_7167,N_7198);
or U7353 (N_7353,N_7078,N_7108);
xor U7354 (N_7354,N_7050,N_7177);
and U7355 (N_7355,N_7083,N_7155);
and U7356 (N_7356,N_7230,N_7037);
and U7357 (N_7357,N_7124,N_7041);
and U7358 (N_7358,N_7126,N_7210);
and U7359 (N_7359,N_7225,N_7191);
nor U7360 (N_7360,N_7101,N_7219);
and U7361 (N_7361,N_7231,N_7203);
nor U7362 (N_7362,N_7048,N_7244);
and U7363 (N_7363,N_7166,N_7119);
or U7364 (N_7364,N_7071,N_7046);
nand U7365 (N_7365,N_7235,N_7011);
nor U7366 (N_7366,N_7184,N_7234);
or U7367 (N_7367,N_7200,N_7113);
nor U7368 (N_7368,N_7024,N_7175);
and U7369 (N_7369,N_7147,N_7181);
or U7370 (N_7370,N_7013,N_7117);
xor U7371 (N_7371,N_7172,N_7098);
nand U7372 (N_7372,N_7240,N_7139);
or U7373 (N_7373,N_7149,N_7018);
nor U7374 (N_7374,N_7179,N_7103);
and U7375 (N_7375,N_7175,N_7074);
nand U7376 (N_7376,N_7180,N_7188);
nor U7377 (N_7377,N_7116,N_7224);
nor U7378 (N_7378,N_7209,N_7013);
and U7379 (N_7379,N_7070,N_7134);
and U7380 (N_7380,N_7103,N_7227);
or U7381 (N_7381,N_7099,N_7043);
or U7382 (N_7382,N_7144,N_7032);
and U7383 (N_7383,N_7093,N_7149);
and U7384 (N_7384,N_7090,N_7100);
or U7385 (N_7385,N_7035,N_7056);
nor U7386 (N_7386,N_7013,N_7213);
and U7387 (N_7387,N_7153,N_7246);
nor U7388 (N_7388,N_7096,N_7053);
nor U7389 (N_7389,N_7185,N_7227);
nand U7390 (N_7390,N_7058,N_7038);
nand U7391 (N_7391,N_7214,N_7026);
nor U7392 (N_7392,N_7052,N_7177);
or U7393 (N_7393,N_7210,N_7041);
or U7394 (N_7394,N_7065,N_7225);
nand U7395 (N_7395,N_7156,N_7084);
nor U7396 (N_7396,N_7117,N_7014);
nand U7397 (N_7397,N_7088,N_7150);
xor U7398 (N_7398,N_7062,N_7045);
nor U7399 (N_7399,N_7063,N_7035);
xor U7400 (N_7400,N_7146,N_7158);
nand U7401 (N_7401,N_7181,N_7028);
and U7402 (N_7402,N_7018,N_7152);
or U7403 (N_7403,N_7154,N_7100);
xor U7404 (N_7404,N_7075,N_7126);
and U7405 (N_7405,N_7075,N_7021);
nand U7406 (N_7406,N_7238,N_7149);
or U7407 (N_7407,N_7153,N_7041);
or U7408 (N_7408,N_7016,N_7156);
nand U7409 (N_7409,N_7068,N_7086);
nand U7410 (N_7410,N_7194,N_7183);
and U7411 (N_7411,N_7209,N_7017);
or U7412 (N_7412,N_7068,N_7052);
nor U7413 (N_7413,N_7019,N_7119);
and U7414 (N_7414,N_7017,N_7016);
and U7415 (N_7415,N_7231,N_7007);
or U7416 (N_7416,N_7035,N_7163);
or U7417 (N_7417,N_7091,N_7082);
and U7418 (N_7418,N_7007,N_7025);
or U7419 (N_7419,N_7205,N_7019);
nor U7420 (N_7420,N_7064,N_7148);
nor U7421 (N_7421,N_7166,N_7127);
nand U7422 (N_7422,N_7143,N_7133);
xnor U7423 (N_7423,N_7061,N_7213);
or U7424 (N_7424,N_7185,N_7119);
or U7425 (N_7425,N_7042,N_7110);
or U7426 (N_7426,N_7183,N_7187);
nand U7427 (N_7427,N_7004,N_7186);
nand U7428 (N_7428,N_7041,N_7084);
and U7429 (N_7429,N_7021,N_7215);
xor U7430 (N_7430,N_7023,N_7026);
nor U7431 (N_7431,N_7066,N_7001);
nand U7432 (N_7432,N_7049,N_7059);
nor U7433 (N_7433,N_7000,N_7190);
or U7434 (N_7434,N_7187,N_7229);
nor U7435 (N_7435,N_7009,N_7125);
or U7436 (N_7436,N_7249,N_7248);
xor U7437 (N_7437,N_7036,N_7219);
nand U7438 (N_7438,N_7029,N_7216);
or U7439 (N_7439,N_7181,N_7170);
nand U7440 (N_7440,N_7127,N_7025);
nand U7441 (N_7441,N_7149,N_7044);
and U7442 (N_7442,N_7149,N_7203);
nor U7443 (N_7443,N_7200,N_7190);
and U7444 (N_7444,N_7152,N_7164);
or U7445 (N_7445,N_7116,N_7192);
or U7446 (N_7446,N_7067,N_7113);
nand U7447 (N_7447,N_7165,N_7016);
nor U7448 (N_7448,N_7166,N_7151);
and U7449 (N_7449,N_7093,N_7123);
xor U7450 (N_7450,N_7095,N_7026);
and U7451 (N_7451,N_7067,N_7152);
nand U7452 (N_7452,N_7242,N_7032);
or U7453 (N_7453,N_7137,N_7049);
and U7454 (N_7454,N_7159,N_7055);
and U7455 (N_7455,N_7137,N_7029);
nand U7456 (N_7456,N_7032,N_7139);
and U7457 (N_7457,N_7116,N_7103);
nand U7458 (N_7458,N_7173,N_7040);
nand U7459 (N_7459,N_7202,N_7063);
or U7460 (N_7460,N_7049,N_7108);
nor U7461 (N_7461,N_7233,N_7187);
nand U7462 (N_7462,N_7006,N_7153);
and U7463 (N_7463,N_7228,N_7083);
nand U7464 (N_7464,N_7226,N_7020);
and U7465 (N_7465,N_7218,N_7230);
or U7466 (N_7466,N_7193,N_7139);
nor U7467 (N_7467,N_7132,N_7155);
nand U7468 (N_7468,N_7058,N_7017);
xor U7469 (N_7469,N_7058,N_7108);
or U7470 (N_7470,N_7090,N_7216);
xnor U7471 (N_7471,N_7043,N_7220);
nand U7472 (N_7472,N_7142,N_7117);
and U7473 (N_7473,N_7009,N_7247);
nand U7474 (N_7474,N_7132,N_7221);
xnor U7475 (N_7475,N_7047,N_7014);
and U7476 (N_7476,N_7092,N_7201);
nand U7477 (N_7477,N_7214,N_7093);
nand U7478 (N_7478,N_7034,N_7207);
or U7479 (N_7479,N_7127,N_7032);
and U7480 (N_7480,N_7039,N_7177);
and U7481 (N_7481,N_7074,N_7102);
and U7482 (N_7482,N_7061,N_7002);
nor U7483 (N_7483,N_7104,N_7132);
nand U7484 (N_7484,N_7071,N_7007);
or U7485 (N_7485,N_7059,N_7003);
nor U7486 (N_7486,N_7053,N_7006);
nand U7487 (N_7487,N_7153,N_7060);
nand U7488 (N_7488,N_7060,N_7015);
xnor U7489 (N_7489,N_7016,N_7000);
or U7490 (N_7490,N_7247,N_7031);
xor U7491 (N_7491,N_7112,N_7248);
nor U7492 (N_7492,N_7064,N_7019);
nand U7493 (N_7493,N_7216,N_7031);
nor U7494 (N_7494,N_7166,N_7101);
and U7495 (N_7495,N_7114,N_7081);
nor U7496 (N_7496,N_7160,N_7059);
and U7497 (N_7497,N_7182,N_7024);
xnor U7498 (N_7498,N_7191,N_7206);
or U7499 (N_7499,N_7124,N_7128);
nand U7500 (N_7500,N_7314,N_7324);
xnor U7501 (N_7501,N_7494,N_7318);
and U7502 (N_7502,N_7355,N_7334);
or U7503 (N_7503,N_7276,N_7275);
nor U7504 (N_7504,N_7406,N_7498);
and U7505 (N_7505,N_7256,N_7317);
nor U7506 (N_7506,N_7356,N_7413);
nor U7507 (N_7507,N_7299,N_7313);
nand U7508 (N_7508,N_7367,N_7373);
or U7509 (N_7509,N_7452,N_7460);
nand U7510 (N_7510,N_7454,N_7496);
nand U7511 (N_7511,N_7285,N_7349);
or U7512 (N_7512,N_7487,N_7440);
or U7513 (N_7513,N_7370,N_7378);
and U7514 (N_7514,N_7469,N_7471);
and U7515 (N_7515,N_7403,N_7447);
and U7516 (N_7516,N_7300,N_7290);
and U7517 (N_7517,N_7338,N_7433);
nand U7518 (N_7518,N_7343,N_7353);
nor U7519 (N_7519,N_7473,N_7287);
nor U7520 (N_7520,N_7493,N_7253);
or U7521 (N_7521,N_7346,N_7341);
nor U7522 (N_7522,N_7280,N_7455);
and U7523 (N_7523,N_7436,N_7450);
nor U7524 (N_7524,N_7263,N_7303);
or U7525 (N_7525,N_7392,N_7427);
nand U7526 (N_7526,N_7422,N_7475);
or U7527 (N_7527,N_7265,N_7307);
nor U7528 (N_7528,N_7289,N_7292);
and U7529 (N_7529,N_7306,N_7371);
xor U7530 (N_7530,N_7463,N_7347);
and U7531 (N_7531,N_7309,N_7298);
xor U7532 (N_7532,N_7474,N_7368);
nor U7533 (N_7533,N_7363,N_7499);
nand U7534 (N_7534,N_7390,N_7385);
xor U7535 (N_7535,N_7483,N_7486);
nand U7536 (N_7536,N_7430,N_7325);
and U7537 (N_7537,N_7416,N_7372);
xnor U7538 (N_7538,N_7464,N_7485);
nand U7539 (N_7539,N_7308,N_7266);
nor U7540 (N_7540,N_7448,N_7302);
and U7541 (N_7541,N_7421,N_7376);
or U7542 (N_7542,N_7365,N_7412);
nand U7543 (N_7543,N_7418,N_7443);
nand U7544 (N_7544,N_7408,N_7482);
nor U7545 (N_7545,N_7260,N_7388);
and U7546 (N_7546,N_7488,N_7348);
nor U7547 (N_7547,N_7295,N_7261);
nor U7548 (N_7548,N_7304,N_7259);
nor U7549 (N_7549,N_7351,N_7291);
nor U7550 (N_7550,N_7366,N_7384);
and U7551 (N_7551,N_7262,N_7411);
or U7552 (N_7552,N_7352,N_7273);
xnor U7553 (N_7553,N_7432,N_7435);
and U7554 (N_7554,N_7495,N_7335);
and U7555 (N_7555,N_7453,N_7410);
and U7556 (N_7556,N_7284,N_7382);
nor U7557 (N_7557,N_7386,N_7319);
nand U7558 (N_7558,N_7254,N_7397);
xor U7559 (N_7559,N_7484,N_7380);
nor U7560 (N_7560,N_7394,N_7350);
xor U7561 (N_7561,N_7282,N_7288);
or U7562 (N_7562,N_7357,N_7477);
or U7563 (N_7563,N_7316,N_7420);
nand U7564 (N_7564,N_7322,N_7437);
or U7565 (N_7565,N_7294,N_7327);
and U7566 (N_7566,N_7362,N_7478);
or U7567 (N_7567,N_7497,N_7490);
and U7568 (N_7568,N_7400,N_7424);
nor U7569 (N_7569,N_7272,N_7377);
or U7570 (N_7570,N_7345,N_7333);
or U7571 (N_7571,N_7489,N_7438);
and U7572 (N_7572,N_7402,N_7344);
and U7573 (N_7573,N_7369,N_7328);
or U7574 (N_7574,N_7423,N_7399);
xor U7575 (N_7575,N_7451,N_7481);
nor U7576 (N_7576,N_7258,N_7431);
and U7577 (N_7577,N_7426,N_7360);
nor U7578 (N_7578,N_7342,N_7472);
or U7579 (N_7579,N_7264,N_7491);
nor U7580 (N_7580,N_7315,N_7329);
nand U7581 (N_7581,N_7359,N_7296);
or U7582 (N_7582,N_7268,N_7336);
or U7583 (N_7583,N_7323,N_7326);
nor U7584 (N_7584,N_7339,N_7251);
nor U7585 (N_7585,N_7414,N_7330);
and U7586 (N_7586,N_7281,N_7257);
and U7587 (N_7587,N_7465,N_7379);
or U7588 (N_7588,N_7405,N_7277);
nand U7589 (N_7589,N_7457,N_7337);
and U7590 (N_7590,N_7417,N_7270);
nor U7591 (N_7591,N_7415,N_7396);
nor U7592 (N_7592,N_7428,N_7391);
nor U7593 (N_7593,N_7429,N_7458);
xor U7594 (N_7594,N_7274,N_7267);
and U7595 (N_7595,N_7404,N_7279);
or U7596 (N_7596,N_7468,N_7381);
nand U7597 (N_7597,N_7383,N_7358);
or U7598 (N_7598,N_7444,N_7278);
xor U7599 (N_7599,N_7283,N_7434);
nand U7600 (N_7600,N_7340,N_7492);
nand U7601 (N_7601,N_7269,N_7393);
and U7602 (N_7602,N_7395,N_7459);
and U7603 (N_7603,N_7456,N_7476);
or U7604 (N_7604,N_7409,N_7301);
nor U7605 (N_7605,N_7331,N_7321);
nand U7606 (N_7606,N_7293,N_7419);
nor U7607 (N_7607,N_7480,N_7354);
or U7608 (N_7608,N_7364,N_7446);
nor U7609 (N_7609,N_7332,N_7305);
xor U7610 (N_7610,N_7425,N_7442);
and U7611 (N_7611,N_7467,N_7470);
nor U7612 (N_7612,N_7286,N_7255);
nand U7613 (N_7613,N_7387,N_7461);
or U7614 (N_7614,N_7312,N_7401);
and U7615 (N_7615,N_7375,N_7271);
nor U7616 (N_7616,N_7439,N_7462);
nand U7617 (N_7617,N_7320,N_7389);
nor U7618 (N_7618,N_7297,N_7466);
xnor U7619 (N_7619,N_7361,N_7250);
nor U7620 (N_7620,N_7407,N_7449);
and U7621 (N_7621,N_7252,N_7398);
or U7622 (N_7622,N_7374,N_7310);
xnor U7623 (N_7623,N_7311,N_7441);
nand U7624 (N_7624,N_7445,N_7479);
or U7625 (N_7625,N_7367,N_7330);
nor U7626 (N_7626,N_7320,N_7468);
or U7627 (N_7627,N_7355,N_7304);
nand U7628 (N_7628,N_7258,N_7419);
and U7629 (N_7629,N_7367,N_7288);
and U7630 (N_7630,N_7465,N_7357);
xor U7631 (N_7631,N_7436,N_7431);
nor U7632 (N_7632,N_7410,N_7280);
nor U7633 (N_7633,N_7462,N_7460);
or U7634 (N_7634,N_7439,N_7385);
or U7635 (N_7635,N_7446,N_7406);
nand U7636 (N_7636,N_7409,N_7267);
xnor U7637 (N_7637,N_7475,N_7326);
nand U7638 (N_7638,N_7347,N_7364);
nor U7639 (N_7639,N_7396,N_7440);
nor U7640 (N_7640,N_7371,N_7478);
nor U7641 (N_7641,N_7410,N_7282);
or U7642 (N_7642,N_7421,N_7321);
nor U7643 (N_7643,N_7261,N_7416);
nor U7644 (N_7644,N_7418,N_7383);
xnor U7645 (N_7645,N_7275,N_7390);
nor U7646 (N_7646,N_7260,N_7269);
xnor U7647 (N_7647,N_7400,N_7497);
nand U7648 (N_7648,N_7286,N_7448);
nand U7649 (N_7649,N_7322,N_7345);
xnor U7650 (N_7650,N_7365,N_7480);
and U7651 (N_7651,N_7439,N_7494);
nand U7652 (N_7652,N_7424,N_7379);
nor U7653 (N_7653,N_7329,N_7333);
and U7654 (N_7654,N_7404,N_7278);
nor U7655 (N_7655,N_7344,N_7355);
or U7656 (N_7656,N_7422,N_7458);
or U7657 (N_7657,N_7399,N_7444);
or U7658 (N_7658,N_7417,N_7271);
or U7659 (N_7659,N_7389,N_7358);
and U7660 (N_7660,N_7288,N_7335);
and U7661 (N_7661,N_7324,N_7498);
and U7662 (N_7662,N_7387,N_7275);
nand U7663 (N_7663,N_7478,N_7430);
and U7664 (N_7664,N_7371,N_7390);
nor U7665 (N_7665,N_7309,N_7472);
nand U7666 (N_7666,N_7251,N_7487);
xor U7667 (N_7667,N_7377,N_7420);
and U7668 (N_7668,N_7323,N_7444);
nor U7669 (N_7669,N_7410,N_7472);
xor U7670 (N_7670,N_7443,N_7444);
nand U7671 (N_7671,N_7481,N_7401);
and U7672 (N_7672,N_7490,N_7468);
and U7673 (N_7673,N_7298,N_7286);
xnor U7674 (N_7674,N_7397,N_7483);
nand U7675 (N_7675,N_7301,N_7278);
or U7676 (N_7676,N_7257,N_7443);
nand U7677 (N_7677,N_7350,N_7419);
nor U7678 (N_7678,N_7355,N_7305);
xnor U7679 (N_7679,N_7316,N_7304);
nand U7680 (N_7680,N_7284,N_7347);
and U7681 (N_7681,N_7327,N_7421);
nor U7682 (N_7682,N_7315,N_7481);
and U7683 (N_7683,N_7431,N_7481);
and U7684 (N_7684,N_7407,N_7360);
or U7685 (N_7685,N_7363,N_7468);
nand U7686 (N_7686,N_7440,N_7377);
xor U7687 (N_7687,N_7272,N_7311);
nor U7688 (N_7688,N_7441,N_7349);
nand U7689 (N_7689,N_7261,N_7434);
nor U7690 (N_7690,N_7273,N_7476);
and U7691 (N_7691,N_7252,N_7400);
nand U7692 (N_7692,N_7453,N_7333);
or U7693 (N_7693,N_7443,N_7263);
and U7694 (N_7694,N_7267,N_7492);
or U7695 (N_7695,N_7412,N_7359);
or U7696 (N_7696,N_7434,N_7421);
and U7697 (N_7697,N_7454,N_7480);
and U7698 (N_7698,N_7305,N_7495);
nand U7699 (N_7699,N_7262,N_7298);
and U7700 (N_7700,N_7494,N_7461);
or U7701 (N_7701,N_7308,N_7353);
nor U7702 (N_7702,N_7279,N_7488);
nand U7703 (N_7703,N_7340,N_7432);
and U7704 (N_7704,N_7280,N_7395);
nand U7705 (N_7705,N_7449,N_7426);
xnor U7706 (N_7706,N_7402,N_7371);
or U7707 (N_7707,N_7250,N_7362);
nor U7708 (N_7708,N_7435,N_7460);
nand U7709 (N_7709,N_7382,N_7250);
nor U7710 (N_7710,N_7406,N_7324);
nand U7711 (N_7711,N_7428,N_7325);
nor U7712 (N_7712,N_7284,N_7306);
nor U7713 (N_7713,N_7296,N_7429);
or U7714 (N_7714,N_7482,N_7464);
or U7715 (N_7715,N_7270,N_7290);
and U7716 (N_7716,N_7414,N_7327);
xor U7717 (N_7717,N_7338,N_7294);
xor U7718 (N_7718,N_7478,N_7391);
and U7719 (N_7719,N_7481,N_7385);
nand U7720 (N_7720,N_7417,N_7343);
nor U7721 (N_7721,N_7480,N_7415);
nand U7722 (N_7722,N_7395,N_7374);
nor U7723 (N_7723,N_7455,N_7364);
nand U7724 (N_7724,N_7489,N_7498);
nor U7725 (N_7725,N_7477,N_7348);
or U7726 (N_7726,N_7336,N_7258);
xnor U7727 (N_7727,N_7494,N_7284);
nor U7728 (N_7728,N_7343,N_7405);
nor U7729 (N_7729,N_7459,N_7336);
and U7730 (N_7730,N_7417,N_7447);
nor U7731 (N_7731,N_7494,N_7403);
and U7732 (N_7732,N_7317,N_7449);
and U7733 (N_7733,N_7340,N_7469);
nand U7734 (N_7734,N_7306,N_7301);
or U7735 (N_7735,N_7311,N_7259);
and U7736 (N_7736,N_7423,N_7392);
nor U7737 (N_7737,N_7263,N_7368);
and U7738 (N_7738,N_7479,N_7449);
or U7739 (N_7739,N_7320,N_7418);
nor U7740 (N_7740,N_7379,N_7268);
nand U7741 (N_7741,N_7471,N_7369);
xnor U7742 (N_7742,N_7313,N_7343);
or U7743 (N_7743,N_7406,N_7412);
nand U7744 (N_7744,N_7431,N_7292);
xnor U7745 (N_7745,N_7289,N_7434);
nand U7746 (N_7746,N_7294,N_7335);
and U7747 (N_7747,N_7400,N_7360);
or U7748 (N_7748,N_7364,N_7427);
and U7749 (N_7749,N_7379,N_7415);
and U7750 (N_7750,N_7697,N_7595);
or U7751 (N_7751,N_7607,N_7645);
nand U7752 (N_7752,N_7589,N_7629);
nor U7753 (N_7753,N_7503,N_7704);
nand U7754 (N_7754,N_7612,N_7513);
or U7755 (N_7755,N_7640,N_7530);
or U7756 (N_7756,N_7714,N_7743);
nand U7757 (N_7757,N_7570,N_7529);
nor U7758 (N_7758,N_7559,N_7680);
and U7759 (N_7759,N_7655,N_7539);
or U7760 (N_7760,N_7521,N_7730);
nor U7761 (N_7761,N_7581,N_7641);
nand U7762 (N_7762,N_7644,N_7511);
and U7763 (N_7763,N_7627,N_7542);
nor U7764 (N_7764,N_7574,N_7546);
nand U7765 (N_7765,N_7507,N_7715);
or U7766 (N_7766,N_7593,N_7667);
nand U7767 (N_7767,N_7603,N_7737);
or U7768 (N_7768,N_7558,N_7555);
or U7769 (N_7769,N_7693,N_7514);
nor U7770 (N_7770,N_7720,N_7648);
and U7771 (N_7771,N_7524,N_7748);
nor U7772 (N_7772,N_7545,N_7738);
xor U7773 (N_7773,N_7597,N_7668);
nand U7774 (N_7774,N_7518,N_7703);
nor U7775 (N_7775,N_7653,N_7532);
and U7776 (N_7776,N_7501,N_7652);
and U7777 (N_7777,N_7508,N_7531);
and U7778 (N_7778,N_7642,N_7684);
or U7779 (N_7779,N_7624,N_7636);
nor U7780 (N_7780,N_7585,N_7637);
nor U7781 (N_7781,N_7614,N_7575);
nand U7782 (N_7782,N_7660,N_7576);
nor U7783 (N_7783,N_7691,N_7553);
or U7784 (N_7784,N_7634,N_7600);
nand U7785 (N_7785,N_7541,N_7702);
nor U7786 (N_7786,N_7734,N_7599);
and U7787 (N_7787,N_7698,N_7661);
xnor U7788 (N_7788,N_7623,N_7618);
xor U7789 (N_7789,N_7708,N_7606);
xor U7790 (N_7790,N_7540,N_7538);
xor U7791 (N_7791,N_7741,N_7608);
and U7792 (N_7792,N_7650,N_7674);
nand U7793 (N_7793,N_7675,N_7617);
nor U7794 (N_7794,N_7745,N_7592);
nand U7795 (N_7795,N_7610,N_7727);
nor U7796 (N_7796,N_7632,N_7721);
or U7797 (N_7797,N_7573,N_7725);
nand U7798 (N_7798,N_7709,N_7579);
nand U7799 (N_7799,N_7525,N_7664);
or U7800 (N_7800,N_7515,N_7561);
and U7801 (N_7801,N_7519,N_7547);
and U7802 (N_7802,N_7517,N_7688);
nand U7803 (N_7803,N_7582,N_7583);
nand U7804 (N_7804,N_7662,N_7735);
nand U7805 (N_7805,N_7651,N_7732);
or U7806 (N_7806,N_7659,N_7695);
nor U7807 (N_7807,N_7685,N_7565);
or U7808 (N_7808,N_7520,N_7587);
xor U7809 (N_7809,N_7591,N_7686);
or U7810 (N_7810,N_7543,N_7628);
or U7811 (N_7811,N_7689,N_7718);
and U7812 (N_7812,N_7665,N_7504);
or U7813 (N_7813,N_7556,N_7669);
nand U7814 (N_7814,N_7588,N_7616);
nand U7815 (N_7815,N_7742,N_7649);
and U7816 (N_7816,N_7722,N_7699);
or U7817 (N_7817,N_7656,N_7707);
nor U7818 (N_7818,N_7749,N_7694);
xor U7819 (N_7819,N_7598,N_7569);
or U7820 (N_7820,N_7638,N_7554);
nand U7821 (N_7821,N_7673,N_7621);
xnor U7822 (N_7822,N_7671,N_7724);
or U7823 (N_7823,N_7550,N_7716);
and U7824 (N_7824,N_7590,N_7663);
nor U7825 (N_7825,N_7705,N_7647);
and U7826 (N_7826,N_7562,N_7571);
nand U7827 (N_7827,N_7620,N_7625);
nand U7828 (N_7828,N_7635,N_7700);
and U7829 (N_7829,N_7643,N_7526);
nand U7830 (N_7830,N_7633,N_7731);
nor U7831 (N_7831,N_7602,N_7596);
xor U7832 (N_7832,N_7717,N_7615);
xor U7833 (N_7833,N_7677,N_7577);
nor U7834 (N_7834,N_7601,N_7692);
nor U7835 (N_7835,N_7534,N_7564);
nor U7836 (N_7836,N_7605,N_7578);
nor U7837 (N_7837,N_7522,N_7523);
and U7838 (N_7838,N_7744,N_7683);
and U7839 (N_7839,N_7631,N_7622);
or U7840 (N_7840,N_7566,N_7657);
and U7841 (N_7841,N_7736,N_7563);
xor U7842 (N_7842,N_7676,N_7646);
nand U7843 (N_7843,N_7604,N_7711);
nor U7844 (N_7844,N_7533,N_7516);
nor U7845 (N_7845,N_7548,N_7696);
nand U7846 (N_7846,N_7505,N_7747);
and U7847 (N_7847,N_7681,N_7557);
nand U7848 (N_7848,N_7580,N_7594);
nor U7849 (N_7849,N_7512,N_7723);
nor U7850 (N_7850,N_7572,N_7733);
nor U7851 (N_7851,N_7670,N_7746);
or U7852 (N_7852,N_7568,N_7611);
and U7853 (N_7853,N_7506,N_7710);
nand U7854 (N_7854,N_7560,N_7679);
nor U7855 (N_7855,N_7619,N_7527);
nor U7856 (N_7856,N_7740,N_7502);
nor U7857 (N_7857,N_7672,N_7535);
and U7858 (N_7858,N_7609,N_7551);
nand U7859 (N_7859,N_7706,N_7626);
and U7860 (N_7860,N_7701,N_7613);
xor U7861 (N_7861,N_7552,N_7728);
nor U7862 (N_7862,N_7509,N_7528);
or U7863 (N_7863,N_7536,N_7654);
and U7864 (N_7864,N_7630,N_7687);
and U7865 (N_7865,N_7544,N_7678);
or U7866 (N_7866,N_7500,N_7739);
xor U7867 (N_7867,N_7658,N_7666);
nand U7868 (N_7868,N_7719,N_7584);
nor U7869 (N_7869,N_7713,N_7537);
nand U7870 (N_7870,N_7549,N_7690);
and U7871 (N_7871,N_7726,N_7729);
xnor U7872 (N_7872,N_7510,N_7682);
or U7873 (N_7873,N_7567,N_7712);
xnor U7874 (N_7874,N_7639,N_7586);
nor U7875 (N_7875,N_7679,N_7515);
xnor U7876 (N_7876,N_7732,N_7622);
or U7877 (N_7877,N_7722,N_7514);
nand U7878 (N_7878,N_7704,N_7666);
nor U7879 (N_7879,N_7600,N_7730);
or U7880 (N_7880,N_7719,N_7516);
and U7881 (N_7881,N_7562,N_7626);
and U7882 (N_7882,N_7500,N_7740);
nor U7883 (N_7883,N_7599,N_7675);
nand U7884 (N_7884,N_7538,N_7584);
nor U7885 (N_7885,N_7749,N_7564);
or U7886 (N_7886,N_7711,N_7692);
nand U7887 (N_7887,N_7580,N_7678);
or U7888 (N_7888,N_7612,N_7749);
nor U7889 (N_7889,N_7585,N_7525);
nor U7890 (N_7890,N_7617,N_7672);
nor U7891 (N_7891,N_7549,N_7561);
or U7892 (N_7892,N_7730,N_7718);
nand U7893 (N_7893,N_7586,N_7640);
nand U7894 (N_7894,N_7505,N_7625);
and U7895 (N_7895,N_7572,N_7688);
and U7896 (N_7896,N_7607,N_7647);
and U7897 (N_7897,N_7614,N_7737);
or U7898 (N_7898,N_7735,N_7708);
xnor U7899 (N_7899,N_7535,N_7653);
or U7900 (N_7900,N_7560,N_7600);
and U7901 (N_7901,N_7550,N_7612);
nor U7902 (N_7902,N_7515,N_7516);
and U7903 (N_7903,N_7607,N_7673);
and U7904 (N_7904,N_7664,N_7642);
nor U7905 (N_7905,N_7700,N_7537);
nand U7906 (N_7906,N_7647,N_7526);
nand U7907 (N_7907,N_7600,N_7697);
and U7908 (N_7908,N_7528,N_7749);
nor U7909 (N_7909,N_7652,N_7691);
xnor U7910 (N_7910,N_7653,N_7566);
xnor U7911 (N_7911,N_7551,N_7644);
nand U7912 (N_7912,N_7516,N_7617);
nand U7913 (N_7913,N_7607,N_7689);
or U7914 (N_7914,N_7729,N_7629);
nor U7915 (N_7915,N_7501,N_7654);
or U7916 (N_7916,N_7645,N_7535);
nand U7917 (N_7917,N_7725,N_7537);
xor U7918 (N_7918,N_7594,N_7503);
and U7919 (N_7919,N_7701,N_7669);
nor U7920 (N_7920,N_7688,N_7662);
nand U7921 (N_7921,N_7680,N_7560);
nand U7922 (N_7922,N_7554,N_7675);
or U7923 (N_7923,N_7500,N_7624);
and U7924 (N_7924,N_7593,N_7699);
xor U7925 (N_7925,N_7666,N_7605);
and U7926 (N_7926,N_7707,N_7738);
nor U7927 (N_7927,N_7669,N_7697);
xor U7928 (N_7928,N_7680,N_7695);
and U7929 (N_7929,N_7749,N_7729);
nor U7930 (N_7930,N_7675,N_7710);
nand U7931 (N_7931,N_7574,N_7571);
and U7932 (N_7932,N_7687,N_7731);
and U7933 (N_7933,N_7720,N_7522);
and U7934 (N_7934,N_7621,N_7575);
and U7935 (N_7935,N_7655,N_7727);
and U7936 (N_7936,N_7560,N_7668);
or U7937 (N_7937,N_7558,N_7615);
or U7938 (N_7938,N_7570,N_7604);
nand U7939 (N_7939,N_7686,N_7712);
nor U7940 (N_7940,N_7571,N_7747);
nand U7941 (N_7941,N_7718,N_7726);
nand U7942 (N_7942,N_7535,N_7722);
or U7943 (N_7943,N_7607,N_7542);
and U7944 (N_7944,N_7689,N_7519);
or U7945 (N_7945,N_7689,N_7501);
xor U7946 (N_7946,N_7615,N_7563);
nor U7947 (N_7947,N_7508,N_7577);
xor U7948 (N_7948,N_7580,N_7531);
nand U7949 (N_7949,N_7727,N_7699);
xnor U7950 (N_7950,N_7704,N_7555);
or U7951 (N_7951,N_7714,N_7591);
nor U7952 (N_7952,N_7538,N_7512);
and U7953 (N_7953,N_7719,N_7574);
nand U7954 (N_7954,N_7683,N_7685);
and U7955 (N_7955,N_7665,N_7563);
and U7956 (N_7956,N_7572,N_7625);
nand U7957 (N_7957,N_7514,N_7715);
nor U7958 (N_7958,N_7721,N_7521);
nor U7959 (N_7959,N_7696,N_7633);
xor U7960 (N_7960,N_7748,N_7580);
nand U7961 (N_7961,N_7691,N_7650);
xor U7962 (N_7962,N_7664,N_7515);
or U7963 (N_7963,N_7536,N_7684);
nand U7964 (N_7964,N_7619,N_7683);
or U7965 (N_7965,N_7637,N_7738);
xor U7966 (N_7966,N_7500,N_7598);
xor U7967 (N_7967,N_7625,N_7579);
or U7968 (N_7968,N_7513,N_7664);
xnor U7969 (N_7969,N_7725,N_7600);
and U7970 (N_7970,N_7556,N_7561);
and U7971 (N_7971,N_7659,N_7580);
and U7972 (N_7972,N_7627,N_7664);
and U7973 (N_7973,N_7505,N_7610);
nand U7974 (N_7974,N_7749,N_7716);
and U7975 (N_7975,N_7583,N_7683);
or U7976 (N_7976,N_7741,N_7601);
nor U7977 (N_7977,N_7579,N_7744);
or U7978 (N_7978,N_7587,N_7578);
nand U7979 (N_7979,N_7565,N_7697);
or U7980 (N_7980,N_7703,N_7657);
nor U7981 (N_7981,N_7524,N_7542);
nor U7982 (N_7982,N_7747,N_7726);
or U7983 (N_7983,N_7588,N_7609);
nand U7984 (N_7984,N_7539,N_7719);
nor U7985 (N_7985,N_7505,N_7708);
nor U7986 (N_7986,N_7561,N_7660);
and U7987 (N_7987,N_7716,N_7522);
nor U7988 (N_7988,N_7596,N_7608);
or U7989 (N_7989,N_7713,N_7699);
xor U7990 (N_7990,N_7614,N_7532);
and U7991 (N_7991,N_7718,N_7656);
nand U7992 (N_7992,N_7718,N_7707);
nand U7993 (N_7993,N_7618,N_7507);
and U7994 (N_7994,N_7605,N_7657);
nor U7995 (N_7995,N_7591,N_7534);
and U7996 (N_7996,N_7709,N_7521);
and U7997 (N_7997,N_7509,N_7553);
xnor U7998 (N_7998,N_7716,N_7567);
nand U7999 (N_7999,N_7629,N_7668);
and U8000 (N_8000,N_7834,N_7927);
and U8001 (N_8001,N_7928,N_7976);
nor U8002 (N_8002,N_7869,N_7915);
and U8003 (N_8003,N_7892,N_7874);
or U8004 (N_8004,N_7838,N_7996);
nand U8005 (N_8005,N_7905,N_7969);
or U8006 (N_8006,N_7978,N_7889);
nor U8007 (N_8007,N_7799,N_7858);
nor U8008 (N_8008,N_7902,N_7800);
nor U8009 (N_8009,N_7820,N_7998);
nand U8010 (N_8010,N_7796,N_7877);
or U8011 (N_8011,N_7842,N_7941);
nor U8012 (N_8012,N_7980,N_7752);
or U8013 (N_8013,N_7979,N_7822);
or U8014 (N_8014,N_7910,N_7772);
or U8015 (N_8015,N_7801,N_7984);
nor U8016 (N_8016,N_7992,N_7850);
nand U8017 (N_8017,N_7863,N_7895);
nand U8018 (N_8018,N_7964,N_7848);
or U8019 (N_8019,N_7782,N_7844);
or U8020 (N_8020,N_7898,N_7845);
xnor U8021 (N_8021,N_7788,N_7816);
nor U8022 (N_8022,N_7839,N_7954);
and U8023 (N_8023,N_7963,N_7826);
or U8024 (N_8024,N_7911,N_7950);
nor U8025 (N_8025,N_7878,N_7864);
or U8026 (N_8026,N_7897,N_7775);
nand U8027 (N_8027,N_7906,N_7994);
xor U8028 (N_8028,N_7764,N_7919);
nor U8029 (N_8029,N_7993,N_7935);
or U8030 (N_8030,N_7865,N_7870);
or U8031 (N_8031,N_7811,N_7912);
and U8032 (N_8032,N_7989,N_7991);
or U8033 (N_8033,N_7757,N_7968);
nor U8034 (N_8034,N_7948,N_7867);
xor U8035 (N_8035,N_7781,N_7854);
nand U8036 (N_8036,N_7824,N_7908);
and U8037 (N_8037,N_7828,N_7955);
and U8038 (N_8038,N_7756,N_7953);
nand U8039 (N_8039,N_7815,N_7841);
nand U8040 (N_8040,N_7923,N_7931);
nand U8041 (N_8041,N_7789,N_7967);
nor U8042 (N_8042,N_7862,N_7977);
and U8043 (N_8043,N_7766,N_7860);
xnor U8044 (N_8044,N_7833,N_7830);
or U8045 (N_8045,N_7888,N_7790);
or U8046 (N_8046,N_7804,N_7893);
and U8047 (N_8047,N_7840,N_7945);
and U8048 (N_8048,N_7872,N_7985);
and U8049 (N_8049,N_7783,N_7965);
nor U8050 (N_8050,N_7805,N_7988);
nor U8051 (N_8051,N_7939,N_7929);
and U8052 (N_8052,N_7938,N_7855);
xnor U8053 (N_8053,N_7852,N_7983);
nor U8054 (N_8054,N_7760,N_7932);
nand U8055 (N_8055,N_7982,N_7999);
nor U8056 (N_8056,N_7966,N_7847);
nor U8057 (N_8057,N_7827,N_7750);
or U8058 (N_8058,N_7777,N_7758);
nand U8059 (N_8059,N_7887,N_7930);
nand U8060 (N_8060,N_7916,N_7861);
nor U8061 (N_8061,N_7885,N_7890);
nor U8062 (N_8062,N_7934,N_7917);
nand U8063 (N_8063,N_7924,N_7856);
nand U8064 (N_8064,N_7880,N_7926);
nand U8065 (N_8065,N_7960,N_7975);
or U8066 (N_8066,N_7821,N_7785);
and U8067 (N_8067,N_7997,N_7794);
and U8068 (N_8068,N_7846,N_7761);
nand U8069 (N_8069,N_7900,N_7759);
nand U8070 (N_8070,N_7971,N_7894);
or U8071 (N_8071,N_7774,N_7798);
nor U8072 (N_8072,N_7810,N_7836);
xor U8073 (N_8073,N_7868,N_7891);
or U8074 (N_8074,N_7809,N_7883);
or U8075 (N_8075,N_7956,N_7763);
and U8076 (N_8076,N_7914,N_7973);
and U8077 (N_8077,N_7806,N_7918);
nor U8078 (N_8078,N_7871,N_7949);
nand U8079 (N_8079,N_7990,N_7831);
or U8080 (N_8080,N_7808,N_7857);
nand U8081 (N_8081,N_7778,N_7904);
and U8082 (N_8082,N_7936,N_7853);
nand U8083 (N_8083,N_7754,N_7951);
and U8084 (N_8084,N_7803,N_7921);
nand U8085 (N_8085,N_7959,N_7818);
nor U8086 (N_8086,N_7957,N_7769);
or U8087 (N_8087,N_7823,N_7768);
or U8088 (N_8088,N_7851,N_7802);
xor U8089 (N_8089,N_7755,N_7946);
and U8090 (N_8090,N_7962,N_7797);
nand U8091 (N_8091,N_7813,N_7765);
nand U8092 (N_8092,N_7792,N_7943);
and U8093 (N_8093,N_7812,N_7786);
and U8094 (N_8094,N_7753,N_7986);
nor U8095 (N_8095,N_7779,N_7995);
nand U8096 (N_8096,N_7884,N_7787);
nand U8097 (N_8097,N_7814,N_7767);
and U8098 (N_8098,N_7751,N_7817);
or U8099 (N_8099,N_7832,N_7940);
nor U8100 (N_8100,N_7922,N_7849);
or U8101 (N_8101,N_7901,N_7875);
and U8102 (N_8102,N_7952,N_7947);
or U8103 (N_8103,N_7907,N_7843);
and U8104 (N_8104,N_7795,N_7903);
nand U8105 (N_8105,N_7882,N_7920);
nand U8106 (N_8106,N_7961,N_7987);
nor U8107 (N_8107,N_7944,N_7762);
and U8108 (N_8108,N_7837,N_7819);
nor U8109 (N_8109,N_7825,N_7886);
xor U8110 (N_8110,N_7770,N_7958);
or U8111 (N_8111,N_7899,N_7793);
xor U8112 (N_8112,N_7972,N_7791);
or U8113 (N_8113,N_7807,N_7937);
xnor U8114 (N_8114,N_7876,N_7835);
nand U8115 (N_8115,N_7771,N_7896);
and U8116 (N_8116,N_7970,N_7909);
nor U8117 (N_8117,N_7776,N_7933);
nor U8118 (N_8118,N_7780,N_7974);
nand U8119 (N_8119,N_7942,N_7829);
nor U8120 (N_8120,N_7879,N_7784);
nand U8121 (N_8121,N_7913,N_7925);
nor U8122 (N_8122,N_7881,N_7866);
xor U8123 (N_8123,N_7859,N_7873);
xnor U8124 (N_8124,N_7981,N_7773);
and U8125 (N_8125,N_7929,N_7800);
or U8126 (N_8126,N_7780,N_7754);
or U8127 (N_8127,N_7832,N_7991);
nor U8128 (N_8128,N_7910,N_7758);
nor U8129 (N_8129,N_7837,N_7858);
nand U8130 (N_8130,N_7801,N_7888);
nor U8131 (N_8131,N_7833,N_7765);
xnor U8132 (N_8132,N_7766,N_7808);
and U8133 (N_8133,N_7867,N_7831);
and U8134 (N_8134,N_7836,N_7936);
nand U8135 (N_8135,N_7778,N_7897);
nand U8136 (N_8136,N_7861,N_7950);
nand U8137 (N_8137,N_7773,N_7982);
nor U8138 (N_8138,N_7970,N_7924);
nor U8139 (N_8139,N_7778,N_7783);
and U8140 (N_8140,N_7771,N_7997);
nor U8141 (N_8141,N_7903,N_7890);
xnor U8142 (N_8142,N_7940,N_7903);
xor U8143 (N_8143,N_7945,N_7815);
nand U8144 (N_8144,N_7807,N_7794);
and U8145 (N_8145,N_7980,N_7957);
or U8146 (N_8146,N_7974,N_7796);
nor U8147 (N_8147,N_7895,N_7762);
or U8148 (N_8148,N_7977,N_7799);
nand U8149 (N_8149,N_7824,N_7939);
or U8150 (N_8150,N_7873,N_7779);
nand U8151 (N_8151,N_7776,N_7982);
or U8152 (N_8152,N_7996,N_7866);
or U8153 (N_8153,N_7817,N_7972);
nand U8154 (N_8154,N_7762,N_7760);
nor U8155 (N_8155,N_7846,N_7870);
nor U8156 (N_8156,N_7871,N_7906);
or U8157 (N_8157,N_7834,N_7985);
nor U8158 (N_8158,N_7991,N_7847);
nor U8159 (N_8159,N_7816,N_7964);
nor U8160 (N_8160,N_7877,N_7992);
nor U8161 (N_8161,N_7901,N_7868);
or U8162 (N_8162,N_7925,N_7945);
and U8163 (N_8163,N_7759,N_7761);
xor U8164 (N_8164,N_7972,N_7921);
nand U8165 (N_8165,N_7943,N_7855);
and U8166 (N_8166,N_7941,N_7902);
xor U8167 (N_8167,N_7888,N_7796);
xnor U8168 (N_8168,N_7952,N_7791);
nand U8169 (N_8169,N_7848,N_7856);
nor U8170 (N_8170,N_7956,N_7809);
and U8171 (N_8171,N_7999,N_7968);
nor U8172 (N_8172,N_7826,N_7762);
or U8173 (N_8173,N_7834,N_7813);
or U8174 (N_8174,N_7773,N_7829);
nor U8175 (N_8175,N_7912,N_7804);
nand U8176 (N_8176,N_7924,N_7941);
or U8177 (N_8177,N_7901,N_7861);
or U8178 (N_8178,N_7986,N_7804);
or U8179 (N_8179,N_7968,N_7785);
or U8180 (N_8180,N_7983,N_7776);
xnor U8181 (N_8181,N_7843,N_7799);
and U8182 (N_8182,N_7782,N_7923);
nor U8183 (N_8183,N_7934,N_7940);
or U8184 (N_8184,N_7990,N_7847);
nor U8185 (N_8185,N_7989,N_7982);
and U8186 (N_8186,N_7826,N_7871);
nand U8187 (N_8187,N_7842,N_7795);
nand U8188 (N_8188,N_7753,N_7817);
nand U8189 (N_8189,N_7809,N_7993);
xnor U8190 (N_8190,N_7799,N_7912);
nand U8191 (N_8191,N_7851,N_7971);
and U8192 (N_8192,N_7780,N_7841);
xnor U8193 (N_8193,N_7835,N_7750);
nor U8194 (N_8194,N_7827,N_7787);
or U8195 (N_8195,N_7756,N_7982);
or U8196 (N_8196,N_7803,N_7939);
and U8197 (N_8197,N_7909,N_7975);
and U8198 (N_8198,N_7778,N_7815);
xnor U8199 (N_8199,N_7805,N_7917);
and U8200 (N_8200,N_7790,N_7894);
nor U8201 (N_8201,N_7954,N_7840);
nand U8202 (N_8202,N_7885,N_7916);
nand U8203 (N_8203,N_7880,N_7800);
and U8204 (N_8204,N_7834,N_7971);
nor U8205 (N_8205,N_7876,N_7938);
nor U8206 (N_8206,N_7850,N_7888);
and U8207 (N_8207,N_7867,N_7792);
xor U8208 (N_8208,N_7902,N_7778);
or U8209 (N_8209,N_7853,N_7966);
or U8210 (N_8210,N_7973,N_7759);
nor U8211 (N_8211,N_7758,N_7903);
nand U8212 (N_8212,N_7819,N_7884);
nand U8213 (N_8213,N_7834,N_7966);
xnor U8214 (N_8214,N_7811,N_7983);
and U8215 (N_8215,N_7753,N_7907);
nor U8216 (N_8216,N_7765,N_7899);
or U8217 (N_8217,N_7974,N_7956);
nand U8218 (N_8218,N_7821,N_7804);
nor U8219 (N_8219,N_7765,N_7967);
nand U8220 (N_8220,N_7786,N_7796);
nand U8221 (N_8221,N_7775,N_7902);
or U8222 (N_8222,N_7806,N_7930);
or U8223 (N_8223,N_7852,N_7930);
nor U8224 (N_8224,N_7835,N_7929);
or U8225 (N_8225,N_7930,N_7908);
nand U8226 (N_8226,N_7819,N_7898);
nand U8227 (N_8227,N_7854,N_7753);
or U8228 (N_8228,N_7869,N_7792);
or U8229 (N_8229,N_7785,N_7998);
nand U8230 (N_8230,N_7843,N_7873);
and U8231 (N_8231,N_7985,N_7899);
and U8232 (N_8232,N_7938,N_7929);
and U8233 (N_8233,N_7934,N_7986);
xor U8234 (N_8234,N_7879,N_7751);
and U8235 (N_8235,N_7817,N_7758);
nand U8236 (N_8236,N_7952,N_7860);
and U8237 (N_8237,N_7853,N_7873);
nand U8238 (N_8238,N_7811,N_7896);
nand U8239 (N_8239,N_7955,N_7836);
and U8240 (N_8240,N_7876,N_7889);
and U8241 (N_8241,N_7844,N_7883);
and U8242 (N_8242,N_7934,N_7833);
nand U8243 (N_8243,N_7946,N_7992);
or U8244 (N_8244,N_7922,N_7799);
nand U8245 (N_8245,N_7963,N_7774);
nor U8246 (N_8246,N_7872,N_7845);
xnor U8247 (N_8247,N_7752,N_7844);
nand U8248 (N_8248,N_7864,N_7857);
or U8249 (N_8249,N_7861,N_7893);
nand U8250 (N_8250,N_8028,N_8106);
and U8251 (N_8251,N_8161,N_8241);
and U8252 (N_8252,N_8011,N_8200);
nor U8253 (N_8253,N_8180,N_8187);
nand U8254 (N_8254,N_8160,N_8085);
nand U8255 (N_8255,N_8236,N_8232);
or U8256 (N_8256,N_8063,N_8091);
and U8257 (N_8257,N_8179,N_8052);
and U8258 (N_8258,N_8110,N_8002);
or U8259 (N_8259,N_8222,N_8000);
and U8260 (N_8260,N_8020,N_8165);
nor U8261 (N_8261,N_8005,N_8202);
nor U8262 (N_8262,N_8040,N_8051);
nand U8263 (N_8263,N_8074,N_8158);
and U8264 (N_8264,N_8134,N_8031);
and U8265 (N_8265,N_8095,N_8194);
and U8266 (N_8266,N_8188,N_8067);
and U8267 (N_8267,N_8159,N_8226);
nor U8268 (N_8268,N_8178,N_8077);
or U8269 (N_8269,N_8039,N_8141);
and U8270 (N_8270,N_8065,N_8054);
nor U8271 (N_8271,N_8068,N_8172);
nand U8272 (N_8272,N_8007,N_8173);
nor U8273 (N_8273,N_8092,N_8162);
nand U8274 (N_8274,N_8197,N_8125);
nand U8275 (N_8275,N_8151,N_8069);
nand U8276 (N_8276,N_8071,N_8216);
or U8277 (N_8277,N_8100,N_8073);
or U8278 (N_8278,N_8057,N_8088);
or U8279 (N_8279,N_8062,N_8212);
nand U8280 (N_8280,N_8131,N_8247);
and U8281 (N_8281,N_8220,N_8041);
nor U8282 (N_8282,N_8117,N_8083);
and U8283 (N_8283,N_8034,N_8013);
and U8284 (N_8284,N_8234,N_8227);
nand U8285 (N_8285,N_8029,N_8056);
xor U8286 (N_8286,N_8030,N_8006);
nor U8287 (N_8287,N_8219,N_8127);
nand U8288 (N_8288,N_8072,N_8102);
nand U8289 (N_8289,N_8199,N_8104);
or U8290 (N_8290,N_8167,N_8113);
nor U8291 (N_8291,N_8023,N_8132);
nand U8292 (N_8292,N_8093,N_8145);
or U8293 (N_8293,N_8025,N_8129);
or U8294 (N_8294,N_8055,N_8097);
and U8295 (N_8295,N_8017,N_8218);
and U8296 (N_8296,N_8205,N_8148);
nor U8297 (N_8297,N_8045,N_8012);
nand U8298 (N_8298,N_8246,N_8175);
nor U8299 (N_8299,N_8130,N_8208);
xor U8300 (N_8300,N_8243,N_8137);
xor U8301 (N_8301,N_8181,N_8024);
nor U8302 (N_8302,N_8064,N_8214);
or U8303 (N_8303,N_8115,N_8033);
nand U8304 (N_8304,N_8168,N_8107);
or U8305 (N_8305,N_8143,N_8231);
and U8306 (N_8306,N_8182,N_8174);
or U8307 (N_8307,N_8066,N_8036);
and U8308 (N_8308,N_8209,N_8101);
nor U8309 (N_8309,N_8108,N_8044);
xor U8310 (N_8310,N_8022,N_8230);
or U8311 (N_8311,N_8076,N_8223);
nand U8312 (N_8312,N_8103,N_8150);
or U8313 (N_8313,N_8001,N_8136);
nor U8314 (N_8314,N_8099,N_8164);
or U8315 (N_8315,N_8050,N_8058);
nor U8316 (N_8316,N_8035,N_8098);
xnor U8317 (N_8317,N_8154,N_8075);
nor U8318 (N_8318,N_8153,N_8018);
nand U8319 (N_8319,N_8242,N_8215);
nor U8320 (N_8320,N_8121,N_8133);
nor U8321 (N_8321,N_8149,N_8147);
and U8322 (N_8322,N_8163,N_8026);
nand U8323 (N_8323,N_8084,N_8116);
nand U8324 (N_8324,N_8217,N_8128);
nand U8325 (N_8325,N_8224,N_8244);
and U8326 (N_8326,N_8225,N_8176);
and U8327 (N_8327,N_8003,N_8221);
nand U8328 (N_8328,N_8139,N_8177);
or U8329 (N_8329,N_8112,N_8239);
nand U8330 (N_8330,N_8185,N_8032);
xnor U8331 (N_8331,N_8015,N_8123);
nand U8332 (N_8332,N_8211,N_8120);
or U8333 (N_8333,N_8037,N_8157);
and U8334 (N_8334,N_8027,N_8061);
or U8335 (N_8335,N_8248,N_8060);
and U8336 (N_8336,N_8048,N_8094);
nand U8337 (N_8337,N_8191,N_8043);
nand U8338 (N_8338,N_8195,N_8124);
nand U8339 (N_8339,N_8078,N_8118);
and U8340 (N_8340,N_8169,N_8019);
or U8341 (N_8341,N_8146,N_8122);
nand U8342 (N_8342,N_8237,N_8196);
nor U8343 (N_8343,N_8081,N_8190);
nand U8344 (N_8344,N_8119,N_8166);
xor U8345 (N_8345,N_8016,N_8142);
nand U8346 (N_8346,N_8171,N_8204);
or U8347 (N_8347,N_8046,N_8082);
nor U8348 (N_8348,N_8009,N_8152);
xnor U8349 (N_8349,N_8245,N_8126);
nand U8350 (N_8350,N_8086,N_8203);
or U8351 (N_8351,N_8087,N_8053);
or U8352 (N_8352,N_8014,N_8206);
and U8353 (N_8353,N_8189,N_8144);
nand U8354 (N_8354,N_8207,N_8109);
or U8355 (N_8355,N_8156,N_8047);
nor U8356 (N_8356,N_8021,N_8249);
nand U8357 (N_8357,N_8183,N_8186);
and U8358 (N_8358,N_8010,N_8089);
nor U8359 (N_8359,N_8235,N_8140);
nand U8360 (N_8360,N_8240,N_8090);
or U8361 (N_8361,N_8192,N_8184);
nand U8362 (N_8362,N_8038,N_8070);
and U8363 (N_8363,N_8138,N_8135);
or U8364 (N_8364,N_8201,N_8105);
nor U8365 (N_8365,N_8238,N_8228);
nor U8366 (N_8366,N_8198,N_8213);
and U8367 (N_8367,N_8080,N_8008);
nor U8368 (N_8368,N_8229,N_8170);
nand U8369 (N_8369,N_8059,N_8079);
and U8370 (N_8370,N_8004,N_8096);
xnor U8371 (N_8371,N_8114,N_8042);
or U8372 (N_8372,N_8111,N_8210);
xnor U8373 (N_8373,N_8233,N_8049);
nand U8374 (N_8374,N_8155,N_8193);
and U8375 (N_8375,N_8236,N_8153);
and U8376 (N_8376,N_8216,N_8247);
nor U8377 (N_8377,N_8193,N_8082);
nor U8378 (N_8378,N_8048,N_8122);
or U8379 (N_8379,N_8093,N_8193);
xnor U8380 (N_8380,N_8193,N_8072);
nand U8381 (N_8381,N_8166,N_8128);
and U8382 (N_8382,N_8133,N_8013);
and U8383 (N_8383,N_8051,N_8178);
nor U8384 (N_8384,N_8134,N_8132);
nor U8385 (N_8385,N_8216,N_8091);
nand U8386 (N_8386,N_8131,N_8160);
nor U8387 (N_8387,N_8029,N_8237);
nand U8388 (N_8388,N_8247,N_8179);
or U8389 (N_8389,N_8144,N_8127);
or U8390 (N_8390,N_8217,N_8178);
nand U8391 (N_8391,N_8004,N_8076);
nand U8392 (N_8392,N_8136,N_8095);
xor U8393 (N_8393,N_8043,N_8000);
nand U8394 (N_8394,N_8123,N_8022);
and U8395 (N_8395,N_8100,N_8239);
xor U8396 (N_8396,N_8035,N_8194);
and U8397 (N_8397,N_8056,N_8115);
and U8398 (N_8398,N_8239,N_8217);
nand U8399 (N_8399,N_8223,N_8015);
and U8400 (N_8400,N_8112,N_8187);
and U8401 (N_8401,N_8190,N_8217);
nand U8402 (N_8402,N_8134,N_8210);
or U8403 (N_8403,N_8135,N_8161);
or U8404 (N_8404,N_8050,N_8212);
nand U8405 (N_8405,N_8237,N_8009);
nor U8406 (N_8406,N_8085,N_8046);
nand U8407 (N_8407,N_8139,N_8169);
and U8408 (N_8408,N_8141,N_8070);
xnor U8409 (N_8409,N_8062,N_8112);
nor U8410 (N_8410,N_8122,N_8236);
or U8411 (N_8411,N_8220,N_8024);
nand U8412 (N_8412,N_8041,N_8013);
nor U8413 (N_8413,N_8193,N_8054);
and U8414 (N_8414,N_8191,N_8078);
nor U8415 (N_8415,N_8140,N_8133);
and U8416 (N_8416,N_8083,N_8188);
nor U8417 (N_8417,N_8057,N_8171);
nor U8418 (N_8418,N_8182,N_8204);
nand U8419 (N_8419,N_8097,N_8018);
nor U8420 (N_8420,N_8176,N_8206);
nor U8421 (N_8421,N_8110,N_8198);
nor U8422 (N_8422,N_8118,N_8180);
nor U8423 (N_8423,N_8066,N_8120);
and U8424 (N_8424,N_8018,N_8241);
or U8425 (N_8425,N_8151,N_8134);
nand U8426 (N_8426,N_8046,N_8107);
and U8427 (N_8427,N_8114,N_8117);
nand U8428 (N_8428,N_8046,N_8227);
nand U8429 (N_8429,N_8011,N_8003);
nor U8430 (N_8430,N_8088,N_8106);
xor U8431 (N_8431,N_8088,N_8103);
nand U8432 (N_8432,N_8088,N_8237);
and U8433 (N_8433,N_8048,N_8110);
or U8434 (N_8434,N_8008,N_8248);
nor U8435 (N_8435,N_8126,N_8113);
nand U8436 (N_8436,N_8052,N_8071);
nor U8437 (N_8437,N_8215,N_8131);
or U8438 (N_8438,N_8047,N_8244);
nand U8439 (N_8439,N_8148,N_8021);
and U8440 (N_8440,N_8132,N_8022);
nor U8441 (N_8441,N_8148,N_8045);
and U8442 (N_8442,N_8148,N_8163);
and U8443 (N_8443,N_8112,N_8070);
and U8444 (N_8444,N_8179,N_8110);
xor U8445 (N_8445,N_8109,N_8214);
nand U8446 (N_8446,N_8244,N_8246);
nor U8447 (N_8447,N_8211,N_8092);
or U8448 (N_8448,N_8208,N_8096);
xnor U8449 (N_8449,N_8106,N_8248);
or U8450 (N_8450,N_8153,N_8042);
or U8451 (N_8451,N_8239,N_8054);
and U8452 (N_8452,N_8236,N_8112);
xnor U8453 (N_8453,N_8195,N_8172);
nand U8454 (N_8454,N_8158,N_8193);
and U8455 (N_8455,N_8068,N_8185);
nor U8456 (N_8456,N_8057,N_8158);
nand U8457 (N_8457,N_8127,N_8145);
or U8458 (N_8458,N_8145,N_8097);
and U8459 (N_8459,N_8121,N_8105);
xnor U8460 (N_8460,N_8169,N_8213);
and U8461 (N_8461,N_8115,N_8049);
and U8462 (N_8462,N_8014,N_8229);
and U8463 (N_8463,N_8061,N_8113);
nor U8464 (N_8464,N_8035,N_8092);
and U8465 (N_8465,N_8203,N_8027);
nor U8466 (N_8466,N_8052,N_8108);
nand U8467 (N_8467,N_8007,N_8126);
xnor U8468 (N_8468,N_8128,N_8117);
and U8469 (N_8469,N_8104,N_8232);
or U8470 (N_8470,N_8127,N_8050);
nand U8471 (N_8471,N_8116,N_8115);
nor U8472 (N_8472,N_8138,N_8075);
xor U8473 (N_8473,N_8150,N_8156);
nand U8474 (N_8474,N_8185,N_8150);
nand U8475 (N_8475,N_8229,N_8114);
nand U8476 (N_8476,N_8055,N_8154);
nor U8477 (N_8477,N_8100,N_8054);
and U8478 (N_8478,N_8059,N_8128);
xor U8479 (N_8479,N_8243,N_8095);
nor U8480 (N_8480,N_8222,N_8183);
nor U8481 (N_8481,N_8210,N_8151);
nand U8482 (N_8482,N_8049,N_8183);
or U8483 (N_8483,N_8044,N_8171);
or U8484 (N_8484,N_8168,N_8157);
and U8485 (N_8485,N_8130,N_8166);
or U8486 (N_8486,N_8003,N_8185);
and U8487 (N_8487,N_8157,N_8215);
nor U8488 (N_8488,N_8038,N_8235);
or U8489 (N_8489,N_8173,N_8169);
or U8490 (N_8490,N_8242,N_8047);
nand U8491 (N_8491,N_8095,N_8019);
nor U8492 (N_8492,N_8007,N_8032);
and U8493 (N_8493,N_8103,N_8049);
nor U8494 (N_8494,N_8085,N_8089);
nor U8495 (N_8495,N_8242,N_8095);
nor U8496 (N_8496,N_8054,N_8018);
and U8497 (N_8497,N_8231,N_8087);
xnor U8498 (N_8498,N_8022,N_8140);
xnor U8499 (N_8499,N_8065,N_8085);
nor U8500 (N_8500,N_8449,N_8337);
nand U8501 (N_8501,N_8324,N_8321);
nor U8502 (N_8502,N_8290,N_8378);
nor U8503 (N_8503,N_8459,N_8494);
nand U8504 (N_8504,N_8358,N_8373);
and U8505 (N_8505,N_8316,N_8456);
nand U8506 (N_8506,N_8294,N_8278);
or U8507 (N_8507,N_8424,N_8377);
nor U8508 (N_8508,N_8437,N_8401);
nor U8509 (N_8509,N_8417,N_8491);
nand U8510 (N_8510,N_8385,N_8258);
and U8511 (N_8511,N_8260,N_8383);
xnor U8512 (N_8512,N_8404,N_8419);
nor U8513 (N_8513,N_8403,N_8416);
nand U8514 (N_8514,N_8349,N_8405);
and U8515 (N_8515,N_8472,N_8261);
or U8516 (N_8516,N_8473,N_8361);
or U8517 (N_8517,N_8259,N_8423);
nor U8518 (N_8518,N_8484,N_8394);
nand U8519 (N_8519,N_8395,N_8436);
nor U8520 (N_8520,N_8334,N_8276);
or U8521 (N_8521,N_8350,N_8285);
nor U8522 (N_8522,N_8289,N_8482);
or U8523 (N_8523,N_8270,N_8420);
nand U8524 (N_8524,N_8400,N_8384);
and U8525 (N_8525,N_8453,N_8267);
nor U8526 (N_8526,N_8268,N_8412);
nor U8527 (N_8527,N_8271,N_8431);
xor U8528 (N_8528,N_8365,N_8359);
or U8529 (N_8529,N_8310,N_8355);
and U8530 (N_8530,N_8388,N_8435);
nand U8531 (N_8531,N_8446,N_8425);
or U8532 (N_8532,N_8369,N_8256);
and U8533 (N_8533,N_8430,N_8280);
and U8534 (N_8534,N_8340,N_8477);
or U8535 (N_8535,N_8468,N_8342);
or U8536 (N_8536,N_8467,N_8432);
nor U8537 (N_8537,N_8406,N_8341);
nor U8538 (N_8538,N_8442,N_8462);
and U8539 (N_8539,N_8458,N_8262);
nor U8540 (N_8540,N_8486,N_8314);
xnor U8541 (N_8541,N_8252,N_8499);
nor U8542 (N_8542,N_8460,N_8371);
nand U8543 (N_8543,N_8269,N_8327);
or U8544 (N_8544,N_8360,N_8330);
nand U8545 (N_8545,N_8292,N_8346);
nor U8546 (N_8546,N_8318,N_8315);
or U8547 (N_8547,N_8376,N_8426);
and U8548 (N_8548,N_8387,N_8362);
or U8549 (N_8549,N_8332,N_8374);
nor U8550 (N_8550,N_8264,N_8463);
and U8551 (N_8551,N_8254,N_8303);
and U8552 (N_8552,N_8397,N_8380);
nand U8553 (N_8553,N_8287,N_8344);
nand U8554 (N_8554,N_8398,N_8296);
nor U8555 (N_8555,N_8301,N_8452);
or U8556 (N_8556,N_8345,N_8409);
nand U8557 (N_8557,N_8495,N_8338);
xnor U8558 (N_8558,N_8266,N_8393);
nor U8559 (N_8559,N_8288,N_8443);
nand U8560 (N_8560,N_8451,N_8354);
nor U8561 (N_8561,N_8323,N_8421);
nand U8562 (N_8562,N_8379,N_8311);
or U8563 (N_8563,N_8429,N_8312);
and U8564 (N_8564,N_8381,N_8480);
or U8565 (N_8565,N_8251,N_8366);
nand U8566 (N_8566,N_8336,N_8461);
or U8567 (N_8567,N_8402,N_8253);
and U8568 (N_8568,N_8319,N_8304);
nand U8569 (N_8569,N_8433,N_8447);
or U8570 (N_8570,N_8281,N_8367);
or U8571 (N_8571,N_8302,N_8471);
nor U8572 (N_8572,N_8438,N_8454);
or U8573 (N_8573,N_8368,N_8485);
nand U8574 (N_8574,N_8257,N_8396);
nor U8575 (N_8575,N_8291,N_8496);
nand U8576 (N_8576,N_8279,N_8493);
and U8577 (N_8577,N_8450,N_8487);
nor U8578 (N_8578,N_8283,N_8255);
nand U8579 (N_8579,N_8295,N_8466);
and U8580 (N_8580,N_8313,N_8414);
nor U8581 (N_8581,N_8434,N_8490);
and U8582 (N_8582,N_8422,N_8299);
or U8583 (N_8583,N_8474,N_8488);
nand U8584 (N_8584,N_8465,N_8320);
nand U8585 (N_8585,N_8326,N_8335);
or U8586 (N_8586,N_8386,N_8250);
nand U8587 (N_8587,N_8445,N_8439);
nand U8588 (N_8588,N_8455,N_8410);
xor U8589 (N_8589,N_8328,N_8444);
and U8590 (N_8590,N_8448,N_8317);
nor U8591 (N_8591,N_8489,N_8382);
or U8592 (N_8592,N_8322,N_8339);
xor U8593 (N_8593,N_8277,N_8356);
xor U8594 (N_8594,N_8305,N_8351);
nand U8595 (N_8595,N_8263,N_8352);
or U8596 (N_8596,N_8375,N_8427);
nor U8597 (N_8597,N_8333,N_8469);
nand U8598 (N_8598,N_8413,N_8478);
nand U8599 (N_8599,N_8411,N_8390);
nor U8600 (N_8600,N_8457,N_8329);
or U8601 (N_8601,N_8492,N_8440);
or U8602 (N_8602,N_8309,N_8307);
or U8603 (N_8603,N_8391,N_8274);
nand U8604 (N_8604,N_8286,N_8498);
nor U8605 (N_8605,N_8475,N_8483);
and U8606 (N_8606,N_8343,N_8325);
nand U8607 (N_8607,N_8298,N_8415);
nor U8608 (N_8608,N_8470,N_8407);
and U8609 (N_8609,N_8265,N_8300);
or U8610 (N_8610,N_8479,N_8481);
and U8611 (N_8611,N_8331,N_8464);
xnor U8612 (N_8612,N_8399,N_8297);
nor U8613 (N_8613,N_8441,N_8306);
or U8614 (N_8614,N_8347,N_8293);
nor U8615 (N_8615,N_8282,N_8272);
nand U8616 (N_8616,N_8275,N_8497);
nand U8617 (N_8617,N_8348,N_8408);
nand U8618 (N_8618,N_8372,N_8284);
nand U8619 (N_8619,N_8273,N_8418);
nor U8620 (N_8620,N_8308,N_8353);
and U8621 (N_8621,N_8364,N_8370);
or U8622 (N_8622,N_8389,N_8428);
or U8623 (N_8623,N_8476,N_8392);
and U8624 (N_8624,N_8363,N_8357);
nor U8625 (N_8625,N_8407,N_8380);
or U8626 (N_8626,N_8414,N_8295);
or U8627 (N_8627,N_8481,N_8346);
xnor U8628 (N_8628,N_8382,N_8477);
nor U8629 (N_8629,N_8291,N_8423);
and U8630 (N_8630,N_8433,N_8409);
xnor U8631 (N_8631,N_8451,N_8482);
nand U8632 (N_8632,N_8439,N_8314);
and U8633 (N_8633,N_8289,N_8479);
and U8634 (N_8634,N_8381,N_8266);
or U8635 (N_8635,N_8464,N_8337);
or U8636 (N_8636,N_8452,N_8258);
or U8637 (N_8637,N_8378,N_8351);
and U8638 (N_8638,N_8297,N_8351);
or U8639 (N_8639,N_8305,N_8490);
nor U8640 (N_8640,N_8393,N_8356);
and U8641 (N_8641,N_8455,N_8288);
nand U8642 (N_8642,N_8379,N_8302);
and U8643 (N_8643,N_8256,N_8451);
and U8644 (N_8644,N_8361,N_8414);
nor U8645 (N_8645,N_8352,N_8449);
nand U8646 (N_8646,N_8366,N_8294);
and U8647 (N_8647,N_8454,N_8322);
nand U8648 (N_8648,N_8336,N_8435);
and U8649 (N_8649,N_8252,N_8327);
nor U8650 (N_8650,N_8316,N_8292);
xor U8651 (N_8651,N_8439,N_8482);
or U8652 (N_8652,N_8430,N_8263);
nor U8653 (N_8653,N_8499,N_8313);
xnor U8654 (N_8654,N_8467,N_8469);
and U8655 (N_8655,N_8349,N_8367);
and U8656 (N_8656,N_8317,N_8461);
and U8657 (N_8657,N_8438,N_8397);
nand U8658 (N_8658,N_8277,N_8263);
and U8659 (N_8659,N_8447,N_8409);
and U8660 (N_8660,N_8464,N_8279);
or U8661 (N_8661,N_8437,N_8498);
and U8662 (N_8662,N_8475,N_8390);
nor U8663 (N_8663,N_8455,N_8361);
nand U8664 (N_8664,N_8252,N_8431);
nor U8665 (N_8665,N_8368,N_8413);
and U8666 (N_8666,N_8399,N_8413);
xnor U8667 (N_8667,N_8368,N_8375);
xnor U8668 (N_8668,N_8459,N_8416);
xnor U8669 (N_8669,N_8494,N_8401);
nor U8670 (N_8670,N_8334,N_8479);
and U8671 (N_8671,N_8336,N_8469);
nand U8672 (N_8672,N_8469,N_8345);
or U8673 (N_8673,N_8416,N_8462);
nor U8674 (N_8674,N_8459,N_8348);
nand U8675 (N_8675,N_8311,N_8395);
or U8676 (N_8676,N_8498,N_8363);
nor U8677 (N_8677,N_8280,N_8261);
nor U8678 (N_8678,N_8398,N_8266);
nand U8679 (N_8679,N_8416,N_8411);
nor U8680 (N_8680,N_8476,N_8281);
nor U8681 (N_8681,N_8446,N_8369);
nor U8682 (N_8682,N_8325,N_8412);
or U8683 (N_8683,N_8406,N_8424);
nand U8684 (N_8684,N_8391,N_8272);
xnor U8685 (N_8685,N_8309,N_8497);
or U8686 (N_8686,N_8377,N_8497);
and U8687 (N_8687,N_8479,N_8478);
and U8688 (N_8688,N_8277,N_8390);
nand U8689 (N_8689,N_8324,N_8355);
or U8690 (N_8690,N_8288,N_8419);
and U8691 (N_8691,N_8478,N_8331);
and U8692 (N_8692,N_8470,N_8301);
xor U8693 (N_8693,N_8253,N_8491);
nor U8694 (N_8694,N_8350,N_8412);
nand U8695 (N_8695,N_8361,N_8445);
and U8696 (N_8696,N_8493,N_8442);
and U8697 (N_8697,N_8496,N_8438);
or U8698 (N_8698,N_8465,N_8331);
or U8699 (N_8699,N_8343,N_8462);
nor U8700 (N_8700,N_8427,N_8460);
and U8701 (N_8701,N_8388,N_8260);
or U8702 (N_8702,N_8420,N_8252);
and U8703 (N_8703,N_8294,N_8323);
or U8704 (N_8704,N_8446,N_8274);
xor U8705 (N_8705,N_8416,N_8464);
nand U8706 (N_8706,N_8340,N_8278);
or U8707 (N_8707,N_8304,N_8294);
or U8708 (N_8708,N_8255,N_8495);
and U8709 (N_8709,N_8305,N_8273);
or U8710 (N_8710,N_8355,N_8490);
xnor U8711 (N_8711,N_8281,N_8270);
or U8712 (N_8712,N_8326,N_8499);
and U8713 (N_8713,N_8371,N_8461);
or U8714 (N_8714,N_8371,N_8339);
and U8715 (N_8715,N_8377,N_8389);
nor U8716 (N_8716,N_8358,N_8418);
nor U8717 (N_8717,N_8464,N_8399);
nand U8718 (N_8718,N_8351,N_8352);
nand U8719 (N_8719,N_8448,N_8467);
nor U8720 (N_8720,N_8250,N_8443);
nand U8721 (N_8721,N_8454,N_8448);
nand U8722 (N_8722,N_8320,N_8259);
nand U8723 (N_8723,N_8425,N_8304);
nor U8724 (N_8724,N_8419,N_8458);
nand U8725 (N_8725,N_8366,N_8288);
or U8726 (N_8726,N_8348,N_8490);
and U8727 (N_8727,N_8374,N_8443);
nand U8728 (N_8728,N_8381,N_8487);
xnor U8729 (N_8729,N_8461,N_8350);
nor U8730 (N_8730,N_8330,N_8384);
or U8731 (N_8731,N_8475,N_8292);
nor U8732 (N_8732,N_8452,N_8479);
nor U8733 (N_8733,N_8325,N_8310);
nand U8734 (N_8734,N_8378,N_8356);
and U8735 (N_8735,N_8419,N_8366);
and U8736 (N_8736,N_8328,N_8442);
nand U8737 (N_8737,N_8360,N_8310);
nor U8738 (N_8738,N_8368,N_8397);
or U8739 (N_8739,N_8359,N_8388);
and U8740 (N_8740,N_8286,N_8434);
nor U8741 (N_8741,N_8307,N_8356);
nand U8742 (N_8742,N_8341,N_8320);
or U8743 (N_8743,N_8429,N_8328);
and U8744 (N_8744,N_8371,N_8307);
or U8745 (N_8745,N_8452,N_8252);
and U8746 (N_8746,N_8348,N_8392);
or U8747 (N_8747,N_8283,N_8300);
nand U8748 (N_8748,N_8472,N_8419);
and U8749 (N_8749,N_8258,N_8428);
nand U8750 (N_8750,N_8679,N_8501);
nor U8751 (N_8751,N_8631,N_8709);
nand U8752 (N_8752,N_8684,N_8635);
nand U8753 (N_8753,N_8523,N_8680);
nor U8754 (N_8754,N_8639,N_8506);
nand U8755 (N_8755,N_8691,N_8651);
nor U8756 (N_8756,N_8510,N_8606);
or U8757 (N_8757,N_8749,N_8723);
or U8758 (N_8758,N_8740,N_8505);
and U8759 (N_8759,N_8683,N_8507);
and U8760 (N_8760,N_8634,N_8707);
nor U8761 (N_8761,N_8669,N_8736);
and U8762 (N_8762,N_8732,N_8554);
or U8763 (N_8763,N_8564,N_8706);
nor U8764 (N_8764,N_8672,N_8549);
nor U8765 (N_8765,N_8745,N_8689);
nor U8766 (N_8766,N_8663,N_8722);
nand U8767 (N_8767,N_8581,N_8734);
or U8768 (N_8768,N_8547,N_8648);
and U8769 (N_8769,N_8699,N_8571);
nand U8770 (N_8770,N_8644,N_8695);
and U8771 (N_8771,N_8696,N_8517);
nand U8772 (N_8772,N_8595,N_8608);
nand U8773 (N_8773,N_8519,N_8637);
nor U8774 (N_8774,N_8682,N_8604);
nand U8775 (N_8775,N_8530,N_8588);
xnor U8776 (N_8776,N_8605,N_8693);
nor U8777 (N_8777,N_8671,N_8703);
or U8778 (N_8778,N_8711,N_8526);
and U8779 (N_8779,N_8529,N_8552);
nor U8780 (N_8780,N_8642,N_8586);
xnor U8781 (N_8781,N_8565,N_8596);
nor U8782 (N_8782,N_8597,N_8576);
xnor U8783 (N_8783,N_8533,N_8551);
xnor U8784 (N_8784,N_8641,N_8717);
nor U8785 (N_8785,N_8583,N_8704);
nor U8786 (N_8786,N_8624,N_8666);
or U8787 (N_8787,N_8578,N_8591);
nor U8788 (N_8788,N_8603,N_8544);
nand U8789 (N_8789,N_8646,N_8582);
nor U8790 (N_8790,N_8559,N_8548);
or U8791 (N_8791,N_8725,N_8555);
nand U8792 (N_8792,N_8613,N_8710);
xnor U8793 (N_8793,N_8658,N_8527);
nor U8794 (N_8794,N_8744,N_8577);
or U8795 (N_8795,N_8649,N_8701);
and U8796 (N_8796,N_8626,N_8739);
or U8797 (N_8797,N_8513,N_8515);
nand U8798 (N_8798,N_8567,N_8667);
nor U8799 (N_8799,N_8538,N_8558);
and U8800 (N_8800,N_8676,N_8647);
nor U8801 (N_8801,N_8585,N_8569);
and U8802 (N_8802,N_8628,N_8503);
xor U8803 (N_8803,N_8747,N_8654);
and U8804 (N_8804,N_8623,N_8590);
nor U8805 (N_8805,N_8550,N_8620);
and U8806 (N_8806,N_8500,N_8625);
nor U8807 (N_8807,N_8668,N_8516);
or U8808 (N_8808,N_8617,N_8560);
or U8809 (N_8809,N_8720,N_8645);
nand U8810 (N_8810,N_8575,N_8580);
xnor U8811 (N_8811,N_8545,N_8528);
nor U8812 (N_8812,N_8661,N_8735);
or U8813 (N_8813,N_8543,N_8572);
or U8814 (N_8814,N_8686,N_8705);
nand U8815 (N_8815,N_8708,N_8630);
nor U8816 (N_8816,N_8643,N_8607);
xor U8817 (N_8817,N_8594,N_8601);
or U8818 (N_8818,N_8685,N_8562);
and U8819 (N_8819,N_8525,N_8633);
xnor U8820 (N_8820,N_8566,N_8598);
and U8821 (N_8821,N_8573,N_8593);
or U8822 (N_8822,N_8719,N_8553);
or U8823 (N_8823,N_8748,N_8531);
nand U8824 (N_8824,N_8638,N_8561);
nand U8825 (N_8825,N_8728,N_8713);
or U8826 (N_8826,N_8664,N_8539);
nand U8827 (N_8827,N_8502,N_8690);
and U8828 (N_8828,N_8688,N_8615);
nor U8829 (N_8829,N_8622,N_8694);
xnor U8830 (N_8830,N_8721,N_8737);
and U8831 (N_8831,N_8599,N_8640);
and U8832 (N_8832,N_8652,N_8592);
and U8833 (N_8833,N_8653,N_8512);
and U8834 (N_8834,N_8718,N_8662);
and U8835 (N_8835,N_8665,N_8697);
or U8836 (N_8836,N_8618,N_8504);
nand U8837 (N_8837,N_8675,N_8520);
nand U8838 (N_8838,N_8714,N_8521);
or U8839 (N_8839,N_8678,N_8535);
or U8840 (N_8840,N_8574,N_8698);
or U8841 (N_8841,N_8609,N_8570);
and U8842 (N_8842,N_8746,N_8579);
nor U8843 (N_8843,N_8587,N_8532);
or U8844 (N_8844,N_8632,N_8741);
or U8845 (N_8845,N_8738,N_8534);
nor U8846 (N_8846,N_8681,N_8656);
and U8847 (N_8847,N_8629,N_8568);
and U8848 (N_8848,N_8729,N_8659);
nand U8849 (N_8849,N_8674,N_8619);
nor U8850 (N_8850,N_8556,N_8610);
and U8851 (N_8851,N_8508,N_8509);
or U8852 (N_8852,N_8677,N_8700);
nand U8853 (N_8853,N_8542,N_8612);
and U8854 (N_8854,N_8524,N_8650);
and U8855 (N_8855,N_8726,N_8602);
and U8856 (N_8856,N_8673,N_8742);
nand U8857 (N_8857,N_8716,N_8692);
or U8858 (N_8858,N_8636,N_8731);
or U8859 (N_8859,N_8557,N_8621);
or U8860 (N_8860,N_8687,N_8727);
nand U8861 (N_8861,N_8611,N_8660);
or U8862 (N_8862,N_8743,N_8514);
nand U8863 (N_8863,N_8511,N_8712);
nand U8864 (N_8864,N_8657,N_8600);
xnor U8865 (N_8865,N_8537,N_8627);
and U8866 (N_8866,N_8655,N_8724);
nor U8867 (N_8867,N_8536,N_8546);
nand U8868 (N_8868,N_8589,N_8616);
nor U8869 (N_8869,N_8584,N_8540);
and U8870 (N_8870,N_8730,N_8715);
and U8871 (N_8871,N_8541,N_8670);
nor U8872 (N_8872,N_8563,N_8522);
nor U8873 (N_8873,N_8518,N_8702);
nor U8874 (N_8874,N_8614,N_8733);
nand U8875 (N_8875,N_8523,N_8726);
nand U8876 (N_8876,N_8543,N_8724);
and U8877 (N_8877,N_8639,N_8643);
and U8878 (N_8878,N_8595,N_8507);
nand U8879 (N_8879,N_8605,N_8500);
nor U8880 (N_8880,N_8711,N_8577);
nor U8881 (N_8881,N_8649,N_8512);
nand U8882 (N_8882,N_8629,N_8713);
and U8883 (N_8883,N_8597,N_8748);
and U8884 (N_8884,N_8575,N_8616);
and U8885 (N_8885,N_8580,N_8749);
xnor U8886 (N_8886,N_8708,N_8521);
nor U8887 (N_8887,N_8597,N_8630);
or U8888 (N_8888,N_8671,N_8660);
and U8889 (N_8889,N_8625,N_8504);
nand U8890 (N_8890,N_8521,N_8716);
xor U8891 (N_8891,N_8735,N_8580);
or U8892 (N_8892,N_8520,N_8580);
nor U8893 (N_8893,N_8679,N_8571);
nand U8894 (N_8894,N_8550,N_8658);
nand U8895 (N_8895,N_8563,N_8611);
nor U8896 (N_8896,N_8623,N_8661);
and U8897 (N_8897,N_8728,N_8738);
or U8898 (N_8898,N_8620,N_8603);
or U8899 (N_8899,N_8674,N_8590);
or U8900 (N_8900,N_8600,N_8652);
or U8901 (N_8901,N_8597,N_8588);
nor U8902 (N_8902,N_8528,N_8659);
nor U8903 (N_8903,N_8573,N_8543);
nor U8904 (N_8904,N_8621,N_8520);
nand U8905 (N_8905,N_8540,N_8603);
nand U8906 (N_8906,N_8720,N_8739);
nor U8907 (N_8907,N_8692,N_8544);
xor U8908 (N_8908,N_8679,N_8732);
xnor U8909 (N_8909,N_8667,N_8563);
or U8910 (N_8910,N_8705,N_8697);
and U8911 (N_8911,N_8619,N_8519);
nand U8912 (N_8912,N_8747,N_8658);
nor U8913 (N_8913,N_8613,N_8716);
and U8914 (N_8914,N_8619,N_8620);
nor U8915 (N_8915,N_8607,N_8586);
and U8916 (N_8916,N_8671,N_8675);
nor U8917 (N_8917,N_8698,N_8702);
and U8918 (N_8918,N_8723,N_8636);
and U8919 (N_8919,N_8511,N_8744);
xor U8920 (N_8920,N_8714,N_8533);
nor U8921 (N_8921,N_8626,N_8601);
nand U8922 (N_8922,N_8624,N_8513);
nand U8923 (N_8923,N_8599,N_8542);
or U8924 (N_8924,N_8525,N_8723);
and U8925 (N_8925,N_8686,N_8562);
or U8926 (N_8926,N_8652,N_8632);
or U8927 (N_8927,N_8500,N_8651);
and U8928 (N_8928,N_8506,N_8618);
and U8929 (N_8929,N_8728,N_8654);
or U8930 (N_8930,N_8592,N_8644);
and U8931 (N_8931,N_8647,N_8711);
nand U8932 (N_8932,N_8593,N_8540);
nand U8933 (N_8933,N_8609,N_8717);
xor U8934 (N_8934,N_8525,N_8695);
or U8935 (N_8935,N_8748,N_8652);
nor U8936 (N_8936,N_8509,N_8628);
and U8937 (N_8937,N_8590,N_8681);
xor U8938 (N_8938,N_8724,N_8590);
or U8939 (N_8939,N_8713,N_8611);
or U8940 (N_8940,N_8700,N_8643);
nand U8941 (N_8941,N_8714,N_8563);
and U8942 (N_8942,N_8558,N_8608);
nand U8943 (N_8943,N_8526,N_8523);
or U8944 (N_8944,N_8557,N_8503);
nor U8945 (N_8945,N_8714,N_8653);
nand U8946 (N_8946,N_8535,N_8623);
nand U8947 (N_8947,N_8715,N_8685);
nand U8948 (N_8948,N_8528,N_8673);
xor U8949 (N_8949,N_8639,N_8592);
and U8950 (N_8950,N_8694,N_8565);
and U8951 (N_8951,N_8748,N_8705);
nand U8952 (N_8952,N_8707,N_8551);
or U8953 (N_8953,N_8516,N_8732);
and U8954 (N_8954,N_8638,N_8651);
nand U8955 (N_8955,N_8671,N_8683);
nand U8956 (N_8956,N_8590,N_8553);
nor U8957 (N_8957,N_8688,N_8692);
and U8958 (N_8958,N_8618,N_8587);
nand U8959 (N_8959,N_8687,N_8538);
and U8960 (N_8960,N_8652,N_8660);
nand U8961 (N_8961,N_8512,N_8613);
or U8962 (N_8962,N_8703,N_8749);
nor U8963 (N_8963,N_8502,N_8565);
nor U8964 (N_8964,N_8536,N_8722);
nand U8965 (N_8965,N_8703,N_8721);
nand U8966 (N_8966,N_8554,N_8704);
and U8967 (N_8967,N_8648,N_8528);
nor U8968 (N_8968,N_8627,N_8591);
or U8969 (N_8969,N_8575,N_8604);
and U8970 (N_8970,N_8545,N_8518);
or U8971 (N_8971,N_8669,N_8659);
or U8972 (N_8972,N_8502,N_8701);
nor U8973 (N_8973,N_8748,N_8685);
nand U8974 (N_8974,N_8581,N_8714);
nand U8975 (N_8975,N_8675,N_8746);
nand U8976 (N_8976,N_8582,N_8608);
xor U8977 (N_8977,N_8711,N_8553);
and U8978 (N_8978,N_8544,N_8504);
or U8979 (N_8979,N_8685,N_8507);
nand U8980 (N_8980,N_8735,N_8593);
and U8981 (N_8981,N_8513,N_8569);
xor U8982 (N_8982,N_8533,N_8573);
nor U8983 (N_8983,N_8554,N_8709);
or U8984 (N_8984,N_8652,N_8651);
nand U8985 (N_8985,N_8560,N_8515);
nor U8986 (N_8986,N_8671,N_8508);
nor U8987 (N_8987,N_8634,N_8628);
or U8988 (N_8988,N_8574,N_8637);
or U8989 (N_8989,N_8631,N_8534);
nand U8990 (N_8990,N_8584,N_8515);
and U8991 (N_8991,N_8553,N_8743);
and U8992 (N_8992,N_8666,N_8553);
xor U8993 (N_8993,N_8623,N_8723);
and U8994 (N_8994,N_8673,N_8599);
nand U8995 (N_8995,N_8690,N_8707);
nor U8996 (N_8996,N_8698,N_8741);
and U8997 (N_8997,N_8608,N_8524);
and U8998 (N_8998,N_8657,N_8683);
or U8999 (N_8999,N_8505,N_8508);
and U9000 (N_9000,N_8987,N_8979);
xnor U9001 (N_9001,N_8822,N_8773);
and U9002 (N_9002,N_8946,N_8969);
nand U9003 (N_9003,N_8967,N_8999);
nor U9004 (N_9004,N_8845,N_8847);
or U9005 (N_9005,N_8952,N_8913);
nand U9006 (N_9006,N_8980,N_8947);
and U9007 (N_9007,N_8857,N_8977);
and U9008 (N_9008,N_8965,N_8821);
and U9009 (N_9009,N_8799,N_8852);
nand U9010 (N_9010,N_8992,N_8915);
xnor U9011 (N_9011,N_8775,N_8751);
and U9012 (N_9012,N_8990,N_8968);
and U9013 (N_9013,N_8837,N_8794);
nand U9014 (N_9014,N_8966,N_8762);
nor U9015 (N_9015,N_8875,N_8774);
nor U9016 (N_9016,N_8991,N_8940);
nand U9017 (N_9017,N_8939,N_8972);
nand U9018 (N_9018,N_8772,N_8783);
nand U9019 (N_9019,N_8923,N_8959);
and U9020 (N_9020,N_8846,N_8807);
and U9021 (N_9021,N_8872,N_8825);
and U9022 (N_9022,N_8973,N_8912);
nand U9023 (N_9023,N_8771,N_8860);
and U9024 (N_9024,N_8963,N_8817);
xor U9025 (N_9025,N_8917,N_8756);
and U9026 (N_9026,N_8922,N_8841);
and U9027 (N_9027,N_8752,N_8903);
and U9028 (N_9028,N_8826,N_8862);
and U9029 (N_9029,N_8948,N_8938);
and U9030 (N_9030,N_8865,N_8777);
xor U9031 (N_9031,N_8907,N_8827);
xnor U9032 (N_9032,N_8927,N_8871);
nand U9033 (N_9033,N_8882,N_8844);
nand U9034 (N_9034,N_8819,N_8881);
and U9035 (N_9035,N_8975,N_8905);
and U9036 (N_9036,N_8823,N_8893);
or U9037 (N_9037,N_8949,N_8970);
nand U9038 (N_9038,N_8870,N_8884);
nor U9039 (N_9039,N_8902,N_8850);
xor U9040 (N_9040,N_8820,N_8778);
nor U9041 (N_9041,N_8818,N_8957);
nand U9042 (N_9042,N_8754,N_8788);
nor U9043 (N_9043,N_8765,N_8998);
nand U9044 (N_9044,N_8802,N_8801);
and U9045 (N_9045,N_8876,N_8858);
nand U9046 (N_9046,N_8892,N_8839);
or U9047 (N_9047,N_8928,N_8945);
nand U9048 (N_9048,N_8950,N_8830);
nor U9049 (N_9049,N_8868,N_8925);
and U9050 (N_9050,N_8889,N_8853);
nand U9051 (N_9051,N_8758,N_8931);
and U9052 (N_9052,N_8908,N_8763);
and U9053 (N_9053,N_8986,N_8916);
nor U9054 (N_9054,N_8974,N_8842);
xor U9055 (N_9055,N_8981,N_8770);
and U9056 (N_9056,N_8929,N_8955);
nor U9057 (N_9057,N_8899,N_8909);
or U9058 (N_9058,N_8895,N_8937);
nor U9059 (N_9059,N_8795,N_8943);
nor U9060 (N_9060,N_8787,N_8835);
nand U9061 (N_9061,N_8873,N_8806);
or U9062 (N_9062,N_8918,N_8985);
nand U9063 (N_9063,N_8932,N_8869);
nor U9064 (N_9064,N_8798,N_8888);
nand U9065 (N_9065,N_8964,N_8800);
or U9066 (N_9066,N_8894,N_8933);
or U9067 (N_9067,N_8934,N_8956);
and U9068 (N_9068,N_8891,N_8936);
or U9069 (N_9069,N_8851,N_8759);
xor U9070 (N_9070,N_8811,N_8942);
nand U9071 (N_9071,N_8831,N_8780);
or U9072 (N_9072,N_8791,N_8878);
and U9073 (N_9073,N_8833,N_8886);
nor U9074 (N_9074,N_8988,N_8813);
nor U9075 (N_9075,N_8750,N_8815);
nand U9076 (N_9076,N_8867,N_8789);
nand U9077 (N_9077,N_8843,N_8782);
or U9078 (N_9078,N_8849,N_8834);
and U9079 (N_9079,N_8760,N_8824);
and U9080 (N_9080,N_8861,N_8761);
or U9081 (N_9081,N_8753,N_8962);
or U9082 (N_9082,N_8914,N_8983);
or U9083 (N_9083,N_8951,N_8994);
nand U9084 (N_9084,N_8890,N_8879);
or U9085 (N_9085,N_8785,N_8896);
and U9086 (N_9086,N_8809,N_8779);
nand U9087 (N_9087,N_8803,N_8814);
and U9088 (N_9088,N_8808,N_8920);
and U9089 (N_9089,N_8805,N_8828);
nand U9090 (N_9090,N_8816,N_8900);
nand U9091 (N_9091,N_8960,N_8995);
nor U9092 (N_9092,N_8784,N_8954);
and U9093 (N_9093,N_8953,N_8901);
and U9094 (N_9094,N_8769,N_8885);
and U9095 (N_9095,N_8887,N_8911);
nand U9096 (N_9096,N_8944,N_8978);
or U9097 (N_9097,N_8855,N_8792);
nand U9098 (N_9098,N_8919,N_8982);
or U9099 (N_9099,N_8921,N_8863);
nor U9100 (N_9100,N_8930,N_8781);
nand U9101 (N_9101,N_8904,N_8786);
nand U9102 (N_9102,N_8976,N_8848);
or U9103 (N_9103,N_8997,N_8961);
or U9104 (N_9104,N_8880,N_8859);
nand U9105 (N_9105,N_8883,N_8935);
nor U9106 (N_9106,N_8854,N_8790);
nand U9107 (N_9107,N_8864,N_8804);
nor U9108 (N_9108,N_8755,N_8958);
nand U9109 (N_9109,N_8797,N_8810);
nor U9110 (N_9110,N_8796,N_8924);
and U9111 (N_9111,N_8838,N_8764);
nor U9112 (N_9112,N_8984,N_8993);
nand U9113 (N_9113,N_8996,N_8989);
xor U9114 (N_9114,N_8941,N_8898);
nor U9115 (N_9115,N_8926,N_8906);
nor U9116 (N_9116,N_8832,N_8767);
nand U9117 (N_9117,N_8910,N_8793);
and U9118 (N_9118,N_8829,N_8768);
nand U9119 (N_9119,N_8757,N_8776);
nor U9120 (N_9120,N_8836,N_8840);
or U9121 (N_9121,N_8877,N_8971);
nand U9122 (N_9122,N_8856,N_8897);
or U9123 (N_9123,N_8766,N_8874);
nor U9124 (N_9124,N_8812,N_8866);
and U9125 (N_9125,N_8823,N_8861);
or U9126 (N_9126,N_8877,N_8755);
nor U9127 (N_9127,N_8975,N_8944);
or U9128 (N_9128,N_8900,N_8861);
nor U9129 (N_9129,N_8983,N_8821);
nor U9130 (N_9130,N_8857,N_8932);
nand U9131 (N_9131,N_8875,N_8892);
and U9132 (N_9132,N_8822,N_8879);
or U9133 (N_9133,N_8900,N_8844);
xor U9134 (N_9134,N_8832,N_8818);
nand U9135 (N_9135,N_8851,N_8804);
and U9136 (N_9136,N_8841,N_8986);
and U9137 (N_9137,N_8838,N_8950);
nor U9138 (N_9138,N_8820,N_8895);
and U9139 (N_9139,N_8934,N_8921);
nor U9140 (N_9140,N_8838,N_8983);
nor U9141 (N_9141,N_8881,N_8754);
nand U9142 (N_9142,N_8950,N_8824);
xor U9143 (N_9143,N_8778,N_8993);
nor U9144 (N_9144,N_8889,N_8981);
and U9145 (N_9145,N_8789,N_8901);
nor U9146 (N_9146,N_8952,N_8934);
and U9147 (N_9147,N_8971,N_8929);
xnor U9148 (N_9148,N_8753,N_8958);
nand U9149 (N_9149,N_8851,N_8971);
xor U9150 (N_9150,N_8858,N_8869);
nor U9151 (N_9151,N_8821,N_8809);
or U9152 (N_9152,N_8866,N_8805);
nor U9153 (N_9153,N_8759,N_8775);
and U9154 (N_9154,N_8769,N_8936);
and U9155 (N_9155,N_8978,N_8949);
nand U9156 (N_9156,N_8849,N_8782);
nor U9157 (N_9157,N_8864,N_8849);
and U9158 (N_9158,N_8764,N_8983);
nand U9159 (N_9159,N_8809,N_8892);
xnor U9160 (N_9160,N_8775,N_8839);
nor U9161 (N_9161,N_8796,N_8975);
xor U9162 (N_9162,N_8980,N_8906);
and U9163 (N_9163,N_8932,N_8844);
nor U9164 (N_9164,N_8965,N_8789);
and U9165 (N_9165,N_8771,N_8872);
nand U9166 (N_9166,N_8915,N_8810);
or U9167 (N_9167,N_8814,N_8788);
xor U9168 (N_9168,N_8928,N_8876);
and U9169 (N_9169,N_8906,N_8856);
nor U9170 (N_9170,N_8957,N_8854);
nand U9171 (N_9171,N_8947,N_8787);
nor U9172 (N_9172,N_8852,N_8802);
xnor U9173 (N_9173,N_8867,N_8934);
nand U9174 (N_9174,N_8982,N_8777);
xor U9175 (N_9175,N_8785,N_8973);
and U9176 (N_9176,N_8980,N_8784);
nor U9177 (N_9177,N_8859,N_8874);
nand U9178 (N_9178,N_8966,N_8792);
nand U9179 (N_9179,N_8980,N_8956);
nand U9180 (N_9180,N_8960,N_8973);
nor U9181 (N_9181,N_8943,N_8961);
or U9182 (N_9182,N_8845,N_8778);
or U9183 (N_9183,N_8955,N_8916);
and U9184 (N_9184,N_8934,N_8932);
nor U9185 (N_9185,N_8816,N_8893);
xnor U9186 (N_9186,N_8886,N_8793);
xnor U9187 (N_9187,N_8996,N_8892);
or U9188 (N_9188,N_8966,N_8980);
nor U9189 (N_9189,N_8993,N_8825);
or U9190 (N_9190,N_8761,N_8793);
and U9191 (N_9191,N_8875,N_8807);
nor U9192 (N_9192,N_8777,N_8866);
nand U9193 (N_9193,N_8750,N_8937);
or U9194 (N_9194,N_8782,N_8975);
or U9195 (N_9195,N_8938,N_8813);
xor U9196 (N_9196,N_8975,N_8967);
or U9197 (N_9197,N_8885,N_8961);
nand U9198 (N_9198,N_8784,N_8807);
xnor U9199 (N_9199,N_8828,N_8793);
nand U9200 (N_9200,N_8997,N_8914);
or U9201 (N_9201,N_8939,N_8778);
or U9202 (N_9202,N_8782,N_8930);
or U9203 (N_9203,N_8868,N_8796);
xor U9204 (N_9204,N_8969,N_8810);
and U9205 (N_9205,N_8821,N_8777);
xor U9206 (N_9206,N_8848,N_8767);
or U9207 (N_9207,N_8976,N_8985);
or U9208 (N_9208,N_8868,N_8814);
or U9209 (N_9209,N_8914,N_8878);
and U9210 (N_9210,N_8808,N_8818);
nand U9211 (N_9211,N_8854,N_8974);
xor U9212 (N_9212,N_8910,N_8999);
nor U9213 (N_9213,N_8924,N_8757);
nor U9214 (N_9214,N_8772,N_8900);
and U9215 (N_9215,N_8797,N_8801);
and U9216 (N_9216,N_8791,N_8818);
nand U9217 (N_9217,N_8900,N_8817);
xnor U9218 (N_9218,N_8856,N_8865);
nor U9219 (N_9219,N_8952,N_8964);
nand U9220 (N_9220,N_8836,N_8889);
nand U9221 (N_9221,N_8931,N_8767);
nand U9222 (N_9222,N_8769,N_8796);
and U9223 (N_9223,N_8954,N_8842);
nor U9224 (N_9224,N_8968,N_8917);
nor U9225 (N_9225,N_8860,N_8839);
and U9226 (N_9226,N_8758,N_8981);
or U9227 (N_9227,N_8948,N_8757);
nor U9228 (N_9228,N_8975,N_8823);
xor U9229 (N_9229,N_8832,N_8940);
nand U9230 (N_9230,N_8970,N_8941);
nand U9231 (N_9231,N_8919,N_8921);
nor U9232 (N_9232,N_8907,N_8901);
and U9233 (N_9233,N_8896,N_8983);
nor U9234 (N_9234,N_8762,N_8935);
nand U9235 (N_9235,N_8989,N_8857);
nand U9236 (N_9236,N_8836,N_8892);
nor U9237 (N_9237,N_8848,N_8922);
or U9238 (N_9238,N_8810,N_8809);
or U9239 (N_9239,N_8904,N_8770);
nor U9240 (N_9240,N_8987,N_8888);
and U9241 (N_9241,N_8892,N_8857);
or U9242 (N_9242,N_8971,N_8867);
nand U9243 (N_9243,N_8899,N_8941);
or U9244 (N_9244,N_8908,N_8903);
and U9245 (N_9245,N_8914,N_8988);
and U9246 (N_9246,N_8987,N_8881);
or U9247 (N_9247,N_8854,N_8895);
or U9248 (N_9248,N_8920,N_8908);
or U9249 (N_9249,N_8785,N_8862);
nor U9250 (N_9250,N_9181,N_9024);
nor U9251 (N_9251,N_9071,N_9136);
nand U9252 (N_9252,N_9065,N_9089);
xor U9253 (N_9253,N_9000,N_9111);
nand U9254 (N_9254,N_9161,N_9045);
nor U9255 (N_9255,N_9222,N_9162);
xnor U9256 (N_9256,N_9150,N_9060);
or U9257 (N_9257,N_9221,N_9123);
nor U9258 (N_9258,N_9068,N_9105);
nand U9259 (N_9259,N_9114,N_9242);
nand U9260 (N_9260,N_9048,N_9165);
nor U9261 (N_9261,N_9056,N_9118);
and U9262 (N_9262,N_9113,N_9037);
nor U9263 (N_9263,N_9189,N_9217);
or U9264 (N_9264,N_9128,N_9053);
nand U9265 (N_9265,N_9127,N_9085);
nor U9266 (N_9266,N_9104,N_9244);
nand U9267 (N_9267,N_9173,N_9070);
nor U9268 (N_9268,N_9015,N_9022);
nand U9269 (N_9269,N_9094,N_9072);
xnor U9270 (N_9270,N_9036,N_9207);
nand U9271 (N_9271,N_9112,N_9144);
nor U9272 (N_9272,N_9027,N_9204);
nor U9273 (N_9273,N_9023,N_9038);
nor U9274 (N_9274,N_9223,N_9074);
nand U9275 (N_9275,N_9055,N_9176);
nor U9276 (N_9276,N_9168,N_9021);
and U9277 (N_9277,N_9073,N_9218);
and U9278 (N_9278,N_9014,N_9077);
and U9279 (N_9279,N_9028,N_9232);
and U9280 (N_9280,N_9140,N_9248);
or U9281 (N_9281,N_9109,N_9210);
nand U9282 (N_9282,N_9230,N_9231);
nor U9283 (N_9283,N_9097,N_9175);
nor U9284 (N_9284,N_9209,N_9115);
and U9285 (N_9285,N_9198,N_9029);
nand U9286 (N_9286,N_9069,N_9083);
nand U9287 (N_9287,N_9125,N_9229);
or U9288 (N_9288,N_9146,N_9008);
nor U9289 (N_9289,N_9110,N_9228);
nand U9290 (N_9290,N_9117,N_9092);
and U9291 (N_9291,N_9195,N_9238);
nor U9292 (N_9292,N_9017,N_9066);
or U9293 (N_9293,N_9169,N_9177);
and U9294 (N_9294,N_9001,N_9216);
nand U9295 (N_9295,N_9172,N_9167);
xnor U9296 (N_9296,N_9240,N_9103);
and U9297 (N_9297,N_9050,N_9180);
or U9298 (N_9298,N_9011,N_9234);
nand U9299 (N_9299,N_9211,N_9208);
or U9300 (N_9300,N_9200,N_9163);
nand U9301 (N_9301,N_9054,N_9081);
nand U9302 (N_9302,N_9026,N_9202);
nor U9303 (N_9303,N_9170,N_9057);
nand U9304 (N_9304,N_9199,N_9035);
nand U9305 (N_9305,N_9033,N_9213);
xnor U9306 (N_9306,N_9133,N_9122);
or U9307 (N_9307,N_9201,N_9040);
or U9308 (N_9308,N_9062,N_9061);
nand U9309 (N_9309,N_9143,N_9154);
and U9310 (N_9310,N_9239,N_9149);
or U9311 (N_9311,N_9119,N_9020);
and U9312 (N_9312,N_9013,N_9205);
and U9313 (N_9313,N_9031,N_9091);
or U9314 (N_9314,N_9245,N_9043);
and U9315 (N_9315,N_9241,N_9005);
nor U9316 (N_9316,N_9009,N_9227);
nand U9317 (N_9317,N_9134,N_9039);
and U9318 (N_9318,N_9183,N_9247);
and U9319 (N_9319,N_9206,N_9166);
nor U9320 (N_9320,N_9246,N_9160);
nand U9321 (N_9321,N_9093,N_9156);
and U9322 (N_9322,N_9203,N_9196);
and U9323 (N_9323,N_9137,N_9191);
or U9324 (N_9324,N_9012,N_9032);
and U9325 (N_9325,N_9116,N_9030);
or U9326 (N_9326,N_9059,N_9100);
nand U9327 (N_9327,N_9010,N_9025);
and U9328 (N_9328,N_9226,N_9046);
nand U9329 (N_9329,N_9047,N_9186);
xnor U9330 (N_9330,N_9124,N_9016);
nand U9331 (N_9331,N_9159,N_9184);
xnor U9332 (N_9332,N_9132,N_9214);
and U9333 (N_9333,N_9224,N_9084);
nor U9334 (N_9334,N_9237,N_9096);
nand U9335 (N_9335,N_9235,N_9138);
nor U9336 (N_9336,N_9004,N_9108);
and U9337 (N_9337,N_9148,N_9076);
xnor U9338 (N_9338,N_9106,N_9190);
and U9339 (N_9339,N_9041,N_9233);
and U9340 (N_9340,N_9236,N_9193);
nand U9341 (N_9341,N_9178,N_9019);
nand U9342 (N_9342,N_9052,N_9007);
or U9343 (N_9343,N_9147,N_9042);
xnor U9344 (N_9344,N_9157,N_9135);
and U9345 (N_9345,N_9212,N_9142);
nand U9346 (N_9346,N_9155,N_9129);
nor U9347 (N_9347,N_9063,N_9139);
and U9348 (N_9348,N_9145,N_9087);
xnor U9349 (N_9349,N_9130,N_9194);
nor U9350 (N_9350,N_9088,N_9192);
nor U9351 (N_9351,N_9095,N_9243);
and U9352 (N_9352,N_9171,N_9099);
and U9353 (N_9353,N_9121,N_9220);
or U9354 (N_9354,N_9002,N_9075);
nand U9355 (N_9355,N_9179,N_9141);
nor U9356 (N_9356,N_9120,N_9086);
nand U9357 (N_9357,N_9080,N_9102);
xor U9358 (N_9358,N_9003,N_9131);
and U9359 (N_9359,N_9018,N_9090);
or U9360 (N_9360,N_9249,N_9064);
or U9361 (N_9361,N_9152,N_9051);
nand U9362 (N_9362,N_9219,N_9174);
and U9363 (N_9363,N_9107,N_9182);
and U9364 (N_9364,N_9034,N_9079);
nor U9365 (N_9365,N_9098,N_9225);
xnor U9366 (N_9366,N_9197,N_9187);
and U9367 (N_9367,N_9164,N_9126);
or U9368 (N_9368,N_9101,N_9006);
xnor U9369 (N_9369,N_9078,N_9188);
nor U9370 (N_9370,N_9151,N_9158);
or U9371 (N_9371,N_9215,N_9153);
or U9372 (N_9372,N_9185,N_9044);
and U9373 (N_9373,N_9049,N_9058);
and U9374 (N_9374,N_9067,N_9082);
nor U9375 (N_9375,N_9208,N_9244);
nand U9376 (N_9376,N_9197,N_9109);
nand U9377 (N_9377,N_9145,N_9036);
and U9378 (N_9378,N_9129,N_9176);
nor U9379 (N_9379,N_9043,N_9218);
nor U9380 (N_9380,N_9099,N_9100);
nand U9381 (N_9381,N_9241,N_9150);
nand U9382 (N_9382,N_9137,N_9171);
nand U9383 (N_9383,N_9212,N_9114);
nor U9384 (N_9384,N_9170,N_9142);
or U9385 (N_9385,N_9070,N_9213);
nand U9386 (N_9386,N_9166,N_9212);
and U9387 (N_9387,N_9172,N_9027);
nor U9388 (N_9388,N_9088,N_9076);
xor U9389 (N_9389,N_9106,N_9121);
nor U9390 (N_9390,N_9231,N_9211);
nor U9391 (N_9391,N_9030,N_9215);
or U9392 (N_9392,N_9124,N_9194);
nand U9393 (N_9393,N_9128,N_9039);
nand U9394 (N_9394,N_9219,N_9101);
xnor U9395 (N_9395,N_9178,N_9010);
and U9396 (N_9396,N_9195,N_9208);
and U9397 (N_9397,N_9068,N_9205);
nand U9398 (N_9398,N_9060,N_9171);
or U9399 (N_9399,N_9196,N_9192);
nor U9400 (N_9400,N_9211,N_9064);
nor U9401 (N_9401,N_9201,N_9215);
xnor U9402 (N_9402,N_9042,N_9024);
and U9403 (N_9403,N_9065,N_9047);
or U9404 (N_9404,N_9018,N_9170);
and U9405 (N_9405,N_9236,N_9059);
nand U9406 (N_9406,N_9021,N_9052);
or U9407 (N_9407,N_9222,N_9177);
and U9408 (N_9408,N_9040,N_9211);
or U9409 (N_9409,N_9215,N_9041);
and U9410 (N_9410,N_9151,N_9062);
and U9411 (N_9411,N_9036,N_9234);
nand U9412 (N_9412,N_9025,N_9180);
or U9413 (N_9413,N_9122,N_9028);
nor U9414 (N_9414,N_9064,N_9183);
or U9415 (N_9415,N_9170,N_9108);
nand U9416 (N_9416,N_9036,N_9200);
and U9417 (N_9417,N_9132,N_9162);
nor U9418 (N_9418,N_9037,N_9148);
xnor U9419 (N_9419,N_9086,N_9236);
nand U9420 (N_9420,N_9107,N_9044);
nor U9421 (N_9421,N_9126,N_9193);
nand U9422 (N_9422,N_9176,N_9182);
nand U9423 (N_9423,N_9187,N_9190);
nor U9424 (N_9424,N_9135,N_9204);
nor U9425 (N_9425,N_9181,N_9180);
or U9426 (N_9426,N_9232,N_9047);
nand U9427 (N_9427,N_9143,N_9056);
nand U9428 (N_9428,N_9078,N_9125);
or U9429 (N_9429,N_9009,N_9232);
nor U9430 (N_9430,N_9026,N_9206);
nor U9431 (N_9431,N_9126,N_9212);
nor U9432 (N_9432,N_9015,N_9184);
or U9433 (N_9433,N_9135,N_9210);
nor U9434 (N_9434,N_9029,N_9181);
and U9435 (N_9435,N_9034,N_9127);
nor U9436 (N_9436,N_9069,N_9198);
and U9437 (N_9437,N_9028,N_9216);
and U9438 (N_9438,N_9082,N_9208);
and U9439 (N_9439,N_9022,N_9036);
nand U9440 (N_9440,N_9011,N_9031);
and U9441 (N_9441,N_9166,N_9011);
or U9442 (N_9442,N_9110,N_9088);
nor U9443 (N_9443,N_9245,N_9191);
or U9444 (N_9444,N_9059,N_9004);
and U9445 (N_9445,N_9128,N_9022);
nor U9446 (N_9446,N_9133,N_9119);
and U9447 (N_9447,N_9169,N_9105);
and U9448 (N_9448,N_9007,N_9081);
nand U9449 (N_9449,N_9019,N_9011);
nor U9450 (N_9450,N_9021,N_9111);
and U9451 (N_9451,N_9070,N_9117);
and U9452 (N_9452,N_9034,N_9073);
and U9453 (N_9453,N_9033,N_9037);
nor U9454 (N_9454,N_9004,N_9186);
nand U9455 (N_9455,N_9245,N_9138);
nor U9456 (N_9456,N_9134,N_9000);
and U9457 (N_9457,N_9161,N_9073);
nand U9458 (N_9458,N_9184,N_9029);
and U9459 (N_9459,N_9240,N_9164);
or U9460 (N_9460,N_9114,N_9008);
and U9461 (N_9461,N_9193,N_9145);
and U9462 (N_9462,N_9146,N_9225);
and U9463 (N_9463,N_9128,N_9077);
and U9464 (N_9464,N_9226,N_9249);
xnor U9465 (N_9465,N_9123,N_9238);
nor U9466 (N_9466,N_9107,N_9230);
and U9467 (N_9467,N_9022,N_9192);
nand U9468 (N_9468,N_9167,N_9016);
nand U9469 (N_9469,N_9116,N_9121);
nand U9470 (N_9470,N_9033,N_9092);
and U9471 (N_9471,N_9042,N_9106);
nand U9472 (N_9472,N_9211,N_9038);
or U9473 (N_9473,N_9160,N_9115);
or U9474 (N_9474,N_9227,N_9019);
or U9475 (N_9475,N_9081,N_9018);
or U9476 (N_9476,N_9061,N_9082);
or U9477 (N_9477,N_9071,N_9031);
nor U9478 (N_9478,N_9064,N_9173);
or U9479 (N_9479,N_9043,N_9101);
nand U9480 (N_9480,N_9029,N_9240);
nor U9481 (N_9481,N_9134,N_9048);
nor U9482 (N_9482,N_9106,N_9117);
and U9483 (N_9483,N_9113,N_9243);
nor U9484 (N_9484,N_9181,N_9225);
nor U9485 (N_9485,N_9203,N_9066);
nand U9486 (N_9486,N_9004,N_9065);
nand U9487 (N_9487,N_9014,N_9020);
nand U9488 (N_9488,N_9022,N_9231);
nand U9489 (N_9489,N_9246,N_9100);
xnor U9490 (N_9490,N_9062,N_9076);
and U9491 (N_9491,N_9215,N_9187);
or U9492 (N_9492,N_9215,N_9019);
nand U9493 (N_9493,N_9067,N_9069);
nand U9494 (N_9494,N_9089,N_9239);
xnor U9495 (N_9495,N_9177,N_9009);
or U9496 (N_9496,N_9051,N_9209);
or U9497 (N_9497,N_9023,N_9011);
and U9498 (N_9498,N_9096,N_9118);
nor U9499 (N_9499,N_9206,N_9212);
or U9500 (N_9500,N_9286,N_9280);
and U9501 (N_9501,N_9465,N_9306);
nand U9502 (N_9502,N_9257,N_9284);
nor U9503 (N_9503,N_9303,N_9485);
xor U9504 (N_9504,N_9266,N_9481);
nand U9505 (N_9505,N_9335,N_9398);
nand U9506 (N_9506,N_9403,N_9352);
xnor U9507 (N_9507,N_9293,N_9262);
or U9508 (N_9508,N_9498,N_9448);
or U9509 (N_9509,N_9353,N_9288);
nand U9510 (N_9510,N_9349,N_9384);
or U9511 (N_9511,N_9310,N_9442);
nand U9512 (N_9512,N_9468,N_9460);
xnor U9513 (N_9513,N_9263,N_9368);
and U9514 (N_9514,N_9260,N_9490);
nor U9515 (N_9515,N_9371,N_9315);
xnor U9516 (N_9516,N_9324,N_9411);
nor U9517 (N_9517,N_9258,N_9289);
nand U9518 (N_9518,N_9499,N_9254);
and U9519 (N_9519,N_9430,N_9359);
nand U9520 (N_9520,N_9357,N_9304);
nand U9521 (N_9521,N_9432,N_9462);
nor U9522 (N_9522,N_9278,N_9358);
nor U9523 (N_9523,N_9261,N_9483);
or U9524 (N_9524,N_9424,N_9287);
nor U9525 (N_9525,N_9351,N_9362);
xor U9526 (N_9526,N_9441,N_9457);
and U9527 (N_9527,N_9376,N_9299);
xor U9528 (N_9528,N_9425,N_9433);
nand U9529 (N_9529,N_9305,N_9328);
nand U9530 (N_9530,N_9484,N_9283);
nand U9531 (N_9531,N_9395,N_9379);
xnor U9532 (N_9532,N_9334,N_9354);
and U9533 (N_9533,N_9370,N_9443);
or U9534 (N_9534,N_9418,N_9453);
xor U9535 (N_9535,N_9300,N_9330);
or U9536 (N_9536,N_9340,N_9292);
xnor U9537 (N_9537,N_9365,N_9265);
and U9538 (N_9538,N_9426,N_9273);
and U9539 (N_9539,N_9389,N_9329);
or U9540 (N_9540,N_9461,N_9367);
nand U9541 (N_9541,N_9440,N_9458);
and U9542 (N_9542,N_9489,N_9476);
nor U9543 (N_9543,N_9495,N_9291);
nand U9544 (N_9544,N_9355,N_9420);
nor U9545 (N_9545,N_9343,N_9270);
nand U9546 (N_9546,N_9323,N_9393);
nand U9547 (N_9547,N_9374,N_9346);
or U9548 (N_9548,N_9282,N_9382);
and U9549 (N_9549,N_9471,N_9437);
nor U9550 (N_9550,N_9251,N_9264);
or U9551 (N_9551,N_9332,N_9477);
and U9552 (N_9552,N_9439,N_9488);
or U9553 (N_9553,N_9322,N_9331);
xor U9554 (N_9554,N_9455,N_9327);
nor U9555 (N_9555,N_9445,N_9388);
nand U9556 (N_9556,N_9467,N_9491);
nand U9557 (N_9557,N_9405,N_9321);
xnor U9558 (N_9558,N_9482,N_9285);
and U9559 (N_9559,N_9383,N_9345);
nand U9560 (N_9560,N_9372,N_9377);
xor U9561 (N_9561,N_9313,N_9309);
and U9562 (N_9562,N_9302,N_9369);
and U9563 (N_9563,N_9279,N_9401);
nand U9564 (N_9564,N_9421,N_9456);
nand U9565 (N_9565,N_9336,N_9276);
and U9566 (N_9566,N_9429,N_9271);
nor U9567 (N_9567,N_9259,N_9480);
nor U9568 (N_9568,N_9378,N_9452);
nor U9569 (N_9569,N_9385,N_9318);
xor U9570 (N_9570,N_9496,N_9294);
and U9571 (N_9571,N_9423,N_9360);
or U9572 (N_9572,N_9339,N_9338);
nor U9573 (N_9573,N_9444,N_9447);
or U9574 (N_9574,N_9256,N_9399);
nand U9575 (N_9575,N_9394,N_9348);
and U9576 (N_9576,N_9414,N_9449);
and U9577 (N_9577,N_9347,N_9312);
or U9578 (N_9578,N_9373,N_9386);
nand U9579 (N_9579,N_9415,N_9446);
nor U9580 (N_9580,N_9400,N_9297);
nand U9581 (N_9581,N_9469,N_9341);
or U9582 (N_9582,N_9290,N_9275);
or U9583 (N_9583,N_9474,N_9326);
nor U9584 (N_9584,N_9366,N_9408);
and U9585 (N_9585,N_9434,N_9428);
nor U9586 (N_9586,N_9308,N_9487);
and U9587 (N_9587,N_9466,N_9409);
xor U9588 (N_9588,N_9407,N_9311);
and U9589 (N_9589,N_9295,N_9250);
xor U9590 (N_9590,N_9272,N_9274);
and U9591 (N_9591,N_9479,N_9463);
and U9592 (N_9592,N_9281,N_9412);
nand U9593 (N_9593,N_9301,N_9435);
or U9594 (N_9594,N_9494,N_9450);
nand U9595 (N_9595,N_9296,N_9298);
or U9596 (N_9596,N_9337,N_9497);
nand U9597 (N_9597,N_9473,N_9390);
or U9598 (N_9598,N_9397,N_9470);
or U9599 (N_9599,N_9472,N_9317);
or U9600 (N_9600,N_9320,N_9431);
or U9601 (N_9601,N_9252,N_9307);
nor U9602 (N_9602,N_9364,N_9387);
nor U9603 (N_9603,N_9380,N_9319);
nor U9604 (N_9604,N_9277,N_9255);
nor U9605 (N_9605,N_9396,N_9493);
or U9606 (N_9606,N_9269,N_9350);
nand U9607 (N_9607,N_9454,N_9459);
nand U9608 (N_9608,N_9402,N_9406);
nor U9609 (N_9609,N_9375,N_9486);
xor U9610 (N_9610,N_9267,N_9314);
or U9611 (N_9611,N_9422,N_9325);
and U9612 (N_9612,N_9316,N_9361);
nor U9613 (N_9613,N_9451,N_9404);
nand U9614 (N_9614,N_9253,N_9464);
and U9615 (N_9615,N_9410,N_9419);
and U9616 (N_9616,N_9492,N_9344);
xnor U9617 (N_9617,N_9478,N_9416);
nor U9618 (N_9618,N_9381,N_9392);
or U9619 (N_9619,N_9333,N_9475);
or U9620 (N_9620,N_9391,N_9268);
nor U9621 (N_9621,N_9436,N_9417);
and U9622 (N_9622,N_9427,N_9363);
nor U9623 (N_9623,N_9438,N_9413);
or U9624 (N_9624,N_9342,N_9356);
or U9625 (N_9625,N_9401,N_9271);
or U9626 (N_9626,N_9274,N_9376);
and U9627 (N_9627,N_9308,N_9392);
nor U9628 (N_9628,N_9443,N_9262);
xor U9629 (N_9629,N_9412,N_9316);
xnor U9630 (N_9630,N_9361,N_9452);
nand U9631 (N_9631,N_9492,N_9415);
xor U9632 (N_9632,N_9259,N_9363);
nand U9633 (N_9633,N_9286,N_9359);
or U9634 (N_9634,N_9466,N_9374);
nor U9635 (N_9635,N_9386,N_9369);
nor U9636 (N_9636,N_9275,N_9265);
nor U9637 (N_9637,N_9460,N_9384);
nand U9638 (N_9638,N_9455,N_9440);
or U9639 (N_9639,N_9462,N_9308);
nand U9640 (N_9640,N_9283,N_9443);
nor U9641 (N_9641,N_9250,N_9270);
and U9642 (N_9642,N_9300,N_9257);
and U9643 (N_9643,N_9319,N_9257);
nor U9644 (N_9644,N_9278,N_9275);
nand U9645 (N_9645,N_9452,N_9253);
nand U9646 (N_9646,N_9365,N_9350);
nor U9647 (N_9647,N_9251,N_9392);
or U9648 (N_9648,N_9449,N_9329);
nor U9649 (N_9649,N_9346,N_9281);
nor U9650 (N_9650,N_9496,N_9460);
or U9651 (N_9651,N_9314,N_9441);
and U9652 (N_9652,N_9479,N_9310);
and U9653 (N_9653,N_9406,N_9490);
nor U9654 (N_9654,N_9314,N_9482);
nand U9655 (N_9655,N_9295,N_9314);
and U9656 (N_9656,N_9459,N_9262);
or U9657 (N_9657,N_9495,N_9390);
nand U9658 (N_9658,N_9474,N_9387);
nor U9659 (N_9659,N_9272,N_9494);
and U9660 (N_9660,N_9280,N_9479);
nand U9661 (N_9661,N_9453,N_9301);
or U9662 (N_9662,N_9497,N_9408);
xnor U9663 (N_9663,N_9440,N_9359);
xnor U9664 (N_9664,N_9299,N_9475);
nand U9665 (N_9665,N_9402,N_9388);
nand U9666 (N_9666,N_9253,N_9348);
xor U9667 (N_9667,N_9273,N_9347);
nand U9668 (N_9668,N_9297,N_9293);
and U9669 (N_9669,N_9304,N_9380);
and U9670 (N_9670,N_9378,N_9375);
nand U9671 (N_9671,N_9319,N_9423);
nor U9672 (N_9672,N_9379,N_9321);
and U9673 (N_9673,N_9481,N_9269);
and U9674 (N_9674,N_9303,N_9338);
or U9675 (N_9675,N_9364,N_9423);
or U9676 (N_9676,N_9306,N_9420);
nor U9677 (N_9677,N_9309,N_9331);
and U9678 (N_9678,N_9451,N_9290);
nor U9679 (N_9679,N_9370,N_9360);
nand U9680 (N_9680,N_9453,N_9444);
or U9681 (N_9681,N_9498,N_9364);
xor U9682 (N_9682,N_9376,N_9472);
and U9683 (N_9683,N_9428,N_9251);
nand U9684 (N_9684,N_9274,N_9337);
or U9685 (N_9685,N_9313,N_9262);
nor U9686 (N_9686,N_9330,N_9338);
nand U9687 (N_9687,N_9250,N_9410);
and U9688 (N_9688,N_9419,N_9258);
or U9689 (N_9689,N_9428,N_9288);
and U9690 (N_9690,N_9262,N_9371);
nand U9691 (N_9691,N_9482,N_9421);
and U9692 (N_9692,N_9411,N_9251);
xor U9693 (N_9693,N_9470,N_9467);
nand U9694 (N_9694,N_9472,N_9347);
xnor U9695 (N_9695,N_9399,N_9308);
or U9696 (N_9696,N_9262,N_9372);
or U9697 (N_9697,N_9325,N_9324);
nor U9698 (N_9698,N_9250,N_9306);
nand U9699 (N_9699,N_9329,N_9412);
or U9700 (N_9700,N_9264,N_9375);
and U9701 (N_9701,N_9395,N_9478);
nand U9702 (N_9702,N_9294,N_9288);
nand U9703 (N_9703,N_9440,N_9385);
xor U9704 (N_9704,N_9479,N_9359);
nor U9705 (N_9705,N_9481,N_9251);
or U9706 (N_9706,N_9256,N_9483);
nand U9707 (N_9707,N_9253,N_9339);
nor U9708 (N_9708,N_9424,N_9312);
nand U9709 (N_9709,N_9478,N_9368);
or U9710 (N_9710,N_9342,N_9268);
and U9711 (N_9711,N_9289,N_9477);
and U9712 (N_9712,N_9324,N_9283);
or U9713 (N_9713,N_9349,N_9465);
and U9714 (N_9714,N_9493,N_9473);
nor U9715 (N_9715,N_9414,N_9454);
and U9716 (N_9716,N_9356,N_9371);
or U9717 (N_9717,N_9334,N_9481);
or U9718 (N_9718,N_9360,N_9309);
nand U9719 (N_9719,N_9483,N_9444);
or U9720 (N_9720,N_9271,N_9435);
xnor U9721 (N_9721,N_9286,N_9352);
or U9722 (N_9722,N_9357,N_9497);
nor U9723 (N_9723,N_9393,N_9289);
or U9724 (N_9724,N_9304,N_9331);
and U9725 (N_9725,N_9366,N_9362);
or U9726 (N_9726,N_9387,N_9349);
nor U9727 (N_9727,N_9392,N_9252);
nand U9728 (N_9728,N_9309,N_9398);
nand U9729 (N_9729,N_9422,N_9359);
nor U9730 (N_9730,N_9494,N_9373);
nand U9731 (N_9731,N_9336,N_9484);
nor U9732 (N_9732,N_9313,N_9419);
or U9733 (N_9733,N_9477,N_9417);
and U9734 (N_9734,N_9398,N_9419);
nor U9735 (N_9735,N_9329,N_9476);
xor U9736 (N_9736,N_9450,N_9329);
nor U9737 (N_9737,N_9430,N_9272);
nand U9738 (N_9738,N_9316,N_9375);
xnor U9739 (N_9739,N_9347,N_9345);
nor U9740 (N_9740,N_9404,N_9280);
or U9741 (N_9741,N_9486,N_9464);
nand U9742 (N_9742,N_9273,N_9442);
or U9743 (N_9743,N_9486,N_9439);
nor U9744 (N_9744,N_9420,N_9274);
nor U9745 (N_9745,N_9362,N_9382);
or U9746 (N_9746,N_9411,N_9332);
or U9747 (N_9747,N_9424,N_9326);
nor U9748 (N_9748,N_9395,N_9381);
nor U9749 (N_9749,N_9297,N_9443);
nand U9750 (N_9750,N_9687,N_9525);
nor U9751 (N_9751,N_9629,N_9705);
and U9752 (N_9752,N_9729,N_9524);
and U9753 (N_9753,N_9505,N_9554);
or U9754 (N_9754,N_9741,N_9711);
and U9755 (N_9755,N_9562,N_9551);
or U9756 (N_9756,N_9580,N_9529);
xnor U9757 (N_9757,N_9647,N_9544);
nor U9758 (N_9758,N_9506,N_9689);
and U9759 (N_9759,N_9575,N_9556);
nor U9760 (N_9760,N_9582,N_9628);
and U9761 (N_9761,N_9720,N_9590);
nand U9762 (N_9762,N_9514,N_9614);
nand U9763 (N_9763,N_9521,N_9737);
nor U9764 (N_9764,N_9644,N_9716);
nand U9765 (N_9765,N_9728,N_9583);
nand U9766 (N_9766,N_9567,N_9504);
and U9767 (N_9767,N_9704,N_9593);
nand U9768 (N_9768,N_9684,N_9730);
nand U9769 (N_9769,N_9513,N_9589);
or U9770 (N_9770,N_9641,N_9561);
and U9771 (N_9771,N_9616,N_9745);
nor U9772 (N_9772,N_9606,N_9527);
nor U9773 (N_9773,N_9530,N_9618);
nor U9774 (N_9774,N_9748,N_9631);
and U9775 (N_9775,N_9546,N_9611);
or U9776 (N_9776,N_9626,N_9653);
nor U9777 (N_9777,N_9643,N_9630);
and U9778 (N_9778,N_9648,N_9501);
nand U9779 (N_9779,N_9636,N_9671);
nand U9780 (N_9780,N_9665,N_9727);
nor U9781 (N_9781,N_9552,N_9654);
or U9782 (N_9782,N_9700,N_9591);
nand U9783 (N_9783,N_9739,N_9717);
or U9784 (N_9784,N_9634,N_9685);
nand U9785 (N_9785,N_9668,N_9651);
nor U9786 (N_9786,N_9608,N_9602);
or U9787 (N_9787,N_9541,N_9646);
nor U9788 (N_9788,N_9573,N_9662);
xor U9789 (N_9789,N_9579,N_9587);
nor U9790 (N_9790,N_9706,N_9528);
and U9791 (N_9791,N_9693,N_9678);
and U9792 (N_9792,N_9718,N_9661);
and U9793 (N_9793,N_9568,N_9663);
nor U9794 (N_9794,N_9533,N_9534);
nor U9795 (N_9795,N_9566,N_9586);
nand U9796 (N_9796,N_9564,N_9694);
nor U9797 (N_9797,N_9681,N_9613);
and U9798 (N_9798,N_9547,N_9701);
or U9799 (N_9799,N_9633,N_9682);
xnor U9800 (N_9800,N_9601,N_9597);
or U9801 (N_9801,N_9569,N_9742);
nand U9802 (N_9802,N_9531,N_9537);
nand U9803 (N_9803,N_9707,N_9596);
and U9804 (N_9804,N_9675,N_9683);
nand U9805 (N_9805,N_9598,N_9714);
or U9806 (N_9806,N_9540,N_9736);
and U9807 (N_9807,N_9518,N_9622);
nor U9808 (N_9808,N_9511,N_9725);
and U9809 (N_9809,N_9592,N_9545);
or U9810 (N_9810,N_9523,N_9732);
or U9811 (N_9811,N_9603,N_9627);
nor U9812 (N_9812,N_9617,N_9657);
and U9813 (N_9813,N_9659,N_9734);
xnor U9814 (N_9814,N_9522,N_9708);
or U9815 (N_9815,N_9609,N_9571);
xor U9816 (N_9816,N_9624,N_9666);
nand U9817 (N_9817,N_9667,N_9555);
and U9818 (N_9818,N_9600,N_9610);
and U9819 (N_9819,N_9558,N_9690);
and U9820 (N_9820,N_9519,N_9721);
and U9821 (N_9821,N_9508,N_9553);
nor U9822 (N_9822,N_9584,N_9686);
and U9823 (N_9823,N_9536,N_9563);
or U9824 (N_9824,N_9510,N_9565);
nor U9825 (N_9825,N_9503,N_9516);
xnor U9826 (N_9826,N_9543,N_9559);
xor U9827 (N_9827,N_9570,N_9672);
or U9828 (N_9828,N_9695,N_9703);
nor U9829 (N_9829,N_9673,N_9577);
or U9830 (N_9830,N_9743,N_9604);
nor U9831 (N_9831,N_9676,N_9747);
xor U9832 (N_9832,N_9637,N_9697);
nor U9833 (N_9833,N_9652,N_9702);
or U9834 (N_9834,N_9699,N_9615);
nand U9835 (N_9835,N_9632,N_9680);
and U9836 (N_9836,N_9621,N_9625);
or U9837 (N_9837,N_9639,N_9538);
or U9838 (N_9838,N_9594,N_9549);
nand U9839 (N_9839,N_9535,N_9712);
or U9840 (N_9840,N_9655,N_9640);
nand U9841 (N_9841,N_9500,N_9688);
xnor U9842 (N_9842,N_9515,N_9724);
nand U9843 (N_9843,N_9557,N_9595);
nand U9844 (N_9844,N_9581,N_9746);
or U9845 (N_9845,N_9526,N_9517);
nand U9846 (N_9846,N_9649,N_9635);
nand U9847 (N_9847,N_9638,N_9660);
or U9848 (N_9848,N_9715,N_9520);
nor U9849 (N_9849,N_9670,N_9674);
xnor U9850 (N_9850,N_9542,N_9619);
nand U9851 (N_9851,N_9669,N_9578);
nor U9852 (N_9852,N_9709,N_9623);
nor U9853 (N_9853,N_9698,N_9572);
nor U9854 (N_9854,N_9512,N_9588);
nand U9855 (N_9855,N_9656,N_9607);
and U9856 (N_9856,N_9550,N_9749);
nor U9857 (N_9857,N_9507,N_9560);
nor U9858 (N_9858,N_9664,N_9509);
nand U9859 (N_9859,N_9599,N_9722);
and U9860 (N_9860,N_9539,N_9658);
nand U9861 (N_9861,N_9642,N_9696);
or U9862 (N_9862,N_9692,N_9723);
or U9863 (N_9863,N_9719,N_9744);
nand U9864 (N_9864,N_9735,N_9620);
nand U9865 (N_9865,N_9645,N_9733);
and U9866 (N_9866,N_9585,N_9731);
or U9867 (N_9867,N_9605,N_9679);
and U9868 (N_9868,N_9726,N_9740);
or U9869 (N_9869,N_9691,N_9650);
nand U9870 (N_9870,N_9677,N_9612);
nor U9871 (N_9871,N_9574,N_9576);
or U9872 (N_9872,N_9710,N_9502);
nand U9873 (N_9873,N_9713,N_9532);
and U9874 (N_9874,N_9738,N_9548);
nor U9875 (N_9875,N_9547,N_9744);
nor U9876 (N_9876,N_9577,N_9550);
or U9877 (N_9877,N_9545,N_9670);
and U9878 (N_9878,N_9656,N_9625);
and U9879 (N_9879,N_9573,N_9531);
or U9880 (N_9880,N_9616,N_9621);
nand U9881 (N_9881,N_9537,N_9587);
or U9882 (N_9882,N_9572,N_9647);
nor U9883 (N_9883,N_9589,N_9632);
and U9884 (N_9884,N_9737,N_9528);
nand U9885 (N_9885,N_9676,N_9708);
or U9886 (N_9886,N_9618,N_9545);
xor U9887 (N_9887,N_9699,N_9501);
or U9888 (N_9888,N_9662,N_9543);
nand U9889 (N_9889,N_9738,N_9702);
and U9890 (N_9890,N_9635,N_9505);
or U9891 (N_9891,N_9633,N_9513);
xnor U9892 (N_9892,N_9601,N_9586);
and U9893 (N_9893,N_9569,N_9725);
nor U9894 (N_9894,N_9648,N_9586);
nor U9895 (N_9895,N_9500,N_9691);
nor U9896 (N_9896,N_9704,N_9725);
nor U9897 (N_9897,N_9707,N_9558);
and U9898 (N_9898,N_9607,N_9599);
and U9899 (N_9899,N_9667,N_9623);
nand U9900 (N_9900,N_9572,N_9731);
xor U9901 (N_9901,N_9559,N_9578);
xor U9902 (N_9902,N_9687,N_9664);
or U9903 (N_9903,N_9681,N_9606);
nor U9904 (N_9904,N_9547,N_9585);
or U9905 (N_9905,N_9722,N_9522);
nand U9906 (N_9906,N_9592,N_9604);
or U9907 (N_9907,N_9684,N_9632);
nor U9908 (N_9908,N_9676,N_9525);
xor U9909 (N_9909,N_9588,N_9649);
nand U9910 (N_9910,N_9520,N_9688);
nor U9911 (N_9911,N_9694,N_9620);
nor U9912 (N_9912,N_9550,N_9543);
xor U9913 (N_9913,N_9566,N_9543);
xnor U9914 (N_9914,N_9636,N_9587);
nand U9915 (N_9915,N_9565,N_9623);
or U9916 (N_9916,N_9600,N_9624);
nor U9917 (N_9917,N_9701,N_9714);
and U9918 (N_9918,N_9602,N_9638);
nor U9919 (N_9919,N_9586,N_9541);
nor U9920 (N_9920,N_9529,N_9609);
and U9921 (N_9921,N_9606,N_9747);
xnor U9922 (N_9922,N_9713,N_9624);
and U9923 (N_9923,N_9665,N_9527);
nand U9924 (N_9924,N_9554,N_9672);
nor U9925 (N_9925,N_9627,N_9578);
nand U9926 (N_9926,N_9651,N_9679);
nand U9927 (N_9927,N_9737,N_9698);
or U9928 (N_9928,N_9590,N_9602);
nand U9929 (N_9929,N_9589,N_9716);
or U9930 (N_9930,N_9744,N_9738);
nor U9931 (N_9931,N_9582,N_9679);
or U9932 (N_9932,N_9567,N_9609);
nor U9933 (N_9933,N_9578,N_9672);
xnor U9934 (N_9934,N_9713,N_9552);
nor U9935 (N_9935,N_9680,N_9606);
xnor U9936 (N_9936,N_9743,N_9628);
nor U9937 (N_9937,N_9585,N_9509);
nand U9938 (N_9938,N_9636,N_9661);
nor U9939 (N_9939,N_9718,N_9642);
and U9940 (N_9940,N_9575,N_9516);
nor U9941 (N_9941,N_9628,N_9671);
or U9942 (N_9942,N_9693,N_9616);
and U9943 (N_9943,N_9520,N_9653);
xor U9944 (N_9944,N_9583,N_9642);
nor U9945 (N_9945,N_9547,N_9641);
nor U9946 (N_9946,N_9631,N_9522);
nand U9947 (N_9947,N_9567,N_9562);
nor U9948 (N_9948,N_9572,N_9686);
nor U9949 (N_9949,N_9662,N_9609);
nand U9950 (N_9950,N_9657,N_9521);
and U9951 (N_9951,N_9701,N_9619);
and U9952 (N_9952,N_9738,N_9534);
and U9953 (N_9953,N_9714,N_9596);
and U9954 (N_9954,N_9600,N_9644);
or U9955 (N_9955,N_9623,N_9713);
or U9956 (N_9956,N_9713,N_9569);
nand U9957 (N_9957,N_9705,N_9553);
nor U9958 (N_9958,N_9672,N_9594);
xor U9959 (N_9959,N_9688,N_9668);
nand U9960 (N_9960,N_9668,N_9549);
nor U9961 (N_9961,N_9690,N_9623);
or U9962 (N_9962,N_9716,N_9739);
nand U9963 (N_9963,N_9525,N_9683);
xor U9964 (N_9964,N_9592,N_9555);
or U9965 (N_9965,N_9685,N_9642);
and U9966 (N_9966,N_9511,N_9652);
and U9967 (N_9967,N_9729,N_9669);
nand U9968 (N_9968,N_9713,N_9593);
nand U9969 (N_9969,N_9713,N_9606);
and U9970 (N_9970,N_9732,N_9702);
xor U9971 (N_9971,N_9745,N_9645);
nand U9972 (N_9972,N_9581,N_9640);
and U9973 (N_9973,N_9588,N_9582);
or U9974 (N_9974,N_9542,N_9686);
or U9975 (N_9975,N_9698,N_9678);
and U9976 (N_9976,N_9551,N_9738);
and U9977 (N_9977,N_9533,N_9505);
or U9978 (N_9978,N_9566,N_9520);
and U9979 (N_9979,N_9648,N_9678);
or U9980 (N_9980,N_9658,N_9506);
or U9981 (N_9981,N_9660,N_9698);
xnor U9982 (N_9982,N_9568,N_9500);
nor U9983 (N_9983,N_9548,N_9706);
or U9984 (N_9984,N_9659,N_9518);
nor U9985 (N_9985,N_9743,N_9569);
and U9986 (N_9986,N_9691,N_9622);
or U9987 (N_9987,N_9615,N_9548);
and U9988 (N_9988,N_9723,N_9719);
nand U9989 (N_9989,N_9533,N_9594);
and U9990 (N_9990,N_9636,N_9735);
nor U9991 (N_9991,N_9702,N_9685);
or U9992 (N_9992,N_9657,N_9615);
or U9993 (N_9993,N_9567,N_9638);
or U9994 (N_9994,N_9639,N_9535);
and U9995 (N_9995,N_9568,N_9592);
and U9996 (N_9996,N_9732,N_9637);
nor U9997 (N_9997,N_9749,N_9675);
nand U9998 (N_9998,N_9549,N_9681);
nor U9999 (N_9999,N_9714,N_9631);
nor U10000 (N_10000,N_9886,N_9804);
and U10001 (N_10001,N_9761,N_9856);
nand U10002 (N_10002,N_9842,N_9829);
nor U10003 (N_10003,N_9758,N_9961);
and U10004 (N_10004,N_9750,N_9935);
nand U10005 (N_10005,N_9902,N_9756);
nor U10006 (N_10006,N_9808,N_9910);
or U10007 (N_10007,N_9795,N_9903);
or U10008 (N_10008,N_9970,N_9922);
and U10009 (N_10009,N_9850,N_9861);
nand U10010 (N_10010,N_9784,N_9981);
nand U10011 (N_10011,N_9941,N_9852);
nand U10012 (N_10012,N_9928,N_9917);
xor U10013 (N_10013,N_9796,N_9989);
nor U10014 (N_10014,N_9958,N_9759);
and U10015 (N_10015,N_9813,N_9789);
nor U10016 (N_10016,N_9879,N_9968);
xnor U10017 (N_10017,N_9919,N_9840);
nor U10018 (N_10018,N_9899,N_9959);
xor U10019 (N_10019,N_9755,N_9925);
or U10020 (N_10020,N_9931,N_9839);
xnor U10021 (N_10021,N_9984,N_9848);
nand U10022 (N_10022,N_9912,N_9977);
and U10023 (N_10023,N_9907,N_9763);
or U10024 (N_10024,N_9983,N_9859);
or U10025 (N_10025,N_9832,N_9851);
or U10026 (N_10026,N_9869,N_9971);
nand U10027 (N_10027,N_9947,N_9969);
nand U10028 (N_10028,N_9817,N_9858);
or U10029 (N_10029,N_9849,N_9788);
and U10030 (N_10030,N_9943,N_9976);
and U10031 (N_10031,N_9798,N_9887);
and U10032 (N_10032,N_9927,N_9866);
and U10033 (N_10033,N_9883,N_9787);
nand U10034 (N_10034,N_9982,N_9993);
and U10035 (N_10035,N_9894,N_9831);
nor U10036 (N_10036,N_9884,N_9998);
nor U10037 (N_10037,N_9822,N_9945);
and U10038 (N_10038,N_9791,N_9882);
and U10039 (N_10039,N_9771,N_9891);
and U10040 (N_10040,N_9860,N_9853);
nand U10041 (N_10041,N_9888,N_9876);
nor U10042 (N_10042,N_9870,N_9948);
or U10043 (N_10043,N_9929,N_9769);
and U10044 (N_10044,N_9833,N_9871);
and U10045 (N_10045,N_9834,N_9914);
and U10046 (N_10046,N_9942,N_9785);
nand U10047 (N_10047,N_9868,N_9986);
nor U10048 (N_10048,N_9938,N_9807);
nand U10049 (N_10049,N_9826,N_9994);
or U10050 (N_10050,N_9889,N_9827);
nor U10051 (N_10051,N_9939,N_9843);
or U10052 (N_10052,N_9892,N_9898);
nor U10053 (N_10053,N_9965,N_9957);
or U10054 (N_10054,N_9885,N_9801);
nor U10055 (N_10055,N_9897,N_9824);
nand U10056 (N_10056,N_9999,N_9814);
nand U10057 (N_10057,N_9823,N_9954);
nand U10058 (N_10058,N_9995,N_9776);
or U10059 (N_10059,N_9778,N_9974);
nor U10060 (N_10060,N_9864,N_9915);
xor U10061 (N_10061,N_9905,N_9786);
xnor U10062 (N_10062,N_9760,N_9881);
nor U10063 (N_10063,N_9920,N_9997);
and U10064 (N_10064,N_9867,N_9781);
nor U10065 (N_10065,N_9956,N_9790);
nand U10066 (N_10066,N_9990,N_9835);
or U10067 (N_10067,N_9792,N_9775);
nand U10068 (N_10068,N_9799,N_9777);
nand U10069 (N_10069,N_9854,N_9819);
nand U10070 (N_10070,N_9923,N_9766);
nand U10071 (N_10071,N_9900,N_9855);
and U10072 (N_10072,N_9937,N_9762);
xnor U10073 (N_10073,N_9909,N_9874);
or U10074 (N_10074,N_9930,N_9774);
and U10075 (N_10075,N_9955,N_9991);
nor U10076 (N_10076,N_9825,N_9967);
or U10077 (N_10077,N_9809,N_9895);
nor U10078 (N_10078,N_9890,N_9896);
nand U10079 (N_10079,N_9985,N_9770);
or U10080 (N_10080,N_9802,N_9810);
nor U10081 (N_10081,N_9966,N_9793);
xor U10082 (N_10082,N_9812,N_9773);
nand U10083 (N_10083,N_9805,N_9988);
nand U10084 (N_10084,N_9960,N_9800);
or U10085 (N_10085,N_9863,N_9949);
and U10086 (N_10086,N_9913,N_9973);
or U10087 (N_10087,N_9828,N_9846);
and U10088 (N_10088,N_9797,N_9873);
nor U10089 (N_10089,N_9944,N_9904);
nand U10090 (N_10090,N_9901,N_9821);
or U10091 (N_10091,N_9975,N_9768);
and U10092 (N_10092,N_9753,N_9767);
or U10093 (N_10093,N_9962,N_9934);
nor U10094 (N_10094,N_9830,N_9765);
and U10095 (N_10095,N_9847,N_9950);
nor U10096 (N_10096,N_9872,N_9951);
or U10097 (N_10097,N_9811,N_9972);
nor U10098 (N_10098,N_9880,N_9979);
xor U10099 (N_10099,N_9816,N_9924);
xor U10100 (N_10100,N_9841,N_9836);
or U10101 (N_10101,N_9980,N_9857);
xor U10102 (N_10102,N_9963,N_9940);
nand U10103 (N_10103,N_9751,N_9911);
or U10104 (N_10104,N_9877,N_9878);
nor U10105 (N_10105,N_9921,N_9779);
xnor U10106 (N_10106,N_9782,N_9996);
or U10107 (N_10107,N_9908,N_9752);
nand U10108 (N_10108,N_9865,N_9918);
and U10109 (N_10109,N_9875,N_9806);
nand U10110 (N_10110,N_9926,N_9987);
nand U10111 (N_10111,N_9862,N_9794);
xor U10112 (N_10112,N_9772,N_9754);
xnor U10113 (N_10113,N_9818,N_9845);
and U10114 (N_10114,N_9906,N_9764);
nand U10115 (N_10115,N_9803,N_9783);
nor U10116 (N_10116,N_9844,N_9932);
nor U10117 (N_10117,N_9992,N_9933);
and U10118 (N_10118,N_9757,N_9964);
or U10119 (N_10119,N_9838,N_9936);
and U10120 (N_10120,N_9916,N_9952);
nand U10121 (N_10121,N_9815,N_9953);
or U10122 (N_10122,N_9946,N_9837);
nand U10123 (N_10123,N_9893,N_9978);
nand U10124 (N_10124,N_9780,N_9820);
or U10125 (N_10125,N_9976,N_9789);
and U10126 (N_10126,N_9842,N_9990);
nand U10127 (N_10127,N_9837,N_9840);
and U10128 (N_10128,N_9946,N_9874);
or U10129 (N_10129,N_9801,N_9889);
nand U10130 (N_10130,N_9756,N_9858);
or U10131 (N_10131,N_9801,N_9928);
and U10132 (N_10132,N_9864,N_9844);
and U10133 (N_10133,N_9814,N_9780);
xnor U10134 (N_10134,N_9911,N_9933);
nand U10135 (N_10135,N_9876,N_9765);
nand U10136 (N_10136,N_9931,N_9767);
nor U10137 (N_10137,N_9826,N_9910);
or U10138 (N_10138,N_9771,N_9791);
nand U10139 (N_10139,N_9844,N_9889);
or U10140 (N_10140,N_9810,N_9768);
xnor U10141 (N_10141,N_9846,N_9781);
or U10142 (N_10142,N_9918,N_9881);
or U10143 (N_10143,N_9765,N_9882);
or U10144 (N_10144,N_9864,N_9753);
and U10145 (N_10145,N_9831,N_9764);
nand U10146 (N_10146,N_9988,N_9750);
xor U10147 (N_10147,N_9984,N_9874);
nand U10148 (N_10148,N_9940,N_9924);
xor U10149 (N_10149,N_9961,N_9969);
nor U10150 (N_10150,N_9910,N_9889);
or U10151 (N_10151,N_9835,N_9874);
and U10152 (N_10152,N_9917,N_9987);
or U10153 (N_10153,N_9889,N_9979);
nor U10154 (N_10154,N_9773,N_9837);
nand U10155 (N_10155,N_9934,N_9904);
and U10156 (N_10156,N_9911,N_9946);
nor U10157 (N_10157,N_9912,N_9783);
or U10158 (N_10158,N_9876,N_9819);
or U10159 (N_10159,N_9790,N_9863);
nor U10160 (N_10160,N_9809,N_9829);
or U10161 (N_10161,N_9906,N_9889);
nor U10162 (N_10162,N_9810,N_9839);
nand U10163 (N_10163,N_9965,N_9950);
nand U10164 (N_10164,N_9959,N_9982);
xnor U10165 (N_10165,N_9807,N_9850);
nor U10166 (N_10166,N_9913,N_9809);
nand U10167 (N_10167,N_9815,N_9907);
nor U10168 (N_10168,N_9812,N_9976);
or U10169 (N_10169,N_9924,N_9923);
nand U10170 (N_10170,N_9779,N_9847);
nand U10171 (N_10171,N_9791,N_9901);
or U10172 (N_10172,N_9961,N_9947);
or U10173 (N_10173,N_9820,N_9879);
nor U10174 (N_10174,N_9894,N_9798);
or U10175 (N_10175,N_9826,N_9868);
or U10176 (N_10176,N_9889,N_9770);
and U10177 (N_10177,N_9832,N_9835);
and U10178 (N_10178,N_9898,N_9864);
and U10179 (N_10179,N_9755,N_9840);
nor U10180 (N_10180,N_9812,N_9768);
or U10181 (N_10181,N_9851,N_9836);
nand U10182 (N_10182,N_9993,N_9795);
nand U10183 (N_10183,N_9847,N_9966);
and U10184 (N_10184,N_9859,N_9999);
and U10185 (N_10185,N_9849,N_9878);
or U10186 (N_10186,N_9917,N_9910);
nor U10187 (N_10187,N_9971,N_9836);
nor U10188 (N_10188,N_9978,N_9779);
nor U10189 (N_10189,N_9827,N_9818);
and U10190 (N_10190,N_9754,N_9854);
and U10191 (N_10191,N_9937,N_9976);
nor U10192 (N_10192,N_9805,N_9877);
nand U10193 (N_10193,N_9906,N_9845);
and U10194 (N_10194,N_9950,N_9921);
nor U10195 (N_10195,N_9812,N_9791);
nor U10196 (N_10196,N_9911,N_9943);
nor U10197 (N_10197,N_9788,N_9848);
xor U10198 (N_10198,N_9761,N_9774);
nand U10199 (N_10199,N_9952,N_9860);
xnor U10200 (N_10200,N_9937,N_9897);
and U10201 (N_10201,N_9849,N_9781);
nor U10202 (N_10202,N_9775,N_9757);
and U10203 (N_10203,N_9830,N_9769);
and U10204 (N_10204,N_9826,N_9955);
and U10205 (N_10205,N_9820,N_9943);
or U10206 (N_10206,N_9816,N_9889);
xor U10207 (N_10207,N_9908,N_9949);
or U10208 (N_10208,N_9758,N_9805);
or U10209 (N_10209,N_9853,N_9770);
and U10210 (N_10210,N_9841,N_9837);
nor U10211 (N_10211,N_9813,N_9804);
and U10212 (N_10212,N_9923,N_9778);
and U10213 (N_10213,N_9986,N_9772);
nor U10214 (N_10214,N_9974,N_9878);
and U10215 (N_10215,N_9792,N_9765);
and U10216 (N_10216,N_9826,N_9924);
nor U10217 (N_10217,N_9784,N_9980);
nor U10218 (N_10218,N_9903,N_9927);
and U10219 (N_10219,N_9987,N_9923);
xnor U10220 (N_10220,N_9907,N_9900);
nor U10221 (N_10221,N_9801,N_9905);
and U10222 (N_10222,N_9864,N_9822);
nand U10223 (N_10223,N_9986,N_9800);
xnor U10224 (N_10224,N_9938,N_9985);
and U10225 (N_10225,N_9872,N_9993);
and U10226 (N_10226,N_9807,N_9856);
or U10227 (N_10227,N_9796,N_9883);
and U10228 (N_10228,N_9926,N_9918);
or U10229 (N_10229,N_9989,N_9888);
nand U10230 (N_10230,N_9961,N_9750);
nand U10231 (N_10231,N_9763,N_9872);
nor U10232 (N_10232,N_9931,N_9920);
nor U10233 (N_10233,N_9857,N_9815);
or U10234 (N_10234,N_9949,N_9979);
xnor U10235 (N_10235,N_9876,N_9904);
nor U10236 (N_10236,N_9777,N_9948);
and U10237 (N_10237,N_9803,N_9844);
or U10238 (N_10238,N_9786,N_9925);
or U10239 (N_10239,N_9777,N_9802);
nand U10240 (N_10240,N_9786,N_9859);
nand U10241 (N_10241,N_9768,N_9967);
nand U10242 (N_10242,N_9920,N_9967);
or U10243 (N_10243,N_9906,N_9847);
xnor U10244 (N_10244,N_9994,N_9937);
or U10245 (N_10245,N_9873,N_9790);
nor U10246 (N_10246,N_9926,N_9961);
or U10247 (N_10247,N_9878,N_9770);
nand U10248 (N_10248,N_9938,N_9843);
or U10249 (N_10249,N_9925,N_9828);
xnor U10250 (N_10250,N_10029,N_10035);
and U10251 (N_10251,N_10120,N_10146);
nand U10252 (N_10252,N_10058,N_10000);
or U10253 (N_10253,N_10102,N_10134);
and U10254 (N_10254,N_10076,N_10160);
or U10255 (N_10255,N_10182,N_10159);
xor U10256 (N_10256,N_10226,N_10130);
or U10257 (N_10257,N_10087,N_10141);
or U10258 (N_10258,N_10106,N_10037);
nand U10259 (N_10259,N_10062,N_10121);
and U10260 (N_10260,N_10154,N_10158);
nor U10261 (N_10261,N_10186,N_10008);
nand U10262 (N_10262,N_10225,N_10021);
or U10263 (N_10263,N_10017,N_10208);
or U10264 (N_10264,N_10211,N_10227);
nand U10265 (N_10265,N_10192,N_10103);
and U10266 (N_10266,N_10046,N_10041);
nor U10267 (N_10267,N_10082,N_10170);
nand U10268 (N_10268,N_10236,N_10163);
or U10269 (N_10269,N_10197,N_10094);
and U10270 (N_10270,N_10171,N_10059);
and U10271 (N_10271,N_10177,N_10230);
or U10272 (N_10272,N_10195,N_10239);
xor U10273 (N_10273,N_10105,N_10080);
and U10274 (N_10274,N_10173,N_10248);
and U10275 (N_10275,N_10193,N_10093);
nor U10276 (N_10276,N_10201,N_10150);
nor U10277 (N_10277,N_10142,N_10061);
nor U10278 (N_10278,N_10075,N_10157);
nand U10279 (N_10279,N_10242,N_10005);
nand U10280 (N_10280,N_10219,N_10016);
xor U10281 (N_10281,N_10210,N_10131);
nand U10282 (N_10282,N_10036,N_10033);
or U10283 (N_10283,N_10156,N_10113);
and U10284 (N_10284,N_10012,N_10085);
nand U10285 (N_10285,N_10006,N_10188);
nor U10286 (N_10286,N_10065,N_10235);
nor U10287 (N_10287,N_10100,N_10009);
and U10288 (N_10288,N_10233,N_10084);
nor U10289 (N_10289,N_10051,N_10136);
nor U10290 (N_10290,N_10191,N_10181);
nor U10291 (N_10291,N_10234,N_10054);
xor U10292 (N_10292,N_10111,N_10176);
nor U10293 (N_10293,N_10206,N_10042);
nand U10294 (N_10294,N_10125,N_10229);
xnor U10295 (N_10295,N_10089,N_10144);
and U10296 (N_10296,N_10222,N_10180);
and U10297 (N_10297,N_10028,N_10138);
nand U10298 (N_10298,N_10224,N_10243);
and U10299 (N_10299,N_10043,N_10143);
nor U10300 (N_10300,N_10174,N_10056);
or U10301 (N_10301,N_10246,N_10088);
nand U10302 (N_10302,N_10018,N_10090);
and U10303 (N_10303,N_10072,N_10161);
nor U10304 (N_10304,N_10108,N_10169);
or U10305 (N_10305,N_10139,N_10026);
or U10306 (N_10306,N_10027,N_10055);
and U10307 (N_10307,N_10073,N_10123);
and U10308 (N_10308,N_10133,N_10116);
or U10309 (N_10309,N_10014,N_10019);
and U10310 (N_10310,N_10038,N_10162);
and U10311 (N_10311,N_10097,N_10119);
nand U10312 (N_10312,N_10147,N_10221);
and U10313 (N_10313,N_10137,N_10241);
nand U10314 (N_10314,N_10011,N_10124);
and U10315 (N_10315,N_10066,N_10127);
nor U10316 (N_10316,N_10081,N_10175);
nand U10317 (N_10317,N_10183,N_10207);
nor U10318 (N_10318,N_10115,N_10140);
nor U10319 (N_10319,N_10245,N_10099);
and U10320 (N_10320,N_10194,N_10047);
nand U10321 (N_10321,N_10128,N_10053);
nor U10322 (N_10322,N_10003,N_10214);
nor U10323 (N_10323,N_10020,N_10034);
nand U10324 (N_10324,N_10096,N_10117);
xnor U10325 (N_10325,N_10045,N_10198);
and U10326 (N_10326,N_10165,N_10068);
nand U10327 (N_10327,N_10199,N_10238);
nor U10328 (N_10328,N_10232,N_10240);
nor U10329 (N_10329,N_10228,N_10007);
or U10330 (N_10330,N_10215,N_10004);
nand U10331 (N_10331,N_10074,N_10220);
xnor U10332 (N_10332,N_10217,N_10212);
or U10333 (N_10333,N_10178,N_10050);
and U10334 (N_10334,N_10164,N_10083);
or U10335 (N_10335,N_10010,N_10209);
nor U10336 (N_10336,N_10118,N_10092);
and U10337 (N_10337,N_10031,N_10101);
nand U10338 (N_10338,N_10184,N_10132);
and U10339 (N_10339,N_10040,N_10032);
and U10340 (N_10340,N_10247,N_10002);
and U10341 (N_10341,N_10064,N_10189);
nor U10342 (N_10342,N_10196,N_10187);
or U10343 (N_10343,N_10024,N_10071);
nor U10344 (N_10344,N_10129,N_10145);
xor U10345 (N_10345,N_10200,N_10044);
or U10346 (N_10346,N_10152,N_10172);
xnor U10347 (N_10347,N_10237,N_10069);
nor U10348 (N_10348,N_10104,N_10025);
or U10349 (N_10349,N_10190,N_10166);
nand U10350 (N_10350,N_10052,N_10110);
nand U10351 (N_10351,N_10112,N_10135);
or U10352 (N_10352,N_10167,N_10231);
and U10353 (N_10353,N_10223,N_10023);
or U10354 (N_10354,N_10013,N_10079);
nand U10355 (N_10355,N_10030,N_10149);
or U10356 (N_10356,N_10151,N_10148);
or U10357 (N_10357,N_10107,N_10001);
and U10358 (N_10358,N_10179,N_10095);
and U10359 (N_10359,N_10168,N_10039);
xor U10360 (N_10360,N_10202,N_10213);
nor U10361 (N_10361,N_10249,N_10063);
nor U10362 (N_10362,N_10216,N_10060);
or U10363 (N_10363,N_10205,N_10122);
nor U10364 (N_10364,N_10091,N_10098);
or U10365 (N_10365,N_10022,N_10204);
and U10366 (N_10366,N_10086,N_10153);
xnor U10367 (N_10367,N_10126,N_10077);
nor U10368 (N_10368,N_10078,N_10067);
or U10369 (N_10369,N_10155,N_10070);
nand U10370 (N_10370,N_10057,N_10049);
nor U10371 (N_10371,N_10218,N_10244);
and U10372 (N_10372,N_10114,N_10015);
xnor U10373 (N_10373,N_10185,N_10203);
and U10374 (N_10374,N_10048,N_10109);
nor U10375 (N_10375,N_10035,N_10219);
nand U10376 (N_10376,N_10097,N_10240);
or U10377 (N_10377,N_10204,N_10088);
nor U10378 (N_10378,N_10159,N_10106);
nor U10379 (N_10379,N_10192,N_10173);
nor U10380 (N_10380,N_10109,N_10055);
or U10381 (N_10381,N_10149,N_10231);
nand U10382 (N_10382,N_10224,N_10220);
nand U10383 (N_10383,N_10201,N_10125);
or U10384 (N_10384,N_10162,N_10068);
and U10385 (N_10385,N_10140,N_10074);
or U10386 (N_10386,N_10070,N_10103);
nand U10387 (N_10387,N_10124,N_10024);
nand U10388 (N_10388,N_10150,N_10236);
xor U10389 (N_10389,N_10236,N_10247);
and U10390 (N_10390,N_10038,N_10195);
or U10391 (N_10391,N_10015,N_10021);
and U10392 (N_10392,N_10091,N_10245);
nor U10393 (N_10393,N_10194,N_10108);
or U10394 (N_10394,N_10122,N_10160);
nor U10395 (N_10395,N_10060,N_10215);
nand U10396 (N_10396,N_10008,N_10169);
and U10397 (N_10397,N_10158,N_10014);
nor U10398 (N_10398,N_10207,N_10199);
xnor U10399 (N_10399,N_10112,N_10039);
and U10400 (N_10400,N_10090,N_10094);
xnor U10401 (N_10401,N_10190,N_10136);
nand U10402 (N_10402,N_10220,N_10046);
nand U10403 (N_10403,N_10080,N_10127);
and U10404 (N_10404,N_10189,N_10061);
or U10405 (N_10405,N_10160,N_10001);
xnor U10406 (N_10406,N_10063,N_10226);
or U10407 (N_10407,N_10097,N_10089);
and U10408 (N_10408,N_10220,N_10073);
or U10409 (N_10409,N_10080,N_10021);
nor U10410 (N_10410,N_10060,N_10006);
and U10411 (N_10411,N_10134,N_10200);
xnor U10412 (N_10412,N_10220,N_10059);
nor U10413 (N_10413,N_10080,N_10161);
nor U10414 (N_10414,N_10053,N_10234);
nor U10415 (N_10415,N_10126,N_10063);
nor U10416 (N_10416,N_10197,N_10190);
nand U10417 (N_10417,N_10172,N_10010);
nor U10418 (N_10418,N_10013,N_10003);
and U10419 (N_10419,N_10197,N_10040);
or U10420 (N_10420,N_10013,N_10098);
or U10421 (N_10421,N_10056,N_10084);
nor U10422 (N_10422,N_10093,N_10108);
or U10423 (N_10423,N_10103,N_10001);
and U10424 (N_10424,N_10166,N_10235);
nand U10425 (N_10425,N_10070,N_10116);
nand U10426 (N_10426,N_10031,N_10069);
nor U10427 (N_10427,N_10034,N_10170);
and U10428 (N_10428,N_10230,N_10065);
nor U10429 (N_10429,N_10195,N_10053);
xnor U10430 (N_10430,N_10009,N_10030);
or U10431 (N_10431,N_10225,N_10007);
nor U10432 (N_10432,N_10163,N_10143);
nand U10433 (N_10433,N_10146,N_10154);
nor U10434 (N_10434,N_10171,N_10185);
nand U10435 (N_10435,N_10160,N_10229);
nor U10436 (N_10436,N_10213,N_10117);
or U10437 (N_10437,N_10174,N_10239);
nand U10438 (N_10438,N_10099,N_10098);
or U10439 (N_10439,N_10089,N_10222);
and U10440 (N_10440,N_10227,N_10135);
or U10441 (N_10441,N_10231,N_10115);
or U10442 (N_10442,N_10152,N_10220);
nand U10443 (N_10443,N_10053,N_10013);
and U10444 (N_10444,N_10126,N_10079);
nor U10445 (N_10445,N_10140,N_10215);
or U10446 (N_10446,N_10016,N_10067);
xnor U10447 (N_10447,N_10080,N_10177);
nor U10448 (N_10448,N_10191,N_10096);
nand U10449 (N_10449,N_10121,N_10075);
nor U10450 (N_10450,N_10017,N_10137);
nor U10451 (N_10451,N_10227,N_10025);
nor U10452 (N_10452,N_10230,N_10245);
or U10453 (N_10453,N_10086,N_10043);
or U10454 (N_10454,N_10036,N_10023);
nor U10455 (N_10455,N_10030,N_10218);
nand U10456 (N_10456,N_10080,N_10099);
and U10457 (N_10457,N_10207,N_10034);
and U10458 (N_10458,N_10038,N_10233);
and U10459 (N_10459,N_10132,N_10050);
or U10460 (N_10460,N_10132,N_10064);
or U10461 (N_10461,N_10053,N_10057);
nand U10462 (N_10462,N_10104,N_10177);
and U10463 (N_10463,N_10246,N_10090);
nand U10464 (N_10464,N_10038,N_10144);
nand U10465 (N_10465,N_10106,N_10049);
or U10466 (N_10466,N_10228,N_10070);
nand U10467 (N_10467,N_10135,N_10156);
or U10468 (N_10468,N_10133,N_10016);
and U10469 (N_10469,N_10110,N_10244);
nand U10470 (N_10470,N_10066,N_10101);
nor U10471 (N_10471,N_10008,N_10124);
and U10472 (N_10472,N_10077,N_10088);
xor U10473 (N_10473,N_10184,N_10047);
or U10474 (N_10474,N_10048,N_10062);
or U10475 (N_10475,N_10040,N_10144);
xor U10476 (N_10476,N_10058,N_10203);
nor U10477 (N_10477,N_10248,N_10148);
nand U10478 (N_10478,N_10232,N_10043);
nand U10479 (N_10479,N_10133,N_10015);
or U10480 (N_10480,N_10094,N_10008);
or U10481 (N_10481,N_10137,N_10244);
or U10482 (N_10482,N_10118,N_10160);
and U10483 (N_10483,N_10037,N_10105);
nand U10484 (N_10484,N_10123,N_10028);
or U10485 (N_10485,N_10233,N_10007);
and U10486 (N_10486,N_10202,N_10103);
nor U10487 (N_10487,N_10005,N_10169);
or U10488 (N_10488,N_10114,N_10107);
nor U10489 (N_10489,N_10094,N_10010);
xor U10490 (N_10490,N_10074,N_10042);
nor U10491 (N_10491,N_10180,N_10027);
and U10492 (N_10492,N_10120,N_10152);
and U10493 (N_10493,N_10056,N_10051);
xor U10494 (N_10494,N_10187,N_10219);
and U10495 (N_10495,N_10191,N_10075);
nand U10496 (N_10496,N_10101,N_10190);
nor U10497 (N_10497,N_10077,N_10193);
and U10498 (N_10498,N_10012,N_10019);
and U10499 (N_10499,N_10168,N_10215);
nand U10500 (N_10500,N_10447,N_10342);
and U10501 (N_10501,N_10328,N_10486);
nand U10502 (N_10502,N_10297,N_10429);
and U10503 (N_10503,N_10267,N_10368);
nand U10504 (N_10504,N_10417,N_10490);
and U10505 (N_10505,N_10413,N_10469);
and U10506 (N_10506,N_10268,N_10262);
nand U10507 (N_10507,N_10437,N_10340);
or U10508 (N_10508,N_10364,N_10336);
or U10509 (N_10509,N_10441,N_10420);
or U10510 (N_10510,N_10325,N_10397);
nor U10511 (N_10511,N_10471,N_10444);
nor U10512 (N_10512,N_10485,N_10306);
or U10513 (N_10513,N_10341,N_10299);
and U10514 (N_10514,N_10388,N_10307);
and U10515 (N_10515,N_10439,N_10335);
or U10516 (N_10516,N_10292,N_10457);
and U10517 (N_10517,N_10472,N_10373);
nor U10518 (N_10518,N_10293,N_10301);
nand U10519 (N_10519,N_10319,N_10255);
nor U10520 (N_10520,N_10465,N_10464);
or U10521 (N_10521,N_10354,N_10374);
and U10522 (N_10522,N_10492,N_10452);
xnor U10523 (N_10523,N_10454,N_10488);
nand U10524 (N_10524,N_10385,N_10321);
or U10525 (N_10525,N_10251,N_10445);
or U10526 (N_10526,N_10264,N_10367);
or U10527 (N_10527,N_10481,N_10280);
nand U10528 (N_10528,N_10381,N_10463);
xnor U10529 (N_10529,N_10257,N_10269);
nand U10530 (N_10530,N_10433,N_10432);
nand U10531 (N_10531,N_10270,N_10440);
xnor U10532 (N_10532,N_10379,N_10357);
or U10533 (N_10533,N_10384,N_10311);
nor U10534 (N_10534,N_10499,N_10329);
nor U10535 (N_10535,N_10313,N_10315);
nor U10536 (N_10536,N_10496,N_10322);
nand U10537 (N_10537,N_10460,N_10347);
nor U10538 (N_10538,N_10473,N_10320);
nand U10539 (N_10539,N_10304,N_10375);
and U10540 (N_10540,N_10380,N_10250);
nor U10541 (N_10541,N_10318,N_10482);
or U10542 (N_10542,N_10431,N_10398);
or U10543 (N_10543,N_10273,N_10310);
and U10544 (N_10544,N_10468,N_10491);
xor U10545 (N_10545,N_10324,N_10284);
or U10546 (N_10546,N_10494,N_10344);
or U10547 (N_10547,N_10461,N_10451);
nor U10548 (N_10548,N_10275,N_10434);
and U10549 (N_10549,N_10355,N_10430);
nand U10550 (N_10550,N_10416,N_10300);
or U10551 (N_10551,N_10288,N_10308);
or U10552 (N_10552,N_10415,N_10419);
or U10553 (N_10553,N_10421,N_10286);
nand U10554 (N_10554,N_10309,N_10386);
nor U10555 (N_10555,N_10402,N_10408);
and U10556 (N_10556,N_10462,N_10276);
nand U10557 (N_10557,N_10351,N_10418);
nor U10558 (N_10558,N_10389,N_10303);
and U10559 (N_10559,N_10378,N_10298);
nand U10560 (N_10560,N_10391,N_10317);
or U10561 (N_10561,N_10339,N_10396);
and U10562 (N_10562,N_10281,N_10495);
and U10563 (N_10563,N_10370,N_10338);
nand U10564 (N_10564,N_10424,N_10393);
nand U10565 (N_10565,N_10345,N_10287);
and U10566 (N_10566,N_10356,N_10448);
or U10567 (N_10567,N_10456,N_10400);
nor U10568 (N_10568,N_10478,N_10266);
nand U10569 (N_10569,N_10450,N_10265);
and U10570 (N_10570,N_10332,N_10363);
nand U10571 (N_10571,N_10395,N_10467);
or U10572 (N_10572,N_10372,N_10259);
nand U10573 (N_10573,N_10474,N_10289);
xnor U10574 (N_10574,N_10366,N_10382);
nor U10575 (N_10575,N_10305,N_10483);
nand U10576 (N_10576,N_10428,N_10409);
nor U10577 (N_10577,N_10283,N_10333);
or U10578 (N_10578,N_10302,N_10295);
nor U10579 (N_10579,N_10480,N_10403);
xor U10580 (N_10580,N_10279,N_10487);
or U10581 (N_10581,N_10414,N_10272);
nor U10582 (N_10582,N_10442,N_10412);
and U10583 (N_10583,N_10404,N_10387);
nor U10584 (N_10584,N_10369,N_10476);
nand U10585 (N_10585,N_10405,N_10479);
and U10586 (N_10586,N_10365,N_10326);
and U10587 (N_10587,N_10376,N_10410);
and U10588 (N_10588,N_10498,N_10290);
or U10589 (N_10589,N_10358,N_10453);
nor U10590 (N_10590,N_10263,N_10359);
nand U10591 (N_10591,N_10377,N_10277);
and U10592 (N_10592,N_10425,N_10316);
nor U10593 (N_10593,N_10466,N_10349);
xnor U10594 (N_10594,N_10436,N_10353);
or U10595 (N_10595,N_10252,N_10282);
and U10596 (N_10596,N_10352,N_10362);
or U10597 (N_10597,N_10274,N_10271);
nor U10598 (N_10598,N_10446,N_10477);
or U10599 (N_10599,N_10458,N_10443);
or U10600 (N_10600,N_10406,N_10470);
nand U10601 (N_10601,N_10256,N_10330);
nor U10602 (N_10602,N_10423,N_10296);
nor U10603 (N_10603,N_10348,N_10426);
nor U10604 (N_10604,N_10254,N_10489);
xnor U10605 (N_10605,N_10449,N_10285);
nand U10606 (N_10606,N_10435,N_10371);
nor U10607 (N_10607,N_10360,N_10383);
or U10608 (N_10608,N_10334,N_10343);
nand U10609 (N_10609,N_10392,N_10484);
nor U10610 (N_10610,N_10350,N_10455);
and U10611 (N_10611,N_10312,N_10346);
or U10612 (N_10612,N_10390,N_10407);
or U10613 (N_10613,N_10438,N_10323);
nor U10614 (N_10614,N_10327,N_10258);
and U10615 (N_10615,N_10331,N_10260);
and U10616 (N_10616,N_10291,N_10261);
and U10617 (N_10617,N_10497,N_10493);
and U10618 (N_10618,N_10278,N_10253);
nand U10619 (N_10619,N_10314,N_10361);
nor U10620 (N_10620,N_10422,N_10459);
or U10621 (N_10621,N_10337,N_10294);
or U10622 (N_10622,N_10411,N_10401);
and U10623 (N_10623,N_10399,N_10427);
and U10624 (N_10624,N_10394,N_10475);
and U10625 (N_10625,N_10484,N_10256);
nor U10626 (N_10626,N_10411,N_10367);
nor U10627 (N_10627,N_10334,N_10322);
nand U10628 (N_10628,N_10269,N_10265);
nand U10629 (N_10629,N_10283,N_10393);
nor U10630 (N_10630,N_10384,N_10325);
or U10631 (N_10631,N_10384,N_10386);
or U10632 (N_10632,N_10442,N_10339);
and U10633 (N_10633,N_10380,N_10466);
and U10634 (N_10634,N_10334,N_10357);
or U10635 (N_10635,N_10265,N_10393);
or U10636 (N_10636,N_10266,N_10414);
nor U10637 (N_10637,N_10431,N_10441);
xor U10638 (N_10638,N_10393,N_10474);
and U10639 (N_10639,N_10346,N_10450);
nand U10640 (N_10640,N_10364,N_10394);
nor U10641 (N_10641,N_10274,N_10319);
nor U10642 (N_10642,N_10424,N_10408);
and U10643 (N_10643,N_10493,N_10275);
nand U10644 (N_10644,N_10442,N_10474);
or U10645 (N_10645,N_10312,N_10325);
and U10646 (N_10646,N_10267,N_10482);
or U10647 (N_10647,N_10347,N_10321);
or U10648 (N_10648,N_10369,N_10485);
xnor U10649 (N_10649,N_10379,N_10404);
nand U10650 (N_10650,N_10366,N_10422);
nand U10651 (N_10651,N_10375,N_10366);
nand U10652 (N_10652,N_10401,N_10313);
and U10653 (N_10653,N_10416,N_10353);
nor U10654 (N_10654,N_10375,N_10353);
or U10655 (N_10655,N_10479,N_10489);
or U10656 (N_10656,N_10451,N_10362);
and U10657 (N_10657,N_10450,N_10408);
nand U10658 (N_10658,N_10441,N_10294);
and U10659 (N_10659,N_10475,N_10362);
nor U10660 (N_10660,N_10367,N_10498);
nand U10661 (N_10661,N_10353,N_10271);
nor U10662 (N_10662,N_10493,N_10269);
xnor U10663 (N_10663,N_10476,N_10256);
nor U10664 (N_10664,N_10250,N_10485);
nand U10665 (N_10665,N_10431,N_10396);
nor U10666 (N_10666,N_10354,N_10463);
nand U10667 (N_10667,N_10329,N_10456);
or U10668 (N_10668,N_10439,N_10269);
and U10669 (N_10669,N_10270,N_10295);
nand U10670 (N_10670,N_10485,N_10275);
xor U10671 (N_10671,N_10462,N_10267);
and U10672 (N_10672,N_10474,N_10396);
or U10673 (N_10673,N_10273,N_10308);
nand U10674 (N_10674,N_10371,N_10451);
and U10675 (N_10675,N_10368,N_10482);
xnor U10676 (N_10676,N_10328,N_10436);
and U10677 (N_10677,N_10373,N_10483);
or U10678 (N_10678,N_10308,N_10345);
or U10679 (N_10679,N_10342,N_10387);
and U10680 (N_10680,N_10437,N_10435);
or U10681 (N_10681,N_10283,N_10311);
nand U10682 (N_10682,N_10479,N_10444);
and U10683 (N_10683,N_10455,N_10462);
nor U10684 (N_10684,N_10454,N_10396);
or U10685 (N_10685,N_10490,N_10412);
xnor U10686 (N_10686,N_10315,N_10470);
xor U10687 (N_10687,N_10324,N_10362);
nand U10688 (N_10688,N_10352,N_10376);
xnor U10689 (N_10689,N_10402,N_10253);
nor U10690 (N_10690,N_10346,N_10270);
xor U10691 (N_10691,N_10492,N_10443);
nor U10692 (N_10692,N_10474,N_10303);
or U10693 (N_10693,N_10352,N_10436);
or U10694 (N_10694,N_10320,N_10477);
nand U10695 (N_10695,N_10417,N_10406);
and U10696 (N_10696,N_10491,N_10256);
xnor U10697 (N_10697,N_10373,N_10328);
nor U10698 (N_10698,N_10324,N_10454);
or U10699 (N_10699,N_10458,N_10362);
and U10700 (N_10700,N_10335,N_10487);
and U10701 (N_10701,N_10458,N_10366);
nand U10702 (N_10702,N_10339,N_10492);
and U10703 (N_10703,N_10307,N_10375);
nand U10704 (N_10704,N_10253,N_10259);
or U10705 (N_10705,N_10337,N_10479);
or U10706 (N_10706,N_10321,N_10307);
nor U10707 (N_10707,N_10296,N_10408);
and U10708 (N_10708,N_10427,N_10364);
nor U10709 (N_10709,N_10495,N_10375);
nor U10710 (N_10710,N_10419,N_10350);
or U10711 (N_10711,N_10446,N_10361);
and U10712 (N_10712,N_10355,N_10294);
or U10713 (N_10713,N_10499,N_10254);
nand U10714 (N_10714,N_10484,N_10405);
nor U10715 (N_10715,N_10471,N_10273);
nand U10716 (N_10716,N_10431,N_10261);
xnor U10717 (N_10717,N_10373,N_10414);
xor U10718 (N_10718,N_10427,N_10371);
or U10719 (N_10719,N_10333,N_10257);
nor U10720 (N_10720,N_10314,N_10432);
and U10721 (N_10721,N_10418,N_10342);
or U10722 (N_10722,N_10491,N_10364);
xor U10723 (N_10723,N_10447,N_10297);
xnor U10724 (N_10724,N_10388,N_10411);
or U10725 (N_10725,N_10277,N_10484);
or U10726 (N_10726,N_10250,N_10393);
nand U10727 (N_10727,N_10302,N_10279);
and U10728 (N_10728,N_10388,N_10264);
nor U10729 (N_10729,N_10313,N_10378);
nor U10730 (N_10730,N_10424,N_10360);
nor U10731 (N_10731,N_10473,N_10381);
or U10732 (N_10732,N_10348,N_10275);
nor U10733 (N_10733,N_10365,N_10485);
or U10734 (N_10734,N_10472,N_10435);
and U10735 (N_10735,N_10401,N_10468);
or U10736 (N_10736,N_10400,N_10387);
or U10737 (N_10737,N_10286,N_10402);
or U10738 (N_10738,N_10303,N_10449);
nand U10739 (N_10739,N_10309,N_10320);
xnor U10740 (N_10740,N_10267,N_10279);
xor U10741 (N_10741,N_10392,N_10409);
or U10742 (N_10742,N_10397,N_10416);
nor U10743 (N_10743,N_10305,N_10425);
nor U10744 (N_10744,N_10368,N_10465);
or U10745 (N_10745,N_10259,N_10471);
or U10746 (N_10746,N_10424,N_10299);
and U10747 (N_10747,N_10481,N_10402);
or U10748 (N_10748,N_10408,N_10327);
nor U10749 (N_10749,N_10446,N_10297);
xor U10750 (N_10750,N_10684,N_10681);
and U10751 (N_10751,N_10542,N_10706);
or U10752 (N_10752,N_10677,N_10553);
or U10753 (N_10753,N_10733,N_10630);
or U10754 (N_10754,N_10705,N_10722);
and U10755 (N_10755,N_10683,N_10697);
xor U10756 (N_10756,N_10587,N_10664);
or U10757 (N_10757,N_10564,N_10600);
xnor U10758 (N_10758,N_10682,N_10624);
nor U10759 (N_10759,N_10583,N_10736);
nand U10760 (N_10760,N_10525,N_10535);
or U10761 (N_10761,N_10709,N_10640);
and U10762 (N_10762,N_10718,N_10744);
nand U10763 (N_10763,N_10719,N_10698);
nor U10764 (N_10764,N_10612,N_10531);
nor U10765 (N_10765,N_10580,N_10659);
nor U10766 (N_10766,N_10575,N_10685);
and U10767 (N_10767,N_10721,N_10549);
nor U10768 (N_10768,N_10699,N_10579);
nor U10769 (N_10769,N_10539,N_10732);
or U10770 (N_10770,N_10626,N_10691);
nand U10771 (N_10771,N_10550,N_10712);
nor U10772 (N_10772,N_10651,N_10572);
nand U10773 (N_10773,N_10545,N_10582);
and U10774 (N_10774,N_10599,N_10704);
or U10775 (N_10775,N_10703,N_10638);
xor U10776 (N_10776,N_10688,N_10506);
xnor U10777 (N_10777,N_10660,N_10727);
or U10778 (N_10778,N_10653,N_10510);
nand U10779 (N_10779,N_10577,N_10538);
and U10780 (N_10780,N_10696,N_10647);
nor U10781 (N_10781,N_10594,N_10505);
and U10782 (N_10782,N_10522,N_10708);
or U10783 (N_10783,N_10702,N_10657);
or U10784 (N_10784,N_10578,N_10745);
nor U10785 (N_10785,N_10610,N_10687);
nand U10786 (N_10786,N_10556,N_10649);
or U10787 (N_10787,N_10526,N_10738);
or U10788 (N_10788,N_10536,N_10500);
and U10789 (N_10789,N_10734,N_10631);
nor U10790 (N_10790,N_10748,N_10590);
or U10791 (N_10791,N_10723,N_10670);
nor U10792 (N_10792,N_10547,N_10554);
nand U10793 (N_10793,N_10747,N_10606);
nor U10794 (N_10794,N_10637,N_10715);
nand U10795 (N_10795,N_10707,N_10695);
nand U10796 (N_10796,N_10509,N_10596);
and U10797 (N_10797,N_10552,N_10743);
nand U10798 (N_10798,N_10532,N_10728);
nand U10799 (N_10799,N_10650,N_10585);
nand U10800 (N_10800,N_10725,N_10665);
nand U10801 (N_10801,N_10669,N_10543);
or U10802 (N_10802,N_10571,N_10645);
nand U10803 (N_10803,N_10513,N_10512);
nand U10804 (N_10804,N_10658,N_10690);
or U10805 (N_10805,N_10740,N_10518);
nand U10806 (N_10806,N_10666,N_10652);
xnor U10807 (N_10807,N_10613,N_10678);
nand U10808 (N_10808,N_10668,N_10636);
and U10809 (N_10809,N_10559,N_10676);
and U10810 (N_10810,N_10726,N_10591);
nand U10811 (N_10811,N_10656,N_10546);
or U10812 (N_10812,N_10621,N_10633);
nor U10813 (N_10813,N_10581,N_10604);
and U10814 (N_10814,N_10503,N_10551);
and U10815 (N_10815,N_10517,N_10627);
nand U10816 (N_10816,N_10662,N_10735);
xor U10817 (N_10817,N_10573,N_10502);
xor U10818 (N_10818,N_10739,N_10720);
nand U10819 (N_10819,N_10516,N_10584);
nand U10820 (N_10820,N_10729,N_10618);
and U10821 (N_10821,N_10561,N_10701);
or U10822 (N_10822,N_10615,N_10567);
nand U10823 (N_10823,N_10574,N_10616);
and U10824 (N_10824,N_10519,N_10614);
or U10825 (N_10825,N_10557,N_10528);
xnor U10826 (N_10826,N_10661,N_10529);
and U10827 (N_10827,N_10592,N_10694);
or U10828 (N_10828,N_10537,N_10501);
and U10829 (N_10829,N_10540,N_10623);
and U10830 (N_10830,N_10597,N_10511);
and U10831 (N_10831,N_10741,N_10639);
or U10832 (N_10832,N_10541,N_10524);
or U10833 (N_10833,N_10625,N_10686);
nand U10834 (N_10834,N_10504,N_10544);
or U10835 (N_10835,N_10566,N_10737);
nand U10836 (N_10836,N_10731,N_10565);
and U10837 (N_10837,N_10634,N_10742);
nor U10838 (N_10838,N_10508,N_10643);
xnor U10839 (N_10839,N_10560,N_10558);
and U10840 (N_10840,N_10534,N_10632);
nor U10841 (N_10841,N_10588,N_10679);
or U10842 (N_10842,N_10689,N_10514);
xnor U10843 (N_10843,N_10644,N_10622);
nand U10844 (N_10844,N_10555,N_10716);
nand U10845 (N_10845,N_10602,N_10680);
nor U10846 (N_10846,N_10717,N_10533);
nand U10847 (N_10847,N_10654,N_10607);
and U10848 (N_10848,N_10724,N_10609);
nor U10849 (N_10849,N_10713,N_10507);
nand U10850 (N_10850,N_10730,N_10593);
nor U10851 (N_10851,N_10675,N_10629);
nor U10852 (N_10852,N_10749,N_10562);
xnor U10853 (N_10853,N_10628,N_10673);
or U10854 (N_10854,N_10521,N_10548);
nor U10855 (N_10855,N_10586,N_10601);
nand U10856 (N_10856,N_10527,N_10563);
nand U10857 (N_10857,N_10692,N_10611);
and U10858 (N_10858,N_10605,N_10710);
nor U10859 (N_10859,N_10520,N_10570);
and U10860 (N_10860,N_10569,N_10648);
or U10861 (N_10861,N_10619,N_10603);
and U10862 (N_10862,N_10693,N_10714);
or U10863 (N_10863,N_10700,N_10617);
nand U10864 (N_10864,N_10711,N_10646);
and U10865 (N_10865,N_10746,N_10576);
nor U10866 (N_10866,N_10620,N_10671);
nand U10867 (N_10867,N_10530,N_10608);
nand U10868 (N_10868,N_10667,N_10663);
or U10869 (N_10869,N_10635,N_10642);
or U10870 (N_10870,N_10515,N_10595);
nand U10871 (N_10871,N_10589,N_10674);
nor U10872 (N_10872,N_10523,N_10655);
xnor U10873 (N_10873,N_10598,N_10672);
nand U10874 (N_10874,N_10641,N_10568);
or U10875 (N_10875,N_10730,N_10599);
and U10876 (N_10876,N_10705,N_10553);
and U10877 (N_10877,N_10666,N_10539);
nand U10878 (N_10878,N_10517,N_10689);
and U10879 (N_10879,N_10504,N_10567);
nand U10880 (N_10880,N_10507,N_10728);
nor U10881 (N_10881,N_10618,N_10684);
or U10882 (N_10882,N_10683,N_10667);
or U10883 (N_10883,N_10576,N_10610);
or U10884 (N_10884,N_10526,N_10510);
or U10885 (N_10885,N_10530,N_10615);
and U10886 (N_10886,N_10639,N_10580);
and U10887 (N_10887,N_10564,N_10541);
nand U10888 (N_10888,N_10614,N_10511);
nor U10889 (N_10889,N_10656,N_10601);
xor U10890 (N_10890,N_10532,N_10525);
or U10891 (N_10891,N_10687,N_10547);
xor U10892 (N_10892,N_10541,N_10631);
xnor U10893 (N_10893,N_10520,N_10579);
nor U10894 (N_10894,N_10611,N_10660);
or U10895 (N_10895,N_10554,N_10524);
or U10896 (N_10896,N_10510,N_10545);
or U10897 (N_10897,N_10556,N_10523);
or U10898 (N_10898,N_10646,N_10601);
nand U10899 (N_10899,N_10692,N_10653);
nor U10900 (N_10900,N_10742,N_10679);
nor U10901 (N_10901,N_10604,N_10729);
or U10902 (N_10902,N_10503,N_10502);
or U10903 (N_10903,N_10513,N_10595);
and U10904 (N_10904,N_10568,N_10655);
nor U10905 (N_10905,N_10579,N_10555);
nand U10906 (N_10906,N_10605,N_10611);
and U10907 (N_10907,N_10602,N_10641);
nor U10908 (N_10908,N_10508,N_10666);
nand U10909 (N_10909,N_10517,N_10732);
nand U10910 (N_10910,N_10699,N_10562);
xnor U10911 (N_10911,N_10727,N_10587);
nand U10912 (N_10912,N_10527,N_10660);
or U10913 (N_10913,N_10721,N_10527);
or U10914 (N_10914,N_10731,N_10605);
nor U10915 (N_10915,N_10708,N_10639);
or U10916 (N_10916,N_10637,N_10557);
nor U10917 (N_10917,N_10661,N_10579);
nor U10918 (N_10918,N_10541,N_10565);
and U10919 (N_10919,N_10524,N_10594);
nor U10920 (N_10920,N_10692,N_10629);
nor U10921 (N_10921,N_10573,N_10653);
nor U10922 (N_10922,N_10544,N_10547);
or U10923 (N_10923,N_10531,N_10742);
xor U10924 (N_10924,N_10544,N_10737);
nand U10925 (N_10925,N_10585,N_10644);
and U10926 (N_10926,N_10571,N_10511);
xor U10927 (N_10927,N_10662,N_10641);
nor U10928 (N_10928,N_10678,N_10562);
xor U10929 (N_10929,N_10555,N_10715);
nand U10930 (N_10930,N_10744,N_10612);
nand U10931 (N_10931,N_10668,N_10665);
nand U10932 (N_10932,N_10514,N_10583);
xnor U10933 (N_10933,N_10657,N_10558);
or U10934 (N_10934,N_10605,N_10728);
and U10935 (N_10935,N_10532,N_10566);
and U10936 (N_10936,N_10505,N_10652);
and U10937 (N_10937,N_10748,N_10517);
or U10938 (N_10938,N_10547,N_10526);
and U10939 (N_10939,N_10537,N_10707);
and U10940 (N_10940,N_10676,N_10598);
and U10941 (N_10941,N_10735,N_10669);
nand U10942 (N_10942,N_10574,N_10729);
nand U10943 (N_10943,N_10566,N_10702);
and U10944 (N_10944,N_10671,N_10581);
or U10945 (N_10945,N_10572,N_10646);
nor U10946 (N_10946,N_10550,N_10614);
or U10947 (N_10947,N_10642,N_10588);
nand U10948 (N_10948,N_10584,N_10740);
or U10949 (N_10949,N_10608,N_10714);
xnor U10950 (N_10950,N_10567,N_10565);
nand U10951 (N_10951,N_10638,N_10510);
xor U10952 (N_10952,N_10729,N_10683);
or U10953 (N_10953,N_10591,N_10548);
nand U10954 (N_10954,N_10677,N_10562);
or U10955 (N_10955,N_10651,N_10696);
or U10956 (N_10956,N_10672,N_10601);
nand U10957 (N_10957,N_10603,N_10672);
or U10958 (N_10958,N_10585,N_10573);
and U10959 (N_10959,N_10722,N_10664);
nor U10960 (N_10960,N_10597,N_10631);
and U10961 (N_10961,N_10518,N_10583);
and U10962 (N_10962,N_10653,N_10532);
nand U10963 (N_10963,N_10573,N_10725);
nor U10964 (N_10964,N_10575,N_10594);
and U10965 (N_10965,N_10699,N_10615);
nor U10966 (N_10966,N_10676,N_10605);
or U10967 (N_10967,N_10588,N_10568);
and U10968 (N_10968,N_10557,N_10609);
or U10969 (N_10969,N_10748,N_10539);
and U10970 (N_10970,N_10631,N_10569);
nor U10971 (N_10971,N_10586,N_10505);
and U10972 (N_10972,N_10529,N_10623);
or U10973 (N_10973,N_10502,N_10730);
nand U10974 (N_10974,N_10570,N_10692);
or U10975 (N_10975,N_10659,N_10555);
or U10976 (N_10976,N_10559,N_10522);
and U10977 (N_10977,N_10605,N_10659);
nor U10978 (N_10978,N_10568,N_10525);
or U10979 (N_10979,N_10626,N_10715);
or U10980 (N_10980,N_10647,N_10610);
and U10981 (N_10981,N_10732,N_10688);
nand U10982 (N_10982,N_10736,N_10574);
or U10983 (N_10983,N_10520,N_10686);
nor U10984 (N_10984,N_10643,N_10627);
xnor U10985 (N_10985,N_10686,N_10585);
nand U10986 (N_10986,N_10713,N_10689);
nor U10987 (N_10987,N_10707,N_10574);
nand U10988 (N_10988,N_10580,N_10719);
and U10989 (N_10989,N_10607,N_10590);
nand U10990 (N_10990,N_10500,N_10623);
and U10991 (N_10991,N_10715,N_10550);
or U10992 (N_10992,N_10630,N_10679);
or U10993 (N_10993,N_10605,N_10570);
or U10994 (N_10994,N_10581,N_10542);
or U10995 (N_10995,N_10692,N_10598);
nand U10996 (N_10996,N_10723,N_10592);
nor U10997 (N_10997,N_10538,N_10593);
nor U10998 (N_10998,N_10703,N_10568);
or U10999 (N_10999,N_10533,N_10695);
xnor U11000 (N_11000,N_10908,N_10791);
nor U11001 (N_11001,N_10949,N_10947);
nand U11002 (N_11002,N_10801,N_10961);
or U11003 (N_11003,N_10829,N_10965);
nand U11004 (N_11004,N_10865,N_10782);
nand U11005 (N_11005,N_10983,N_10786);
nor U11006 (N_11006,N_10846,N_10996);
or U11007 (N_11007,N_10939,N_10906);
nor U11008 (N_11008,N_10836,N_10884);
or U11009 (N_11009,N_10752,N_10938);
nand U11010 (N_11010,N_10942,N_10788);
nor U11011 (N_11011,N_10831,N_10826);
or U11012 (N_11012,N_10835,N_10860);
nor U11013 (N_11013,N_10819,N_10794);
nand U11014 (N_11014,N_10844,N_10963);
and U11015 (N_11015,N_10785,N_10857);
nand U11016 (N_11016,N_10759,N_10795);
nand U11017 (N_11017,N_10951,N_10837);
nor U11018 (N_11018,N_10799,N_10764);
and U11019 (N_11019,N_10883,N_10854);
and U11020 (N_11020,N_10851,N_10888);
nand U11021 (N_11021,N_10910,N_10903);
and U11022 (N_11022,N_10989,N_10870);
nand U11023 (N_11023,N_10887,N_10962);
nor U11024 (N_11024,N_10978,N_10976);
nand U11025 (N_11025,N_10885,N_10789);
xor U11026 (N_11026,N_10915,N_10967);
xnor U11027 (N_11027,N_10895,N_10891);
nor U11028 (N_11028,N_10973,N_10850);
nor U11029 (N_11029,N_10918,N_10800);
xor U11030 (N_11030,N_10867,N_10925);
nor U11031 (N_11031,N_10838,N_10928);
and U11032 (N_11032,N_10796,N_10950);
nand U11033 (N_11033,N_10769,N_10761);
xnor U11034 (N_11034,N_10811,N_10827);
or U11035 (N_11035,N_10899,N_10964);
xnor U11036 (N_11036,N_10790,N_10913);
nor U11037 (N_11037,N_10914,N_10817);
nand U11038 (N_11038,N_10856,N_10970);
and U11039 (N_11039,N_10815,N_10926);
nor U11040 (N_11040,N_10999,N_10921);
nor U11041 (N_11041,N_10853,N_10905);
or U11042 (N_11042,N_10880,N_10927);
and U11043 (N_11043,N_10841,N_10936);
nor U11044 (N_11044,N_10784,N_10992);
nor U11045 (N_11045,N_10776,N_10832);
and U11046 (N_11046,N_10792,N_10974);
nor U11047 (N_11047,N_10798,N_10855);
nand U11048 (N_11048,N_10787,N_10802);
and U11049 (N_11049,N_10988,N_10783);
nor U11050 (N_11050,N_10822,N_10881);
nand U11051 (N_11051,N_10772,N_10842);
and U11052 (N_11052,N_10780,N_10893);
and U11053 (N_11053,N_10966,N_10777);
nand U11054 (N_11054,N_10773,N_10755);
and U11055 (N_11055,N_10944,N_10872);
or U11056 (N_11056,N_10991,N_10753);
nor U11057 (N_11057,N_10808,N_10863);
and U11058 (N_11058,N_10882,N_10834);
xor U11059 (N_11059,N_10980,N_10797);
nand U11060 (N_11060,N_10778,N_10843);
and U11061 (N_11061,N_10848,N_10897);
nand U11062 (N_11062,N_10852,N_10806);
and U11063 (N_11063,N_10859,N_10960);
and U11064 (N_11064,N_10821,N_10902);
xor U11065 (N_11065,N_10779,N_10953);
nand U11066 (N_11066,N_10775,N_10941);
nand U11067 (N_11067,N_10833,N_10985);
nand U11068 (N_11068,N_10820,N_10824);
and U11069 (N_11069,N_10896,N_10898);
xor U11070 (N_11070,N_10793,N_10760);
nand U11071 (N_11071,N_10814,N_10876);
and U11072 (N_11072,N_10758,N_10868);
nor U11073 (N_11073,N_10892,N_10931);
and U11074 (N_11074,N_10968,N_10877);
nor U11075 (N_11075,N_10917,N_10981);
and U11076 (N_11076,N_10809,N_10803);
nand U11077 (N_11077,N_10889,N_10957);
or U11078 (N_11078,N_10812,N_10971);
xor U11079 (N_11079,N_10932,N_10823);
or U11080 (N_11080,N_10750,N_10767);
and U11081 (N_11081,N_10924,N_10945);
nor U11082 (N_11082,N_10756,N_10904);
and U11083 (N_11083,N_10858,N_10922);
nor U11084 (N_11084,N_10886,N_10804);
and U11085 (N_11085,N_10975,N_10986);
nor U11086 (N_11086,N_10982,N_10977);
or U11087 (N_11087,N_10940,N_10900);
nand U11088 (N_11088,N_10781,N_10825);
and U11089 (N_11089,N_10762,N_10816);
or U11090 (N_11090,N_10879,N_10774);
nor U11091 (N_11091,N_10768,N_10770);
and U11092 (N_11092,N_10923,N_10845);
and U11093 (N_11093,N_10861,N_10765);
nand U11094 (N_11094,N_10955,N_10813);
xnor U11095 (N_11095,N_10956,N_10995);
nor U11096 (N_11096,N_10912,N_10890);
and U11097 (N_11097,N_10958,N_10840);
or U11098 (N_11098,N_10935,N_10934);
nand U11099 (N_11099,N_10972,N_10993);
nand U11100 (N_11100,N_10839,N_10997);
and U11101 (N_11101,N_10771,N_10866);
nor U11102 (N_11102,N_10828,N_10984);
nor U11103 (N_11103,N_10937,N_10959);
and U11104 (N_11104,N_10849,N_10919);
nor U11105 (N_11105,N_10990,N_10871);
nand U11106 (N_11106,N_10763,N_10979);
nand U11107 (N_11107,N_10916,N_10907);
nor U11108 (N_11108,N_10930,N_10754);
nor U11109 (N_11109,N_10869,N_10998);
or U11110 (N_11110,N_10911,N_10873);
nor U11111 (N_11111,N_10994,N_10818);
nor U11112 (N_11112,N_10954,N_10952);
or U11113 (N_11113,N_10757,N_10943);
and U11114 (N_11114,N_10807,N_10987);
nand U11115 (N_11115,N_10969,N_10810);
nand U11116 (N_11116,N_10948,N_10946);
and U11117 (N_11117,N_10901,N_10864);
nor U11118 (N_11118,N_10847,N_10894);
xor U11119 (N_11119,N_10874,N_10751);
nor U11120 (N_11120,N_10805,N_10875);
nand U11121 (N_11121,N_10929,N_10920);
nor U11122 (N_11122,N_10830,N_10933);
nor U11123 (N_11123,N_10909,N_10766);
and U11124 (N_11124,N_10878,N_10862);
nand U11125 (N_11125,N_10960,N_10966);
nor U11126 (N_11126,N_10904,N_10853);
or U11127 (N_11127,N_10979,N_10757);
and U11128 (N_11128,N_10865,N_10904);
or U11129 (N_11129,N_10963,N_10765);
and U11130 (N_11130,N_10835,N_10866);
nor U11131 (N_11131,N_10971,N_10827);
nand U11132 (N_11132,N_10757,N_10949);
nor U11133 (N_11133,N_10782,N_10768);
or U11134 (N_11134,N_10988,N_10794);
or U11135 (N_11135,N_10961,N_10953);
nand U11136 (N_11136,N_10970,N_10880);
nand U11137 (N_11137,N_10771,N_10864);
or U11138 (N_11138,N_10821,N_10792);
nand U11139 (N_11139,N_10794,N_10772);
nor U11140 (N_11140,N_10794,N_10853);
xor U11141 (N_11141,N_10971,N_10985);
or U11142 (N_11142,N_10967,N_10964);
and U11143 (N_11143,N_10837,N_10986);
nand U11144 (N_11144,N_10996,N_10797);
and U11145 (N_11145,N_10883,N_10976);
nor U11146 (N_11146,N_10775,N_10883);
and U11147 (N_11147,N_10775,N_10906);
or U11148 (N_11148,N_10960,N_10951);
nand U11149 (N_11149,N_10757,N_10904);
or U11150 (N_11150,N_10790,N_10856);
nand U11151 (N_11151,N_10934,N_10796);
nor U11152 (N_11152,N_10914,N_10944);
nand U11153 (N_11153,N_10841,N_10863);
and U11154 (N_11154,N_10940,N_10920);
nand U11155 (N_11155,N_10800,N_10923);
nor U11156 (N_11156,N_10774,N_10965);
nand U11157 (N_11157,N_10793,N_10843);
and U11158 (N_11158,N_10924,N_10931);
xnor U11159 (N_11159,N_10976,N_10874);
xnor U11160 (N_11160,N_10786,N_10882);
nor U11161 (N_11161,N_10949,N_10930);
nand U11162 (N_11162,N_10830,N_10805);
or U11163 (N_11163,N_10996,N_10995);
or U11164 (N_11164,N_10958,N_10841);
or U11165 (N_11165,N_10892,N_10859);
or U11166 (N_11166,N_10879,N_10983);
nor U11167 (N_11167,N_10769,N_10921);
nor U11168 (N_11168,N_10871,N_10960);
nor U11169 (N_11169,N_10859,N_10905);
xor U11170 (N_11170,N_10938,N_10846);
nand U11171 (N_11171,N_10981,N_10776);
nor U11172 (N_11172,N_10855,N_10842);
xnor U11173 (N_11173,N_10763,N_10946);
and U11174 (N_11174,N_10915,N_10903);
nand U11175 (N_11175,N_10780,N_10960);
nor U11176 (N_11176,N_10955,N_10843);
and U11177 (N_11177,N_10754,N_10761);
nor U11178 (N_11178,N_10862,N_10920);
and U11179 (N_11179,N_10900,N_10897);
nor U11180 (N_11180,N_10798,N_10994);
and U11181 (N_11181,N_10795,N_10944);
or U11182 (N_11182,N_10873,N_10895);
or U11183 (N_11183,N_10940,N_10925);
nor U11184 (N_11184,N_10944,N_10762);
and U11185 (N_11185,N_10788,N_10777);
or U11186 (N_11186,N_10966,N_10766);
or U11187 (N_11187,N_10981,N_10957);
and U11188 (N_11188,N_10958,N_10801);
nor U11189 (N_11189,N_10868,N_10898);
nor U11190 (N_11190,N_10752,N_10935);
xor U11191 (N_11191,N_10982,N_10961);
and U11192 (N_11192,N_10863,N_10801);
or U11193 (N_11193,N_10977,N_10756);
and U11194 (N_11194,N_10770,N_10803);
or U11195 (N_11195,N_10786,N_10795);
nand U11196 (N_11196,N_10994,N_10754);
nor U11197 (N_11197,N_10982,N_10930);
nand U11198 (N_11198,N_10752,N_10956);
xor U11199 (N_11199,N_10956,N_10886);
or U11200 (N_11200,N_10766,N_10841);
nor U11201 (N_11201,N_10767,N_10923);
nand U11202 (N_11202,N_10843,N_10988);
xnor U11203 (N_11203,N_10983,N_10849);
nand U11204 (N_11204,N_10868,N_10982);
and U11205 (N_11205,N_10934,N_10871);
xnor U11206 (N_11206,N_10788,N_10803);
nor U11207 (N_11207,N_10868,N_10958);
and U11208 (N_11208,N_10961,N_10846);
nand U11209 (N_11209,N_10772,N_10824);
and U11210 (N_11210,N_10948,N_10863);
nand U11211 (N_11211,N_10950,N_10953);
nor U11212 (N_11212,N_10876,N_10919);
nand U11213 (N_11213,N_10752,N_10876);
nor U11214 (N_11214,N_10877,N_10937);
or U11215 (N_11215,N_10928,N_10888);
or U11216 (N_11216,N_10979,N_10929);
nand U11217 (N_11217,N_10972,N_10776);
and U11218 (N_11218,N_10953,N_10945);
or U11219 (N_11219,N_10889,N_10926);
nand U11220 (N_11220,N_10954,N_10797);
nand U11221 (N_11221,N_10997,N_10931);
nand U11222 (N_11222,N_10918,N_10929);
nand U11223 (N_11223,N_10843,N_10860);
and U11224 (N_11224,N_10971,N_10942);
nor U11225 (N_11225,N_10758,N_10883);
nand U11226 (N_11226,N_10877,N_10868);
or U11227 (N_11227,N_10948,N_10857);
and U11228 (N_11228,N_10871,N_10767);
nor U11229 (N_11229,N_10878,N_10814);
or U11230 (N_11230,N_10915,N_10895);
or U11231 (N_11231,N_10907,N_10765);
or U11232 (N_11232,N_10828,N_10768);
and U11233 (N_11233,N_10870,N_10903);
or U11234 (N_11234,N_10750,N_10817);
or U11235 (N_11235,N_10931,N_10915);
or U11236 (N_11236,N_10780,N_10924);
and U11237 (N_11237,N_10850,N_10843);
nand U11238 (N_11238,N_10944,N_10800);
nand U11239 (N_11239,N_10818,N_10949);
and U11240 (N_11240,N_10828,N_10779);
nand U11241 (N_11241,N_10819,N_10877);
or U11242 (N_11242,N_10825,N_10797);
and U11243 (N_11243,N_10976,N_10955);
or U11244 (N_11244,N_10937,N_10764);
xor U11245 (N_11245,N_10934,N_10835);
xnor U11246 (N_11246,N_10846,N_10759);
nor U11247 (N_11247,N_10800,N_10901);
or U11248 (N_11248,N_10788,N_10933);
or U11249 (N_11249,N_10782,N_10853);
and U11250 (N_11250,N_11094,N_11047);
nor U11251 (N_11251,N_11230,N_11079);
or U11252 (N_11252,N_11063,N_11195);
xor U11253 (N_11253,N_11081,N_11090);
or U11254 (N_11254,N_11169,N_11035);
and U11255 (N_11255,N_11186,N_11159);
xnor U11256 (N_11256,N_11241,N_11140);
and U11257 (N_11257,N_11189,N_11158);
or U11258 (N_11258,N_11232,N_11043);
or U11259 (N_11259,N_11089,N_11190);
nand U11260 (N_11260,N_11045,N_11187);
nand U11261 (N_11261,N_11068,N_11072);
and U11262 (N_11262,N_11175,N_11226);
or U11263 (N_11263,N_11182,N_11016);
nand U11264 (N_11264,N_11152,N_11073);
or U11265 (N_11265,N_11174,N_11212);
or U11266 (N_11266,N_11000,N_11070);
nand U11267 (N_11267,N_11021,N_11117);
nor U11268 (N_11268,N_11123,N_11141);
nor U11269 (N_11269,N_11163,N_11139);
and U11270 (N_11270,N_11246,N_11065);
nor U11271 (N_11271,N_11151,N_11106);
xnor U11272 (N_11272,N_11233,N_11091);
nor U11273 (N_11273,N_11087,N_11059);
nand U11274 (N_11274,N_11040,N_11207);
or U11275 (N_11275,N_11206,N_11228);
or U11276 (N_11276,N_11054,N_11034);
and U11277 (N_11277,N_11166,N_11044);
and U11278 (N_11278,N_11014,N_11067);
and U11279 (N_11279,N_11080,N_11027);
or U11280 (N_11280,N_11099,N_11135);
nand U11281 (N_11281,N_11053,N_11064);
nor U11282 (N_11282,N_11240,N_11078);
nand U11283 (N_11283,N_11062,N_11136);
and U11284 (N_11284,N_11013,N_11172);
nand U11285 (N_11285,N_11126,N_11235);
or U11286 (N_11286,N_11179,N_11180);
or U11287 (N_11287,N_11196,N_11248);
nand U11288 (N_11288,N_11008,N_11088);
nand U11289 (N_11289,N_11096,N_11191);
nor U11290 (N_11290,N_11120,N_11066);
xnor U11291 (N_11291,N_11029,N_11109);
or U11292 (N_11292,N_11074,N_11007);
and U11293 (N_11293,N_11222,N_11188);
or U11294 (N_11294,N_11161,N_11092);
and U11295 (N_11295,N_11134,N_11162);
nand U11296 (N_11296,N_11153,N_11198);
nor U11297 (N_11297,N_11076,N_11193);
xnor U11298 (N_11298,N_11102,N_11024);
or U11299 (N_11299,N_11224,N_11055);
or U11300 (N_11300,N_11133,N_11015);
nor U11301 (N_11301,N_11083,N_11234);
or U11302 (N_11302,N_11002,N_11142);
and U11303 (N_11303,N_11049,N_11150);
or U11304 (N_11304,N_11113,N_11143);
nor U11305 (N_11305,N_11114,N_11071);
and U11306 (N_11306,N_11243,N_11157);
or U11307 (N_11307,N_11116,N_11184);
nand U11308 (N_11308,N_11178,N_11130);
nor U11309 (N_11309,N_11156,N_11108);
or U11310 (N_11310,N_11165,N_11085);
nor U11311 (N_11311,N_11192,N_11218);
or U11312 (N_11312,N_11170,N_11009);
xor U11313 (N_11313,N_11038,N_11220);
xor U11314 (N_11314,N_11176,N_11125);
and U11315 (N_11315,N_11075,N_11211);
nor U11316 (N_11316,N_11118,N_11046);
nor U11317 (N_11317,N_11204,N_11030);
nand U11318 (N_11318,N_11115,N_11041);
and U11319 (N_11319,N_11048,N_11105);
nand U11320 (N_11320,N_11210,N_11132);
or U11321 (N_11321,N_11237,N_11214);
nand U11322 (N_11322,N_11229,N_11056);
and U11323 (N_11323,N_11127,N_11011);
or U11324 (N_11324,N_11112,N_11052);
nor U11325 (N_11325,N_11095,N_11148);
nor U11326 (N_11326,N_11242,N_11205);
xnor U11327 (N_11327,N_11168,N_11203);
nand U11328 (N_11328,N_11051,N_11098);
and U11329 (N_11329,N_11208,N_11181);
nand U11330 (N_11330,N_11122,N_11005);
nand U11331 (N_11331,N_11171,N_11032);
nand U11332 (N_11332,N_11057,N_11017);
and U11333 (N_11333,N_11003,N_11202);
nand U11334 (N_11334,N_11145,N_11209);
or U11335 (N_11335,N_11238,N_11033);
and U11336 (N_11336,N_11215,N_11037);
nor U11337 (N_11337,N_11042,N_11110);
and U11338 (N_11338,N_11077,N_11197);
and U11339 (N_11339,N_11001,N_11167);
or U11340 (N_11340,N_11213,N_11023);
nand U11341 (N_11341,N_11050,N_11173);
nor U11342 (N_11342,N_11147,N_11177);
or U11343 (N_11343,N_11058,N_11039);
nand U11344 (N_11344,N_11100,N_11154);
and U11345 (N_11345,N_11216,N_11144);
xor U11346 (N_11346,N_11138,N_11101);
or U11347 (N_11347,N_11061,N_11128);
or U11348 (N_11348,N_11103,N_11107);
nand U11349 (N_11349,N_11119,N_11146);
and U11350 (N_11350,N_11164,N_11244);
and U11351 (N_11351,N_11006,N_11239);
or U11352 (N_11352,N_11086,N_11084);
nor U11353 (N_11353,N_11149,N_11010);
xnor U11354 (N_11354,N_11111,N_11247);
nor U11355 (N_11355,N_11160,N_11225);
and U11356 (N_11356,N_11022,N_11245);
nor U11357 (N_11357,N_11185,N_11227);
xor U11358 (N_11358,N_11137,N_11082);
and U11359 (N_11359,N_11201,N_11236);
nor U11360 (N_11360,N_11129,N_11012);
nor U11361 (N_11361,N_11097,N_11018);
or U11362 (N_11362,N_11249,N_11231);
nor U11363 (N_11363,N_11200,N_11026);
nand U11364 (N_11364,N_11019,N_11155);
xnor U11365 (N_11365,N_11036,N_11028);
nand U11366 (N_11366,N_11217,N_11093);
or U11367 (N_11367,N_11223,N_11069);
or U11368 (N_11368,N_11183,N_11219);
and U11369 (N_11369,N_11194,N_11060);
nand U11370 (N_11370,N_11199,N_11131);
and U11371 (N_11371,N_11025,N_11104);
or U11372 (N_11372,N_11031,N_11121);
or U11373 (N_11373,N_11004,N_11124);
and U11374 (N_11374,N_11221,N_11020);
nor U11375 (N_11375,N_11123,N_11046);
nand U11376 (N_11376,N_11058,N_11134);
nand U11377 (N_11377,N_11015,N_11230);
xnor U11378 (N_11378,N_11085,N_11156);
and U11379 (N_11379,N_11242,N_11101);
or U11380 (N_11380,N_11055,N_11178);
xor U11381 (N_11381,N_11043,N_11013);
and U11382 (N_11382,N_11149,N_11186);
xnor U11383 (N_11383,N_11132,N_11238);
nand U11384 (N_11384,N_11049,N_11129);
or U11385 (N_11385,N_11104,N_11042);
or U11386 (N_11386,N_11245,N_11204);
and U11387 (N_11387,N_11093,N_11120);
nand U11388 (N_11388,N_11174,N_11111);
or U11389 (N_11389,N_11023,N_11162);
nand U11390 (N_11390,N_11030,N_11027);
and U11391 (N_11391,N_11152,N_11063);
and U11392 (N_11392,N_11024,N_11060);
or U11393 (N_11393,N_11087,N_11039);
nand U11394 (N_11394,N_11187,N_11123);
nand U11395 (N_11395,N_11084,N_11168);
or U11396 (N_11396,N_11218,N_11038);
nor U11397 (N_11397,N_11180,N_11197);
and U11398 (N_11398,N_11216,N_11073);
nor U11399 (N_11399,N_11044,N_11240);
and U11400 (N_11400,N_11025,N_11182);
and U11401 (N_11401,N_11142,N_11189);
nand U11402 (N_11402,N_11206,N_11212);
and U11403 (N_11403,N_11171,N_11119);
or U11404 (N_11404,N_11133,N_11167);
nor U11405 (N_11405,N_11174,N_11242);
or U11406 (N_11406,N_11158,N_11141);
and U11407 (N_11407,N_11094,N_11218);
and U11408 (N_11408,N_11249,N_11011);
or U11409 (N_11409,N_11238,N_11065);
or U11410 (N_11410,N_11149,N_11157);
nand U11411 (N_11411,N_11125,N_11037);
nor U11412 (N_11412,N_11042,N_11209);
nor U11413 (N_11413,N_11157,N_11207);
nor U11414 (N_11414,N_11090,N_11144);
or U11415 (N_11415,N_11221,N_11038);
nor U11416 (N_11416,N_11101,N_11104);
nor U11417 (N_11417,N_11180,N_11158);
nand U11418 (N_11418,N_11236,N_11041);
and U11419 (N_11419,N_11160,N_11148);
nand U11420 (N_11420,N_11234,N_11189);
nand U11421 (N_11421,N_11111,N_11027);
nand U11422 (N_11422,N_11164,N_11089);
nor U11423 (N_11423,N_11109,N_11232);
nand U11424 (N_11424,N_11216,N_11191);
or U11425 (N_11425,N_11230,N_11168);
nor U11426 (N_11426,N_11162,N_11039);
nand U11427 (N_11427,N_11215,N_11042);
nand U11428 (N_11428,N_11009,N_11217);
xnor U11429 (N_11429,N_11249,N_11002);
and U11430 (N_11430,N_11034,N_11216);
xor U11431 (N_11431,N_11154,N_11177);
nand U11432 (N_11432,N_11044,N_11114);
or U11433 (N_11433,N_11194,N_11164);
or U11434 (N_11434,N_11222,N_11142);
or U11435 (N_11435,N_11132,N_11153);
or U11436 (N_11436,N_11101,N_11047);
or U11437 (N_11437,N_11023,N_11066);
or U11438 (N_11438,N_11001,N_11084);
and U11439 (N_11439,N_11209,N_11175);
or U11440 (N_11440,N_11219,N_11065);
nand U11441 (N_11441,N_11020,N_11004);
nand U11442 (N_11442,N_11018,N_11106);
or U11443 (N_11443,N_11116,N_11159);
or U11444 (N_11444,N_11015,N_11070);
or U11445 (N_11445,N_11107,N_11222);
and U11446 (N_11446,N_11225,N_11248);
nand U11447 (N_11447,N_11126,N_11037);
and U11448 (N_11448,N_11182,N_11190);
nor U11449 (N_11449,N_11162,N_11009);
and U11450 (N_11450,N_11103,N_11184);
and U11451 (N_11451,N_11137,N_11241);
nor U11452 (N_11452,N_11201,N_11191);
nor U11453 (N_11453,N_11037,N_11102);
or U11454 (N_11454,N_11193,N_11130);
nor U11455 (N_11455,N_11129,N_11199);
or U11456 (N_11456,N_11217,N_11131);
nor U11457 (N_11457,N_11040,N_11136);
nor U11458 (N_11458,N_11094,N_11188);
nor U11459 (N_11459,N_11220,N_11056);
xnor U11460 (N_11460,N_11226,N_11020);
xor U11461 (N_11461,N_11200,N_11169);
and U11462 (N_11462,N_11049,N_11076);
nand U11463 (N_11463,N_11021,N_11089);
and U11464 (N_11464,N_11049,N_11059);
nand U11465 (N_11465,N_11156,N_11038);
and U11466 (N_11466,N_11160,N_11085);
xnor U11467 (N_11467,N_11026,N_11125);
nor U11468 (N_11468,N_11094,N_11120);
nor U11469 (N_11469,N_11194,N_11212);
and U11470 (N_11470,N_11081,N_11234);
nand U11471 (N_11471,N_11072,N_11228);
nand U11472 (N_11472,N_11176,N_11054);
and U11473 (N_11473,N_11031,N_11064);
or U11474 (N_11474,N_11155,N_11214);
nand U11475 (N_11475,N_11025,N_11244);
nor U11476 (N_11476,N_11234,N_11239);
nor U11477 (N_11477,N_11205,N_11222);
and U11478 (N_11478,N_11095,N_11180);
or U11479 (N_11479,N_11054,N_11221);
xor U11480 (N_11480,N_11012,N_11218);
nand U11481 (N_11481,N_11095,N_11133);
xnor U11482 (N_11482,N_11225,N_11247);
or U11483 (N_11483,N_11174,N_11021);
and U11484 (N_11484,N_11194,N_11181);
nand U11485 (N_11485,N_11040,N_11100);
and U11486 (N_11486,N_11057,N_11000);
nand U11487 (N_11487,N_11124,N_11040);
and U11488 (N_11488,N_11166,N_11189);
and U11489 (N_11489,N_11050,N_11008);
or U11490 (N_11490,N_11109,N_11156);
nor U11491 (N_11491,N_11164,N_11095);
and U11492 (N_11492,N_11230,N_11118);
nor U11493 (N_11493,N_11047,N_11121);
nor U11494 (N_11494,N_11134,N_11247);
nand U11495 (N_11495,N_11129,N_11024);
xnor U11496 (N_11496,N_11036,N_11121);
nand U11497 (N_11497,N_11081,N_11078);
and U11498 (N_11498,N_11244,N_11040);
nand U11499 (N_11499,N_11196,N_11155);
and U11500 (N_11500,N_11334,N_11275);
or U11501 (N_11501,N_11399,N_11499);
nand U11502 (N_11502,N_11273,N_11310);
and U11503 (N_11503,N_11440,N_11250);
or U11504 (N_11504,N_11422,N_11442);
and U11505 (N_11505,N_11402,N_11487);
or U11506 (N_11506,N_11360,N_11471);
xnor U11507 (N_11507,N_11337,N_11267);
nand U11508 (N_11508,N_11465,N_11414);
or U11509 (N_11509,N_11287,N_11394);
and U11510 (N_11510,N_11293,N_11466);
nand U11511 (N_11511,N_11362,N_11482);
xnor U11512 (N_11512,N_11305,N_11332);
nor U11513 (N_11513,N_11354,N_11307);
nand U11514 (N_11514,N_11411,N_11285);
and U11515 (N_11515,N_11484,N_11406);
xor U11516 (N_11516,N_11387,N_11451);
nor U11517 (N_11517,N_11283,N_11377);
or U11518 (N_11518,N_11476,N_11381);
nand U11519 (N_11519,N_11308,N_11404);
nand U11520 (N_11520,N_11265,N_11398);
xnor U11521 (N_11521,N_11468,N_11461);
nand U11522 (N_11522,N_11369,N_11376);
or U11523 (N_11523,N_11481,N_11258);
nand U11524 (N_11524,N_11346,N_11251);
nor U11525 (N_11525,N_11426,N_11493);
or U11526 (N_11526,N_11445,N_11455);
and U11527 (N_11527,N_11252,N_11313);
and U11528 (N_11528,N_11338,N_11450);
xor U11529 (N_11529,N_11435,N_11384);
or U11530 (N_11530,N_11311,N_11254);
nor U11531 (N_11531,N_11460,N_11412);
or U11532 (N_11532,N_11457,N_11361);
nor U11533 (N_11533,N_11424,N_11456);
and U11534 (N_11534,N_11486,N_11474);
or U11535 (N_11535,N_11470,N_11320);
xnor U11536 (N_11536,N_11292,N_11357);
or U11537 (N_11537,N_11453,N_11423);
nand U11538 (N_11538,N_11255,N_11278);
nand U11539 (N_11539,N_11301,N_11359);
nor U11540 (N_11540,N_11467,N_11421);
nor U11541 (N_11541,N_11400,N_11336);
and U11542 (N_11542,N_11295,N_11473);
and U11543 (N_11543,N_11356,N_11304);
nand U11544 (N_11544,N_11492,N_11444);
nand U11545 (N_11545,N_11291,N_11419);
and U11546 (N_11546,N_11259,N_11438);
xor U11547 (N_11547,N_11270,N_11284);
or U11548 (N_11548,N_11389,N_11347);
and U11549 (N_11549,N_11317,N_11345);
nand U11550 (N_11550,N_11319,N_11263);
or U11551 (N_11551,N_11396,N_11318);
and U11552 (N_11552,N_11316,N_11328);
nor U11553 (N_11553,N_11405,N_11324);
and U11554 (N_11554,N_11418,N_11430);
nor U11555 (N_11555,N_11358,N_11483);
nor U11556 (N_11556,N_11416,N_11350);
nand U11557 (N_11557,N_11459,N_11458);
and U11558 (N_11558,N_11296,N_11323);
and U11559 (N_11559,N_11397,N_11367);
nand U11560 (N_11560,N_11299,N_11410);
nor U11561 (N_11561,N_11441,N_11490);
or U11562 (N_11562,N_11344,N_11371);
xnor U11563 (N_11563,N_11428,N_11447);
and U11564 (N_11564,N_11494,N_11348);
and U11565 (N_11565,N_11335,N_11298);
nor U11566 (N_11566,N_11495,N_11463);
nor U11567 (N_11567,N_11409,N_11443);
and U11568 (N_11568,N_11480,N_11253);
nand U11569 (N_11569,N_11417,N_11448);
nand U11570 (N_11570,N_11407,N_11368);
nor U11571 (N_11571,N_11329,N_11330);
or U11572 (N_11572,N_11326,N_11327);
and U11573 (N_11573,N_11322,N_11390);
nand U11574 (N_11574,N_11341,N_11333);
nand U11575 (N_11575,N_11446,N_11268);
xnor U11576 (N_11576,N_11439,N_11365);
nand U11577 (N_11577,N_11343,N_11286);
nand U11578 (N_11578,N_11314,N_11415);
or U11579 (N_11579,N_11437,N_11498);
xnor U11580 (N_11580,N_11478,N_11432);
and U11581 (N_11581,N_11315,N_11372);
xor U11582 (N_11582,N_11454,N_11276);
and U11583 (N_11583,N_11256,N_11289);
nor U11584 (N_11584,N_11279,N_11385);
xor U11585 (N_11585,N_11366,N_11340);
or U11586 (N_11586,N_11271,N_11420);
and U11587 (N_11587,N_11373,N_11272);
or U11588 (N_11588,N_11370,N_11325);
nand U11589 (N_11589,N_11485,N_11434);
nand U11590 (N_11590,N_11374,N_11294);
and U11591 (N_11591,N_11309,N_11331);
and U11592 (N_11592,N_11477,N_11302);
and U11593 (N_11593,N_11306,N_11469);
nand U11594 (N_11594,N_11433,N_11497);
nor U11595 (N_11595,N_11408,N_11277);
nor U11596 (N_11596,N_11452,N_11393);
nand U11597 (N_11597,N_11349,N_11281);
nor U11598 (N_11598,N_11431,N_11378);
and U11599 (N_11599,N_11363,N_11262);
and U11600 (N_11600,N_11403,N_11479);
nand U11601 (N_11601,N_11472,N_11496);
or U11602 (N_11602,N_11489,N_11383);
and U11603 (N_11603,N_11475,N_11364);
nand U11604 (N_11604,N_11355,N_11375);
and U11605 (N_11605,N_11464,N_11392);
and U11606 (N_11606,N_11342,N_11266);
nor U11607 (N_11607,N_11257,N_11395);
and U11608 (N_11608,N_11339,N_11351);
or U11609 (N_11609,N_11401,N_11462);
nor U11610 (N_11610,N_11282,N_11386);
nand U11611 (N_11611,N_11321,N_11413);
nand U11612 (N_11612,N_11427,N_11379);
nor U11613 (N_11613,N_11449,N_11382);
xor U11614 (N_11614,N_11269,N_11391);
nand U11615 (N_11615,N_11425,N_11290);
and U11616 (N_11616,N_11436,N_11353);
and U11617 (N_11617,N_11380,N_11303);
xor U11618 (N_11618,N_11300,N_11280);
xor U11619 (N_11619,N_11264,N_11297);
nor U11620 (N_11620,N_11274,N_11260);
nor U11621 (N_11621,N_11261,N_11491);
or U11622 (N_11622,N_11352,N_11388);
xnor U11623 (N_11623,N_11429,N_11312);
and U11624 (N_11624,N_11488,N_11288);
nand U11625 (N_11625,N_11487,N_11380);
nand U11626 (N_11626,N_11384,N_11432);
nand U11627 (N_11627,N_11264,N_11405);
nand U11628 (N_11628,N_11497,N_11392);
nor U11629 (N_11629,N_11371,N_11359);
nand U11630 (N_11630,N_11483,N_11399);
and U11631 (N_11631,N_11395,N_11414);
nand U11632 (N_11632,N_11306,N_11395);
or U11633 (N_11633,N_11468,N_11276);
nand U11634 (N_11634,N_11278,N_11475);
or U11635 (N_11635,N_11379,N_11327);
or U11636 (N_11636,N_11302,N_11468);
nor U11637 (N_11637,N_11468,N_11319);
xnor U11638 (N_11638,N_11298,N_11278);
or U11639 (N_11639,N_11349,N_11352);
xnor U11640 (N_11640,N_11425,N_11453);
nand U11641 (N_11641,N_11339,N_11385);
or U11642 (N_11642,N_11327,N_11335);
nand U11643 (N_11643,N_11373,N_11296);
and U11644 (N_11644,N_11324,N_11393);
nand U11645 (N_11645,N_11422,N_11250);
or U11646 (N_11646,N_11283,N_11375);
nand U11647 (N_11647,N_11471,N_11409);
or U11648 (N_11648,N_11429,N_11278);
and U11649 (N_11649,N_11345,N_11404);
nor U11650 (N_11650,N_11266,N_11268);
nor U11651 (N_11651,N_11365,N_11460);
xor U11652 (N_11652,N_11429,N_11263);
nor U11653 (N_11653,N_11348,N_11394);
and U11654 (N_11654,N_11477,N_11296);
and U11655 (N_11655,N_11322,N_11400);
nand U11656 (N_11656,N_11449,N_11463);
or U11657 (N_11657,N_11452,N_11272);
and U11658 (N_11658,N_11438,N_11470);
nor U11659 (N_11659,N_11450,N_11461);
nand U11660 (N_11660,N_11404,N_11275);
and U11661 (N_11661,N_11348,N_11285);
nand U11662 (N_11662,N_11459,N_11349);
nand U11663 (N_11663,N_11433,N_11292);
or U11664 (N_11664,N_11351,N_11390);
nor U11665 (N_11665,N_11342,N_11322);
nand U11666 (N_11666,N_11491,N_11359);
xnor U11667 (N_11667,N_11405,N_11378);
or U11668 (N_11668,N_11491,N_11304);
nand U11669 (N_11669,N_11311,N_11271);
nor U11670 (N_11670,N_11434,N_11254);
nor U11671 (N_11671,N_11298,N_11301);
and U11672 (N_11672,N_11427,N_11421);
and U11673 (N_11673,N_11462,N_11429);
and U11674 (N_11674,N_11257,N_11393);
and U11675 (N_11675,N_11489,N_11392);
nor U11676 (N_11676,N_11254,N_11408);
nor U11677 (N_11677,N_11496,N_11495);
or U11678 (N_11678,N_11368,N_11319);
nor U11679 (N_11679,N_11431,N_11401);
or U11680 (N_11680,N_11426,N_11429);
nand U11681 (N_11681,N_11337,N_11251);
and U11682 (N_11682,N_11347,N_11250);
and U11683 (N_11683,N_11490,N_11419);
nor U11684 (N_11684,N_11277,N_11264);
or U11685 (N_11685,N_11320,N_11256);
nand U11686 (N_11686,N_11454,N_11467);
and U11687 (N_11687,N_11331,N_11365);
xor U11688 (N_11688,N_11449,N_11259);
or U11689 (N_11689,N_11255,N_11340);
nand U11690 (N_11690,N_11324,N_11312);
and U11691 (N_11691,N_11268,N_11344);
nor U11692 (N_11692,N_11268,N_11280);
or U11693 (N_11693,N_11427,N_11269);
xor U11694 (N_11694,N_11478,N_11467);
nand U11695 (N_11695,N_11470,N_11445);
nor U11696 (N_11696,N_11434,N_11336);
or U11697 (N_11697,N_11473,N_11381);
nand U11698 (N_11698,N_11447,N_11339);
nor U11699 (N_11699,N_11430,N_11453);
nor U11700 (N_11700,N_11452,N_11370);
nor U11701 (N_11701,N_11388,N_11337);
xor U11702 (N_11702,N_11365,N_11318);
nor U11703 (N_11703,N_11498,N_11399);
and U11704 (N_11704,N_11418,N_11340);
xor U11705 (N_11705,N_11340,N_11498);
and U11706 (N_11706,N_11481,N_11409);
or U11707 (N_11707,N_11343,N_11386);
nand U11708 (N_11708,N_11316,N_11438);
and U11709 (N_11709,N_11495,N_11492);
or U11710 (N_11710,N_11443,N_11375);
xor U11711 (N_11711,N_11265,N_11403);
and U11712 (N_11712,N_11364,N_11262);
nor U11713 (N_11713,N_11432,N_11409);
nor U11714 (N_11714,N_11380,N_11273);
and U11715 (N_11715,N_11388,N_11376);
nor U11716 (N_11716,N_11484,N_11382);
nor U11717 (N_11717,N_11362,N_11473);
nor U11718 (N_11718,N_11429,N_11371);
nand U11719 (N_11719,N_11310,N_11340);
nand U11720 (N_11720,N_11379,N_11410);
nand U11721 (N_11721,N_11261,N_11321);
or U11722 (N_11722,N_11344,N_11316);
nor U11723 (N_11723,N_11379,N_11484);
nand U11724 (N_11724,N_11381,N_11317);
nand U11725 (N_11725,N_11477,N_11412);
nand U11726 (N_11726,N_11417,N_11432);
or U11727 (N_11727,N_11380,N_11460);
or U11728 (N_11728,N_11258,N_11485);
and U11729 (N_11729,N_11431,N_11487);
nand U11730 (N_11730,N_11399,N_11269);
or U11731 (N_11731,N_11393,N_11384);
and U11732 (N_11732,N_11421,N_11436);
nor U11733 (N_11733,N_11481,N_11331);
or U11734 (N_11734,N_11472,N_11300);
or U11735 (N_11735,N_11427,N_11317);
nor U11736 (N_11736,N_11453,N_11495);
nand U11737 (N_11737,N_11269,N_11499);
and U11738 (N_11738,N_11421,N_11447);
nor U11739 (N_11739,N_11457,N_11412);
or U11740 (N_11740,N_11398,N_11498);
and U11741 (N_11741,N_11418,N_11328);
or U11742 (N_11742,N_11252,N_11292);
xnor U11743 (N_11743,N_11449,N_11491);
or U11744 (N_11744,N_11354,N_11469);
nand U11745 (N_11745,N_11498,N_11371);
or U11746 (N_11746,N_11406,N_11316);
or U11747 (N_11747,N_11434,N_11348);
nand U11748 (N_11748,N_11408,N_11419);
nor U11749 (N_11749,N_11495,N_11396);
and U11750 (N_11750,N_11507,N_11595);
nand U11751 (N_11751,N_11566,N_11710);
or U11752 (N_11752,N_11689,N_11702);
and U11753 (N_11753,N_11735,N_11630);
nand U11754 (N_11754,N_11746,N_11587);
or U11755 (N_11755,N_11502,N_11637);
nand U11756 (N_11756,N_11600,N_11680);
and U11757 (N_11757,N_11516,N_11576);
nand U11758 (N_11758,N_11557,N_11588);
nand U11759 (N_11759,N_11635,N_11552);
nor U11760 (N_11760,N_11596,N_11504);
xor U11761 (N_11761,N_11603,N_11733);
or U11762 (N_11762,N_11741,N_11505);
and U11763 (N_11763,N_11738,N_11580);
nor U11764 (N_11764,N_11568,N_11619);
nor U11765 (N_11765,N_11565,N_11695);
nand U11766 (N_11766,N_11511,N_11650);
nand U11767 (N_11767,N_11656,N_11701);
nand U11768 (N_11768,N_11717,N_11745);
and U11769 (N_11769,N_11744,N_11612);
nand U11770 (N_11770,N_11642,N_11697);
and U11771 (N_11771,N_11714,N_11520);
nor U11772 (N_11772,N_11524,N_11513);
or U11773 (N_11773,N_11669,N_11626);
nor U11774 (N_11774,N_11665,N_11657);
nand U11775 (N_11775,N_11547,N_11724);
nand U11776 (N_11776,N_11574,N_11641);
or U11777 (N_11777,N_11748,N_11616);
or U11778 (N_11778,N_11585,N_11549);
and U11779 (N_11779,N_11518,N_11737);
xor U11780 (N_11780,N_11571,N_11646);
nand U11781 (N_11781,N_11655,N_11506);
nor U11782 (N_11782,N_11608,N_11685);
and U11783 (N_11783,N_11601,N_11698);
nor U11784 (N_11784,N_11525,N_11592);
and U11785 (N_11785,N_11584,N_11562);
nand U11786 (N_11786,N_11666,N_11614);
nor U11787 (N_11787,N_11687,N_11602);
and U11788 (N_11788,N_11621,N_11530);
and U11789 (N_11789,N_11572,N_11540);
nor U11790 (N_11790,N_11720,N_11501);
or U11791 (N_11791,N_11664,N_11703);
nor U11792 (N_11792,N_11629,N_11672);
nand U11793 (N_11793,N_11545,N_11747);
nand U11794 (N_11794,N_11509,N_11597);
and U11795 (N_11795,N_11648,N_11719);
nand U11796 (N_11796,N_11712,N_11508);
nand U11797 (N_11797,N_11512,N_11654);
or U11798 (N_11798,N_11586,N_11681);
nand U11799 (N_11799,N_11716,N_11636);
xnor U11800 (N_11800,N_11652,N_11613);
nand U11801 (N_11801,N_11644,N_11628);
nor U11802 (N_11802,N_11688,N_11554);
nand U11803 (N_11803,N_11734,N_11618);
and U11804 (N_11804,N_11573,N_11694);
nor U11805 (N_11805,N_11544,N_11531);
nor U11806 (N_11806,N_11532,N_11667);
nor U11807 (N_11807,N_11577,N_11670);
nand U11808 (N_11808,N_11503,N_11625);
or U11809 (N_11809,N_11591,N_11740);
or U11810 (N_11810,N_11742,N_11521);
nor U11811 (N_11811,N_11709,N_11707);
and U11812 (N_11812,N_11539,N_11510);
xnor U11813 (N_11813,N_11555,N_11711);
xor U11814 (N_11814,N_11677,N_11522);
and U11815 (N_11815,N_11564,N_11579);
xnor U11816 (N_11816,N_11556,N_11583);
nor U11817 (N_11817,N_11668,N_11643);
nor U11818 (N_11818,N_11634,N_11721);
and U11819 (N_11819,N_11699,N_11682);
nand U11820 (N_11820,N_11627,N_11684);
nand U11821 (N_11821,N_11558,N_11663);
or U11822 (N_11822,N_11623,N_11693);
or U11823 (N_11823,N_11610,N_11582);
or U11824 (N_11824,N_11659,N_11599);
nor U11825 (N_11825,N_11569,N_11514);
xor U11826 (N_11826,N_11575,N_11683);
nand U11827 (N_11827,N_11671,N_11723);
or U11828 (N_11828,N_11662,N_11515);
and U11829 (N_11829,N_11749,N_11728);
or U11830 (N_11830,N_11686,N_11611);
xor U11831 (N_11831,N_11551,N_11606);
and U11832 (N_11832,N_11624,N_11675);
nand U11833 (N_11833,N_11739,N_11553);
and U11834 (N_11834,N_11559,N_11560);
or U11835 (N_11835,N_11543,N_11632);
or U11836 (N_11836,N_11658,N_11535);
nand U11837 (N_11837,N_11528,N_11718);
nor U11838 (N_11838,N_11526,N_11651);
and U11839 (N_11839,N_11519,N_11696);
nor U11840 (N_11840,N_11639,N_11529);
nand U11841 (N_11841,N_11722,N_11660);
nand U11842 (N_11842,N_11607,N_11645);
or U11843 (N_11843,N_11700,N_11534);
and U11844 (N_11844,N_11638,N_11715);
nand U11845 (N_11845,N_11609,N_11673);
xnor U11846 (N_11846,N_11726,N_11500);
and U11847 (N_11847,N_11620,N_11713);
nand U11848 (N_11848,N_11548,N_11706);
nand U11849 (N_11849,N_11589,N_11676);
or U11850 (N_11850,N_11705,N_11615);
nor U11851 (N_11851,N_11727,N_11550);
nand U11852 (N_11852,N_11640,N_11536);
or U11853 (N_11853,N_11725,N_11537);
or U11854 (N_11854,N_11661,N_11593);
nand U11855 (N_11855,N_11679,N_11729);
nor U11856 (N_11856,N_11563,N_11736);
nor U11857 (N_11857,N_11570,N_11567);
nand U11858 (N_11858,N_11517,N_11598);
nor U11859 (N_11859,N_11743,N_11578);
and U11860 (N_11860,N_11581,N_11617);
and U11861 (N_11861,N_11542,N_11546);
nor U11862 (N_11862,N_11594,N_11674);
or U11863 (N_11863,N_11732,N_11647);
nand U11864 (N_11864,N_11631,N_11523);
nor U11865 (N_11865,N_11538,N_11692);
xnor U11866 (N_11866,N_11541,N_11622);
and U11867 (N_11867,N_11704,N_11690);
xor U11868 (N_11868,N_11649,N_11633);
nor U11869 (N_11869,N_11533,N_11590);
xor U11870 (N_11870,N_11678,N_11731);
nand U11871 (N_11871,N_11691,N_11527);
and U11872 (N_11872,N_11730,N_11653);
or U11873 (N_11873,N_11604,N_11708);
and U11874 (N_11874,N_11561,N_11605);
and U11875 (N_11875,N_11581,N_11586);
nand U11876 (N_11876,N_11698,N_11575);
xnor U11877 (N_11877,N_11692,N_11504);
or U11878 (N_11878,N_11688,N_11686);
nand U11879 (N_11879,N_11730,N_11648);
or U11880 (N_11880,N_11606,N_11628);
nor U11881 (N_11881,N_11561,N_11737);
nand U11882 (N_11882,N_11664,N_11686);
xor U11883 (N_11883,N_11683,N_11612);
nor U11884 (N_11884,N_11622,N_11702);
and U11885 (N_11885,N_11656,N_11703);
nor U11886 (N_11886,N_11564,N_11729);
and U11887 (N_11887,N_11682,N_11617);
nand U11888 (N_11888,N_11644,N_11526);
nand U11889 (N_11889,N_11691,N_11525);
and U11890 (N_11890,N_11734,N_11580);
or U11891 (N_11891,N_11678,N_11728);
and U11892 (N_11892,N_11561,N_11744);
or U11893 (N_11893,N_11609,N_11528);
xnor U11894 (N_11894,N_11512,N_11671);
or U11895 (N_11895,N_11664,N_11506);
or U11896 (N_11896,N_11729,N_11617);
nor U11897 (N_11897,N_11627,N_11727);
and U11898 (N_11898,N_11736,N_11599);
and U11899 (N_11899,N_11541,N_11554);
nor U11900 (N_11900,N_11608,N_11509);
or U11901 (N_11901,N_11630,N_11548);
nor U11902 (N_11902,N_11603,N_11681);
nand U11903 (N_11903,N_11564,N_11508);
nor U11904 (N_11904,N_11713,N_11699);
nor U11905 (N_11905,N_11738,N_11577);
or U11906 (N_11906,N_11621,N_11548);
or U11907 (N_11907,N_11668,N_11591);
nor U11908 (N_11908,N_11670,N_11671);
nor U11909 (N_11909,N_11666,N_11516);
and U11910 (N_11910,N_11532,N_11689);
nand U11911 (N_11911,N_11726,N_11589);
and U11912 (N_11912,N_11560,N_11640);
nand U11913 (N_11913,N_11647,N_11648);
nor U11914 (N_11914,N_11713,N_11568);
and U11915 (N_11915,N_11541,N_11546);
xor U11916 (N_11916,N_11567,N_11719);
and U11917 (N_11917,N_11591,N_11546);
or U11918 (N_11918,N_11639,N_11701);
nand U11919 (N_11919,N_11583,N_11635);
nor U11920 (N_11920,N_11601,N_11576);
nand U11921 (N_11921,N_11620,N_11612);
or U11922 (N_11922,N_11562,N_11645);
nand U11923 (N_11923,N_11595,N_11512);
or U11924 (N_11924,N_11543,N_11703);
and U11925 (N_11925,N_11554,N_11675);
or U11926 (N_11926,N_11576,N_11558);
and U11927 (N_11927,N_11704,N_11566);
and U11928 (N_11928,N_11586,N_11646);
and U11929 (N_11929,N_11613,N_11582);
nand U11930 (N_11930,N_11737,N_11732);
and U11931 (N_11931,N_11705,N_11574);
nand U11932 (N_11932,N_11604,N_11726);
xnor U11933 (N_11933,N_11740,N_11674);
xnor U11934 (N_11934,N_11556,N_11590);
nand U11935 (N_11935,N_11706,N_11500);
or U11936 (N_11936,N_11538,N_11543);
nand U11937 (N_11937,N_11659,N_11638);
xnor U11938 (N_11938,N_11570,N_11558);
nand U11939 (N_11939,N_11605,N_11707);
nor U11940 (N_11940,N_11618,N_11727);
or U11941 (N_11941,N_11547,N_11548);
or U11942 (N_11942,N_11746,N_11618);
nor U11943 (N_11943,N_11633,N_11674);
or U11944 (N_11944,N_11577,N_11594);
and U11945 (N_11945,N_11735,N_11708);
or U11946 (N_11946,N_11713,N_11520);
nand U11947 (N_11947,N_11657,N_11656);
nand U11948 (N_11948,N_11602,N_11685);
nor U11949 (N_11949,N_11628,N_11702);
nor U11950 (N_11950,N_11702,N_11505);
or U11951 (N_11951,N_11631,N_11709);
and U11952 (N_11952,N_11656,N_11535);
nor U11953 (N_11953,N_11610,N_11630);
nand U11954 (N_11954,N_11643,N_11531);
xor U11955 (N_11955,N_11580,N_11639);
or U11956 (N_11956,N_11559,N_11747);
or U11957 (N_11957,N_11586,N_11527);
xor U11958 (N_11958,N_11639,N_11629);
xnor U11959 (N_11959,N_11675,N_11690);
or U11960 (N_11960,N_11648,N_11620);
nor U11961 (N_11961,N_11610,N_11651);
or U11962 (N_11962,N_11708,N_11722);
nor U11963 (N_11963,N_11674,N_11716);
and U11964 (N_11964,N_11693,N_11592);
nor U11965 (N_11965,N_11692,N_11712);
and U11966 (N_11966,N_11535,N_11540);
or U11967 (N_11967,N_11637,N_11700);
nand U11968 (N_11968,N_11658,N_11614);
nor U11969 (N_11969,N_11646,N_11585);
xor U11970 (N_11970,N_11642,N_11573);
or U11971 (N_11971,N_11663,N_11729);
and U11972 (N_11972,N_11555,N_11553);
or U11973 (N_11973,N_11707,N_11501);
nand U11974 (N_11974,N_11653,N_11549);
or U11975 (N_11975,N_11700,N_11738);
nor U11976 (N_11976,N_11648,N_11518);
nor U11977 (N_11977,N_11727,N_11528);
nand U11978 (N_11978,N_11727,N_11743);
and U11979 (N_11979,N_11606,N_11739);
xnor U11980 (N_11980,N_11584,N_11606);
nand U11981 (N_11981,N_11548,N_11624);
nand U11982 (N_11982,N_11600,N_11630);
nand U11983 (N_11983,N_11674,N_11707);
or U11984 (N_11984,N_11721,N_11743);
or U11985 (N_11985,N_11545,N_11671);
nor U11986 (N_11986,N_11528,N_11546);
or U11987 (N_11987,N_11562,N_11726);
and U11988 (N_11988,N_11537,N_11637);
or U11989 (N_11989,N_11645,N_11564);
and U11990 (N_11990,N_11718,N_11653);
nor U11991 (N_11991,N_11501,N_11744);
and U11992 (N_11992,N_11703,N_11583);
and U11993 (N_11993,N_11596,N_11588);
nand U11994 (N_11994,N_11543,N_11519);
and U11995 (N_11995,N_11563,N_11588);
nor U11996 (N_11996,N_11552,N_11711);
and U11997 (N_11997,N_11526,N_11538);
and U11998 (N_11998,N_11677,N_11739);
and U11999 (N_11999,N_11614,N_11644);
and U12000 (N_12000,N_11883,N_11856);
nor U12001 (N_12001,N_11898,N_11851);
or U12002 (N_12002,N_11817,N_11795);
and U12003 (N_12003,N_11997,N_11879);
nor U12004 (N_12004,N_11855,N_11853);
and U12005 (N_12005,N_11822,N_11917);
or U12006 (N_12006,N_11774,N_11801);
or U12007 (N_12007,N_11869,N_11874);
and U12008 (N_12008,N_11836,N_11779);
nor U12009 (N_12009,N_11842,N_11990);
or U12010 (N_12010,N_11937,N_11957);
and U12011 (N_12011,N_11992,N_11766);
and U12012 (N_12012,N_11888,N_11909);
nand U12013 (N_12013,N_11803,N_11929);
nand U12014 (N_12014,N_11945,N_11861);
or U12015 (N_12015,N_11982,N_11828);
xor U12016 (N_12016,N_11981,N_11897);
nor U12017 (N_12017,N_11802,N_11798);
nor U12018 (N_12018,N_11872,N_11931);
xor U12019 (N_12019,N_11833,N_11991);
and U12020 (N_12020,N_11913,N_11846);
or U12021 (N_12021,N_11885,N_11860);
xor U12022 (N_12022,N_11960,N_11811);
or U12023 (N_12023,N_11791,N_11995);
or U12024 (N_12024,N_11825,N_11865);
nand U12025 (N_12025,N_11938,N_11902);
nor U12026 (N_12026,N_11771,N_11948);
nand U12027 (N_12027,N_11764,N_11984);
and U12028 (N_12028,N_11841,N_11914);
or U12029 (N_12029,N_11763,N_11788);
nand U12030 (N_12030,N_11958,N_11889);
nor U12031 (N_12031,N_11829,N_11906);
nor U12032 (N_12032,N_11893,N_11794);
and U12033 (N_12033,N_11873,N_11904);
or U12034 (N_12034,N_11839,N_11975);
nor U12035 (N_12035,N_11890,N_11800);
and U12036 (N_12036,N_11778,N_11963);
nand U12037 (N_12037,N_11993,N_11980);
or U12038 (N_12038,N_11934,N_11949);
nor U12039 (N_12039,N_11767,N_11773);
nor U12040 (N_12040,N_11910,N_11866);
nand U12041 (N_12041,N_11871,N_11759);
nand U12042 (N_12042,N_11862,N_11810);
or U12043 (N_12043,N_11988,N_11944);
nand U12044 (N_12044,N_11940,N_11790);
or U12045 (N_12045,N_11837,N_11813);
or U12046 (N_12046,N_11905,N_11830);
or U12047 (N_12047,N_11849,N_11930);
and U12048 (N_12048,N_11881,N_11911);
nor U12049 (N_12049,N_11953,N_11932);
nor U12050 (N_12050,N_11775,N_11924);
and U12051 (N_12051,N_11952,N_11915);
nand U12052 (N_12052,N_11947,N_11877);
and U12053 (N_12053,N_11859,N_11820);
nand U12054 (N_12054,N_11935,N_11776);
and U12055 (N_12055,N_11827,N_11812);
or U12056 (N_12056,N_11781,N_11816);
or U12057 (N_12057,N_11956,N_11989);
or U12058 (N_12058,N_11760,N_11782);
xor U12059 (N_12059,N_11756,N_11899);
and U12060 (N_12060,N_11863,N_11765);
or U12061 (N_12061,N_11946,N_11754);
nand U12062 (N_12062,N_11927,N_11974);
nand U12063 (N_12063,N_11920,N_11850);
and U12064 (N_12064,N_11826,N_11780);
or U12065 (N_12065,N_11808,N_11959);
or U12066 (N_12066,N_11887,N_11784);
and U12067 (N_12067,N_11923,N_11806);
and U12068 (N_12068,N_11796,N_11857);
nor U12069 (N_12069,N_11854,N_11950);
nand U12070 (N_12070,N_11831,N_11939);
or U12071 (N_12071,N_11891,N_11818);
nor U12072 (N_12072,N_11965,N_11921);
or U12073 (N_12073,N_11976,N_11815);
nor U12074 (N_12074,N_11844,N_11908);
nand U12075 (N_12075,N_11972,N_11977);
and U12076 (N_12076,N_11814,N_11783);
nand U12077 (N_12077,N_11912,N_11799);
nand U12078 (N_12078,N_11903,N_11999);
nor U12079 (N_12079,N_11755,N_11951);
nor U12080 (N_12080,N_11805,N_11882);
nor U12081 (N_12081,N_11973,N_11750);
or U12082 (N_12082,N_11848,N_11916);
and U12083 (N_12083,N_11884,N_11880);
or U12084 (N_12084,N_11970,N_11926);
nand U12085 (N_12085,N_11770,N_11996);
or U12086 (N_12086,N_11769,N_11966);
or U12087 (N_12087,N_11994,N_11786);
nor U12088 (N_12088,N_11971,N_11858);
nor U12089 (N_12089,N_11824,N_11758);
and U12090 (N_12090,N_11942,N_11875);
nor U12091 (N_12091,N_11955,N_11777);
nor U12092 (N_12092,N_11907,N_11928);
and U12093 (N_12093,N_11793,N_11840);
xnor U12094 (N_12094,N_11787,N_11954);
and U12095 (N_12095,N_11838,N_11964);
xor U12096 (N_12096,N_11900,N_11789);
xnor U12097 (N_12097,N_11876,N_11807);
nor U12098 (N_12098,N_11752,N_11979);
nand U12099 (N_12099,N_11772,N_11864);
or U12100 (N_12100,N_11998,N_11922);
nand U12101 (N_12101,N_11792,N_11797);
nor U12102 (N_12102,N_11809,N_11983);
nand U12103 (N_12103,N_11868,N_11867);
nand U12104 (N_12104,N_11978,N_11933);
nand U12105 (N_12105,N_11757,N_11936);
or U12106 (N_12106,N_11968,N_11886);
xor U12107 (N_12107,N_11987,N_11961);
and U12108 (N_12108,N_11834,N_11901);
or U12109 (N_12109,N_11892,N_11804);
nand U12110 (N_12110,N_11761,N_11847);
and U12111 (N_12111,N_11962,N_11852);
or U12112 (N_12112,N_11819,N_11918);
nor U12113 (N_12113,N_11878,N_11821);
nand U12114 (N_12114,N_11753,N_11751);
nand U12115 (N_12115,N_11894,N_11762);
nand U12116 (N_12116,N_11986,N_11845);
nor U12117 (N_12117,N_11832,N_11895);
or U12118 (N_12118,N_11843,N_11969);
nand U12119 (N_12119,N_11768,N_11823);
or U12120 (N_12120,N_11870,N_11941);
nand U12121 (N_12121,N_11785,N_11967);
nor U12122 (N_12122,N_11985,N_11919);
nand U12123 (N_12123,N_11896,N_11943);
nor U12124 (N_12124,N_11925,N_11835);
xor U12125 (N_12125,N_11787,N_11791);
and U12126 (N_12126,N_11758,N_11822);
or U12127 (N_12127,N_11843,N_11936);
nor U12128 (N_12128,N_11936,N_11841);
and U12129 (N_12129,N_11940,N_11975);
nand U12130 (N_12130,N_11773,N_11957);
and U12131 (N_12131,N_11804,N_11965);
nand U12132 (N_12132,N_11860,N_11899);
and U12133 (N_12133,N_11922,N_11901);
and U12134 (N_12134,N_11932,N_11922);
xnor U12135 (N_12135,N_11912,N_11903);
and U12136 (N_12136,N_11778,N_11993);
and U12137 (N_12137,N_11994,N_11944);
or U12138 (N_12138,N_11893,N_11858);
nand U12139 (N_12139,N_11954,N_11893);
nand U12140 (N_12140,N_11931,N_11844);
nand U12141 (N_12141,N_11956,N_11900);
nand U12142 (N_12142,N_11844,N_11874);
or U12143 (N_12143,N_11892,N_11772);
nand U12144 (N_12144,N_11978,N_11837);
xor U12145 (N_12145,N_11848,N_11974);
xor U12146 (N_12146,N_11990,N_11826);
or U12147 (N_12147,N_11929,N_11907);
or U12148 (N_12148,N_11758,N_11795);
nand U12149 (N_12149,N_11931,N_11980);
and U12150 (N_12150,N_11958,N_11849);
xor U12151 (N_12151,N_11843,N_11950);
or U12152 (N_12152,N_11800,N_11904);
nand U12153 (N_12153,N_11998,N_11805);
and U12154 (N_12154,N_11946,N_11814);
or U12155 (N_12155,N_11973,N_11830);
nor U12156 (N_12156,N_11940,N_11869);
nand U12157 (N_12157,N_11843,N_11881);
nand U12158 (N_12158,N_11925,N_11872);
or U12159 (N_12159,N_11767,N_11884);
nor U12160 (N_12160,N_11858,N_11941);
nor U12161 (N_12161,N_11774,N_11847);
or U12162 (N_12162,N_11826,N_11870);
nand U12163 (N_12163,N_11843,N_11844);
and U12164 (N_12164,N_11972,N_11893);
or U12165 (N_12165,N_11856,N_11845);
or U12166 (N_12166,N_11905,N_11755);
nand U12167 (N_12167,N_11825,N_11976);
nand U12168 (N_12168,N_11916,N_11951);
nor U12169 (N_12169,N_11916,N_11953);
xnor U12170 (N_12170,N_11935,N_11767);
nor U12171 (N_12171,N_11961,N_11847);
xor U12172 (N_12172,N_11761,N_11864);
and U12173 (N_12173,N_11862,N_11884);
or U12174 (N_12174,N_11973,N_11976);
nand U12175 (N_12175,N_11993,N_11964);
or U12176 (N_12176,N_11927,N_11767);
or U12177 (N_12177,N_11848,N_11805);
and U12178 (N_12178,N_11981,N_11783);
or U12179 (N_12179,N_11783,N_11953);
or U12180 (N_12180,N_11891,N_11939);
nor U12181 (N_12181,N_11842,N_11847);
and U12182 (N_12182,N_11805,N_11945);
nand U12183 (N_12183,N_11794,N_11883);
and U12184 (N_12184,N_11835,N_11908);
or U12185 (N_12185,N_11789,N_11834);
and U12186 (N_12186,N_11761,N_11758);
nor U12187 (N_12187,N_11973,N_11817);
and U12188 (N_12188,N_11927,N_11840);
nand U12189 (N_12189,N_11967,N_11898);
xnor U12190 (N_12190,N_11897,N_11894);
nand U12191 (N_12191,N_11832,N_11834);
or U12192 (N_12192,N_11810,N_11963);
nor U12193 (N_12193,N_11890,N_11812);
nand U12194 (N_12194,N_11797,N_11853);
nor U12195 (N_12195,N_11972,N_11995);
nand U12196 (N_12196,N_11994,N_11843);
xor U12197 (N_12197,N_11961,N_11919);
or U12198 (N_12198,N_11920,N_11894);
nor U12199 (N_12199,N_11913,N_11783);
and U12200 (N_12200,N_11873,N_11881);
nand U12201 (N_12201,N_11862,N_11855);
nor U12202 (N_12202,N_11930,N_11859);
and U12203 (N_12203,N_11798,N_11929);
and U12204 (N_12204,N_11899,N_11770);
xor U12205 (N_12205,N_11982,N_11772);
nor U12206 (N_12206,N_11906,N_11763);
nor U12207 (N_12207,N_11787,N_11840);
or U12208 (N_12208,N_11836,N_11941);
or U12209 (N_12209,N_11978,N_11924);
nand U12210 (N_12210,N_11925,N_11973);
or U12211 (N_12211,N_11816,N_11973);
nor U12212 (N_12212,N_11844,N_11839);
nor U12213 (N_12213,N_11942,N_11787);
and U12214 (N_12214,N_11980,N_11802);
and U12215 (N_12215,N_11836,N_11800);
and U12216 (N_12216,N_11988,N_11859);
nand U12217 (N_12217,N_11768,N_11764);
xor U12218 (N_12218,N_11922,N_11950);
and U12219 (N_12219,N_11779,N_11768);
or U12220 (N_12220,N_11773,N_11907);
nand U12221 (N_12221,N_11921,N_11825);
nor U12222 (N_12222,N_11767,N_11952);
xor U12223 (N_12223,N_11899,N_11784);
and U12224 (N_12224,N_11896,N_11964);
or U12225 (N_12225,N_11972,N_11967);
and U12226 (N_12226,N_11876,N_11834);
nor U12227 (N_12227,N_11963,N_11868);
nor U12228 (N_12228,N_11984,N_11948);
nor U12229 (N_12229,N_11972,N_11872);
and U12230 (N_12230,N_11806,N_11792);
xor U12231 (N_12231,N_11997,N_11809);
and U12232 (N_12232,N_11763,N_11758);
or U12233 (N_12233,N_11909,N_11813);
or U12234 (N_12234,N_11754,N_11759);
nand U12235 (N_12235,N_11799,N_11947);
xor U12236 (N_12236,N_11805,N_11776);
nor U12237 (N_12237,N_11865,N_11801);
xnor U12238 (N_12238,N_11962,N_11899);
and U12239 (N_12239,N_11986,N_11869);
and U12240 (N_12240,N_11931,N_11781);
nor U12241 (N_12241,N_11769,N_11909);
or U12242 (N_12242,N_11830,N_11936);
and U12243 (N_12243,N_11752,N_11924);
nand U12244 (N_12244,N_11965,N_11934);
nor U12245 (N_12245,N_11878,N_11769);
nor U12246 (N_12246,N_11904,N_11862);
nor U12247 (N_12247,N_11987,N_11814);
or U12248 (N_12248,N_11903,N_11867);
nor U12249 (N_12249,N_11859,N_11945);
and U12250 (N_12250,N_12221,N_12235);
nand U12251 (N_12251,N_12214,N_12091);
or U12252 (N_12252,N_12150,N_12060);
nor U12253 (N_12253,N_12016,N_12094);
nor U12254 (N_12254,N_12172,N_12102);
xor U12255 (N_12255,N_12165,N_12058);
or U12256 (N_12256,N_12181,N_12115);
nor U12257 (N_12257,N_12128,N_12160);
and U12258 (N_12258,N_12050,N_12074);
xnor U12259 (N_12259,N_12053,N_12105);
and U12260 (N_12260,N_12122,N_12240);
nand U12261 (N_12261,N_12171,N_12180);
xnor U12262 (N_12262,N_12008,N_12145);
and U12263 (N_12263,N_12049,N_12107);
nand U12264 (N_12264,N_12238,N_12175);
nor U12265 (N_12265,N_12051,N_12021);
or U12266 (N_12266,N_12041,N_12228);
nand U12267 (N_12267,N_12029,N_12056);
xnor U12268 (N_12268,N_12007,N_12118);
xor U12269 (N_12269,N_12133,N_12210);
or U12270 (N_12270,N_12183,N_12163);
xor U12271 (N_12271,N_12218,N_12138);
or U12272 (N_12272,N_12001,N_12025);
or U12273 (N_12273,N_12002,N_12249);
nand U12274 (N_12274,N_12075,N_12103);
xnor U12275 (N_12275,N_12174,N_12045);
nor U12276 (N_12276,N_12077,N_12222);
and U12277 (N_12277,N_12042,N_12035);
or U12278 (N_12278,N_12095,N_12036);
and U12279 (N_12279,N_12113,N_12018);
nor U12280 (N_12280,N_12032,N_12028);
or U12281 (N_12281,N_12031,N_12124);
nand U12282 (N_12282,N_12213,N_12081);
xor U12283 (N_12283,N_12179,N_12186);
or U12284 (N_12284,N_12040,N_12088);
nand U12285 (N_12285,N_12038,N_12080);
nor U12286 (N_12286,N_12223,N_12151);
nor U12287 (N_12287,N_12022,N_12127);
or U12288 (N_12288,N_12026,N_12116);
xnor U12289 (N_12289,N_12166,N_12068);
nor U12290 (N_12290,N_12147,N_12247);
or U12291 (N_12291,N_12152,N_12211);
or U12292 (N_12292,N_12090,N_12108);
or U12293 (N_12293,N_12069,N_12061);
and U12294 (N_12294,N_12248,N_12059);
or U12295 (N_12295,N_12190,N_12131);
or U12296 (N_12296,N_12104,N_12157);
nand U12297 (N_12297,N_12188,N_12246);
nor U12298 (N_12298,N_12054,N_12207);
or U12299 (N_12299,N_12212,N_12197);
nand U12300 (N_12300,N_12071,N_12083);
xnor U12301 (N_12301,N_12215,N_12195);
nor U12302 (N_12302,N_12132,N_12048);
xor U12303 (N_12303,N_12010,N_12136);
or U12304 (N_12304,N_12189,N_12201);
xnor U12305 (N_12305,N_12110,N_12065);
and U12306 (N_12306,N_12027,N_12137);
nor U12307 (N_12307,N_12044,N_12226);
nor U12308 (N_12308,N_12141,N_12125);
and U12309 (N_12309,N_12158,N_12243);
nor U12310 (N_12310,N_12046,N_12084);
and U12311 (N_12311,N_12154,N_12167);
nor U12312 (N_12312,N_12164,N_12052);
nand U12313 (N_12313,N_12193,N_12097);
nor U12314 (N_12314,N_12230,N_12196);
or U12315 (N_12315,N_12209,N_12191);
nand U12316 (N_12316,N_12089,N_12194);
xnor U12317 (N_12317,N_12192,N_12078);
or U12318 (N_12318,N_12184,N_12079);
nand U12319 (N_12319,N_12009,N_12126);
nand U12320 (N_12320,N_12208,N_12015);
and U12321 (N_12321,N_12011,N_12030);
or U12322 (N_12322,N_12143,N_12047);
or U12323 (N_12323,N_12144,N_12224);
xnor U12324 (N_12324,N_12245,N_12135);
or U12325 (N_12325,N_12204,N_12233);
or U12326 (N_12326,N_12216,N_12155);
nor U12327 (N_12327,N_12123,N_12085);
and U12328 (N_12328,N_12063,N_12004);
or U12329 (N_12329,N_12006,N_12202);
or U12330 (N_12330,N_12017,N_12129);
xor U12331 (N_12331,N_12130,N_12112);
or U12332 (N_12332,N_12037,N_12064);
and U12333 (N_12333,N_12134,N_12217);
nand U12334 (N_12334,N_12225,N_12087);
or U12335 (N_12335,N_12206,N_12234);
or U12336 (N_12336,N_12176,N_12003);
or U12337 (N_12337,N_12149,N_12169);
nand U12338 (N_12338,N_12098,N_12231);
nand U12339 (N_12339,N_12055,N_12034);
and U12340 (N_12340,N_12066,N_12067);
xor U12341 (N_12341,N_12062,N_12111);
nor U12342 (N_12342,N_12073,N_12200);
or U12343 (N_12343,N_12013,N_12242);
or U12344 (N_12344,N_12148,N_12239);
and U12345 (N_12345,N_12153,N_12100);
and U12346 (N_12346,N_12082,N_12024);
and U12347 (N_12347,N_12177,N_12146);
or U12348 (N_12348,N_12241,N_12178);
or U12349 (N_12349,N_12023,N_12072);
nor U12350 (N_12350,N_12161,N_12057);
nand U12351 (N_12351,N_12117,N_12120);
nor U12352 (N_12352,N_12106,N_12092);
and U12353 (N_12353,N_12139,N_12227);
or U12354 (N_12354,N_12086,N_12244);
xor U12355 (N_12355,N_12162,N_12114);
or U12356 (N_12356,N_12205,N_12096);
nor U12357 (N_12357,N_12185,N_12142);
nor U12358 (N_12358,N_12203,N_12020);
nand U12359 (N_12359,N_12168,N_12033);
and U12360 (N_12360,N_12076,N_12159);
and U12361 (N_12361,N_12014,N_12236);
or U12362 (N_12362,N_12099,N_12000);
and U12363 (N_12363,N_12187,N_12070);
nor U12364 (N_12364,N_12119,N_12199);
or U12365 (N_12365,N_12019,N_12229);
or U12366 (N_12366,N_12173,N_12198);
or U12367 (N_12367,N_12093,N_12109);
or U12368 (N_12368,N_12012,N_12219);
or U12369 (N_12369,N_12101,N_12005);
xor U12370 (N_12370,N_12043,N_12156);
nor U12371 (N_12371,N_12170,N_12039);
or U12372 (N_12372,N_12121,N_12182);
or U12373 (N_12373,N_12237,N_12140);
and U12374 (N_12374,N_12220,N_12232);
nor U12375 (N_12375,N_12015,N_12149);
nor U12376 (N_12376,N_12069,N_12026);
nor U12377 (N_12377,N_12096,N_12155);
nor U12378 (N_12378,N_12169,N_12114);
and U12379 (N_12379,N_12052,N_12016);
and U12380 (N_12380,N_12239,N_12135);
nor U12381 (N_12381,N_12032,N_12070);
and U12382 (N_12382,N_12112,N_12174);
nor U12383 (N_12383,N_12059,N_12242);
or U12384 (N_12384,N_12075,N_12215);
and U12385 (N_12385,N_12155,N_12003);
or U12386 (N_12386,N_12041,N_12014);
and U12387 (N_12387,N_12101,N_12171);
or U12388 (N_12388,N_12038,N_12131);
nor U12389 (N_12389,N_12053,N_12083);
nand U12390 (N_12390,N_12213,N_12118);
nand U12391 (N_12391,N_12042,N_12195);
nor U12392 (N_12392,N_12013,N_12057);
or U12393 (N_12393,N_12177,N_12076);
nand U12394 (N_12394,N_12177,N_12133);
nor U12395 (N_12395,N_12067,N_12034);
nand U12396 (N_12396,N_12017,N_12201);
nor U12397 (N_12397,N_12206,N_12195);
and U12398 (N_12398,N_12166,N_12121);
and U12399 (N_12399,N_12182,N_12036);
and U12400 (N_12400,N_12054,N_12227);
or U12401 (N_12401,N_12100,N_12006);
or U12402 (N_12402,N_12223,N_12237);
or U12403 (N_12403,N_12130,N_12148);
nand U12404 (N_12404,N_12079,N_12226);
nand U12405 (N_12405,N_12203,N_12194);
nor U12406 (N_12406,N_12198,N_12131);
nor U12407 (N_12407,N_12008,N_12096);
or U12408 (N_12408,N_12042,N_12161);
nand U12409 (N_12409,N_12088,N_12219);
and U12410 (N_12410,N_12132,N_12094);
nor U12411 (N_12411,N_12139,N_12195);
or U12412 (N_12412,N_12021,N_12243);
nor U12413 (N_12413,N_12148,N_12199);
nor U12414 (N_12414,N_12055,N_12008);
and U12415 (N_12415,N_12248,N_12160);
or U12416 (N_12416,N_12123,N_12022);
and U12417 (N_12417,N_12007,N_12073);
and U12418 (N_12418,N_12049,N_12008);
nand U12419 (N_12419,N_12191,N_12199);
or U12420 (N_12420,N_12000,N_12024);
nand U12421 (N_12421,N_12017,N_12090);
nor U12422 (N_12422,N_12148,N_12048);
nor U12423 (N_12423,N_12032,N_12122);
nand U12424 (N_12424,N_12132,N_12170);
nand U12425 (N_12425,N_12231,N_12225);
nor U12426 (N_12426,N_12048,N_12216);
and U12427 (N_12427,N_12028,N_12086);
or U12428 (N_12428,N_12021,N_12210);
nor U12429 (N_12429,N_12227,N_12046);
or U12430 (N_12430,N_12163,N_12153);
nand U12431 (N_12431,N_12137,N_12059);
nor U12432 (N_12432,N_12203,N_12113);
or U12433 (N_12433,N_12222,N_12083);
and U12434 (N_12434,N_12187,N_12051);
nand U12435 (N_12435,N_12218,N_12111);
or U12436 (N_12436,N_12086,N_12227);
or U12437 (N_12437,N_12205,N_12004);
nand U12438 (N_12438,N_12171,N_12043);
nor U12439 (N_12439,N_12061,N_12003);
nor U12440 (N_12440,N_12075,N_12158);
or U12441 (N_12441,N_12153,N_12039);
xor U12442 (N_12442,N_12200,N_12117);
nand U12443 (N_12443,N_12051,N_12072);
or U12444 (N_12444,N_12177,N_12088);
nor U12445 (N_12445,N_12037,N_12143);
nor U12446 (N_12446,N_12244,N_12047);
nor U12447 (N_12447,N_12093,N_12035);
or U12448 (N_12448,N_12089,N_12021);
or U12449 (N_12449,N_12041,N_12100);
nor U12450 (N_12450,N_12171,N_12036);
nor U12451 (N_12451,N_12187,N_12193);
nor U12452 (N_12452,N_12144,N_12037);
nor U12453 (N_12453,N_12235,N_12244);
nand U12454 (N_12454,N_12132,N_12019);
nand U12455 (N_12455,N_12143,N_12011);
nor U12456 (N_12456,N_12208,N_12229);
or U12457 (N_12457,N_12057,N_12131);
and U12458 (N_12458,N_12224,N_12239);
nor U12459 (N_12459,N_12194,N_12222);
or U12460 (N_12460,N_12210,N_12073);
or U12461 (N_12461,N_12207,N_12063);
or U12462 (N_12462,N_12150,N_12039);
xnor U12463 (N_12463,N_12045,N_12186);
and U12464 (N_12464,N_12246,N_12076);
nand U12465 (N_12465,N_12102,N_12095);
nand U12466 (N_12466,N_12244,N_12139);
or U12467 (N_12467,N_12043,N_12222);
xor U12468 (N_12468,N_12055,N_12214);
nand U12469 (N_12469,N_12025,N_12008);
or U12470 (N_12470,N_12132,N_12161);
nor U12471 (N_12471,N_12206,N_12101);
or U12472 (N_12472,N_12043,N_12135);
nand U12473 (N_12473,N_12183,N_12241);
nand U12474 (N_12474,N_12248,N_12177);
nand U12475 (N_12475,N_12020,N_12243);
or U12476 (N_12476,N_12224,N_12031);
nor U12477 (N_12477,N_12082,N_12085);
nor U12478 (N_12478,N_12022,N_12103);
nand U12479 (N_12479,N_12019,N_12183);
nor U12480 (N_12480,N_12192,N_12242);
nand U12481 (N_12481,N_12218,N_12210);
and U12482 (N_12482,N_12112,N_12116);
nor U12483 (N_12483,N_12048,N_12007);
or U12484 (N_12484,N_12152,N_12104);
nor U12485 (N_12485,N_12240,N_12089);
nand U12486 (N_12486,N_12012,N_12177);
and U12487 (N_12487,N_12146,N_12244);
nor U12488 (N_12488,N_12051,N_12058);
nor U12489 (N_12489,N_12188,N_12215);
nor U12490 (N_12490,N_12231,N_12028);
and U12491 (N_12491,N_12064,N_12077);
nand U12492 (N_12492,N_12008,N_12136);
or U12493 (N_12493,N_12228,N_12024);
xnor U12494 (N_12494,N_12171,N_12081);
or U12495 (N_12495,N_12030,N_12081);
xnor U12496 (N_12496,N_12141,N_12043);
nand U12497 (N_12497,N_12030,N_12104);
nor U12498 (N_12498,N_12052,N_12179);
nor U12499 (N_12499,N_12065,N_12202);
and U12500 (N_12500,N_12383,N_12398);
or U12501 (N_12501,N_12361,N_12410);
nor U12502 (N_12502,N_12308,N_12314);
nor U12503 (N_12503,N_12342,N_12389);
and U12504 (N_12504,N_12441,N_12403);
and U12505 (N_12505,N_12268,N_12411);
or U12506 (N_12506,N_12254,N_12488);
or U12507 (N_12507,N_12307,N_12365);
xnor U12508 (N_12508,N_12256,N_12315);
nor U12509 (N_12509,N_12323,N_12355);
nor U12510 (N_12510,N_12435,N_12421);
nor U12511 (N_12511,N_12391,N_12294);
nor U12512 (N_12512,N_12362,N_12352);
nor U12513 (N_12513,N_12266,N_12485);
nor U12514 (N_12514,N_12311,N_12261);
nor U12515 (N_12515,N_12399,N_12340);
xor U12516 (N_12516,N_12334,N_12487);
nand U12517 (N_12517,N_12439,N_12369);
nor U12518 (N_12518,N_12394,N_12446);
or U12519 (N_12519,N_12289,N_12499);
nand U12520 (N_12520,N_12346,N_12466);
nor U12521 (N_12521,N_12449,N_12364);
and U12522 (N_12522,N_12276,N_12288);
nand U12523 (N_12523,N_12408,N_12468);
nand U12524 (N_12524,N_12335,N_12444);
and U12525 (N_12525,N_12345,N_12448);
and U12526 (N_12526,N_12430,N_12453);
nand U12527 (N_12527,N_12416,N_12328);
and U12528 (N_12528,N_12472,N_12393);
xnor U12529 (N_12529,N_12338,N_12324);
nor U12530 (N_12530,N_12486,N_12373);
or U12531 (N_12531,N_12400,N_12291);
or U12532 (N_12532,N_12458,N_12258);
or U12533 (N_12533,N_12343,N_12437);
and U12534 (N_12534,N_12490,N_12496);
or U12535 (N_12535,N_12303,N_12427);
nor U12536 (N_12536,N_12379,N_12385);
or U12537 (N_12537,N_12321,N_12269);
xnor U12538 (N_12538,N_12319,N_12498);
nand U12539 (N_12539,N_12406,N_12341);
or U12540 (N_12540,N_12386,N_12360);
xnor U12541 (N_12541,N_12283,N_12265);
nor U12542 (N_12542,N_12442,N_12368);
nor U12543 (N_12543,N_12380,N_12257);
or U12544 (N_12544,N_12409,N_12372);
nor U12545 (N_12545,N_12282,N_12378);
and U12546 (N_12546,N_12418,N_12279);
nor U12547 (N_12547,N_12290,N_12310);
and U12548 (N_12548,N_12447,N_12425);
and U12549 (N_12549,N_12339,N_12297);
nand U12550 (N_12550,N_12489,N_12274);
nand U12551 (N_12551,N_12417,N_12415);
or U12552 (N_12552,N_12358,N_12312);
or U12553 (N_12553,N_12454,N_12428);
and U12554 (N_12554,N_12464,N_12250);
or U12555 (N_12555,N_12267,N_12337);
nor U12556 (N_12556,N_12484,N_12359);
or U12557 (N_12557,N_12434,N_12493);
nand U12558 (N_12558,N_12285,N_12480);
and U12559 (N_12559,N_12262,N_12420);
nand U12560 (N_12560,N_12419,N_12405);
and U12561 (N_12561,N_12348,N_12280);
nand U12562 (N_12562,N_12473,N_12450);
or U12563 (N_12563,N_12443,N_12465);
or U12564 (N_12564,N_12251,N_12366);
or U12565 (N_12565,N_12327,N_12374);
or U12566 (N_12566,N_12281,N_12482);
xor U12567 (N_12567,N_12371,N_12470);
nor U12568 (N_12568,N_12357,N_12436);
nand U12569 (N_12569,N_12356,N_12497);
xnor U12570 (N_12570,N_12286,N_12476);
nor U12571 (N_12571,N_12271,N_12301);
and U12572 (N_12572,N_12325,N_12332);
nand U12573 (N_12573,N_12309,N_12330);
and U12574 (N_12574,N_12467,N_12349);
nor U12575 (N_12575,N_12494,N_12431);
or U12576 (N_12576,N_12384,N_12333);
or U12577 (N_12577,N_12397,N_12272);
and U12578 (N_12578,N_12295,N_12304);
nand U12579 (N_12579,N_12392,N_12396);
nand U12580 (N_12580,N_12459,N_12376);
and U12581 (N_12581,N_12463,N_12273);
and U12582 (N_12582,N_12481,N_12255);
or U12583 (N_12583,N_12375,N_12433);
xnor U12584 (N_12584,N_12306,N_12456);
xor U12585 (N_12585,N_12460,N_12370);
nand U12586 (N_12586,N_12347,N_12452);
nor U12587 (N_12587,N_12432,N_12275);
or U12588 (N_12588,N_12412,N_12475);
nor U12589 (N_12589,N_12302,N_12351);
xor U12590 (N_12590,N_12426,N_12483);
nand U12591 (N_12591,N_12377,N_12445);
or U12592 (N_12592,N_12331,N_12264);
and U12593 (N_12593,N_12317,N_12451);
nor U12594 (N_12594,N_12471,N_12353);
xor U12595 (N_12595,N_12401,N_12495);
xnor U12596 (N_12596,N_12424,N_12455);
and U12597 (N_12597,N_12423,N_12479);
or U12598 (N_12598,N_12322,N_12320);
nand U12599 (N_12599,N_12491,N_12253);
nor U12600 (N_12600,N_12284,N_12382);
or U12601 (N_12601,N_12296,N_12422);
and U12602 (N_12602,N_12492,N_12277);
or U12603 (N_12603,N_12407,N_12429);
and U12604 (N_12604,N_12263,N_12300);
nor U12605 (N_12605,N_12318,N_12478);
nor U12606 (N_12606,N_12278,N_12367);
nor U12607 (N_12607,N_12413,N_12387);
nand U12608 (N_12608,N_12313,N_12299);
and U12609 (N_12609,N_12404,N_12316);
xnor U12610 (N_12610,N_12402,N_12388);
nand U12611 (N_12611,N_12326,N_12252);
and U12612 (N_12612,N_12461,N_12293);
or U12613 (N_12613,N_12440,N_12395);
and U12614 (N_12614,N_12292,N_12469);
xnor U12615 (N_12615,N_12298,N_12477);
nor U12616 (N_12616,N_12260,N_12354);
nor U12617 (N_12617,N_12381,N_12305);
and U12618 (N_12618,N_12414,N_12390);
nand U12619 (N_12619,N_12438,N_12259);
or U12620 (N_12620,N_12344,N_12350);
or U12621 (N_12621,N_12270,N_12363);
and U12622 (N_12622,N_12462,N_12287);
nor U12623 (N_12623,N_12336,N_12457);
or U12624 (N_12624,N_12474,N_12329);
and U12625 (N_12625,N_12470,N_12282);
and U12626 (N_12626,N_12286,N_12256);
or U12627 (N_12627,N_12320,N_12294);
nor U12628 (N_12628,N_12351,N_12424);
nor U12629 (N_12629,N_12275,N_12374);
nor U12630 (N_12630,N_12251,N_12319);
nor U12631 (N_12631,N_12388,N_12335);
or U12632 (N_12632,N_12353,N_12386);
or U12633 (N_12633,N_12332,N_12286);
or U12634 (N_12634,N_12406,N_12451);
and U12635 (N_12635,N_12269,N_12481);
nand U12636 (N_12636,N_12425,N_12304);
nand U12637 (N_12637,N_12392,N_12366);
nor U12638 (N_12638,N_12314,N_12397);
nor U12639 (N_12639,N_12374,N_12298);
nand U12640 (N_12640,N_12399,N_12314);
and U12641 (N_12641,N_12296,N_12414);
and U12642 (N_12642,N_12251,N_12362);
xor U12643 (N_12643,N_12357,N_12483);
nand U12644 (N_12644,N_12339,N_12420);
or U12645 (N_12645,N_12325,N_12337);
or U12646 (N_12646,N_12351,N_12393);
nor U12647 (N_12647,N_12280,N_12350);
nand U12648 (N_12648,N_12320,N_12376);
nand U12649 (N_12649,N_12347,N_12370);
or U12650 (N_12650,N_12383,N_12310);
nand U12651 (N_12651,N_12455,N_12262);
or U12652 (N_12652,N_12369,N_12370);
nand U12653 (N_12653,N_12362,N_12471);
or U12654 (N_12654,N_12429,N_12440);
nand U12655 (N_12655,N_12283,N_12466);
nand U12656 (N_12656,N_12488,N_12422);
or U12657 (N_12657,N_12289,N_12265);
and U12658 (N_12658,N_12353,N_12305);
nand U12659 (N_12659,N_12485,N_12383);
and U12660 (N_12660,N_12348,N_12443);
nand U12661 (N_12661,N_12310,N_12379);
or U12662 (N_12662,N_12332,N_12363);
nor U12663 (N_12663,N_12424,N_12482);
nor U12664 (N_12664,N_12387,N_12428);
or U12665 (N_12665,N_12498,N_12466);
and U12666 (N_12666,N_12272,N_12474);
nand U12667 (N_12667,N_12293,N_12443);
or U12668 (N_12668,N_12354,N_12338);
nand U12669 (N_12669,N_12499,N_12381);
nand U12670 (N_12670,N_12363,N_12464);
nand U12671 (N_12671,N_12439,N_12334);
and U12672 (N_12672,N_12373,N_12435);
or U12673 (N_12673,N_12326,N_12253);
nor U12674 (N_12674,N_12351,N_12263);
or U12675 (N_12675,N_12465,N_12354);
nor U12676 (N_12676,N_12430,N_12339);
nor U12677 (N_12677,N_12479,N_12275);
and U12678 (N_12678,N_12380,N_12291);
and U12679 (N_12679,N_12448,N_12481);
or U12680 (N_12680,N_12446,N_12261);
nor U12681 (N_12681,N_12252,N_12419);
or U12682 (N_12682,N_12361,N_12481);
and U12683 (N_12683,N_12432,N_12476);
nor U12684 (N_12684,N_12394,N_12349);
or U12685 (N_12685,N_12338,N_12491);
nand U12686 (N_12686,N_12292,N_12495);
or U12687 (N_12687,N_12344,N_12464);
nand U12688 (N_12688,N_12346,N_12471);
nand U12689 (N_12689,N_12395,N_12333);
or U12690 (N_12690,N_12482,N_12382);
or U12691 (N_12691,N_12356,N_12416);
or U12692 (N_12692,N_12465,N_12399);
or U12693 (N_12693,N_12351,N_12391);
and U12694 (N_12694,N_12476,N_12371);
or U12695 (N_12695,N_12322,N_12343);
nor U12696 (N_12696,N_12460,N_12278);
and U12697 (N_12697,N_12433,N_12485);
or U12698 (N_12698,N_12341,N_12376);
or U12699 (N_12699,N_12318,N_12432);
nor U12700 (N_12700,N_12392,N_12479);
xor U12701 (N_12701,N_12387,N_12395);
or U12702 (N_12702,N_12447,N_12379);
nor U12703 (N_12703,N_12260,N_12370);
xor U12704 (N_12704,N_12449,N_12354);
nor U12705 (N_12705,N_12284,N_12469);
or U12706 (N_12706,N_12364,N_12251);
and U12707 (N_12707,N_12385,N_12455);
or U12708 (N_12708,N_12284,N_12436);
or U12709 (N_12709,N_12351,N_12352);
nor U12710 (N_12710,N_12312,N_12378);
nor U12711 (N_12711,N_12352,N_12430);
nand U12712 (N_12712,N_12391,N_12381);
nor U12713 (N_12713,N_12357,N_12333);
nor U12714 (N_12714,N_12497,N_12423);
or U12715 (N_12715,N_12446,N_12360);
nor U12716 (N_12716,N_12295,N_12255);
and U12717 (N_12717,N_12272,N_12305);
or U12718 (N_12718,N_12327,N_12322);
nand U12719 (N_12719,N_12424,N_12464);
nor U12720 (N_12720,N_12479,N_12456);
nor U12721 (N_12721,N_12316,N_12474);
xnor U12722 (N_12722,N_12432,N_12384);
and U12723 (N_12723,N_12403,N_12404);
nand U12724 (N_12724,N_12265,N_12401);
and U12725 (N_12725,N_12351,N_12250);
and U12726 (N_12726,N_12446,N_12469);
nand U12727 (N_12727,N_12399,N_12369);
or U12728 (N_12728,N_12293,N_12470);
nand U12729 (N_12729,N_12455,N_12329);
nand U12730 (N_12730,N_12324,N_12442);
xnor U12731 (N_12731,N_12354,N_12473);
and U12732 (N_12732,N_12422,N_12453);
xor U12733 (N_12733,N_12268,N_12478);
nor U12734 (N_12734,N_12407,N_12267);
xor U12735 (N_12735,N_12357,N_12287);
nand U12736 (N_12736,N_12480,N_12412);
nand U12737 (N_12737,N_12473,N_12416);
nor U12738 (N_12738,N_12290,N_12432);
nor U12739 (N_12739,N_12385,N_12423);
and U12740 (N_12740,N_12289,N_12331);
and U12741 (N_12741,N_12480,N_12297);
nor U12742 (N_12742,N_12388,N_12350);
and U12743 (N_12743,N_12496,N_12451);
xnor U12744 (N_12744,N_12413,N_12300);
and U12745 (N_12745,N_12446,N_12370);
or U12746 (N_12746,N_12446,N_12353);
nor U12747 (N_12747,N_12420,N_12457);
xnor U12748 (N_12748,N_12464,N_12443);
or U12749 (N_12749,N_12312,N_12399);
nand U12750 (N_12750,N_12707,N_12696);
or U12751 (N_12751,N_12511,N_12575);
or U12752 (N_12752,N_12676,N_12527);
and U12753 (N_12753,N_12641,N_12704);
or U12754 (N_12754,N_12669,N_12556);
nor U12755 (N_12755,N_12686,N_12591);
nand U12756 (N_12756,N_12744,N_12725);
and U12757 (N_12757,N_12507,N_12694);
or U12758 (N_12758,N_12630,N_12510);
nand U12759 (N_12759,N_12623,N_12710);
and U12760 (N_12760,N_12682,N_12528);
nand U12761 (N_12761,N_12701,N_12746);
nand U12762 (N_12762,N_12632,N_12554);
nand U12763 (N_12763,N_12559,N_12541);
or U12764 (N_12764,N_12693,N_12702);
nand U12765 (N_12765,N_12628,N_12708);
and U12766 (N_12766,N_12520,N_12657);
or U12767 (N_12767,N_12537,N_12736);
and U12768 (N_12768,N_12618,N_12664);
nor U12769 (N_12769,N_12519,N_12599);
or U12770 (N_12770,N_12579,N_12561);
nand U12771 (N_12771,N_12550,N_12518);
nor U12772 (N_12772,N_12622,N_12563);
nand U12773 (N_12773,N_12582,N_12670);
nor U12774 (N_12774,N_12601,N_12724);
or U12775 (N_12775,N_12516,N_12723);
nor U12776 (N_12776,N_12648,N_12583);
or U12777 (N_12777,N_12740,N_12592);
nor U12778 (N_12778,N_12739,N_12692);
xor U12779 (N_12779,N_12674,N_12569);
or U12780 (N_12780,N_12726,N_12580);
or U12781 (N_12781,N_12689,N_12524);
xnor U12782 (N_12782,N_12566,N_12568);
nand U12783 (N_12783,N_12544,N_12607);
nor U12784 (N_12784,N_12522,N_12699);
and U12785 (N_12785,N_12558,N_12646);
nand U12786 (N_12786,N_12578,N_12735);
and U12787 (N_12787,N_12645,N_12548);
nand U12788 (N_12788,N_12517,N_12616);
nor U12789 (N_12789,N_12668,N_12508);
or U12790 (N_12790,N_12617,N_12546);
or U12791 (N_12791,N_12504,N_12594);
xnor U12792 (N_12792,N_12531,N_12593);
xor U12793 (N_12793,N_12747,N_12659);
nor U12794 (N_12794,N_12529,N_12712);
nor U12795 (N_12795,N_12613,N_12612);
nand U12796 (N_12796,N_12715,N_12631);
and U12797 (N_12797,N_12545,N_12567);
and U12798 (N_12798,N_12539,N_12691);
or U12799 (N_12799,N_12738,N_12643);
or U12800 (N_12800,N_12625,N_12698);
nor U12801 (N_12801,N_12653,N_12502);
and U12802 (N_12802,N_12637,N_12614);
xor U12803 (N_12803,N_12671,N_12611);
or U12804 (N_12804,N_12733,N_12576);
xor U12805 (N_12805,N_12737,N_12722);
nand U12806 (N_12806,N_12572,N_12705);
nand U12807 (N_12807,N_12655,N_12596);
and U12808 (N_12808,N_12602,N_12680);
or U12809 (N_12809,N_12512,N_12662);
nand U12810 (N_12810,N_12562,N_12719);
and U12811 (N_12811,N_12731,N_12703);
nor U12812 (N_12812,N_12711,N_12642);
nand U12813 (N_12813,N_12714,N_12577);
and U12814 (N_12814,N_12745,N_12585);
and U12815 (N_12815,N_12672,N_12748);
or U12816 (N_12816,N_12581,N_12564);
or U12817 (N_12817,N_12673,N_12649);
and U12818 (N_12818,N_12526,N_12521);
or U12819 (N_12819,N_12535,N_12729);
nand U12820 (N_12820,N_12685,N_12660);
xnor U12821 (N_12821,N_12678,N_12640);
nand U12822 (N_12822,N_12652,N_12589);
or U12823 (N_12823,N_12633,N_12624);
xor U12824 (N_12824,N_12536,N_12675);
nor U12825 (N_12825,N_12540,N_12684);
nor U12826 (N_12826,N_12718,N_12565);
and U12827 (N_12827,N_12663,N_12634);
and U12828 (N_12828,N_12621,N_12650);
and U12829 (N_12829,N_12721,N_12629);
xor U12830 (N_12830,N_12555,N_12501);
or U12831 (N_12831,N_12690,N_12500);
nand U12832 (N_12832,N_12584,N_12620);
or U12833 (N_12833,N_12627,N_12534);
nor U12834 (N_12834,N_12709,N_12720);
nand U12835 (N_12835,N_12727,N_12598);
nor U12836 (N_12836,N_12551,N_12588);
and U12837 (N_12837,N_12547,N_12728);
and U12838 (N_12838,N_12635,N_12717);
or U12839 (N_12839,N_12542,N_12654);
xnor U12840 (N_12840,N_12570,N_12647);
and U12841 (N_12841,N_12679,N_12557);
nand U12842 (N_12842,N_12741,N_12687);
nor U12843 (N_12843,N_12626,N_12665);
nor U12844 (N_12844,N_12523,N_12514);
and U12845 (N_12845,N_12560,N_12608);
xor U12846 (N_12846,N_12749,N_12609);
nor U12847 (N_12847,N_12734,N_12677);
and U12848 (N_12848,N_12573,N_12636);
nor U12849 (N_12849,N_12615,N_12590);
or U12850 (N_12850,N_12700,N_12553);
xnor U12851 (N_12851,N_12730,N_12658);
nand U12852 (N_12852,N_12538,N_12595);
and U12853 (N_12853,N_12532,N_12549);
xor U12854 (N_12854,N_12605,N_12587);
nand U12855 (N_12855,N_12530,N_12552);
and U12856 (N_12856,N_12656,N_12533);
nor U12857 (N_12857,N_12666,N_12515);
and U12858 (N_12858,N_12713,N_12505);
nor U12859 (N_12859,N_12697,N_12574);
xor U12860 (N_12860,N_12597,N_12716);
nand U12861 (N_12861,N_12509,N_12603);
nor U12862 (N_12862,N_12661,N_12651);
and U12863 (N_12863,N_12606,N_12619);
nand U12864 (N_12864,N_12543,N_12706);
nor U12865 (N_12865,N_12742,N_12681);
and U12866 (N_12866,N_12688,N_12683);
nor U12867 (N_12867,N_12525,N_12667);
or U12868 (N_12868,N_12506,N_12513);
or U12869 (N_12869,N_12639,N_12610);
nor U12870 (N_12870,N_12695,N_12604);
xnor U12871 (N_12871,N_12503,N_12586);
or U12872 (N_12872,N_12743,N_12644);
and U12873 (N_12873,N_12732,N_12638);
or U12874 (N_12874,N_12600,N_12571);
or U12875 (N_12875,N_12517,N_12558);
and U12876 (N_12876,N_12742,N_12749);
or U12877 (N_12877,N_12729,N_12603);
or U12878 (N_12878,N_12685,N_12590);
nand U12879 (N_12879,N_12743,N_12669);
or U12880 (N_12880,N_12707,N_12512);
or U12881 (N_12881,N_12734,N_12669);
nand U12882 (N_12882,N_12725,N_12674);
nor U12883 (N_12883,N_12503,N_12664);
and U12884 (N_12884,N_12726,N_12591);
nor U12885 (N_12885,N_12563,N_12541);
xnor U12886 (N_12886,N_12690,N_12646);
nor U12887 (N_12887,N_12642,N_12621);
xor U12888 (N_12888,N_12546,N_12611);
or U12889 (N_12889,N_12679,N_12682);
xor U12890 (N_12890,N_12597,N_12675);
xor U12891 (N_12891,N_12541,N_12640);
and U12892 (N_12892,N_12744,N_12718);
nor U12893 (N_12893,N_12575,N_12611);
nor U12894 (N_12894,N_12616,N_12579);
xor U12895 (N_12895,N_12528,N_12742);
and U12896 (N_12896,N_12711,N_12539);
xnor U12897 (N_12897,N_12504,N_12738);
nor U12898 (N_12898,N_12542,N_12522);
or U12899 (N_12899,N_12621,N_12584);
or U12900 (N_12900,N_12723,N_12581);
xnor U12901 (N_12901,N_12556,N_12648);
nor U12902 (N_12902,N_12574,N_12618);
xor U12903 (N_12903,N_12581,N_12714);
nor U12904 (N_12904,N_12673,N_12641);
and U12905 (N_12905,N_12678,N_12689);
nand U12906 (N_12906,N_12615,N_12685);
or U12907 (N_12907,N_12629,N_12569);
nor U12908 (N_12908,N_12622,N_12533);
and U12909 (N_12909,N_12617,N_12659);
nor U12910 (N_12910,N_12727,N_12522);
nor U12911 (N_12911,N_12514,N_12621);
and U12912 (N_12912,N_12670,N_12569);
nand U12913 (N_12913,N_12582,N_12608);
or U12914 (N_12914,N_12632,N_12716);
or U12915 (N_12915,N_12651,N_12531);
and U12916 (N_12916,N_12595,N_12521);
nand U12917 (N_12917,N_12551,N_12539);
nor U12918 (N_12918,N_12507,N_12719);
or U12919 (N_12919,N_12631,N_12602);
nand U12920 (N_12920,N_12504,N_12505);
nand U12921 (N_12921,N_12553,N_12748);
and U12922 (N_12922,N_12665,N_12534);
or U12923 (N_12923,N_12605,N_12727);
or U12924 (N_12924,N_12522,N_12583);
nor U12925 (N_12925,N_12519,N_12605);
xnor U12926 (N_12926,N_12661,N_12735);
or U12927 (N_12927,N_12609,N_12510);
or U12928 (N_12928,N_12711,N_12738);
or U12929 (N_12929,N_12513,N_12700);
or U12930 (N_12930,N_12586,N_12614);
nand U12931 (N_12931,N_12548,N_12564);
and U12932 (N_12932,N_12721,N_12637);
or U12933 (N_12933,N_12626,N_12537);
or U12934 (N_12934,N_12506,N_12544);
nand U12935 (N_12935,N_12572,N_12546);
nand U12936 (N_12936,N_12578,N_12731);
nor U12937 (N_12937,N_12728,N_12607);
nand U12938 (N_12938,N_12549,N_12508);
and U12939 (N_12939,N_12740,N_12670);
nor U12940 (N_12940,N_12637,N_12590);
or U12941 (N_12941,N_12745,N_12557);
or U12942 (N_12942,N_12626,N_12728);
nand U12943 (N_12943,N_12631,N_12644);
or U12944 (N_12944,N_12668,N_12500);
and U12945 (N_12945,N_12631,N_12619);
or U12946 (N_12946,N_12626,N_12647);
or U12947 (N_12947,N_12747,N_12506);
or U12948 (N_12948,N_12719,N_12608);
nor U12949 (N_12949,N_12694,N_12731);
nor U12950 (N_12950,N_12718,N_12649);
nand U12951 (N_12951,N_12695,N_12728);
and U12952 (N_12952,N_12545,N_12594);
xnor U12953 (N_12953,N_12572,N_12505);
or U12954 (N_12954,N_12748,N_12720);
or U12955 (N_12955,N_12555,N_12629);
nand U12956 (N_12956,N_12545,N_12654);
nor U12957 (N_12957,N_12652,N_12505);
nor U12958 (N_12958,N_12679,N_12717);
nand U12959 (N_12959,N_12673,N_12595);
or U12960 (N_12960,N_12581,N_12605);
nand U12961 (N_12961,N_12671,N_12577);
nand U12962 (N_12962,N_12515,N_12536);
or U12963 (N_12963,N_12718,N_12652);
nand U12964 (N_12964,N_12601,N_12547);
nor U12965 (N_12965,N_12685,N_12728);
or U12966 (N_12966,N_12600,N_12586);
xor U12967 (N_12967,N_12626,N_12614);
xnor U12968 (N_12968,N_12665,N_12509);
nor U12969 (N_12969,N_12508,N_12548);
nand U12970 (N_12970,N_12613,N_12608);
nor U12971 (N_12971,N_12577,N_12545);
and U12972 (N_12972,N_12591,N_12508);
nand U12973 (N_12973,N_12706,N_12617);
nor U12974 (N_12974,N_12524,N_12677);
or U12975 (N_12975,N_12629,N_12653);
nor U12976 (N_12976,N_12640,N_12595);
or U12977 (N_12977,N_12729,N_12631);
nor U12978 (N_12978,N_12679,N_12675);
or U12979 (N_12979,N_12684,N_12630);
or U12980 (N_12980,N_12658,N_12731);
nand U12981 (N_12981,N_12708,N_12654);
nand U12982 (N_12982,N_12602,N_12555);
and U12983 (N_12983,N_12667,N_12664);
nor U12984 (N_12984,N_12644,N_12653);
nor U12985 (N_12985,N_12702,N_12704);
nor U12986 (N_12986,N_12740,N_12565);
and U12987 (N_12987,N_12501,N_12672);
and U12988 (N_12988,N_12663,N_12652);
and U12989 (N_12989,N_12722,N_12513);
or U12990 (N_12990,N_12741,N_12562);
and U12991 (N_12991,N_12552,N_12508);
xor U12992 (N_12992,N_12634,N_12545);
and U12993 (N_12993,N_12647,N_12602);
nand U12994 (N_12994,N_12748,N_12516);
xnor U12995 (N_12995,N_12553,N_12665);
nor U12996 (N_12996,N_12610,N_12516);
or U12997 (N_12997,N_12732,N_12670);
xor U12998 (N_12998,N_12718,N_12538);
nor U12999 (N_12999,N_12549,N_12719);
and U13000 (N_13000,N_12882,N_12900);
nor U13001 (N_13001,N_12974,N_12935);
and U13002 (N_13002,N_12881,N_12993);
and U13003 (N_13003,N_12962,N_12978);
nor U13004 (N_13004,N_12893,N_12791);
nand U13005 (N_13005,N_12856,N_12906);
nand U13006 (N_13006,N_12909,N_12777);
and U13007 (N_13007,N_12865,N_12968);
nand U13008 (N_13008,N_12901,N_12822);
nor U13009 (N_13009,N_12982,N_12778);
or U13010 (N_13010,N_12789,N_12939);
or U13011 (N_13011,N_12927,N_12899);
and U13012 (N_13012,N_12798,N_12894);
nand U13013 (N_13013,N_12889,N_12902);
nand U13014 (N_13014,N_12815,N_12760);
or U13015 (N_13015,N_12945,N_12776);
nor U13016 (N_13016,N_12753,N_12774);
xnor U13017 (N_13017,N_12884,N_12771);
nand U13018 (N_13018,N_12885,N_12796);
nor U13019 (N_13019,N_12892,N_12792);
nand U13020 (N_13020,N_12840,N_12886);
and U13021 (N_13021,N_12763,N_12952);
nor U13022 (N_13022,N_12977,N_12936);
and U13023 (N_13023,N_12752,N_12836);
nor U13024 (N_13024,N_12869,N_12844);
and U13025 (N_13025,N_12960,N_12929);
nor U13026 (N_13026,N_12958,N_12898);
nand U13027 (N_13027,N_12756,N_12891);
nand U13028 (N_13028,N_12808,N_12827);
and U13029 (N_13029,N_12975,N_12852);
nand U13030 (N_13030,N_12970,N_12768);
nor U13031 (N_13031,N_12911,N_12951);
or U13032 (N_13032,N_12766,N_12941);
or U13033 (N_13033,N_12956,N_12913);
xnor U13034 (N_13034,N_12924,N_12751);
nand U13035 (N_13035,N_12821,N_12839);
nand U13036 (N_13036,N_12938,N_12866);
nand U13037 (N_13037,N_12969,N_12834);
nor U13038 (N_13038,N_12876,N_12971);
or U13039 (N_13039,N_12787,N_12918);
nand U13040 (N_13040,N_12942,N_12785);
and U13041 (N_13041,N_12795,N_12926);
or U13042 (N_13042,N_12813,N_12930);
or U13043 (N_13043,N_12861,N_12803);
and U13044 (N_13044,N_12950,N_12843);
xnor U13045 (N_13045,N_12878,N_12880);
xnor U13046 (N_13046,N_12954,N_12860);
and U13047 (N_13047,N_12987,N_12758);
or U13048 (N_13048,N_12804,N_12750);
or U13049 (N_13049,N_12805,N_12767);
nand U13050 (N_13050,N_12830,N_12967);
nor U13051 (N_13051,N_12863,N_12986);
nor U13052 (N_13052,N_12985,N_12921);
xnor U13053 (N_13053,N_12991,N_12990);
nand U13054 (N_13054,N_12794,N_12838);
or U13055 (N_13055,N_12928,N_12849);
nor U13056 (N_13056,N_12995,N_12997);
nand U13057 (N_13057,N_12769,N_12920);
nand U13058 (N_13058,N_12932,N_12961);
xor U13059 (N_13059,N_12980,N_12999);
nor U13060 (N_13060,N_12829,N_12887);
nor U13061 (N_13061,N_12755,N_12896);
nor U13062 (N_13062,N_12915,N_12841);
nand U13063 (N_13063,N_12850,N_12966);
nand U13064 (N_13064,N_12957,N_12964);
nor U13065 (N_13065,N_12855,N_12802);
and U13066 (N_13066,N_12761,N_12870);
nor U13067 (N_13067,N_12790,N_12875);
nand U13068 (N_13068,N_12972,N_12989);
nand U13069 (N_13069,N_12871,N_12937);
nand U13070 (N_13070,N_12811,N_12963);
nand U13071 (N_13071,N_12879,N_12888);
nor U13072 (N_13072,N_12994,N_12933);
xor U13073 (N_13073,N_12917,N_12782);
nor U13074 (N_13074,N_12773,N_12903);
and U13075 (N_13075,N_12890,N_12818);
nor U13076 (N_13076,N_12820,N_12809);
nand U13077 (N_13077,N_12877,N_12810);
or U13078 (N_13078,N_12946,N_12944);
and U13079 (N_13079,N_12959,N_12853);
or U13080 (N_13080,N_12943,N_12925);
or U13081 (N_13081,N_12784,N_12859);
or U13082 (N_13082,N_12797,N_12786);
nand U13083 (N_13083,N_12883,N_12828);
nand U13084 (N_13084,N_12757,N_12953);
or U13085 (N_13085,N_12848,N_12922);
nand U13086 (N_13086,N_12765,N_12992);
and U13087 (N_13087,N_12779,N_12812);
nor U13088 (N_13088,N_12823,N_12772);
nor U13089 (N_13089,N_12832,N_12831);
or U13090 (N_13090,N_12908,N_12806);
xnor U13091 (N_13091,N_12955,N_12916);
nor U13092 (N_13092,N_12910,N_12912);
nand U13093 (N_13093,N_12754,N_12846);
xor U13094 (N_13094,N_12931,N_12948);
and U13095 (N_13095,N_12897,N_12940);
and U13096 (N_13096,N_12780,N_12907);
or U13097 (N_13097,N_12770,N_12775);
xor U13098 (N_13098,N_12835,N_12872);
xnor U13099 (N_13099,N_12923,N_12814);
nor U13100 (N_13100,N_12873,N_12793);
nand U13101 (N_13101,N_12914,N_12867);
nor U13102 (N_13102,N_12949,N_12842);
and U13103 (N_13103,N_12919,N_12998);
and U13104 (N_13104,N_12799,N_12816);
or U13105 (N_13105,N_12825,N_12979);
nand U13106 (N_13106,N_12764,N_12819);
nor U13107 (N_13107,N_12965,N_12807);
xor U13108 (N_13108,N_12973,N_12895);
nand U13109 (N_13109,N_12858,N_12868);
nand U13110 (N_13110,N_12854,N_12845);
and U13111 (N_13111,N_12904,N_12826);
or U13112 (N_13112,N_12817,N_12857);
nand U13113 (N_13113,N_12983,N_12874);
xnor U13114 (N_13114,N_12788,N_12981);
nand U13115 (N_13115,N_12862,N_12984);
nand U13116 (N_13116,N_12837,N_12996);
nand U13117 (N_13117,N_12833,N_12783);
xor U13118 (N_13118,N_12988,N_12800);
nor U13119 (N_13119,N_12851,N_12976);
or U13120 (N_13120,N_12905,N_12947);
nor U13121 (N_13121,N_12801,N_12934);
nand U13122 (N_13122,N_12759,N_12824);
or U13123 (N_13123,N_12847,N_12781);
nor U13124 (N_13124,N_12864,N_12762);
xnor U13125 (N_13125,N_12996,N_12966);
and U13126 (N_13126,N_12788,N_12946);
nor U13127 (N_13127,N_12930,N_12774);
nand U13128 (N_13128,N_12854,N_12791);
nand U13129 (N_13129,N_12906,N_12902);
or U13130 (N_13130,N_12838,N_12895);
nand U13131 (N_13131,N_12767,N_12757);
and U13132 (N_13132,N_12889,N_12948);
nand U13133 (N_13133,N_12868,N_12768);
and U13134 (N_13134,N_12772,N_12939);
nor U13135 (N_13135,N_12820,N_12765);
or U13136 (N_13136,N_12923,N_12767);
nor U13137 (N_13137,N_12992,N_12962);
and U13138 (N_13138,N_12959,N_12856);
xor U13139 (N_13139,N_12774,N_12984);
nand U13140 (N_13140,N_12989,N_12960);
nand U13141 (N_13141,N_12930,N_12871);
or U13142 (N_13142,N_12766,N_12998);
xor U13143 (N_13143,N_12846,N_12836);
and U13144 (N_13144,N_12925,N_12824);
and U13145 (N_13145,N_12779,N_12862);
and U13146 (N_13146,N_12972,N_12871);
and U13147 (N_13147,N_12761,N_12878);
nand U13148 (N_13148,N_12993,N_12996);
and U13149 (N_13149,N_12967,N_12768);
or U13150 (N_13150,N_12974,N_12931);
or U13151 (N_13151,N_12862,N_12996);
or U13152 (N_13152,N_12974,N_12976);
nand U13153 (N_13153,N_12885,N_12757);
nor U13154 (N_13154,N_12766,N_12796);
nand U13155 (N_13155,N_12810,N_12751);
or U13156 (N_13156,N_12945,N_12801);
or U13157 (N_13157,N_12761,N_12807);
and U13158 (N_13158,N_12843,N_12769);
xnor U13159 (N_13159,N_12937,N_12841);
or U13160 (N_13160,N_12961,N_12762);
or U13161 (N_13161,N_12989,N_12918);
nor U13162 (N_13162,N_12859,N_12988);
and U13163 (N_13163,N_12758,N_12755);
or U13164 (N_13164,N_12767,N_12955);
nor U13165 (N_13165,N_12908,N_12942);
or U13166 (N_13166,N_12891,N_12873);
nor U13167 (N_13167,N_12918,N_12846);
and U13168 (N_13168,N_12988,N_12946);
nand U13169 (N_13169,N_12799,N_12814);
nand U13170 (N_13170,N_12785,N_12787);
nand U13171 (N_13171,N_12795,N_12844);
nand U13172 (N_13172,N_12909,N_12941);
xor U13173 (N_13173,N_12796,N_12846);
nor U13174 (N_13174,N_12910,N_12750);
and U13175 (N_13175,N_12872,N_12822);
nor U13176 (N_13176,N_12790,N_12996);
and U13177 (N_13177,N_12769,N_12821);
or U13178 (N_13178,N_12903,N_12876);
nand U13179 (N_13179,N_12917,N_12950);
or U13180 (N_13180,N_12927,N_12865);
nor U13181 (N_13181,N_12848,N_12934);
nor U13182 (N_13182,N_12769,N_12941);
nand U13183 (N_13183,N_12751,N_12767);
or U13184 (N_13184,N_12830,N_12983);
or U13185 (N_13185,N_12866,N_12807);
or U13186 (N_13186,N_12866,N_12819);
and U13187 (N_13187,N_12869,N_12831);
or U13188 (N_13188,N_12879,N_12847);
nand U13189 (N_13189,N_12873,N_12808);
nor U13190 (N_13190,N_12937,N_12866);
and U13191 (N_13191,N_12915,N_12966);
nor U13192 (N_13192,N_12776,N_12839);
and U13193 (N_13193,N_12791,N_12934);
nor U13194 (N_13194,N_12980,N_12898);
and U13195 (N_13195,N_12898,N_12977);
or U13196 (N_13196,N_12863,N_12971);
or U13197 (N_13197,N_12866,N_12946);
nand U13198 (N_13198,N_12950,N_12769);
nor U13199 (N_13199,N_12964,N_12976);
nor U13200 (N_13200,N_12902,N_12964);
nand U13201 (N_13201,N_12811,N_12752);
or U13202 (N_13202,N_12817,N_12977);
nand U13203 (N_13203,N_12928,N_12807);
xnor U13204 (N_13204,N_12759,N_12942);
nand U13205 (N_13205,N_12789,N_12776);
and U13206 (N_13206,N_12939,N_12877);
nor U13207 (N_13207,N_12800,N_12752);
nand U13208 (N_13208,N_12827,N_12937);
xnor U13209 (N_13209,N_12891,N_12977);
nand U13210 (N_13210,N_12815,N_12988);
or U13211 (N_13211,N_12850,N_12942);
and U13212 (N_13212,N_12767,N_12954);
nand U13213 (N_13213,N_12975,N_12988);
and U13214 (N_13214,N_12795,N_12951);
and U13215 (N_13215,N_12934,N_12964);
and U13216 (N_13216,N_12980,N_12955);
nand U13217 (N_13217,N_12793,N_12865);
xnor U13218 (N_13218,N_12937,N_12957);
xnor U13219 (N_13219,N_12892,N_12901);
nand U13220 (N_13220,N_12763,N_12872);
nor U13221 (N_13221,N_12786,N_12916);
or U13222 (N_13222,N_12951,N_12782);
or U13223 (N_13223,N_12759,N_12845);
nand U13224 (N_13224,N_12796,N_12919);
or U13225 (N_13225,N_12985,N_12984);
nor U13226 (N_13226,N_12999,N_12832);
or U13227 (N_13227,N_12773,N_12756);
xnor U13228 (N_13228,N_12953,N_12810);
or U13229 (N_13229,N_12767,N_12836);
nor U13230 (N_13230,N_12815,N_12980);
and U13231 (N_13231,N_12961,N_12852);
nand U13232 (N_13232,N_12756,N_12943);
xnor U13233 (N_13233,N_12784,N_12845);
and U13234 (N_13234,N_12988,N_12970);
nor U13235 (N_13235,N_12935,N_12808);
nand U13236 (N_13236,N_12965,N_12836);
nor U13237 (N_13237,N_12849,N_12783);
nand U13238 (N_13238,N_12806,N_12865);
nor U13239 (N_13239,N_12841,N_12911);
or U13240 (N_13240,N_12776,N_12858);
xnor U13241 (N_13241,N_12960,N_12756);
and U13242 (N_13242,N_12939,N_12757);
nor U13243 (N_13243,N_12891,N_12957);
nor U13244 (N_13244,N_12934,N_12969);
and U13245 (N_13245,N_12886,N_12804);
xor U13246 (N_13246,N_12917,N_12902);
nand U13247 (N_13247,N_12880,N_12894);
and U13248 (N_13248,N_12972,N_12770);
or U13249 (N_13249,N_12926,N_12830);
nand U13250 (N_13250,N_13145,N_13168);
nor U13251 (N_13251,N_13171,N_13102);
or U13252 (N_13252,N_13069,N_13243);
and U13253 (N_13253,N_13178,N_13101);
and U13254 (N_13254,N_13244,N_13239);
nand U13255 (N_13255,N_13127,N_13113);
nor U13256 (N_13256,N_13216,N_13128);
xnor U13257 (N_13257,N_13176,N_13172);
nor U13258 (N_13258,N_13029,N_13035);
or U13259 (N_13259,N_13068,N_13215);
or U13260 (N_13260,N_13241,N_13236);
or U13261 (N_13261,N_13193,N_13249);
or U13262 (N_13262,N_13135,N_13198);
and U13263 (N_13263,N_13201,N_13003);
nor U13264 (N_13264,N_13018,N_13206);
nor U13265 (N_13265,N_13081,N_13235);
nor U13266 (N_13266,N_13186,N_13119);
or U13267 (N_13267,N_13188,N_13051);
nor U13268 (N_13268,N_13149,N_13017);
and U13269 (N_13269,N_13181,N_13247);
or U13270 (N_13270,N_13213,N_13191);
and U13271 (N_13271,N_13082,N_13173);
or U13272 (N_13272,N_13057,N_13103);
nor U13273 (N_13273,N_13166,N_13008);
or U13274 (N_13274,N_13152,N_13070);
nand U13275 (N_13275,N_13210,N_13059);
and U13276 (N_13276,N_13220,N_13025);
xnor U13277 (N_13277,N_13091,N_13159);
or U13278 (N_13278,N_13009,N_13015);
and U13279 (N_13279,N_13155,N_13169);
and U13280 (N_13280,N_13074,N_13170);
and U13281 (N_13281,N_13162,N_13089);
nand U13282 (N_13282,N_13163,N_13177);
or U13283 (N_13283,N_13217,N_13161);
or U13284 (N_13284,N_13233,N_13147);
nor U13285 (N_13285,N_13046,N_13086);
or U13286 (N_13286,N_13043,N_13019);
nor U13287 (N_13287,N_13246,N_13223);
nand U13288 (N_13288,N_13121,N_13197);
xor U13289 (N_13289,N_13125,N_13066);
xor U13290 (N_13290,N_13150,N_13148);
nand U13291 (N_13291,N_13061,N_13226);
or U13292 (N_13292,N_13180,N_13208);
and U13293 (N_13293,N_13054,N_13242);
nand U13294 (N_13294,N_13189,N_13209);
nand U13295 (N_13295,N_13122,N_13211);
and U13296 (N_13296,N_13134,N_13062);
nor U13297 (N_13297,N_13144,N_13165);
nor U13298 (N_13298,N_13240,N_13232);
or U13299 (N_13299,N_13117,N_13084);
and U13300 (N_13300,N_13027,N_13204);
and U13301 (N_13301,N_13228,N_13196);
nand U13302 (N_13302,N_13199,N_13065);
and U13303 (N_13303,N_13092,N_13112);
and U13304 (N_13304,N_13049,N_13120);
nor U13305 (N_13305,N_13079,N_13229);
or U13306 (N_13306,N_13090,N_13230);
nor U13307 (N_13307,N_13225,N_13158);
nor U13308 (N_13308,N_13023,N_13203);
nand U13309 (N_13309,N_13221,N_13037);
nand U13310 (N_13310,N_13205,N_13004);
and U13311 (N_13311,N_13234,N_13187);
nand U13312 (N_13312,N_13021,N_13028);
or U13313 (N_13313,N_13108,N_13156);
and U13314 (N_13314,N_13093,N_13100);
or U13315 (N_13315,N_13000,N_13096);
or U13316 (N_13316,N_13099,N_13055);
nor U13317 (N_13317,N_13056,N_13073);
nor U13318 (N_13318,N_13105,N_13040);
nand U13319 (N_13319,N_13227,N_13106);
nand U13320 (N_13320,N_13248,N_13031);
nand U13321 (N_13321,N_13110,N_13131);
and U13322 (N_13322,N_13080,N_13047);
xnor U13323 (N_13323,N_13116,N_13001);
nand U13324 (N_13324,N_13067,N_13077);
nor U13325 (N_13325,N_13095,N_13164);
nand U13326 (N_13326,N_13151,N_13050);
and U13327 (N_13327,N_13041,N_13042);
or U13328 (N_13328,N_13111,N_13130);
nand U13329 (N_13329,N_13032,N_13142);
or U13330 (N_13330,N_13154,N_13052);
nor U13331 (N_13331,N_13034,N_13139);
nand U13332 (N_13332,N_13011,N_13076);
or U13333 (N_13333,N_13140,N_13184);
or U13334 (N_13334,N_13022,N_13048);
or U13335 (N_13335,N_13072,N_13219);
and U13336 (N_13336,N_13207,N_13114);
or U13337 (N_13337,N_13174,N_13195);
nand U13338 (N_13338,N_13238,N_13013);
nor U13339 (N_13339,N_13104,N_13020);
nor U13340 (N_13340,N_13097,N_13094);
and U13341 (N_13341,N_13146,N_13123);
xnor U13342 (N_13342,N_13045,N_13007);
and U13343 (N_13343,N_13024,N_13214);
and U13344 (N_13344,N_13129,N_13194);
nor U13345 (N_13345,N_13085,N_13064);
or U13346 (N_13346,N_13016,N_13118);
nor U13347 (N_13347,N_13138,N_13087);
and U13348 (N_13348,N_13083,N_13115);
or U13349 (N_13349,N_13014,N_13039);
nand U13350 (N_13350,N_13190,N_13237);
or U13351 (N_13351,N_13044,N_13132);
nor U13352 (N_13352,N_13109,N_13141);
and U13353 (N_13353,N_13036,N_13218);
nand U13354 (N_13354,N_13192,N_13136);
and U13355 (N_13355,N_13075,N_13124);
and U13356 (N_13356,N_13005,N_13183);
xnor U13357 (N_13357,N_13212,N_13060);
nand U13358 (N_13358,N_13179,N_13098);
and U13359 (N_13359,N_13058,N_13143);
nor U13360 (N_13360,N_13010,N_13160);
and U13361 (N_13361,N_13063,N_13126);
and U13362 (N_13362,N_13030,N_13012);
and U13363 (N_13363,N_13071,N_13078);
or U13364 (N_13364,N_13137,N_13107);
nor U13365 (N_13365,N_13002,N_13245);
nor U13366 (N_13366,N_13038,N_13153);
nand U13367 (N_13367,N_13006,N_13231);
nor U13368 (N_13368,N_13222,N_13053);
nor U13369 (N_13369,N_13033,N_13185);
nor U13370 (N_13370,N_13224,N_13202);
nor U13371 (N_13371,N_13200,N_13182);
nand U13372 (N_13372,N_13167,N_13157);
nor U13373 (N_13373,N_13175,N_13026);
nand U13374 (N_13374,N_13133,N_13088);
nor U13375 (N_13375,N_13077,N_13171);
nand U13376 (N_13376,N_13034,N_13138);
nor U13377 (N_13377,N_13080,N_13115);
xnor U13378 (N_13378,N_13170,N_13033);
or U13379 (N_13379,N_13180,N_13101);
or U13380 (N_13380,N_13140,N_13070);
or U13381 (N_13381,N_13097,N_13069);
and U13382 (N_13382,N_13081,N_13244);
nand U13383 (N_13383,N_13196,N_13175);
nand U13384 (N_13384,N_13001,N_13052);
nand U13385 (N_13385,N_13145,N_13119);
nor U13386 (N_13386,N_13059,N_13053);
and U13387 (N_13387,N_13141,N_13034);
and U13388 (N_13388,N_13035,N_13131);
and U13389 (N_13389,N_13141,N_13002);
and U13390 (N_13390,N_13232,N_13134);
nor U13391 (N_13391,N_13208,N_13044);
xor U13392 (N_13392,N_13186,N_13244);
nor U13393 (N_13393,N_13107,N_13044);
or U13394 (N_13394,N_13112,N_13248);
or U13395 (N_13395,N_13025,N_13074);
nand U13396 (N_13396,N_13121,N_13027);
or U13397 (N_13397,N_13222,N_13074);
or U13398 (N_13398,N_13139,N_13143);
and U13399 (N_13399,N_13152,N_13027);
or U13400 (N_13400,N_13032,N_13117);
and U13401 (N_13401,N_13038,N_13062);
and U13402 (N_13402,N_13193,N_13057);
or U13403 (N_13403,N_13228,N_13045);
and U13404 (N_13404,N_13121,N_13196);
xor U13405 (N_13405,N_13189,N_13106);
and U13406 (N_13406,N_13040,N_13072);
nand U13407 (N_13407,N_13181,N_13025);
nand U13408 (N_13408,N_13137,N_13110);
nor U13409 (N_13409,N_13056,N_13075);
nor U13410 (N_13410,N_13222,N_13099);
or U13411 (N_13411,N_13190,N_13162);
and U13412 (N_13412,N_13116,N_13005);
nor U13413 (N_13413,N_13241,N_13153);
or U13414 (N_13414,N_13198,N_13136);
or U13415 (N_13415,N_13106,N_13199);
nand U13416 (N_13416,N_13040,N_13066);
nor U13417 (N_13417,N_13148,N_13198);
and U13418 (N_13418,N_13157,N_13116);
nand U13419 (N_13419,N_13127,N_13220);
nand U13420 (N_13420,N_13211,N_13077);
nor U13421 (N_13421,N_13217,N_13002);
xnor U13422 (N_13422,N_13125,N_13028);
nand U13423 (N_13423,N_13022,N_13133);
or U13424 (N_13424,N_13249,N_13062);
and U13425 (N_13425,N_13233,N_13001);
or U13426 (N_13426,N_13038,N_13227);
nor U13427 (N_13427,N_13008,N_13035);
nor U13428 (N_13428,N_13207,N_13013);
or U13429 (N_13429,N_13204,N_13235);
nor U13430 (N_13430,N_13231,N_13226);
or U13431 (N_13431,N_13084,N_13051);
nand U13432 (N_13432,N_13199,N_13248);
nor U13433 (N_13433,N_13047,N_13161);
and U13434 (N_13434,N_13163,N_13115);
nor U13435 (N_13435,N_13135,N_13120);
nand U13436 (N_13436,N_13087,N_13021);
or U13437 (N_13437,N_13200,N_13169);
or U13438 (N_13438,N_13108,N_13181);
nor U13439 (N_13439,N_13167,N_13026);
nand U13440 (N_13440,N_13112,N_13014);
nand U13441 (N_13441,N_13219,N_13005);
xor U13442 (N_13442,N_13136,N_13070);
nand U13443 (N_13443,N_13063,N_13173);
nand U13444 (N_13444,N_13106,N_13116);
or U13445 (N_13445,N_13248,N_13222);
nor U13446 (N_13446,N_13191,N_13093);
nand U13447 (N_13447,N_13040,N_13131);
nand U13448 (N_13448,N_13105,N_13129);
or U13449 (N_13449,N_13224,N_13091);
and U13450 (N_13450,N_13114,N_13008);
nor U13451 (N_13451,N_13139,N_13132);
or U13452 (N_13452,N_13194,N_13082);
or U13453 (N_13453,N_13202,N_13108);
nand U13454 (N_13454,N_13007,N_13203);
and U13455 (N_13455,N_13248,N_13167);
and U13456 (N_13456,N_13176,N_13118);
or U13457 (N_13457,N_13162,N_13170);
nand U13458 (N_13458,N_13054,N_13247);
nor U13459 (N_13459,N_13149,N_13125);
nand U13460 (N_13460,N_13054,N_13039);
nor U13461 (N_13461,N_13204,N_13046);
nand U13462 (N_13462,N_13072,N_13022);
and U13463 (N_13463,N_13236,N_13071);
and U13464 (N_13464,N_13215,N_13020);
nand U13465 (N_13465,N_13100,N_13194);
nand U13466 (N_13466,N_13090,N_13149);
or U13467 (N_13467,N_13213,N_13236);
or U13468 (N_13468,N_13205,N_13238);
nor U13469 (N_13469,N_13092,N_13236);
and U13470 (N_13470,N_13120,N_13127);
nand U13471 (N_13471,N_13238,N_13115);
or U13472 (N_13472,N_13131,N_13175);
and U13473 (N_13473,N_13198,N_13178);
nor U13474 (N_13474,N_13043,N_13221);
or U13475 (N_13475,N_13176,N_13098);
and U13476 (N_13476,N_13062,N_13166);
and U13477 (N_13477,N_13163,N_13078);
or U13478 (N_13478,N_13152,N_13125);
or U13479 (N_13479,N_13246,N_13055);
nand U13480 (N_13480,N_13025,N_13235);
nor U13481 (N_13481,N_13000,N_13173);
nor U13482 (N_13482,N_13164,N_13092);
or U13483 (N_13483,N_13066,N_13087);
nor U13484 (N_13484,N_13000,N_13162);
or U13485 (N_13485,N_13146,N_13128);
nor U13486 (N_13486,N_13224,N_13148);
nor U13487 (N_13487,N_13226,N_13018);
and U13488 (N_13488,N_13127,N_13060);
or U13489 (N_13489,N_13120,N_13145);
and U13490 (N_13490,N_13006,N_13159);
or U13491 (N_13491,N_13035,N_13013);
nand U13492 (N_13492,N_13217,N_13031);
nor U13493 (N_13493,N_13118,N_13084);
nor U13494 (N_13494,N_13102,N_13106);
xor U13495 (N_13495,N_13050,N_13134);
nand U13496 (N_13496,N_13158,N_13189);
nand U13497 (N_13497,N_13099,N_13204);
nand U13498 (N_13498,N_13115,N_13087);
and U13499 (N_13499,N_13240,N_13246);
or U13500 (N_13500,N_13254,N_13412);
and U13501 (N_13501,N_13405,N_13463);
xor U13502 (N_13502,N_13380,N_13329);
and U13503 (N_13503,N_13324,N_13437);
nor U13504 (N_13504,N_13394,N_13481);
nor U13505 (N_13505,N_13343,N_13474);
nor U13506 (N_13506,N_13383,N_13363);
nand U13507 (N_13507,N_13339,N_13453);
nor U13508 (N_13508,N_13422,N_13365);
nand U13509 (N_13509,N_13425,N_13390);
nor U13510 (N_13510,N_13299,N_13288);
nand U13511 (N_13511,N_13452,N_13350);
or U13512 (N_13512,N_13421,N_13284);
nor U13513 (N_13513,N_13456,N_13472);
or U13514 (N_13514,N_13256,N_13257);
xor U13515 (N_13515,N_13478,N_13389);
nand U13516 (N_13516,N_13443,N_13442);
nand U13517 (N_13517,N_13308,N_13417);
or U13518 (N_13518,N_13351,N_13419);
or U13519 (N_13519,N_13427,N_13346);
nand U13520 (N_13520,N_13325,N_13263);
nand U13521 (N_13521,N_13391,N_13496);
nor U13522 (N_13522,N_13468,N_13392);
or U13523 (N_13523,N_13440,N_13438);
nor U13524 (N_13524,N_13447,N_13337);
nand U13525 (N_13525,N_13251,N_13345);
nand U13526 (N_13526,N_13295,N_13262);
xnor U13527 (N_13527,N_13276,N_13283);
and U13528 (N_13528,N_13287,N_13471);
nor U13529 (N_13529,N_13489,N_13282);
and U13530 (N_13530,N_13448,N_13432);
nor U13531 (N_13531,N_13445,N_13358);
nor U13532 (N_13532,N_13255,N_13398);
or U13533 (N_13533,N_13498,N_13424);
xnor U13534 (N_13534,N_13364,N_13483);
or U13535 (N_13535,N_13289,N_13428);
xor U13536 (N_13536,N_13435,N_13334);
nand U13537 (N_13537,N_13371,N_13367);
or U13538 (N_13538,N_13356,N_13261);
xnor U13539 (N_13539,N_13355,N_13477);
nand U13540 (N_13540,N_13304,N_13436);
nand U13541 (N_13541,N_13354,N_13279);
nor U13542 (N_13542,N_13401,N_13360);
nand U13543 (N_13543,N_13485,N_13488);
nand U13544 (N_13544,N_13273,N_13476);
or U13545 (N_13545,N_13470,N_13395);
and U13546 (N_13546,N_13451,N_13396);
xnor U13547 (N_13547,N_13497,N_13321);
and U13548 (N_13548,N_13366,N_13306);
xor U13549 (N_13549,N_13336,N_13335);
nor U13550 (N_13550,N_13397,N_13480);
and U13551 (N_13551,N_13406,N_13313);
or U13552 (N_13552,N_13423,N_13487);
or U13553 (N_13553,N_13409,N_13384);
and U13554 (N_13554,N_13326,N_13449);
nor U13555 (N_13555,N_13332,N_13490);
and U13556 (N_13556,N_13466,N_13331);
xor U13557 (N_13557,N_13382,N_13333);
or U13558 (N_13558,N_13362,N_13462);
nor U13559 (N_13559,N_13265,N_13312);
or U13560 (N_13560,N_13486,N_13464);
or U13561 (N_13561,N_13361,N_13385);
nor U13562 (N_13562,N_13387,N_13274);
xor U13563 (N_13563,N_13297,N_13270);
nand U13564 (N_13564,N_13266,N_13376);
xor U13565 (N_13565,N_13473,N_13340);
or U13566 (N_13566,N_13482,N_13374);
nor U13567 (N_13567,N_13375,N_13402);
xor U13568 (N_13568,N_13353,N_13441);
or U13569 (N_13569,N_13431,N_13311);
and U13570 (N_13570,N_13458,N_13260);
nor U13571 (N_13571,N_13454,N_13357);
or U13572 (N_13572,N_13269,N_13281);
nor U13573 (N_13573,N_13352,N_13460);
and U13574 (N_13574,N_13268,N_13399);
and U13575 (N_13575,N_13475,N_13479);
and U13576 (N_13576,N_13317,N_13416);
nor U13577 (N_13577,N_13264,N_13393);
and U13578 (N_13578,N_13259,N_13323);
or U13579 (N_13579,N_13450,N_13499);
nand U13580 (N_13580,N_13495,N_13293);
nand U13581 (N_13581,N_13258,N_13444);
nor U13582 (N_13582,N_13461,N_13408);
nor U13583 (N_13583,N_13400,N_13338);
and U13584 (N_13584,N_13349,N_13253);
and U13585 (N_13585,N_13347,N_13280);
nor U13586 (N_13586,N_13301,N_13348);
or U13587 (N_13587,N_13314,N_13373);
nor U13588 (N_13588,N_13493,N_13369);
and U13589 (N_13589,N_13344,N_13403);
or U13590 (N_13590,N_13286,N_13319);
nor U13591 (N_13591,N_13309,N_13429);
nand U13592 (N_13592,N_13252,N_13418);
or U13593 (N_13593,N_13302,N_13250);
nor U13594 (N_13594,N_13320,N_13469);
nor U13595 (N_13595,N_13410,N_13491);
and U13596 (N_13596,N_13372,N_13420);
nand U13597 (N_13597,N_13272,N_13315);
and U13598 (N_13598,N_13296,N_13271);
nand U13599 (N_13599,N_13341,N_13434);
nor U13600 (N_13600,N_13298,N_13379);
and U13601 (N_13601,N_13430,N_13381);
and U13602 (N_13602,N_13414,N_13307);
or U13603 (N_13603,N_13492,N_13411);
nand U13604 (N_13604,N_13404,N_13327);
and U13605 (N_13605,N_13328,N_13310);
nor U13606 (N_13606,N_13292,N_13316);
nand U13607 (N_13607,N_13370,N_13285);
and U13608 (N_13608,N_13368,N_13457);
nand U13609 (N_13609,N_13465,N_13407);
nor U13610 (N_13610,N_13330,N_13386);
nor U13611 (N_13611,N_13277,N_13388);
xnor U13612 (N_13612,N_13494,N_13342);
or U13613 (N_13613,N_13294,N_13267);
or U13614 (N_13614,N_13318,N_13433);
and U13615 (N_13615,N_13290,N_13359);
nor U13616 (N_13616,N_13378,N_13322);
xor U13617 (N_13617,N_13305,N_13415);
nor U13618 (N_13618,N_13439,N_13275);
nand U13619 (N_13619,N_13467,N_13291);
xor U13620 (N_13620,N_13377,N_13300);
nor U13621 (N_13621,N_13455,N_13446);
nor U13622 (N_13622,N_13484,N_13303);
nand U13623 (N_13623,N_13413,N_13459);
nand U13624 (N_13624,N_13426,N_13278);
and U13625 (N_13625,N_13293,N_13358);
or U13626 (N_13626,N_13362,N_13473);
nor U13627 (N_13627,N_13385,N_13444);
nand U13628 (N_13628,N_13475,N_13486);
nor U13629 (N_13629,N_13286,N_13450);
or U13630 (N_13630,N_13454,N_13322);
nand U13631 (N_13631,N_13481,N_13456);
or U13632 (N_13632,N_13304,N_13292);
and U13633 (N_13633,N_13435,N_13259);
nor U13634 (N_13634,N_13468,N_13257);
nand U13635 (N_13635,N_13280,N_13283);
nand U13636 (N_13636,N_13475,N_13313);
and U13637 (N_13637,N_13330,N_13305);
nor U13638 (N_13638,N_13474,N_13490);
or U13639 (N_13639,N_13332,N_13265);
and U13640 (N_13640,N_13372,N_13289);
nand U13641 (N_13641,N_13404,N_13263);
nor U13642 (N_13642,N_13492,N_13283);
and U13643 (N_13643,N_13349,N_13341);
xor U13644 (N_13644,N_13492,N_13276);
or U13645 (N_13645,N_13393,N_13359);
or U13646 (N_13646,N_13443,N_13364);
nor U13647 (N_13647,N_13322,N_13331);
or U13648 (N_13648,N_13469,N_13328);
nor U13649 (N_13649,N_13393,N_13491);
nand U13650 (N_13650,N_13321,N_13468);
xor U13651 (N_13651,N_13497,N_13451);
nor U13652 (N_13652,N_13310,N_13383);
and U13653 (N_13653,N_13289,N_13407);
nor U13654 (N_13654,N_13272,N_13367);
nor U13655 (N_13655,N_13317,N_13307);
and U13656 (N_13656,N_13373,N_13263);
nand U13657 (N_13657,N_13467,N_13274);
and U13658 (N_13658,N_13300,N_13474);
nand U13659 (N_13659,N_13386,N_13406);
nor U13660 (N_13660,N_13405,N_13413);
nand U13661 (N_13661,N_13340,N_13258);
nand U13662 (N_13662,N_13280,N_13281);
and U13663 (N_13663,N_13318,N_13391);
nand U13664 (N_13664,N_13468,N_13493);
nor U13665 (N_13665,N_13270,N_13324);
nor U13666 (N_13666,N_13380,N_13307);
nor U13667 (N_13667,N_13374,N_13330);
and U13668 (N_13668,N_13309,N_13341);
nor U13669 (N_13669,N_13282,N_13431);
nand U13670 (N_13670,N_13392,N_13345);
nor U13671 (N_13671,N_13462,N_13400);
or U13672 (N_13672,N_13296,N_13471);
nand U13673 (N_13673,N_13334,N_13360);
or U13674 (N_13674,N_13356,N_13337);
nand U13675 (N_13675,N_13316,N_13267);
nand U13676 (N_13676,N_13256,N_13367);
or U13677 (N_13677,N_13381,N_13303);
and U13678 (N_13678,N_13454,N_13498);
or U13679 (N_13679,N_13417,N_13470);
nand U13680 (N_13680,N_13327,N_13439);
nand U13681 (N_13681,N_13327,N_13300);
and U13682 (N_13682,N_13491,N_13300);
and U13683 (N_13683,N_13375,N_13440);
and U13684 (N_13684,N_13463,N_13389);
and U13685 (N_13685,N_13413,N_13452);
and U13686 (N_13686,N_13342,N_13442);
nand U13687 (N_13687,N_13270,N_13277);
and U13688 (N_13688,N_13279,N_13267);
nand U13689 (N_13689,N_13478,N_13462);
or U13690 (N_13690,N_13375,N_13429);
nor U13691 (N_13691,N_13432,N_13400);
and U13692 (N_13692,N_13319,N_13274);
or U13693 (N_13693,N_13493,N_13437);
xnor U13694 (N_13694,N_13278,N_13292);
and U13695 (N_13695,N_13307,N_13365);
nand U13696 (N_13696,N_13338,N_13286);
nor U13697 (N_13697,N_13369,N_13404);
xor U13698 (N_13698,N_13414,N_13263);
and U13699 (N_13699,N_13397,N_13279);
or U13700 (N_13700,N_13252,N_13459);
and U13701 (N_13701,N_13334,N_13414);
or U13702 (N_13702,N_13343,N_13303);
nand U13703 (N_13703,N_13405,N_13494);
or U13704 (N_13704,N_13407,N_13487);
nand U13705 (N_13705,N_13255,N_13357);
nand U13706 (N_13706,N_13289,N_13432);
nand U13707 (N_13707,N_13392,N_13477);
xnor U13708 (N_13708,N_13265,N_13325);
and U13709 (N_13709,N_13346,N_13420);
nand U13710 (N_13710,N_13343,N_13440);
nor U13711 (N_13711,N_13420,N_13395);
and U13712 (N_13712,N_13398,N_13361);
or U13713 (N_13713,N_13419,N_13337);
xor U13714 (N_13714,N_13287,N_13486);
and U13715 (N_13715,N_13367,N_13389);
or U13716 (N_13716,N_13388,N_13295);
xor U13717 (N_13717,N_13477,N_13277);
and U13718 (N_13718,N_13333,N_13486);
nand U13719 (N_13719,N_13391,N_13421);
nand U13720 (N_13720,N_13434,N_13263);
nor U13721 (N_13721,N_13322,N_13264);
xnor U13722 (N_13722,N_13304,N_13302);
nor U13723 (N_13723,N_13284,N_13433);
nor U13724 (N_13724,N_13330,N_13422);
or U13725 (N_13725,N_13488,N_13315);
and U13726 (N_13726,N_13257,N_13459);
nor U13727 (N_13727,N_13489,N_13378);
nand U13728 (N_13728,N_13320,N_13297);
nor U13729 (N_13729,N_13307,N_13484);
nor U13730 (N_13730,N_13463,N_13310);
and U13731 (N_13731,N_13481,N_13342);
or U13732 (N_13732,N_13326,N_13406);
and U13733 (N_13733,N_13372,N_13453);
nand U13734 (N_13734,N_13409,N_13395);
or U13735 (N_13735,N_13488,N_13405);
and U13736 (N_13736,N_13297,N_13373);
and U13737 (N_13737,N_13291,N_13476);
nor U13738 (N_13738,N_13494,N_13377);
nand U13739 (N_13739,N_13293,N_13291);
nor U13740 (N_13740,N_13459,N_13458);
or U13741 (N_13741,N_13289,N_13350);
nor U13742 (N_13742,N_13266,N_13324);
nand U13743 (N_13743,N_13320,N_13433);
or U13744 (N_13744,N_13428,N_13268);
and U13745 (N_13745,N_13354,N_13361);
nor U13746 (N_13746,N_13336,N_13250);
or U13747 (N_13747,N_13331,N_13256);
or U13748 (N_13748,N_13483,N_13286);
nor U13749 (N_13749,N_13323,N_13421);
and U13750 (N_13750,N_13694,N_13529);
nand U13751 (N_13751,N_13622,N_13562);
xor U13752 (N_13752,N_13651,N_13636);
nand U13753 (N_13753,N_13702,N_13656);
nor U13754 (N_13754,N_13717,N_13723);
nor U13755 (N_13755,N_13524,N_13688);
nor U13756 (N_13756,N_13720,N_13658);
nand U13757 (N_13757,N_13510,N_13654);
nand U13758 (N_13758,N_13724,N_13737);
nor U13759 (N_13759,N_13729,N_13508);
and U13760 (N_13760,N_13674,N_13744);
nor U13761 (N_13761,N_13573,N_13578);
nand U13762 (N_13762,N_13697,N_13610);
nor U13763 (N_13763,N_13653,N_13617);
nor U13764 (N_13764,N_13568,N_13725);
nand U13765 (N_13765,N_13649,N_13684);
nand U13766 (N_13766,N_13618,N_13671);
nand U13767 (N_13767,N_13582,N_13629);
nor U13768 (N_13768,N_13619,N_13580);
nand U13769 (N_13769,N_13544,N_13687);
and U13770 (N_13770,N_13650,N_13581);
or U13771 (N_13771,N_13552,N_13545);
nand U13772 (N_13772,N_13594,N_13696);
nor U13773 (N_13773,N_13706,N_13742);
nor U13774 (N_13774,N_13728,N_13634);
xor U13775 (N_13775,N_13563,N_13628);
or U13776 (N_13776,N_13553,N_13519);
and U13777 (N_13777,N_13556,N_13741);
xnor U13778 (N_13778,N_13542,N_13588);
nor U13779 (N_13779,N_13716,N_13539);
nor U13780 (N_13780,N_13740,N_13596);
nor U13781 (N_13781,N_13565,N_13743);
nand U13782 (N_13782,N_13733,N_13685);
or U13783 (N_13783,N_13527,N_13583);
xnor U13784 (N_13784,N_13659,N_13749);
or U13785 (N_13785,N_13615,N_13730);
and U13786 (N_13786,N_13734,N_13567);
nand U13787 (N_13787,N_13709,N_13576);
or U13788 (N_13788,N_13599,N_13558);
nand U13789 (N_13789,N_13536,N_13606);
or U13790 (N_13790,N_13712,N_13708);
xnor U13791 (N_13791,N_13526,N_13623);
or U13792 (N_13792,N_13633,N_13661);
xnor U13793 (N_13793,N_13603,N_13630);
and U13794 (N_13794,N_13589,N_13555);
nor U13795 (N_13795,N_13604,N_13745);
nand U13796 (N_13796,N_13692,N_13640);
or U13797 (N_13797,N_13657,N_13520);
nor U13798 (N_13798,N_13531,N_13530);
nand U13799 (N_13799,N_13516,N_13592);
xnor U13800 (N_13800,N_13572,N_13523);
or U13801 (N_13801,N_13501,N_13509);
nor U13802 (N_13802,N_13597,N_13655);
or U13803 (N_13803,N_13566,N_13505);
or U13804 (N_13804,N_13705,N_13593);
nor U13805 (N_13805,N_13660,N_13718);
xnor U13806 (N_13806,N_13550,N_13626);
nor U13807 (N_13807,N_13643,N_13605);
and U13808 (N_13808,N_13500,N_13665);
nand U13809 (N_13809,N_13642,N_13514);
nor U13810 (N_13810,N_13574,N_13504);
and U13811 (N_13811,N_13675,N_13631);
nor U13812 (N_13812,N_13732,N_13584);
and U13813 (N_13813,N_13731,N_13557);
nand U13814 (N_13814,N_13561,N_13746);
or U13815 (N_13815,N_13513,N_13644);
and U13816 (N_13816,N_13736,N_13739);
or U13817 (N_13817,N_13602,N_13668);
nor U13818 (N_13818,N_13662,N_13543);
or U13819 (N_13819,N_13595,N_13547);
nor U13820 (N_13820,N_13652,N_13548);
nor U13821 (N_13821,N_13707,N_13682);
nand U13822 (N_13822,N_13637,N_13699);
nand U13823 (N_13823,N_13598,N_13546);
nor U13824 (N_13824,N_13689,N_13667);
and U13825 (N_13825,N_13669,N_13620);
or U13826 (N_13826,N_13535,N_13570);
and U13827 (N_13827,N_13683,N_13738);
nor U13828 (N_13828,N_13735,N_13616);
nand U13829 (N_13829,N_13673,N_13710);
nor U13830 (N_13830,N_13502,N_13571);
nor U13831 (N_13831,N_13690,N_13612);
or U13832 (N_13832,N_13635,N_13569);
and U13833 (N_13833,N_13511,N_13506);
and U13834 (N_13834,N_13704,N_13670);
or U13835 (N_13835,N_13666,N_13621);
xnor U13836 (N_13836,N_13693,N_13715);
nor U13837 (N_13837,N_13577,N_13638);
nand U13838 (N_13838,N_13686,N_13517);
or U13839 (N_13839,N_13522,N_13645);
nand U13840 (N_13840,N_13528,N_13721);
or U13841 (N_13841,N_13679,N_13714);
or U13842 (N_13842,N_13691,N_13747);
xnor U13843 (N_13843,N_13538,N_13680);
nand U13844 (N_13844,N_13719,N_13587);
or U13845 (N_13845,N_13575,N_13559);
and U13846 (N_13846,N_13541,N_13512);
nand U13847 (N_13847,N_13611,N_13534);
or U13848 (N_13848,N_13678,N_13601);
nor U13849 (N_13849,N_13532,N_13748);
nor U13850 (N_13850,N_13701,N_13591);
nand U13851 (N_13851,N_13560,N_13681);
and U13852 (N_13852,N_13607,N_13549);
nor U13853 (N_13853,N_13585,N_13663);
nor U13854 (N_13854,N_13722,N_13537);
and U13855 (N_13855,N_13727,N_13700);
and U13856 (N_13856,N_13521,N_13627);
or U13857 (N_13857,N_13518,N_13503);
nand U13858 (N_13858,N_13713,N_13507);
xor U13859 (N_13859,N_13590,N_13726);
nand U13860 (N_13860,N_13609,N_13608);
xnor U13861 (N_13861,N_13600,N_13641);
and U13862 (N_13862,N_13540,N_13647);
nor U13863 (N_13863,N_13632,N_13672);
nand U13864 (N_13864,N_13551,N_13646);
nor U13865 (N_13865,N_13676,N_13613);
nand U13866 (N_13866,N_13703,N_13698);
and U13867 (N_13867,N_13614,N_13525);
nor U13868 (N_13868,N_13648,N_13624);
nand U13869 (N_13869,N_13564,N_13515);
nand U13870 (N_13870,N_13711,N_13586);
nand U13871 (N_13871,N_13554,N_13579);
or U13872 (N_13872,N_13639,N_13677);
and U13873 (N_13873,N_13664,N_13695);
or U13874 (N_13874,N_13625,N_13533);
or U13875 (N_13875,N_13593,N_13508);
xnor U13876 (N_13876,N_13583,N_13668);
nand U13877 (N_13877,N_13643,N_13600);
nand U13878 (N_13878,N_13594,N_13522);
or U13879 (N_13879,N_13586,N_13710);
and U13880 (N_13880,N_13566,N_13518);
nand U13881 (N_13881,N_13614,N_13682);
nand U13882 (N_13882,N_13518,N_13660);
and U13883 (N_13883,N_13706,N_13741);
nor U13884 (N_13884,N_13621,N_13517);
and U13885 (N_13885,N_13523,N_13605);
xor U13886 (N_13886,N_13525,N_13557);
or U13887 (N_13887,N_13618,N_13564);
nand U13888 (N_13888,N_13676,N_13706);
and U13889 (N_13889,N_13722,N_13522);
nand U13890 (N_13890,N_13575,N_13639);
and U13891 (N_13891,N_13615,N_13662);
or U13892 (N_13892,N_13507,N_13739);
xor U13893 (N_13893,N_13619,N_13584);
nor U13894 (N_13894,N_13715,N_13625);
nand U13895 (N_13895,N_13667,N_13575);
nand U13896 (N_13896,N_13749,N_13522);
nand U13897 (N_13897,N_13577,N_13707);
and U13898 (N_13898,N_13687,N_13516);
or U13899 (N_13899,N_13630,N_13715);
or U13900 (N_13900,N_13690,N_13530);
or U13901 (N_13901,N_13568,N_13536);
nand U13902 (N_13902,N_13715,N_13686);
nand U13903 (N_13903,N_13582,N_13655);
nor U13904 (N_13904,N_13605,N_13510);
nor U13905 (N_13905,N_13696,N_13610);
or U13906 (N_13906,N_13533,N_13637);
nand U13907 (N_13907,N_13664,N_13619);
nor U13908 (N_13908,N_13508,N_13643);
and U13909 (N_13909,N_13569,N_13702);
and U13910 (N_13910,N_13687,N_13517);
and U13911 (N_13911,N_13524,N_13572);
nor U13912 (N_13912,N_13714,N_13560);
and U13913 (N_13913,N_13606,N_13555);
and U13914 (N_13914,N_13552,N_13699);
or U13915 (N_13915,N_13522,N_13634);
or U13916 (N_13916,N_13619,N_13655);
nand U13917 (N_13917,N_13654,N_13675);
and U13918 (N_13918,N_13572,N_13529);
or U13919 (N_13919,N_13535,N_13669);
nand U13920 (N_13920,N_13579,N_13523);
and U13921 (N_13921,N_13682,N_13548);
nor U13922 (N_13922,N_13710,N_13681);
nand U13923 (N_13923,N_13694,N_13637);
or U13924 (N_13924,N_13619,N_13642);
or U13925 (N_13925,N_13602,N_13656);
or U13926 (N_13926,N_13714,N_13525);
nand U13927 (N_13927,N_13560,N_13579);
or U13928 (N_13928,N_13666,N_13524);
nand U13929 (N_13929,N_13739,N_13660);
and U13930 (N_13930,N_13735,N_13708);
nand U13931 (N_13931,N_13667,N_13583);
xnor U13932 (N_13932,N_13673,N_13533);
or U13933 (N_13933,N_13615,N_13572);
and U13934 (N_13934,N_13710,N_13620);
nand U13935 (N_13935,N_13729,N_13678);
xor U13936 (N_13936,N_13587,N_13645);
xnor U13937 (N_13937,N_13584,N_13749);
or U13938 (N_13938,N_13688,N_13744);
nand U13939 (N_13939,N_13571,N_13504);
or U13940 (N_13940,N_13687,N_13525);
and U13941 (N_13941,N_13669,N_13681);
or U13942 (N_13942,N_13596,N_13540);
and U13943 (N_13943,N_13598,N_13577);
and U13944 (N_13944,N_13536,N_13520);
or U13945 (N_13945,N_13726,N_13532);
nor U13946 (N_13946,N_13742,N_13539);
or U13947 (N_13947,N_13621,N_13606);
or U13948 (N_13948,N_13718,N_13739);
nor U13949 (N_13949,N_13682,N_13665);
nand U13950 (N_13950,N_13604,N_13569);
and U13951 (N_13951,N_13512,N_13685);
xnor U13952 (N_13952,N_13734,N_13561);
nor U13953 (N_13953,N_13516,N_13590);
nand U13954 (N_13954,N_13505,N_13609);
nand U13955 (N_13955,N_13672,N_13673);
nor U13956 (N_13956,N_13543,N_13747);
xor U13957 (N_13957,N_13680,N_13600);
or U13958 (N_13958,N_13749,N_13689);
nor U13959 (N_13959,N_13727,N_13541);
and U13960 (N_13960,N_13546,N_13513);
xor U13961 (N_13961,N_13532,N_13682);
and U13962 (N_13962,N_13606,N_13741);
or U13963 (N_13963,N_13622,N_13535);
and U13964 (N_13964,N_13560,N_13500);
nor U13965 (N_13965,N_13631,N_13619);
or U13966 (N_13966,N_13611,N_13586);
xnor U13967 (N_13967,N_13741,N_13733);
nand U13968 (N_13968,N_13736,N_13554);
nor U13969 (N_13969,N_13594,N_13679);
or U13970 (N_13970,N_13519,N_13612);
xnor U13971 (N_13971,N_13530,N_13668);
or U13972 (N_13972,N_13740,N_13609);
xnor U13973 (N_13973,N_13738,N_13730);
xnor U13974 (N_13974,N_13611,N_13558);
nor U13975 (N_13975,N_13747,N_13650);
nand U13976 (N_13976,N_13578,N_13693);
and U13977 (N_13977,N_13579,N_13662);
xnor U13978 (N_13978,N_13650,N_13628);
and U13979 (N_13979,N_13693,N_13528);
or U13980 (N_13980,N_13503,N_13566);
nand U13981 (N_13981,N_13616,N_13530);
nand U13982 (N_13982,N_13707,N_13580);
nand U13983 (N_13983,N_13576,N_13605);
and U13984 (N_13984,N_13619,N_13657);
nor U13985 (N_13985,N_13645,N_13636);
and U13986 (N_13986,N_13637,N_13658);
nor U13987 (N_13987,N_13547,N_13535);
or U13988 (N_13988,N_13684,N_13645);
nor U13989 (N_13989,N_13665,N_13743);
nand U13990 (N_13990,N_13631,N_13706);
nand U13991 (N_13991,N_13694,N_13743);
xnor U13992 (N_13992,N_13543,N_13632);
xor U13993 (N_13993,N_13749,N_13504);
nor U13994 (N_13994,N_13527,N_13611);
xor U13995 (N_13995,N_13733,N_13598);
and U13996 (N_13996,N_13651,N_13548);
and U13997 (N_13997,N_13712,N_13688);
xor U13998 (N_13998,N_13559,N_13672);
nor U13999 (N_13999,N_13549,N_13584);
nor U14000 (N_14000,N_13975,N_13992);
nand U14001 (N_14001,N_13857,N_13783);
nand U14002 (N_14002,N_13972,N_13938);
and U14003 (N_14003,N_13912,N_13796);
nand U14004 (N_14004,N_13990,N_13988);
xor U14005 (N_14005,N_13757,N_13911);
nand U14006 (N_14006,N_13883,N_13995);
nor U14007 (N_14007,N_13895,N_13901);
and U14008 (N_14008,N_13773,N_13834);
xnor U14009 (N_14009,N_13921,N_13758);
xor U14010 (N_14010,N_13801,N_13944);
nor U14011 (N_14011,N_13900,N_13769);
or U14012 (N_14012,N_13787,N_13891);
nand U14013 (N_14013,N_13963,N_13851);
nand U14014 (N_14014,N_13937,N_13925);
nor U14015 (N_14015,N_13914,N_13767);
nor U14016 (N_14016,N_13752,N_13967);
nand U14017 (N_14017,N_13951,N_13952);
or U14018 (N_14018,N_13922,N_13755);
nor U14019 (N_14019,N_13751,N_13961);
nand U14020 (N_14020,N_13909,N_13887);
and U14021 (N_14021,N_13933,N_13780);
and U14022 (N_14022,N_13776,N_13807);
or U14023 (N_14023,N_13879,N_13794);
nor U14024 (N_14024,N_13945,N_13835);
and U14025 (N_14025,N_13955,N_13971);
or U14026 (N_14026,N_13763,N_13927);
or U14027 (N_14027,N_13765,N_13778);
and U14028 (N_14028,N_13840,N_13903);
xnor U14029 (N_14029,N_13991,N_13826);
xnor U14030 (N_14030,N_13997,N_13756);
nor U14031 (N_14031,N_13973,N_13848);
nor U14032 (N_14032,N_13885,N_13888);
nor U14033 (N_14033,N_13799,N_13941);
nor U14034 (N_14034,N_13978,N_13808);
nor U14035 (N_14035,N_13761,N_13790);
nor U14036 (N_14036,N_13868,N_13965);
nor U14037 (N_14037,N_13764,N_13797);
nand U14038 (N_14038,N_13788,N_13779);
nand U14039 (N_14039,N_13960,N_13999);
nor U14040 (N_14040,N_13828,N_13775);
nand U14041 (N_14041,N_13985,N_13817);
and U14042 (N_14042,N_13820,N_13917);
or U14043 (N_14043,N_13935,N_13760);
nor U14044 (N_14044,N_13898,N_13753);
nand U14045 (N_14045,N_13873,N_13754);
nand U14046 (N_14046,N_13982,N_13822);
nor U14047 (N_14047,N_13876,N_13860);
nor U14048 (N_14048,N_13994,N_13866);
and U14049 (N_14049,N_13855,N_13926);
and U14050 (N_14050,N_13913,N_13825);
or U14051 (N_14051,N_13789,N_13948);
nor U14052 (N_14052,N_13849,N_13907);
nor U14053 (N_14053,N_13814,N_13929);
nor U14054 (N_14054,N_13821,N_13812);
nand U14055 (N_14055,N_13934,N_13916);
xnor U14056 (N_14056,N_13894,N_13956);
xor U14057 (N_14057,N_13804,N_13844);
nand U14058 (N_14058,N_13806,N_13810);
xor U14059 (N_14059,N_13792,N_13953);
nor U14060 (N_14060,N_13892,N_13986);
nand U14061 (N_14061,N_13928,N_13939);
xnor U14062 (N_14062,N_13981,N_13899);
or U14063 (N_14063,N_13819,N_13993);
and U14064 (N_14064,N_13870,N_13896);
nor U14065 (N_14065,N_13932,N_13946);
and U14066 (N_14066,N_13877,N_13824);
or U14067 (N_14067,N_13793,N_13869);
xnor U14068 (N_14068,N_13839,N_13847);
and U14069 (N_14069,N_13947,N_13831);
nor U14070 (N_14070,N_13915,N_13750);
and U14071 (N_14071,N_13852,N_13987);
and U14072 (N_14072,N_13964,N_13970);
and U14073 (N_14073,N_13983,N_13800);
nor U14074 (N_14074,N_13998,N_13950);
nor U14075 (N_14075,N_13889,N_13818);
and U14076 (N_14076,N_13943,N_13781);
xnor U14077 (N_14077,N_13918,N_13864);
or U14078 (N_14078,N_13862,N_13803);
and U14079 (N_14079,N_13962,N_13786);
nand U14080 (N_14080,N_13874,N_13968);
nor U14081 (N_14081,N_13771,N_13798);
nor U14082 (N_14082,N_13897,N_13910);
xnor U14083 (N_14083,N_13853,N_13811);
and U14084 (N_14084,N_13777,N_13832);
nor U14085 (N_14085,N_13958,N_13930);
nor U14086 (N_14086,N_13957,N_13875);
nand U14087 (N_14087,N_13906,N_13871);
xor U14088 (N_14088,N_13774,N_13861);
nand U14089 (N_14089,N_13902,N_13845);
and U14090 (N_14090,N_13890,N_13886);
xnor U14091 (N_14091,N_13795,N_13836);
or U14092 (N_14092,N_13880,N_13977);
or U14093 (N_14093,N_13859,N_13949);
nor U14094 (N_14094,N_13989,N_13878);
nor U14095 (N_14095,N_13829,N_13863);
or U14096 (N_14096,N_13904,N_13816);
or U14097 (N_14097,N_13842,N_13846);
or U14098 (N_14098,N_13830,N_13805);
and U14099 (N_14099,N_13920,N_13770);
and U14100 (N_14100,N_13974,N_13768);
and U14101 (N_14101,N_13843,N_13827);
nor U14102 (N_14102,N_13850,N_13954);
or U14103 (N_14103,N_13791,N_13782);
and U14104 (N_14104,N_13837,N_13984);
and U14105 (N_14105,N_13802,N_13908);
and U14106 (N_14106,N_13959,N_13784);
or U14107 (N_14107,N_13766,N_13856);
xnor U14108 (N_14108,N_13919,N_13884);
and U14109 (N_14109,N_13841,N_13882);
nand U14110 (N_14110,N_13905,N_13854);
or U14111 (N_14111,N_13969,N_13940);
nor U14112 (N_14112,N_13923,N_13893);
nand U14113 (N_14113,N_13815,N_13980);
nor U14114 (N_14114,N_13881,N_13942);
and U14115 (N_14115,N_13809,N_13936);
nor U14116 (N_14116,N_13996,N_13867);
and U14117 (N_14117,N_13785,N_13966);
nand U14118 (N_14118,N_13813,N_13924);
or U14119 (N_14119,N_13762,N_13858);
nor U14120 (N_14120,N_13931,N_13772);
nor U14121 (N_14121,N_13833,N_13872);
and U14122 (N_14122,N_13976,N_13759);
and U14123 (N_14123,N_13823,N_13979);
nand U14124 (N_14124,N_13865,N_13838);
nor U14125 (N_14125,N_13868,N_13964);
or U14126 (N_14126,N_13970,N_13784);
and U14127 (N_14127,N_13933,N_13816);
xor U14128 (N_14128,N_13856,N_13777);
nor U14129 (N_14129,N_13806,N_13875);
nor U14130 (N_14130,N_13860,N_13772);
nor U14131 (N_14131,N_13904,N_13922);
or U14132 (N_14132,N_13878,N_13782);
and U14133 (N_14133,N_13773,N_13796);
xor U14134 (N_14134,N_13834,N_13928);
xor U14135 (N_14135,N_13805,N_13965);
or U14136 (N_14136,N_13858,N_13972);
nor U14137 (N_14137,N_13757,N_13829);
and U14138 (N_14138,N_13802,N_13753);
xor U14139 (N_14139,N_13883,N_13770);
nor U14140 (N_14140,N_13919,N_13936);
xnor U14141 (N_14141,N_13931,N_13751);
nand U14142 (N_14142,N_13812,N_13899);
and U14143 (N_14143,N_13870,N_13997);
nand U14144 (N_14144,N_13869,N_13972);
and U14145 (N_14145,N_13805,N_13754);
nor U14146 (N_14146,N_13947,N_13759);
or U14147 (N_14147,N_13870,N_13947);
nand U14148 (N_14148,N_13791,N_13803);
nand U14149 (N_14149,N_13883,N_13998);
nor U14150 (N_14150,N_13760,N_13877);
nand U14151 (N_14151,N_13880,N_13968);
and U14152 (N_14152,N_13837,N_13874);
nand U14153 (N_14153,N_13828,N_13797);
and U14154 (N_14154,N_13832,N_13929);
or U14155 (N_14155,N_13880,N_13992);
and U14156 (N_14156,N_13994,N_13757);
and U14157 (N_14157,N_13774,N_13762);
or U14158 (N_14158,N_13756,N_13884);
or U14159 (N_14159,N_13955,N_13952);
or U14160 (N_14160,N_13992,N_13819);
nor U14161 (N_14161,N_13990,N_13907);
nor U14162 (N_14162,N_13886,N_13781);
or U14163 (N_14163,N_13945,N_13801);
or U14164 (N_14164,N_13865,N_13913);
and U14165 (N_14165,N_13931,N_13944);
nor U14166 (N_14166,N_13775,N_13970);
nor U14167 (N_14167,N_13853,N_13838);
and U14168 (N_14168,N_13865,N_13999);
and U14169 (N_14169,N_13914,N_13812);
and U14170 (N_14170,N_13775,N_13830);
or U14171 (N_14171,N_13883,N_13786);
and U14172 (N_14172,N_13908,N_13925);
nand U14173 (N_14173,N_13999,N_13794);
or U14174 (N_14174,N_13844,N_13845);
and U14175 (N_14175,N_13870,N_13813);
nor U14176 (N_14176,N_13840,N_13782);
nand U14177 (N_14177,N_13928,N_13838);
nand U14178 (N_14178,N_13877,N_13954);
nor U14179 (N_14179,N_13941,N_13804);
nand U14180 (N_14180,N_13958,N_13921);
xor U14181 (N_14181,N_13818,N_13955);
and U14182 (N_14182,N_13845,N_13933);
and U14183 (N_14183,N_13787,N_13834);
nor U14184 (N_14184,N_13978,N_13895);
or U14185 (N_14185,N_13846,N_13794);
nand U14186 (N_14186,N_13971,N_13876);
or U14187 (N_14187,N_13765,N_13754);
and U14188 (N_14188,N_13850,N_13763);
or U14189 (N_14189,N_13946,N_13945);
or U14190 (N_14190,N_13857,N_13980);
or U14191 (N_14191,N_13896,N_13904);
nor U14192 (N_14192,N_13935,N_13818);
nand U14193 (N_14193,N_13906,N_13916);
nand U14194 (N_14194,N_13815,N_13854);
nor U14195 (N_14195,N_13840,N_13846);
nor U14196 (N_14196,N_13865,N_13978);
nor U14197 (N_14197,N_13897,N_13970);
nor U14198 (N_14198,N_13777,N_13920);
xor U14199 (N_14199,N_13946,N_13870);
nor U14200 (N_14200,N_13767,N_13996);
nor U14201 (N_14201,N_13917,N_13837);
nand U14202 (N_14202,N_13934,N_13981);
xor U14203 (N_14203,N_13869,N_13883);
nor U14204 (N_14204,N_13946,N_13807);
xnor U14205 (N_14205,N_13868,N_13985);
nand U14206 (N_14206,N_13817,N_13788);
nand U14207 (N_14207,N_13798,N_13979);
and U14208 (N_14208,N_13776,N_13917);
or U14209 (N_14209,N_13908,N_13986);
nand U14210 (N_14210,N_13933,N_13922);
xor U14211 (N_14211,N_13984,N_13847);
and U14212 (N_14212,N_13835,N_13885);
nor U14213 (N_14213,N_13981,N_13880);
or U14214 (N_14214,N_13942,N_13984);
nor U14215 (N_14215,N_13887,N_13972);
nor U14216 (N_14216,N_13901,N_13874);
and U14217 (N_14217,N_13928,N_13972);
nand U14218 (N_14218,N_13972,N_13965);
nand U14219 (N_14219,N_13899,N_13834);
or U14220 (N_14220,N_13866,N_13830);
and U14221 (N_14221,N_13863,N_13765);
or U14222 (N_14222,N_13927,N_13923);
xnor U14223 (N_14223,N_13903,N_13862);
and U14224 (N_14224,N_13903,N_13885);
nor U14225 (N_14225,N_13821,N_13998);
xor U14226 (N_14226,N_13975,N_13972);
or U14227 (N_14227,N_13876,N_13938);
and U14228 (N_14228,N_13905,N_13816);
or U14229 (N_14229,N_13784,N_13980);
or U14230 (N_14230,N_13764,N_13801);
nand U14231 (N_14231,N_13792,N_13976);
nand U14232 (N_14232,N_13854,N_13861);
nor U14233 (N_14233,N_13778,N_13835);
or U14234 (N_14234,N_13982,N_13944);
nand U14235 (N_14235,N_13889,N_13793);
or U14236 (N_14236,N_13934,N_13925);
or U14237 (N_14237,N_13967,N_13817);
or U14238 (N_14238,N_13963,N_13847);
xnor U14239 (N_14239,N_13975,N_13946);
or U14240 (N_14240,N_13918,N_13971);
nand U14241 (N_14241,N_13867,N_13917);
or U14242 (N_14242,N_13800,N_13988);
nand U14243 (N_14243,N_13907,N_13818);
nor U14244 (N_14244,N_13917,N_13949);
and U14245 (N_14245,N_13894,N_13883);
nand U14246 (N_14246,N_13963,N_13753);
nand U14247 (N_14247,N_13800,N_13763);
and U14248 (N_14248,N_13753,N_13982);
or U14249 (N_14249,N_13913,N_13784);
nand U14250 (N_14250,N_14068,N_14104);
nand U14251 (N_14251,N_14137,N_14151);
xnor U14252 (N_14252,N_14067,N_14059);
nand U14253 (N_14253,N_14192,N_14001);
nor U14254 (N_14254,N_14205,N_14027);
and U14255 (N_14255,N_14036,N_14159);
or U14256 (N_14256,N_14106,N_14008);
and U14257 (N_14257,N_14190,N_14145);
or U14258 (N_14258,N_14081,N_14219);
and U14259 (N_14259,N_14168,N_14167);
or U14260 (N_14260,N_14248,N_14209);
nand U14261 (N_14261,N_14127,N_14061);
or U14262 (N_14262,N_14017,N_14011);
or U14263 (N_14263,N_14118,N_14156);
nand U14264 (N_14264,N_14244,N_14089);
or U14265 (N_14265,N_14242,N_14110);
nor U14266 (N_14266,N_14009,N_14071);
nand U14267 (N_14267,N_14003,N_14014);
nand U14268 (N_14268,N_14088,N_14152);
nor U14269 (N_14269,N_14206,N_14176);
nor U14270 (N_14270,N_14047,N_14051);
or U14271 (N_14271,N_14235,N_14180);
nand U14272 (N_14272,N_14087,N_14117);
or U14273 (N_14273,N_14198,N_14125);
nor U14274 (N_14274,N_14130,N_14102);
nor U14275 (N_14275,N_14060,N_14232);
and U14276 (N_14276,N_14070,N_14173);
nand U14277 (N_14277,N_14218,N_14229);
nand U14278 (N_14278,N_14124,N_14058);
nand U14279 (N_14279,N_14210,N_14163);
and U14280 (N_14280,N_14141,N_14233);
nor U14281 (N_14281,N_14048,N_14193);
nand U14282 (N_14282,N_14121,N_14095);
nor U14283 (N_14283,N_14055,N_14054);
or U14284 (N_14284,N_14016,N_14230);
xor U14285 (N_14285,N_14085,N_14245);
and U14286 (N_14286,N_14107,N_14238);
or U14287 (N_14287,N_14021,N_14076);
nand U14288 (N_14288,N_14119,N_14039);
nor U14289 (N_14289,N_14032,N_14155);
xor U14290 (N_14290,N_14227,N_14084);
and U14291 (N_14291,N_14195,N_14090);
nand U14292 (N_14292,N_14083,N_14066);
nand U14293 (N_14293,N_14199,N_14220);
and U14294 (N_14294,N_14063,N_14188);
nand U14295 (N_14295,N_14174,N_14149);
nor U14296 (N_14296,N_14094,N_14018);
nor U14297 (N_14297,N_14128,N_14040);
or U14298 (N_14298,N_14221,N_14165);
and U14299 (N_14299,N_14170,N_14191);
xor U14300 (N_14300,N_14140,N_14042);
nor U14301 (N_14301,N_14237,N_14091);
and U14302 (N_14302,N_14216,N_14109);
nand U14303 (N_14303,N_14160,N_14114);
and U14304 (N_14304,N_14169,N_14241);
and U14305 (N_14305,N_14074,N_14101);
xor U14306 (N_14306,N_14052,N_14019);
nor U14307 (N_14307,N_14080,N_14236);
or U14308 (N_14308,N_14175,N_14208);
or U14309 (N_14309,N_14213,N_14143);
and U14310 (N_14310,N_14164,N_14171);
or U14311 (N_14311,N_14131,N_14093);
nor U14312 (N_14312,N_14225,N_14010);
nor U14313 (N_14313,N_14249,N_14029);
nand U14314 (N_14314,N_14082,N_14239);
or U14315 (N_14315,N_14126,N_14123);
or U14316 (N_14316,N_14187,N_14023);
xor U14317 (N_14317,N_14194,N_14065);
and U14318 (N_14318,N_14006,N_14207);
and U14319 (N_14319,N_14069,N_14211);
or U14320 (N_14320,N_14028,N_14035);
and U14321 (N_14321,N_14024,N_14183);
nand U14322 (N_14322,N_14079,N_14166);
nor U14323 (N_14323,N_14034,N_14002);
and U14324 (N_14324,N_14172,N_14142);
or U14325 (N_14325,N_14072,N_14184);
nand U14326 (N_14326,N_14108,N_14186);
xnor U14327 (N_14327,N_14154,N_14049);
or U14328 (N_14328,N_14147,N_14045);
nor U14329 (N_14329,N_14158,N_14038);
nor U14330 (N_14330,N_14030,N_14138);
nor U14331 (N_14331,N_14231,N_14135);
or U14332 (N_14332,N_14100,N_14077);
nand U14333 (N_14333,N_14223,N_14005);
xor U14334 (N_14334,N_14120,N_14112);
nand U14335 (N_14335,N_14200,N_14007);
xor U14336 (N_14336,N_14224,N_14243);
nand U14337 (N_14337,N_14073,N_14247);
or U14338 (N_14338,N_14111,N_14134);
and U14339 (N_14339,N_14132,N_14103);
nand U14340 (N_14340,N_14022,N_14004);
or U14341 (N_14341,N_14015,N_14092);
nor U14342 (N_14342,N_14098,N_14000);
or U14343 (N_14343,N_14215,N_14116);
nand U14344 (N_14344,N_14031,N_14056);
nor U14345 (N_14345,N_14204,N_14179);
and U14346 (N_14346,N_14115,N_14139);
xor U14347 (N_14347,N_14157,N_14240);
and U14348 (N_14348,N_14234,N_14129);
nand U14349 (N_14349,N_14122,N_14043);
or U14350 (N_14350,N_14214,N_14217);
nand U14351 (N_14351,N_14136,N_14178);
and U14352 (N_14352,N_14150,N_14148);
nand U14353 (N_14353,N_14013,N_14033);
and U14354 (N_14354,N_14097,N_14182);
nand U14355 (N_14355,N_14099,N_14096);
and U14356 (N_14356,N_14012,N_14105);
or U14357 (N_14357,N_14146,N_14203);
nor U14358 (N_14358,N_14113,N_14181);
nand U14359 (N_14359,N_14153,N_14086);
nand U14360 (N_14360,N_14046,N_14050);
nand U14361 (N_14361,N_14026,N_14162);
and U14362 (N_14362,N_14037,N_14246);
nand U14363 (N_14363,N_14185,N_14062);
and U14364 (N_14364,N_14075,N_14177);
and U14365 (N_14365,N_14222,N_14133);
nor U14366 (N_14366,N_14197,N_14212);
nor U14367 (N_14367,N_14078,N_14202);
nor U14368 (N_14368,N_14161,N_14226);
xnor U14369 (N_14369,N_14144,N_14053);
nand U14370 (N_14370,N_14228,N_14020);
nand U14371 (N_14371,N_14064,N_14201);
or U14372 (N_14372,N_14057,N_14196);
and U14373 (N_14373,N_14041,N_14189);
or U14374 (N_14374,N_14044,N_14025);
xnor U14375 (N_14375,N_14014,N_14155);
nor U14376 (N_14376,N_14034,N_14049);
nor U14377 (N_14377,N_14160,N_14067);
nand U14378 (N_14378,N_14060,N_14221);
or U14379 (N_14379,N_14054,N_14185);
nor U14380 (N_14380,N_14172,N_14044);
nor U14381 (N_14381,N_14066,N_14110);
nand U14382 (N_14382,N_14164,N_14138);
and U14383 (N_14383,N_14243,N_14138);
and U14384 (N_14384,N_14246,N_14027);
and U14385 (N_14385,N_14058,N_14015);
nand U14386 (N_14386,N_14233,N_14034);
nand U14387 (N_14387,N_14125,N_14249);
nor U14388 (N_14388,N_14231,N_14170);
nor U14389 (N_14389,N_14110,N_14181);
or U14390 (N_14390,N_14173,N_14168);
or U14391 (N_14391,N_14225,N_14187);
xor U14392 (N_14392,N_14143,N_14166);
or U14393 (N_14393,N_14122,N_14164);
and U14394 (N_14394,N_14216,N_14205);
or U14395 (N_14395,N_14013,N_14090);
nand U14396 (N_14396,N_14063,N_14230);
nor U14397 (N_14397,N_14194,N_14095);
and U14398 (N_14398,N_14129,N_14127);
nor U14399 (N_14399,N_14153,N_14094);
nor U14400 (N_14400,N_14103,N_14039);
or U14401 (N_14401,N_14049,N_14042);
or U14402 (N_14402,N_14097,N_14232);
nor U14403 (N_14403,N_14064,N_14223);
nand U14404 (N_14404,N_14192,N_14184);
xnor U14405 (N_14405,N_14025,N_14116);
nand U14406 (N_14406,N_14061,N_14186);
nand U14407 (N_14407,N_14018,N_14185);
and U14408 (N_14408,N_14191,N_14182);
xor U14409 (N_14409,N_14219,N_14073);
nand U14410 (N_14410,N_14053,N_14038);
nor U14411 (N_14411,N_14112,N_14154);
or U14412 (N_14412,N_14058,N_14177);
nand U14413 (N_14413,N_14224,N_14231);
and U14414 (N_14414,N_14230,N_14095);
or U14415 (N_14415,N_14151,N_14181);
nor U14416 (N_14416,N_14075,N_14069);
nand U14417 (N_14417,N_14200,N_14017);
nor U14418 (N_14418,N_14110,N_14057);
and U14419 (N_14419,N_14029,N_14175);
and U14420 (N_14420,N_14097,N_14093);
or U14421 (N_14421,N_14025,N_14228);
nor U14422 (N_14422,N_14169,N_14107);
nand U14423 (N_14423,N_14021,N_14114);
nor U14424 (N_14424,N_14050,N_14033);
nand U14425 (N_14425,N_14224,N_14022);
and U14426 (N_14426,N_14062,N_14144);
xor U14427 (N_14427,N_14099,N_14209);
or U14428 (N_14428,N_14031,N_14132);
and U14429 (N_14429,N_14162,N_14113);
and U14430 (N_14430,N_14214,N_14220);
nor U14431 (N_14431,N_14220,N_14058);
or U14432 (N_14432,N_14006,N_14018);
and U14433 (N_14433,N_14074,N_14133);
and U14434 (N_14434,N_14101,N_14177);
nand U14435 (N_14435,N_14201,N_14032);
nand U14436 (N_14436,N_14076,N_14136);
nor U14437 (N_14437,N_14244,N_14136);
and U14438 (N_14438,N_14230,N_14132);
nand U14439 (N_14439,N_14126,N_14170);
nor U14440 (N_14440,N_14239,N_14090);
and U14441 (N_14441,N_14161,N_14167);
nor U14442 (N_14442,N_14228,N_14059);
nor U14443 (N_14443,N_14240,N_14241);
nand U14444 (N_14444,N_14055,N_14134);
or U14445 (N_14445,N_14123,N_14028);
and U14446 (N_14446,N_14240,N_14046);
nand U14447 (N_14447,N_14053,N_14199);
and U14448 (N_14448,N_14122,N_14085);
nor U14449 (N_14449,N_14198,N_14179);
nor U14450 (N_14450,N_14236,N_14114);
xor U14451 (N_14451,N_14173,N_14228);
nand U14452 (N_14452,N_14215,N_14178);
nand U14453 (N_14453,N_14236,N_14215);
nand U14454 (N_14454,N_14047,N_14042);
and U14455 (N_14455,N_14148,N_14072);
nand U14456 (N_14456,N_14079,N_14180);
and U14457 (N_14457,N_14229,N_14053);
and U14458 (N_14458,N_14023,N_14072);
nand U14459 (N_14459,N_14029,N_14062);
nand U14460 (N_14460,N_14028,N_14218);
and U14461 (N_14461,N_14106,N_14050);
nand U14462 (N_14462,N_14007,N_14034);
or U14463 (N_14463,N_14088,N_14192);
nor U14464 (N_14464,N_14029,N_14026);
and U14465 (N_14465,N_14243,N_14150);
or U14466 (N_14466,N_14060,N_14134);
or U14467 (N_14467,N_14248,N_14033);
nand U14468 (N_14468,N_14138,N_14045);
and U14469 (N_14469,N_14159,N_14128);
and U14470 (N_14470,N_14075,N_14140);
or U14471 (N_14471,N_14160,N_14184);
xor U14472 (N_14472,N_14047,N_14124);
and U14473 (N_14473,N_14160,N_14201);
and U14474 (N_14474,N_14025,N_14163);
or U14475 (N_14475,N_14084,N_14212);
nand U14476 (N_14476,N_14239,N_14074);
nor U14477 (N_14477,N_14207,N_14094);
and U14478 (N_14478,N_14082,N_14151);
nand U14479 (N_14479,N_14134,N_14221);
nand U14480 (N_14480,N_14244,N_14094);
nor U14481 (N_14481,N_14212,N_14073);
nand U14482 (N_14482,N_14109,N_14125);
or U14483 (N_14483,N_14223,N_14149);
or U14484 (N_14484,N_14177,N_14180);
or U14485 (N_14485,N_14176,N_14163);
or U14486 (N_14486,N_14083,N_14135);
nor U14487 (N_14487,N_14067,N_14157);
or U14488 (N_14488,N_14238,N_14062);
nand U14489 (N_14489,N_14208,N_14029);
or U14490 (N_14490,N_14038,N_14187);
xor U14491 (N_14491,N_14033,N_14216);
and U14492 (N_14492,N_14180,N_14213);
and U14493 (N_14493,N_14014,N_14240);
or U14494 (N_14494,N_14142,N_14103);
nand U14495 (N_14495,N_14037,N_14098);
or U14496 (N_14496,N_14087,N_14016);
nor U14497 (N_14497,N_14236,N_14056);
and U14498 (N_14498,N_14030,N_14225);
nand U14499 (N_14499,N_14059,N_14142);
or U14500 (N_14500,N_14351,N_14492);
or U14501 (N_14501,N_14449,N_14400);
xnor U14502 (N_14502,N_14459,N_14486);
nand U14503 (N_14503,N_14323,N_14474);
nor U14504 (N_14504,N_14307,N_14484);
xnor U14505 (N_14505,N_14252,N_14301);
and U14506 (N_14506,N_14432,N_14457);
and U14507 (N_14507,N_14377,N_14298);
or U14508 (N_14508,N_14314,N_14493);
nor U14509 (N_14509,N_14430,N_14367);
nor U14510 (N_14510,N_14473,N_14409);
nor U14511 (N_14511,N_14332,N_14300);
nand U14512 (N_14512,N_14425,N_14448);
nand U14513 (N_14513,N_14406,N_14263);
nand U14514 (N_14514,N_14280,N_14465);
nand U14515 (N_14515,N_14353,N_14348);
and U14516 (N_14516,N_14397,N_14281);
nor U14517 (N_14517,N_14266,N_14347);
nand U14518 (N_14518,N_14345,N_14384);
nor U14519 (N_14519,N_14490,N_14331);
or U14520 (N_14520,N_14421,N_14309);
nor U14521 (N_14521,N_14335,N_14405);
and U14522 (N_14522,N_14402,N_14325);
nand U14523 (N_14523,N_14251,N_14466);
and U14524 (N_14524,N_14362,N_14291);
nand U14525 (N_14525,N_14338,N_14352);
or U14526 (N_14526,N_14462,N_14464);
or U14527 (N_14527,N_14398,N_14330);
or U14528 (N_14528,N_14388,N_14256);
or U14529 (N_14529,N_14297,N_14305);
nor U14530 (N_14530,N_14477,N_14413);
nand U14531 (N_14531,N_14364,N_14456);
xor U14532 (N_14532,N_14311,N_14316);
or U14533 (N_14533,N_14313,N_14283);
and U14534 (N_14534,N_14312,N_14343);
nor U14535 (N_14535,N_14373,N_14393);
nor U14536 (N_14536,N_14489,N_14470);
xor U14537 (N_14537,N_14395,N_14288);
nand U14538 (N_14538,N_14375,N_14411);
nor U14539 (N_14539,N_14420,N_14438);
and U14540 (N_14540,N_14417,N_14267);
or U14541 (N_14541,N_14404,N_14276);
or U14542 (N_14542,N_14328,N_14356);
xor U14543 (N_14543,N_14446,N_14317);
and U14544 (N_14544,N_14278,N_14396);
and U14545 (N_14545,N_14487,N_14419);
or U14546 (N_14546,N_14416,N_14381);
nor U14547 (N_14547,N_14382,N_14304);
or U14548 (N_14548,N_14467,N_14376);
or U14549 (N_14549,N_14357,N_14310);
or U14550 (N_14550,N_14275,N_14491);
or U14551 (N_14551,N_14440,N_14441);
or U14552 (N_14552,N_14392,N_14410);
or U14553 (N_14553,N_14320,N_14354);
nand U14554 (N_14554,N_14460,N_14431);
nor U14555 (N_14555,N_14424,N_14387);
nor U14556 (N_14556,N_14262,N_14269);
and U14557 (N_14557,N_14482,N_14483);
and U14558 (N_14558,N_14497,N_14469);
nor U14559 (N_14559,N_14401,N_14422);
and U14560 (N_14560,N_14293,N_14289);
nor U14561 (N_14561,N_14306,N_14445);
xor U14562 (N_14562,N_14260,N_14444);
xor U14563 (N_14563,N_14340,N_14250);
and U14564 (N_14564,N_14447,N_14268);
nand U14565 (N_14565,N_14368,N_14472);
nor U14566 (N_14566,N_14326,N_14321);
nand U14567 (N_14567,N_14333,N_14408);
nor U14568 (N_14568,N_14385,N_14427);
nor U14569 (N_14569,N_14350,N_14435);
nand U14570 (N_14570,N_14315,N_14264);
nor U14571 (N_14571,N_14294,N_14371);
nand U14572 (N_14572,N_14258,N_14471);
and U14573 (N_14573,N_14394,N_14443);
and U14574 (N_14574,N_14461,N_14339);
nor U14575 (N_14575,N_14407,N_14302);
nor U14576 (N_14576,N_14403,N_14324);
and U14577 (N_14577,N_14498,N_14277);
and U14578 (N_14578,N_14478,N_14257);
nand U14579 (N_14579,N_14481,N_14329);
nand U14580 (N_14580,N_14374,N_14423);
xnor U14581 (N_14581,N_14418,N_14284);
nor U14582 (N_14582,N_14355,N_14463);
nor U14583 (N_14583,N_14452,N_14454);
nand U14584 (N_14584,N_14414,N_14485);
or U14585 (N_14585,N_14412,N_14363);
or U14586 (N_14586,N_14499,N_14439);
nor U14587 (N_14587,N_14383,N_14265);
xnor U14588 (N_14588,N_14271,N_14475);
nor U14589 (N_14589,N_14327,N_14318);
nor U14590 (N_14590,N_14389,N_14366);
nand U14591 (N_14591,N_14319,N_14434);
and U14592 (N_14592,N_14496,N_14468);
nand U14593 (N_14593,N_14386,N_14286);
nor U14594 (N_14594,N_14322,N_14292);
nand U14595 (N_14595,N_14380,N_14295);
nor U14596 (N_14596,N_14337,N_14361);
nand U14597 (N_14597,N_14436,N_14372);
nand U14598 (N_14598,N_14272,N_14254);
nand U14599 (N_14599,N_14308,N_14426);
and U14600 (N_14600,N_14296,N_14341);
xor U14601 (N_14601,N_14342,N_14279);
nor U14602 (N_14602,N_14253,N_14458);
nand U14603 (N_14603,N_14450,N_14299);
or U14604 (N_14604,N_14399,N_14261);
nor U14605 (N_14605,N_14370,N_14290);
nor U14606 (N_14606,N_14391,N_14365);
and U14607 (N_14607,N_14259,N_14344);
nand U14608 (N_14608,N_14255,N_14451);
or U14609 (N_14609,N_14336,N_14479);
nand U14610 (N_14610,N_14360,N_14415);
and U14611 (N_14611,N_14442,N_14428);
nor U14612 (N_14612,N_14495,N_14429);
or U14613 (N_14613,N_14455,N_14303);
nand U14614 (N_14614,N_14480,N_14390);
or U14615 (N_14615,N_14369,N_14334);
nor U14616 (N_14616,N_14274,N_14488);
nor U14617 (N_14617,N_14453,N_14476);
xnor U14618 (N_14618,N_14358,N_14273);
and U14619 (N_14619,N_14359,N_14285);
and U14620 (N_14620,N_14270,N_14287);
and U14621 (N_14621,N_14433,N_14346);
or U14622 (N_14622,N_14349,N_14437);
nand U14623 (N_14623,N_14494,N_14378);
or U14624 (N_14624,N_14379,N_14282);
nand U14625 (N_14625,N_14355,N_14368);
nor U14626 (N_14626,N_14344,N_14411);
nand U14627 (N_14627,N_14272,N_14261);
xnor U14628 (N_14628,N_14477,N_14376);
or U14629 (N_14629,N_14253,N_14481);
xor U14630 (N_14630,N_14427,N_14270);
nor U14631 (N_14631,N_14277,N_14347);
nand U14632 (N_14632,N_14490,N_14380);
and U14633 (N_14633,N_14283,N_14276);
nor U14634 (N_14634,N_14350,N_14337);
or U14635 (N_14635,N_14424,N_14443);
nor U14636 (N_14636,N_14364,N_14370);
and U14637 (N_14637,N_14270,N_14388);
nor U14638 (N_14638,N_14354,N_14418);
and U14639 (N_14639,N_14485,N_14443);
or U14640 (N_14640,N_14355,N_14352);
and U14641 (N_14641,N_14281,N_14423);
or U14642 (N_14642,N_14402,N_14253);
and U14643 (N_14643,N_14288,N_14275);
nor U14644 (N_14644,N_14261,N_14336);
xnor U14645 (N_14645,N_14455,N_14492);
nand U14646 (N_14646,N_14255,N_14277);
nor U14647 (N_14647,N_14325,N_14365);
and U14648 (N_14648,N_14311,N_14279);
and U14649 (N_14649,N_14386,N_14381);
nand U14650 (N_14650,N_14440,N_14310);
xor U14651 (N_14651,N_14259,N_14413);
nand U14652 (N_14652,N_14315,N_14415);
nor U14653 (N_14653,N_14342,N_14265);
and U14654 (N_14654,N_14376,N_14294);
nand U14655 (N_14655,N_14426,N_14439);
nand U14656 (N_14656,N_14377,N_14344);
and U14657 (N_14657,N_14259,N_14428);
or U14658 (N_14658,N_14419,N_14489);
nand U14659 (N_14659,N_14251,N_14359);
xor U14660 (N_14660,N_14333,N_14362);
nand U14661 (N_14661,N_14269,N_14339);
nor U14662 (N_14662,N_14485,N_14353);
nor U14663 (N_14663,N_14308,N_14494);
nor U14664 (N_14664,N_14315,N_14423);
or U14665 (N_14665,N_14264,N_14493);
nand U14666 (N_14666,N_14450,N_14449);
nor U14667 (N_14667,N_14275,N_14407);
and U14668 (N_14668,N_14453,N_14298);
or U14669 (N_14669,N_14333,N_14260);
nand U14670 (N_14670,N_14458,N_14395);
nor U14671 (N_14671,N_14399,N_14393);
and U14672 (N_14672,N_14309,N_14482);
nor U14673 (N_14673,N_14267,N_14458);
nand U14674 (N_14674,N_14357,N_14412);
nor U14675 (N_14675,N_14353,N_14301);
nor U14676 (N_14676,N_14283,N_14330);
nand U14677 (N_14677,N_14342,N_14263);
and U14678 (N_14678,N_14280,N_14279);
and U14679 (N_14679,N_14436,N_14490);
and U14680 (N_14680,N_14433,N_14327);
nor U14681 (N_14681,N_14423,N_14437);
nor U14682 (N_14682,N_14424,N_14323);
and U14683 (N_14683,N_14336,N_14464);
nor U14684 (N_14684,N_14370,N_14276);
nor U14685 (N_14685,N_14315,N_14364);
and U14686 (N_14686,N_14320,N_14263);
or U14687 (N_14687,N_14294,N_14317);
xnor U14688 (N_14688,N_14351,N_14411);
or U14689 (N_14689,N_14425,N_14285);
or U14690 (N_14690,N_14338,N_14374);
nor U14691 (N_14691,N_14497,N_14433);
nor U14692 (N_14692,N_14495,N_14435);
nor U14693 (N_14693,N_14372,N_14396);
nor U14694 (N_14694,N_14381,N_14441);
and U14695 (N_14695,N_14289,N_14335);
nor U14696 (N_14696,N_14382,N_14452);
nand U14697 (N_14697,N_14335,N_14384);
nand U14698 (N_14698,N_14313,N_14277);
nand U14699 (N_14699,N_14383,N_14254);
nor U14700 (N_14700,N_14416,N_14264);
or U14701 (N_14701,N_14349,N_14359);
xor U14702 (N_14702,N_14455,N_14477);
and U14703 (N_14703,N_14398,N_14493);
and U14704 (N_14704,N_14428,N_14436);
nor U14705 (N_14705,N_14467,N_14313);
nor U14706 (N_14706,N_14337,N_14490);
nor U14707 (N_14707,N_14383,N_14317);
or U14708 (N_14708,N_14315,N_14474);
and U14709 (N_14709,N_14473,N_14415);
nand U14710 (N_14710,N_14332,N_14453);
nand U14711 (N_14711,N_14389,N_14327);
nor U14712 (N_14712,N_14314,N_14362);
nand U14713 (N_14713,N_14426,N_14436);
nand U14714 (N_14714,N_14465,N_14419);
nand U14715 (N_14715,N_14427,N_14340);
and U14716 (N_14716,N_14433,N_14284);
or U14717 (N_14717,N_14470,N_14407);
and U14718 (N_14718,N_14296,N_14251);
and U14719 (N_14719,N_14254,N_14334);
nand U14720 (N_14720,N_14254,N_14368);
and U14721 (N_14721,N_14385,N_14382);
nor U14722 (N_14722,N_14258,N_14381);
or U14723 (N_14723,N_14493,N_14326);
nor U14724 (N_14724,N_14395,N_14388);
nor U14725 (N_14725,N_14368,N_14284);
or U14726 (N_14726,N_14272,N_14398);
nor U14727 (N_14727,N_14328,N_14452);
nor U14728 (N_14728,N_14329,N_14352);
and U14729 (N_14729,N_14445,N_14430);
xnor U14730 (N_14730,N_14368,N_14334);
and U14731 (N_14731,N_14478,N_14298);
xnor U14732 (N_14732,N_14332,N_14255);
xnor U14733 (N_14733,N_14415,N_14486);
or U14734 (N_14734,N_14254,N_14263);
and U14735 (N_14735,N_14361,N_14413);
nor U14736 (N_14736,N_14308,N_14471);
nand U14737 (N_14737,N_14268,N_14291);
and U14738 (N_14738,N_14469,N_14369);
or U14739 (N_14739,N_14290,N_14449);
nor U14740 (N_14740,N_14345,N_14420);
nand U14741 (N_14741,N_14479,N_14470);
xor U14742 (N_14742,N_14447,N_14392);
or U14743 (N_14743,N_14412,N_14419);
nand U14744 (N_14744,N_14431,N_14323);
nand U14745 (N_14745,N_14410,N_14403);
and U14746 (N_14746,N_14362,N_14499);
xor U14747 (N_14747,N_14495,N_14344);
nand U14748 (N_14748,N_14468,N_14352);
or U14749 (N_14749,N_14458,N_14292);
nand U14750 (N_14750,N_14638,N_14643);
or U14751 (N_14751,N_14724,N_14618);
and U14752 (N_14752,N_14529,N_14575);
nand U14753 (N_14753,N_14504,N_14501);
nand U14754 (N_14754,N_14708,N_14702);
and U14755 (N_14755,N_14635,N_14599);
xnor U14756 (N_14756,N_14566,N_14515);
or U14757 (N_14757,N_14502,N_14676);
xor U14758 (N_14758,N_14695,N_14598);
xor U14759 (N_14759,N_14737,N_14668);
nand U14760 (N_14760,N_14659,N_14713);
or U14761 (N_14761,N_14611,N_14583);
and U14762 (N_14762,N_14694,N_14650);
and U14763 (N_14763,N_14621,N_14662);
nor U14764 (N_14764,N_14661,N_14619);
nor U14765 (N_14765,N_14608,N_14538);
xor U14766 (N_14766,N_14574,N_14547);
and U14767 (N_14767,N_14640,N_14688);
nor U14768 (N_14768,N_14548,N_14564);
nor U14769 (N_14769,N_14701,N_14532);
or U14770 (N_14770,N_14531,N_14627);
and U14771 (N_14771,N_14579,N_14645);
xor U14772 (N_14772,N_14723,N_14506);
nand U14773 (N_14773,N_14717,N_14649);
or U14774 (N_14774,N_14587,N_14572);
or U14775 (N_14775,N_14663,N_14729);
and U14776 (N_14776,N_14542,N_14620);
or U14777 (N_14777,N_14716,N_14656);
and U14778 (N_14778,N_14686,N_14591);
nand U14779 (N_14779,N_14639,N_14703);
nor U14780 (N_14780,N_14610,N_14581);
xnor U14781 (N_14781,N_14540,N_14647);
and U14782 (N_14782,N_14633,N_14578);
nor U14783 (N_14783,N_14609,N_14636);
nor U14784 (N_14784,N_14570,N_14519);
or U14785 (N_14785,N_14617,N_14550);
and U14786 (N_14786,N_14730,N_14614);
or U14787 (N_14787,N_14705,N_14718);
and U14788 (N_14788,N_14657,N_14562);
nand U14789 (N_14789,N_14732,N_14741);
or U14790 (N_14790,N_14521,N_14655);
xnor U14791 (N_14791,N_14526,N_14704);
or U14792 (N_14792,N_14664,N_14685);
nor U14793 (N_14793,N_14692,N_14584);
and U14794 (N_14794,N_14518,N_14670);
and U14795 (N_14795,N_14556,N_14585);
and U14796 (N_14796,N_14597,N_14660);
and U14797 (N_14797,N_14600,N_14697);
xnor U14798 (N_14798,N_14545,N_14699);
nor U14799 (N_14799,N_14747,N_14536);
or U14800 (N_14800,N_14721,N_14571);
or U14801 (N_14801,N_14543,N_14679);
nand U14802 (N_14802,N_14646,N_14700);
or U14803 (N_14803,N_14561,N_14606);
nand U14804 (N_14804,N_14588,N_14528);
xnor U14805 (N_14805,N_14565,N_14641);
nor U14806 (N_14806,N_14742,N_14744);
or U14807 (N_14807,N_14678,N_14553);
nor U14808 (N_14808,N_14652,N_14714);
nand U14809 (N_14809,N_14514,N_14669);
xor U14810 (N_14810,N_14625,N_14593);
nand U14811 (N_14811,N_14637,N_14644);
nor U14812 (N_14812,N_14552,N_14706);
xor U14813 (N_14813,N_14616,N_14707);
or U14814 (N_14814,N_14672,N_14623);
and U14815 (N_14815,N_14537,N_14563);
nand U14816 (N_14816,N_14541,N_14683);
nand U14817 (N_14817,N_14677,N_14507);
or U14818 (N_14818,N_14690,N_14634);
xnor U14819 (N_14819,N_14734,N_14624);
and U14820 (N_14820,N_14733,N_14533);
nor U14821 (N_14821,N_14601,N_14689);
xor U14822 (N_14822,N_14727,N_14568);
and U14823 (N_14823,N_14651,N_14712);
and U14824 (N_14824,N_14500,N_14726);
or U14825 (N_14825,N_14505,N_14691);
or U14826 (N_14826,N_14512,N_14569);
nor U14827 (N_14827,N_14632,N_14749);
nor U14828 (N_14828,N_14551,N_14510);
nand U14829 (N_14829,N_14687,N_14513);
nand U14830 (N_14830,N_14648,N_14527);
nand U14831 (N_14831,N_14602,N_14693);
and U14832 (N_14832,N_14674,N_14508);
nand U14833 (N_14833,N_14654,N_14503);
nand U14834 (N_14834,N_14534,N_14516);
nand U14835 (N_14835,N_14509,N_14546);
or U14836 (N_14836,N_14740,N_14719);
xnor U14837 (N_14837,N_14517,N_14560);
nand U14838 (N_14838,N_14653,N_14525);
nand U14839 (N_14839,N_14539,N_14582);
nor U14840 (N_14840,N_14671,N_14595);
nand U14841 (N_14841,N_14681,N_14696);
or U14842 (N_14842,N_14520,N_14715);
xnor U14843 (N_14843,N_14586,N_14522);
and U14844 (N_14844,N_14665,N_14630);
nor U14845 (N_14845,N_14736,N_14680);
or U14846 (N_14846,N_14710,N_14615);
nor U14847 (N_14847,N_14605,N_14622);
and U14848 (N_14848,N_14555,N_14631);
or U14849 (N_14849,N_14612,N_14739);
nand U14850 (N_14850,N_14666,N_14675);
and U14851 (N_14851,N_14567,N_14554);
and U14852 (N_14852,N_14511,N_14684);
nor U14853 (N_14853,N_14682,N_14642);
nor U14854 (N_14854,N_14604,N_14592);
nor U14855 (N_14855,N_14549,N_14735);
or U14856 (N_14856,N_14629,N_14607);
and U14857 (N_14857,N_14667,N_14728);
or U14858 (N_14858,N_14613,N_14577);
xnor U14859 (N_14859,N_14589,N_14580);
nor U14860 (N_14860,N_14558,N_14745);
or U14861 (N_14861,N_14720,N_14746);
or U14862 (N_14862,N_14673,N_14557);
and U14863 (N_14863,N_14573,N_14594);
nand U14864 (N_14864,N_14626,N_14544);
nand U14865 (N_14865,N_14524,N_14722);
nor U14866 (N_14866,N_14535,N_14711);
and U14867 (N_14867,N_14530,N_14590);
and U14868 (N_14868,N_14709,N_14596);
and U14869 (N_14869,N_14603,N_14559);
and U14870 (N_14870,N_14748,N_14738);
nand U14871 (N_14871,N_14725,N_14523);
or U14872 (N_14872,N_14658,N_14698);
nand U14873 (N_14873,N_14743,N_14628);
nand U14874 (N_14874,N_14576,N_14731);
nand U14875 (N_14875,N_14570,N_14586);
nor U14876 (N_14876,N_14572,N_14515);
nand U14877 (N_14877,N_14724,N_14616);
or U14878 (N_14878,N_14603,N_14685);
nand U14879 (N_14879,N_14552,N_14532);
nor U14880 (N_14880,N_14602,N_14673);
nand U14881 (N_14881,N_14718,N_14608);
nand U14882 (N_14882,N_14745,N_14700);
or U14883 (N_14883,N_14677,N_14565);
and U14884 (N_14884,N_14579,N_14641);
and U14885 (N_14885,N_14550,N_14749);
or U14886 (N_14886,N_14524,N_14732);
xor U14887 (N_14887,N_14588,N_14671);
and U14888 (N_14888,N_14655,N_14558);
or U14889 (N_14889,N_14745,N_14513);
and U14890 (N_14890,N_14519,N_14615);
and U14891 (N_14891,N_14738,N_14678);
and U14892 (N_14892,N_14609,N_14543);
and U14893 (N_14893,N_14695,N_14660);
and U14894 (N_14894,N_14628,N_14737);
nand U14895 (N_14895,N_14687,N_14675);
or U14896 (N_14896,N_14686,N_14521);
nor U14897 (N_14897,N_14526,N_14514);
nand U14898 (N_14898,N_14689,N_14714);
nor U14899 (N_14899,N_14650,N_14537);
and U14900 (N_14900,N_14556,N_14746);
nor U14901 (N_14901,N_14663,N_14576);
xor U14902 (N_14902,N_14670,N_14568);
and U14903 (N_14903,N_14629,N_14558);
xnor U14904 (N_14904,N_14685,N_14628);
or U14905 (N_14905,N_14658,N_14592);
or U14906 (N_14906,N_14579,N_14607);
nand U14907 (N_14907,N_14664,N_14665);
and U14908 (N_14908,N_14614,N_14665);
or U14909 (N_14909,N_14620,N_14556);
and U14910 (N_14910,N_14514,N_14668);
xor U14911 (N_14911,N_14651,N_14559);
nor U14912 (N_14912,N_14723,N_14526);
and U14913 (N_14913,N_14728,N_14696);
and U14914 (N_14914,N_14745,N_14626);
xor U14915 (N_14915,N_14517,N_14711);
and U14916 (N_14916,N_14661,N_14687);
and U14917 (N_14917,N_14689,N_14561);
or U14918 (N_14918,N_14610,N_14643);
nor U14919 (N_14919,N_14556,N_14530);
nor U14920 (N_14920,N_14737,N_14654);
nand U14921 (N_14921,N_14744,N_14683);
nor U14922 (N_14922,N_14632,N_14511);
nor U14923 (N_14923,N_14693,N_14735);
nor U14924 (N_14924,N_14513,N_14599);
or U14925 (N_14925,N_14582,N_14748);
or U14926 (N_14926,N_14674,N_14519);
or U14927 (N_14927,N_14641,N_14668);
nand U14928 (N_14928,N_14740,N_14567);
or U14929 (N_14929,N_14542,N_14543);
or U14930 (N_14930,N_14674,N_14615);
nand U14931 (N_14931,N_14625,N_14587);
or U14932 (N_14932,N_14509,N_14705);
nor U14933 (N_14933,N_14542,N_14525);
nor U14934 (N_14934,N_14696,N_14524);
and U14935 (N_14935,N_14550,N_14579);
and U14936 (N_14936,N_14742,N_14694);
nand U14937 (N_14937,N_14654,N_14656);
nand U14938 (N_14938,N_14665,N_14538);
and U14939 (N_14939,N_14549,N_14649);
nand U14940 (N_14940,N_14580,N_14632);
and U14941 (N_14941,N_14654,N_14554);
nand U14942 (N_14942,N_14615,N_14668);
xnor U14943 (N_14943,N_14550,N_14583);
and U14944 (N_14944,N_14614,N_14623);
and U14945 (N_14945,N_14713,N_14509);
or U14946 (N_14946,N_14575,N_14510);
xor U14947 (N_14947,N_14652,N_14731);
and U14948 (N_14948,N_14549,N_14563);
nor U14949 (N_14949,N_14518,N_14579);
nand U14950 (N_14950,N_14738,N_14559);
or U14951 (N_14951,N_14537,N_14697);
xnor U14952 (N_14952,N_14727,N_14572);
and U14953 (N_14953,N_14567,N_14576);
xnor U14954 (N_14954,N_14549,N_14691);
nor U14955 (N_14955,N_14642,N_14748);
nand U14956 (N_14956,N_14675,N_14526);
nand U14957 (N_14957,N_14633,N_14536);
or U14958 (N_14958,N_14581,N_14593);
and U14959 (N_14959,N_14634,N_14721);
nand U14960 (N_14960,N_14697,N_14553);
nand U14961 (N_14961,N_14693,N_14678);
nor U14962 (N_14962,N_14593,N_14616);
and U14963 (N_14963,N_14658,N_14510);
and U14964 (N_14964,N_14623,N_14604);
or U14965 (N_14965,N_14601,N_14598);
and U14966 (N_14966,N_14572,N_14579);
xor U14967 (N_14967,N_14709,N_14688);
nor U14968 (N_14968,N_14516,N_14635);
or U14969 (N_14969,N_14561,N_14747);
or U14970 (N_14970,N_14649,N_14742);
and U14971 (N_14971,N_14660,N_14725);
nand U14972 (N_14972,N_14589,N_14552);
nor U14973 (N_14973,N_14721,N_14580);
nor U14974 (N_14974,N_14710,N_14652);
or U14975 (N_14975,N_14665,N_14672);
and U14976 (N_14976,N_14534,N_14539);
nand U14977 (N_14977,N_14504,N_14603);
nand U14978 (N_14978,N_14677,N_14504);
and U14979 (N_14979,N_14566,N_14603);
or U14980 (N_14980,N_14710,N_14669);
and U14981 (N_14981,N_14655,N_14728);
nand U14982 (N_14982,N_14569,N_14628);
or U14983 (N_14983,N_14567,N_14744);
nand U14984 (N_14984,N_14502,N_14724);
or U14985 (N_14985,N_14519,N_14549);
and U14986 (N_14986,N_14543,N_14562);
nand U14987 (N_14987,N_14590,N_14553);
and U14988 (N_14988,N_14724,N_14705);
nor U14989 (N_14989,N_14620,N_14629);
or U14990 (N_14990,N_14663,N_14582);
and U14991 (N_14991,N_14700,N_14722);
nor U14992 (N_14992,N_14553,N_14568);
or U14993 (N_14993,N_14555,N_14615);
nor U14994 (N_14994,N_14542,N_14721);
nand U14995 (N_14995,N_14640,N_14610);
nor U14996 (N_14996,N_14697,N_14671);
nor U14997 (N_14997,N_14544,N_14735);
nand U14998 (N_14998,N_14504,N_14576);
nand U14999 (N_14999,N_14551,N_14684);
nand UO_0 (O_0,N_14774,N_14820);
nor UO_1 (O_1,N_14880,N_14796);
and UO_2 (O_2,N_14948,N_14860);
nand UO_3 (O_3,N_14910,N_14781);
nor UO_4 (O_4,N_14929,N_14998);
or UO_5 (O_5,N_14761,N_14772);
and UO_6 (O_6,N_14976,N_14852);
or UO_7 (O_7,N_14791,N_14927);
nor UO_8 (O_8,N_14865,N_14939);
and UO_9 (O_9,N_14775,N_14858);
and UO_10 (O_10,N_14978,N_14845);
nor UO_11 (O_11,N_14918,N_14794);
or UO_12 (O_12,N_14790,N_14798);
and UO_13 (O_13,N_14834,N_14766);
nor UO_14 (O_14,N_14871,N_14801);
or UO_15 (O_15,N_14991,N_14968);
nor UO_16 (O_16,N_14993,N_14851);
nand UO_17 (O_17,N_14779,N_14967);
nor UO_18 (O_18,N_14862,N_14857);
nor UO_19 (O_19,N_14827,N_14872);
and UO_20 (O_20,N_14830,N_14979);
nor UO_21 (O_21,N_14934,N_14797);
nand UO_22 (O_22,N_14981,N_14988);
or UO_23 (O_23,N_14756,N_14789);
or UO_24 (O_24,N_14821,N_14754);
nor UO_25 (O_25,N_14914,N_14917);
nor UO_26 (O_26,N_14908,N_14881);
and UO_27 (O_27,N_14937,N_14949);
or UO_28 (O_28,N_14894,N_14902);
nor UO_29 (O_29,N_14780,N_14760);
and UO_30 (O_30,N_14837,N_14888);
xor UO_31 (O_31,N_14813,N_14767);
nor UO_32 (O_32,N_14977,N_14853);
nor UO_33 (O_33,N_14926,N_14973);
nor UO_34 (O_34,N_14953,N_14861);
xor UO_35 (O_35,N_14793,N_14825);
xnor UO_36 (O_36,N_14900,N_14833);
and UO_37 (O_37,N_14922,N_14757);
and UO_38 (O_38,N_14759,N_14810);
or UO_39 (O_39,N_14884,N_14816);
nor UO_40 (O_40,N_14933,N_14782);
and UO_41 (O_41,N_14987,N_14863);
nand UO_42 (O_42,N_14906,N_14975);
nor UO_43 (O_43,N_14959,N_14818);
nand UO_44 (O_44,N_14985,N_14885);
nor UO_45 (O_45,N_14951,N_14905);
nand UO_46 (O_46,N_14855,N_14964);
xor UO_47 (O_47,N_14940,N_14765);
xor UO_48 (O_48,N_14963,N_14823);
nor UO_49 (O_49,N_14836,N_14764);
nor UO_50 (O_50,N_14969,N_14913);
or UO_51 (O_51,N_14895,N_14824);
nor UO_52 (O_52,N_14778,N_14792);
and UO_53 (O_53,N_14974,N_14971);
and UO_54 (O_54,N_14962,N_14912);
nand UO_55 (O_55,N_14864,N_14904);
nor UO_56 (O_56,N_14955,N_14751);
xnor UO_57 (O_57,N_14995,N_14989);
and UO_58 (O_58,N_14839,N_14891);
nand UO_59 (O_59,N_14999,N_14986);
xor UO_60 (O_60,N_14923,N_14965);
xor UO_61 (O_61,N_14882,N_14842);
nand UO_62 (O_62,N_14808,N_14920);
nand UO_63 (O_63,N_14903,N_14982);
and UO_64 (O_64,N_14755,N_14758);
and UO_65 (O_65,N_14896,N_14809);
nand UO_66 (O_66,N_14786,N_14915);
nand UO_67 (O_67,N_14930,N_14856);
or UO_68 (O_68,N_14887,N_14826);
or UO_69 (O_69,N_14784,N_14938);
or UO_70 (O_70,N_14773,N_14990);
and UO_71 (O_71,N_14840,N_14960);
nor UO_72 (O_72,N_14936,N_14867);
nand UO_73 (O_73,N_14983,N_14907);
and UO_74 (O_74,N_14957,N_14901);
and UO_75 (O_75,N_14768,N_14835);
and UO_76 (O_76,N_14970,N_14807);
and UO_77 (O_77,N_14846,N_14817);
or UO_78 (O_78,N_14890,N_14802);
nand UO_79 (O_79,N_14879,N_14873);
and UO_80 (O_80,N_14805,N_14925);
nand UO_81 (O_81,N_14946,N_14942);
and UO_82 (O_82,N_14919,N_14803);
nand UO_83 (O_83,N_14777,N_14994);
nor UO_84 (O_84,N_14889,N_14935);
or UO_85 (O_85,N_14877,N_14752);
nand UO_86 (O_86,N_14961,N_14868);
or UO_87 (O_87,N_14753,N_14776);
nor UO_88 (O_88,N_14893,N_14812);
nand UO_89 (O_89,N_14844,N_14956);
and UO_90 (O_90,N_14952,N_14771);
nand UO_91 (O_91,N_14980,N_14931);
nor UO_92 (O_92,N_14762,N_14941);
nand UO_93 (O_93,N_14854,N_14932);
nand UO_94 (O_94,N_14996,N_14875);
and UO_95 (O_95,N_14831,N_14829);
or UO_96 (O_96,N_14832,N_14876);
nor UO_97 (O_97,N_14997,N_14770);
nor UO_98 (O_98,N_14819,N_14870);
or UO_99 (O_99,N_14966,N_14921);
and UO_100 (O_100,N_14795,N_14947);
and UO_101 (O_101,N_14769,N_14814);
and UO_102 (O_102,N_14763,N_14787);
or UO_103 (O_103,N_14897,N_14899);
and UO_104 (O_104,N_14944,N_14849);
or UO_105 (O_105,N_14886,N_14958);
xnor UO_106 (O_106,N_14909,N_14841);
or UO_107 (O_107,N_14878,N_14799);
nand UO_108 (O_108,N_14800,N_14911);
nand UO_109 (O_109,N_14866,N_14848);
nor UO_110 (O_110,N_14950,N_14806);
nor UO_111 (O_111,N_14972,N_14850);
nor UO_112 (O_112,N_14750,N_14838);
and UO_113 (O_113,N_14859,N_14916);
nand UO_114 (O_114,N_14822,N_14928);
nand UO_115 (O_115,N_14874,N_14828);
nand UO_116 (O_116,N_14883,N_14892);
nand UO_117 (O_117,N_14785,N_14804);
or UO_118 (O_118,N_14815,N_14898);
nand UO_119 (O_119,N_14945,N_14788);
xor UO_120 (O_120,N_14847,N_14992);
nand UO_121 (O_121,N_14869,N_14811);
nand UO_122 (O_122,N_14783,N_14954);
xor UO_123 (O_123,N_14924,N_14984);
or UO_124 (O_124,N_14943,N_14843);
or UO_125 (O_125,N_14942,N_14850);
and UO_126 (O_126,N_14925,N_14848);
nand UO_127 (O_127,N_14933,N_14843);
nor UO_128 (O_128,N_14859,N_14889);
and UO_129 (O_129,N_14911,N_14846);
and UO_130 (O_130,N_14935,N_14954);
xnor UO_131 (O_131,N_14784,N_14816);
and UO_132 (O_132,N_14868,N_14836);
nand UO_133 (O_133,N_14987,N_14803);
nand UO_134 (O_134,N_14906,N_14957);
and UO_135 (O_135,N_14936,N_14888);
or UO_136 (O_136,N_14829,N_14763);
nor UO_137 (O_137,N_14919,N_14774);
nor UO_138 (O_138,N_14965,N_14824);
nor UO_139 (O_139,N_14772,N_14969);
and UO_140 (O_140,N_14899,N_14853);
and UO_141 (O_141,N_14850,N_14789);
or UO_142 (O_142,N_14861,N_14791);
nand UO_143 (O_143,N_14845,N_14959);
or UO_144 (O_144,N_14973,N_14910);
nor UO_145 (O_145,N_14761,N_14951);
xor UO_146 (O_146,N_14861,N_14883);
and UO_147 (O_147,N_14831,N_14818);
and UO_148 (O_148,N_14871,N_14772);
nand UO_149 (O_149,N_14876,N_14955);
nand UO_150 (O_150,N_14898,N_14848);
nor UO_151 (O_151,N_14876,N_14840);
xnor UO_152 (O_152,N_14886,N_14770);
nor UO_153 (O_153,N_14772,N_14904);
and UO_154 (O_154,N_14910,N_14828);
or UO_155 (O_155,N_14838,N_14977);
nor UO_156 (O_156,N_14896,N_14988);
and UO_157 (O_157,N_14996,N_14871);
xnor UO_158 (O_158,N_14803,N_14854);
nand UO_159 (O_159,N_14908,N_14922);
or UO_160 (O_160,N_14762,N_14952);
nor UO_161 (O_161,N_14938,N_14956);
nor UO_162 (O_162,N_14800,N_14766);
or UO_163 (O_163,N_14778,N_14800);
nor UO_164 (O_164,N_14995,N_14984);
nand UO_165 (O_165,N_14875,N_14881);
nor UO_166 (O_166,N_14941,N_14922);
nand UO_167 (O_167,N_14986,N_14935);
or UO_168 (O_168,N_14974,N_14808);
nor UO_169 (O_169,N_14882,N_14850);
or UO_170 (O_170,N_14762,N_14964);
and UO_171 (O_171,N_14813,N_14800);
nor UO_172 (O_172,N_14962,N_14989);
or UO_173 (O_173,N_14913,N_14915);
nor UO_174 (O_174,N_14880,N_14773);
nor UO_175 (O_175,N_14806,N_14947);
or UO_176 (O_176,N_14873,N_14862);
nand UO_177 (O_177,N_14863,N_14856);
nand UO_178 (O_178,N_14834,N_14838);
nand UO_179 (O_179,N_14954,N_14972);
or UO_180 (O_180,N_14836,N_14996);
nor UO_181 (O_181,N_14775,N_14920);
nand UO_182 (O_182,N_14829,N_14875);
or UO_183 (O_183,N_14922,N_14774);
nand UO_184 (O_184,N_14988,N_14989);
and UO_185 (O_185,N_14852,N_14813);
and UO_186 (O_186,N_14828,N_14963);
nor UO_187 (O_187,N_14806,N_14996);
or UO_188 (O_188,N_14767,N_14838);
nand UO_189 (O_189,N_14956,N_14900);
or UO_190 (O_190,N_14880,N_14867);
or UO_191 (O_191,N_14939,N_14944);
or UO_192 (O_192,N_14940,N_14784);
nor UO_193 (O_193,N_14758,N_14961);
or UO_194 (O_194,N_14990,N_14952);
nor UO_195 (O_195,N_14894,N_14913);
or UO_196 (O_196,N_14993,N_14902);
and UO_197 (O_197,N_14994,N_14787);
nor UO_198 (O_198,N_14995,N_14853);
or UO_199 (O_199,N_14803,N_14763);
or UO_200 (O_200,N_14831,N_14869);
and UO_201 (O_201,N_14926,N_14863);
nor UO_202 (O_202,N_14958,N_14792);
nand UO_203 (O_203,N_14859,N_14876);
nand UO_204 (O_204,N_14762,N_14855);
nor UO_205 (O_205,N_14849,N_14837);
and UO_206 (O_206,N_14969,N_14751);
nand UO_207 (O_207,N_14958,N_14941);
nor UO_208 (O_208,N_14922,N_14784);
or UO_209 (O_209,N_14960,N_14874);
and UO_210 (O_210,N_14916,N_14781);
or UO_211 (O_211,N_14909,N_14788);
nor UO_212 (O_212,N_14964,N_14997);
nand UO_213 (O_213,N_14983,N_14758);
or UO_214 (O_214,N_14966,N_14916);
nand UO_215 (O_215,N_14825,N_14914);
nand UO_216 (O_216,N_14788,N_14760);
and UO_217 (O_217,N_14989,N_14755);
or UO_218 (O_218,N_14811,N_14815);
xor UO_219 (O_219,N_14793,N_14846);
and UO_220 (O_220,N_14816,N_14833);
nor UO_221 (O_221,N_14823,N_14775);
xnor UO_222 (O_222,N_14884,N_14896);
or UO_223 (O_223,N_14935,N_14927);
or UO_224 (O_224,N_14856,N_14968);
and UO_225 (O_225,N_14786,N_14968);
and UO_226 (O_226,N_14794,N_14862);
or UO_227 (O_227,N_14841,N_14849);
nand UO_228 (O_228,N_14795,N_14794);
nand UO_229 (O_229,N_14930,N_14974);
nand UO_230 (O_230,N_14938,N_14845);
nor UO_231 (O_231,N_14845,N_14785);
or UO_232 (O_232,N_14827,N_14958);
or UO_233 (O_233,N_14983,N_14835);
nor UO_234 (O_234,N_14782,N_14965);
nand UO_235 (O_235,N_14755,N_14793);
nor UO_236 (O_236,N_14898,N_14875);
nor UO_237 (O_237,N_14874,N_14758);
nor UO_238 (O_238,N_14920,N_14805);
and UO_239 (O_239,N_14928,N_14833);
nor UO_240 (O_240,N_14754,N_14759);
nor UO_241 (O_241,N_14781,N_14772);
nand UO_242 (O_242,N_14989,N_14947);
and UO_243 (O_243,N_14805,N_14844);
and UO_244 (O_244,N_14941,N_14924);
and UO_245 (O_245,N_14777,N_14940);
xnor UO_246 (O_246,N_14758,N_14865);
nand UO_247 (O_247,N_14763,N_14929);
nand UO_248 (O_248,N_14803,N_14955);
nand UO_249 (O_249,N_14798,N_14979);
nor UO_250 (O_250,N_14904,N_14839);
nand UO_251 (O_251,N_14911,N_14927);
nor UO_252 (O_252,N_14879,N_14896);
xnor UO_253 (O_253,N_14820,N_14801);
nand UO_254 (O_254,N_14777,N_14952);
nor UO_255 (O_255,N_14835,N_14902);
and UO_256 (O_256,N_14807,N_14797);
nand UO_257 (O_257,N_14839,N_14750);
or UO_258 (O_258,N_14841,N_14827);
xnor UO_259 (O_259,N_14841,N_14886);
or UO_260 (O_260,N_14864,N_14944);
nor UO_261 (O_261,N_14946,N_14837);
nor UO_262 (O_262,N_14770,N_14761);
nor UO_263 (O_263,N_14874,N_14909);
nand UO_264 (O_264,N_14863,N_14934);
and UO_265 (O_265,N_14976,N_14820);
nor UO_266 (O_266,N_14870,N_14965);
nand UO_267 (O_267,N_14982,N_14842);
xnor UO_268 (O_268,N_14790,N_14750);
or UO_269 (O_269,N_14831,N_14845);
xor UO_270 (O_270,N_14886,N_14982);
or UO_271 (O_271,N_14842,N_14859);
nand UO_272 (O_272,N_14886,N_14971);
and UO_273 (O_273,N_14828,N_14993);
nor UO_274 (O_274,N_14845,N_14951);
or UO_275 (O_275,N_14969,N_14836);
and UO_276 (O_276,N_14985,N_14894);
xor UO_277 (O_277,N_14957,N_14801);
and UO_278 (O_278,N_14958,N_14857);
nand UO_279 (O_279,N_14911,N_14785);
nand UO_280 (O_280,N_14856,N_14876);
xnor UO_281 (O_281,N_14863,N_14842);
nand UO_282 (O_282,N_14956,N_14878);
and UO_283 (O_283,N_14760,N_14895);
or UO_284 (O_284,N_14949,N_14765);
or UO_285 (O_285,N_14951,N_14883);
and UO_286 (O_286,N_14837,N_14825);
nor UO_287 (O_287,N_14762,N_14772);
nor UO_288 (O_288,N_14915,N_14879);
xor UO_289 (O_289,N_14961,N_14852);
nand UO_290 (O_290,N_14769,N_14898);
nor UO_291 (O_291,N_14809,N_14845);
or UO_292 (O_292,N_14935,N_14765);
or UO_293 (O_293,N_14945,N_14800);
nand UO_294 (O_294,N_14800,N_14950);
nor UO_295 (O_295,N_14750,N_14906);
and UO_296 (O_296,N_14759,N_14770);
nand UO_297 (O_297,N_14923,N_14889);
or UO_298 (O_298,N_14784,N_14768);
or UO_299 (O_299,N_14930,N_14954);
nor UO_300 (O_300,N_14894,N_14807);
or UO_301 (O_301,N_14936,N_14933);
xnor UO_302 (O_302,N_14937,N_14892);
and UO_303 (O_303,N_14762,N_14939);
or UO_304 (O_304,N_14949,N_14943);
nor UO_305 (O_305,N_14830,N_14802);
nor UO_306 (O_306,N_14919,N_14940);
nor UO_307 (O_307,N_14926,N_14929);
nand UO_308 (O_308,N_14769,N_14753);
or UO_309 (O_309,N_14997,N_14776);
nand UO_310 (O_310,N_14914,N_14996);
and UO_311 (O_311,N_14796,N_14940);
or UO_312 (O_312,N_14768,N_14984);
or UO_313 (O_313,N_14969,N_14906);
nand UO_314 (O_314,N_14769,N_14999);
or UO_315 (O_315,N_14829,N_14925);
and UO_316 (O_316,N_14972,N_14898);
xnor UO_317 (O_317,N_14991,N_14859);
nor UO_318 (O_318,N_14989,N_14821);
and UO_319 (O_319,N_14817,N_14950);
or UO_320 (O_320,N_14894,N_14820);
or UO_321 (O_321,N_14968,N_14941);
and UO_322 (O_322,N_14801,N_14989);
and UO_323 (O_323,N_14943,N_14955);
nor UO_324 (O_324,N_14825,N_14989);
and UO_325 (O_325,N_14873,N_14867);
and UO_326 (O_326,N_14967,N_14802);
or UO_327 (O_327,N_14994,N_14776);
xor UO_328 (O_328,N_14865,N_14834);
nor UO_329 (O_329,N_14937,N_14905);
nand UO_330 (O_330,N_14855,N_14852);
xnor UO_331 (O_331,N_14812,N_14983);
xnor UO_332 (O_332,N_14981,N_14765);
nand UO_333 (O_333,N_14817,N_14949);
nor UO_334 (O_334,N_14893,N_14980);
or UO_335 (O_335,N_14872,N_14847);
nor UO_336 (O_336,N_14778,N_14822);
xnor UO_337 (O_337,N_14870,N_14881);
nand UO_338 (O_338,N_14916,N_14993);
nand UO_339 (O_339,N_14815,N_14809);
xnor UO_340 (O_340,N_14921,N_14970);
and UO_341 (O_341,N_14882,N_14948);
xnor UO_342 (O_342,N_14954,N_14767);
or UO_343 (O_343,N_14968,N_14949);
nor UO_344 (O_344,N_14850,N_14804);
and UO_345 (O_345,N_14951,N_14914);
or UO_346 (O_346,N_14829,N_14893);
or UO_347 (O_347,N_14807,N_14967);
nor UO_348 (O_348,N_14791,N_14944);
nand UO_349 (O_349,N_14967,N_14987);
nand UO_350 (O_350,N_14771,N_14767);
nor UO_351 (O_351,N_14823,N_14803);
nor UO_352 (O_352,N_14790,N_14803);
nand UO_353 (O_353,N_14800,N_14803);
nor UO_354 (O_354,N_14811,N_14798);
and UO_355 (O_355,N_14797,N_14898);
nor UO_356 (O_356,N_14975,N_14791);
xnor UO_357 (O_357,N_14776,N_14927);
nor UO_358 (O_358,N_14999,N_14906);
nor UO_359 (O_359,N_14784,N_14820);
and UO_360 (O_360,N_14994,N_14752);
and UO_361 (O_361,N_14973,N_14750);
nor UO_362 (O_362,N_14762,N_14765);
nand UO_363 (O_363,N_14859,N_14771);
xnor UO_364 (O_364,N_14902,N_14978);
or UO_365 (O_365,N_14950,N_14896);
xor UO_366 (O_366,N_14862,N_14833);
nor UO_367 (O_367,N_14808,N_14764);
or UO_368 (O_368,N_14877,N_14966);
nor UO_369 (O_369,N_14752,N_14794);
or UO_370 (O_370,N_14768,N_14811);
nor UO_371 (O_371,N_14839,N_14812);
or UO_372 (O_372,N_14966,N_14770);
xor UO_373 (O_373,N_14974,N_14793);
and UO_374 (O_374,N_14887,N_14756);
and UO_375 (O_375,N_14769,N_14940);
xor UO_376 (O_376,N_14962,N_14887);
or UO_377 (O_377,N_14972,N_14976);
and UO_378 (O_378,N_14988,N_14810);
nor UO_379 (O_379,N_14945,N_14955);
nor UO_380 (O_380,N_14905,N_14915);
nand UO_381 (O_381,N_14862,N_14899);
or UO_382 (O_382,N_14843,N_14948);
and UO_383 (O_383,N_14791,N_14794);
nand UO_384 (O_384,N_14918,N_14994);
and UO_385 (O_385,N_14860,N_14879);
nand UO_386 (O_386,N_14755,N_14824);
or UO_387 (O_387,N_14969,N_14962);
or UO_388 (O_388,N_14877,N_14835);
xnor UO_389 (O_389,N_14868,N_14943);
nand UO_390 (O_390,N_14867,N_14844);
or UO_391 (O_391,N_14827,N_14782);
nand UO_392 (O_392,N_14978,N_14933);
and UO_393 (O_393,N_14970,N_14915);
and UO_394 (O_394,N_14937,N_14959);
or UO_395 (O_395,N_14821,N_14920);
nor UO_396 (O_396,N_14933,N_14832);
or UO_397 (O_397,N_14845,N_14776);
and UO_398 (O_398,N_14775,N_14769);
nand UO_399 (O_399,N_14857,N_14880);
nor UO_400 (O_400,N_14888,N_14763);
nor UO_401 (O_401,N_14987,N_14997);
nor UO_402 (O_402,N_14878,N_14847);
nand UO_403 (O_403,N_14949,N_14932);
or UO_404 (O_404,N_14931,N_14873);
nor UO_405 (O_405,N_14822,N_14784);
xor UO_406 (O_406,N_14913,N_14980);
nand UO_407 (O_407,N_14994,N_14824);
or UO_408 (O_408,N_14880,N_14845);
or UO_409 (O_409,N_14859,N_14947);
nor UO_410 (O_410,N_14809,N_14811);
nor UO_411 (O_411,N_14863,N_14884);
or UO_412 (O_412,N_14778,N_14944);
nand UO_413 (O_413,N_14834,N_14812);
nand UO_414 (O_414,N_14980,N_14972);
nand UO_415 (O_415,N_14863,N_14799);
xor UO_416 (O_416,N_14763,N_14802);
nor UO_417 (O_417,N_14770,N_14888);
and UO_418 (O_418,N_14981,N_14845);
nor UO_419 (O_419,N_14836,N_14963);
nand UO_420 (O_420,N_14780,N_14891);
nand UO_421 (O_421,N_14762,N_14950);
and UO_422 (O_422,N_14980,N_14792);
xor UO_423 (O_423,N_14939,N_14840);
nor UO_424 (O_424,N_14976,N_14992);
and UO_425 (O_425,N_14860,N_14885);
nor UO_426 (O_426,N_14876,N_14992);
nand UO_427 (O_427,N_14791,N_14788);
nor UO_428 (O_428,N_14826,N_14841);
or UO_429 (O_429,N_14983,N_14984);
nand UO_430 (O_430,N_14819,N_14987);
nor UO_431 (O_431,N_14946,N_14857);
and UO_432 (O_432,N_14871,N_14786);
and UO_433 (O_433,N_14824,N_14881);
and UO_434 (O_434,N_14754,N_14841);
nor UO_435 (O_435,N_14962,N_14806);
or UO_436 (O_436,N_14908,N_14854);
nor UO_437 (O_437,N_14849,N_14811);
and UO_438 (O_438,N_14925,N_14947);
nor UO_439 (O_439,N_14984,N_14832);
or UO_440 (O_440,N_14961,N_14860);
and UO_441 (O_441,N_14991,N_14823);
or UO_442 (O_442,N_14823,N_14948);
xor UO_443 (O_443,N_14851,N_14840);
or UO_444 (O_444,N_14975,N_14954);
nand UO_445 (O_445,N_14843,N_14975);
and UO_446 (O_446,N_14772,N_14790);
or UO_447 (O_447,N_14990,N_14750);
or UO_448 (O_448,N_14776,N_14774);
xor UO_449 (O_449,N_14762,N_14958);
or UO_450 (O_450,N_14824,N_14889);
nor UO_451 (O_451,N_14908,N_14977);
and UO_452 (O_452,N_14802,N_14950);
and UO_453 (O_453,N_14834,N_14851);
nor UO_454 (O_454,N_14786,N_14971);
nor UO_455 (O_455,N_14987,N_14830);
or UO_456 (O_456,N_14824,N_14962);
nand UO_457 (O_457,N_14898,N_14958);
nand UO_458 (O_458,N_14816,N_14807);
nor UO_459 (O_459,N_14814,N_14765);
nand UO_460 (O_460,N_14920,N_14847);
xor UO_461 (O_461,N_14851,N_14966);
and UO_462 (O_462,N_14962,N_14997);
nor UO_463 (O_463,N_14925,N_14820);
nand UO_464 (O_464,N_14876,N_14810);
nor UO_465 (O_465,N_14899,N_14844);
nand UO_466 (O_466,N_14912,N_14843);
nor UO_467 (O_467,N_14867,N_14843);
nand UO_468 (O_468,N_14971,N_14980);
nand UO_469 (O_469,N_14794,N_14801);
or UO_470 (O_470,N_14946,N_14976);
nand UO_471 (O_471,N_14762,N_14971);
or UO_472 (O_472,N_14850,N_14938);
xnor UO_473 (O_473,N_14908,N_14846);
nand UO_474 (O_474,N_14847,N_14796);
or UO_475 (O_475,N_14795,N_14792);
and UO_476 (O_476,N_14753,N_14756);
nand UO_477 (O_477,N_14971,N_14846);
nor UO_478 (O_478,N_14989,N_14986);
nor UO_479 (O_479,N_14765,N_14983);
nor UO_480 (O_480,N_14851,N_14968);
nand UO_481 (O_481,N_14943,N_14898);
or UO_482 (O_482,N_14935,N_14891);
nor UO_483 (O_483,N_14896,N_14989);
and UO_484 (O_484,N_14869,N_14862);
or UO_485 (O_485,N_14812,N_14777);
xnor UO_486 (O_486,N_14952,N_14923);
nand UO_487 (O_487,N_14794,N_14872);
or UO_488 (O_488,N_14938,N_14901);
xnor UO_489 (O_489,N_14751,N_14895);
nand UO_490 (O_490,N_14864,N_14941);
or UO_491 (O_491,N_14917,N_14808);
or UO_492 (O_492,N_14751,N_14940);
nor UO_493 (O_493,N_14931,N_14955);
and UO_494 (O_494,N_14782,N_14875);
nand UO_495 (O_495,N_14927,N_14796);
xnor UO_496 (O_496,N_14936,N_14859);
nand UO_497 (O_497,N_14884,N_14921);
nor UO_498 (O_498,N_14895,N_14929);
nor UO_499 (O_499,N_14981,N_14942);
or UO_500 (O_500,N_14941,N_14787);
xnor UO_501 (O_501,N_14994,N_14961);
nand UO_502 (O_502,N_14770,N_14858);
nor UO_503 (O_503,N_14942,N_14870);
xor UO_504 (O_504,N_14775,N_14850);
nor UO_505 (O_505,N_14788,N_14796);
xnor UO_506 (O_506,N_14751,N_14947);
or UO_507 (O_507,N_14931,N_14792);
and UO_508 (O_508,N_14838,N_14835);
and UO_509 (O_509,N_14919,N_14996);
nor UO_510 (O_510,N_14983,N_14787);
nor UO_511 (O_511,N_14936,N_14864);
nor UO_512 (O_512,N_14806,N_14902);
nand UO_513 (O_513,N_14972,N_14792);
and UO_514 (O_514,N_14916,N_14977);
or UO_515 (O_515,N_14927,N_14973);
and UO_516 (O_516,N_14825,N_14912);
and UO_517 (O_517,N_14846,N_14775);
or UO_518 (O_518,N_14824,N_14848);
xnor UO_519 (O_519,N_14840,N_14896);
and UO_520 (O_520,N_14761,N_14763);
or UO_521 (O_521,N_14984,N_14989);
or UO_522 (O_522,N_14823,N_14947);
nand UO_523 (O_523,N_14867,N_14798);
xor UO_524 (O_524,N_14791,N_14776);
or UO_525 (O_525,N_14802,N_14823);
nand UO_526 (O_526,N_14939,N_14951);
nand UO_527 (O_527,N_14830,N_14869);
and UO_528 (O_528,N_14919,N_14973);
and UO_529 (O_529,N_14814,N_14859);
and UO_530 (O_530,N_14879,N_14765);
and UO_531 (O_531,N_14776,N_14807);
nor UO_532 (O_532,N_14880,N_14912);
and UO_533 (O_533,N_14946,N_14778);
xnor UO_534 (O_534,N_14957,N_14973);
nand UO_535 (O_535,N_14854,N_14755);
or UO_536 (O_536,N_14838,N_14817);
and UO_537 (O_537,N_14950,N_14884);
nand UO_538 (O_538,N_14930,N_14976);
and UO_539 (O_539,N_14987,N_14806);
xor UO_540 (O_540,N_14876,N_14978);
nand UO_541 (O_541,N_14967,N_14908);
nand UO_542 (O_542,N_14851,N_14804);
xor UO_543 (O_543,N_14750,N_14856);
or UO_544 (O_544,N_14907,N_14943);
xnor UO_545 (O_545,N_14972,N_14979);
nor UO_546 (O_546,N_14762,N_14871);
xnor UO_547 (O_547,N_14930,N_14871);
nor UO_548 (O_548,N_14979,N_14793);
nand UO_549 (O_549,N_14804,N_14815);
and UO_550 (O_550,N_14859,N_14928);
and UO_551 (O_551,N_14868,N_14952);
nor UO_552 (O_552,N_14899,N_14906);
nor UO_553 (O_553,N_14880,N_14841);
and UO_554 (O_554,N_14908,N_14890);
or UO_555 (O_555,N_14773,N_14949);
nand UO_556 (O_556,N_14967,N_14783);
nand UO_557 (O_557,N_14809,N_14972);
and UO_558 (O_558,N_14917,N_14958);
nor UO_559 (O_559,N_14759,N_14855);
or UO_560 (O_560,N_14773,N_14972);
or UO_561 (O_561,N_14914,N_14829);
nand UO_562 (O_562,N_14963,N_14951);
nor UO_563 (O_563,N_14824,N_14871);
or UO_564 (O_564,N_14980,N_14955);
and UO_565 (O_565,N_14851,N_14867);
nor UO_566 (O_566,N_14827,N_14937);
or UO_567 (O_567,N_14931,N_14965);
and UO_568 (O_568,N_14760,N_14803);
xnor UO_569 (O_569,N_14798,N_14960);
nor UO_570 (O_570,N_14790,N_14770);
and UO_571 (O_571,N_14833,N_14962);
nand UO_572 (O_572,N_14767,N_14833);
nand UO_573 (O_573,N_14871,N_14833);
xor UO_574 (O_574,N_14933,N_14836);
nand UO_575 (O_575,N_14916,N_14762);
xor UO_576 (O_576,N_14875,N_14813);
or UO_577 (O_577,N_14783,N_14970);
and UO_578 (O_578,N_14859,N_14871);
xor UO_579 (O_579,N_14873,N_14856);
nor UO_580 (O_580,N_14905,N_14849);
xor UO_581 (O_581,N_14785,N_14999);
or UO_582 (O_582,N_14973,N_14917);
and UO_583 (O_583,N_14940,N_14971);
nand UO_584 (O_584,N_14859,N_14789);
nand UO_585 (O_585,N_14875,N_14858);
nand UO_586 (O_586,N_14982,N_14857);
nor UO_587 (O_587,N_14989,N_14822);
and UO_588 (O_588,N_14834,N_14898);
or UO_589 (O_589,N_14846,N_14809);
and UO_590 (O_590,N_14814,N_14978);
and UO_591 (O_591,N_14922,N_14985);
nor UO_592 (O_592,N_14771,N_14934);
xnor UO_593 (O_593,N_14995,N_14891);
or UO_594 (O_594,N_14976,N_14784);
nor UO_595 (O_595,N_14759,N_14786);
xnor UO_596 (O_596,N_14955,N_14923);
or UO_597 (O_597,N_14923,N_14972);
nor UO_598 (O_598,N_14989,N_14948);
or UO_599 (O_599,N_14866,N_14892);
nor UO_600 (O_600,N_14994,N_14879);
nand UO_601 (O_601,N_14775,N_14880);
nand UO_602 (O_602,N_14877,N_14882);
or UO_603 (O_603,N_14871,N_14909);
or UO_604 (O_604,N_14825,N_14964);
nor UO_605 (O_605,N_14920,N_14845);
nor UO_606 (O_606,N_14787,N_14956);
and UO_607 (O_607,N_14796,N_14930);
nor UO_608 (O_608,N_14822,N_14756);
or UO_609 (O_609,N_14756,N_14910);
nand UO_610 (O_610,N_14849,N_14827);
and UO_611 (O_611,N_14884,N_14932);
or UO_612 (O_612,N_14830,N_14954);
or UO_613 (O_613,N_14873,N_14987);
nor UO_614 (O_614,N_14966,N_14971);
xnor UO_615 (O_615,N_14960,N_14946);
nand UO_616 (O_616,N_14929,N_14791);
and UO_617 (O_617,N_14846,N_14759);
or UO_618 (O_618,N_14873,N_14764);
nor UO_619 (O_619,N_14784,N_14921);
nor UO_620 (O_620,N_14862,N_14847);
or UO_621 (O_621,N_14886,N_14957);
xnor UO_622 (O_622,N_14828,N_14880);
nor UO_623 (O_623,N_14878,N_14767);
xor UO_624 (O_624,N_14960,N_14837);
xnor UO_625 (O_625,N_14939,N_14959);
and UO_626 (O_626,N_14907,N_14819);
nor UO_627 (O_627,N_14787,N_14871);
and UO_628 (O_628,N_14757,N_14917);
nor UO_629 (O_629,N_14757,N_14812);
nand UO_630 (O_630,N_14872,N_14934);
nand UO_631 (O_631,N_14958,N_14990);
or UO_632 (O_632,N_14751,N_14848);
or UO_633 (O_633,N_14829,N_14917);
nand UO_634 (O_634,N_14884,N_14930);
nand UO_635 (O_635,N_14862,N_14907);
and UO_636 (O_636,N_14955,N_14780);
nand UO_637 (O_637,N_14980,N_14833);
nor UO_638 (O_638,N_14960,N_14809);
nand UO_639 (O_639,N_14990,N_14762);
or UO_640 (O_640,N_14897,N_14791);
xor UO_641 (O_641,N_14930,N_14846);
nor UO_642 (O_642,N_14782,N_14800);
or UO_643 (O_643,N_14853,N_14987);
nand UO_644 (O_644,N_14953,N_14806);
nand UO_645 (O_645,N_14989,N_14933);
nor UO_646 (O_646,N_14996,N_14950);
nor UO_647 (O_647,N_14828,N_14797);
nor UO_648 (O_648,N_14834,N_14892);
and UO_649 (O_649,N_14873,N_14816);
nor UO_650 (O_650,N_14898,N_14966);
or UO_651 (O_651,N_14893,N_14818);
nand UO_652 (O_652,N_14877,N_14823);
or UO_653 (O_653,N_14851,N_14841);
or UO_654 (O_654,N_14972,N_14832);
and UO_655 (O_655,N_14810,N_14822);
or UO_656 (O_656,N_14983,N_14951);
and UO_657 (O_657,N_14834,N_14781);
nor UO_658 (O_658,N_14891,N_14924);
nand UO_659 (O_659,N_14958,N_14918);
nor UO_660 (O_660,N_14888,N_14944);
and UO_661 (O_661,N_14863,N_14859);
nand UO_662 (O_662,N_14870,N_14974);
nor UO_663 (O_663,N_14936,N_14788);
and UO_664 (O_664,N_14865,N_14965);
nand UO_665 (O_665,N_14790,N_14884);
nand UO_666 (O_666,N_14810,N_14973);
or UO_667 (O_667,N_14820,N_14753);
nand UO_668 (O_668,N_14755,N_14805);
nor UO_669 (O_669,N_14760,N_14865);
or UO_670 (O_670,N_14897,N_14909);
or UO_671 (O_671,N_14840,N_14856);
nor UO_672 (O_672,N_14918,N_14860);
and UO_673 (O_673,N_14820,N_14836);
or UO_674 (O_674,N_14837,N_14900);
xnor UO_675 (O_675,N_14768,N_14947);
and UO_676 (O_676,N_14925,N_14851);
and UO_677 (O_677,N_14978,N_14851);
and UO_678 (O_678,N_14884,N_14821);
or UO_679 (O_679,N_14764,N_14834);
or UO_680 (O_680,N_14952,N_14750);
nand UO_681 (O_681,N_14938,N_14903);
and UO_682 (O_682,N_14872,N_14806);
and UO_683 (O_683,N_14875,N_14930);
and UO_684 (O_684,N_14859,N_14852);
nor UO_685 (O_685,N_14822,N_14982);
nand UO_686 (O_686,N_14757,N_14916);
xor UO_687 (O_687,N_14890,N_14786);
or UO_688 (O_688,N_14792,N_14805);
nor UO_689 (O_689,N_14841,N_14955);
nand UO_690 (O_690,N_14769,N_14811);
or UO_691 (O_691,N_14989,N_14960);
nor UO_692 (O_692,N_14895,N_14863);
or UO_693 (O_693,N_14998,N_14988);
or UO_694 (O_694,N_14904,N_14796);
nor UO_695 (O_695,N_14809,N_14820);
nand UO_696 (O_696,N_14982,N_14758);
and UO_697 (O_697,N_14876,N_14764);
or UO_698 (O_698,N_14909,N_14955);
nand UO_699 (O_699,N_14856,N_14969);
nand UO_700 (O_700,N_14753,N_14975);
or UO_701 (O_701,N_14952,N_14830);
and UO_702 (O_702,N_14905,N_14993);
nor UO_703 (O_703,N_14819,N_14886);
nand UO_704 (O_704,N_14804,N_14874);
xnor UO_705 (O_705,N_14940,N_14909);
nand UO_706 (O_706,N_14932,N_14885);
nand UO_707 (O_707,N_14826,N_14787);
and UO_708 (O_708,N_14909,N_14959);
nor UO_709 (O_709,N_14973,N_14886);
nor UO_710 (O_710,N_14819,N_14925);
nor UO_711 (O_711,N_14912,N_14934);
and UO_712 (O_712,N_14977,N_14871);
nand UO_713 (O_713,N_14770,N_14791);
or UO_714 (O_714,N_14783,N_14852);
and UO_715 (O_715,N_14990,N_14821);
xnor UO_716 (O_716,N_14804,N_14757);
xnor UO_717 (O_717,N_14822,N_14915);
and UO_718 (O_718,N_14759,N_14765);
nor UO_719 (O_719,N_14894,N_14868);
nand UO_720 (O_720,N_14953,N_14856);
or UO_721 (O_721,N_14992,N_14884);
and UO_722 (O_722,N_14901,N_14944);
and UO_723 (O_723,N_14963,N_14879);
nand UO_724 (O_724,N_14762,N_14825);
and UO_725 (O_725,N_14999,N_14819);
nand UO_726 (O_726,N_14863,N_14844);
nor UO_727 (O_727,N_14791,N_14947);
nand UO_728 (O_728,N_14771,N_14807);
and UO_729 (O_729,N_14979,N_14942);
nor UO_730 (O_730,N_14969,N_14866);
and UO_731 (O_731,N_14876,N_14964);
xnor UO_732 (O_732,N_14858,N_14781);
or UO_733 (O_733,N_14843,N_14825);
nand UO_734 (O_734,N_14762,N_14902);
xor UO_735 (O_735,N_14917,N_14947);
xor UO_736 (O_736,N_14761,N_14756);
or UO_737 (O_737,N_14822,N_14772);
nor UO_738 (O_738,N_14934,N_14853);
or UO_739 (O_739,N_14965,N_14904);
and UO_740 (O_740,N_14931,N_14845);
xor UO_741 (O_741,N_14966,N_14862);
and UO_742 (O_742,N_14786,N_14910);
nor UO_743 (O_743,N_14971,N_14866);
or UO_744 (O_744,N_14786,N_14873);
xnor UO_745 (O_745,N_14943,N_14832);
xnor UO_746 (O_746,N_14767,N_14984);
or UO_747 (O_747,N_14952,N_14793);
nor UO_748 (O_748,N_14841,N_14937);
xor UO_749 (O_749,N_14994,N_14822);
and UO_750 (O_750,N_14994,N_14957);
nor UO_751 (O_751,N_14910,N_14859);
and UO_752 (O_752,N_14878,N_14977);
nor UO_753 (O_753,N_14871,N_14919);
nand UO_754 (O_754,N_14891,N_14827);
nand UO_755 (O_755,N_14775,N_14856);
or UO_756 (O_756,N_14921,N_14764);
or UO_757 (O_757,N_14855,N_14796);
nor UO_758 (O_758,N_14920,N_14977);
nor UO_759 (O_759,N_14922,N_14912);
and UO_760 (O_760,N_14971,N_14970);
xor UO_761 (O_761,N_14997,N_14843);
nand UO_762 (O_762,N_14778,N_14932);
nand UO_763 (O_763,N_14816,N_14910);
nand UO_764 (O_764,N_14882,N_14785);
nor UO_765 (O_765,N_14960,N_14912);
or UO_766 (O_766,N_14928,N_14756);
or UO_767 (O_767,N_14820,N_14777);
or UO_768 (O_768,N_14834,N_14925);
nand UO_769 (O_769,N_14826,N_14795);
xor UO_770 (O_770,N_14753,N_14845);
and UO_771 (O_771,N_14917,N_14932);
nand UO_772 (O_772,N_14953,N_14996);
xnor UO_773 (O_773,N_14964,N_14834);
nor UO_774 (O_774,N_14755,N_14946);
xnor UO_775 (O_775,N_14835,N_14904);
xor UO_776 (O_776,N_14773,N_14894);
nor UO_777 (O_777,N_14887,N_14847);
and UO_778 (O_778,N_14756,N_14971);
nand UO_779 (O_779,N_14983,N_14861);
nand UO_780 (O_780,N_14960,N_14984);
or UO_781 (O_781,N_14975,N_14912);
and UO_782 (O_782,N_14958,N_14874);
nor UO_783 (O_783,N_14784,N_14833);
and UO_784 (O_784,N_14870,N_14849);
nor UO_785 (O_785,N_14798,N_14807);
nor UO_786 (O_786,N_14813,N_14907);
nand UO_787 (O_787,N_14897,N_14888);
nor UO_788 (O_788,N_14895,N_14918);
nand UO_789 (O_789,N_14773,N_14833);
nor UO_790 (O_790,N_14763,N_14801);
and UO_791 (O_791,N_14803,N_14971);
nor UO_792 (O_792,N_14836,N_14814);
nor UO_793 (O_793,N_14829,N_14913);
and UO_794 (O_794,N_14822,N_14932);
nand UO_795 (O_795,N_14944,N_14896);
xnor UO_796 (O_796,N_14817,N_14881);
and UO_797 (O_797,N_14848,N_14883);
nand UO_798 (O_798,N_14964,N_14773);
or UO_799 (O_799,N_14978,N_14808);
nor UO_800 (O_800,N_14818,N_14763);
and UO_801 (O_801,N_14840,N_14931);
xnor UO_802 (O_802,N_14756,N_14821);
nor UO_803 (O_803,N_14836,N_14791);
nor UO_804 (O_804,N_14945,N_14846);
xor UO_805 (O_805,N_14913,N_14853);
nand UO_806 (O_806,N_14770,N_14835);
nand UO_807 (O_807,N_14765,N_14985);
or UO_808 (O_808,N_14782,N_14810);
and UO_809 (O_809,N_14773,N_14914);
xnor UO_810 (O_810,N_14909,N_14850);
nor UO_811 (O_811,N_14988,N_14982);
or UO_812 (O_812,N_14918,N_14967);
nor UO_813 (O_813,N_14949,N_14785);
nand UO_814 (O_814,N_14916,N_14836);
nand UO_815 (O_815,N_14993,N_14853);
and UO_816 (O_816,N_14913,N_14862);
nor UO_817 (O_817,N_14913,N_14970);
nor UO_818 (O_818,N_14877,N_14967);
or UO_819 (O_819,N_14891,N_14945);
and UO_820 (O_820,N_14879,N_14956);
or UO_821 (O_821,N_14769,N_14982);
nand UO_822 (O_822,N_14968,N_14761);
or UO_823 (O_823,N_14832,N_14885);
nor UO_824 (O_824,N_14940,N_14868);
nor UO_825 (O_825,N_14865,N_14943);
or UO_826 (O_826,N_14761,N_14927);
or UO_827 (O_827,N_14946,N_14886);
and UO_828 (O_828,N_14830,N_14951);
xor UO_829 (O_829,N_14932,N_14848);
and UO_830 (O_830,N_14845,N_14997);
nor UO_831 (O_831,N_14901,N_14813);
or UO_832 (O_832,N_14838,N_14815);
or UO_833 (O_833,N_14826,N_14780);
or UO_834 (O_834,N_14876,N_14809);
or UO_835 (O_835,N_14945,N_14943);
nor UO_836 (O_836,N_14866,N_14948);
or UO_837 (O_837,N_14920,N_14951);
and UO_838 (O_838,N_14755,N_14762);
nand UO_839 (O_839,N_14877,N_14869);
nand UO_840 (O_840,N_14813,N_14996);
or UO_841 (O_841,N_14859,N_14993);
and UO_842 (O_842,N_14984,N_14986);
xor UO_843 (O_843,N_14996,N_14981);
or UO_844 (O_844,N_14756,N_14838);
nand UO_845 (O_845,N_14922,N_14862);
xor UO_846 (O_846,N_14814,N_14841);
nor UO_847 (O_847,N_14984,N_14955);
or UO_848 (O_848,N_14797,N_14993);
xnor UO_849 (O_849,N_14868,N_14850);
nand UO_850 (O_850,N_14806,N_14765);
nor UO_851 (O_851,N_14977,N_14870);
nand UO_852 (O_852,N_14999,N_14965);
nor UO_853 (O_853,N_14956,N_14819);
nand UO_854 (O_854,N_14805,N_14993);
nand UO_855 (O_855,N_14990,N_14755);
nor UO_856 (O_856,N_14977,N_14959);
or UO_857 (O_857,N_14856,N_14779);
or UO_858 (O_858,N_14933,N_14881);
xnor UO_859 (O_859,N_14836,N_14950);
nor UO_860 (O_860,N_14764,N_14903);
or UO_861 (O_861,N_14921,N_14891);
xor UO_862 (O_862,N_14912,N_14931);
or UO_863 (O_863,N_14889,N_14911);
nand UO_864 (O_864,N_14774,N_14855);
nand UO_865 (O_865,N_14883,N_14953);
and UO_866 (O_866,N_14930,N_14928);
or UO_867 (O_867,N_14822,N_14842);
xor UO_868 (O_868,N_14843,N_14827);
or UO_869 (O_869,N_14898,N_14914);
or UO_870 (O_870,N_14795,N_14986);
and UO_871 (O_871,N_14832,N_14924);
or UO_872 (O_872,N_14942,N_14802);
nor UO_873 (O_873,N_14863,N_14890);
nand UO_874 (O_874,N_14992,N_14790);
and UO_875 (O_875,N_14934,N_14882);
xnor UO_876 (O_876,N_14880,N_14852);
and UO_877 (O_877,N_14778,N_14781);
nand UO_878 (O_878,N_14863,N_14885);
nand UO_879 (O_879,N_14962,N_14770);
nand UO_880 (O_880,N_14757,N_14864);
and UO_881 (O_881,N_14988,N_14909);
nor UO_882 (O_882,N_14814,N_14944);
nor UO_883 (O_883,N_14857,N_14889);
or UO_884 (O_884,N_14867,N_14847);
nor UO_885 (O_885,N_14840,N_14940);
nand UO_886 (O_886,N_14855,N_14915);
xor UO_887 (O_887,N_14970,N_14786);
or UO_888 (O_888,N_14934,N_14979);
and UO_889 (O_889,N_14928,N_14958);
nand UO_890 (O_890,N_14997,N_14760);
nor UO_891 (O_891,N_14904,N_14901);
nor UO_892 (O_892,N_14930,N_14848);
and UO_893 (O_893,N_14962,N_14951);
and UO_894 (O_894,N_14964,N_14973);
and UO_895 (O_895,N_14843,N_14909);
nor UO_896 (O_896,N_14879,N_14977);
nand UO_897 (O_897,N_14955,N_14892);
nor UO_898 (O_898,N_14891,N_14766);
or UO_899 (O_899,N_14804,N_14845);
or UO_900 (O_900,N_14838,N_14825);
nand UO_901 (O_901,N_14973,N_14785);
nand UO_902 (O_902,N_14804,N_14940);
or UO_903 (O_903,N_14759,N_14768);
and UO_904 (O_904,N_14992,N_14815);
and UO_905 (O_905,N_14792,N_14919);
or UO_906 (O_906,N_14969,N_14883);
and UO_907 (O_907,N_14839,N_14803);
nor UO_908 (O_908,N_14874,N_14823);
and UO_909 (O_909,N_14755,N_14985);
nor UO_910 (O_910,N_14779,N_14783);
nor UO_911 (O_911,N_14818,N_14946);
nor UO_912 (O_912,N_14968,N_14794);
nand UO_913 (O_913,N_14884,N_14853);
xnor UO_914 (O_914,N_14921,N_14986);
or UO_915 (O_915,N_14855,N_14974);
nor UO_916 (O_916,N_14941,N_14763);
or UO_917 (O_917,N_14798,N_14976);
and UO_918 (O_918,N_14763,N_14760);
xnor UO_919 (O_919,N_14815,N_14970);
xor UO_920 (O_920,N_14891,N_14789);
or UO_921 (O_921,N_14959,N_14762);
nor UO_922 (O_922,N_14791,N_14904);
nor UO_923 (O_923,N_14911,N_14914);
nor UO_924 (O_924,N_14921,N_14852);
nor UO_925 (O_925,N_14908,N_14934);
nor UO_926 (O_926,N_14757,N_14914);
and UO_927 (O_927,N_14910,N_14759);
nand UO_928 (O_928,N_14791,N_14916);
or UO_929 (O_929,N_14772,N_14898);
and UO_930 (O_930,N_14921,N_14786);
and UO_931 (O_931,N_14810,N_14792);
nor UO_932 (O_932,N_14827,N_14905);
nor UO_933 (O_933,N_14868,N_14802);
and UO_934 (O_934,N_14857,N_14788);
xnor UO_935 (O_935,N_14821,N_14836);
nor UO_936 (O_936,N_14912,N_14777);
and UO_937 (O_937,N_14958,N_14826);
nand UO_938 (O_938,N_14973,N_14968);
and UO_939 (O_939,N_14949,N_14988);
or UO_940 (O_940,N_14932,N_14899);
or UO_941 (O_941,N_14910,N_14798);
or UO_942 (O_942,N_14827,N_14864);
xor UO_943 (O_943,N_14944,N_14980);
and UO_944 (O_944,N_14966,N_14980);
or UO_945 (O_945,N_14896,N_14802);
and UO_946 (O_946,N_14814,N_14995);
and UO_947 (O_947,N_14893,N_14863);
and UO_948 (O_948,N_14946,N_14972);
nor UO_949 (O_949,N_14787,N_14766);
or UO_950 (O_950,N_14914,N_14967);
nand UO_951 (O_951,N_14759,N_14750);
nand UO_952 (O_952,N_14862,N_14952);
nand UO_953 (O_953,N_14895,N_14900);
and UO_954 (O_954,N_14932,N_14986);
nand UO_955 (O_955,N_14942,N_14917);
nand UO_956 (O_956,N_14979,N_14980);
and UO_957 (O_957,N_14821,N_14933);
nor UO_958 (O_958,N_14955,N_14800);
or UO_959 (O_959,N_14959,N_14972);
nor UO_960 (O_960,N_14830,N_14806);
and UO_961 (O_961,N_14768,N_14891);
or UO_962 (O_962,N_14877,N_14993);
or UO_963 (O_963,N_14989,N_14950);
or UO_964 (O_964,N_14760,N_14767);
nand UO_965 (O_965,N_14999,N_14982);
nor UO_966 (O_966,N_14850,N_14998);
nor UO_967 (O_967,N_14983,N_14981);
nor UO_968 (O_968,N_14890,N_14891);
nor UO_969 (O_969,N_14883,N_14784);
nand UO_970 (O_970,N_14867,N_14801);
nand UO_971 (O_971,N_14973,N_14903);
nor UO_972 (O_972,N_14890,N_14793);
xor UO_973 (O_973,N_14994,N_14804);
nor UO_974 (O_974,N_14832,N_14813);
or UO_975 (O_975,N_14956,N_14916);
or UO_976 (O_976,N_14753,N_14787);
and UO_977 (O_977,N_14993,N_14808);
or UO_978 (O_978,N_14960,N_14895);
and UO_979 (O_979,N_14971,N_14900);
or UO_980 (O_980,N_14783,N_14793);
nand UO_981 (O_981,N_14851,N_14833);
nand UO_982 (O_982,N_14831,N_14777);
and UO_983 (O_983,N_14878,N_14832);
or UO_984 (O_984,N_14854,N_14853);
nand UO_985 (O_985,N_14962,N_14836);
or UO_986 (O_986,N_14898,N_14820);
xnor UO_987 (O_987,N_14941,N_14891);
and UO_988 (O_988,N_14759,N_14826);
nor UO_989 (O_989,N_14822,N_14773);
or UO_990 (O_990,N_14980,N_14860);
and UO_991 (O_991,N_14963,N_14899);
and UO_992 (O_992,N_14777,N_14769);
nor UO_993 (O_993,N_14761,N_14905);
nand UO_994 (O_994,N_14940,N_14878);
nor UO_995 (O_995,N_14860,N_14854);
and UO_996 (O_996,N_14978,N_14982);
nor UO_997 (O_997,N_14985,N_14777);
nand UO_998 (O_998,N_14841,N_14952);
or UO_999 (O_999,N_14782,N_14855);
nor UO_1000 (O_1000,N_14918,N_14889);
and UO_1001 (O_1001,N_14778,N_14973);
or UO_1002 (O_1002,N_14789,N_14925);
nand UO_1003 (O_1003,N_14877,N_14940);
nor UO_1004 (O_1004,N_14823,N_14795);
and UO_1005 (O_1005,N_14809,N_14829);
nor UO_1006 (O_1006,N_14810,N_14956);
or UO_1007 (O_1007,N_14887,N_14853);
nor UO_1008 (O_1008,N_14942,N_14843);
or UO_1009 (O_1009,N_14814,N_14877);
and UO_1010 (O_1010,N_14754,N_14855);
xor UO_1011 (O_1011,N_14801,N_14774);
or UO_1012 (O_1012,N_14948,N_14946);
nor UO_1013 (O_1013,N_14777,N_14896);
or UO_1014 (O_1014,N_14759,N_14971);
or UO_1015 (O_1015,N_14968,N_14819);
nand UO_1016 (O_1016,N_14995,N_14974);
nor UO_1017 (O_1017,N_14755,N_14945);
nand UO_1018 (O_1018,N_14891,N_14973);
or UO_1019 (O_1019,N_14958,N_14764);
nor UO_1020 (O_1020,N_14900,N_14832);
nor UO_1021 (O_1021,N_14877,N_14811);
or UO_1022 (O_1022,N_14897,N_14997);
xor UO_1023 (O_1023,N_14779,N_14756);
nand UO_1024 (O_1024,N_14759,N_14959);
or UO_1025 (O_1025,N_14893,N_14858);
nand UO_1026 (O_1026,N_14885,N_14834);
or UO_1027 (O_1027,N_14986,N_14951);
nor UO_1028 (O_1028,N_14888,N_14761);
or UO_1029 (O_1029,N_14783,N_14752);
or UO_1030 (O_1030,N_14753,N_14863);
or UO_1031 (O_1031,N_14946,N_14907);
nor UO_1032 (O_1032,N_14909,N_14971);
and UO_1033 (O_1033,N_14845,N_14900);
nand UO_1034 (O_1034,N_14883,N_14993);
and UO_1035 (O_1035,N_14815,N_14872);
and UO_1036 (O_1036,N_14994,N_14979);
nand UO_1037 (O_1037,N_14983,N_14923);
or UO_1038 (O_1038,N_14992,N_14832);
or UO_1039 (O_1039,N_14838,N_14871);
and UO_1040 (O_1040,N_14911,N_14945);
or UO_1041 (O_1041,N_14910,N_14844);
or UO_1042 (O_1042,N_14779,N_14880);
nand UO_1043 (O_1043,N_14845,N_14879);
xnor UO_1044 (O_1044,N_14908,N_14978);
nor UO_1045 (O_1045,N_14860,N_14986);
nand UO_1046 (O_1046,N_14847,N_14968);
nor UO_1047 (O_1047,N_14953,N_14767);
nor UO_1048 (O_1048,N_14787,N_14758);
nor UO_1049 (O_1049,N_14795,N_14900);
nand UO_1050 (O_1050,N_14782,N_14915);
or UO_1051 (O_1051,N_14870,N_14888);
xor UO_1052 (O_1052,N_14898,N_14823);
or UO_1053 (O_1053,N_14989,N_14832);
and UO_1054 (O_1054,N_14757,N_14909);
or UO_1055 (O_1055,N_14885,N_14982);
and UO_1056 (O_1056,N_14926,N_14956);
nand UO_1057 (O_1057,N_14928,N_14852);
xnor UO_1058 (O_1058,N_14838,N_14928);
nand UO_1059 (O_1059,N_14871,N_14826);
or UO_1060 (O_1060,N_14885,N_14939);
and UO_1061 (O_1061,N_14947,N_14844);
and UO_1062 (O_1062,N_14901,N_14909);
nor UO_1063 (O_1063,N_14890,N_14932);
nand UO_1064 (O_1064,N_14820,N_14982);
nand UO_1065 (O_1065,N_14870,N_14996);
or UO_1066 (O_1066,N_14932,N_14873);
and UO_1067 (O_1067,N_14824,N_14783);
or UO_1068 (O_1068,N_14795,N_14831);
and UO_1069 (O_1069,N_14845,N_14756);
or UO_1070 (O_1070,N_14974,N_14811);
xnor UO_1071 (O_1071,N_14891,N_14816);
nand UO_1072 (O_1072,N_14933,N_14961);
xnor UO_1073 (O_1073,N_14989,N_14925);
nand UO_1074 (O_1074,N_14801,N_14849);
nor UO_1075 (O_1075,N_14869,N_14832);
or UO_1076 (O_1076,N_14903,N_14925);
or UO_1077 (O_1077,N_14980,N_14905);
or UO_1078 (O_1078,N_14964,N_14928);
xor UO_1079 (O_1079,N_14910,N_14960);
nor UO_1080 (O_1080,N_14930,N_14999);
nand UO_1081 (O_1081,N_14939,N_14932);
or UO_1082 (O_1082,N_14819,N_14761);
and UO_1083 (O_1083,N_14836,N_14939);
or UO_1084 (O_1084,N_14789,N_14824);
nor UO_1085 (O_1085,N_14911,N_14990);
xnor UO_1086 (O_1086,N_14828,N_14757);
nor UO_1087 (O_1087,N_14759,N_14992);
or UO_1088 (O_1088,N_14880,N_14800);
xnor UO_1089 (O_1089,N_14896,N_14922);
nor UO_1090 (O_1090,N_14969,N_14948);
or UO_1091 (O_1091,N_14805,N_14808);
or UO_1092 (O_1092,N_14761,N_14999);
nor UO_1093 (O_1093,N_14981,N_14844);
nand UO_1094 (O_1094,N_14898,N_14762);
xor UO_1095 (O_1095,N_14968,N_14986);
and UO_1096 (O_1096,N_14773,N_14825);
nand UO_1097 (O_1097,N_14752,N_14775);
xor UO_1098 (O_1098,N_14811,N_14851);
or UO_1099 (O_1099,N_14808,N_14905);
nand UO_1100 (O_1100,N_14832,N_14888);
nor UO_1101 (O_1101,N_14884,N_14946);
nor UO_1102 (O_1102,N_14949,N_14844);
nor UO_1103 (O_1103,N_14918,N_14909);
nand UO_1104 (O_1104,N_14801,N_14828);
or UO_1105 (O_1105,N_14809,N_14979);
xor UO_1106 (O_1106,N_14792,N_14812);
nor UO_1107 (O_1107,N_14797,N_14922);
nor UO_1108 (O_1108,N_14828,N_14804);
nor UO_1109 (O_1109,N_14850,N_14891);
nor UO_1110 (O_1110,N_14912,N_14765);
nor UO_1111 (O_1111,N_14916,N_14752);
nor UO_1112 (O_1112,N_14787,N_14937);
and UO_1113 (O_1113,N_14918,N_14956);
nand UO_1114 (O_1114,N_14769,N_14835);
nor UO_1115 (O_1115,N_14862,N_14912);
xnor UO_1116 (O_1116,N_14872,N_14942);
nand UO_1117 (O_1117,N_14774,N_14927);
and UO_1118 (O_1118,N_14843,N_14992);
or UO_1119 (O_1119,N_14900,N_14981);
nor UO_1120 (O_1120,N_14853,N_14918);
nand UO_1121 (O_1121,N_14854,N_14914);
and UO_1122 (O_1122,N_14941,N_14868);
nor UO_1123 (O_1123,N_14882,N_14905);
nor UO_1124 (O_1124,N_14970,N_14789);
xor UO_1125 (O_1125,N_14967,N_14810);
nand UO_1126 (O_1126,N_14754,N_14920);
nand UO_1127 (O_1127,N_14889,N_14871);
nand UO_1128 (O_1128,N_14916,N_14989);
or UO_1129 (O_1129,N_14980,N_14923);
or UO_1130 (O_1130,N_14999,N_14766);
nor UO_1131 (O_1131,N_14913,N_14892);
xor UO_1132 (O_1132,N_14838,N_14811);
nor UO_1133 (O_1133,N_14869,N_14846);
and UO_1134 (O_1134,N_14953,N_14990);
nor UO_1135 (O_1135,N_14973,N_14830);
and UO_1136 (O_1136,N_14793,N_14835);
or UO_1137 (O_1137,N_14832,N_14931);
or UO_1138 (O_1138,N_14923,N_14766);
nand UO_1139 (O_1139,N_14984,N_14987);
or UO_1140 (O_1140,N_14817,N_14800);
xor UO_1141 (O_1141,N_14930,N_14904);
nand UO_1142 (O_1142,N_14957,N_14757);
nor UO_1143 (O_1143,N_14844,N_14974);
nand UO_1144 (O_1144,N_14837,N_14949);
or UO_1145 (O_1145,N_14849,N_14854);
or UO_1146 (O_1146,N_14777,N_14879);
and UO_1147 (O_1147,N_14772,N_14891);
and UO_1148 (O_1148,N_14765,N_14965);
nor UO_1149 (O_1149,N_14993,N_14892);
and UO_1150 (O_1150,N_14796,N_14873);
and UO_1151 (O_1151,N_14953,N_14960);
or UO_1152 (O_1152,N_14795,N_14800);
nor UO_1153 (O_1153,N_14952,N_14839);
xnor UO_1154 (O_1154,N_14910,N_14750);
nand UO_1155 (O_1155,N_14873,N_14820);
nor UO_1156 (O_1156,N_14979,N_14800);
nor UO_1157 (O_1157,N_14967,N_14790);
nor UO_1158 (O_1158,N_14766,N_14893);
nor UO_1159 (O_1159,N_14853,N_14784);
or UO_1160 (O_1160,N_14859,N_14844);
nand UO_1161 (O_1161,N_14764,N_14908);
and UO_1162 (O_1162,N_14762,N_14943);
and UO_1163 (O_1163,N_14993,N_14895);
nand UO_1164 (O_1164,N_14978,N_14783);
or UO_1165 (O_1165,N_14768,N_14761);
nor UO_1166 (O_1166,N_14913,N_14786);
or UO_1167 (O_1167,N_14950,N_14761);
nand UO_1168 (O_1168,N_14773,N_14799);
or UO_1169 (O_1169,N_14957,N_14780);
nor UO_1170 (O_1170,N_14848,N_14888);
nor UO_1171 (O_1171,N_14964,N_14757);
and UO_1172 (O_1172,N_14759,N_14757);
nor UO_1173 (O_1173,N_14857,N_14753);
nand UO_1174 (O_1174,N_14953,N_14752);
nor UO_1175 (O_1175,N_14997,N_14934);
or UO_1176 (O_1176,N_14956,N_14914);
nor UO_1177 (O_1177,N_14907,N_14998);
or UO_1178 (O_1178,N_14909,N_14880);
or UO_1179 (O_1179,N_14803,N_14859);
nor UO_1180 (O_1180,N_14843,N_14790);
nor UO_1181 (O_1181,N_14813,N_14919);
nor UO_1182 (O_1182,N_14909,N_14762);
nor UO_1183 (O_1183,N_14969,N_14981);
nor UO_1184 (O_1184,N_14917,N_14985);
or UO_1185 (O_1185,N_14988,N_14822);
nand UO_1186 (O_1186,N_14757,N_14937);
nand UO_1187 (O_1187,N_14846,N_14993);
nand UO_1188 (O_1188,N_14781,N_14775);
nor UO_1189 (O_1189,N_14908,N_14956);
or UO_1190 (O_1190,N_14857,N_14943);
and UO_1191 (O_1191,N_14820,N_14754);
and UO_1192 (O_1192,N_14810,N_14791);
nand UO_1193 (O_1193,N_14870,N_14869);
nand UO_1194 (O_1194,N_14981,N_14977);
or UO_1195 (O_1195,N_14902,N_14799);
nor UO_1196 (O_1196,N_14766,N_14959);
nand UO_1197 (O_1197,N_14916,N_14844);
xnor UO_1198 (O_1198,N_14919,N_14824);
nand UO_1199 (O_1199,N_14889,N_14775);
or UO_1200 (O_1200,N_14869,N_14922);
nor UO_1201 (O_1201,N_14769,N_14896);
and UO_1202 (O_1202,N_14937,N_14804);
or UO_1203 (O_1203,N_14811,N_14862);
or UO_1204 (O_1204,N_14982,N_14937);
and UO_1205 (O_1205,N_14857,N_14867);
nand UO_1206 (O_1206,N_14840,N_14975);
and UO_1207 (O_1207,N_14903,N_14978);
and UO_1208 (O_1208,N_14867,N_14934);
nand UO_1209 (O_1209,N_14893,N_14953);
nand UO_1210 (O_1210,N_14934,N_14776);
and UO_1211 (O_1211,N_14885,N_14780);
xor UO_1212 (O_1212,N_14970,N_14997);
nand UO_1213 (O_1213,N_14775,N_14814);
or UO_1214 (O_1214,N_14834,N_14796);
nand UO_1215 (O_1215,N_14834,N_14822);
or UO_1216 (O_1216,N_14762,N_14929);
xor UO_1217 (O_1217,N_14811,N_14812);
nor UO_1218 (O_1218,N_14988,N_14825);
or UO_1219 (O_1219,N_14957,N_14997);
xor UO_1220 (O_1220,N_14764,N_14783);
nand UO_1221 (O_1221,N_14814,N_14770);
or UO_1222 (O_1222,N_14772,N_14999);
nand UO_1223 (O_1223,N_14943,N_14819);
nand UO_1224 (O_1224,N_14780,N_14879);
and UO_1225 (O_1225,N_14871,N_14966);
and UO_1226 (O_1226,N_14850,N_14977);
or UO_1227 (O_1227,N_14932,N_14964);
and UO_1228 (O_1228,N_14877,N_14824);
xnor UO_1229 (O_1229,N_14980,N_14993);
xor UO_1230 (O_1230,N_14814,N_14826);
nand UO_1231 (O_1231,N_14826,N_14964);
and UO_1232 (O_1232,N_14833,N_14998);
xnor UO_1233 (O_1233,N_14969,N_14858);
nand UO_1234 (O_1234,N_14803,N_14845);
nor UO_1235 (O_1235,N_14807,N_14898);
nor UO_1236 (O_1236,N_14838,N_14949);
and UO_1237 (O_1237,N_14956,N_14973);
or UO_1238 (O_1238,N_14915,N_14930);
nor UO_1239 (O_1239,N_14818,N_14867);
xor UO_1240 (O_1240,N_14866,N_14910);
or UO_1241 (O_1241,N_14768,N_14806);
or UO_1242 (O_1242,N_14952,N_14941);
or UO_1243 (O_1243,N_14779,N_14973);
nor UO_1244 (O_1244,N_14916,N_14968);
or UO_1245 (O_1245,N_14759,N_14858);
nand UO_1246 (O_1246,N_14825,N_14869);
nand UO_1247 (O_1247,N_14843,N_14782);
xnor UO_1248 (O_1248,N_14775,N_14997);
nor UO_1249 (O_1249,N_14858,N_14834);
or UO_1250 (O_1250,N_14887,N_14987);
nor UO_1251 (O_1251,N_14800,N_14977);
nor UO_1252 (O_1252,N_14918,N_14787);
xor UO_1253 (O_1253,N_14913,N_14990);
nor UO_1254 (O_1254,N_14961,N_14870);
nor UO_1255 (O_1255,N_14970,N_14769);
nor UO_1256 (O_1256,N_14862,N_14985);
nand UO_1257 (O_1257,N_14953,N_14908);
nand UO_1258 (O_1258,N_14807,N_14790);
nand UO_1259 (O_1259,N_14818,N_14970);
or UO_1260 (O_1260,N_14773,N_14916);
nand UO_1261 (O_1261,N_14789,N_14827);
or UO_1262 (O_1262,N_14862,N_14892);
nor UO_1263 (O_1263,N_14812,N_14859);
or UO_1264 (O_1264,N_14899,N_14802);
nand UO_1265 (O_1265,N_14899,N_14964);
xnor UO_1266 (O_1266,N_14987,N_14858);
nor UO_1267 (O_1267,N_14830,N_14833);
or UO_1268 (O_1268,N_14982,N_14998);
and UO_1269 (O_1269,N_14755,N_14955);
and UO_1270 (O_1270,N_14902,N_14944);
or UO_1271 (O_1271,N_14836,N_14877);
nor UO_1272 (O_1272,N_14751,N_14837);
nor UO_1273 (O_1273,N_14966,N_14787);
or UO_1274 (O_1274,N_14806,N_14823);
nor UO_1275 (O_1275,N_14914,N_14888);
nand UO_1276 (O_1276,N_14966,N_14789);
nor UO_1277 (O_1277,N_14992,N_14775);
nor UO_1278 (O_1278,N_14909,N_14848);
nor UO_1279 (O_1279,N_14783,N_14893);
and UO_1280 (O_1280,N_14912,N_14881);
and UO_1281 (O_1281,N_14830,N_14959);
or UO_1282 (O_1282,N_14751,N_14934);
and UO_1283 (O_1283,N_14772,N_14775);
nor UO_1284 (O_1284,N_14757,N_14798);
nor UO_1285 (O_1285,N_14968,N_14859);
nand UO_1286 (O_1286,N_14927,N_14901);
or UO_1287 (O_1287,N_14906,N_14781);
xnor UO_1288 (O_1288,N_14944,N_14855);
nand UO_1289 (O_1289,N_14966,N_14759);
xnor UO_1290 (O_1290,N_14773,N_14876);
or UO_1291 (O_1291,N_14833,N_14845);
nand UO_1292 (O_1292,N_14973,N_14965);
nor UO_1293 (O_1293,N_14957,N_14948);
xor UO_1294 (O_1294,N_14790,N_14752);
and UO_1295 (O_1295,N_14751,N_14882);
nor UO_1296 (O_1296,N_14869,N_14750);
xnor UO_1297 (O_1297,N_14963,N_14761);
and UO_1298 (O_1298,N_14890,N_14942);
nor UO_1299 (O_1299,N_14903,N_14785);
and UO_1300 (O_1300,N_14982,N_14757);
nand UO_1301 (O_1301,N_14806,N_14770);
xor UO_1302 (O_1302,N_14758,N_14923);
and UO_1303 (O_1303,N_14778,N_14768);
nor UO_1304 (O_1304,N_14918,N_14919);
or UO_1305 (O_1305,N_14771,N_14948);
nor UO_1306 (O_1306,N_14834,N_14924);
and UO_1307 (O_1307,N_14979,N_14771);
xnor UO_1308 (O_1308,N_14889,N_14845);
and UO_1309 (O_1309,N_14956,N_14781);
xnor UO_1310 (O_1310,N_14755,N_14821);
or UO_1311 (O_1311,N_14888,N_14986);
nor UO_1312 (O_1312,N_14835,N_14953);
nor UO_1313 (O_1313,N_14790,N_14971);
nor UO_1314 (O_1314,N_14887,N_14946);
nand UO_1315 (O_1315,N_14832,N_14834);
and UO_1316 (O_1316,N_14758,N_14907);
and UO_1317 (O_1317,N_14925,N_14932);
xnor UO_1318 (O_1318,N_14967,N_14890);
nand UO_1319 (O_1319,N_14768,N_14814);
or UO_1320 (O_1320,N_14943,N_14957);
or UO_1321 (O_1321,N_14903,N_14831);
nand UO_1322 (O_1322,N_14892,N_14755);
or UO_1323 (O_1323,N_14993,N_14913);
nor UO_1324 (O_1324,N_14860,N_14758);
xor UO_1325 (O_1325,N_14996,N_14959);
nand UO_1326 (O_1326,N_14767,N_14868);
xor UO_1327 (O_1327,N_14802,N_14788);
and UO_1328 (O_1328,N_14859,N_14949);
nand UO_1329 (O_1329,N_14937,N_14852);
or UO_1330 (O_1330,N_14911,N_14998);
nor UO_1331 (O_1331,N_14930,N_14787);
xnor UO_1332 (O_1332,N_14899,N_14857);
nor UO_1333 (O_1333,N_14830,N_14786);
and UO_1334 (O_1334,N_14782,N_14954);
nor UO_1335 (O_1335,N_14950,N_14923);
or UO_1336 (O_1336,N_14758,N_14913);
nor UO_1337 (O_1337,N_14889,N_14836);
and UO_1338 (O_1338,N_14946,N_14763);
nand UO_1339 (O_1339,N_14955,N_14977);
nor UO_1340 (O_1340,N_14991,N_14818);
and UO_1341 (O_1341,N_14945,N_14993);
nor UO_1342 (O_1342,N_14888,N_14931);
or UO_1343 (O_1343,N_14802,N_14847);
and UO_1344 (O_1344,N_14990,N_14977);
nor UO_1345 (O_1345,N_14802,N_14821);
xnor UO_1346 (O_1346,N_14808,N_14867);
nand UO_1347 (O_1347,N_14785,N_14793);
nor UO_1348 (O_1348,N_14789,N_14792);
or UO_1349 (O_1349,N_14754,N_14956);
nor UO_1350 (O_1350,N_14839,N_14953);
nand UO_1351 (O_1351,N_14962,N_14923);
and UO_1352 (O_1352,N_14930,N_14873);
nor UO_1353 (O_1353,N_14894,N_14754);
or UO_1354 (O_1354,N_14972,N_14940);
xor UO_1355 (O_1355,N_14971,N_14799);
nor UO_1356 (O_1356,N_14856,N_14751);
nor UO_1357 (O_1357,N_14931,N_14769);
and UO_1358 (O_1358,N_14948,N_14890);
or UO_1359 (O_1359,N_14756,N_14752);
or UO_1360 (O_1360,N_14759,N_14908);
xnor UO_1361 (O_1361,N_14826,N_14788);
and UO_1362 (O_1362,N_14823,N_14887);
and UO_1363 (O_1363,N_14835,N_14883);
nor UO_1364 (O_1364,N_14850,N_14919);
nand UO_1365 (O_1365,N_14866,N_14760);
nor UO_1366 (O_1366,N_14923,N_14769);
nand UO_1367 (O_1367,N_14834,N_14932);
or UO_1368 (O_1368,N_14856,N_14855);
and UO_1369 (O_1369,N_14791,N_14816);
nand UO_1370 (O_1370,N_14836,N_14853);
nand UO_1371 (O_1371,N_14829,N_14855);
and UO_1372 (O_1372,N_14866,N_14935);
and UO_1373 (O_1373,N_14830,N_14866);
or UO_1374 (O_1374,N_14914,N_14910);
and UO_1375 (O_1375,N_14750,N_14975);
and UO_1376 (O_1376,N_14949,N_14816);
or UO_1377 (O_1377,N_14885,N_14806);
or UO_1378 (O_1378,N_14775,N_14991);
nand UO_1379 (O_1379,N_14854,N_14760);
or UO_1380 (O_1380,N_14861,N_14937);
or UO_1381 (O_1381,N_14900,N_14950);
nor UO_1382 (O_1382,N_14998,N_14847);
and UO_1383 (O_1383,N_14761,N_14896);
nand UO_1384 (O_1384,N_14846,N_14923);
and UO_1385 (O_1385,N_14893,N_14821);
nand UO_1386 (O_1386,N_14885,N_14859);
and UO_1387 (O_1387,N_14940,N_14993);
and UO_1388 (O_1388,N_14994,N_14938);
nand UO_1389 (O_1389,N_14970,N_14945);
and UO_1390 (O_1390,N_14777,N_14904);
nor UO_1391 (O_1391,N_14923,N_14959);
nor UO_1392 (O_1392,N_14798,N_14814);
and UO_1393 (O_1393,N_14752,N_14830);
nand UO_1394 (O_1394,N_14922,N_14910);
and UO_1395 (O_1395,N_14965,N_14810);
or UO_1396 (O_1396,N_14926,N_14992);
or UO_1397 (O_1397,N_14993,N_14854);
or UO_1398 (O_1398,N_14832,N_14908);
nand UO_1399 (O_1399,N_14770,N_14787);
or UO_1400 (O_1400,N_14915,N_14754);
and UO_1401 (O_1401,N_14863,N_14826);
nand UO_1402 (O_1402,N_14784,N_14810);
nand UO_1403 (O_1403,N_14796,N_14757);
xor UO_1404 (O_1404,N_14816,N_14840);
and UO_1405 (O_1405,N_14958,N_14912);
and UO_1406 (O_1406,N_14965,N_14942);
nand UO_1407 (O_1407,N_14912,N_14764);
and UO_1408 (O_1408,N_14837,N_14912);
and UO_1409 (O_1409,N_14930,N_14777);
nor UO_1410 (O_1410,N_14771,N_14786);
and UO_1411 (O_1411,N_14958,N_14850);
nor UO_1412 (O_1412,N_14854,N_14773);
or UO_1413 (O_1413,N_14932,N_14825);
nor UO_1414 (O_1414,N_14754,N_14867);
or UO_1415 (O_1415,N_14918,N_14990);
xnor UO_1416 (O_1416,N_14974,N_14792);
xor UO_1417 (O_1417,N_14860,N_14853);
nor UO_1418 (O_1418,N_14952,N_14945);
or UO_1419 (O_1419,N_14949,N_14915);
nor UO_1420 (O_1420,N_14879,N_14867);
xnor UO_1421 (O_1421,N_14794,N_14806);
and UO_1422 (O_1422,N_14968,N_14760);
nor UO_1423 (O_1423,N_14874,N_14756);
or UO_1424 (O_1424,N_14994,N_14836);
nor UO_1425 (O_1425,N_14880,N_14882);
nand UO_1426 (O_1426,N_14830,N_14998);
or UO_1427 (O_1427,N_14765,N_14870);
nand UO_1428 (O_1428,N_14777,N_14823);
nand UO_1429 (O_1429,N_14957,N_14777);
and UO_1430 (O_1430,N_14913,N_14893);
and UO_1431 (O_1431,N_14953,N_14790);
nand UO_1432 (O_1432,N_14899,N_14878);
or UO_1433 (O_1433,N_14946,N_14789);
nand UO_1434 (O_1434,N_14917,N_14925);
and UO_1435 (O_1435,N_14781,N_14940);
or UO_1436 (O_1436,N_14793,N_14961);
or UO_1437 (O_1437,N_14968,N_14808);
and UO_1438 (O_1438,N_14948,N_14863);
and UO_1439 (O_1439,N_14909,N_14867);
xnor UO_1440 (O_1440,N_14847,N_14977);
xnor UO_1441 (O_1441,N_14901,N_14751);
and UO_1442 (O_1442,N_14954,N_14823);
nand UO_1443 (O_1443,N_14952,N_14876);
nand UO_1444 (O_1444,N_14914,N_14979);
or UO_1445 (O_1445,N_14997,N_14829);
and UO_1446 (O_1446,N_14944,N_14773);
nand UO_1447 (O_1447,N_14823,N_14797);
nand UO_1448 (O_1448,N_14806,N_14751);
xor UO_1449 (O_1449,N_14759,N_14894);
or UO_1450 (O_1450,N_14893,N_14898);
or UO_1451 (O_1451,N_14813,N_14945);
nand UO_1452 (O_1452,N_14801,N_14923);
or UO_1453 (O_1453,N_14943,N_14982);
or UO_1454 (O_1454,N_14869,N_14851);
and UO_1455 (O_1455,N_14951,N_14918);
or UO_1456 (O_1456,N_14765,N_14898);
nor UO_1457 (O_1457,N_14995,N_14951);
and UO_1458 (O_1458,N_14815,N_14848);
or UO_1459 (O_1459,N_14786,N_14755);
xor UO_1460 (O_1460,N_14858,N_14830);
nand UO_1461 (O_1461,N_14765,N_14909);
or UO_1462 (O_1462,N_14986,N_14875);
nor UO_1463 (O_1463,N_14959,N_14944);
and UO_1464 (O_1464,N_14817,N_14824);
xor UO_1465 (O_1465,N_14829,N_14922);
and UO_1466 (O_1466,N_14903,N_14813);
and UO_1467 (O_1467,N_14815,N_14766);
nand UO_1468 (O_1468,N_14836,N_14818);
xnor UO_1469 (O_1469,N_14989,N_14753);
nor UO_1470 (O_1470,N_14842,N_14890);
xnor UO_1471 (O_1471,N_14784,N_14936);
or UO_1472 (O_1472,N_14907,N_14929);
nor UO_1473 (O_1473,N_14906,N_14976);
xnor UO_1474 (O_1474,N_14829,N_14825);
and UO_1475 (O_1475,N_14821,N_14772);
and UO_1476 (O_1476,N_14773,N_14945);
nand UO_1477 (O_1477,N_14902,N_14860);
and UO_1478 (O_1478,N_14810,N_14771);
nor UO_1479 (O_1479,N_14991,N_14800);
nand UO_1480 (O_1480,N_14892,N_14922);
or UO_1481 (O_1481,N_14836,N_14936);
nand UO_1482 (O_1482,N_14966,N_14981);
or UO_1483 (O_1483,N_14791,N_14890);
nor UO_1484 (O_1484,N_14756,N_14996);
nand UO_1485 (O_1485,N_14840,N_14921);
nand UO_1486 (O_1486,N_14776,N_14978);
nand UO_1487 (O_1487,N_14927,N_14993);
nor UO_1488 (O_1488,N_14756,N_14949);
nor UO_1489 (O_1489,N_14829,N_14808);
nor UO_1490 (O_1490,N_14811,N_14911);
or UO_1491 (O_1491,N_14966,N_14965);
nor UO_1492 (O_1492,N_14919,N_14825);
nand UO_1493 (O_1493,N_14926,N_14800);
and UO_1494 (O_1494,N_14971,N_14873);
nand UO_1495 (O_1495,N_14829,N_14847);
or UO_1496 (O_1496,N_14944,N_14758);
nor UO_1497 (O_1497,N_14834,N_14767);
or UO_1498 (O_1498,N_14829,N_14965);
nand UO_1499 (O_1499,N_14766,N_14771);
nand UO_1500 (O_1500,N_14833,N_14898);
or UO_1501 (O_1501,N_14972,N_14952);
nand UO_1502 (O_1502,N_14923,N_14810);
and UO_1503 (O_1503,N_14813,N_14830);
or UO_1504 (O_1504,N_14862,N_14895);
and UO_1505 (O_1505,N_14876,N_14934);
nand UO_1506 (O_1506,N_14872,N_14999);
or UO_1507 (O_1507,N_14953,N_14963);
nor UO_1508 (O_1508,N_14838,N_14953);
nor UO_1509 (O_1509,N_14997,N_14915);
and UO_1510 (O_1510,N_14799,N_14939);
and UO_1511 (O_1511,N_14838,N_14913);
and UO_1512 (O_1512,N_14809,N_14800);
and UO_1513 (O_1513,N_14926,N_14866);
nor UO_1514 (O_1514,N_14873,N_14996);
nor UO_1515 (O_1515,N_14923,N_14993);
nor UO_1516 (O_1516,N_14756,N_14935);
and UO_1517 (O_1517,N_14785,N_14813);
or UO_1518 (O_1518,N_14950,N_14786);
or UO_1519 (O_1519,N_14903,N_14851);
or UO_1520 (O_1520,N_14961,N_14753);
and UO_1521 (O_1521,N_14958,N_14884);
nand UO_1522 (O_1522,N_14963,N_14857);
nand UO_1523 (O_1523,N_14768,N_14983);
nor UO_1524 (O_1524,N_14887,N_14814);
xor UO_1525 (O_1525,N_14766,N_14986);
xor UO_1526 (O_1526,N_14832,N_14848);
nand UO_1527 (O_1527,N_14916,N_14848);
and UO_1528 (O_1528,N_14996,N_14893);
nand UO_1529 (O_1529,N_14920,N_14997);
and UO_1530 (O_1530,N_14841,N_14766);
nor UO_1531 (O_1531,N_14769,N_14973);
nor UO_1532 (O_1532,N_14804,N_14784);
and UO_1533 (O_1533,N_14993,N_14938);
nor UO_1534 (O_1534,N_14918,N_14875);
nor UO_1535 (O_1535,N_14979,N_14839);
nand UO_1536 (O_1536,N_14941,N_14950);
nor UO_1537 (O_1537,N_14864,N_14991);
or UO_1538 (O_1538,N_14772,N_14895);
nand UO_1539 (O_1539,N_14963,N_14757);
and UO_1540 (O_1540,N_14944,N_14785);
nor UO_1541 (O_1541,N_14876,N_14937);
and UO_1542 (O_1542,N_14764,N_14985);
or UO_1543 (O_1543,N_14835,N_14789);
nor UO_1544 (O_1544,N_14937,N_14891);
or UO_1545 (O_1545,N_14802,N_14971);
or UO_1546 (O_1546,N_14875,N_14847);
nor UO_1547 (O_1547,N_14753,N_14943);
or UO_1548 (O_1548,N_14867,N_14771);
and UO_1549 (O_1549,N_14860,N_14914);
nand UO_1550 (O_1550,N_14977,N_14946);
or UO_1551 (O_1551,N_14928,N_14912);
nor UO_1552 (O_1552,N_14943,N_14806);
nor UO_1553 (O_1553,N_14807,N_14947);
nor UO_1554 (O_1554,N_14843,N_14987);
nor UO_1555 (O_1555,N_14989,N_14773);
xnor UO_1556 (O_1556,N_14882,N_14915);
nand UO_1557 (O_1557,N_14800,N_14864);
nand UO_1558 (O_1558,N_14815,N_14846);
xor UO_1559 (O_1559,N_14772,N_14878);
or UO_1560 (O_1560,N_14990,N_14789);
nand UO_1561 (O_1561,N_14848,N_14811);
nor UO_1562 (O_1562,N_14779,N_14958);
and UO_1563 (O_1563,N_14983,N_14857);
or UO_1564 (O_1564,N_14826,N_14939);
nor UO_1565 (O_1565,N_14849,N_14817);
and UO_1566 (O_1566,N_14774,N_14976);
xnor UO_1567 (O_1567,N_14755,N_14922);
nand UO_1568 (O_1568,N_14887,N_14991);
nor UO_1569 (O_1569,N_14802,N_14822);
nand UO_1570 (O_1570,N_14801,N_14776);
and UO_1571 (O_1571,N_14844,N_14965);
nor UO_1572 (O_1572,N_14858,N_14756);
xor UO_1573 (O_1573,N_14921,N_14796);
and UO_1574 (O_1574,N_14841,N_14941);
or UO_1575 (O_1575,N_14854,N_14996);
and UO_1576 (O_1576,N_14965,N_14945);
nand UO_1577 (O_1577,N_14793,N_14924);
nor UO_1578 (O_1578,N_14836,N_14861);
nand UO_1579 (O_1579,N_14813,N_14766);
and UO_1580 (O_1580,N_14900,N_14940);
xor UO_1581 (O_1581,N_14900,N_14954);
and UO_1582 (O_1582,N_14777,N_14915);
nand UO_1583 (O_1583,N_14943,N_14844);
or UO_1584 (O_1584,N_14796,N_14908);
xnor UO_1585 (O_1585,N_14939,N_14889);
nor UO_1586 (O_1586,N_14834,N_14803);
and UO_1587 (O_1587,N_14962,N_14931);
and UO_1588 (O_1588,N_14835,N_14969);
nand UO_1589 (O_1589,N_14853,N_14936);
and UO_1590 (O_1590,N_14827,N_14984);
nor UO_1591 (O_1591,N_14816,N_14912);
nor UO_1592 (O_1592,N_14851,N_14789);
or UO_1593 (O_1593,N_14985,N_14758);
nor UO_1594 (O_1594,N_14986,N_14814);
and UO_1595 (O_1595,N_14788,N_14842);
nor UO_1596 (O_1596,N_14943,N_14856);
nand UO_1597 (O_1597,N_14763,N_14961);
nand UO_1598 (O_1598,N_14925,N_14956);
or UO_1599 (O_1599,N_14820,N_14828);
or UO_1600 (O_1600,N_14974,N_14801);
and UO_1601 (O_1601,N_14875,N_14965);
nor UO_1602 (O_1602,N_14885,N_14755);
nor UO_1603 (O_1603,N_14996,N_14943);
nor UO_1604 (O_1604,N_14863,N_14807);
and UO_1605 (O_1605,N_14783,N_14883);
or UO_1606 (O_1606,N_14903,N_14977);
and UO_1607 (O_1607,N_14765,N_14865);
nor UO_1608 (O_1608,N_14780,N_14875);
or UO_1609 (O_1609,N_14841,N_14947);
or UO_1610 (O_1610,N_14869,N_14891);
or UO_1611 (O_1611,N_14795,N_14866);
or UO_1612 (O_1612,N_14973,N_14774);
or UO_1613 (O_1613,N_14920,N_14923);
or UO_1614 (O_1614,N_14779,N_14990);
nor UO_1615 (O_1615,N_14863,N_14865);
nand UO_1616 (O_1616,N_14784,N_14769);
nand UO_1617 (O_1617,N_14939,N_14781);
nor UO_1618 (O_1618,N_14991,N_14927);
nor UO_1619 (O_1619,N_14795,N_14889);
nor UO_1620 (O_1620,N_14943,N_14822);
or UO_1621 (O_1621,N_14821,N_14876);
or UO_1622 (O_1622,N_14774,N_14805);
nand UO_1623 (O_1623,N_14780,N_14753);
xnor UO_1624 (O_1624,N_14997,N_14764);
or UO_1625 (O_1625,N_14775,N_14768);
xor UO_1626 (O_1626,N_14904,N_14774);
and UO_1627 (O_1627,N_14905,N_14881);
or UO_1628 (O_1628,N_14889,N_14927);
or UO_1629 (O_1629,N_14838,N_14863);
nor UO_1630 (O_1630,N_14761,N_14964);
and UO_1631 (O_1631,N_14864,N_14901);
nand UO_1632 (O_1632,N_14975,N_14768);
and UO_1633 (O_1633,N_14890,N_14924);
and UO_1634 (O_1634,N_14820,N_14835);
xnor UO_1635 (O_1635,N_14988,N_14767);
and UO_1636 (O_1636,N_14995,N_14795);
and UO_1637 (O_1637,N_14856,N_14888);
and UO_1638 (O_1638,N_14898,N_14757);
or UO_1639 (O_1639,N_14754,N_14950);
or UO_1640 (O_1640,N_14782,N_14957);
or UO_1641 (O_1641,N_14992,N_14827);
nand UO_1642 (O_1642,N_14808,N_14783);
nor UO_1643 (O_1643,N_14915,N_14940);
nand UO_1644 (O_1644,N_14794,N_14838);
or UO_1645 (O_1645,N_14984,N_14801);
nor UO_1646 (O_1646,N_14761,N_14894);
and UO_1647 (O_1647,N_14841,N_14780);
nor UO_1648 (O_1648,N_14780,N_14847);
nand UO_1649 (O_1649,N_14843,N_14759);
nor UO_1650 (O_1650,N_14879,N_14882);
or UO_1651 (O_1651,N_14947,N_14894);
or UO_1652 (O_1652,N_14812,N_14804);
and UO_1653 (O_1653,N_14758,N_14794);
nand UO_1654 (O_1654,N_14901,N_14936);
or UO_1655 (O_1655,N_14826,N_14883);
nand UO_1656 (O_1656,N_14818,N_14823);
and UO_1657 (O_1657,N_14786,N_14807);
nand UO_1658 (O_1658,N_14893,N_14831);
and UO_1659 (O_1659,N_14957,N_14962);
and UO_1660 (O_1660,N_14923,N_14893);
or UO_1661 (O_1661,N_14754,N_14982);
nor UO_1662 (O_1662,N_14819,N_14842);
or UO_1663 (O_1663,N_14911,N_14934);
nand UO_1664 (O_1664,N_14761,N_14908);
nor UO_1665 (O_1665,N_14835,N_14784);
and UO_1666 (O_1666,N_14891,N_14750);
and UO_1667 (O_1667,N_14817,N_14873);
nor UO_1668 (O_1668,N_14763,N_14841);
nor UO_1669 (O_1669,N_14950,N_14840);
nand UO_1670 (O_1670,N_14807,N_14988);
nor UO_1671 (O_1671,N_14777,N_14959);
xor UO_1672 (O_1672,N_14839,N_14801);
nand UO_1673 (O_1673,N_14801,N_14992);
and UO_1674 (O_1674,N_14925,N_14955);
nand UO_1675 (O_1675,N_14983,N_14814);
nor UO_1676 (O_1676,N_14949,N_14846);
nand UO_1677 (O_1677,N_14946,N_14760);
or UO_1678 (O_1678,N_14788,N_14973);
nor UO_1679 (O_1679,N_14801,N_14781);
and UO_1680 (O_1680,N_14894,N_14755);
or UO_1681 (O_1681,N_14854,N_14969);
or UO_1682 (O_1682,N_14973,N_14923);
or UO_1683 (O_1683,N_14850,N_14896);
or UO_1684 (O_1684,N_14931,N_14874);
or UO_1685 (O_1685,N_14952,N_14953);
and UO_1686 (O_1686,N_14752,N_14844);
nand UO_1687 (O_1687,N_14891,N_14922);
nor UO_1688 (O_1688,N_14899,N_14824);
and UO_1689 (O_1689,N_14801,N_14894);
and UO_1690 (O_1690,N_14991,N_14875);
nor UO_1691 (O_1691,N_14904,N_14841);
and UO_1692 (O_1692,N_14935,N_14863);
nor UO_1693 (O_1693,N_14924,N_14919);
or UO_1694 (O_1694,N_14894,N_14797);
or UO_1695 (O_1695,N_14974,N_14881);
nand UO_1696 (O_1696,N_14776,N_14827);
nand UO_1697 (O_1697,N_14780,N_14766);
nand UO_1698 (O_1698,N_14939,N_14943);
and UO_1699 (O_1699,N_14824,N_14797);
nor UO_1700 (O_1700,N_14960,N_14811);
or UO_1701 (O_1701,N_14863,N_14903);
nand UO_1702 (O_1702,N_14779,N_14757);
nor UO_1703 (O_1703,N_14800,N_14989);
and UO_1704 (O_1704,N_14904,N_14979);
nor UO_1705 (O_1705,N_14964,N_14779);
and UO_1706 (O_1706,N_14876,N_14954);
and UO_1707 (O_1707,N_14766,N_14996);
xor UO_1708 (O_1708,N_14894,N_14897);
and UO_1709 (O_1709,N_14899,N_14768);
and UO_1710 (O_1710,N_14926,N_14750);
or UO_1711 (O_1711,N_14989,N_14942);
and UO_1712 (O_1712,N_14800,N_14857);
nand UO_1713 (O_1713,N_14894,N_14906);
nor UO_1714 (O_1714,N_14807,N_14900);
nand UO_1715 (O_1715,N_14986,N_14900);
or UO_1716 (O_1716,N_14910,N_14958);
xnor UO_1717 (O_1717,N_14938,N_14970);
nor UO_1718 (O_1718,N_14786,N_14956);
or UO_1719 (O_1719,N_14989,N_14877);
and UO_1720 (O_1720,N_14887,N_14864);
or UO_1721 (O_1721,N_14906,N_14832);
or UO_1722 (O_1722,N_14948,N_14953);
nand UO_1723 (O_1723,N_14823,N_14812);
and UO_1724 (O_1724,N_14844,N_14848);
xnor UO_1725 (O_1725,N_14973,N_14835);
nor UO_1726 (O_1726,N_14855,N_14867);
nand UO_1727 (O_1727,N_14914,N_14798);
and UO_1728 (O_1728,N_14946,N_14953);
nor UO_1729 (O_1729,N_14794,N_14855);
nand UO_1730 (O_1730,N_14843,N_14897);
nor UO_1731 (O_1731,N_14915,N_14955);
nor UO_1732 (O_1732,N_14992,N_14909);
nand UO_1733 (O_1733,N_14948,N_14968);
nand UO_1734 (O_1734,N_14853,N_14868);
or UO_1735 (O_1735,N_14778,N_14833);
nand UO_1736 (O_1736,N_14831,N_14973);
nand UO_1737 (O_1737,N_14755,N_14753);
xnor UO_1738 (O_1738,N_14897,N_14953);
xnor UO_1739 (O_1739,N_14872,N_14833);
or UO_1740 (O_1740,N_14957,N_14988);
nor UO_1741 (O_1741,N_14803,N_14945);
nand UO_1742 (O_1742,N_14889,N_14819);
or UO_1743 (O_1743,N_14813,N_14786);
nor UO_1744 (O_1744,N_14975,N_14885);
nand UO_1745 (O_1745,N_14963,N_14892);
and UO_1746 (O_1746,N_14974,N_14775);
or UO_1747 (O_1747,N_14857,N_14922);
and UO_1748 (O_1748,N_14895,N_14910);
nor UO_1749 (O_1749,N_14761,N_14781);
nor UO_1750 (O_1750,N_14827,N_14879);
and UO_1751 (O_1751,N_14950,N_14913);
nor UO_1752 (O_1752,N_14795,N_14982);
xnor UO_1753 (O_1753,N_14842,N_14930);
or UO_1754 (O_1754,N_14824,N_14884);
nand UO_1755 (O_1755,N_14860,N_14943);
or UO_1756 (O_1756,N_14859,N_14847);
or UO_1757 (O_1757,N_14900,N_14777);
or UO_1758 (O_1758,N_14889,N_14908);
nand UO_1759 (O_1759,N_14855,N_14924);
nand UO_1760 (O_1760,N_14905,N_14954);
and UO_1761 (O_1761,N_14954,N_14770);
and UO_1762 (O_1762,N_14895,N_14790);
and UO_1763 (O_1763,N_14889,N_14812);
nor UO_1764 (O_1764,N_14985,N_14785);
nand UO_1765 (O_1765,N_14868,N_14962);
or UO_1766 (O_1766,N_14908,N_14994);
nor UO_1767 (O_1767,N_14774,N_14771);
nor UO_1768 (O_1768,N_14859,N_14862);
nor UO_1769 (O_1769,N_14972,N_14852);
and UO_1770 (O_1770,N_14769,N_14855);
nor UO_1771 (O_1771,N_14890,N_14997);
xnor UO_1772 (O_1772,N_14994,N_14843);
and UO_1773 (O_1773,N_14856,N_14950);
nor UO_1774 (O_1774,N_14774,N_14983);
and UO_1775 (O_1775,N_14785,N_14831);
and UO_1776 (O_1776,N_14841,N_14823);
or UO_1777 (O_1777,N_14848,N_14891);
nand UO_1778 (O_1778,N_14787,N_14923);
xor UO_1779 (O_1779,N_14755,N_14941);
or UO_1780 (O_1780,N_14935,N_14899);
xnor UO_1781 (O_1781,N_14917,N_14930);
nand UO_1782 (O_1782,N_14940,N_14922);
xnor UO_1783 (O_1783,N_14914,N_14931);
or UO_1784 (O_1784,N_14907,N_14911);
xor UO_1785 (O_1785,N_14877,N_14984);
or UO_1786 (O_1786,N_14845,N_14771);
and UO_1787 (O_1787,N_14775,N_14955);
nand UO_1788 (O_1788,N_14886,N_14941);
and UO_1789 (O_1789,N_14956,N_14929);
and UO_1790 (O_1790,N_14883,N_14887);
xnor UO_1791 (O_1791,N_14996,N_14821);
nand UO_1792 (O_1792,N_14849,N_14910);
nand UO_1793 (O_1793,N_14892,N_14880);
or UO_1794 (O_1794,N_14762,N_14752);
nand UO_1795 (O_1795,N_14884,N_14860);
and UO_1796 (O_1796,N_14788,N_14836);
and UO_1797 (O_1797,N_14969,N_14923);
nand UO_1798 (O_1798,N_14994,N_14893);
or UO_1799 (O_1799,N_14924,N_14850);
nor UO_1800 (O_1800,N_14976,N_14855);
or UO_1801 (O_1801,N_14768,N_14941);
and UO_1802 (O_1802,N_14804,N_14963);
xnor UO_1803 (O_1803,N_14822,N_14887);
xnor UO_1804 (O_1804,N_14825,N_14854);
nor UO_1805 (O_1805,N_14750,N_14967);
nor UO_1806 (O_1806,N_14797,N_14888);
nor UO_1807 (O_1807,N_14965,N_14899);
nand UO_1808 (O_1808,N_14811,N_14898);
nor UO_1809 (O_1809,N_14797,N_14958);
nand UO_1810 (O_1810,N_14803,N_14928);
and UO_1811 (O_1811,N_14918,N_14891);
nor UO_1812 (O_1812,N_14774,N_14961);
and UO_1813 (O_1813,N_14883,N_14814);
or UO_1814 (O_1814,N_14855,N_14838);
nor UO_1815 (O_1815,N_14855,N_14880);
xnor UO_1816 (O_1816,N_14982,N_14911);
nor UO_1817 (O_1817,N_14868,N_14934);
or UO_1818 (O_1818,N_14806,N_14756);
xnor UO_1819 (O_1819,N_14887,N_14861);
and UO_1820 (O_1820,N_14766,N_14799);
nand UO_1821 (O_1821,N_14905,N_14829);
nor UO_1822 (O_1822,N_14889,N_14891);
or UO_1823 (O_1823,N_14794,N_14813);
nand UO_1824 (O_1824,N_14776,N_14937);
and UO_1825 (O_1825,N_14958,N_14865);
nor UO_1826 (O_1826,N_14793,N_14807);
or UO_1827 (O_1827,N_14884,N_14957);
and UO_1828 (O_1828,N_14801,N_14977);
nand UO_1829 (O_1829,N_14888,N_14950);
and UO_1830 (O_1830,N_14987,N_14836);
or UO_1831 (O_1831,N_14875,N_14985);
and UO_1832 (O_1832,N_14810,N_14907);
nor UO_1833 (O_1833,N_14757,N_14848);
and UO_1834 (O_1834,N_14897,N_14957);
or UO_1835 (O_1835,N_14990,N_14935);
xor UO_1836 (O_1836,N_14752,N_14981);
or UO_1837 (O_1837,N_14947,N_14800);
or UO_1838 (O_1838,N_14930,N_14783);
or UO_1839 (O_1839,N_14817,N_14944);
nand UO_1840 (O_1840,N_14951,N_14793);
nor UO_1841 (O_1841,N_14996,N_14841);
nand UO_1842 (O_1842,N_14897,N_14800);
nor UO_1843 (O_1843,N_14943,N_14862);
nand UO_1844 (O_1844,N_14786,N_14846);
and UO_1845 (O_1845,N_14904,N_14770);
or UO_1846 (O_1846,N_14943,N_14813);
and UO_1847 (O_1847,N_14862,N_14783);
and UO_1848 (O_1848,N_14806,N_14988);
nand UO_1849 (O_1849,N_14960,N_14972);
nor UO_1850 (O_1850,N_14826,N_14753);
xor UO_1851 (O_1851,N_14848,N_14806);
xor UO_1852 (O_1852,N_14980,N_14977);
or UO_1853 (O_1853,N_14764,N_14844);
or UO_1854 (O_1854,N_14901,N_14763);
and UO_1855 (O_1855,N_14989,N_14866);
nor UO_1856 (O_1856,N_14963,N_14971);
nor UO_1857 (O_1857,N_14801,N_14924);
nor UO_1858 (O_1858,N_14927,N_14830);
and UO_1859 (O_1859,N_14856,N_14916);
nand UO_1860 (O_1860,N_14959,N_14933);
nand UO_1861 (O_1861,N_14906,N_14841);
nand UO_1862 (O_1862,N_14983,N_14810);
or UO_1863 (O_1863,N_14948,N_14826);
nor UO_1864 (O_1864,N_14762,N_14781);
or UO_1865 (O_1865,N_14855,N_14823);
nand UO_1866 (O_1866,N_14826,N_14881);
nor UO_1867 (O_1867,N_14967,N_14782);
or UO_1868 (O_1868,N_14772,N_14860);
nor UO_1869 (O_1869,N_14821,N_14935);
nor UO_1870 (O_1870,N_14813,N_14997);
and UO_1871 (O_1871,N_14781,N_14826);
nand UO_1872 (O_1872,N_14959,N_14895);
or UO_1873 (O_1873,N_14786,N_14836);
nor UO_1874 (O_1874,N_14769,N_14817);
and UO_1875 (O_1875,N_14972,N_14883);
nor UO_1876 (O_1876,N_14810,N_14778);
nor UO_1877 (O_1877,N_14941,N_14839);
nor UO_1878 (O_1878,N_14986,N_14780);
nand UO_1879 (O_1879,N_14946,N_14839);
nor UO_1880 (O_1880,N_14841,N_14900);
nand UO_1881 (O_1881,N_14933,N_14929);
and UO_1882 (O_1882,N_14882,N_14750);
or UO_1883 (O_1883,N_14941,N_14979);
nor UO_1884 (O_1884,N_14810,N_14812);
nand UO_1885 (O_1885,N_14802,N_14951);
and UO_1886 (O_1886,N_14889,N_14848);
nand UO_1887 (O_1887,N_14980,N_14848);
nand UO_1888 (O_1888,N_14896,N_14847);
nand UO_1889 (O_1889,N_14833,N_14785);
nand UO_1890 (O_1890,N_14913,N_14826);
nor UO_1891 (O_1891,N_14893,N_14855);
or UO_1892 (O_1892,N_14875,N_14792);
nand UO_1893 (O_1893,N_14804,N_14914);
nor UO_1894 (O_1894,N_14805,N_14883);
nor UO_1895 (O_1895,N_14898,N_14904);
nand UO_1896 (O_1896,N_14854,N_14945);
nand UO_1897 (O_1897,N_14844,N_14803);
nand UO_1898 (O_1898,N_14965,N_14922);
and UO_1899 (O_1899,N_14864,N_14984);
and UO_1900 (O_1900,N_14894,N_14795);
and UO_1901 (O_1901,N_14887,N_14755);
and UO_1902 (O_1902,N_14822,N_14776);
or UO_1903 (O_1903,N_14852,N_14962);
xnor UO_1904 (O_1904,N_14904,N_14975);
and UO_1905 (O_1905,N_14810,N_14946);
nand UO_1906 (O_1906,N_14847,N_14858);
nor UO_1907 (O_1907,N_14879,N_14914);
xor UO_1908 (O_1908,N_14833,N_14985);
or UO_1909 (O_1909,N_14797,N_14995);
or UO_1910 (O_1910,N_14886,N_14882);
xnor UO_1911 (O_1911,N_14885,N_14758);
or UO_1912 (O_1912,N_14945,N_14876);
and UO_1913 (O_1913,N_14823,N_14781);
or UO_1914 (O_1914,N_14866,N_14940);
nand UO_1915 (O_1915,N_14887,N_14844);
xnor UO_1916 (O_1916,N_14886,N_14869);
nand UO_1917 (O_1917,N_14922,N_14990);
nand UO_1918 (O_1918,N_14791,N_14875);
and UO_1919 (O_1919,N_14922,N_14906);
or UO_1920 (O_1920,N_14816,N_14937);
or UO_1921 (O_1921,N_14906,N_14752);
and UO_1922 (O_1922,N_14852,N_14801);
and UO_1923 (O_1923,N_14763,N_14872);
nand UO_1924 (O_1924,N_14967,N_14850);
nand UO_1925 (O_1925,N_14824,N_14976);
nand UO_1926 (O_1926,N_14944,N_14877);
and UO_1927 (O_1927,N_14868,N_14837);
or UO_1928 (O_1928,N_14775,N_14947);
nand UO_1929 (O_1929,N_14790,N_14863);
nor UO_1930 (O_1930,N_14795,N_14962);
nor UO_1931 (O_1931,N_14905,N_14926);
nand UO_1932 (O_1932,N_14762,N_14850);
or UO_1933 (O_1933,N_14762,N_14977);
nor UO_1934 (O_1934,N_14775,N_14765);
nand UO_1935 (O_1935,N_14866,N_14927);
and UO_1936 (O_1936,N_14796,N_14770);
nand UO_1937 (O_1937,N_14838,N_14784);
and UO_1938 (O_1938,N_14756,N_14937);
or UO_1939 (O_1939,N_14838,N_14809);
and UO_1940 (O_1940,N_14944,N_14958);
or UO_1941 (O_1941,N_14842,N_14780);
nand UO_1942 (O_1942,N_14884,N_14798);
nand UO_1943 (O_1943,N_14993,N_14791);
and UO_1944 (O_1944,N_14751,N_14791);
nor UO_1945 (O_1945,N_14899,N_14772);
nand UO_1946 (O_1946,N_14994,N_14806);
nor UO_1947 (O_1947,N_14756,N_14872);
nor UO_1948 (O_1948,N_14850,N_14822);
or UO_1949 (O_1949,N_14823,N_14865);
xnor UO_1950 (O_1950,N_14819,N_14798);
or UO_1951 (O_1951,N_14792,N_14803);
nor UO_1952 (O_1952,N_14859,N_14908);
nor UO_1953 (O_1953,N_14762,N_14997);
or UO_1954 (O_1954,N_14847,N_14890);
nand UO_1955 (O_1955,N_14789,N_14901);
nand UO_1956 (O_1956,N_14787,N_14939);
or UO_1957 (O_1957,N_14970,N_14812);
nor UO_1958 (O_1958,N_14758,N_14827);
and UO_1959 (O_1959,N_14761,N_14757);
nand UO_1960 (O_1960,N_14949,N_14831);
or UO_1961 (O_1961,N_14936,N_14807);
or UO_1962 (O_1962,N_14966,N_14917);
nor UO_1963 (O_1963,N_14807,N_14782);
nand UO_1964 (O_1964,N_14772,N_14836);
nand UO_1965 (O_1965,N_14835,N_14907);
or UO_1966 (O_1966,N_14857,N_14969);
and UO_1967 (O_1967,N_14868,N_14870);
or UO_1968 (O_1968,N_14950,N_14812);
nor UO_1969 (O_1969,N_14982,N_14897);
and UO_1970 (O_1970,N_14938,N_14991);
nand UO_1971 (O_1971,N_14794,N_14995);
or UO_1972 (O_1972,N_14806,N_14843);
and UO_1973 (O_1973,N_14865,N_14963);
and UO_1974 (O_1974,N_14924,N_14851);
nor UO_1975 (O_1975,N_14863,N_14806);
nor UO_1976 (O_1976,N_14752,N_14828);
or UO_1977 (O_1977,N_14986,N_14974);
nand UO_1978 (O_1978,N_14800,N_14942);
nand UO_1979 (O_1979,N_14759,N_14924);
nand UO_1980 (O_1980,N_14810,N_14773);
nand UO_1981 (O_1981,N_14941,N_14856);
or UO_1982 (O_1982,N_14807,N_14982);
and UO_1983 (O_1983,N_14856,N_14790);
nand UO_1984 (O_1984,N_14896,N_14821);
nand UO_1985 (O_1985,N_14881,N_14807);
nor UO_1986 (O_1986,N_14804,N_14781);
nand UO_1987 (O_1987,N_14913,N_14911);
or UO_1988 (O_1988,N_14923,N_14905);
and UO_1989 (O_1989,N_14785,N_14994);
nand UO_1990 (O_1990,N_14946,N_14891);
xor UO_1991 (O_1991,N_14954,N_14826);
xor UO_1992 (O_1992,N_14999,N_14889);
nand UO_1993 (O_1993,N_14877,N_14819);
and UO_1994 (O_1994,N_14857,N_14955);
nand UO_1995 (O_1995,N_14925,N_14804);
or UO_1996 (O_1996,N_14826,N_14810);
xnor UO_1997 (O_1997,N_14797,N_14972);
nand UO_1998 (O_1998,N_14886,N_14897);
and UO_1999 (O_1999,N_14833,N_14957);
endmodule