module basic_2000_20000_2500_4_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_952,In_1837);
and U1 (N_1,In_469,In_1632);
or U2 (N_2,In_473,In_1502);
nand U3 (N_3,In_634,In_1101);
nand U4 (N_4,In_1533,In_1259);
nand U5 (N_5,In_38,In_1759);
nand U6 (N_6,In_116,In_1740);
nor U7 (N_7,In_1854,In_321);
or U8 (N_8,In_1080,In_1076);
nand U9 (N_9,In_13,In_175);
nand U10 (N_10,In_584,In_316);
nor U11 (N_11,In_1399,In_564);
or U12 (N_12,In_1816,In_1771);
or U13 (N_13,In_1321,In_797);
and U14 (N_14,In_260,In_1234);
nor U15 (N_15,In_711,In_544);
nand U16 (N_16,In_1784,In_1249);
and U17 (N_17,In_1901,In_1332);
or U18 (N_18,In_842,In_16);
or U19 (N_19,In_1801,In_747);
and U20 (N_20,In_1810,In_1135);
nand U21 (N_21,In_30,In_1876);
or U22 (N_22,In_1731,In_1229);
xor U23 (N_23,In_1443,In_895);
nor U24 (N_24,In_247,In_1405);
and U25 (N_25,In_1576,In_1956);
nand U26 (N_26,In_1213,In_1573);
or U27 (N_27,In_188,In_1543);
and U28 (N_28,In_306,In_365);
and U29 (N_29,In_1083,In_411);
nor U30 (N_30,In_231,In_796);
nor U31 (N_31,In_1774,In_1808);
xor U32 (N_32,In_309,In_1850);
or U33 (N_33,In_616,In_680);
or U34 (N_34,In_1544,In_1966);
and U35 (N_35,In_1785,In_465);
and U36 (N_36,In_751,In_1115);
nor U37 (N_37,In_1000,In_204);
nor U38 (N_38,In_479,In_1219);
or U39 (N_39,In_613,In_1097);
and U40 (N_40,In_1651,In_1176);
nand U41 (N_41,In_427,In_1335);
nand U42 (N_42,In_1730,In_1839);
nor U43 (N_43,In_72,In_612);
and U44 (N_44,In_1160,In_605);
or U45 (N_45,In_1548,In_445);
or U46 (N_46,In_1471,In_1189);
xor U47 (N_47,In_386,In_658);
nor U48 (N_48,In_970,In_1993);
nand U49 (N_49,In_1001,In_1981);
nor U50 (N_50,In_641,In_755);
xor U51 (N_51,In_665,In_210);
nor U52 (N_52,In_166,In_1346);
nand U53 (N_53,In_1900,In_899);
nand U54 (N_54,In_1647,In_891);
and U55 (N_55,In_481,In_1223);
or U56 (N_56,In_1968,In_1077);
and U57 (N_57,In_1663,In_1032);
nand U58 (N_58,In_1324,In_381);
xor U59 (N_59,In_397,In_1062);
and U60 (N_60,In_829,In_1309);
or U61 (N_61,In_578,In_1407);
or U62 (N_62,In_32,In_1737);
nand U63 (N_63,In_207,In_1211);
or U64 (N_64,In_938,In_1979);
nand U65 (N_65,In_396,In_927);
or U66 (N_66,In_81,In_34);
and U67 (N_67,In_832,In_1939);
or U68 (N_68,In_1949,In_1743);
xnor U69 (N_69,In_1996,In_252);
nor U70 (N_70,In_1387,In_1316);
or U71 (N_71,In_1148,In_1575);
nand U72 (N_72,In_1398,In_663);
nand U73 (N_73,In_1437,In_686);
xor U74 (N_74,In_284,In_1447);
nand U75 (N_75,In_884,In_651);
nand U76 (N_76,In_524,In_698);
nor U77 (N_77,In_319,In_240);
and U78 (N_78,In_1764,In_1403);
nor U79 (N_79,In_111,In_1931);
nor U80 (N_80,In_810,In_1865);
and U81 (N_81,In_881,In_1012);
xor U82 (N_82,In_1216,In_290);
nand U83 (N_83,In_985,In_681);
or U84 (N_84,In_1884,In_967);
nor U85 (N_85,In_323,In_1120);
and U86 (N_86,In_1936,In_898);
nand U87 (N_87,In_901,In_1685);
nand U88 (N_88,In_189,In_1645);
and U89 (N_89,In_1727,In_174);
xnor U90 (N_90,In_569,In_308);
nand U91 (N_91,In_617,In_1087);
nand U92 (N_92,In_1152,In_1819);
and U93 (N_93,In_1442,In_645);
nand U94 (N_94,In_464,In_706);
nor U95 (N_95,In_1440,In_248);
nor U96 (N_96,In_1190,In_1976);
and U97 (N_97,In_1043,In_1869);
or U98 (N_98,In_1519,In_588);
xnor U99 (N_99,In_1756,In_347);
nor U100 (N_100,In_349,In_1380);
or U101 (N_101,In_1674,In_948);
nor U102 (N_102,In_60,In_442);
xor U103 (N_103,In_449,In_1276);
nor U104 (N_104,In_380,In_440);
nand U105 (N_105,In_1297,In_137);
nor U106 (N_106,In_1849,In_114);
and U107 (N_107,In_1497,In_1615);
or U108 (N_108,In_1212,In_1893);
nand U109 (N_109,In_1323,In_1425);
and U110 (N_110,In_1233,In_1796);
nand U111 (N_111,In_1170,In_705);
and U112 (N_112,In_1603,In_275);
nand U113 (N_113,In_1365,In_1953);
or U114 (N_114,In_811,In_1943);
nand U115 (N_115,In_305,In_601);
and U116 (N_116,In_619,In_1776);
and U117 (N_117,In_1593,In_778);
nor U118 (N_118,In_1726,In_932);
nand U119 (N_119,In_1518,In_725);
nor U120 (N_120,In_192,In_483);
or U121 (N_121,In_1495,In_912);
nor U122 (N_122,In_1048,In_693);
or U123 (N_123,In_872,In_656);
nand U124 (N_124,In_905,In_520);
or U125 (N_125,In_1879,In_138);
nand U126 (N_126,In_1070,In_1011);
and U127 (N_127,In_450,In_956);
or U128 (N_128,In_1252,In_1183);
and U129 (N_129,In_550,In_211);
xnor U130 (N_130,In_1227,In_1315);
and U131 (N_131,In_1192,In_1264);
nor U132 (N_132,In_1624,In_1626);
xor U133 (N_133,In_190,In_1988);
nand U134 (N_134,In_1842,In_89);
nand U135 (N_135,In_1618,In_1721);
nand U136 (N_136,In_1684,In_866);
nor U137 (N_137,In_74,In_625);
or U138 (N_138,In_106,In_730);
xor U139 (N_139,In_1374,In_43);
nand U140 (N_140,In_1607,In_103);
and U141 (N_141,In_1421,In_278);
or U142 (N_142,In_1970,In_1975);
nand U143 (N_143,In_1580,In_1178);
or U144 (N_144,In_186,In_598);
or U145 (N_145,In_1058,In_764);
and U146 (N_146,In_1741,In_997);
nand U147 (N_147,In_21,In_406);
nand U148 (N_148,In_1292,In_921);
nand U149 (N_149,In_24,In_1814);
xnor U150 (N_150,In_906,In_48);
nand U151 (N_151,In_592,In_992);
or U152 (N_152,In_262,In_1073);
or U153 (N_153,In_156,In_456);
nand U154 (N_154,In_892,In_1959);
or U155 (N_155,In_1559,In_1706);
xor U156 (N_156,In_1817,In_1751);
nor U157 (N_157,In_1408,In_1824);
xnor U158 (N_158,In_1995,In_707);
and U159 (N_159,In_1286,In_1431);
nand U160 (N_160,In_1017,In_1778);
nor U161 (N_161,In_1605,In_1599);
or U162 (N_162,In_926,In_1830);
nor U163 (N_163,In_1827,In_1753);
and U164 (N_164,In_1551,In_41);
or U165 (N_165,In_1232,In_261);
or U166 (N_166,In_1793,In_990);
or U167 (N_167,In_1415,In_514);
and U168 (N_168,In_1838,In_194);
nor U169 (N_169,In_315,In_461);
and U170 (N_170,In_991,In_903);
nor U171 (N_171,In_80,In_12);
and U172 (N_172,In_947,In_241);
and U173 (N_173,In_1341,In_417);
and U174 (N_174,In_814,In_131);
and U175 (N_175,In_1350,In_1345);
nor U176 (N_176,In_923,In_1973);
or U177 (N_177,In_1504,In_236);
xor U178 (N_178,In_1373,In_225);
or U179 (N_179,In_1794,In_1804);
nand U180 (N_180,In_1111,In_431);
or U181 (N_181,In_324,In_696);
or U182 (N_182,In_1182,In_1283);
nand U183 (N_183,In_1719,In_610);
and U184 (N_184,In_1694,In_945);
or U185 (N_185,In_1485,In_750);
or U186 (N_186,In_1195,In_1840);
nor U187 (N_187,In_420,In_975);
xor U188 (N_188,In_372,In_1466);
nand U189 (N_189,In_1113,In_512);
nand U190 (N_190,In_673,In_1517);
nor U191 (N_191,In_56,In_1265);
and U192 (N_192,In_1298,In_685);
and U193 (N_193,In_1745,In_1285);
nand U194 (N_194,In_1700,In_233);
or U195 (N_195,In_1688,In_142);
or U196 (N_196,In_541,In_1185);
and U197 (N_197,In_1733,In_1263);
xnor U198 (N_198,In_909,In_1649);
xnor U199 (N_199,In_561,In_1646);
or U200 (N_200,In_351,In_82);
xnor U201 (N_201,In_1660,In_1846);
nor U202 (N_202,In_425,In_198);
nor U203 (N_203,In_1456,In_375);
nand U204 (N_204,In_684,In_1319);
nor U205 (N_205,In_1452,In_851);
nor U206 (N_206,In_793,In_503);
and U207 (N_207,In_1567,In_966);
or U208 (N_208,In_476,In_1812);
or U209 (N_209,In_19,In_1037);
or U210 (N_210,In_650,In_1918);
and U211 (N_211,In_232,In_1556);
and U212 (N_212,In_678,In_1457);
or U213 (N_213,In_484,In_1507);
nand U214 (N_214,In_462,In_1678);
nand U215 (N_215,In_1354,In_58);
nand U216 (N_216,In_354,In_1424);
or U217 (N_217,In_1149,In_1029);
nor U218 (N_218,In_1188,In_1867);
nand U219 (N_219,In_1067,In_618);
and U220 (N_220,In_206,In_430);
nand U221 (N_221,In_1873,In_1179);
nand U222 (N_222,In_1811,In_1175);
nor U223 (N_223,In_727,In_558);
nor U224 (N_224,In_1327,In_1041);
nor U225 (N_225,In_1033,In_1522);
xnor U226 (N_226,In_1699,In_127);
nor U227 (N_227,In_1384,In_1308);
or U228 (N_228,In_113,In_91);
nor U229 (N_229,In_890,In_1198);
nand U230 (N_230,In_914,In_1571);
nand U231 (N_231,In_378,In_629);
or U232 (N_232,In_1503,In_1419);
nor U233 (N_233,In_410,In_120);
xor U234 (N_234,In_587,In_1542);
and U235 (N_235,In_129,In_666);
nand U236 (N_236,In_435,In_1617);
and U237 (N_237,In_875,In_1791);
or U238 (N_238,In_1102,In_871);
nor U239 (N_239,In_408,In_245);
nand U240 (N_240,In_243,In_1498);
nor U241 (N_241,In_852,In_766);
and U242 (N_242,In_322,In_969);
nor U243 (N_243,In_653,In_786);
and U244 (N_244,In_459,In_1564);
and U245 (N_245,In_29,In_398);
nor U246 (N_246,In_864,In_830);
or U247 (N_247,In_1402,In_1831);
nand U248 (N_248,In_1171,In_787);
nand U249 (N_249,In_1236,In_489);
nand U250 (N_250,In_1353,In_1271);
and U251 (N_251,In_326,In_1707);
or U252 (N_252,In_212,In_1393);
and U253 (N_253,In_1269,In_862);
nand U254 (N_254,In_1281,In_385);
or U255 (N_255,In_295,In_259);
nor U256 (N_256,In_35,In_1716);
nand U257 (N_257,In_888,In_155);
and U258 (N_258,In_345,In_218);
nand U259 (N_259,In_414,In_1693);
or U260 (N_260,In_159,In_1932);
nand U261 (N_261,In_320,In_1834);
nor U262 (N_262,In_216,In_1557);
nor U263 (N_263,In_1255,In_1347);
nor U264 (N_264,In_533,In_50);
or U265 (N_265,In_1763,In_1206);
nand U266 (N_266,In_1038,In_671);
nand U267 (N_267,In_760,In_158);
nor U268 (N_268,In_615,In_729);
nor U269 (N_269,In_1383,In_1449);
nand U270 (N_270,In_1818,In_1691);
and U271 (N_271,In_500,In_920);
xor U272 (N_272,In_946,In_1018);
and U273 (N_273,In_1366,In_603);
and U274 (N_274,In_807,In_1851);
or U275 (N_275,In_1057,In_1463);
and U276 (N_276,In_1583,In_736);
and U277 (N_277,In_1007,In_1952);
or U278 (N_278,In_1193,In_1585);
xor U279 (N_279,In_1493,In_443);
or U280 (N_280,In_1775,In_602);
xnor U281 (N_281,In_1145,In_105);
nor U282 (N_282,In_1333,In_874);
and U283 (N_283,In_69,In_1406);
and U284 (N_284,In_530,In_1781);
nand U285 (N_285,In_1156,In_1779);
and U286 (N_286,In_1862,In_1967);
nand U287 (N_287,In_1099,In_935);
or U288 (N_288,In_1279,In_1910);
and U289 (N_289,In_1954,In_1060);
nand U290 (N_290,In_1620,In_759);
or U291 (N_291,In_774,In_944);
nand U292 (N_292,In_1124,In_1322);
or U293 (N_293,In_387,In_1307);
or U294 (N_294,In_348,In_229);
nand U295 (N_295,In_715,In_1871);
and U296 (N_296,In_1946,In_998);
and U297 (N_297,In_1301,In_1004);
nor U298 (N_298,In_543,In_694);
or U299 (N_299,In_502,In_203);
or U300 (N_300,In_513,In_1908);
nor U301 (N_301,In_336,In_1116);
nand U302 (N_302,In_1539,In_826);
or U303 (N_303,In_373,In_144);
nor U304 (N_304,In_1377,In_1100);
nand U305 (N_305,In_1250,In_1054);
nor U306 (N_306,In_940,In_963);
and U307 (N_307,In_1205,In_487);
nand U308 (N_308,In_1597,In_1143);
xnor U309 (N_309,In_1983,In_1509);
and U310 (N_310,In_1439,In_1010);
or U311 (N_311,In_767,In_1181);
or U312 (N_312,In_754,In_1467);
nor U313 (N_313,In_1359,In_1653);
and U314 (N_314,In_1065,In_640);
nor U315 (N_315,In_688,In_84);
or U316 (N_316,In_1595,In_813);
xor U317 (N_317,In_1251,In_258);
or U318 (N_318,In_1878,In_1174);
xnor U319 (N_319,In_1072,In_393);
nand U320 (N_320,In_1411,In_1492);
xnor U321 (N_321,In_889,In_1891);
nand U322 (N_322,In_642,In_517);
or U323 (N_323,In_1560,In_1516);
or U324 (N_324,In_1465,In_894);
nand U325 (N_325,In_904,In_734);
xnor U326 (N_326,In_1325,In_434);
nand U327 (N_327,In_1390,In_1698);
and U328 (N_328,In_402,In_1969);
or U329 (N_329,In_1683,In_745);
or U330 (N_330,In_1147,In_1242);
and U331 (N_331,In_107,In_97);
nand U332 (N_332,In_1549,In_1805);
nand U333 (N_333,In_556,In_1627);
nand U334 (N_334,In_96,In_497);
nor U335 (N_335,In_1623,In_820);
nor U336 (N_336,In_572,In_1885);
xnor U337 (N_337,In_1608,In_1562);
xor U338 (N_338,In_1864,In_1534);
nand U339 (N_339,In_1306,In_823);
nor U340 (N_340,In_1362,In_873);
xor U341 (N_341,In_1899,In_1351);
and U342 (N_342,In_1226,In_1270);
nor U343 (N_343,In_1266,In_853);
and U344 (N_344,In_1843,In_758);
nand U345 (N_345,In_1766,In_1880);
nor U346 (N_346,In_1948,In_224);
nand U347 (N_347,In_837,In_1014);
nand U348 (N_348,In_59,In_682);
and U349 (N_349,In_1059,In_1277);
nor U350 (N_350,In_257,In_700);
and U351 (N_351,In_1815,In_1022);
or U352 (N_352,In_528,In_1082);
xor U353 (N_353,In_1146,In_37);
nor U354 (N_354,In_1222,In_1039);
nor U355 (N_355,In_1356,In_600);
nand U356 (N_356,In_539,In_1877);
nand U357 (N_357,In_1882,In_215);
and U358 (N_358,In_547,In_1629);
or U359 (N_359,In_1550,In_827);
or U360 (N_360,In_560,In_292);
nand U361 (N_361,In_646,In_1413);
and U362 (N_362,In_800,In_1273);
nand U363 (N_363,In_1462,In_576);
nand U364 (N_364,In_1600,In_1122);
and U365 (N_365,In_1589,In_636);
xnor U366 (N_366,In_31,In_1888);
and U367 (N_367,In_92,In_761);
nor U368 (N_368,In_1761,In_1809);
xnor U369 (N_369,In_1150,In_1521);
nor U370 (N_370,In_1584,In_104);
nand U371 (N_371,In_1904,In_1246);
nand U372 (N_372,In_1806,In_1566);
nand U373 (N_373,In_1875,In_1933);
xnor U374 (N_374,In_1847,In_1254);
nand U375 (N_375,In_1085,In_1606);
nand U376 (N_376,In_296,In_644);
or U377 (N_377,In_987,In_1244);
or U378 (N_378,In_657,In_1477);
nand U379 (N_379,In_1289,In_993);
or U380 (N_380,In_1758,In_586);
or U381 (N_381,In_263,In_496);
nand U382 (N_382,In_633,In_1527);
nor U383 (N_383,In_1772,In_762);
nand U384 (N_384,In_731,In_317);
or U385 (N_385,In_1529,In_546);
or U386 (N_386,In_128,In_819);
and U387 (N_387,In_1020,In_1302);
xnor U388 (N_388,In_112,In_1381);
or U389 (N_389,In_169,In_1166);
or U390 (N_390,In_1820,In_28);
and U391 (N_391,In_328,In_799);
nor U392 (N_392,In_1395,In_432);
nand U393 (N_393,In_125,In_1228);
nand U394 (N_394,In_209,In_1734);
or U395 (N_395,In_1868,In_630);
nand U396 (N_396,In_1369,In_1639);
nand U397 (N_397,In_220,In_1168);
nor U398 (N_398,In_101,In_358);
nand U399 (N_399,In_62,In_1971);
nor U400 (N_400,In_1505,In_495);
nand U401 (N_401,In_1690,In_357);
and U402 (N_402,In_720,In_1767);
or U403 (N_403,In_749,In_1677);
nor U404 (N_404,In_781,In_1090);
nor U405 (N_405,In_1670,In_1340);
nor U406 (N_406,In_907,In_1538);
nor U407 (N_407,In_519,In_170);
or U408 (N_408,In_669,In_264);
nor U409 (N_409,In_1494,In_1379);
or U410 (N_410,In_1614,In_1616);
nor U411 (N_411,In_1628,In_173);
nor U412 (N_412,In_185,In_1499);
and U413 (N_413,In_1450,In_925);
and U414 (N_414,In_360,In_803);
nand U415 (N_415,In_1655,In_708);
nand U416 (N_416,In_1990,In_157);
or U417 (N_417,In_1787,In_376);
nor U418 (N_418,In_1042,In_1024);
or U419 (N_419,In_861,In_1960);
and U420 (N_420,In_1291,In_1201);
or U421 (N_421,In_954,In_1320);
xnor U422 (N_422,In_33,In_1044);
nor U423 (N_423,In_330,In_860);
and U424 (N_424,In_674,In_458);
and U425 (N_425,In_1780,In_1392);
nor U426 (N_426,In_704,In_1063);
nand U427 (N_427,In_1069,In_99);
or U428 (N_428,In_775,In_1129);
and U429 (N_429,In_716,In_670);
xor U430 (N_430,In_1460,In_516);
or U431 (N_431,In_983,In_1164);
nand U432 (N_432,In_1305,In_937);
nand U433 (N_433,In_250,In_893);
or U434 (N_434,In_858,In_549);
xor U435 (N_435,In_989,In_1955);
or U436 (N_436,In_1797,In_64);
nand U437 (N_437,In_746,In_1487);
nor U438 (N_438,In_222,In_1610);
or U439 (N_439,In_1695,In_1829);
or U440 (N_440,In_167,In_1679);
nand U441 (N_441,In_1235,In_1386);
or U442 (N_442,In_39,In_1261);
nor U443 (N_443,In_585,In_312);
or U444 (N_444,In_1681,In_1375);
nand U445 (N_445,In_1441,In_701);
nand U446 (N_446,In_49,In_44);
and U447 (N_447,In_563,In_54);
nand U448 (N_448,In_1587,In_1105);
and U449 (N_449,In_959,In_559);
nand U450 (N_450,In_1984,In_943);
nor U451 (N_451,In_178,In_1293);
nor U452 (N_452,In_1611,In_119);
nor U453 (N_453,In_1654,In_1747);
xnor U454 (N_454,In_1709,In_726);
and U455 (N_455,In_311,In_3);
nor U456 (N_456,In_573,In_1574);
and U457 (N_457,In_597,In_457);
or U458 (N_458,In_1664,In_1930);
nand U459 (N_459,In_335,In_1427);
or U460 (N_460,In_302,In_333);
or U461 (N_461,In_1397,In_980);
or U462 (N_462,In_1015,In_1112);
or U463 (N_463,In_1673,In_647);
nand U464 (N_464,In_423,In_608);
and U465 (N_465,In_499,In_313);
nor U466 (N_466,In_1601,In_249);
and U467 (N_467,In_1723,In_460);
xnor U468 (N_468,In_87,In_208);
nand U469 (N_469,In_659,In_353);
nor U470 (N_470,In_1652,In_643);
xor U471 (N_471,In_1546,In_1312);
nand U472 (N_472,In_1500,In_46);
nor U473 (N_473,In_1053,In_1712);
and U474 (N_474,In_1874,In_1659);
nor U475 (N_475,In_1897,In_824);
nor U476 (N_476,In_1895,In_1991);
nor U477 (N_477,In_1098,In_140);
nor U478 (N_478,In_395,In_57);
or U479 (N_479,In_964,In_817);
nand U480 (N_480,In_83,In_1777);
and U481 (N_481,In_692,In_1974);
nor U482 (N_482,In_1890,In_565);
nand U483 (N_483,In_783,In_1468);
or U484 (N_484,In_702,In_555);
and U485 (N_485,In_409,In_620);
nor U486 (N_486,In_883,In_1453);
or U487 (N_487,In_1414,In_865);
or U488 (N_488,In_147,In_623);
xnor U489 (N_489,In_1472,In_374);
and U490 (N_490,In_534,In_1330);
nor U491 (N_491,In_867,In_1448);
and U492 (N_492,In_1750,In_1328);
xor U493 (N_493,In_283,In_538);
nand U494 (N_494,In_815,In_477);
and U495 (N_495,In_1803,In_132);
and U496 (N_496,In_1945,In_974);
nand U497 (N_497,In_255,In_1861);
nor U498 (N_498,In_63,In_1672);
or U499 (N_499,In_67,In_1376);
and U500 (N_500,In_5,In_280);
xor U501 (N_501,In_1071,In_223);
nor U502 (N_502,In_366,In_294);
nor U503 (N_503,In_235,In_1568);
nand U504 (N_504,In_1857,In_1385);
nor U505 (N_505,In_1138,In_471);
and U506 (N_506,In_679,In_878);
nor U507 (N_507,In_1096,In_1360);
nor U508 (N_508,In_1592,In_1718);
or U509 (N_509,In_788,In_1262);
and U510 (N_510,In_428,In_929);
nand U511 (N_511,In_453,In_770);
nor U512 (N_512,In_802,In_982);
nor U513 (N_513,In_269,In_1121);
and U514 (N_514,In_593,In_1410);
or U515 (N_515,In_1056,In_1896);
and U516 (N_516,In_1558,In_581);
or U517 (N_517,In_86,In_1903);
nand U518 (N_518,In_370,In_1355);
nor U519 (N_519,In_994,In_1125);
nand U520 (N_520,In_1735,In_117);
and U521 (N_521,In_1378,In_340);
nor U522 (N_522,In_1088,In_1641);
and U523 (N_523,In_467,In_1537);
and U524 (N_524,In_273,In_1714);
or U525 (N_525,In_379,In_631);
nor U526 (N_526,In_145,In_1520);
nor U527 (N_527,In_789,In_1977);
or U528 (N_528,In_1144,In_822);
or U529 (N_529,In_1963,In_1525);
or U530 (N_530,In_438,In_661);
nor U531 (N_531,In_540,In_1886);
and U532 (N_532,In_1926,In_299);
or U533 (N_533,In_924,In_859);
or U534 (N_534,In_1613,In_1907);
nor U535 (N_535,In_1079,In_1922);
nor U536 (N_536,In_1528,In_522);
or U537 (N_537,In_1086,In_654);
or U538 (N_538,In_621,In_752);
nand U539 (N_539,In_568,In_66);
or U540 (N_540,In_896,In_1489);
nor U541 (N_541,In_1091,In_535);
xnor U542 (N_542,In_1303,In_768);
or U543 (N_543,In_1760,In_902);
nor U544 (N_544,In_1095,In_677);
nor U545 (N_545,In_844,In_908);
nor U546 (N_546,In_868,In_1339);
nand U547 (N_547,In_1515,In_1640);
or U548 (N_548,In_234,In_1540);
nor U549 (N_549,In_371,In_1940);
xnor U550 (N_550,In_1496,In_548);
or U551 (N_551,In_352,In_1935);
nor U552 (N_552,In_582,In_798);
nand U553 (N_553,In_1417,In_607);
and U554 (N_554,In_933,In_426);
nor U555 (N_555,In_1469,In_337);
nor U556 (N_556,In_1972,In_532);
nor U557 (N_557,In_304,In_492);
nand U558 (N_558,In_1184,In_415);
nor U559 (N_559,In_668,In_196);
nor U560 (N_560,In_1807,In_1581);
nand U561 (N_561,In_849,In_1795);
or U562 (N_562,In_739,In_136);
or U563 (N_563,In_551,In_1128);
nand U564 (N_564,In_331,In_272);
and U565 (N_565,In_1635,In_356);
nand U566 (N_566,In_782,In_1161);
or U567 (N_567,In_1980,In_737);
nand U568 (N_568,In_1326,In_1074);
nand U569 (N_569,In_1866,In_1169);
or U570 (N_570,In_1582,In_447);
and U571 (N_571,In_1506,In_575);
and U572 (N_572,In_1591,In_1118);
and U573 (N_573,In_75,In_237);
nand U574 (N_574,In_1482,In_191);
nor U575 (N_575,In_288,In_1898);
xor U576 (N_576,In_525,In_1009);
or U577 (N_577,In_1370,In_845);
and U578 (N_578,In_88,In_1268);
and U579 (N_579,In_675,In_960);
nor U580 (N_580,In_4,In_772);
nor U581 (N_581,In_553,In_1633);
nor U582 (N_582,In_1430,In_161);
nor U583 (N_583,In_291,In_1371);
and U584 (N_584,In_1158,In_1314);
and U585 (N_585,In_687,In_595);
or U586 (N_586,In_554,In_419);
nand U587 (N_587,In_1770,In_1987);
and U588 (N_588,In_809,In_1925);
nor U589 (N_589,In_795,In_1662);
and U590 (N_590,In_298,In_1045);
or U591 (N_591,In_199,In_808);
or U592 (N_592,In_1713,In_79);
or U593 (N_593,In_1196,In_1428);
or U594 (N_594,In_1965,In_1892);
or U595 (N_595,In_1692,In_804);
nor U596 (N_596,In_949,In_1746);
and U597 (N_597,In_401,In_1363);
and U598 (N_598,In_100,In_6);
or U599 (N_599,In_1650,In_361);
nand U600 (N_600,In_1026,In_1941);
and U601 (N_601,In_1950,In_327);
nand U602 (N_602,In_1081,In_286);
and U603 (N_603,In_1142,In_1224);
nor U604 (N_604,In_171,In_1207);
nand U605 (N_605,In_15,In_1409);
and U606 (N_606,In_254,In_486);
or U607 (N_607,In_1982,In_470);
nand U608 (N_608,In_639,In_1642);
xnor U609 (N_609,In_1648,In_652);
or U610 (N_610,In_1177,In_1909);
nor U611 (N_611,In_165,In_490);
nor U612 (N_612,In_1686,In_1511);
nand U613 (N_613,In_1172,In_452);
and U614 (N_614,In_1075,In_1400);
nor U615 (N_615,In_1401,In_1738);
nor U616 (N_616,In_146,In_339);
or U617 (N_617,In_1295,In_1790);
xor U618 (N_618,In_879,In_400);
or U619 (N_619,In_1768,In_1258);
and U620 (N_620,In_856,In_391);
nand U621 (N_621,In_805,In_529);
and U622 (N_622,In_1028,In_1636);
and U623 (N_623,In_76,In_98);
and U624 (N_624,In_1555,In_149);
nand U625 (N_625,In_662,In_1241);
and U626 (N_626,In_1526,In_279);
and U627 (N_627,In_968,In_466);
nor U628 (N_628,In_256,In_979);
and U629 (N_629,In_1300,In_162);
xor U630 (N_630,In_880,In_297);
or U631 (N_631,In_53,In_1438);
and U632 (N_632,In_1724,In_1331);
or U633 (N_633,In_1221,In_270);
or U634 (N_634,In_1123,In_183);
xor U635 (N_635,In_816,In_1786);
or U636 (N_636,In_1284,In_510);
xor U637 (N_637,In_493,In_433);
or U638 (N_638,In_506,In_509);
and U639 (N_639,In_742,In_1924);
xnor U640 (N_640,In_1051,In_801);
nand U641 (N_641,In_124,In_1962);
nor U642 (N_642,In_1214,In_61);
or U643 (N_643,In_1047,In_1396);
nor U644 (N_644,In_1906,In_1203);
nor U645 (N_645,In_118,In_965);
xor U646 (N_646,In_1513,In_1119);
or U647 (N_647,In_1154,In_1202);
or U648 (N_648,In_1913,In_1696);
nor U649 (N_649,In_300,In_1434);
xnor U650 (N_650,In_205,In_771);
nor U651 (N_651,In_709,In_628);
or U652 (N_652,In_870,In_999);
or U653 (N_653,In_121,In_78);
nor U654 (N_654,In_1491,In_835);
or U655 (N_655,In_246,In_1773);
or U656 (N_656,In_115,In_455);
or U657 (N_657,In_1986,In_1025);
and U658 (N_658,In_1682,In_1199);
and U659 (N_659,In_1501,In_1357);
nand U660 (N_660,In_1631,In_404);
xnor U661 (N_661,In_776,In_722);
nand U662 (N_662,In_367,In_1133);
or U663 (N_663,In_1288,In_168);
nor U664 (N_664,In_251,In_648);
nand U665 (N_665,In_1050,In_1132);
and U666 (N_666,In_743,In_1958);
or U667 (N_667,In_1535,In_1313);
and U668 (N_668,In_580,In_1103);
and U669 (N_669,In_672,In_1416);
nand U670 (N_670,In_936,In_285);
and U671 (N_671,In_986,In_1915);
or U672 (N_672,In_265,In_1749);
and U673 (N_673,In_910,In_1708);
xnor U674 (N_674,In_1828,In_536);
nand U675 (N_675,In_271,In_1141);
nand U676 (N_676,In_1887,In_887);
nand U677 (N_677,In_193,In_537);
or U678 (N_678,In_436,In_26);
nand U679 (N_679,In_735,In_266);
nand U680 (N_680,In_1554,In_1570);
xnor U681 (N_681,In_1563,In_70);
nor U682 (N_682,In_507,In_472);
and U683 (N_683,In_1036,In_717);
xor U684 (N_684,In_1272,In_1588);
nand U685 (N_685,In_343,In_531);
nand U686 (N_686,In_638,In_85);
and U687 (N_687,In_1689,In_1167);
or U688 (N_688,In_570,In_1464);
xor U689 (N_689,In_769,In_916);
and U690 (N_690,In_1136,In_1137);
or U691 (N_691,In_1094,In_150);
nor U692 (N_692,In_1225,In_785);
or U693 (N_693,In_1703,In_599);
nand U694 (N_694,In_133,In_40);
or U695 (N_695,In_1577,In_579);
nor U696 (N_696,In_1093,In_7);
nor U697 (N_697,In_995,In_1078);
xor U698 (N_698,In_821,In_624);
xnor U699 (N_699,In_1789,In_448);
or U700 (N_700,In_1274,In_1013);
and U701 (N_701,In_482,In_915);
and U702 (N_702,In_939,In_1919);
xor U703 (N_703,In_429,In_377);
nor U704 (N_704,In_383,In_451);
or U705 (N_705,In_413,In_972);
nor U706 (N_706,In_1243,In_289);
and U707 (N_707,In_840,In_1792);
nor U708 (N_708,In_958,In_130);
nor U709 (N_709,In_1478,In_931);
or U710 (N_710,In_1002,In_757);
and U711 (N_711,In_863,In_622);
and U712 (N_712,In_1210,In_1030);
nand U713 (N_713,In_344,In_1368);
nor U714 (N_714,In_1479,In_1016);
nand U715 (N_715,In_143,In_981);
or U716 (N_716,In_421,In_36);
nor U717 (N_717,In_342,In_1998);
or U718 (N_718,In_1151,In_1267);
nand U719 (N_719,In_17,In_139);
or U720 (N_720,In_42,In_1134);
nor U721 (N_721,In_1938,In_1429);
or U722 (N_722,In_1841,In_1204);
and U723 (N_723,In_1569,In_690);
or U724 (N_724,In_1622,In_1619);
nor U725 (N_725,In_825,In_854);
nor U726 (N_726,In_1348,In_664);
nor U727 (N_727,In_1928,In_833);
or U728 (N_728,In_494,In_1055);
nand U729 (N_729,In_1832,In_221);
nand U730 (N_730,In_1643,In_1657);
or U731 (N_731,In_346,In_267);
nor U732 (N_732,In_163,In_1609);
xnor U733 (N_733,In_1826,In_1344);
or U734 (N_734,In_1006,In_846);
nand U735 (N_735,In_1461,In_562);
xnor U736 (N_736,In_791,In_1475);
and U737 (N_737,In_748,In_388);
nor U738 (N_738,In_527,In_1621);
nor U739 (N_739,In_1473,In_876);
and U740 (N_740,In_187,In_697);
nor U741 (N_741,In_90,In_474);
or U742 (N_742,In_1736,In_1389);
nor U743 (N_743,In_504,In_1697);
nor U744 (N_744,In_1231,In_1294);
or U745 (N_745,In_282,In_1765);
nand U746 (N_746,In_18,In_1068);
or U747 (N_747,In_399,In_1338);
nand U748 (N_748,In_1310,In_1994);
or U749 (N_749,In_869,In_1131);
xor U750 (N_750,In_122,In_744);
nor U751 (N_751,In_738,In_134);
nand U752 (N_752,In_971,In_407);
and U753 (N_753,In_885,In_918);
xor U754 (N_754,In_984,In_1848);
nor U755 (N_755,In_703,In_1420);
and U756 (N_756,In_596,In_1604);
nor U757 (N_757,In_1139,In_649);
and U758 (N_758,In_1412,In_1257);
nor U759 (N_759,In_1126,In_710);
nand U760 (N_760,In_1187,In_1432);
nand U761 (N_761,In_8,In_94);
or U762 (N_762,In_201,In_913);
xnor U763 (N_763,In_1547,In_1114);
or U764 (N_764,In_1658,In_1239);
and U765 (N_765,In_253,In_1256);
nor U766 (N_766,In_1799,In_1107);
and U767 (N_767,In_1046,In_1);
or U768 (N_768,In_996,In_1422);
nand U769 (N_769,In_164,In_1917);
nor U770 (N_770,In_52,In_1863);
or U771 (N_771,In_1667,In_363);
nor U772 (N_772,In_779,In_1092);
and U773 (N_773,In_2,In_691);
and U774 (N_774,In_51,In_721);
and U775 (N_775,In_160,In_355);
or U776 (N_776,In_1732,In_1844);
or U777 (N_777,In_1218,In_1989);
nand U778 (N_778,In_733,In_604);
and U779 (N_779,In_491,In_545);
or U780 (N_780,In_1858,In_1701);
or U781 (N_781,In_73,In_1754);
or U782 (N_782,In_521,In_77);
and U783 (N_783,In_1578,In_1426);
and U784 (N_784,In_405,In_526);
and U785 (N_785,In_1311,In_1194);
or U786 (N_786,In_1927,In_1349);
nand U787 (N_787,In_1705,In_1937);
and U788 (N_788,In_14,In_784);
nand U789 (N_789,In_1836,In_179);
nor U790 (N_790,In_515,In_184);
and U791 (N_791,In_740,In_325);
or U792 (N_792,In_1602,In_1852);
nand U793 (N_793,In_1027,In_110);
or U794 (N_794,In_594,In_928);
nor U795 (N_795,In_850,In_1680);
or U796 (N_796,In_1480,In_1524);
nor U797 (N_797,In_153,In_1744);
nand U798 (N_798,In_1835,In_818);
and U799 (N_799,In_1717,In_1590);
nor U800 (N_800,In_389,In_847);
and U801 (N_801,In_1755,In_557);
nand U802 (N_802,In_418,In_955);
nand U803 (N_803,In_1883,In_714);
nand U804 (N_804,In_571,In_268);
and U805 (N_805,In_338,In_1748);
nor U806 (N_806,In_828,In_1275);
xnor U807 (N_807,In_609,In_329);
or U808 (N_808,In_1317,In_1404);
nand U809 (N_809,In_723,In_790);
and U810 (N_810,In_542,In_1008);
nor U811 (N_811,In_444,In_577);
and U812 (N_812,In_314,In_1436);
and U813 (N_813,In_1372,In_446);
xor U814 (N_814,In_1661,In_1444);
nand U815 (N_815,In_362,In_1586);
xnor U816 (N_816,In_177,In_911);
nand U817 (N_817,In_437,In_468);
nor U818 (N_818,In_1612,In_1367);
or U819 (N_819,In_68,In_412);
or U820 (N_820,In_219,In_1565);
and U821 (N_821,In_200,In_95);
nor U822 (N_822,In_422,In_65);
and U823 (N_823,In_1536,In_518);
nor U824 (N_824,In_839,In_773);
nor U825 (N_825,In_1418,In_1318);
nand U826 (N_826,In_977,In_359);
or U827 (N_827,In_1035,In_831);
and U828 (N_828,In_27,In_1725);
nand U829 (N_829,In_392,In_281);
or U830 (N_830,In_1455,In_1488);
xnor U831 (N_831,In_463,In_1157);
xnor U832 (N_832,In_202,In_403);
and U833 (N_833,In_976,In_1561);
nor U834 (N_834,In_382,In_1364);
or U835 (N_835,In_390,In_1382);
nor U836 (N_836,In_1752,In_1089);
nor U837 (N_837,In_485,In_897);
nand U838 (N_838,In_877,In_334);
and U839 (N_839,In_1061,In_368);
and U840 (N_840,In_838,In_857);
nor U841 (N_841,In_1066,In_765);
or U842 (N_842,In_1579,In_1108);
and U843 (N_843,In_699,In_1474);
nor U844 (N_844,In_1675,In_1530);
nand U845 (N_845,In_1220,In_1870);
and U846 (N_846,In_180,In_1783);
nor U847 (N_847,In_741,In_611);
nor U848 (N_848,In_1215,In_1914);
nor U849 (N_849,In_1729,In_109);
nor U850 (N_850,In_942,In_1021);
and U851 (N_851,In_919,In_1911);
or U852 (N_852,In_1304,In_1514);
and U853 (N_853,In_9,In_1757);
nor U854 (N_854,In_1833,In_1034);
xor U855 (N_855,In_1019,In_900);
nor U856 (N_856,In_1625,In_1961);
or U857 (N_857,In_384,In_480);
nor U858 (N_858,In_1802,In_0);
nand U859 (N_859,In_1905,In_718);
and U860 (N_860,In_1788,In_478);
nand U861 (N_861,In_843,In_148);
or U862 (N_862,In_1230,In_195);
or U863 (N_863,In_1117,In_1110);
nor U864 (N_864,In_1470,In_11);
and U865 (N_865,In_55,In_780);
nor U866 (N_866,In_941,In_683);
and U867 (N_867,In_276,In_552);
and U868 (N_868,In_1247,In_1352);
nor U869 (N_869,In_973,In_655);
xor U870 (N_870,In_719,In_606);
or U871 (N_871,In_1637,In_1782);
or U872 (N_872,In_1180,In_1005);
nand U873 (N_873,In_1130,In_1388);
nand U874 (N_874,In_1822,In_834);
or U875 (N_875,In_23,In_1508);
xor U876 (N_876,In_154,In_957);
nor U877 (N_877,In_1040,In_1902);
nand U878 (N_878,In_1159,In_301);
nand U879 (N_879,In_1248,In_1127);
xor U880 (N_880,In_667,In_1728);
and U881 (N_881,In_242,In_1253);
nand U882 (N_882,In_141,In_1490);
and U883 (N_883,In_1476,In_1859);
or U884 (N_884,In_1912,In_332);
and U885 (N_885,In_930,In_505);
and U886 (N_886,In_794,In_1800);
and U887 (N_887,In_1999,In_1337);
xnor U888 (N_888,In_1458,In_1278);
nor U889 (N_889,In_93,In_1934);
or U890 (N_890,In_632,In_1162);
xor U891 (N_891,In_1296,In_1923);
xnor U892 (N_892,In_1049,In_1872);
and U893 (N_893,In_213,In_566);
nor U894 (N_894,In_45,In_1334);
or U895 (N_895,In_922,In_1676);
or U896 (N_896,In_1361,In_1209);
nand U897 (N_897,In_1845,In_501);
nand U898 (N_898,In_1186,In_724);
or U899 (N_899,In_1739,In_1997);
nand U900 (N_900,In_812,In_1512);
nand U901 (N_901,In_350,In_917);
and U902 (N_902,In_1545,In_950);
nand U903 (N_903,In_1163,In_614);
and U904 (N_904,In_239,In_988);
nor U905 (N_905,In_806,In_732);
nor U906 (N_906,In_713,In_589);
and U907 (N_907,In_1964,In_1715);
nor U908 (N_908,In_1240,In_1687);
xor U909 (N_909,In_47,In_318);
nor U910 (N_910,In_1299,In_1454);
nor U911 (N_911,In_498,In_369);
xnor U912 (N_912,In_962,In_1260);
and U913 (N_913,In_1762,In_1208);
or U914 (N_914,In_1644,In_1153);
xor U915 (N_915,In_1916,In_1481);
or U916 (N_916,In_1484,In_475);
nand U917 (N_917,In_123,In_1391);
nand U918 (N_918,In_1084,In_1003);
xor U919 (N_919,In_1342,In_102);
or U920 (N_920,In_1671,In_1853);
and U921 (N_921,In_1483,In_848);
nor U922 (N_922,In_951,In_637);
nor U923 (N_923,In_1031,In_1704);
or U924 (N_924,In_567,In_836);
and U925 (N_925,In_1523,In_1951);
xor U926 (N_926,In_792,In_1666);
xnor U927 (N_927,In_151,In_1200);
nand U928 (N_928,In_1769,In_763);
xor U929 (N_929,In_1894,In_1237);
or U930 (N_930,In_583,In_511);
or U931 (N_931,In_1921,In_841);
nand U932 (N_932,In_1634,In_424);
nand U933 (N_933,In_1165,In_22);
nand U934 (N_934,In_676,In_303);
or U935 (N_935,In_1813,In_197);
nand U936 (N_936,In_1106,In_1668);
or U937 (N_937,In_287,In_1394);
and U938 (N_938,In_627,In_307);
and U939 (N_939,In_1821,In_416);
nor U940 (N_940,In_176,In_364);
nand U941 (N_941,In_1282,In_1598);
and U942 (N_942,In_274,In_1336);
nand U943 (N_943,In_961,In_1722);
xnor U944 (N_944,In_20,In_1711);
or U945 (N_945,In_1329,In_1109);
nand U946 (N_946,In_753,In_695);
and U947 (N_947,In_1358,In_230);
xnor U948 (N_948,In_244,In_1553);
or U949 (N_949,In_214,In_1023);
and U950 (N_950,In_135,In_454);
nor U951 (N_951,In_1992,In_1486);
and U952 (N_952,In_1572,In_1855);
nand U953 (N_953,In_1155,In_1978);
nor U954 (N_954,In_689,In_523);
nand U955 (N_955,In_660,In_277);
nor U956 (N_956,In_1423,In_441);
nor U957 (N_957,In_1541,In_1140);
or U958 (N_958,In_1957,In_1552);
nor U959 (N_959,In_1742,In_1217);
or U960 (N_960,In_1445,In_1532);
and U961 (N_961,In_591,In_488);
xor U962 (N_962,In_1459,In_293);
nand U963 (N_963,In_1881,In_1710);
or U964 (N_964,In_1510,In_1942);
nand U965 (N_965,In_1944,In_1856);
xnor U966 (N_966,In_152,In_1594);
and U967 (N_967,In_1435,In_508);
or U968 (N_968,In_1238,In_934);
nand U969 (N_969,In_1245,In_1669);
nor U970 (N_970,In_882,In_1280);
and U971 (N_971,In_1197,In_1860);
and U972 (N_972,In_1798,In_1638);
xnor U973 (N_973,In_341,In_182);
nand U974 (N_974,In_1191,In_1823);
or U975 (N_975,In_728,In_574);
and U976 (N_976,In_978,In_1596);
and U977 (N_977,In_1531,In_25);
and U978 (N_978,In_777,In_1889);
nand U979 (N_979,In_1920,In_439);
and U980 (N_980,In_1720,In_590);
and U981 (N_981,In_228,In_1343);
nor U982 (N_982,In_953,In_1446);
or U983 (N_983,In_756,In_1929);
nor U984 (N_984,In_1433,In_181);
and U985 (N_985,In_1451,In_886);
nand U986 (N_986,In_1287,In_238);
xor U987 (N_987,In_310,In_394);
xor U988 (N_988,In_1173,In_712);
xor U989 (N_989,In_1947,In_217);
nand U990 (N_990,In_10,In_1064);
nand U991 (N_991,In_855,In_1052);
or U992 (N_992,In_226,In_626);
nor U993 (N_993,In_71,In_172);
nor U994 (N_994,In_1630,In_227);
or U995 (N_995,In_108,In_1665);
and U996 (N_996,In_1290,In_126);
nand U997 (N_997,In_1104,In_1985);
or U998 (N_998,In_1702,In_635);
or U999 (N_999,In_1656,In_1825);
nand U1000 (N_1000,In_1951,In_911);
or U1001 (N_1001,In_710,In_1205);
nand U1002 (N_1002,In_1531,In_1920);
and U1003 (N_1003,In_476,In_1356);
or U1004 (N_1004,In_95,In_516);
or U1005 (N_1005,In_1551,In_560);
nand U1006 (N_1006,In_136,In_1688);
or U1007 (N_1007,In_678,In_1599);
and U1008 (N_1008,In_784,In_272);
xnor U1009 (N_1009,In_1676,In_1694);
or U1010 (N_1010,In_1085,In_1301);
xor U1011 (N_1011,In_53,In_914);
or U1012 (N_1012,In_432,In_582);
and U1013 (N_1013,In_899,In_1873);
or U1014 (N_1014,In_1422,In_811);
and U1015 (N_1015,In_1337,In_603);
nor U1016 (N_1016,In_1548,In_1715);
and U1017 (N_1017,In_647,In_677);
nand U1018 (N_1018,In_1422,In_1085);
or U1019 (N_1019,In_1708,In_564);
and U1020 (N_1020,In_1015,In_825);
nor U1021 (N_1021,In_149,In_1027);
and U1022 (N_1022,In_73,In_967);
nor U1023 (N_1023,In_520,In_317);
nor U1024 (N_1024,In_1217,In_659);
nor U1025 (N_1025,In_1313,In_709);
xor U1026 (N_1026,In_1464,In_422);
nand U1027 (N_1027,In_1814,In_780);
or U1028 (N_1028,In_637,In_1004);
nand U1029 (N_1029,In_1674,In_1071);
nor U1030 (N_1030,In_381,In_1396);
nor U1031 (N_1031,In_1967,In_1139);
nor U1032 (N_1032,In_1476,In_1761);
or U1033 (N_1033,In_590,In_1228);
nand U1034 (N_1034,In_1112,In_215);
nand U1035 (N_1035,In_1646,In_312);
and U1036 (N_1036,In_71,In_1577);
or U1037 (N_1037,In_578,In_1378);
or U1038 (N_1038,In_1132,In_1160);
and U1039 (N_1039,In_1059,In_928);
nor U1040 (N_1040,In_1678,In_696);
or U1041 (N_1041,In_773,In_1873);
nand U1042 (N_1042,In_648,In_1946);
xor U1043 (N_1043,In_1745,In_496);
nor U1044 (N_1044,In_831,In_99);
or U1045 (N_1045,In_10,In_1431);
and U1046 (N_1046,In_1768,In_295);
nor U1047 (N_1047,In_69,In_1945);
nor U1048 (N_1048,In_748,In_383);
nand U1049 (N_1049,In_301,In_1430);
nor U1050 (N_1050,In_1222,In_912);
or U1051 (N_1051,In_29,In_489);
or U1052 (N_1052,In_1248,In_1608);
nand U1053 (N_1053,In_326,In_680);
xnor U1054 (N_1054,In_1463,In_1754);
and U1055 (N_1055,In_868,In_951);
and U1056 (N_1056,In_380,In_1122);
nand U1057 (N_1057,In_588,In_1007);
nand U1058 (N_1058,In_1466,In_820);
nand U1059 (N_1059,In_129,In_1608);
or U1060 (N_1060,In_1182,In_1009);
nand U1061 (N_1061,In_1838,In_1845);
or U1062 (N_1062,In_1398,In_1328);
nor U1063 (N_1063,In_810,In_1900);
or U1064 (N_1064,In_831,In_539);
or U1065 (N_1065,In_1101,In_1036);
or U1066 (N_1066,In_1455,In_991);
nor U1067 (N_1067,In_1620,In_228);
or U1068 (N_1068,In_1483,In_161);
nor U1069 (N_1069,In_554,In_1821);
and U1070 (N_1070,In_1431,In_1246);
or U1071 (N_1071,In_1422,In_581);
nand U1072 (N_1072,In_154,In_431);
nor U1073 (N_1073,In_1019,In_1184);
nor U1074 (N_1074,In_1578,In_139);
or U1075 (N_1075,In_1891,In_1414);
and U1076 (N_1076,In_1153,In_1356);
and U1077 (N_1077,In_557,In_625);
nand U1078 (N_1078,In_1035,In_567);
nor U1079 (N_1079,In_1829,In_1463);
nand U1080 (N_1080,In_627,In_541);
and U1081 (N_1081,In_1921,In_724);
or U1082 (N_1082,In_1239,In_873);
or U1083 (N_1083,In_1284,In_440);
nand U1084 (N_1084,In_213,In_1340);
xnor U1085 (N_1085,In_64,In_1613);
or U1086 (N_1086,In_992,In_1713);
nand U1087 (N_1087,In_519,In_334);
nand U1088 (N_1088,In_1158,In_180);
and U1089 (N_1089,In_314,In_398);
nor U1090 (N_1090,In_1356,In_394);
nor U1091 (N_1091,In_1050,In_212);
and U1092 (N_1092,In_1866,In_1444);
or U1093 (N_1093,In_1538,In_53);
nand U1094 (N_1094,In_536,In_430);
and U1095 (N_1095,In_502,In_1994);
nand U1096 (N_1096,In_1041,In_1982);
nand U1097 (N_1097,In_1171,In_688);
nand U1098 (N_1098,In_411,In_1695);
nor U1099 (N_1099,In_1320,In_735);
nand U1100 (N_1100,In_1548,In_86);
and U1101 (N_1101,In_423,In_1960);
nand U1102 (N_1102,In_1880,In_1796);
nand U1103 (N_1103,In_1462,In_1754);
or U1104 (N_1104,In_1438,In_647);
nor U1105 (N_1105,In_1970,In_1520);
xor U1106 (N_1106,In_202,In_1577);
nand U1107 (N_1107,In_128,In_727);
nand U1108 (N_1108,In_1417,In_36);
xor U1109 (N_1109,In_100,In_185);
or U1110 (N_1110,In_1230,In_1183);
or U1111 (N_1111,In_701,In_1863);
and U1112 (N_1112,In_65,In_1488);
and U1113 (N_1113,In_496,In_1666);
xor U1114 (N_1114,In_269,In_696);
and U1115 (N_1115,In_1152,In_78);
nand U1116 (N_1116,In_801,In_486);
or U1117 (N_1117,In_260,In_1831);
nand U1118 (N_1118,In_1198,In_1041);
nor U1119 (N_1119,In_1340,In_158);
or U1120 (N_1120,In_69,In_725);
or U1121 (N_1121,In_1544,In_36);
nor U1122 (N_1122,In_1265,In_114);
nand U1123 (N_1123,In_1047,In_1725);
and U1124 (N_1124,In_1769,In_1617);
nand U1125 (N_1125,In_58,In_269);
nor U1126 (N_1126,In_1110,In_188);
nor U1127 (N_1127,In_796,In_1083);
and U1128 (N_1128,In_605,In_1807);
and U1129 (N_1129,In_586,In_1312);
or U1130 (N_1130,In_1912,In_343);
nor U1131 (N_1131,In_105,In_202);
nor U1132 (N_1132,In_1554,In_583);
and U1133 (N_1133,In_1458,In_493);
xnor U1134 (N_1134,In_508,In_1501);
nor U1135 (N_1135,In_55,In_1616);
and U1136 (N_1136,In_1066,In_1230);
nand U1137 (N_1137,In_197,In_478);
and U1138 (N_1138,In_1247,In_610);
and U1139 (N_1139,In_497,In_1829);
nand U1140 (N_1140,In_635,In_1160);
and U1141 (N_1141,In_799,In_1738);
or U1142 (N_1142,In_1489,In_1382);
xnor U1143 (N_1143,In_677,In_1323);
nor U1144 (N_1144,In_951,In_814);
nand U1145 (N_1145,In_588,In_110);
nand U1146 (N_1146,In_97,In_261);
nand U1147 (N_1147,In_925,In_1572);
nor U1148 (N_1148,In_815,In_293);
nor U1149 (N_1149,In_366,In_1487);
nor U1150 (N_1150,In_1015,In_1836);
or U1151 (N_1151,In_583,In_200);
xnor U1152 (N_1152,In_1787,In_480);
xnor U1153 (N_1153,In_1036,In_735);
or U1154 (N_1154,In_1864,In_247);
and U1155 (N_1155,In_1709,In_463);
and U1156 (N_1156,In_1386,In_910);
nand U1157 (N_1157,In_327,In_1901);
xnor U1158 (N_1158,In_935,In_1747);
xor U1159 (N_1159,In_401,In_327);
or U1160 (N_1160,In_3,In_499);
nand U1161 (N_1161,In_1618,In_1146);
and U1162 (N_1162,In_196,In_433);
or U1163 (N_1163,In_1006,In_517);
xor U1164 (N_1164,In_1025,In_885);
nor U1165 (N_1165,In_1173,In_1468);
and U1166 (N_1166,In_726,In_2);
or U1167 (N_1167,In_1468,In_1987);
xor U1168 (N_1168,In_1820,In_1437);
nand U1169 (N_1169,In_1434,In_261);
nand U1170 (N_1170,In_618,In_533);
xor U1171 (N_1171,In_360,In_1797);
nand U1172 (N_1172,In_1555,In_1880);
and U1173 (N_1173,In_622,In_1182);
or U1174 (N_1174,In_1351,In_1442);
and U1175 (N_1175,In_1964,In_580);
nand U1176 (N_1176,In_1455,In_193);
or U1177 (N_1177,In_82,In_1559);
and U1178 (N_1178,In_259,In_215);
nor U1179 (N_1179,In_517,In_1561);
nor U1180 (N_1180,In_1344,In_1363);
nand U1181 (N_1181,In_1162,In_1929);
or U1182 (N_1182,In_545,In_958);
nand U1183 (N_1183,In_37,In_1231);
nand U1184 (N_1184,In_1574,In_1084);
nand U1185 (N_1185,In_68,In_353);
nor U1186 (N_1186,In_558,In_1318);
and U1187 (N_1187,In_188,In_949);
or U1188 (N_1188,In_993,In_1630);
and U1189 (N_1189,In_224,In_983);
or U1190 (N_1190,In_876,In_186);
xor U1191 (N_1191,In_580,In_872);
nand U1192 (N_1192,In_1517,In_657);
xor U1193 (N_1193,In_1336,In_1444);
and U1194 (N_1194,In_1010,In_73);
nand U1195 (N_1195,In_133,In_4);
nor U1196 (N_1196,In_1968,In_208);
or U1197 (N_1197,In_925,In_138);
nor U1198 (N_1198,In_1340,In_403);
and U1199 (N_1199,In_1915,In_1351);
or U1200 (N_1200,In_1403,In_1063);
nor U1201 (N_1201,In_1657,In_298);
and U1202 (N_1202,In_523,In_1114);
or U1203 (N_1203,In_908,In_1074);
or U1204 (N_1204,In_457,In_192);
nor U1205 (N_1205,In_1283,In_435);
or U1206 (N_1206,In_1124,In_1857);
and U1207 (N_1207,In_1279,In_1147);
nor U1208 (N_1208,In_677,In_775);
and U1209 (N_1209,In_73,In_1074);
and U1210 (N_1210,In_278,In_221);
or U1211 (N_1211,In_1073,In_1653);
nand U1212 (N_1212,In_846,In_1567);
and U1213 (N_1213,In_785,In_1394);
nand U1214 (N_1214,In_577,In_472);
or U1215 (N_1215,In_620,In_809);
or U1216 (N_1216,In_956,In_1647);
nand U1217 (N_1217,In_1385,In_1574);
nor U1218 (N_1218,In_569,In_182);
or U1219 (N_1219,In_731,In_1257);
and U1220 (N_1220,In_814,In_298);
xnor U1221 (N_1221,In_522,In_1555);
or U1222 (N_1222,In_1034,In_326);
and U1223 (N_1223,In_1391,In_1981);
nor U1224 (N_1224,In_890,In_214);
nand U1225 (N_1225,In_448,In_1523);
nor U1226 (N_1226,In_1075,In_50);
or U1227 (N_1227,In_70,In_502);
or U1228 (N_1228,In_467,In_1569);
nand U1229 (N_1229,In_1243,In_1229);
and U1230 (N_1230,In_1354,In_512);
or U1231 (N_1231,In_1290,In_759);
nand U1232 (N_1232,In_1991,In_1596);
or U1233 (N_1233,In_1122,In_661);
nor U1234 (N_1234,In_1859,In_709);
nor U1235 (N_1235,In_1930,In_658);
nor U1236 (N_1236,In_206,In_610);
and U1237 (N_1237,In_1490,In_1741);
nand U1238 (N_1238,In_1023,In_1652);
and U1239 (N_1239,In_62,In_1441);
nand U1240 (N_1240,In_1778,In_990);
nand U1241 (N_1241,In_756,In_1187);
and U1242 (N_1242,In_773,In_227);
nor U1243 (N_1243,In_252,In_1833);
nor U1244 (N_1244,In_618,In_836);
nor U1245 (N_1245,In_287,In_1040);
nor U1246 (N_1246,In_1285,In_1216);
or U1247 (N_1247,In_228,In_1458);
or U1248 (N_1248,In_1467,In_1023);
nand U1249 (N_1249,In_1478,In_1801);
or U1250 (N_1250,In_1742,In_1896);
and U1251 (N_1251,In_1820,In_1343);
nor U1252 (N_1252,In_995,In_1769);
nor U1253 (N_1253,In_45,In_1694);
and U1254 (N_1254,In_316,In_290);
nand U1255 (N_1255,In_699,In_1601);
and U1256 (N_1256,In_593,In_1273);
or U1257 (N_1257,In_808,In_683);
or U1258 (N_1258,In_1385,In_341);
and U1259 (N_1259,In_92,In_1573);
nand U1260 (N_1260,In_407,In_1425);
and U1261 (N_1261,In_101,In_20);
or U1262 (N_1262,In_211,In_1693);
nand U1263 (N_1263,In_1389,In_153);
nor U1264 (N_1264,In_1276,In_1493);
nor U1265 (N_1265,In_816,In_1343);
nand U1266 (N_1266,In_1099,In_1706);
nand U1267 (N_1267,In_817,In_812);
and U1268 (N_1268,In_1106,In_1805);
nor U1269 (N_1269,In_28,In_1220);
nand U1270 (N_1270,In_789,In_1761);
nor U1271 (N_1271,In_793,In_1791);
nor U1272 (N_1272,In_483,In_369);
nor U1273 (N_1273,In_922,In_1635);
and U1274 (N_1274,In_1544,In_1660);
and U1275 (N_1275,In_1326,In_1761);
nand U1276 (N_1276,In_724,In_1247);
or U1277 (N_1277,In_941,In_1606);
xor U1278 (N_1278,In_935,In_956);
and U1279 (N_1279,In_782,In_525);
nand U1280 (N_1280,In_1970,In_1997);
and U1281 (N_1281,In_540,In_660);
nor U1282 (N_1282,In_1247,In_322);
xor U1283 (N_1283,In_1663,In_1225);
xor U1284 (N_1284,In_1201,In_1962);
and U1285 (N_1285,In_481,In_775);
nor U1286 (N_1286,In_164,In_45);
xor U1287 (N_1287,In_1859,In_658);
or U1288 (N_1288,In_1851,In_505);
or U1289 (N_1289,In_1601,In_967);
and U1290 (N_1290,In_1661,In_509);
and U1291 (N_1291,In_1551,In_1331);
nand U1292 (N_1292,In_310,In_1571);
xnor U1293 (N_1293,In_1212,In_232);
and U1294 (N_1294,In_544,In_902);
nand U1295 (N_1295,In_1156,In_281);
xor U1296 (N_1296,In_876,In_312);
nand U1297 (N_1297,In_455,In_1569);
or U1298 (N_1298,In_208,In_82);
and U1299 (N_1299,In_703,In_348);
and U1300 (N_1300,In_1960,In_818);
and U1301 (N_1301,In_749,In_1324);
or U1302 (N_1302,In_753,In_595);
nor U1303 (N_1303,In_1855,In_309);
or U1304 (N_1304,In_1626,In_730);
and U1305 (N_1305,In_1551,In_1752);
or U1306 (N_1306,In_1393,In_1683);
nand U1307 (N_1307,In_1708,In_1572);
or U1308 (N_1308,In_1056,In_1724);
or U1309 (N_1309,In_722,In_1219);
nor U1310 (N_1310,In_1510,In_1743);
and U1311 (N_1311,In_1929,In_1258);
nor U1312 (N_1312,In_473,In_171);
or U1313 (N_1313,In_1171,In_404);
xor U1314 (N_1314,In_421,In_840);
xor U1315 (N_1315,In_181,In_662);
nor U1316 (N_1316,In_1288,In_656);
and U1317 (N_1317,In_9,In_1662);
and U1318 (N_1318,In_275,In_1949);
and U1319 (N_1319,In_16,In_1237);
and U1320 (N_1320,In_221,In_1911);
nor U1321 (N_1321,In_29,In_1176);
nand U1322 (N_1322,In_1941,In_1704);
or U1323 (N_1323,In_948,In_168);
or U1324 (N_1324,In_851,In_958);
xnor U1325 (N_1325,In_1810,In_5);
nor U1326 (N_1326,In_505,In_1378);
and U1327 (N_1327,In_1768,In_1681);
xor U1328 (N_1328,In_52,In_1890);
nor U1329 (N_1329,In_1161,In_928);
or U1330 (N_1330,In_1969,In_491);
or U1331 (N_1331,In_1265,In_291);
and U1332 (N_1332,In_1516,In_1394);
xor U1333 (N_1333,In_1635,In_21);
or U1334 (N_1334,In_348,In_169);
nor U1335 (N_1335,In_1350,In_993);
nor U1336 (N_1336,In_648,In_1492);
nand U1337 (N_1337,In_1790,In_179);
and U1338 (N_1338,In_930,In_1784);
and U1339 (N_1339,In_1526,In_1951);
and U1340 (N_1340,In_335,In_1558);
and U1341 (N_1341,In_15,In_83);
or U1342 (N_1342,In_330,In_1326);
or U1343 (N_1343,In_1878,In_1231);
nor U1344 (N_1344,In_363,In_649);
nand U1345 (N_1345,In_950,In_602);
xnor U1346 (N_1346,In_1175,In_1083);
or U1347 (N_1347,In_1532,In_827);
nand U1348 (N_1348,In_785,In_937);
nand U1349 (N_1349,In_619,In_1691);
nand U1350 (N_1350,In_901,In_1345);
nand U1351 (N_1351,In_537,In_249);
and U1352 (N_1352,In_945,In_1865);
or U1353 (N_1353,In_432,In_1461);
nor U1354 (N_1354,In_475,In_825);
xnor U1355 (N_1355,In_804,In_698);
nor U1356 (N_1356,In_1384,In_1773);
or U1357 (N_1357,In_1989,In_1534);
xor U1358 (N_1358,In_1876,In_1511);
or U1359 (N_1359,In_339,In_114);
nand U1360 (N_1360,In_293,In_1657);
or U1361 (N_1361,In_1266,In_981);
xnor U1362 (N_1362,In_247,In_1576);
nand U1363 (N_1363,In_123,In_1365);
or U1364 (N_1364,In_254,In_123);
or U1365 (N_1365,In_812,In_191);
nor U1366 (N_1366,In_1156,In_172);
or U1367 (N_1367,In_968,In_1868);
nor U1368 (N_1368,In_1833,In_695);
or U1369 (N_1369,In_147,In_1831);
or U1370 (N_1370,In_1674,In_261);
nor U1371 (N_1371,In_197,In_417);
nand U1372 (N_1372,In_707,In_1568);
or U1373 (N_1373,In_1851,In_1123);
xor U1374 (N_1374,In_1168,In_184);
nand U1375 (N_1375,In_1281,In_1932);
and U1376 (N_1376,In_1747,In_1417);
nor U1377 (N_1377,In_669,In_1066);
nor U1378 (N_1378,In_1367,In_1717);
nand U1379 (N_1379,In_148,In_581);
or U1380 (N_1380,In_766,In_846);
or U1381 (N_1381,In_1403,In_1763);
or U1382 (N_1382,In_1368,In_464);
xnor U1383 (N_1383,In_1325,In_1863);
or U1384 (N_1384,In_926,In_1034);
nand U1385 (N_1385,In_715,In_1236);
nand U1386 (N_1386,In_866,In_670);
or U1387 (N_1387,In_1723,In_1391);
or U1388 (N_1388,In_1699,In_1613);
nand U1389 (N_1389,In_579,In_1771);
or U1390 (N_1390,In_633,In_1490);
and U1391 (N_1391,In_183,In_591);
and U1392 (N_1392,In_450,In_1222);
or U1393 (N_1393,In_1454,In_273);
and U1394 (N_1394,In_444,In_1158);
and U1395 (N_1395,In_44,In_747);
and U1396 (N_1396,In_730,In_848);
nand U1397 (N_1397,In_1282,In_1584);
nor U1398 (N_1398,In_1440,In_1489);
nor U1399 (N_1399,In_737,In_1201);
nor U1400 (N_1400,In_1384,In_920);
xor U1401 (N_1401,In_1516,In_1554);
nand U1402 (N_1402,In_715,In_1811);
or U1403 (N_1403,In_217,In_1469);
or U1404 (N_1404,In_748,In_1549);
nor U1405 (N_1405,In_1070,In_1360);
and U1406 (N_1406,In_1380,In_1889);
nand U1407 (N_1407,In_1507,In_1755);
and U1408 (N_1408,In_1514,In_1161);
or U1409 (N_1409,In_806,In_846);
and U1410 (N_1410,In_1799,In_1326);
xor U1411 (N_1411,In_662,In_341);
and U1412 (N_1412,In_1679,In_603);
and U1413 (N_1413,In_1733,In_1265);
nor U1414 (N_1414,In_647,In_978);
or U1415 (N_1415,In_808,In_1489);
nor U1416 (N_1416,In_984,In_1763);
and U1417 (N_1417,In_1578,In_915);
or U1418 (N_1418,In_517,In_1756);
and U1419 (N_1419,In_1770,In_1580);
nand U1420 (N_1420,In_903,In_367);
nand U1421 (N_1421,In_404,In_1170);
nand U1422 (N_1422,In_1329,In_372);
nor U1423 (N_1423,In_859,In_585);
and U1424 (N_1424,In_79,In_1404);
nor U1425 (N_1425,In_1224,In_163);
xor U1426 (N_1426,In_1240,In_1059);
nor U1427 (N_1427,In_169,In_952);
nand U1428 (N_1428,In_1072,In_1141);
and U1429 (N_1429,In_1284,In_981);
nand U1430 (N_1430,In_1506,In_446);
xnor U1431 (N_1431,In_1997,In_1062);
and U1432 (N_1432,In_269,In_1898);
or U1433 (N_1433,In_357,In_911);
xnor U1434 (N_1434,In_487,In_492);
or U1435 (N_1435,In_1405,In_1948);
nand U1436 (N_1436,In_985,In_407);
nor U1437 (N_1437,In_1292,In_672);
and U1438 (N_1438,In_814,In_1098);
or U1439 (N_1439,In_491,In_327);
or U1440 (N_1440,In_347,In_1360);
or U1441 (N_1441,In_225,In_1251);
nor U1442 (N_1442,In_199,In_1244);
and U1443 (N_1443,In_826,In_1590);
nand U1444 (N_1444,In_1603,In_1409);
and U1445 (N_1445,In_1730,In_1161);
xnor U1446 (N_1446,In_1593,In_1776);
or U1447 (N_1447,In_836,In_560);
and U1448 (N_1448,In_596,In_1804);
nor U1449 (N_1449,In_238,In_1027);
nand U1450 (N_1450,In_1701,In_1062);
and U1451 (N_1451,In_406,In_814);
and U1452 (N_1452,In_1107,In_1728);
nand U1453 (N_1453,In_1908,In_225);
and U1454 (N_1454,In_925,In_1613);
and U1455 (N_1455,In_1664,In_1200);
nor U1456 (N_1456,In_196,In_8);
and U1457 (N_1457,In_548,In_1339);
and U1458 (N_1458,In_1910,In_818);
nor U1459 (N_1459,In_1322,In_850);
and U1460 (N_1460,In_1256,In_639);
nor U1461 (N_1461,In_1501,In_525);
nor U1462 (N_1462,In_1241,In_1731);
nand U1463 (N_1463,In_524,In_1475);
nand U1464 (N_1464,In_598,In_614);
xnor U1465 (N_1465,In_1454,In_1322);
xor U1466 (N_1466,In_541,In_207);
nor U1467 (N_1467,In_808,In_1188);
nor U1468 (N_1468,In_296,In_40);
xnor U1469 (N_1469,In_1263,In_1710);
nand U1470 (N_1470,In_38,In_1562);
and U1471 (N_1471,In_923,In_1264);
xnor U1472 (N_1472,In_1485,In_1829);
nand U1473 (N_1473,In_960,In_1055);
or U1474 (N_1474,In_350,In_158);
nand U1475 (N_1475,In_671,In_1502);
and U1476 (N_1476,In_1973,In_1921);
xnor U1477 (N_1477,In_954,In_1866);
xor U1478 (N_1478,In_627,In_1147);
and U1479 (N_1479,In_1782,In_413);
xnor U1480 (N_1480,In_887,In_1198);
nand U1481 (N_1481,In_1806,In_1489);
nor U1482 (N_1482,In_205,In_1042);
nor U1483 (N_1483,In_315,In_1649);
nand U1484 (N_1484,In_551,In_560);
nor U1485 (N_1485,In_253,In_1155);
nand U1486 (N_1486,In_1368,In_715);
or U1487 (N_1487,In_219,In_396);
nand U1488 (N_1488,In_1911,In_565);
and U1489 (N_1489,In_1397,In_1477);
nor U1490 (N_1490,In_311,In_531);
or U1491 (N_1491,In_1523,In_153);
nor U1492 (N_1492,In_1795,In_786);
or U1493 (N_1493,In_1480,In_1278);
and U1494 (N_1494,In_1649,In_611);
and U1495 (N_1495,In_352,In_1206);
nand U1496 (N_1496,In_539,In_1030);
or U1497 (N_1497,In_830,In_466);
or U1498 (N_1498,In_1227,In_458);
and U1499 (N_1499,In_1515,In_1837);
nor U1500 (N_1500,In_1325,In_2);
and U1501 (N_1501,In_402,In_404);
xor U1502 (N_1502,In_98,In_1959);
or U1503 (N_1503,In_222,In_798);
nand U1504 (N_1504,In_130,In_24);
nand U1505 (N_1505,In_854,In_1619);
or U1506 (N_1506,In_151,In_1446);
nor U1507 (N_1507,In_666,In_519);
nor U1508 (N_1508,In_1383,In_1993);
and U1509 (N_1509,In_384,In_1974);
and U1510 (N_1510,In_1205,In_1271);
nor U1511 (N_1511,In_288,In_1182);
nor U1512 (N_1512,In_631,In_1154);
or U1513 (N_1513,In_1372,In_1428);
and U1514 (N_1514,In_1741,In_672);
nor U1515 (N_1515,In_1663,In_1097);
and U1516 (N_1516,In_39,In_401);
or U1517 (N_1517,In_1901,In_711);
and U1518 (N_1518,In_1935,In_1081);
nand U1519 (N_1519,In_1867,In_1173);
and U1520 (N_1520,In_348,In_796);
or U1521 (N_1521,In_1881,In_831);
nor U1522 (N_1522,In_1359,In_488);
nor U1523 (N_1523,In_166,In_1045);
or U1524 (N_1524,In_1612,In_336);
xor U1525 (N_1525,In_1177,In_643);
or U1526 (N_1526,In_1342,In_614);
xnor U1527 (N_1527,In_1301,In_1441);
nor U1528 (N_1528,In_1289,In_407);
nor U1529 (N_1529,In_1976,In_426);
and U1530 (N_1530,In_1227,In_1880);
or U1531 (N_1531,In_908,In_265);
and U1532 (N_1532,In_1482,In_1288);
nor U1533 (N_1533,In_930,In_758);
and U1534 (N_1534,In_1271,In_908);
nor U1535 (N_1535,In_957,In_1464);
or U1536 (N_1536,In_656,In_1715);
nand U1537 (N_1537,In_1214,In_1374);
nand U1538 (N_1538,In_472,In_526);
and U1539 (N_1539,In_1184,In_998);
xnor U1540 (N_1540,In_535,In_1105);
nor U1541 (N_1541,In_1453,In_871);
nand U1542 (N_1542,In_480,In_1972);
or U1543 (N_1543,In_1862,In_506);
nand U1544 (N_1544,In_1344,In_1891);
and U1545 (N_1545,In_897,In_1700);
nor U1546 (N_1546,In_606,In_766);
nand U1547 (N_1547,In_1136,In_1622);
and U1548 (N_1548,In_624,In_940);
nand U1549 (N_1549,In_506,In_270);
nand U1550 (N_1550,In_276,In_196);
nor U1551 (N_1551,In_844,In_1888);
and U1552 (N_1552,In_313,In_895);
and U1553 (N_1553,In_332,In_438);
and U1554 (N_1554,In_1636,In_1171);
xnor U1555 (N_1555,In_816,In_1947);
nand U1556 (N_1556,In_846,In_1378);
nor U1557 (N_1557,In_1920,In_1516);
and U1558 (N_1558,In_872,In_1844);
xnor U1559 (N_1559,In_1394,In_1785);
nand U1560 (N_1560,In_966,In_1027);
or U1561 (N_1561,In_1341,In_1101);
and U1562 (N_1562,In_142,In_1626);
or U1563 (N_1563,In_401,In_224);
nand U1564 (N_1564,In_518,In_532);
nor U1565 (N_1565,In_1579,In_205);
and U1566 (N_1566,In_48,In_1890);
nor U1567 (N_1567,In_1493,In_726);
nor U1568 (N_1568,In_495,In_1449);
nand U1569 (N_1569,In_326,In_882);
or U1570 (N_1570,In_329,In_1047);
and U1571 (N_1571,In_63,In_1244);
nand U1572 (N_1572,In_1323,In_1424);
or U1573 (N_1573,In_1307,In_120);
xnor U1574 (N_1574,In_1768,In_374);
or U1575 (N_1575,In_1932,In_1477);
or U1576 (N_1576,In_175,In_173);
and U1577 (N_1577,In_1344,In_1158);
and U1578 (N_1578,In_1554,In_808);
and U1579 (N_1579,In_1322,In_247);
and U1580 (N_1580,In_1458,In_551);
nor U1581 (N_1581,In_657,In_683);
and U1582 (N_1582,In_1043,In_931);
or U1583 (N_1583,In_1484,In_307);
nor U1584 (N_1584,In_1472,In_1326);
or U1585 (N_1585,In_1491,In_1033);
nor U1586 (N_1586,In_952,In_897);
and U1587 (N_1587,In_1638,In_227);
nand U1588 (N_1588,In_87,In_912);
nor U1589 (N_1589,In_1391,In_601);
xor U1590 (N_1590,In_1624,In_623);
or U1591 (N_1591,In_1155,In_288);
nand U1592 (N_1592,In_1985,In_1761);
or U1593 (N_1593,In_1725,In_1876);
or U1594 (N_1594,In_1577,In_781);
nand U1595 (N_1595,In_1401,In_1964);
and U1596 (N_1596,In_228,In_1755);
nand U1597 (N_1597,In_1685,In_1896);
and U1598 (N_1598,In_1752,In_1046);
nand U1599 (N_1599,In_501,In_891);
nor U1600 (N_1600,In_1782,In_955);
and U1601 (N_1601,In_64,In_423);
or U1602 (N_1602,In_1858,In_1528);
nor U1603 (N_1603,In_956,In_695);
nand U1604 (N_1604,In_882,In_1220);
nor U1605 (N_1605,In_1801,In_1002);
nand U1606 (N_1606,In_68,In_477);
nor U1607 (N_1607,In_1486,In_558);
nand U1608 (N_1608,In_975,In_111);
nand U1609 (N_1609,In_980,In_38);
nand U1610 (N_1610,In_814,In_1473);
nand U1611 (N_1611,In_24,In_1904);
nand U1612 (N_1612,In_1139,In_1405);
and U1613 (N_1613,In_412,In_16);
and U1614 (N_1614,In_1240,In_333);
xnor U1615 (N_1615,In_461,In_692);
or U1616 (N_1616,In_334,In_765);
nor U1617 (N_1617,In_6,In_1710);
nand U1618 (N_1618,In_1715,In_1132);
or U1619 (N_1619,In_1105,In_597);
or U1620 (N_1620,In_364,In_631);
nor U1621 (N_1621,In_1934,In_790);
nor U1622 (N_1622,In_452,In_410);
nand U1623 (N_1623,In_1933,In_1091);
nor U1624 (N_1624,In_622,In_1932);
nor U1625 (N_1625,In_1735,In_1820);
or U1626 (N_1626,In_860,In_379);
or U1627 (N_1627,In_1666,In_1621);
nor U1628 (N_1628,In_956,In_1989);
nand U1629 (N_1629,In_1962,In_448);
or U1630 (N_1630,In_1759,In_447);
and U1631 (N_1631,In_1480,In_1223);
nor U1632 (N_1632,In_872,In_993);
nand U1633 (N_1633,In_843,In_1307);
or U1634 (N_1634,In_644,In_945);
or U1635 (N_1635,In_1681,In_1645);
or U1636 (N_1636,In_115,In_1347);
or U1637 (N_1637,In_554,In_1660);
nor U1638 (N_1638,In_1567,In_926);
nand U1639 (N_1639,In_794,In_1912);
and U1640 (N_1640,In_503,In_1947);
nand U1641 (N_1641,In_55,In_1398);
or U1642 (N_1642,In_376,In_411);
nand U1643 (N_1643,In_1562,In_898);
and U1644 (N_1644,In_677,In_829);
nor U1645 (N_1645,In_1813,In_1996);
and U1646 (N_1646,In_1365,In_1633);
nor U1647 (N_1647,In_984,In_1985);
nor U1648 (N_1648,In_1087,In_297);
or U1649 (N_1649,In_1939,In_1560);
or U1650 (N_1650,In_719,In_100);
or U1651 (N_1651,In_27,In_1918);
or U1652 (N_1652,In_1123,In_630);
xor U1653 (N_1653,In_1028,In_1661);
and U1654 (N_1654,In_1868,In_1500);
nand U1655 (N_1655,In_699,In_1552);
nand U1656 (N_1656,In_160,In_1201);
nor U1657 (N_1657,In_1844,In_1153);
and U1658 (N_1658,In_1444,In_1177);
or U1659 (N_1659,In_826,In_1880);
nand U1660 (N_1660,In_1795,In_319);
or U1661 (N_1661,In_760,In_152);
or U1662 (N_1662,In_214,In_612);
or U1663 (N_1663,In_1778,In_1168);
and U1664 (N_1664,In_1803,In_436);
nor U1665 (N_1665,In_89,In_331);
and U1666 (N_1666,In_1433,In_120);
nor U1667 (N_1667,In_1642,In_1444);
nor U1668 (N_1668,In_1693,In_331);
and U1669 (N_1669,In_513,In_1512);
and U1670 (N_1670,In_1275,In_1254);
nand U1671 (N_1671,In_40,In_199);
nand U1672 (N_1672,In_192,In_1970);
or U1673 (N_1673,In_542,In_87);
or U1674 (N_1674,In_1784,In_1544);
and U1675 (N_1675,In_1835,In_1395);
nand U1676 (N_1676,In_698,In_1385);
nor U1677 (N_1677,In_1039,In_247);
xor U1678 (N_1678,In_921,In_1995);
xor U1679 (N_1679,In_1234,In_559);
xnor U1680 (N_1680,In_261,In_1312);
and U1681 (N_1681,In_1253,In_1999);
xnor U1682 (N_1682,In_1811,In_570);
or U1683 (N_1683,In_528,In_581);
nor U1684 (N_1684,In_1625,In_1963);
or U1685 (N_1685,In_252,In_1908);
xnor U1686 (N_1686,In_1545,In_1743);
nand U1687 (N_1687,In_1759,In_1468);
or U1688 (N_1688,In_1587,In_791);
nand U1689 (N_1689,In_499,In_348);
or U1690 (N_1690,In_438,In_874);
nand U1691 (N_1691,In_1775,In_517);
nor U1692 (N_1692,In_563,In_1296);
or U1693 (N_1693,In_738,In_514);
or U1694 (N_1694,In_1145,In_704);
nor U1695 (N_1695,In_1898,In_986);
nand U1696 (N_1696,In_1966,In_1434);
or U1697 (N_1697,In_1911,In_1558);
or U1698 (N_1698,In_409,In_1103);
nand U1699 (N_1699,In_1826,In_799);
nor U1700 (N_1700,In_1076,In_707);
xnor U1701 (N_1701,In_990,In_1917);
or U1702 (N_1702,In_719,In_995);
nand U1703 (N_1703,In_197,In_659);
nand U1704 (N_1704,In_1717,In_72);
nand U1705 (N_1705,In_540,In_1891);
xnor U1706 (N_1706,In_1838,In_1380);
and U1707 (N_1707,In_735,In_1027);
nand U1708 (N_1708,In_1339,In_1657);
or U1709 (N_1709,In_700,In_675);
or U1710 (N_1710,In_574,In_599);
xor U1711 (N_1711,In_1876,In_1430);
nor U1712 (N_1712,In_812,In_750);
and U1713 (N_1713,In_689,In_236);
or U1714 (N_1714,In_1881,In_1714);
xor U1715 (N_1715,In_1137,In_1581);
and U1716 (N_1716,In_1210,In_961);
nor U1717 (N_1717,In_375,In_749);
and U1718 (N_1718,In_1211,In_1715);
nand U1719 (N_1719,In_1631,In_1761);
or U1720 (N_1720,In_1009,In_1851);
xnor U1721 (N_1721,In_101,In_1224);
nand U1722 (N_1722,In_51,In_609);
and U1723 (N_1723,In_1008,In_618);
and U1724 (N_1724,In_621,In_656);
or U1725 (N_1725,In_572,In_864);
xor U1726 (N_1726,In_1457,In_1030);
nand U1727 (N_1727,In_4,In_1227);
or U1728 (N_1728,In_42,In_1771);
xnor U1729 (N_1729,In_162,In_1502);
and U1730 (N_1730,In_687,In_1524);
and U1731 (N_1731,In_1648,In_174);
nand U1732 (N_1732,In_1007,In_949);
and U1733 (N_1733,In_1146,In_1821);
or U1734 (N_1734,In_219,In_85);
nor U1735 (N_1735,In_610,In_929);
nor U1736 (N_1736,In_848,In_208);
nor U1737 (N_1737,In_1757,In_661);
nor U1738 (N_1738,In_1173,In_531);
nand U1739 (N_1739,In_680,In_705);
nand U1740 (N_1740,In_308,In_796);
nor U1741 (N_1741,In_1715,In_1277);
or U1742 (N_1742,In_1442,In_1846);
or U1743 (N_1743,In_355,In_102);
nand U1744 (N_1744,In_1688,In_1915);
or U1745 (N_1745,In_537,In_1368);
nand U1746 (N_1746,In_791,In_766);
nand U1747 (N_1747,In_1471,In_965);
and U1748 (N_1748,In_1705,In_818);
and U1749 (N_1749,In_1812,In_1503);
and U1750 (N_1750,In_376,In_1770);
and U1751 (N_1751,In_1061,In_976);
and U1752 (N_1752,In_187,In_1362);
xor U1753 (N_1753,In_1216,In_880);
nor U1754 (N_1754,In_452,In_166);
nand U1755 (N_1755,In_155,In_379);
or U1756 (N_1756,In_294,In_503);
and U1757 (N_1757,In_1945,In_177);
nand U1758 (N_1758,In_1947,In_1680);
and U1759 (N_1759,In_497,In_1912);
nand U1760 (N_1760,In_101,In_877);
or U1761 (N_1761,In_1241,In_1544);
nor U1762 (N_1762,In_1370,In_30);
nand U1763 (N_1763,In_254,In_690);
nor U1764 (N_1764,In_1327,In_1287);
xnor U1765 (N_1765,In_1988,In_1342);
and U1766 (N_1766,In_179,In_843);
and U1767 (N_1767,In_557,In_830);
or U1768 (N_1768,In_565,In_1963);
nor U1769 (N_1769,In_1145,In_1113);
nand U1770 (N_1770,In_134,In_962);
nor U1771 (N_1771,In_1635,In_1102);
xnor U1772 (N_1772,In_1753,In_485);
xnor U1773 (N_1773,In_1354,In_1861);
nor U1774 (N_1774,In_947,In_1518);
xor U1775 (N_1775,In_1931,In_1552);
and U1776 (N_1776,In_1009,In_431);
or U1777 (N_1777,In_1241,In_1176);
nand U1778 (N_1778,In_967,In_1126);
or U1779 (N_1779,In_1982,In_327);
xor U1780 (N_1780,In_726,In_1101);
or U1781 (N_1781,In_1121,In_1055);
nand U1782 (N_1782,In_448,In_1814);
or U1783 (N_1783,In_1791,In_1592);
and U1784 (N_1784,In_161,In_1590);
or U1785 (N_1785,In_1889,In_242);
or U1786 (N_1786,In_828,In_1855);
or U1787 (N_1787,In_1496,In_1113);
nand U1788 (N_1788,In_1914,In_1028);
and U1789 (N_1789,In_775,In_920);
and U1790 (N_1790,In_1778,In_1566);
nand U1791 (N_1791,In_988,In_529);
nand U1792 (N_1792,In_545,In_84);
nor U1793 (N_1793,In_763,In_1775);
or U1794 (N_1794,In_722,In_1285);
and U1795 (N_1795,In_504,In_88);
nand U1796 (N_1796,In_1349,In_903);
nand U1797 (N_1797,In_1172,In_103);
nand U1798 (N_1798,In_1073,In_189);
and U1799 (N_1799,In_1157,In_1160);
and U1800 (N_1800,In_1199,In_220);
and U1801 (N_1801,In_819,In_64);
nor U1802 (N_1802,In_1354,In_1013);
or U1803 (N_1803,In_745,In_793);
or U1804 (N_1804,In_1381,In_1830);
nor U1805 (N_1805,In_356,In_1024);
xor U1806 (N_1806,In_1623,In_486);
and U1807 (N_1807,In_1663,In_1291);
or U1808 (N_1808,In_1925,In_72);
or U1809 (N_1809,In_655,In_1932);
nor U1810 (N_1810,In_997,In_682);
or U1811 (N_1811,In_1915,In_1531);
or U1812 (N_1812,In_1331,In_1315);
nand U1813 (N_1813,In_1363,In_905);
or U1814 (N_1814,In_495,In_1063);
xor U1815 (N_1815,In_1306,In_1524);
xnor U1816 (N_1816,In_312,In_1835);
xnor U1817 (N_1817,In_1227,In_1899);
and U1818 (N_1818,In_13,In_765);
or U1819 (N_1819,In_1083,In_878);
nor U1820 (N_1820,In_1328,In_287);
or U1821 (N_1821,In_695,In_1251);
nor U1822 (N_1822,In_173,In_136);
xnor U1823 (N_1823,In_1267,In_454);
xnor U1824 (N_1824,In_190,In_1619);
and U1825 (N_1825,In_786,In_272);
nor U1826 (N_1826,In_877,In_1292);
or U1827 (N_1827,In_404,In_1599);
nand U1828 (N_1828,In_1309,In_1403);
nor U1829 (N_1829,In_313,In_512);
or U1830 (N_1830,In_1878,In_1578);
nand U1831 (N_1831,In_663,In_1205);
or U1832 (N_1832,In_1486,In_1974);
and U1833 (N_1833,In_1220,In_1473);
and U1834 (N_1834,In_558,In_1491);
nand U1835 (N_1835,In_1295,In_1822);
or U1836 (N_1836,In_91,In_822);
and U1837 (N_1837,In_1959,In_611);
nand U1838 (N_1838,In_861,In_232);
nor U1839 (N_1839,In_1319,In_635);
nand U1840 (N_1840,In_270,In_1758);
and U1841 (N_1841,In_1826,In_73);
nor U1842 (N_1842,In_443,In_1215);
or U1843 (N_1843,In_1153,In_791);
and U1844 (N_1844,In_1405,In_442);
nand U1845 (N_1845,In_723,In_1133);
and U1846 (N_1846,In_914,In_394);
nor U1847 (N_1847,In_1008,In_443);
and U1848 (N_1848,In_460,In_350);
and U1849 (N_1849,In_1637,In_1805);
nor U1850 (N_1850,In_1175,In_1068);
nand U1851 (N_1851,In_1614,In_429);
nand U1852 (N_1852,In_1806,In_553);
and U1853 (N_1853,In_120,In_329);
xnor U1854 (N_1854,In_462,In_85);
and U1855 (N_1855,In_439,In_724);
nor U1856 (N_1856,In_1581,In_1241);
or U1857 (N_1857,In_126,In_401);
xor U1858 (N_1858,In_1173,In_1687);
xnor U1859 (N_1859,In_1897,In_822);
nand U1860 (N_1860,In_799,In_589);
and U1861 (N_1861,In_1503,In_661);
xnor U1862 (N_1862,In_235,In_554);
nor U1863 (N_1863,In_1119,In_187);
nand U1864 (N_1864,In_411,In_1733);
and U1865 (N_1865,In_1383,In_1247);
nor U1866 (N_1866,In_1686,In_1614);
nor U1867 (N_1867,In_1101,In_44);
nand U1868 (N_1868,In_197,In_1264);
and U1869 (N_1869,In_1888,In_655);
and U1870 (N_1870,In_1994,In_1115);
nand U1871 (N_1871,In_1625,In_1323);
nor U1872 (N_1872,In_1011,In_747);
or U1873 (N_1873,In_1253,In_437);
nand U1874 (N_1874,In_140,In_812);
nor U1875 (N_1875,In_314,In_1008);
nor U1876 (N_1876,In_1289,In_1825);
and U1877 (N_1877,In_501,In_1549);
xor U1878 (N_1878,In_879,In_1371);
and U1879 (N_1879,In_1928,In_973);
or U1880 (N_1880,In_739,In_1756);
nand U1881 (N_1881,In_140,In_1516);
or U1882 (N_1882,In_718,In_1185);
or U1883 (N_1883,In_1824,In_253);
and U1884 (N_1884,In_1655,In_951);
and U1885 (N_1885,In_1883,In_81);
or U1886 (N_1886,In_1791,In_98);
or U1887 (N_1887,In_1735,In_898);
and U1888 (N_1888,In_390,In_1682);
nand U1889 (N_1889,In_972,In_1604);
and U1890 (N_1890,In_1204,In_724);
or U1891 (N_1891,In_199,In_1219);
and U1892 (N_1892,In_486,In_1649);
or U1893 (N_1893,In_1642,In_552);
and U1894 (N_1894,In_513,In_1958);
nand U1895 (N_1895,In_298,In_1193);
nand U1896 (N_1896,In_1135,In_1031);
or U1897 (N_1897,In_1157,In_1326);
nor U1898 (N_1898,In_605,In_503);
nand U1899 (N_1899,In_1567,In_57);
and U1900 (N_1900,In_225,In_1127);
and U1901 (N_1901,In_524,In_369);
nand U1902 (N_1902,In_1206,In_73);
or U1903 (N_1903,In_763,In_1111);
nand U1904 (N_1904,In_458,In_1310);
nand U1905 (N_1905,In_1128,In_1321);
xor U1906 (N_1906,In_1052,In_1210);
nor U1907 (N_1907,In_529,In_430);
and U1908 (N_1908,In_1899,In_1083);
nand U1909 (N_1909,In_37,In_381);
nor U1910 (N_1910,In_1742,In_1403);
and U1911 (N_1911,In_896,In_130);
or U1912 (N_1912,In_1339,In_30);
nor U1913 (N_1913,In_283,In_618);
nand U1914 (N_1914,In_1648,In_112);
nor U1915 (N_1915,In_1493,In_1850);
and U1916 (N_1916,In_0,In_1277);
nand U1917 (N_1917,In_1613,In_164);
nand U1918 (N_1918,In_365,In_1963);
and U1919 (N_1919,In_428,In_1041);
or U1920 (N_1920,In_525,In_1296);
or U1921 (N_1921,In_1616,In_984);
nand U1922 (N_1922,In_759,In_1157);
nand U1923 (N_1923,In_321,In_314);
nor U1924 (N_1924,In_285,In_1613);
nor U1925 (N_1925,In_1919,In_538);
and U1926 (N_1926,In_687,In_1491);
nand U1927 (N_1927,In_231,In_1255);
nand U1928 (N_1928,In_734,In_605);
or U1929 (N_1929,In_409,In_1225);
nor U1930 (N_1930,In_1158,In_1773);
or U1931 (N_1931,In_763,In_325);
and U1932 (N_1932,In_1859,In_1949);
or U1933 (N_1933,In_496,In_1973);
nor U1934 (N_1934,In_710,In_1235);
and U1935 (N_1935,In_1520,In_1698);
nand U1936 (N_1936,In_293,In_297);
nand U1937 (N_1937,In_144,In_781);
nor U1938 (N_1938,In_728,In_761);
nor U1939 (N_1939,In_1199,In_966);
xor U1940 (N_1940,In_603,In_1383);
xor U1941 (N_1941,In_906,In_370);
nor U1942 (N_1942,In_952,In_1394);
nand U1943 (N_1943,In_1047,In_528);
nand U1944 (N_1944,In_279,In_325);
nand U1945 (N_1945,In_1840,In_160);
or U1946 (N_1946,In_1235,In_1701);
nor U1947 (N_1947,In_1215,In_173);
nor U1948 (N_1948,In_464,In_774);
nand U1949 (N_1949,In_1480,In_884);
nor U1950 (N_1950,In_1611,In_1262);
or U1951 (N_1951,In_1469,In_677);
and U1952 (N_1952,In_824,In_1558);
xor U1953 (N_1953,In_1772,In_1572);
nand U1954 (N_1954,In_1635,In_1631);
xnor U1955 (N_1955,In_101,In_530);
nand U1956 (N_1956,In_1299,In_4);
nor U1957 (N_1957,In_1956,In_1990);
nand U1958 (N_1958,In_764,In_589);
nor U1959 (N_1959,In_1058,In_810);
xnor U1960 (N_1960,In_1017,In_1075);
and U1961 (N_1961,In_1978,In_900);
nor U1962 (N_1962,In_1776,In_186);
nand U1963 (N_1963,In_326,In_398);
nor U1964 (N_1964,In_742,In_1174);
or U1965 (N_1965,In_1636,In_1881);
or U1966 (N_1966,In_336,In_1054);
nand U1967 (N_1967,In_1076,In_1574);
nor U1968 (N_1968,In_1503,In_1102);
and U1969 (N_1969,In_501,In_832);
nand U1970 (N_1970,In_969,In_728);
nor U1971 (N_1971,In_120,In_1766);
or U1972 (N_1972,In_617,In_154);
nor U1973 (N_1973,In_922,In_1377);
nand U1974 (N_1974,In_165,In_1146);
or U1975 (N_1975,In_1578,In_1088);
nand U1976 (N_1976,In_224,In_1166);
nand U1977 (N_1977,In_1969,In_233);
xor U1978 (N_1978,In_1480,In_271);
and U1979 (N_1979,In_381,In_907);
nor U1980 (N_1980,In_469,In_1302);
and U1981 (N_1981,In_1172,In_1788);
nor U1982 (N_1982,In_1475,In_422);
xor U1983 (N_1983,In_1365,In_966);
nand U1984 (N_1984,In_740,In_1926);
or U1985 (N_1985,In_899,In_1141);
nand U1986 (N_1986,In_1209,In_1302);
nor U1987 (N_1987,In_1896,In_545);
nor U1988 (N_1988,In_630,In_49);
or U1989 (N_1989,In_483,In_950);
or U1990 (N_1990,In_351,In_687);
nor U1991 (N_1991,In_557,In_1086);
and U1992 (N_1992,In_998,In_1603);
and U1993 (N_1993,In_853,In_234);
xor U1994 (N_1994,In_157,In_1927);
nor U1995 (N_1995,In_201,In_969);
nor U1996 (N_1996,In_440,In_186);
or U1997 (N_1997,In_602,In_1561);
nand U1998 (N_1998,In_1315,In_168);
nand U1999 (N_1999,In_1704,In_1567);
and U2000 (N_2000,In_529,In_1842);
nor U2001 (N_2001,In_1643,In_375);
and U2002 (N_2002,In_514,In_1405);
xnor U2003 (N_2003,In_1185,In_431);
nor U2004 (N_2004,In_1680,In_1126);
or U2005 (N_2005,In_1802,In_1430);
and U2006 (N_2006,In_1411,In_1522);
nor U2007 (N_2007,In_9,In_1524);
and U2008 (N_2008,In_248,In_1042);
or U2009 (N_2009,In_33,In_388);
nor U2010 (N_2010,In_25,In_478);
nand U2011 (N_2011,In_194,In_665);
and U2012 (N_2012,In_908,In_856);
nor U2013 (N_2013,In_1125,In_80);
xnor U2014 (N_2014,In_917,In_95);
xor U2015 (N_2015,In_1253,In_578);
and U2016 (N_2016,In_1689,In_114);
nor U2017 (N_2017,In_1044,In_1154);
nor U2018 (N_2018,In_49,In_1114);
and U2019 (N_2019,In_1341,In_1592);
or U2020 (N_2020,In_1310,In_1502);
or U2021 (N_2021,In_623,In_795);
nand U2022 (N_2022,In_122,In_1748);
nor U2023 (N_2023,In_1283,In_1167);
and U2024 (N_2024,In_344,In_975);
and U2025 (N_2025,In_353,In_1802);
or U2026 (N_2026,In_1867,In_741);
nand U2027 (N_2027,In_1368,In_1071);
nor U2028 (N_2028,In_300,In_808);
and U2029 (N_2029,In_1564,In_244);
nor U2030 (N_2030,In_1074,In_567);
nor U2031 (N_2031,In_783,In_192);
xor U2032 (N_2032,In_220,In_1078);
nand U2033 (N_2033,In_1247,In_1052);
xor U2034 (N_2034,In_1621,In_1140);
xnor U2035 (N_2035,In_748,In_629);
or U2036 (N_2036,In_1012,In_1407);
nor U2037 (N_2037,In_1982,In_1507);
and U2038 (N_2038,In_530,In_1292);
xor U2039 (N_2039,In_82,In_216);
or U2040 (N_2040,In_542,In_1573);
and U2041 (N_2041,In_1060,In_423);
and U2042 (N_2042,In_172,In_608);
nor U2043 (N_2043,In_25,In_37);
nor U2044 (N_2044,In_1550,In_663);
nor U2045 (N_2045,In_320,In_1537);
xnor U2046 (N_2046,In_616,In_685);
nand U2047 (N_2047,In_1562,In_306);
nor U2048 (N_2048,In_535,In_1405);
and U2049 (N_2049,In_470,In_870);
and U2050 (N_2050,In_1706,In_1155);
nor U2051 (N_2051,In_971,In_660);
nor U2052 (N_2052,In_1905,In_1830);
and U2053 (N_2053,In_1898,In_1332);
nand U2054 (N_2054,In_981,In_877);
nand U2055 (N_2055,In_84,In_1893);
nor U2056 (N_2056,In_1012,In_1899);
xnor U2057 (N_2057,In_371,In_724);
nand U2058 (N_2058,In_132,In_3);
xnor U2059 (N_2059,In_48,In_830);
or U2060 (N_2060,In_1140,In_1334);
nand U2061 (N_2061,In_571,In_341);
nand U2062 (N_2062,In_1842,In_493);
nor U2063 (N_2063,In_1331,In_774);
or U2064 (N_2064,In_1337,In_1812);
and U2065 (N_2065,In_357,In_1312);
and U2066 (N_2066,In_218,In_1223);
nand U2067 (N_2067,In_321,In_1374);
or U2068 (N_2068,In_1886,In_437);
nor U2069 (N_2069,In_922,In_265);
or U2070 (N_2070,In_1842,In_1248);
and U2071 (N_2071,In_316,In_815);
or U2072 (N_2072,In_926,In_1520);
and U2073 (N_2073,In_577,In_121);
or U2074 (N_2074,In_720,In_32);
nor U2075 (N_2075,In_1774,In_938);
and U2076 (N_2076,In_879,In_1438);
and U2077 (N_2077,In_855,In_559);
nor U2078 (N_2078,In_1278,In_33);
and U2079 (N_2079,In_1169,In_488);
nand U2080 (N_2080,In_1868,In_458);
or U2081 (N_2081,In_1356,In_934);
xnor U2082 (N_2082,In_985,In_991);
nor U2083 (N_2083,In_1260,In_143);
and U2084 (N_2084,In_1475,In_188);
xor U2085 (N_2085,In_1394,In_772);
xnor U2086 (N_2086,In_1914,In_1670);
xnor U2087 (N_2087,In_1496,In_923);
and U2088 (N_2088,In_835,In_603);
nor U2089 (N_2089,In_1815,In_1509);
nor U2090 (N_2090,In_138,In_1652);
or U2091 (N_2091,In_1704,In_616);
xor U2092 (N_2092,In_1399,In_162);
nand U2093 (N_2093,In_1693,In_1420);
or U2094 (N_2094,In_276,In_270);
and U2095 (N_2095,In_1259,In_44);
and U2096 (N_2096,In_1134,In_1477);
nand U2097 (N_2097,In_475,In_1847);
and U2098 (N_2098,In_463,In_397);
and U2099 (N_2099,In_1171,In_1407);
xor U2100 (N_2100,In_1696,In_1990);
nor U2101 (N_2101,In_572,In_843);
and U2102 (N_2102,In_718,In_1602);
and U2103 (N_2103,In_118,In_374);
nand U2104 (N_2104,In_1913,In_1998);
nor U2105 (N_2105,In_1295,In_1097);
nand U2106 (N_2106,In_1702,In_99);
nor U2107 (N_2107,In_1874,In_1385);
and U2108 (N_2108,In_1323,In_575);
or U2109 (N_2109,In_1831,In_1713);
or U2110 (N_2110,In_568,In_1083);
xnor U2111 (N_2111,In_1100,In_1843);
or U2112 (N_2112,In_300,In_1971);
and U2113 (N_2113,In_1619,In_1915);
nor U2114 (N_2114,In_1510,In_1013);
or U2115 (N_2115,In_394,In_320);
nor U2116 (N_2116,In_39,In_527);
nand U2117 (N_2117,In_1250,In_1191);
or U2118 (N_2118,In_443,In_824);
nor U2119 (N_2119,In_1681,In_1043);
nand U2120 (N_2120,In_1118,In_515);
or U2121 (N_2121,In_1787,In_704);
or U2122 (N_2122,In_1106,In_1038);
nor U2123 (N_2123,In_291,In_438);
nor U2124 (N_2124,In_1451,In_727);
and U2125 (N_2125,In_605,In_1922);
nand U2126 (N_2126,In_1340,In_1146);
and U2127 (N_2127,In_1536,In_1166);
nand U2128 (N_2128,In_247,In_198);
nand U2129 (N_2129,In_566,In_456);
or U2130 (N_2130,In_628,In_1594);
nor U2131 (N_2131,In_658,In_1839);
and U2132 (N_2132,In_58,In_1974);
or U2133 (N_2133,In_1734,In_1332);
nand U2134 (N_2134,In_411,In_1772);
nand U2135 (N_2135,In_757,In_645);
nand U2136 (N_2136,In_1874,In_277);
nand U2137 (N_2137,In_531,In_1938);
nand U2138 (N_2138,In_526,In_1019);
or U2139 (N_2139,In_1540,In_1501);
or U2140 (N_2140,In_1330,In_1818);
and U2141 (N_2141,In_1496,In_944);
nand U2142 (N_2142,In_1815,In_683);
nor U2143 (N_2143,In_1719,In_1934);
or U2144 (N_2144,In_1191,In_1545);
or U2145 (N_2145,In_1412,In_1000);
nand U2146 (N_2146,In_1991,In_1119);
nor U2147 (N_2147,In_1347,In_387);
nand U2148 (N_2148,In_1870,In_1294);
nand U2149 (N_2149,In_931,In_347);
nor U2150 (N_2150,In_13,In_1483);
nand U2151 (N_2151,In_897,In_308);
and U2152 (N_2152,In_1289,In_559);
nor U2153 (N_2153,In_1911,In_1618);
or U2154 (N_2154,In_637,In_1905);
or U2155 (N_2155,In_1450,In_1725);
and U2156 (N_2156,In_28,In_779);
nor U2157 (N_2157,In_1445,In_905);
and U2158 (N_2158,In_843,In_1356);
and U2159 (N_2159,In_73,In_1436);
xnor U2160 (N_2160,In_226,In_1260);
or U2161 (N_2161,In_969,In_605);
nor U2162 (N_2162,In_817,In_1627);
xnor U2163 (N_2163,In_177,In_1850);
nor U2164 (N_2164,In_1355,In_819);
nand U2165 (N_2165,In_832,In_175);
or U2166 (N_2166,In_358,In_1195);
or U2167 (N_2167,In_416,In_1987);
and U2168 (N_2168,In_83,In_1555);
nor U2169 (N_2169,In_962,In_600);
nand U2170 (N_2170,In_106,In_1247);
or U2171 (N_2171,In_1487,In_1730);
nor U2172 (N_2172,In_767,In_567);
nor U2173 (N_2173,In_1367,In_1573);
nor U2174 (N_2174,In_1448,In_745);
and U2175 (N_2175,In_1254,In_177);
nor U2176 (N_2176,In_1623,In_711);
nor U2177 (N_2177,In_566,In_1379);
nand U2178 (N_2178,In_1677,In_1028);
and U2179 (N_2179,In_1566,In_1997);
nand U2180 (N_2180,In_143,In_196);
xnor U2181 (N_2181,In_817,In_927);
xor U2182 (N_2182,In_338,In_1553);
and U2183 (N_2183,In_1374,In_186);
nor U2184 (N_2184,In_1841,In_1975);
nand U2185 (N_2185,In_200,In_1521);
or U2186 (N_2186,In_637,In_88);
nor U2187 (N_2187,In_1491,In_1090);
or U2188 (N_2188,In_360,In_842);
nand U2189 (N_2189,In_1501,In_1767);
nand U2190 (N_2190,In_338,In_1745);
or U2191 (N_2191,In_1275,In_394);
or U2192 (N_2192,In_828,In_1892);
and U2193 (N_2193,In_835,In_880);
or U2194 (N_2194,In_1614,In_114);
nand U2195 (N_2195,In_904,In_1848);
or U2196 (N_2196,In_1237,In_1908);
nand U2197 (N_2197,In_1837,In_1907);
nor U2198 (N_2198,In_1905,In_1759);
and U2199 (N_2199,In_465,In_1649);
or U2200 (N_2200,In_1868,In_109);
or U2201 (N_2201,In_729,In_199);
and U2202 (N_2202,In_308,In_142);
and U2203 (N_2203,In_893,In_653);
nand U2204 (N_2204,In_1238,In_1270);
and U2205 (N_2205,In_1953,In_552);
and U2206 (N_2206,In_1385,In_1030);
and U2207 (N_2207,In_705,In_662);
nand U2208 (N_2208,In_1822,In_1593);
nand U2209 (N_2209,In_74,In_892);
xnor U2210 (N_2210,In_984,In_1578);
xor U2211 (N_2211,In_968,In_505);
xnor U2212 (N_2212,In_51,In_1456);
or U2213 (N_2213,In_1143,In_203);
xor U2214 (N_2214,In_1661,In_868);
nor U2215 (N_2215,In_872,In_1874);
nand U2216 (N_2216,In_217,In_790);
or U2217 (N_2217,In_1206,In_883);
nand U2218 (N_2218,In_178,In_425);
and U2219 (N_2219,In_1177,In_599);
xor U2220 (N_2220,In_1206,In_248);
or U2221 (N_2221,In_1309,In_1036);
or U2222 (N_2222,In_736,In_437);
and U2223 (N_2223,In_622,In_318);
and U2224 (N_2224,In_1817,In_1305);
nand U2225 (N_2225,In_1892,In_1319);
xnor U2226 (N_2226,In_35,In_1875);
xnor U2227 (N_2227,In_1799,In_1389);
nor U2228 (N_2228,In_77,In_1979);
nor U2229 (N_2229,In_803,In_974);
nand U2230 (N_2230,In_893,In_1196);
or U2231 (N_2231,In_1297,In_970);
nand U2232 (N_2232,In_1771,In_75);
nand U2233 (N_2233,In_266,In_1951);
nand U2234 (N_2234,In_886,In_1676);
or U2235 (N_2235,In_182,In_1249);
or U2236 (N_2236,In_706,In_904);
and U2237 (N_2237,In_176,In_726);
and U2238 (N_2238,In_246,In_1574);
nor U2239 (N_2239,In_1734,In_446);
nand U2240 (N_2240,In_1734,In_555);
nor U2241 (N_2241,In_1349,In_220);
or U2242 (N_2242,In_1947,In_1587);
nor U2243 (N_2243,In_1966,In_168);
nand U2244 (N_2244,In_546,In_441);
and U2245 (N_2245,In_50,In_789);
and U2246 (N_2246,In_681,In_702);
nor U2247 (N_2247,In_921,In_1369);
or U2248 (N_2248,In_1214,In_390);
and U2249 (N_2249,In_1369,In_1881);
or U2250 (N_2250,In_188,In_1219);
nand U2251 (N_2251,In_839,In_1174);
or U2252 (N_2252,In_898,In_1803);
nor U2253 (N_2253,In_619,In_1391);
xnor U2254 (N_2254,In_897,In_456);
and U2255 (N_2255,In_1872,In_679);
nor U2256 (N_2256,In_1402,In_1842);
nand U2257 (N_2257,In_1430,In_1425);
nor U2258 (N_2258,In_579,In_153);
or U2259 (N_2259,In_816,In_1936);
nand U2260 (N_2260,In_1606,In_142);
and U2261 (N_2261,In_482,In_979);
and U2262 (N_2262,In_1548,In_1347);
and U2263 (N_2263,In_624,In_1725);
nor U2264 (N_2264,In_1236,In_349);
or U2265 (N_2265,In_516,In_1973);
nand U2266 (N_2266,In_1839,In_1046);
or U2267 (N_2267,In_830,In_1954);
or U2268 (N_2268,In_466,In_478);
or U2269 (N_2269,In_587,In_24);
nand U2270 (N_2270,In_1613,In_1738);
and U2271 (N_2271,In_531,In_1645);
and U2272 (N_2272,In_791,In_1842);
or U2273 (N_2273,In_1634,In_1728);
xor U2274 (N_2274,In_1556,In_1367);
or U2275 (N_2275,In_625,In_429);
nand U2276 (N_2276,In_404,In_1575);
and U2277 (N_2277,In_222,In_446);
or U2278 (N_2278,In_1719,In_1646);
or U2279 (N_2279,In_1305,In_1496);
nand U2280 (N_2280,In_1618,In_209);
or U2281 (N_2281,In_857,In_1905);
nand U2282 (N_2282,In_448,In_1283);
or U2283 (N_2283,In_1965,In_1878);
nand U2284 (N_2284,In_548,In_1509);
and U2285 (N_2285,In_850,In_1357);
and U2286 (N_2286,In_702,In_1050);
nand U2287 (N_2287,In_1634,In_111);
nor U2288 (N_2288,In_87,In_860);
and U2289 (N_2289,In_970,In_202);
nor U2290 (N_2290,In_706,In_852);
nor U2291 (N_2291,In_1916,In_1878);
nor U2292 (N_2292,In_1898,In_1501);
nand U2293 (N_2293,In_437,In_1311);
or U2294 (N_2294,In_283,In_29);
nand U2295 (N_2295,In_1312,In_1280);
nor U2296 (N_2296,In_1862,In_847);
nand U2297 (N_2297,In_105,In_285);
or U2298 (N_2298,In_1784,In_996);
and U2299 (N_2299,In_358,In_1961);
or U2300 (N_2300,In_1999,In_625);
nor U2301 (N_2301,In_772,In_1629);
and U2302 (N_2302,In_470,In_1692);
nor U2303 (N_2303,In_1760,In_483);
or U2304 (N_2304,In_791,In_1276);
xor U2305 (N_2305,In_408,In_483);
or U2306 (N_2306,In_371,In_1548);
or U2307 (N_2307,In_104,In_619);
nand U2308 (N_2308,In_721,In_40);
xor U2309 (N_2309,In_823,In_1138);
or U2310 (N_2310,In_1891,In_518);
or U2311 (N_2311,In_2,In_681);
and U2312 (N_2312,In_1548,In_466);
nand U2313 (N_2313,In_202,In_1671);
nor U2314 (N_2314,In_1158,In_14);
and U2315 (N_2315,In_1114,In_952);
and U2316 (N_2316,In_456,In_443);
or U2317 (N_2317,In_1156,In_1634);
or U2318 (N_2318,In_369,In_167);
or U2319 (N_2319,In_972,In_866);
nand U2320 (N_2320,In_1463,In_1814);
xor U2321 (N_2321,In_137,In_1985);
and U2322 (N_2322,In_1116,In_1714);
and U2323 (N_2323,In_414,In_1816);
or U2324 (N_2324,In_616,In_571);
or U2325 (N_2325,In_875,In_1201);
nor U2326 (N_2326,In_106,In_1439);
and U2327 (N_2327,In_615,In_1839);
and U2328 (N_2328,In_576,In_1422);
xnor U2329 (N_2329,In_774,In_852);
nand U2330 (N_2330,In_1035,In_202);
and U2331 (N_2331,In_1270,In_1781);
and U2332 (N_2332,In_568,In_617);
nor U2333 (N_2333,In_18,In_1430);
nor U2334 (N_2334,In_244,In_1431);
xnor U2335 (N_2335,In_802,In_1279);
xor U2336 (N_2336,In_1626,In_593);
nand U2337 (N_2337,In_77,In_1010);
nor U2338 (N_2338,In_715,In_473);
and U2339 (N_2339,In_930,In_291);
nand U2340 (N_2340,In_1432,In_1826);
nand U2341 (N_2341,In_1159,In_170);
or U2342 (N_2342,In_497,In_1694);
nand U2343 (N_2343,In_688,In_1882);
nand U2344 (N_2344,In_1121,In_1782);
xor U2345 (N_2345,In_444,In_840);
nand U2346 (N_2346,In_1470,In_1604);
xor U2347 (N_2347,In_1853,In_133);
nand U2348 (N_2348,In_1877,In_1498);
and U2349 (N_2349,In_1129,In_1092);
nand U2350 (N_2350,In_76,In_1896);
or U2351 (N_2351,In_1386,In_151);
nor U2352 (N_2352,In_430,In_1521);
nand U2353 (N_2353,In_243,In_1386);
nor U2354 (N_2354,In_404,In_1788);
nand U2355 (N_2355,In_499,In_908);
nor U2356 (N_2356,In_917,In_861);
nor U2357 (N_2357,In_1434,In_1609);
and U2358 (N_2358,In_1922,In_382);
nor U2359 (N_2359,In_1675,In_730);
and U2360 (N_2360,In_1825,In_621);
nor U2361 (N_2361,In_1021,In_1031);
and U2362 (N_2362,In_1743,In_234);
or U2363 (N_2363,In_764,In_1727);
or U2364 (N_2364,In_667,In_850);
nand U2365 (N_2365,In_1493,In_1331);
or U2366 (N_2366,In_753,In_1775);
and U2367 (N_2367,In_1537,In_1240);
and U2368 (N_2368,In_1193,In_1116);
or U2369 (N_2369,In_1481,In_1680);
nand U2370 (N_2370,In_140,In_1502);
nor U2371 (N_2371,In_905,In_281);
nand U2372 (N_2372,In_863,In_184);
nand U2373 (N_2373,In_1721,In_1439);
or U2374 (N_2374,In_1810,In_845);
xnor U2375 (N_2375,In_1148,In_54);
and U2376 (N_2376,In_1313,In_108);
and U2377 (N_2377,In_1875,In_1648);
nand U2378 (N_2378,In_394,In_1568);
nor U2379 (N_2379,In_182,In_1446);
nor U2380 (N_2380,In_1706,In_955);
or U2381 (N_2381,In_796,In_1015);
nand U2382 (N_2382,In_246,In_781);
and U2383 (N_2383,In_293,In_61);
nor U2384 (N_2384,In_1661,In_631);
or U2385 (N_2385,In_1545,In_1313);
and U2386 (N_2386,In_0,In_999);
and U2387 (N_2387,In_805,In_471);
nor U2388 (N_2388,In_1688,In_1741);
nand U2389 (N_2389,In_1334,In_217);
or U2390 (N_2390,In_925,In_796);
or U2391 (N_2391,In_130,In_908);
nor U2392 (N_2392,In_826,In_1017);
nor U2393 (N_2393,In_836,In_661);
nand U2394 (N_2394,In_1277,In_281);
xor U2395 (N_2395,In_1191,In_1764);
or U2396 (N_2396,In_917,In_1522);
or U2397 (N_2397,In_757,In_932);
and U2398 (N_2398,In_789,In_1782);
nand U2399 (N_2399,In_1978,In_288);
xnor U2400 (N_2400,In_868,In_420);
xor U2401 (N_2401,In_234,In_113);
or U2402 (N_2402,In_596,In_634);
nand U2403 (N_2403,In_604,In_1556);
or U2404 (N_2404,In_852,In_509);
or U2405 (N_2405,In_1700,In_18);
nand U2406 (N_2406,In_1527,In_731);
and U2407 (N_2407,In_91,In_753);
nand U2408 (N_2408,In_1948,In_491);
or U2409 (N_2409,In_613,In_211);
xor U2410 (N_2410,In_1445,In_1303);
and U2411 (N_2411,In_910,In_1485);
nor U2412 (N_2412,In_1496,In_20);
nor U2413 (N_2413,In_1158,In_1715);
nor U2414 (N_2414,In_1666,In_103);
nor U2415 (N_2415,In_1487,In_1124);
nand U2416 (N_2416,In_1913,In_89);
nor U2417 (N_2417,In_737,In_1512);
nand U2418 (N_2418,In_1952,In_1178);
nand U2419 (N_2419,In_8,In_1710);
and U2420 (N_2420,In_644,In_1998);
and U2421 (N_2421,In_1411,In_651);
and U2422 (N_2422,In_486,In_563);
nor U2423 (N_2423,In_1286,In_219);
or U2424 (N_2424,In_689,In_943);
and U2425 (N_2425,In_530,In_1040);
nor U2426 (N_2426,In_1358,In_275);
nor U2427 (N_2427,In_1593,In_1264);
and U2428 (N_2428,In_1564,In_425);
and U2429 (N_2429,In_679,In_643);
xnor U2430 (N_2430,In_757,In_1720);
or U2431 (N_2431,In_609,In_688);
and U2432 (N_2432,In_101,In_1036);
nor U2433 (N_2433,In_1838,In_1963);
xor U2434 (N_2434,In_1053,In_1716);
nand U2435 (N_2435,In_158,In_864);
and U2436 (N_2436,In_1684,In_272);
xnor U2437 (N_2437,In_152,In_1316);
nor U2438 (N_2438,In_1723,In_290);
and U2439 (N_2439,In_336,In_688);
and U2440 (N_2440,In_345,In_1820);
nor U2441 (N_2441,In_1526,In_999);
nor U2442 (N_2442,In_1605,In_1483);
nand U2443 (N_2443,In_184,In_871);
nor U2444 (N_2444,In_1787,In_1712);
or U2445 (N_2445,In_577,In_1171);
or U2446 (N_2446,In_1895,In_150);
xnor U2447 (N_2447,In_584,In_1055);
and U2448 (N_2448,In_756,In_167);
and U2449 (N_2449,In_1054,In_683);
nor U2450 (N_2450,In_538,In_1567);
nor U2451 (N_2451,In_1865,In_1568);
nor U2452 (N_2452,In_542,In_367);
xnor U2453 (N_2453,In_1931,In_1430);
or U2454 (N_2454,In_1439,In_357);
and U2455 (N_2455,In_1775,In_1465);
or U2456 (N_2456,In_337,In_729);
nor U2457 (N_2457,In_567,In_1732);
nand U2458 (N_2458,In_206,In_721);
nand U2459 (N_2459,In_1758,In_1795);
or U2460 (N_2460,In_22,In_903);
nand U2461 (N_2461,In_701,In_129);
nand U2462 (N_2462,In_173,In_1113);
or U2463 (N_2463,In_701,In_1300);
nand U2464 (N_2464,In_870,In_979);
or U2465 (N_2465,In_705,In_1954);
nor U2466 (N_2466,In_1430,In_1831);
nor U2467 (N_2467,In_300,In_388);
nand U2468 (N_2468,In_1320,In_1619);
xor U2469 (N_2469,In_874,In_735);
nand U2470 (N_2470,In_353,In_1824);
and U2471 (N_2471,In_1949,In_825);
nand U2472 (N_2472,In_1466,In_1947);
nand U2473 (N_2473,In_1724,In_1087);
and U2474 (N_2474,In_1732,In_252);
xnor U2475 (N_2475,In_1546,In_945);
nor U2476 (N_2476,In_1251,In_474);
and U2477 (N_2477,In_1467,In_1883);
nand U2478 (N_2478,In_170,In_1966);
and U2479 (N_2479,In_308,In_1950);
nand U2480 (N_2480,In_1614,In_1870);
nand U2481 (N_2481,In_466,In_1555);
or U2482 (N_2482,In_1777,In_574);
and U2483 (N_2483,In_281,In_1796);
and U2484 (N_2484,In_1064,In_1718);
nand U2485 (N_2485,In_1188,In_795);
nor U2486 (N_2486,In_1506,In_726);
nor U2487 (N_2487,In_1227,In_964);
and U2488 (N_2488,In_376,In_1378);
nor U2489 (N_2489,In_1751,In_975);
or U2490 (N_2490,In_1480,In_1358);
nor U2491 (N_2491,In_193,In_442);
and U2492 (N_2492,In_1322,In_1354);
or U2493 (N_2493,In_426,In_1155);
and U2494 (N_2494,In_1696,In_150);
nor U2495 (N_2495,In_814,In_496);
xor U2496 (N_2496,In_796,In_1534);
nor U2497 (N_2497,In_670,In_1318);
or U2498 (N_2498,In_1279,In_1937);
nor U2499 (N_2499,In_1291,In_1235);
nor U2500 (N_2500,In_1910,In_174);
and U2501 (N_2501,In_694,In_1620);
nand U2502 (N_2502,In_390,In_1684);
nor U2503 (N_2503,In_878,In_868);
and U2504 (N_2504,In_1997,In_738);
and U2505 (N_2505,In_1372,In_898);
and U2506 (N_2506,In_1138,In_403);
xnor U2507 (N_2507,In_879,In_6);
and U2508 (N_2508,In_248,In_282);
xnor U2509 (N_2509,In_732,In_356);
nand U2510 (N_2510,In_227,In_889);
or U2511 (N_2511,In_1922,In_289);
nor U2512 (N_2512,In_478,In_347);
xor U2513 (N_2513,In_1115,In_1711);
or U2514 (N_2514,In_1192,In_391);
nor U2515 (N_2515,In_368,In_1076);
xnor U2516 (N_2516,In_259,In_1590);
xor U2517 (N_2517,In_1617,In_24);
and U2518 (N_2518,In_1814,In_565);
and U2519 (N_2519,In_1595,In_588);
nand U2520 (N_2520,In_34,In_1025);
or U2521 (N_2521,In_1079,In_1966);
xor U2522 (N_2522,In_460,In_666);
nand U2523 (N_2523,In_1915,In_1121);
xnor U2524 (N_2524,In_669,In_777);
nor U2525 (N_2525,In_353,In_1598);
nand U2526 (N_2526,In_1872,In_1326);
nor U2527 (N_2527,In_1823,In_1211);
nor U2528 (N_2528,In_649,In_834);
nand U2529 (N_2529,In_1872,In_1114);
nor U2530 (N_2530,In_562,In_418);
nor U2531 (N_2531,In_573,In_133);
nor U2532 (N_2532,In_468,In_1096);
nand U2533 (N_2533,In_1329,In_1172);
nand U2534 (N_2534,In_666,In_269);
xnor U2535 (N_2535,In_478,In_1671);
or U2536 (N_2536,In_1154,In_709);
nor U2537 (N_2537,In_1501,In_1555);
and U2538 (N_2538,In_266,In_1635);
and U2539 (N_2539,In_1299,In_1040);
xnor U2540 (N_2540,In_1029,In_287);
and U2541 (N_2541,In_1666,In_1377);
or U2542 (N_2542,In_450,In_569);
nand U2543 (N_2543,In_1323,In_1109);
nand U2544 (N_2544,In_280,In_1644);
nand U2545 (N_2545,In_91,In_1751);
or U2546 (N_2546,In_1283,In_728);
or U2547 (N_2547,In_737,In_1473);
nand U2548 (N_2548,In_1964,In_122);
or U2549 (N_2549,In_1042,In_605);
nand U2550 (N_2550,In_131,In_973);
nand U2551 (N_2551,In_1451,In_1538);
or U2552 (N_2552,In_579,In_1811);
or U2553 (N_2553,In_1655,In_1492);
nor U2554 (N_2554,In_489,In_1089);
and U2555 (N_2555,In_1650,In_120);
nor U2556 (N_2556,In_1460,In_769);
xor U2557 (N_2557,In_256,In_221);
xor U2558 (N_2558,In_1380,In_303);
and U2559 (N_2559,In_1647,In_700);
xnor U2560 (N_2560,In_347,In_979);
or U2561 (N_2561,In_1617,In_1459);
or U2562 (N_2562,In_1104,In_980);
nor U2563 (N_2563,In_1760,In_568);
nand U2564 (N_2564,In_1684,In_578);
or U2565 (N_2565,In_1514,In_130);
or U2566 (N_2566,In_1943,In_422);
or U2567 (N_2567,In_1618,In_446);
nand U2568 (N_2568,In_1548,In_402);
and U2569 (N_2569,In_830,In_252);
and U2570 (N_2570,In_988,In_653);
nand U2571 (N_2571,In_1957,In_1556);
nor U2572 (N_2572,In_186,In_52);
nor U2573 (N_2573,In_1485,In_1442);
nand U2574 (N_2574,In_1028,In_459);
nand U2575 (N_2575,In_110,In_1934);
nor U2576 (N_2576,In_1229,In_412);
and U2577 (N_2577,In_1834,In_390);
or U2578 (N_2578,In_311,In_1394);
nor U2579 (N_2579,In_1296,In_231);
nor U2580 (N_2580,In_142,In_1836);
and U2581 (N_2581,In_1582,In_793);
or U2582 (N_2582,In_1852,In_1701);
xor U2583 (N_2583,In_92,In_829);
or U2584 (N_2584,In_524,In_344);
or U2585 (N_2585,In_1373,In_251);
nand U2586 (N_2586,In_46,In_807);
and U2587 (N_2587,In_1016,In_1975);
nand U2588 (N_2588,In_765,In_562);
nor U2589 (N_2589,In_1927,In_760);
and U2590 (N_2590,In_1295,In_1891);
or U2591 (N_2591,In_358,In_909);
nor U2592 (N_2592,In_1055,In_997);
nand U2593 (N_2593,In_1608,In_1705);
and U2594 (N_2594,In_1790,In_371);
nand U2595 (N_2595,In_1491,In_622);
nand U2596 (N_2596,In_302,In_1539);
and U2597 (N_2597,In_713,In_955);
and U2598 (N_2598,In_1833,In_1481);
nand U2599 (N_2599,In_241,In_993);
nor U2600 (N_2600,In_1545,In_1488);
nand U2601 (N_2601,In_1447,In_908);
or U2602 (N_2602,In_221,In_1620);
and U2603 (N_2603,In_1148,In_1316);
nand U2604 (N_2604,In_98,In_1891);
or U2605 (N_2605,In_1550,In_1078);
and U2606 (N_2606,In_1771,In_1467);
or U2607 (N_2607,In_516,In_868);
nor U2608 (N_2608,In_1743,In_478);
xor U2609 (N_2609,In_1837,In_698);
or U2610 (N_2610,In_960,In_921);
nand U2611 (N_2611,In_1416,In_1665);
and U2612 (N_2612,In_230,In_1192);
and U2613 (N_2613,In_863,In_993);
nor U2614 (N_2614,In_996,In_961);
and U2615 (N_2615,In_251,In_778);
nand U2616 (N_2616,In_46,In_1521);
and U2617 (N_2617,In_1447,In_1717);
xor U2618 (N_2618,In_1560,In_679);
or U2619 (N_2619,In_268,In_1640);
nand U2620 (N_2620,In_309,In_1280);
xnor U2621 (N_2621,In_1235,In_1955);
nor U2622 (N_2622,In_1494,In_347);
or U2623 (N_2623,In_865,In_91);
xor U2624 (N_2624,In_148,In_943);
nor U2625 (N_2625,In_559,In_1042);
and U2626 (N_2626,In_725,In_1861);
or U2627 (N_2627,In_588,In_513);
nor U2628 (N_2628,In_613,In_1540);
nor U2629 (N_2629,In_824,In_68);
nor U2630 (N_2630,In_280,In_1476);
or U2631 (N_2631,In_102,In_1638);
nor U2632 (N_2632,In_1182,In_696);
nand U2633 (N_2633,In_1446,In_911);
or U2634 (N_2634,In_47,In_1231);
nor U2635 (N_2635,In_125,In_638);
nand U2636 (N_2636,In_1424,In_707);
nand U2637 (N_2637,In_14,In_1247);
nor U2638 (N_2638,In_1400,In_1328);
nor U2639 (N_2639,In_1024,In_273);
nand U2640 (N_2640,In_351,In_757);
or U2641 (N_2641,In_537,In_782);
nor U2642 (N_2642,In_1977,In_603);
nor U2643 (N_2643,In_1236,In_1341);
and U2644 (N_2644,In_516,In_462);
or U2645 (N_2645,In_1720,In_637);
nand U2646 (N_2646,In_1631,In_1777);
nand U2647 (N_2647,In_1837,In_948);
nand U2648 (N_2648,In_294,In_767);
or U2649 (N_2649,In_934,In_888);
nor U2650 (N_2650,In_182,In_88);
nor U2651 (N_2651,In_1558,In_999);
nand U2652 (N_2652,In_705,In_1860);
nor U2653 (N_2653,In_1351,In_180);
and U2654 (N_2654,In_1409,In_564);
nand U2655 (N_2655,In_1309,In_491);
or U2656 (N_2656,In_602,In_269);
xnor U2657 (N_2657,In_427,In_1499);
and U2658 (N_2658,In_198,In_1834);
nor U2659 (N_2659,In_1370,In_471);
and U2660 (N_2660,In_1582,In_1147);
or U2661 (N_2661,In_1783,In_514);
nor U2662 (N_2662,In_1276,In_304);
nor U2663 (N_2663,In_1740,In_1542);
or U2664 (N_2664,In_1538,In_1296);
xnor U2665 (N_2665,In_606,In_1464);
nand U2666 (N_2666,In_1863,In_1406);
or U2667 (N_2667,In_1459,In_237);
and U2668 (N_2668,In_1124,In_1740);
nor U2669 (N_2669,In_1602,In_564);
xor U2670 (N_2670,In_807,In_1548);
or U2671 (N_2671,In_1392,In_1277);
nor U2672 (N_2672,In_1976,In_285);
nor U2673 (N_2673,In_310,In_1660);
or U2674 (N_2674,In_738,In_1483);
and U2675 (N_2675,In_1908,In_397);
and U2676 (N_2676,In_1542,In_653);
nand U2677 (N_2677,In_1424,In_1076);
nand U2678 (N_2678,In_33,In_1181);
nor U2679 (N_2679,In_172,In_985);
xor U2680 (N_2680,In_573,In_192);
nand U2681 (N_2681,In_501,In_329);
nand U2682 (N_2682,In_789,In_809);
nor U2683 (N_2683,In_915,In_78);
and U2684 (N_2684,In_981,In_637);
nand U2685 (N_2685,In_333,In_308);
nand U2686 (N_2686,In_90,In_716);
or U2687 (N_2687,In_94,In_1035);
nand U2688 (N_2688,In_1746,In_1796);
and U2689 (N_2689,In_1961,In_247);
and U2690 (N_2690,In_154,In_159);
or U2691 (N_2691,In_449,In_1416);
or U2692 (N_2692,In_1069,In_619);
or U2693 (N_2693,In_1259,In_1653);
nor U2694 (N_2694,In_1411,In_425);
and U2695 (N_2695,In_884,In_1425);
and U2696 (N_2696,In_1875,In_740);
xnor U2697 (N_2697,In_1639,In_1605);
and U2698 (N_2698,In_781,In_707);
nand U2699 (N_2699,In_432,In_1597);
nor U2700 (N_2700,In_176,In_1939);
nor U2701 (N_2701,In_544,In_1885);
nand U2702 (N_2702,In_1522,In_887);
and U2703 (N_2703,In_871,In_1624);
or U2704 (N_2704,In_13,In_538);
nor U2705 (N_2705,In_387,In_85);
xor U2706 (N_2706,In_1435,In_158);
nand U2707 (N_2707,In_302,In_1431);
nor U2708 (N_2708,In_776,In_1553);
nor U2709 (N_2709,In_1019,In_1407);
or U2710 (N_2710,In_1903,In_114);
nor U2711 (N_2711,In_475,In_1009);
nand U2712 (N_2712,In_1215,In_1011);
and U2713 (N_2713,In_517,In_1296);
or U2714 (N_2714,In_843,In_1453);
or U2715 (N_2715,In_126,In_1316);
nand U2716 (N_2716,In_1618,In_1690);
nor U2717 (N_2717,In_1071,In_1468);
or U2718 (N_2718,In_655,In_883);
and U2719 (N_2719,In_609,In_1138);
or U2720 (N_2720,In_113,In_180);
nor U2721 (N_2721,In_1817,In_275);
or U2722 (N_2722,In_1535,In_1350);
nor U2723 (N_2723,In_577,In_346);
and U2724 (N_2724,In_1354,In_280);
or U2725 (N_2725,In_1743,In_662);
xnor U2726 (N_2726,In_492,In_447);
or U2727 (N_2727,In_449,In_763);
nand U2728 (N_2728,In_1527,In_170);
nand U2729 (N_2729,In_60,In_560);
or U2730 (N_2730,In_849,In_1139);
nand U2731 (N_2731,In_1195,In_655);
nor U2732 (N_2732,In_1211,In_633);
nand U2733 (N_2733,In_704,In_1788);
or U2734 (N_2734,In_969,In_1155);
nor U2735 (N_2735,In_1295,In_1134);
or U2736 (N_2736,In_1151,In_6);
xor U2737 (N_2737,In_281,In_1429);
xnor U2738 (N_2738,In_899,In_646);
nand U2739 (N_2739,In_1412,In_492);
xor U2740 (N_2740,In_1803,In_1436);
or U2741 (N_2741,In_473,In_1928);
or U2742 (N_2742,In_1168,In_813);
or U2743 (N_2743,In_1285,In_1143);
nand U2744 (N_2744,In_1478,In_978);
nand U2745 (N_2745,In_952,In_1543);
or U2746 (N_2746,In_1317,In_245);
or U2747 (N_2747,In_1208,In_1046);
and U2748 (N_2748,In_1684,In_1806);
and U2749 (N_2749,In_437,In_899);
or U2750 (N_2750,In_1688,In_1663);
nor U2751 (N_2751,In_111,In_1656);
nand U2752 (N_2752,In_1168,In_1207);
nand U2753 (N_2753,In_888,In_387);
xor U2754 (N_2754,In_1055,In_312);
nor U2755 (N_2755,In_266,In_1439);
nor U2756 (N_2756,In_1075,In_398);
nor U2757 (N_2757,In_1356,In_254);
nor U2758 (N_2758,In_1444,In_392);
and U2759 (N_2759,In_1192,In_764);
xor U2760 (N_2760,In_1304,In_1269);
or U2761 (N_2761,In_1943,In_1124);
and U2762 (N_2762,In_353,In_1027);
nand U2763 (N_2763,In_1960,In_1917);
and U2764 (N_2764,In_902,In_1745);
nand U2765 (N_2765,In_722,In_1582);
nand U2766 (N_2766,In_409,In_1474);
xor U2767 (N_2767,In_835,In_369);
xor U2768 (N_2768,In_677,In_1318);
and U2769 (N_2769,In_1305,In_1933);
and U2770 (N_2770,In_1360,In_494);
nor U2771 (N_2771,In_1250,In_1153);
nor U2772 (N_2772,In_152,In_595);
or U2773 (N_2773,In_354,In_714);
nand U2774 (N_2774,In_106,In_1521);
nand U2775 (N_2775,In_43,In_883);
or U2776 (N_2776,In_1653,In_1749);
xor U2777 (N_2777,In_1749,In_1262);
nor U2778 (N_2778,In_639,In_702);
and U2779 (N_2779,In_1357,In_1883);
nand U2780 (N_2780,In_224,In_1243);
or U2781 (N_2781,In_1468,In_930);
nand U2782 (N_2782,In_834,In_389);
and U2783 (N_2783,In_179,In_1408);
nor U2784 (N_2784,In_1849,In_1266);
and U2785 (N_2785,In_369,In_1669);
and U2786 (N_2786,In_1168,In_170);
or U2787 (N_2787,In_392,In_1730);
nor U2788 (N_2788,In_339,In_333);
and U2789 (N_2789,In_482,In_315);
or U2790 (N_2790,In_1245,In_1836);
nor U2791 (N_2791,In_127,In_162);
nor U2792 (N_2792,In_350,In_610);
nor U2793 (N_2793,In_187,In_1295);
or U2794 (N_2794,In_896,In_696);
nor U2795 (N_2795,In_100,In_1864);
nor U2796 (N_2796,In_707,In_1521);
nand U2797 (N_2797,In_1013,In_1228);
nand U2798 (N_2798,In_1908,In_735);
or U2799 (N_2799,In_217,In_1010);
nand U2800 (N_2800,In_923,In_712);
and U2801 (N_2801,In_530,In_340);
and U2802 (N_2802,In_1927,In_1421);
nor U2803 (N_2803,In_1771,In_297);
and U2804 (N_2804,In_1823,In_517);
or U2805 (N_2805,In_834,In_829);
nor U2806 (N_2806,In_1674,In_1318);
nand U2807 (N_2807,In_446,In_215);
or U2808 (N_2808,In_1583,In_933);
nand U2809 (N_2809,In_1669,In_1520);
nand U2810 (N_2810,In_537,In_1654);
xnor U2811 (N_2811,In_817,In_1223);
or U2812 (N_2812,In_1919,In_1376);
nand U2813 (N_2813,In_1984,In_1425);
and U2814 (N_2814,In_792,In_1249);
or U2815 (N_2815,In_756,In_1451);
and U2816 (N_2816,In_683,In_1052);
or U2817 (N_2817,In_363,In_515);
nand U2818 (N_2818,In_1249,In_1357);
nor U2819 (N_2819,In_1525,In_1988);
nor U2820 (N_2820,In_647,In_101);
and U2821 (N_2821,In_1430,In_729);
nor U2822 (N_2822,In_1394,In_722);
or U2823 (N_2823,In_716,In_1286);
or U2824 (N_2824,In_1797,In_637);
nand U2825 (N_2825,In_1850,In_1504);
nand U2826 (N_2826,In_105,In_115);
nand U2827 (N_2827,In_1642,In_1882);
or U2828 (N_2828,In_53,In_463);
and U2829 (N_2829,In_808,In_952);
nand U2830 (N_2830,In_1310,In_59);
and U2831 (N_2831,In_194,In_1048);
nor U2832 (N_2832,In_1875,In_380);
or U2833 (N_2833,In_1490,In_290);
nand U2834 (N_2834,In_1921,In_1598);
nand U2835 (N_2835,In_1470,In_1949);
nor U2836 (N_2836,In_1745,In_673);
or U2837 (N_2837,In_511,In_840);
or U2838 (N_2838,In_140,In_1467);
nand U2839 (N_2839,In_900,In_1014);
or U2840 (N_2840,In_1749,In_645);
and U2841 (N_2841,In_563,In_1151);
or U2842 (N_2842,In_200,In_679);
xor U2843 (N_2843,In_465,In_1738);
or U2844 (N_2844,In_347,In_1917);
nand U2845 (N_2845,In_1166,In_1943);
nor U2846 (N_2846,In_1501,In_1095);
and U2847 (N_2847,In_1026,In_35);
nand U2848 (N_2848,In_1631,In_841);
or U2849 (N_2849,In_253,In_262);
or U2850 (N_2850,In_1291,In_732);
nand U2851 (N_2851,In_112,In_591);
nor U2852 (N_2852,In_1411,In_6);
and U2853 (N_2853,In_457,In_992);
nor U2854 (N_2854,In_1323,In_633);
nand U2855 (N_2855,In_612,In_108);
nor U2856 (N_2856,In_1891,In_14);
or U2857 (N_2857,In_1297,In_23);
or U2858 (N_2858,In_332,In_678);
nor U2859 (N_2859,In_1982,In_862);
nand U2860 (N_2860,In_549,In_37);
and U2861 (N_2861,In_349,In_465);
xor U2862 (N_2862,In_1686,In_1837);
nor U2863 (N_2863,In_717,In_468);
nor U2864 (N_2864,In_1552,In_912);
or U2865 (N_2865,In_1039,In_1987);
and U2866 (N_2866,In_1097,In_913);
nand U2867 (N_2867,In_905,In_1813);
nor U2868 (N_2868,In_491,In_965);
nor U2869 (N_2869,In_571,In_7);
and U2870 (N_2870,In_1076,In_546);
or U2871 (N_2871,In_1584,In_1432);
and U2872 (N_2872,In_560,In_643);
or U2873 (N_2873,In_450,In_511);
nand U2874 (N_2874,In_1183,In_414);
nand U2875 (N_2875,In_730,In_1772);
and U2876 (N_2876,In_270,In_576);
and U2877 (N_2877,In_913,In_949);
and U2878 (N_2878,In_1165,In_258);
and U2879 (N_2879,In_1117,In_312);
or U2880 (N_2880,In_333,In_1174);
or U2881 (N_2881,In_680,In_823);
nand U2882 (N_2882,In_933,In_642);
and U2883 (N_2883,In_1562,In_33);
nand U2884 (N_2884,In_1390,In_526);
nor U2885 (N_2885,In_519,In_1626);
nor U2886 (N_2886,In_1534,In_41);
or U2887 (N_2887,In_810,In_1449);
nor U2888 (N_2888,In_1832,In_231);
nand U2889 (N_2889,In_1366,In_693);
nand U2890 (N_2890,In_1114,In_426);
and U2891 (N_2891,In_530,In_179);
and U2892 (N_2892,In_1743,In_1482);
nor U2893 (N_2893,In_1133,In_1947);
xor U2894 (N_2894,In_1837,In_1741);
and U2895 (N_2895,In_1390,In_498);
nor U2896 (N_2896,In_1120,In_127);
nand U2897 (N_2897,In_1641,In_1155);
nor U2898 (N_2898,In_541,In_362);
or U2899 (N_2899,In_1051,In_1029);
and U2900 (N_2900,In_1137,In_1052);
nand U2901 (N_2901,In_1494,In_748);
nand U2902 (N_2902,In_943,In_992);
nor U2903 (N_2903,In_1269,In_1183);
or U2904 (N_2904,In_17,In_115);
nand U2905 (N_2905,In_1792,In_82);
nor U2906 (N_2906,In_405,In_1681);
or U2907 (N_2907,In_124,In_1877);
and U2908 (N_2908,In_1356,In_1043);
or U2909 (N_2909,In_1818,In_452);
and U2910 (N_2910,In_1957,In_847);
nand U2911 (N_2911,In_1444,In_730);
nand U2912 (N_2912,In_776,In_321);
and U2913 (N_2913,In_1085,In_375);
nand U2914 (N_2914,In_1298,In_385);
or U2915 (N_2915,In_1910,In_1298);
nor U2916 (N_2916,In_1656,In_1795);
xor U2917 (N_2917,In_1710,In_1266);
and U2918 (N_2918,In_1803,In_1560);
or U2919 (N_2919,In_251,In_313);
nor U2920 (N_2920,In_520,In_753);
and U2921 (N_2921,In_1259,In_107);
nand U2922 (N_2922,In_174,In_1829);
and U2923 (N_2923,In_474,In_1477);
xnor U2924 (N_2924,In_1533,In_357);
or U2925 (N_2925,In_1292,In_1412);
or U2926 (N_2926,In_756,In_899);
nand U2927 (N_2927,In_470,In_688);
nand U2928 (N_2928,In_809,In_1042);
nand U2929 (N_2929,In_1571,In_1587);
nor U2930 (N_2930,In_701,In_194);
nand U2931 (N_2931,In_184,In_409);
or U2932 (N_2932,In_1195,In_1629);
and U2933 (N_2933,In_1718,In_628);
nor U2934 (N_2934,In_598,In_1309);
and U2935 (N_2935,In_1157,In_805);
nor U2936 (N_2936,In_1517,In_1652);
nor U2937 (N_2937,In_802,In_1403);
or U2938 (N_2938,In_1494,In_1510);
nand U2939 (N_2939,In_1193,In_539);
nor U2940 (N_2940,In_1268,In_818);
and U2941 (N_2941,In_852,In_1046);
and U2942 (N_2942,In_8,In_1288);
xor U2943 (N_2943,In_1555,In_230);
and U2944 (N_2944,In_1502,In_591);
nor U2945 (N_2945,In_779,In_569);
or U2946 (N_2946,In_1212,In_1686);
nor U2947 (N_2947,In_1674,In_1312);
or U2948 (N_2948,In_598,In_1383);
nand U2949 (N_2949,In_1587,In_702);
nand U2950 (N_2950,In_1581,In_767);
or U2951 (N_2951,In_234,In_684);
or U2952 (N_2952,In_1782,In_1639);
or U2953 (N_2953,In_91,In_1860);
and U2954 (N_2954,In_919,In_1175);
nor U2955 (N_2955,In_1601,In_1203);
xnor U2956 (N_2956,In_579,In_1049);
or U2957 (N_2957,In_1495,In_1616);
and U2958 (N_2958,In_516,In_215);
or U2959 (N_2959,In_1040,In_1409);
xnor U2960 (N_2960,In_1099,In_167);
nand U2961 (N_2961,In_699,In_1633);
nor U2962 (N_2962,In_406,In_793);
nand U2963 (N_2963,In_1670,In_1237);
xnor U2964 (N_2964,In_331,In_1164);
and U2965 (N_2965,In_1666,In_1681);
and U2966 (N_2966,In_1469,In_268);
and U2967 (N_2967,In_1473,In_1084);
nand U2968 (N_2968,In_934,In_1835);
xnor U2969 (N_2969,In_1860,In_507);
or U2970 (N_2970,In_1325,In_589);
xor U2971 (N_2971,In_403,In_154);
or U2972 (N_2972,In_1896,In_150);
nand U2973 (N_2973,In_1614,In_1280);
and U2974 (N_2974,In_1949,In_1126);
xnor U2975 (N_2975,In_865,In_129);
and U2976 (N_2976,In_1032,In_1789);
or U2977 (N_2977,In_438,In_1946);
xnor U2978 (N_2978,In_284,In_944);
nor U2979 (N_2979,In_1138,In_852);
nand U2980 (N_2980,In_1257,In_213);
nand U2981 (N_2981,In_1248,In_1065);
and U2982 (N_2982,In_1637,In_1978);
and U2983 (N_2983,In_316,In_206);
nand U2984 (N_2984,In_872,In_871);
nand U2985 (N_2985,In_520,In_617);
nor U2986 (N_2986,In_906,In_815);
nand U2987 (N_2987,In_106,In_957);
xor U2988 (N_2988,In_1454,In_200);
or U2989 (N_2989,In_993,In_1357);
xor U2990 (N_2990,In_334,In_525);
nor U2991 (N_2991,In_1839,In_1609);
nand U2992 (N_2992,In_1358,In_1815);
or U2993 (N_2993,In_588,In_1744);
and U2994 (N_2994,In_1541,In_1276);
or U2995 (N_2995,In_976,In_1887);
nand U2996 (N_2996,In_10,In_86);
nand U2997 (N_2997,In_247,In_998);
nor U2998 (N_2998,In_677,In_478);
nor U2999 (N_2999,In_27,In_661);
nand U3000 (N_3000,In_1990,In_991);
or U3001 (N_3001,In_6,In_600);
xnor U3002 (N_3002,In_952,In_1805);
nor U3003 (N_3003,In_812,In_480);
nor U3004 (N_3004,In_997,In_215);
xor U3005 (N_3005,In_696,In_1304);
and U3006 (N_3006,In_793,In_1743);
xnor U3007 (N_3007,In_1109,In_856);
nor U3008 (N_3008,In_1141,In_1777);
nor U3009 (N_3009,In_811,In_925);
nor U3010 (N_3010,In_748,In_590);
nand U3011 (N_3011,In_534,In_1806);
xor U3012 (N_3012,In_1972,In_166);
nor U3013 (N_3013,In_519,In_470);
nand U3014 (N_3014,In_1326,In_866);
nor U3015 (N_3015,In_1810,In_97);
nor U3016 (N_3016,In_1845,In_1699);
xor U3017 (N_3017,In_943,In_113);
nor U3018 (N_3018,In_1702,In_315);
and U3019 (N_3019,In_942,In_1531);
nor U3020 (N_3020,In_121,In_1586);
xnor U3021 (N_3021,In_1474,In_1246);
nand U3022 (N_3022,In_295,In_888);
nor U3023 (N_3023,In_345,In_259);
or U3024 (N_3024,In_61,In_1670);
nand U3025 (N_3025,In_1193,In_1770);
nand U3026 (N_3026,In_684,In_918);
nor U3027 (N_3027,In_604,In_151);
xor U3028 (N_3028,In_960,In_1038);
or U3029 (N_3029,In_1499,In_1352);
nand U3030 (N_3030,In_564,In_1242);
or U3031 (N_3031,In_338,In_828);
nor U3032 (N_3032,In_1693,In_452);
or U3033 (N_3033,In_383,In_930);
and U3034 (N_3034,In_1225,In_60);
nor U3035 (N_3035,In_952,In_1043);
xor U3036 (N_3036,In_1140,In_464);
xnor U3037 (N_3037,In_1850,In_1362);
and U3038 (N_3038,In_1845,In_446);
nand U3039 (N_3039,In_485,In_1468);
nor U3040 (N_3040,In_823,In_32);
xnor U3041 (N_3041,In_1891,In_328);
xor U3042 (N_3042,In_1504,In_1529);
and U3043 (N_3043,In_1687,In_352);
and U3044 (N_3044,In_1222,In_952);
nand U3045 (N_3045,In_1886,In_410);
nor U3046 (N_3046,In_461,In_1721);
xnor U3047 (N_3047,In_861,In_868);
and U3048 (N_3048,In_128,In_231);
xor U3049 (N_3049,In_1445,In_553);
and U3050 (N_3050,In_880,In_1961);
or U3051 (N_3051,In_782,In_1836);
or U3052 (N_3052,In_1022,In_1153);
nor U3053 (N_3053,In_1499,In_1092);
or U3054 (N_3054,In_1592,In_825);
and U3055 (N_3055,In_529,In_143);
nor U3056 (N_3056,In_1305,In_38);
and U3057 (N_3057,In_403,In_682);
nor U3058 (N_3058,In_1224,In_819);
or U3059 (N_3059,In_1908,In_1502);
nor U3060 (N_3060,In_1464,In_1020);
and U3061 (N_3061,In_711,In_1694);
nor U3062 (N_3062,In_459,In_1470);
or U3063 (N_3063,In_1059,In_1649);
nor U3064 (N_3064,In_373,In_767);
and U3065 (N_3065,In_293,In_383);
nand U3066 (N_3066,In_131,In_653);
and U3067 (N_3067,In_948,In_1392);
or U3068 (N_3068,In_362,In_1134);
or U3069 (N_3069,In_1471,In_418);
or U3070 (N_3070,In_954,In_10);
nand U3071 (N_3071,In_1081,In_1818);
or U3072 (N_3072,In_1102,In_1034);
nand U3073 (N_3073,In_908,In_437);
or U3074 (N_3074,In_1956,In_1675);
nand U3075 (N_3075,In_1678,In_307);
nand U3076 (N_3076,In_674,In_692);
or U3077 (N_3077,In_862,In_320);
nor U3078 (N_3078,In_263,In_17);
and U3079 (N_3079,In_1283,In_955);
nand U3080 (N_3080,In_89,In_699);
nor U3081 (N_3081,In_1921,In_1596);
and U3082 (N_3082,In_1426,In_631);
xnor U3083 (N_3083,In_571,In_531);
nand U3084 (N_3084,In_1385,In_802);
or U3085 (N_3085,In_1248,In_302);
nor U3086 (N_3086,In_244,In_1454);
nand U3087 (N_3087,In_4,In_223);
and U3088 (N_3088,In_1068,In_490);
xor U3089 (N_3089,In_1980,In_1618);
and U3090 (N_3090,In_855,In_980);
nor U3091 (N_3091,In_1990,In_1804);
nor U3092 (N_3092,In_715,In_1549);
nor U3093 (N_3093,In_1918,In_613);
nand U3094 (N_3094,In_1586,In_1119);
and U3095 (N_3095,In_1590,In_321);
or U3096 (N_3096,In_740,In_1868);
or U3097 (N_3097,In_928,In_1100);
nand U3098 (N_3098,In_1172,In_805);
and U3099 (N_3099,In_1217,In_1777);
and U3100 (N_3100,In_1313,In_1931);
and U3101 (N_3101,In_1322,In_116);
nand U3102 (N_3102,In_1486,In_984);
nor U3103 (N_3103,In_499,In_752);
or U3104 (N_3104,In_1694,In_36);
nor U3105 (N_3105,In_1871,In_534);
and U3106 (N_3106,In_1177,In_1632);
or U3107 (N_3107,In_809,In_1257);
nor U3108 (N_3108,In_62,In_726);
nor U3109 (N_3109,In_1573,In_1010);
nand U3110 (N_3110,In_1351,In_840);
nand U3111 (N_3111,In_728,In_161);
nand U3112 (N_3112,In_1881,In_458);
nor U3113 (N_3113,In_1685,In_834);
nand U3114 (N_3114,In_578,In_1222);
or U3115 (N_3115,In_1115,In_685);
nor U3116 (N_3116,In_430,In_1961);
or U3117 (N_3117,In_159,In_402);
nand U3118 (N_3118,In_1770,In_1720);
nand U3119 (N_3119,In_27,In_133);
nand U3120 (N_3120,In_45,In_580);
nand U3121 (N_3121,In_1445,In_848);
and U3122 (N_3122,In_1905,In_1243);
or U3123 (N_3123,In_653,In_871);
nand U3124 (N_3124,In_537,In_1202);
and U3125 (N_3125,In_117,In_1985);
nor U3126 (N_3126,In_1510,In_1632);
and U3127 (N_3127,In_667,In_1898);
nor U3128 (N_3128,In_1815,In_331);
nand U3129 (N_3129,In_1013,In_914);
nand U3130 (N_3130,In_1352,In_589);
or U3131 (N_3131,In_478,In_1142);
nor U3132 (N_3132,In_131,In_1157);
and U3133 (N_3133,In_1996,In_456);
and U3134 (N_3134,In_654,In_1149);
or U3135 (N_3135,In_36,In_197);
nand U3136 (N_3136,In_1296,In_1814);
and U3137 (N_3137,In_1987,In_105);
nor U3138 (N_3138,In_1068,In_1239);
nor U3139 (N_3139,In_207,In_637);
nor U3140 (N_3140,In_1826,In_1327);
and U3141 (N_3141,In_1734,In_1121);
xnor U3142 (N_3142,In_1178,In_1094);
nor U3143 (N_3143,In_99,In_817);
or U3144 (N_3144,In_1186,In_1157);
and U3145 (N_3145,In_1738,In_948);
and U3146 (N_3146,In_836,In_418);
or U3147 (N_3147,In_196,In_810);
or U3148 (N_3148,In_927,In_1263);
nor U3149 (N_3149,In_1180,In_1009);
or U3150 (N_3150,In_662,In_1362);
and U3151 (N_3151,In_1563,In_885);
or U3152 (N_3152,In_159,In_529);
or U3153 (N_3153,In_87,In_807);
xnor U3154 (N_3154,In_721,In_1358);
nor U3155 (N_3155,In_1669,In_1950);
and U3156 (N_3156,In_343,In_633);
nor U3157 (N_3157,In_365,In_106);
xor U3158 (N_3158,In_1822,In_887);
nor U3159 (N_3159,In_106,In_1322);
and U3160 (N_3160,In_1481,In_1220);
nor U3161 (N_3161,In_1218,In_836);
xnor U3162 (N_3162,In_1456,In_1121);
nand U3163 (N_3163,In_1927,In_90);
or U3164 (N_3164,In_152,In_609);
or U3165 (N_3165,In_697,In_1530);
xor U3166 (N_3166,In_1766,In_990);
and U3167 (N_3167,In_995,In_1255);
nand U3168 (N_3168,In_1407,In_772);
nor U3169 (N_3169,In_469,In_300);
nand U3170 (N_3170,In_1546,In_773);
nor U3171 (N_3171,In_128,In_893);
and U3172 (N_3172,In_528,In_489);
and U3173 (N_3173,In_848,In_1702);
nor U3174 (N_3174,In_1825,In_1263);
or U3175 (N_3175,In_1946,In_589);
or U3176 (N_3176,In_493,In_764);
nor U3177 (N_3177,In_655,In_336);
and U3178 (N_3178,In_1654,In_954);
and U3179 (N_3179,In_765,In_1692);
and U3180 (N_3180,In_853,In_978);
nand U3181 (N_3181,In_420,In_354);
and U3182 (N_3182,In_763,In_1594);
nand U3183 (N_3183,In_1131,In_1804);
or U3184 (N_3184,In_960,In_510);
nand U3185 (N_3185,In_1808,In_347);
or U3186 (N_3186,In_1483,In_890);
nor U3187 (N_3187,In_601,In_1124);
and U3188 (N_3188,In_50,In_560);
nor U3189 (N_3189,In_1641,In_543);
nor U3190 (N_3190,In_425,In_1034);
nor U3191 (N_3191,In_148,In_32);
nor U3192 (N_3192,In_76,In_1757);
nor U3193 (N_3193,In_1448,In_53);
nand U3194 (N_3194,In_218,In_1975);
nor U3195 (N_3195,In_1077,In_725);
or U3196 (N_3196,In_507,In_1974);
or U3197 (N_3197,In_528,In_1440);
xor U3198 (N_3198,In_1096,In_478);
and U3199 (N_3199,In_1079,In_583);
and U3200 (N_3200,In_445,In_456);
nand U3201 (N_3201,In_1584,In_388);
and U3202 (N_3202,In_1049,In_773);
nand U3203 (N_3203,In_436,In_868);
nand U3204 (N_3204,In_117,In_408);
xor U3205 (N_3205,In_246,In_269);
nand U3206 (N_3206,In_398,In_1492);
and U3207 (N_3207,In_969,In_45);
and U3208 (N_3208,In_1199,In_702);
and U3209 (N_3209,In_1326,In_373);
or U3210 (N_3210,In_1079,In_1539);
nor U3211 (N_3211,In_112,In_877);
nand U3212 (N_3212,In_1438,In_479);
nor U3213 (N_3213,In_116,In_522);
nand U3214 (N_3214,In_359,In_605);
nand U3215 (N_3215,In_1996,In_1746);
or U3216 (N_3216,In_669,In_1250);
nand U3217 (N_3217,In_286,In_1802);
and U3218 (N_3218,In_1960,In_31);
and U3219 (N_3219,In_126,In_1465);
xnor U3220 (N_3220,In_1104,In_197);
nand U3221 (N_3221,In_882,In_1132);
nand U3222 (N_3222,In_1257,In_349);
and U3223 (N_3223,In_1094,In_345);
and U3224 (N_3224,In_464,In_532);
nand U3225 (N_3225,In_482,In_1751);
nor U3226 (N_3226,In_1892,In_1891);
nand U3227 (N_3227,In_316,In_1460);
nor U3228 (N_3228,In_1424,In_693);
nand U3229 (N_3229,In_412,In_1194);
and U3230 (N_3230,In_803,In_196);
and U3231 (N_3231,In_11,In_323);
and U3232 (N_3232,In_1163,In_1205);
nand U3233 (N_3233,In_277,In_614);
and U3234 (N_3234,In_1035,In_1965);
or U3235 (N_3235,In_202,In_1516);
and U3236 (N_3236,In_1768,In_1304);
nand U3237 (N_3237,In_1578,In_672);
nor U3238 (N_3238,In_1128,In_813);
nor U3239 (N_3239,In_425,In_1537);
nor U3240 (N_3240,In_670,In_1565);
nand U3241 (N_3241,In_1027,In_982);
nor U3242 (N_3242,In_519,In_840);
and U3243 (N_3243,In_1509,In_667);
and U3244 (N_3244,In_884,In_1239);
or U3245 (N_3245,In_1181,In_261);
and U3246 (N_3246,In_1654,In_1599);
xnor U3247 (N_3247,In_1495,In_891);
nor U3248 (N_3248,In_1283,In_269);
or U3249 (N_3249,In_1334,In_1328);
nor U3250 (N_3250,In_987,In_1649);
nand U3251 (N_3251,In_1290,In_1652);
and U3252 (N_3252,In_896,In_461);
nand U3253 (N_3253,In_514,In_367);
or U3254 (N_3254,In_572,In_691);
xnor U3255 (N_3255,In_268,In_166);
nor U3256 (N_3256,In_260,In_1990);
nor U3257 (N_3257,In_1326,In_76);
and U3258 (N_3258,In_1121,In_1520);
nand U3259 (N_3259,In_1529,In_865);
nand U3260 (N_3260,In_1266,In_1537);
and U3261 (N_3261,In_1914,In_1038);
and U3262 (N_3262,In_12,In_1189);
nor U3263 (N_3263,In_998,In_1974);
nand U3264 (N_3264,In_394,In_1325);
and U3265 (N_3265,In_1946,In_1414);
and U3266 (N_3266,In_77,In_1832);
and U3267 (N_3267,In_878,In_315);
nand U3268 (N_3268,In_1856,In_1402);
and U3269 (N_3269,In_624,In_1403);
nand U3270 (N_3270,In_1876,In_79);
xnor U3271 (N_3271,In_1598,In_1621);
nand U3272 (N_3272,In_1257,In_1695);
nand U3273 (N_3273,In_878,In_352);
or U3274 (N_3274,In_635,In_763);
nor U3275 (N_3275,In_260,In_192);
nand U3276 (N_3276,In_1873,In_631);
and U3277 (N_3277,In_1010,In_663);
and U3278 (N_3278,In_1711,In_627);
or U3279 (N_3279,In_377,In_1288);
nor U3280 (N_3280,In_1888,In_491);
nor U3281 (N_3281,In_1487,In_1628);
and U3282 (N_3282,In_1098,In_920);
nand U3283 (N_3283,In_475,In_1977);
and U3284 (N_3284,In_152,In_1964);
and U3285 (N_3285,In_1783,In_1375);
nand U3286 (N_3286,In_1138,In_814);
and U3287 (N_3287,In_1361,In_878);
or U3288 (N_3288,In_1727,In_439);
xor U3289 (N_3289,In_1313,In_294);
or U3290 (N_3290,In_1316,In_1893);
and U3291 (N_3291,In_728,In_1405);
nand U3292 (N_3292,In_1446,In_314);
nor U3293 (N_3293,In_540,In_442);
and U3294 (N_3294,In_1952,In_1611);
nand U3295 (N_3295,In_832,In_865);
nand U3296 (N_3296,In_1462,In_1400);
nand U3297 (N_3297,In_792,In_106);
nor U3298 (N_3298,In_427,In_1723);
nand U3299 (N_3299,In_1436,In_409);
nand U3300 (N_3300,In_769,In_417);
and U3301 (N_3301,In_229,In_1173);
nand U3302 (N_3302,In_1074,In_1983);
xor U3303 (N_3303,In_1937,In_954);
nand U3304 (N_3304,In_812,In_756);
xnor U3305 (N_3305,In_478,In_247);
and U3306 (N_3306,In_1316,In_1529);
or U3307 (N_3307,In_658,In_1674);
or U3308 (N_3308,In_38,In_1680);
nor U3309 (N_3309,In_540,In_641);
nand U3310 (N_3310,In_1517,In_1816);
and U3311 (N_3311,In_1837,In_1354);
nor U3312 (N_3312,In_1707,In_136);
or U3313 (N_3313,In_1804,In_953);
xor U3314 (N_3314,In_593,In_1959);
xor U3315 (N_3315,In_1751,In_1413);
nor U3316 (N_3316,In_417,In_327);
nor U3317 (N_3317,In_392,In_1414);
xnor U3318 (N_3318,In_1374,In_1654);
and U3319 (N_3319,In_1686,In_1230);
and U3320 (N_3320,In_136,In_388);
nand U3321 (N_3321,In_151,In_1641);
nor U3322 (N_3322,In_1009,In_1724);
nor U3323 (N_3323,In_1432,In_569);
or U3324 (N_3324,In_304,In_446);
nand U3325 (N_3325,In_273,In_1219);
nor U3326 (N_3326,In_661,In_577);
or U3327 (N_3327,In_886,In_922);
nand U3328 (N_3328,In_1912,In_546);
nand U3329 (N_3329,In_1179,In_644);
nor U3330 (N_3330,In_443,In_696);
nand U3331 (N_3331,In_959,In_198);
nand U3332 (N_3332,In_1353,In_257);
and U3333 (N_3333,In_584,In_368);
nor U3334 (N_3334,In_731,In_1505);
or U3335 (N_3335,In_1892,In_1816);
or U3336 (N_3336,In_606,In_207);
or U3337 (N_3337,In_1761,In_117);
nand U3338 (N_3338,In_125,In_1500);
xor U3339 (N_3339,In_371,In_1236);
and U3340 (N_3340,In_1754,In_639);
nand U3341 (N_3341,In_1054,In_198);
nor U3342 (N_3342,In_1646,In_869);
xor U3343 (N_3343,In_1210,In_1222);
xor U3344 (N_3344,In_764,In_787);
xor U3345 (N_3345,In_772,In_692);
nor U3346 (N_3346,In_1936,In_574);
and U3347 (N_3347,In_1593,In_675);
and U3348 (N_3348,In_1974,In_1436);
and U3349 (N_3349,In_413,In_551);
nor U3350 (N_3350,In_869,In_417);
nand U3351 (N_3351,In_1622,In_408);
nor U3352 (N_3352,In_487,In_801);
or U3353 (N_3353,In_265,In_1610);
and U3354 (N_3354,In_1295,In_1481);
xnor U3355 (N_3355,In_1212,In_1539);
nor U3356 (N_3356,In_244,In_1165);
or U3357 (N_3357,In_1511,In_1910);
nand U3358 (N_3358,In_1492,In_1215);
and U3359 (N_3359,In_896,In_1752);
nor U3360 (N_3360,In_585,In_445);
and U3361 (N_3361,In_1547,In_848);
nor U3362 (N_3362,In_352,In_1070);
nor U3363 (N_3363,In_772,In_380);
and U3364 (N_3364,In_1,In_102);
nor U3365 (N_3365,In_962,In_1666);
nand U3366 (N_3366,In_693,In_1683);
or U3367 (N_3367,In_1044,In_953);
nor U3368 (N_3368,In_877,In_1310);
or U3369 (N_3369,In_474,In_952);
and U3370 (N_3370,In_1305,In_1100);
nor U3371 (N_3371,In_545,In_1868);
nor U3372 (N_3372,In_730,In_1465);
xor U3373 (N_3373,In_1563,In_1769);
or U3374 (N_3374,In_1829,In_1130);
or U3375 (N_3375,In_1705,In_1804);
and U3376 (N_3376,In_1146,In_124);
xnor U3377 (N_3377,In_1074,In_391);
nand U3378 (N_3378,In_1647,In_833);
and U3379 (N_3379,In_930,In_49);
and U3380 (N_3380,In_90,In_881);
and U3381 (N_3381,In_1284,In_1847);
and U3382 (N_3382,In_339,In_1262);
or U3383 (N_3383,In_776,In_1444);
xor U3384 (N_3384,In_915,In_1576);
nand U3385 (N_3385,In_82,In_662);
nand U3386 (N_3386,In_1298,In_313);
nor U3387 (N_3387,In_1312,In_279);
xor U3388 (N_3388,In_847,In_1689);
nor U3389 (N_3389,In_1826,In_1064);
nor U3390 (N_3390,In_1197,In_579);
or U3391 (N_3391,In_1434,In_1535);
and U3392 (N_3392,In_394,In_1764);
nand U3393 (N_3393,In_629,In_19);
nor U3394 (N_3394,In_1968,In_857);
nand U3395 (N_3395,In_478,In_312);
and U3396 (N_3396,In_724,In_384);
nand U3397 (N_3397,In_235,In_1823);
nor U3398 (N_3398,In_351,In_1656);
nand U3399 (N_3399,In_577,In_320);
and U3400 (N_3400,In_852,In_688);
xnor U3401 (N_3401,In_416,In_45);
or U3402 (N_3402,In_1320,In_1773);
or U3403 (N_3403,In_1078,In_1443);
or U3404 (N_3404,In_770,In_569);
nand U3405 (N_3405,In_1604,In_1016);
or U3406 (N_3406,In_1796,In_1359);
or U3407 (N_3407,In_498,In_1588);
xor U3408 (N_3408,In_1807,In_1393);
nor U3409 (N_3409,In_1210,In_831);
and U3410 (N_3410,In_26,In_1586);
and U3411 (N_3411,In_253,In_1081);
nor U3412 (N_3412,In_1294,In_1673);
nor U3413 (N_3413,In_1217,In_152);
nor U3414 (N_3414,In_1821,In_372);
nor U3415 (N_3415,In_859,In_1623);
nand U3416 (N_3416,In_587,In_569);
nand U3417 (N_3417,In_1546,In_447);
or U3418 (N_3418,In_138,In_688);
or U3419 (N_3419,In_1519,In_418);
and U3420 (N_3420,In_520,In_346);
nand U3421 (N_3421,In_188,In_94);
and U3422 (N_3422,In_637,In_1576);
or U3423 (N_3423,In_1489,In_1977);
xnor U3424 (N_3424,In_1558,In_1417);
or U3425 (N_3425,In_1628,In_341);
or U3426 (N_3426,In_8,In_1002);
nor U3427 (N_3427,In_625,In_655);
or U3428 (N_3428,In_1834,In_223);
nand U3429 (N_3429,In_1385,In_549);
nor U3430 (N_3430,In_610,In_1113);
or U3431 (N_3431,In_1731,In_1393);
nor U3432 (N_3432,In_810,In_595);
xnor U3433 (N_3433,In_183,In_1045);
nor U3434 (N_3434,In_1953,In_205);
or U3435 (N_3435,In_42,In_1165);
or U3436 (N_3436,In_1876,In_751);
and U3437 (N_3437,In_162,In_979);
nand U3438 (N_3438,In_1260,In_1760);
and U3439 (N_3439,In_1559,In_1362);
or U3440 (N_3440,In_1630,In_1600);
nand U3441 (N_3441,In_5,In_1226);
and U3442 (N_3442,In_95,In_952);
and U3443 (N_3443,In_1581,In_1164);
xnor U3444 (N_3444,In_17,In_1263);
or U3445 (N_3445,In_984,In_1582);
and U3446 (N_3446,In_1500,In_123);
and U3447 (N_3447,In_781,In_1094);
or U3448 (N_3448,In_132,In_125);
or U3449 (N_3449,In_1980,In_1597);
nor U3450 (N_3450,In_1753,In_1850);
and U3451 (N_3451,In_1352,In_1738);
and U3452 (N_3452,In_322,In_471);
nand U3453 (N_3453,In_402,In_1189);
or U3454 (N_3454,In_965,In_1173);
nor U3455 (N_3455,In_1417,In_645);
and U3456 (N_3456,In_89,In_996);
or U3457 (N_3457,In_338,In_1778);
nor U3458 (N_3458,In_1375,In_592);
xor U3459 (N_3459,In_1975,In_1822);
or U3460 (N_3460,In_1865,In_1988);
and U3461 (N_3461,In_172,In_1017);
nor U3462 (N_3462,In_352,In_1615);
and U3463 (N_3463,In_451,In_1237);
or U3464 (N_3464,In_1100,In_1209);
or U3465 (N_3465,In_354,In_1103);
or U3466 (N_3466,In_1173,In_252);
and U3467 (N_3467,In_209,In_268);
or U3468 (N_3468,In_1237,In_1212);
nor U3469 (N_3469,In_273,In_881);
and U3470 (N_3470,In_625,In_7);
or U3471 (N_3471,In_971,In_230);
nand U3472 (N_3472,In_1855,In_1961);
nor U3473 (N_3473,In_1469,In_1615);
and U3474 (N_3474,In_1509,In_1050);
nor U3475 (N_3475,In_680,In_795);
nand U3476 (N_3476,In_990,In_328);
nor U3477 (N_3477,In_1256,In_1436);
nor U3478 (N_3478,In_1127,In_1190);
and U3479 (N_3479,In_383,In_1378);
nand U3480 (N_3480,In_1492,In_905);
nand U3481 (N_3481,In_295,In_1178);
and U3482 (N_3482,In_473,In_739);
nor U3483 (N_3483,In_1283,In_601);
nor U3484 (N_3484,In_1247,In_1406);
and U3485 (N_3485,In_1056,In_1334);
nor U3486 (N_3486,In_1606,In_114);
or U3487 (N_3487,In_1934,In_426);
nand U3488 (N_3488,In_313,In_1840);
and U3489 (N_3489,In_656,In_1994);
nand U3490 (N_3490,In_939,In_633);
and U3491 (N_3491,In_311,In_511);
or U3492 (N_3492,In_1901,In_1653);
nor U3493 (N_3493,In_342,In_60);
or U3494 (N_3494,In_1563,In_1040);
xnor U3495 (N_3495,In_493,In_1965);
nand U3496 (N_3496,In_1220,In_1121);
or U3497 (N_3497,In_68,In_1069);
xnor U3498 (N_3498,In_280,In_1600);
or U3499 (N_3499,In_763,In_443);
nor U3500 (N_3500,In_952,In_1956);
nand U3501 (N_3501,In_433,In_1982);
and U3502 (N_3502,In_162,In_408);
and U3503 (N_3503,In_387,In_18);
nand U3504 (N_3504,In_1722,In_1727);
and U3505 (N_3505,In_1437,In_88);
or U3506 (N_3506,In_175,In_954);
xnor U3507 (N_3507,In_255,In_739);
nor U3508 (N_3508,In_992,In_272);
nor U3509 (N_3509,In_1688,In_931);
nor U3510 (N_3510,In_1092,In_550);
or U3511 (N_3511,In_938,In_1128);
or U3512 (N_3512,In_1649,In_957);
nand U3513 (N_3513,In_1619,In_882);
and U3514 (N_3514,In_76,In_623);
and U3515 (N_3515,In_1817,In_137);
nor U3516 (N_3516,In_917,In_1294);
nor U3517 (N_3517,In_1845,In_1681);
nor U3518 (N_3518,In_1278,In_1036);
nor U3519 (N_3519,In_70,In_257);
and U3520 (N_3520,In_1263,In_1517);
xor U3521 (N_3521,In_1551,In_1359);
and U3522 (N_3522,In_1740,In_1031);
and U3523 (N_3523,In_57,In_1250);
and U3524 (N_3524,In_1497,In_1520);
nor U3525 (N_3525,In_692,In_1425);
nand U3526 (N_3526,In_373,In_1115);
and U3527 (N_3527,In_1190,In_9);
nand U3528 (N_3528,In_1147,In_463);
nand U3529 (N_3529,In_1600,In_732);
nor U3530 (N_3530,In_441,In_303);
nor U3531 (N_3531,In_1924,In_1369);
nand U3532 (N_3532,In_2,In_917);
or U3533 (N_3533,In_971,In_650);
nand U3534 (N_3534,In_55,In_831);
nor U3535 (N_3535,In_799,In_1265);
nor U3536 (N_3536,In_756,In_1723);
and U3537 (N_3537,In_329,In_1507);
and U3538 (N_3538,In_397,In_1790);
nand U3539 (N_3539,In_219,In_431);
or U3540 (N_3540,In_1326,In_988);
nor U3541 (N_3541,In_1493,In_1293);
or U3542 (N_3542,In_1285,In_115);
or U3543 (N_3543,In_707,In_1777);
nor U3544 (N_3544,In_1673,In_480);
or U3545 (N_3545,In_956,In_878);
and U3546 (N_3546,In_1415,In_427);
xor U3547 (N_3547,In_1341,In_1429);
and U3548 (N_3548,In_379,In_1883);
nand U3549 (N_3549,In_1973,In_1861);
xor U3550 (N_3550,In_751,In_89);
and U3551 (N_3551,In_145,In_55);
and U3552 (N_3552,In_368,In_1784);
or U3553 (N_3553,In_982,In_1102);
or U3554 (N_3554,In_1620,In_1452);
and U3555 (N_3555,In_700,In_537);
and U3556 (N_3556,In_1193,In_1488);
nor U3557 (N_3557,In_1605,In_841);
and U3558 (N_3558,In_1537,In_172);
and U3559 (N_3559,In_684,In_354);
nor U3560 (N_3560,In_1243,In_1694);
nand U3561 (N_3561,In_594,In_1104);
xor U3562 (N_3562,In_177,In_363);
nand U3563 (N_3563,In_455,In_410);
nand U3564 (N_3564,In_966,In_669);
nor U3565 (N_3565,In_1235,In_241);
and U3566 (N_3566,In_1657,In_1083);
nand U3567 (N_3567,In_1039,In_1970);
nand U3568 (N_3568,In_1087,In_1120);
and U3569 (N_3569,In_345,In_1705);
nor U3570 (N_3570,In_1253,In_1222);
nor U3571 (N_3571,In_1595,In_270);
and U3572 (N_3572,In_1359,In_763);
and U3573 (N_3573,In_1140,In_493);
xor U3574 (N_3574,In_47,In_1935);
and U3575 (N_3575,In_507,In_1212);
nor U3576 (N_3576,In_931,In_1058);
or U3577 (N_3577,In_195,In_352);
nand U3578 (N_3578,In_710,In_551);
or U3579 (N_3579,In_1877,In_1131);
nor U3580 (N_3580,In_754,In_793);
xnor U3581 (N_3581,In_1368,In_1311);
nand U3582 (N_3582,In_1223,In_428);
and U3583 (N_3583,In_1077,In_335);
nor U3584 (N_3584,In_1487,In_964);
nand U3585 (N_3585,In_1930,In_1781);
nor U3586 (N_3586,In_1407,In_1554);
and U3587 (N_3587,In_410,In_530);
nand U3588 (N_3588,In_921,In_485);
nor U3589 (N_3589,In_1425,In_665);
or U3590 (N_3590,In_423,In_1241);
or U3591 (N_3591,In_156,In_402);
nand U3592 (N_3592,In_1856,In_1069);
xnor U3593 (N_3593,In_1451,In_382);
and U3594 (N_3594,In_345,In_58);
nor U3595 (N_3595,In_1063,In_1035);
nor U3596 (N_3596,In_544,In_854);
nand U3597 (N_3597,In_1958,In_705);
xor U3598 (N_3598,In_547,In_1822);
nand U3599 (N_3599,In_1714,In_1456);
nand U3600 (N_3600,In_385,In_1036);
nor U3601 (N_3601,In_497,In_126);
or U3602 (N_3602,In_266,In_527);
or U3603 (N_3603,In_605,In_1177);
and U3604 (N_3604,In_649,In_338);
nor U3605 (N_3605,In_719,In_959);
and U3606 (N_3606,In_1292,In_973);
nor U3607 (N_3607,In_1453,In_1894);
and U3608 (N_3608,In_285,In_215);
xnor U3609 (N_3609,In_1998,In_296);
nand U3610 (N_3610,In_164,In_602);
nand U3611 (N_3611,In_605,In_1781);
nand U3612 (N_3612,In_263,In_1959);
and U3613 (N_3613,In_1001,In_1100);
nand U3614 (N_3614,In_948,In_1798);
and U3615 (N_3615,In_1775,In_893);
xor U3616 (N_3616,In_538,In_571);
nand U3617 (N_3617,In_284,In_90);
and U3618 (N_3618,In_68,In_636);
nand U3619 (N_3619,In_1474,In_495);
nand U3620 (N_3620,In_953,In_568);
nand U3621 (N_3621,In_904,In_859);
or U3622 (N_3622,In_1697,In_522);
nor U3623 (N_3623,In_445,In_1776);
or U3624 (N_3624,In_1482,In_1488);
or U3625 (N_3625,In_1389,In_1242);
or U3626 (N_3626,In_1436,In_1173);
nand U3627 (N_3627,In_1940,In_1888);
and U3628 (N_3628,In_1278,In_541);
and U3629 (N_3629,In_762,In_1573);
or U3630 (N_3630,In_1588,In_1798);
xor U3631 (N_3631,In_1409,In_1071);
nor U3632 (N_3632,In_1566,In_175);
and U3633 (N_3633,In_1227,In_1895);
nor U3634 (N_3634,In_1235,In_943);
nand U3635 (N_3635,In_1291,In_819);
nand U3636 (N_3636,In_197,In_918);
or U3637 (N_3637,In_114,In_733);
nor U3638 (N_3638,In_167,In_4);
and U3639 (N_3639,In_1273,In_1668);
xor U3640 (N_3640,In_328,In_933);
nor U3641 (N_3641,In_647,In_252);
or U3642 (N_3642,In_217,In_103);
xnor U3643 (N_3643,In_1427,In_1774);
xor U3644 (N_3644,In_228,In_488);
nand U3645 (N_3645,In_772,In_1818);
or U3646 (N_3646,In_1140,In_1076);
nor U3647 (N_3647,In_597,In_493);
xor U3648 (N_3648,In_61,In_1248);
nand U3649 (N_3649,In_1259,In_168);
nor U3650 (N_3650,In_169,In_634);
and U3651 (N_3651,In_884,In_1418);
and U3652 (N_3652,In_1800,In_1091);
nor U3653 (N_3653,In_1593,In_1664);
nor U3654 (N_3654,In_448,In_973);
or U3655 (N_3655,In_1385,In_1991);
nand U3656 (N_3656,In_131,In_301);
or U3657 (N_3657,In_31,In_443);
nand U3658 (N_3658,In_137,In_1442);
and U3659 (N_3659,In_1613,In_591);
and U3660 (N_3660,In_221,In_864);
or U3661 (N_3661,In_1849,In_1139);
nor U3662 (N_3662,In_409,In_869);
and U3663 (N_3663,In_1658,In_1369);
nand U3664 (N_3664,In_1082,In_669);
nand U3665 (N_3665,In_1297,In_1992);
and U3666 (N_3666,In_1314,In_1928);
nor U3667 (N_3667,In_587,In_1530);
nor U3668 (N_3668,In_1039,In_1124);
and U3669 (N_3669,In_1074,In_1241);
nand U3670 (N_3670,In_866,In_1497);
xnor U3671 (N_3671,In_1187,In_459);
nand U3672 (N_3672,In_472,In_513);
nand U3673 (N_3673,In_1543,In_1801);
nor U3674 (N_3674,In_1193,In_1833);
nand U3675 (N_3675,In_636,In_1716);
nand U3676 (N_3676,In_1592,In_1354);
and U3677 (N_3677,In_1000,In_1115);
xnor U3678 (N_3678,In_1860,In_219);
nand U3679 (N_3679,In_1034,In_554);
xor U3680 (N_3680,In_884,In_47);
nand U3681 (N_3681,In_472,In_401);
xor U3682 (N_3682,In_1529,In_76);
and U3683 (N_3683,In_848,In_365);
nor U3684 (N_3684,In_876,In_1009);
or U3685 (N_3685,In_1294,In_1997);
nand U3686 (N_3686,In_1107,In_490);
or U3687 (N_3687,In_1585,In_299);
or U3688 (N_3688,In_1708,In_638);
nor U3689 (N_3689,In_1062,In_83);
and U3690 (N_3690,In_602,In_790);
or U3691 (N_3691,In_1030,In_1709);
and U3692 (N_3692,In_947,In_192);
nor U3693 (N_3693,In_815,In_375);
nand U3694 (N_3694,In_224,In_1484);
xor U3695 (N_3695,In_559,In_417);
and U3696 (N_3696,In_541,In_173);
nor U3697 (N_3697,In_334,In_1150);
xor U3698 (N_3698,In_1545,In_1319);
or U3699 (N_3699,In_311,In_419);
or U3700 (N_3700,In_1292,In_55);
or U3701 (N_3701,In_1888,In_1272);
or U3702 (N_3702,In_674,In_1443);
nor U3703 (N_3703,In_502,In_29);
nor U3704 (N_3704,In_1656,In_1061);
nand U3705 (N_3705,In_1237,In_1997);
and U3706 (N_3706,In_655,In_1021);
and U3707 (N_3707,In_428,In_1381);
nand U3708 (N_3708,In_1664,In_292);
xnor U3709 (N_3709,In_1878,In_1314);
or U3710 (N_3710,In_983,In_1275);
nor U3711 (N_3711,In_162,In_1319);
or U3712 (N_3712,In_277,In_1140);
nand U3713 (N_3713,In_1642,In_658);
or U3714 (N_3714,In_316,In_1430);
nand U3715 (N_3715,In_332,In_466);
xnor U3716 (N_3716,In_1028,In_423);
or U3717 (N_3717,In_609,In_499);
or U3718 (N_3718,In_1215,In_632);
and U3719 (N_3719,In_1565,In_1056);
xnor U3720 (N_3720,In_427,In_1389);
or U3721 (N_3721,In_1224,In_392);
or U3722 (N_3722,In_252,In_1877);
or U3723 (N_3723,In_1710,In_1123);
xnor U3724 (N_3724,In_553,In_1732);
or U3725 (N_3725,In_1734,In_489);
and U3726 (N_3726,In_293,In_424);
and U3727 (N_3727,In_429,In_1038);
xor U3728 (N_3728,In_1955,In_1219);
or U3729 (N_3729,In_1239,In_1524);
nor U3730 (N_3730,In_1624,In_849);
nor U3731 (N_3731,In_1330,In_1404);
nand U3732 (N_3732,In_1409,In_642);
nor U3733 (N_3733,In_239,In_1246);
nor U3734 (N_3734,In_991,In_1806);
and U3735 (N_3735,In_1875,In_1887);
nand U3736 (N_3736,In_970,In_956);
nand U3737 (N_3737,In_1345,In_1581);
or U3738 (N_3738,In_1021,In_651);
nor U3739 (N_3739,In_909,In_730);
nor U3740 (N_3740,In_63,In_1372);
nor U3741 (N_3741,In_1929,In_572);
or U3742 (N_3742,In_1820,In_1697);
nand U3743 (N_3743,In_723,In_1105);
nor U3744 (N_3744,In_339,In_1352);
and U3745 (N_3745,In_1701,In_1214);
or U3746 (N_3746,In_1315,In_1327);
or U3747 (N_3747,In_1053,In_956);
nand U3748 (N_3748,In_1656,In_1712);
and U3749 (N_3749,In_997,In_1454);
nor U3750 (N_3750,In_566,In_698);
nand U3751 (N_3751,In_1661,In_426);
nor U3752 (N_3752,In_71,In_1543);
nand U3753 (N_3753,In_1954,In_911);
nor U3754 (N_3754,In_1640,In_1525);
and U3755 (N_3755,In_571,In_805);
and U3756 (N_3756,In_823,In_9);
nand U3757 (N_3757,In_1696,In_1644);
or U3758 (N_3758,In_1774,In_913);
and U3759 (N_3759,In_105,In_1961);
and U3760 (N_3760,In_357,In_1932);
nor U3761 (N_3761,In_634,In_1065);
and U3762 (N_3762,In_419,In_1474);
or U3763 (N_3763,In_299,In_653);
or U3764 (N_3764,In_1286,In_1202);
nor U3765 (N_3765,In_33,In_1665);
and U3766 (N_3766,In_847,In_366);
nor U3767 (N_3767,In_976,In_675);
nand U3768 (N_3768,In_949,In_655);
nor U3769 (N_3769,In_1111,In_328);
xnor U3770 (N_3770,In_1740,In_485);
nand U3771 (N_3771,In_0,In_1994);
nor U3772 (N_3772,In_1683,In_1928);
nor U3773 (N_3773,In_763,In_836);
nor U3774 (N_3774,In_1736,In_997);
and U3775 (N_3775,In_1786,In_220);
and U3776 (N_3776,In_1598,In_692);
or U3777 (N_3777,In_465,In_97);
nor U3778 (N_3778,In_200,In_1097);
nand U3779 (N_3779,In_766,In_66);
and U3780 (N_3780,In_1132,In_81);
and U3781 (N_3781,In_1640,In_552);
nor U3782 (N_3782,In_797,In_67);
or U3783 (N_3783,In_1889,In_104);
xor U3784 (N_3784,In_918,In_206);
xor U3785 (N_3785,In_1781,In_1134);
or U3786 (N_3786,In_1310,In_718);
nor U3787 (N_3787,In_516,In_1968);
and U3788 (N_3788,In_1802,In_1573);
and U3789 (N_3789,In_787,In_128);
or U3790 (N_3790,In_1376,In_156);
or U3791 (N_3791,In_1591,In_813);
and U3792 (N_3792,In_1519,In_75);
nor U3793 (N_3793,In_1358,In_426);
xor U3794 (N_3794,In_1345,In_1489);
or U3795 (N_3795,In_500,In_1991);
or U3796 (N_3796,In_19,In_513);
nor U3797 (N_3797,In_631,In_1592);
and U3798 (N_3798,In_559,In_346);
or U3799 (N_3799,In_908,In_1332);
nor U3800 (N_3800,In_709,In_240);
and U3801 (N_3801,In_860,In_1753);
or U3802 (N_3802,In_975,In_911);
nor U3803 (N_3803,In_1631,In_1613);
and U3804 (N_3804,In_1507,In_1443);
nor U3805 (N_3805,In_1328,In_270);
nor U3806 (N_3806,In_1338,In_1001);
or U3807 (N_3807,In_683,In_126);
xnor U3808 (N_3808,In_45,In_22);
or U3809 (N_3809,In_921,In_1244);
nand U3810 (N_3810,In_1187,In_563);
nand U3811 (N_3811,In_842,In_1603);
or U3812 (N_3812,In_1588,In_930);
and U3813 (N_3813,In_3,In_1507);
nor U3814 (N_3814,In_1896,In_1065);
and U3815 (N_3815,In_1280,In_690);
xor U3816 (N_3816,In_12,In_1446);
nand U3817 (N_3817,In_1823,In_731);
xor U3818 (N_3818,In_908,In_1006);
nand U3819 (N_3819,In_251,In_261);
nand U3820 (N_3820,In_235,In_917);
and U3821 (N_3821,In_1286,In_702);
nand U3822 (N_3822,In_993,In_1413);
and U3823 (N_3823,In_802,In_640);
or U3824 (N_3824,In_135,In_795);
and U3825 (N_3825,In_1960,In_1125);
nor U3826 (N_3826,In_1437,In_902);
nor U3827 (N_3827,In_1732,In_1006);
and U3828 (N_3828,In_755,In_599);
nor U3829 (N_3829,In_1040,In_1355);
nand U3830 (N_3830,In_1902,In_513);
or U3831 (N_3831,In_375,In_1274);
nand U3832 (N_3832,In_948,In_1476);
and U3833 (N_3833,In_1466,In_1663);
or U3834 (N_3834,In_629,In_768);
xnor U3835 (N_3835,In_1316,In_483);
nor U3836 (N_3836,In_1726,In_1799);
and U3837 (N_3837,In_1981,In_71);
nor U3838 (N_3838,In_88,In_537);
or U3839 (N_3839,In_478,In_746);
nor U3840 (N_3840,In_7,In_683);
nor U3841 (N_3841,In_297,In_740);
or U3842 (N_3842,In_1621,In_902);
nand U3843 (N_3843,In_469,In_1158);
and U3844 (N_3844,In_1260,In_1814);
nand U3845 (N_3845,In_1203,In_1958);
nor U3846 (N_3846,In_1913,In_1361);
and U3847 (N_3847,In_419,In_986);
and U3848 (N_3848,In_841,In_1042);
or U3849 (N_3849,In_1815,In_1228);
nand U3850 (N_3850,In_1045,In_1682);
nand U3851 (N_3851,In_1697,In_692);
nor U3852 (N_3852,In_1919,In_272);
and U3853 (N_3853,In_440,In_1859);
and U3854 (N_3854,In_1899,In_1613);
and U3855 (N_3855,In_831,In_1230);
xnor U3856 (N_3856,In_1754,In_491);
nand U3857 (N_3857,In_192,In_1722);
nor U3858 (N_3858,In_778,In_1858);
xor U3859 (N_3859,In_436,In_685);
or U3860 (N_3860,In_958,In_412);
nand U3861 (N_3861,In_261,In_1015);
nor U3862 (N_3862,In_119,In_528);
nor U3863 (N_3863,In_277,In_1178);
nand U3864 (N_3864,In_1476,In_712);
nor U3865 (N_3865,In_1341,In_305);
and U3866 (N_3866,In_1194,In_894);
or U3867 (N_3867,In_579,In_891);
nor U3868 (N_3868,In_555,In_383);
nand U3869 (N_3869,In_1894,In_617);
or U3870 (N_3870,In_308,In_728);
nand U3871 (N_3871,In_1352,In_393);
xnor U3872 (N_3872,In_798,In_982);
or U3873 (N_3873,In_897,In_1582);
nand U3874 (N_3874,In_1990,In_398);
or U3875 (N_3875,In_1365,In_1351);
or U3876 (N_3876,In_1905,In_1184);
and U3877 (N_3877,In_1428,In_641);
nand U3878 (N_3878,In_1336,In_1530);
or U3879 (N_3879,In_1334,In_1038);
nand U3880 (N_3880,In_1157,In_1353);
nor U3881 (N_3881,In_1657,In_609);
nand U3882 (N_3882,In_693,In_506);
nand U3883 (N_3883,In_1669,In_1919);
nand U3884 (N_3884,In_679,In_362);
or U3885 (N_3885,In_459,In_377);
and U3886 (N_3886,In_1065,In_329);
nor U3887 (N_3887,In_1529,In_1807);
nor U3888 (N_3888,In_18,In_728);
nor U3889 (N_3889,In_879,In_958);
or U3890 (N_3890,In_1455,In_757);
or U3891 (N_3891,In_529,In_1098);
and U3892 (N_3892,In_1593,In_1794);
nand U3893 (N_3893,In_1675,In_1582);
and U3894 (N_3894,In_512,In_1002);
nor U3895 (N_3895,In_886,In_709);
or U3896 (N_3896,In_717,In_550);
or U3897 (N_3897,In_170,In_1272);
nor U3898 (N_3898,In_706,In_996);
nor U3899 (N_3899,In_1482,In_399);
and U3900 (N_3900,In_947,In_485);
or U3901 (N_3901,In_1416,In_101);
nor U3902 (N_3902,In_344,In_368);
nand U3903 (N_3903,In_245,In_1839);
or U3904 (N_3904,In_1078,In_1650);
nand U3905 (N_3905,In_212,In_1168);
nor U3906 (N_3906,In_1046,In_1431);
or U3907 (N_3907,In_1131,In_765);
and U3908 (N_3908,In_1133,In_83);
and U3909 (N_3909,In_199,In_1465);
nand U3910 (N_3910,In_1120,In_263);
and U3911 (N_3911,In_1022,In_1286);
nand U3912 (N_3912,In_1130,In_590);
nand U3913 (N_3913,In_1665,In_290);
nand U3914 (N_3914,In_368,In_1534);
nand U3915 (N_3915,In_1372,In_832);
xnor U3916 (N_3916,In_53,In_343);
nand U3917 (N_3917,In_674,In_558);
or U3918 (N_3918,In_1809,In_1952);
nor U3919 (N_3919,In_1071,In_713);
xor U3920 (N_3920,In_1238,In_1893);
or U3921 (N_3921,In_1736,In_1172);
and U3922 (N_3922,In_1116,In_1243);
and U3923 (N_3923,In_1519,In_1789);
or U3924 (N_3924,In_1876,In_1974);
nor U3925 (N_3925,In_1614,In_15);
and U3926 (N_3926,In_1567,In_587);
nor U3927 (N_3927,In_1234,In_1469);
xor U3928 (N_3928,In_1908,In_931);
nor U3929 (N_3929,In_1248,In_1296);
and U3930 (N_3930,In_1860,In_1757);
nand U3931 (N_3931,In_1935,In_96);
nand U3932 (N_3932,In_307,In_1453);
nor U3933 (N_3933,In_1681,In_902);
or U3934 (N_3934,In_417,In_1818);
and U3935 (N_3935,In_160,In_1823);
nor U3936 (N_3936,In_1893,In_1627);
nand U3937 (N_3937,In_1907,In_237);
nand U3938 (N_3938,In_1451,In_455);
and U3939 (N_3939,In_1995,In_139);
nand U3940 (N_3940,In_209,In_47);
nand U3941 (N_3941,In_522,In_830);
nand U3942 (N_3942,In_841,In_198);
nor U3943 (N_3943,In_775,In_1217);
xor U3944 (N_3944,In_335,In_368);
or U3945 (N_3945,In_281,In_1789);
nand U3946 (N_3946,In_575,In_810);
nand U3947 (N_3947,In_1448,In_1080);
and U3948 (N_3948,In_450,In_1876);
and U3949 (N_3949,In_1655,In_79);
or U3950 (N_3950,In_508,In_1829);
nor U3951 (N_3951,In_617,In_736);
nor U3952 (N_3952,In_1909,In_646);
nor U3953 (N_3953,In_426,In_752);
nand U3954 (N_3954,In_1469,In_1637);
and U3955 (N_3955,In_1982,In_916);
and U3956 (N_3956,In_385,In_112);
and U3957 (N_3957,In_1022,In_1824);
nor U3958 (N_3958,In_1747,In_955);
nor U3959 (N_3959,In_1408,In_997);
or U3960 (N_3960,In_1206,In_1793);
or U3961 (N_3961,In_53,In_1311);
or U3962 (N_3962,In_1191,In_1886);
or U3963 (N_3963,In_755,In_357);
xor U3964 (N_3964,In_1383,In_473);
nand U3965 (N_3965,In_1975,In_1790);
or U3966 (N_3966,In_1787,In_658);
nor U3967 (N_3967,In_970,In_896);
nand U3968 (N_3968,In_457,In_517);
nand U3969 (N_3969,In_1161,In_710);
xor U3970 (N_3970,In_290,In_1074);
nor U3971 (N_3971,In_859,In_1315);
or U3972 (N_3972,In_457,In_173);
or U3973 (N_3973,In_877,In_1810);
and U3974 (N_3974,In_1602,In_1769);
nor U3975 (N_3975,In_17,In_402);
nor U3976 (N_3976,In_713,In_355);
or U3977 (N_3977,In_1764,In_65);
and U3978 (N_3978,In_353,In_1248);
nand U3979 (N_3979,In_32,In_847);
nor U3980 (N_3980,In_1430,In_1912);
nor U3981 (N_3981,In_1902,In_1752);
nor U3982 (N_3982,In_1771,In_307);
nand U3983 (N_3983,In_506,In_346);
nor U3984 (N_3984,In_1257,In_652);
nand U3985 (N_3985,In_27,In_1661);
nor U3986 (N_3986,In_1619,In_1798);
nor U3987 (N_3987,In_1732,In_63);
or U3988 (N_3988,In_1451,In_1685);
nand U3989 (N_3989,In_1455,In_926);
and U3990 (N_3990,In_1114,In_118);
nand U3991 (N_3991,In_819,In_1939);
and U3992 (N_3992,In_813,In_340);
or U3993 (N_3993,In_1011,In_656);
or U3994 (N_3994,In_863,In_526);
nand U3995 (N_3995,In_1498,In_1639);
and U3996 (N_3996,In_1129,In_1956);
or U3997 (N_3997,In_1556,In_508);
nand U3998 (N_3998,In_57,In_990);
and U3999 (N_3999,In_1828,In_1986);
and U4000 (N_4000,In_1291,In_922);
or U4001 (N_4001,In_472,In_678);
nor U4002 (N_4002,In_1304,In_775);
nor U4003 (N_4003,In_553,In_1334);
nor U4004 (N_4004,In_434,In_659);
nor U4005 (N_4005,In_1336,In_1875);
nand U4006 (N_4006,In_453,In_1547);
and U4007 (N_4007,In_1516,In_1461);
xor U4008 (N_4008,In_686,In_1334);
or U4009 (N_4009,In_1435,In_954);
or U4010 (N_4010,In_1545,In_1485);
nor U4011 (N_4011,In_598,In_57);
nand U4012 (N_4012,In_137,In_210);
nor U4013 (N_4013,In_1155,In_1834);
or U4014 (N_4014,In_1086,In_1521);
xor U4015 (N_4015,In_1545,In_1312);
nor U4016 (N_4016,In_1166,In_1367);
or U4017 (N_4017,In_1705,In_552);
nand U4018 (N_4018,In_1623,In_596);
nor U4019 (N_4019,In_155,In_1278);
nor U4020 (N_4020,In_83,In_1763);
or U4021 (N_4021,In_1864,In_709);
nor U4022 (N_4022,In_832,In_1122);
nor U4023 (N_4023,In_829,In_1273);
nand U4024 (N_4024,In_1717,In_580);
or U4025 (N_4025,In_684,In_1167);
xor U4026 (N_4026,In_124,In_1155);
nand U4027 (N_4027,In_1713,In_974);
nand U4028 (N_4028,In_1344,In_179);
xor U4029 (N_4029,In_413,In_827);
nand U4030 (N_4030,In_667,In_1309);
or U4031 (N_4031,In_650,In_618);
nor U4032 (N_4032,In_183,In_220);
xor U4033 (N_4033,In_1496,In_1030);
or U4034 (N_4034,In_669,In_13);
or U4035 (N_4035,In_246,In_1485);
or U4036 (N_4036,In_621,In_1970);
and U4037 (N_4037,In_774,In_404);
nor U4038 (N_4038,In_179,In_735);
and U4039 (N_4039,In_1282,In_148);
or U4040 (N_4040,In_1584,In_210);
or U4041 (N_4041,In_168,In_1419);
or U4042 (N_4042,In_644,In_1014);
nor U4043 (N_4043,In_1895,In_834);
nand U4044 (N_4044,In_1899,In_868);
nor U4045 (N_4045,In_736,In_1145);
nand U4046 (N_4046,In_1050,In_1186);
nand U4047 (N_4047,In_1019,In_1321);
and U4048 (N_4048,In_1662,In_1107);
nand U4049 (N_4049,In_230,In_705);
and U4050 (N_4050,In_925,In_1344);
nand U4051 (N_4051,In_1854,In_657);
or U4052 (N_4052,In_788,In_1992);
nand U4053 (N_4053,In_523,In_351);
nand U4054 (N_4054,In_124,In_1998);
and U4055 (N_4055,In_1774,In_399);
and U4056 (N_4056,In_1922,In_855);
xnor U4057 (N_4057,In_1966,In_218);
and U4058 (N_4058,In_1602,In_695);
and U4059 (N_4059,In_859,In_848);
or U4060 (N_4060,In_123,In_301);
nand U4061 (N_4061,In_1142,In_1659);
nand U4062 (N_4062,In_937,In_1452);
and U4063 (N_4063,In_412,In_688);
nor U4064 (N_4064,In_1291,In_984);
xor U4065 (N_4065,In_1436,In_1158);
nor U4066 (N_4066,In_977,In_205);
or U4067 (N_4067,In_1122,In_1176);
nand U4068 (N_4068,In_1971,In_1683);
and U4069 (N_4069,In_1734,In_1011);
and U4070 (N_4070,In_1310,In_1241);
or U4071 (N_4071,In_755,In_1455);
xor U4072 (N_4072,In_1847,In_1769);
nor U4073 (N_4073,In_585,In_1276);
nor U4074 (N_4074,In_554,In_1769);
and U4075 (N_4075,In_1398,In_1578);
and U4076 (N_4076,In_1221,In_69);
and U4077 (N_4077,In_1624,In_1673);
nand U4078 (N_4078,In_706,In_1244);
xnor U4079 (N_4079,In_1931,In_1222);
and U4080 (N_4080,In_475,In_388);
xor U4081 (N_4081,In_234,In_1623);
or U4082 (N_4082,In_1468,In_1532);
nand U4083 (N_4083,In_1071,In_920);
nor U4084 (N_4084,In_726,In_857);
and U4085 (N_4085,In_162,In_1107);
nor U4086 (N_4086,In_1038,In_42);
or U4087 (N_4087,In_1601,In_1045);
or U4088 (N_4088,In_1329,In_530);
and U4089 (N_4089,In_692,In_528);
and U4090 (N_4090,In_1694,In_901);
xnor U4091 (N_4091,In_807,In_1874);
and U4092 (N_4092,In_1144,In_1007);
nand U4093 (N_4093,In_1937,In_1575);
and U4094 (N_4094,In_1429,In_1960);
xnor U4095 (N_4095,In_1625,In_811);
and U4096 (N_4096,In_825,In_232);
xnor U4097 (N_4097,In_528,In_1915);
xnor U4098 (N_4098,In_1365,In_1820);
and U4099 (N_4099,In_1587,In_234);
or U4100 (N_4100,In_766,In_108);
and U4101 (N_4101,In_889,In_679);
xnor U4102 (N_4102,In_290,In_512);
or U4103 (N_4103,In_549,In_1662);
nor U4104 (N_4104,In_253,In_1188);
xor U4105 (N_4105,In_944,In_462);
or U4106 (N_4106,In_825,In_400);
nor U4107 (N_4107,In_500,In_1223);
nor U4108 (N_4108,In_195,In_32);
or U4109 (N_4109,In_62,In_1567);
nand U4110 (N_4110,In_177,In_521);
and U4111 (N_4111,In_986,In_522);
or U4112 (N_4112,In_41,In_639);
and U4113 (N_4113,In_474,In_508);
and U4114 (N_4114,In_966,In_1264);
nand U4115 (N_4115,In_58,In_919);
nor U4116 (N_4116,In_413,In_1579);
nand U4117 (N_4117,In_771,In_1521);
nor U4118 (N_4118,In_1916,In_1512);
nor U4119 (N_4119,In_220,In_1644);
xnor U4120 (N_4120,In_565,In_167);
nand U4121 (N_4121,In_976,In_1169);
or U4122 (N_4122,In_1260,In_1985);
and U4123 (N_4123,In_325,In_911);
nor U4124 (N_4124,In_1789,In_1954);
xnor U4125 (N_4125,In_1697,In_1288);
and U4126 (N_4126,In_108,In_1435);
nand U4127 (N_4127,In_918,In_1779);
and U4128 (N_4128,In_744,In_1233);
nand U4129 (N_4129,In_135,In_92);
or U4130 (N_4130,In_1658,In_250);
or U4131 (N_4131,In_1797,In_813);
xnor U4132 (N_4132,In_467,In_579);
and U4133 (N_4133,In_1971,In_279);
xnor U4134 (N_4134,In_1377,In_77);
and U4135 (N_4135,In_572,In_732);
nor U4136 (N_4136,In_910,In_1727);
nor U4137 (N_4137,In_1970,In_1673);
or U4138 (N_4138,In_1634,In_1451);
and U4139 (N_4139,In_1092,In_1944);
or U4140 (N_4140,In_336,In_1479);
or U4141 (N_4141,In_1614,In_167);
nand U4142 (N_4142,In_1139,In_1877);
or U4143 (N_4143,In_1671,In_1847);
nand U4144 (N_4144,In_914,In_1031);
nor U4145 (N_4145,In_59,In_825);
or U4146 (N_4146,In_1203,In_602);
nand U4147 (N_4147,In_1623,In_1995);
nand U4148 (N_4148,In_841,In_861);
xnor U4149 (N_4149,In_386,In_100);
and U4150 (N_4150,In_1017,In_1827);
and U4151 (N_4151,In_1446,In_1093);
xor U4152 (N_4152,In_135,In_965);
nand U4153 (N_4153,In_1190,In_1517);
or U4154 (N_4154,In_1326,In_1632);
nand U4155 (N_4155,In_1370,In_1649);
nand U4156 (N_4156,In_820,In_76);
nor U4157 (N_4157,In_1908,In_674);
nand U4158 (N_4158,In_1441,In_909);
nand U4159 (N_4159,In_914,In_1153);
nor U4160 (N_4160,In_1005,In_1274);
xnor U4161 (N_4161,In_174,In_541);
nand U4162 (N_4162,In_485,In_1829);
nand U4163 (N_4163,In_461,In_81);
nor U4164 (N_4164,In_1266,In_615);
nor U4165 (N_4165,In_770,In_663);
nand U4166 (N_4166,In_529,In_1379);
nand U4167 (N_4167,In_440,In_1714);
and U4168 (N_4168,In_1135,In_114);
xnor U4169 (N_4169,In_1846,In_347);
or U4170 (N_4170,In_882,In_832);
nor U4171 (N_4171,In_1742,In_1368);
and U4172 (N_4172,In_1572,In_1714);
and U4173 (N_4173,In_1772,In_1781);
and U4174 (N_4174,In_537,In_1500);
or U4175 (N_4175,In_1413,In_1902);
or U4176 (N_4176,In_1871,In_1218);
nand U4177 (N_4177,In_804,In_990);
xnor U4178 (N_4178,In_520,In_1913);
or U4179 (N_4179,In_1453,In_353);
or U4180 (N_4180,In_1883,In_1707);
nand U4181 (N_4181,In_44,In_1397);
nand U4182 (N_4182,In_1730,In_685);
and U4183 (N_4183,In_566,In_618);
nor U4184 (N_4184,In_1827,In_1328);
nor U4185 (N_4185,In_1161,In_183);
nor U4186 (N_4186,In_250,In_1088);
or U4187 (N_4187,In_60,In_189);
or U4188 (N_4188,In_4,In_1874);
and U4189 (N_4189,In_1859,In_619);
nor U4190 (N_4190,In_1148,In_1827);
and U4191 (N_4191,In_355,In_1724);
nand U4192 (N_4192,In_1939,In_623);
nor U4193 (N_4193,In_1384,In_849);
and U4194 (N_4194,In_206,In_484);
or U4195 (N_4195,In_644,In_1440);
or U4196 (N_4196,In_1467,In_1192);
or U4197 (N_4197,In_715,In_30);
nand U4198 (N_4198,In_377,In_1189);
or U4199 (N_4199,In_899,In_321);
nand U4200 (N_4200,In_57,In_1325);
nand U4201 (N_4201,In_1905,In_1792);
and U4202 (N_4202,In_511,In_1228);
nor U4203 (N_4203,In_177,In_1454);
nor U4204 (N_4204,In_1439,In_747);
xnor U4205 (N_4205,In_983,In_1707);
or U4206 (N_4206,In_66,In_44);
or U4207 (N_4207,In_1069,In_118);
nor U4208 (N_4208,In_1535,In_347);
nor U4209 (N_4209,In_1134,In_1867);
or U4210 (N_4210,In_1722,In_1702);
nor U4211 (N_4211,In_299,In_1558);
and U4212 (N_4212,In_1535,In_1269);
nand U4213 (N_4213,In_1436,In_34);
or U4214 (N_4214,In_197,In_667);
or U4215 (N_4215,In_1291,In_1375);
or U4216 (N_4216,In_1156,In_300);
nand U4217 (N_4217,In_1974,In_562);
nand U4218 (N_4218,In_743,In_1510);
nand U4219 (N_4219,In_1921,In_1569);
xnor U4220 (N_4220,In_985,In_805);
xor U4221 (N_4221,In_1874,In_1578);
nor U4222 (N_4222,In_1579,In_1402);
nand U4223 (N_4223,In_356,In_1428);
or U4224 (N_4224,In_671,In_728);
or U4225 (N_4225,In_1107,In_1807);
nor U4226 (N_4226,In_66,In_575);
and U4227 (N_4227,In_596,In_1496);
and U4228 (N_4228,In_1057,In_334);
nand U4229 (N_4229,In_1179,In_380);
and U4230 (N_4230,In_1882,In_483);
and U4231 (N_4231,In_503,In_3);
nand U4232 (N_4232,In_1945,In_729);
xor U4233 (N_4233,In_214,In_667);
or U4234 (N_4234,In_833,In_1386);
nand U4235 (N_4235,In_859,In_1280);
nor U4236 (N_4236,In_566,In_1440);
or U4237 (N_4237,In_861,In_1944);
and U4238 (N_4238,In_1629,In_735);
xor U4239 (N_4239,In_549,In_1029);
nor U4240 (N_4240,In_1052,In_15);
nor U4241 (N_4241,In_752,In_1279);
or U4242 (N_4242,In_712,In_1887);
nand U4243 (N_4243,In_744,In_1470);
nor U4244 (N_4244,In_979,In_286);
nand U4245 (N_4245,In_633,In_1839);
xnor U4246 (N_4246,In_1740,In_1366);
nor U4247 (N_4247,In_1135,In_403);
nand U4248 (N_4248,In_664,In_61);
xnor U4249 (N_4249,In_1845,In_712);
nand U4250 (N_4250,In_1962,In_1772);
or U4251 (N_4251,In_699,In_1400);
and U4252 (N_4252,In_108,In_1027);
xor U4253 (N_4253,In_650,In_391);
nand U4254 (N_4254,In_1445,In_1318);
nor U4255 (N_4255,In_574,In_314);
or U4256 (N_4256,In_646,In_1456);
or U4257 (N_4257,In_1502,In_1202);
and U4258 (N_4258,In_1182,In_1145);
xor U4259 (N_4259,In_893,In_1091);
nor U4260 (N_4260,In_1955,In_1546);
or U4261 (N_4261,In_483,In_1288);
nor U4262 (N_4262,In_898,In_1596);
nor U4263 (N_4263,In_10,In_1129);
nand U4264 (N_4264,In_747,In_1966);
nand U4265 (N_4265,In_1065,In_430);
nand U4266 (N_4266,In_1742,In_646);
and U4267 (N_4267,In_284,In_34);
or U4268 (N_4268,In_1537,In_279);
or U4269 (N_4269,In_1894,In_1969);
and U4270 (N_4270,In_1839,In_308);
nor U4271 (N_4271,In_1749,In_584);
nand U4272 (N_4272,In_1795,In_883);
nor U4273 (N_4273,In_545,In_1707);
nor U4274 (N_4274,In_1687,In_204);
nand U4275 (N_4275,In_701,In_1170);
and U4276 (N_4276,In_1927,In_98);
nand U4277 (N_4277,In_1315,In_1694);
and U4278 (N_4278,In_464,In_1212);
xor U4279 (N_4279,In_1133,In_514);
nor U4280 (N_4280,In_1791,In_635);
nand U4281 (N_4281,In_515,In_1343);
or U4282 (N_4282,In_1996,In_1658);
nor U4283 (N_4283,In_1801,In_1681);
nand U4284 (N_4284,In_1188,In_261);
or U4285 (N_4285,In_233,In_454);
or U4286 (N_4286,In_53,In_710);
and U4287 (N_4287,In_1747,In_1003);
nand U4288 (N_4288,In_1384,In_1733);
and U4289 (N_4289,In_1598,In_1047);
nand U4290 (N_4290,In_1272,In_569);
or U4291 (N_4291,In_355,In_1894);
or U4292 (N_4292,In_1367,In_1239);
and U4293 (N_4293,In_1523,In_1706);
or U4294 (N_4294,In_974,In_170);
nor U4295 (N_4295,In_113,In_547);
nor U4296 (N_4296,In_999,In_577);
xor U4297 (N_4297,In_991,In_230);
and U4298 (N_4298,In_803,In_801);
nand U4299 (N_4299,In_929,In_253);
and U4300 (N_4300,In_1138,In_1956);
nand U4301 (N_4301,In_803,In_358);
nand U4302 (N_4302,In_1095,In_1611);
or U4303 (N_4303,In_1419,In_384);
nor U4304 (N_4304,In_241,In_1706);
and U4305 (N_4305,In_297,In_384);
and U4306 (N_4306,In_1941,In_618);
nand U4307 (N_4307,In_74,In_632);
nand U4308 (N_4308,In_1863,In_90);
and U4309 (N_4309,In_621,In_1936);
and U4310 (N_4310,In_566,In_1486);
and U4311 (N_4311,In_1150,In_911);
and U4312 (N_4312,In_1778,In_1524);
or U4313 (N_4313,In_1617,In_1149);
nand U4314 (N_4314,In_302,In_1326);
nand U4315 (N_4315,In_1795,In_1092);
or U4316 (N_4316,In_1384,In_1534);
nor U4317 (N_4317,In_111,In_821);
nand U4318 (N_4318,In_1989,In_1058);
nand U4319 (N_4319,In_1123,In_484);
nor U4320 (N_4320,In_747,In_391);
nor U4321 (N_4321,In_1908,In_1651);
nor U4322 (N_4322,In_973,In_283);
or U4323 (N_4323,In_62,In_1652);
xnor U4324 (N_4324,In_208,In_945);
and U4325 (N_4325,In_915,In_179);
or U4326 (N_4326,In_0,In_1844);
and U4327 (N_4327,In_1422,In_950);
nor U4328 (N_4328,In_1094,In_1691);
nand U4329 (N_4329,In_848,In_1842);
and U4330 (N_4330,In_1748,In_938);
or U4331 (N_4331,In_376,In_931);
or U4332 (N_4332,In_665,In_1265);
nor U4333 (N_4333,In_22,In_1356);
nor U4334 (N_4334,In_1434,In_225);
and U4335 (N_4335,In_1021,In_498);
nand U4336 (N_4336,In_1769,In_1412);
or U4337 (N_4337,In_1776,In_633);
or U4338 (N_4338,In_1751,In_201);
nor U4339 (N_4339,In_1974,In_1151);
or U4340 (N_4340,In_903,In_370);
or U4341 (N_4341,In_263,In_698);
nand U4342 (N_4342,In_1467,In_1535);
nor U4343 (N_4343,In_1139,In_1170);
or U4344 (N_4344,In_44,In_702);
nand U4345 (N_4345,In_1332,In_1627);
or U4346 (N_4346,In_96,In_1554);
nor U4347 (N_4347,In_445,In_909);
xnor U4348 (N_4348,In_77,In_1840);
nand U4349 (N_4349,In_822,In_1147);
and U4350 (N_4350,In_511,In_1486);
or U4351 (N_4351,In_593,In_262);
nand U4352 (N_4352,In_1672,In_1599);
xor U4353 (N_4353,In_1029,In_646);
or U4354 (N_4354,In_1112,In_1910);
and U4355 (N_4355,In_1621,In_838);
and U4356 (N_4356,In_459,In_1619);
or U4357 (N_4357,In_107,In_164);
and U4358 (N_4358,In_672,In_42);
nand U4359 (N_4359,In_1375,In_604);
or U4360 (N_4360,In_1044,In_1671);
xor U4361 (N_4361,In_1869,In_1405);
nor U4362 (N_4362,In_526,In_1142);
or U4363 (N_4363,In_1190,In_359);
and U4364 (N_4364,In_249,In_1961);
nand U4365 (N_4365,In_952,In_429);
nor U4366 (N_4366,In_1290,In_1431);
and U4367 (N_4367,In_883,In_1488);
and U4368 (N_4368,In_1224,In_1961);
nand U4369 (N_4369,In_1003,In_497);
and U4370 (N_4370,In_1068,In_924);
xnor U4371 (N_4371,In_670,In_1032);
or U4372 (N_4372,In_947,In_276);
and U4373 (N_4373,In_1912,In_715);
or U4374 (N_4374,In_727,In_602);
and U4375 (N_4375,In_1478,In_1886);
or U4376 (N_4376,In_765,In_786);
and U4377 (N_4377,In_425,In_302);
nand U4378 (N_4378,In_1968,In_1366);
xor U4379 (N_4379,In_95,In_1223);
nand U4380 (N_4380,In_1091,In_1407);
or U4381 (N_4381,In_113,In_1818);
nor U4382 (N_4382,In_193,In_1190);
and U4383 (N_4383,In_824,In_405);
nor U4384 (N_4384,In_1811,In_332);
and U4385 (N_4385,In_1819,In_179);
nand U4386 (N_4386,In_374,In_1619);
or U4387 (N_4387,In_1669,In_1531);
nand U4388 (N_4388,In_708,In_475);
xnor U4389 (N_4389,In_1963,In_1377);
nor U4390 (N_4390,In_1892,In_502);
nor U4391 (N_4391,In_1669,In_1583);
nand U4392 (N_4392,In_63,In_1339);
and U4393 (N_4393,In_1629,In_1178);
or U4394 (N_4394,In_787,In_86);
or U4395 (N_4395,In_27,In_743);
nor U4396 (N_4396,In_1844,In_1384);
xnor U4397 (N_4397,In_298,In_466);
and U4398 (N_4398,In_1743,In_1458);
nand U4399 (N_4399,In_1126,In_1760);
or U4400 (N_4400,In_117,In_443);
and U4401 (N_4401,In_1969,In_598);
nand U4402 (N_4402,In_632,In_1213);
nor U4403 (N_4403,In_1095,In_1719);
or U4404 (N_4404,In_326,In_1608);
or U4405 (N_4405,In_766,In_1885);
or U4406 (N_4406,In_819,In_578);
xnor U4407 (N_4407,In_66,In_1744);
or U4408 (N_4408,In_849,In_1723);
and U4409 (N_4409,In_489,In_349);
nor U4410 (N_4410,In_1674,In_1183);
nand U4411 (N_4411,In_557,In_489);
nand U4412 (N_4412,In_1405,In_1992);
nor U4413 (N_4413,In_1957,In_535);
nand U4414 (N_4414,In_1038,In_88);
xnor U4415 (N_4415,In_109,In_420);
nor U4416 (N_4416,In_1217,In_591);
nor U4417 (N_4417,In_252,In_595);
or U4418 (N_4418,In_928,In_736);
nand U4419 (N_4419,In_1824,In_668);
and U4420 (N_4420,In_1231,In_1170);
nand U4421 (N_4421,In_1947,In_1021);
xor U4422 (N_4422,In_212,In_311);
nand U4423 (N_4423,In_265,In_829);
or U4424 (N_4424,In_406,In_343);
and U4425 (N_4425,In_474,In_1567);
nor U4426 (N_4426,In_1593,In_245);
and U4427 (N_4427,In_958,In_358);
nor U4428 (N_4428,In_902,In_1478);
nand U4429 (N_4429,In_1529,In_1935);
nand U4430 (N_4430,In_1613,In_391);
and U4431 (N_4431,In_698,In_1599);
and U4432 (N_4432,In_1484,In_284);
nand U4433 (N_4433,In_826,In_1393);
nor U4434 (N_4434,In_1297,In_77);
and U4435 (N_4435,In_1293,In_613);
and U4436 (N_4436,In_456,In_407);
or U4437 (N_4437,In_837,In_1627);
or U4438 (N_4438,In_162,In_316);
nor U4439 (N_4439,In_319,In_1245);
nand U4440 (N_4440,In_1312,In_1246);
nand U4441 (N_4441,In_500,In_983);
nor U4442 (N_4442,In_218,In_1530);
and U4443 (N_4443,In_1271,In_1146);
xor U4444 (N_4444,In_831,In_1868);
nor U4445 (N_4445,In_1490,In_616);
nand U4446 (N_4446,In_1531,In_1016);
nor U4447 (N_4447,In_233,In_245);
nor U4448 (N_4448,In_1875,In_1594);
or U4449 (N_4449,In_1212,In_1928);
nand U4450 (N_4450,In_260,In_1701);
or U4451 (N_4451,In_1569,In_1164);
nand U4452 (N_4452,In_1134,In_220);
or U4453 (N_4453,In_593,In_1714);
nand U4454 (N_4454,In_310,In_7);
nand U4455 (N_4455,In_713,In_34);
nand U4456 (N_4456,In_453,In_246);
and U4457 (N_4457,In_1626,In_387);
and U4458 (N_4458,In_1917,In_1889);
or U4459 (N_4459,In_280,In_673);
xor U4460 (N_4460,In_1946,In_680);
nor U4461 (N_4461,In_996,In_1729);
and U4462 (N_4462,In_1569,In_1637);
or U4463 (N_4463,In_1520,In_1897);
nand U4464 (N_4464,In_1812,In_1141);
or U4465 (N_4465,In_392,In_719);
nand U4466 (N_4466,In_1382,In_97);
nor U4467 (N_4467,In_834,In_1095);
or U4468 (N_4468,In_267,In_1819);
and U4469 (N_4469,In_1900,In_689);
and U4470 (N_4470,In_1374,In_1737);
or U4471 (N_4471,In_1121,In_1242);
and U4472 (N_4472,In_1723,In_1827);
nand U4473 (N_4473,In_1617,In_1184);
or U4474 (N_4474,In_71,In_640);
and U4475 (N_4475,In_6,In_249);
or U4476 (N_4476,In_1081,In_1417);
nand U4477 (N_4477,In_1732,In_54);
nand U4478 (N_4478,In_778,In_1551);
nor U4479 (N_4479,In_1664,In_318);
or U4480 (N_4480,In_959,In_318);
nand U4481 (N_4481,In_1501,In_968);
or U4482 (N_4482,In_1115,In_1492);
and U4483 (N_4483,In_827,In_684);
nor U4484 (N_4484,In_437,In_1313);
nand U4485 (N_4485,In_169,In_791);
nand U4486 (N_4486,In_1390,In_1144);
or U4487 (N_4487,In_1304,In_921);
nand U4488 (N_4488,In_803,In_935);
or U4489 (N_4489,In_1294,In_909);
or U4490 (N_4490,In_1941,In_251);
and U4491 (N_4491,In_263,In_1998);
xnor U4492 (N_4492,In_718,In_427);
nor U4493 (N_4493,In_746,In_1440);
and U4494 (N_4494,In_470,In_195);
or U4495 (N_4495,In_966,In_1184);
and U4496 (N_4496,In_1056,In_1304);
or U4497 (N_4497,In_200,In_534);
nor U4498 (N_4498,In_718,In_1046);
nor U4499 (N_4499,In_1152,In_776);
or U4500 (N_4500,In_1632,In_867);
nor U4501 (N_4501,In_960,In_328);
or U4502 (N_4502,In_794,In_1324);
or U4503 (N_4503,In_888,In_1127);
nor U4504 (N_4504,In_1474,In_1576);
xor U4505 (N_4505,In_220,In_1464);
and U4506 (N_4506,In_407,In_1212);
nor U4507 (N_4507,In_1469,In_1674);
nor U4508 (N_4508,In_1316,In_1901);
and U4509 (N_4509,In_720,In_74);
and U4510 (N_4510,In_539,In_1041);
and U4511 (N_4511,In_1189,In_354);
or U4512 (N_4512,In_1313,In_1768);
nor U4513 (N_4513,In_349,In_1347);
or U4514 (N_4514,In_127,In_536);
or U4515 (N_4515,In_1387,In_648);
xor U4516 (N_4516,In_808,In_948);
nor U4517 (N_4517,In_26,In_532);
nand U4518 (N_4518,In_1234,In_262);
nor U4519 (N_4519,In_212,In_656);
nand U4520 (N_4520,In_612,In_1014);
or U4521 (N_4521,In_1375,In_1373);
nor U4522 (N_4522,In_1857,In_453);
and U4523 (N_4523,In_1294,In_67);
or U4524 (N_4524,In_1534,In_409);
and U4525 (N_4525,In_1269,In_663);
nor U4526 (N_4526,In_848,In_632);
and U4527 (N_4527,In_1484,In_1764);
and U4528 (N_4528,In_1580,In_1810);
nand U4529 (N_4529,In_1997,In_1587);
nand U4530 (N_4530,In_1665,In_638);
or U4531 (N_4531,In_852,In_110);
and U4532 (N_4532,In_696,In_1729);
nor U4533 (N_4533,In_1587,In_213);
nand U4534 (N_4534,In_1772,In_74);
or U4535 (N_4535,In_968,In_1513);
nand U4536 (N_4536,In_236,In_984);
nor U4537 (N_4537,In_713,In_1606);
nor U4538 (N_4538,In_1721,In_1589);
or U4539 (N_4539,In_1560,In_636);
nand U4540 (N_4540,In_853,In_773);
or U4541 (N_4541,In_302,In_1420);
nand U4542 (N_4542,In_1912,In_1544);
xnor U4543 (N_4543,In_1822,In_331);
and U4544 (N_4544,In_439,In_1995);
nand U4545 (N_4545,In_116,In_700);
nand U4546 (N_4546,In_347,In_1895);
nand U4547 (N_4547,In_284,In_1790);
nand U4548 (N_4548,In_1701,In_290);
or U4549 (N_4549,In_355,In_391);
and U4550 (N_4550,In_1476,In_1104);
nand U4551 (N_4551,In_552,In_335);
nor U4552 (N_4552,In_813,In_94);
nor U4553 (N_4553,In_1735,In_1533);
or U4554 (N_4554,In_1596,In_745);
xor U4555 (N_4555,In_416,In_648);
and U4556 (N_4556,In_913,In_850);
and U4557 (N_4557,In_245,In_765);
and U4558 (N_4558,In_1270,In_1927);
or U4559 (N_4559,In_1076,In_729);
xor U4560 (N_4560,In_205,In_975);
nor U4561 (N_4561,In_1607,In_826);
nor U4562 (N_4562,In_1039,In_1650);
and U4563 (N_4563,In_584,In_738);
or U4564 (N_4564,In_777,In_1443);
nor U4565 (N_4565,In_903,In_1889);
nor U4566 (N_4566,In_166,In_353);
nor U4567 (N_4567,In_12,In_628);
nand U4568 (N_4568,In_1903,In_953);
or U4569 (N_4569,In_1899,In_557);
nand U4570 (N_4570,In_843,In_29);
or U4571 (N_4571,In_812,In_1593);
and U4572 (N_4572,In_520,In_1194);
and U4573 (N_4573,In_948,In_1657);
or U4574 (N_4574,In_833,In_1493);
nand U4575 (N_4575,In_1188,In_1080);
nor U4576 (N_4576,In_833,In_1796);
nand U4577 (N_4577,In_1820,In_392);
or U4578 (N_4578,In_957,In_431);
nor U4579 (N_4579,In_502,In_885);
or U4580 (N_4580,In_6,In_1753);
nor U4581 (N_4581,In_1404,In_1438);
nor U4582 (N_4582,In_1990,In_636);
or U4583 (N_4583,In_899,In_1591);
nor U4584 (N_4584,In_231,In_658);
and U4585 (N_4585,In_1585,In_817);
and U4586 (N_4586,In_451,In_886);
nand U4587 (N_4587,In_1555,In_1101);
nor U4588 (N_4588,In_872,In_151);
nor U4589 (N_4589,In_1877,In_733);
or U4590 (N_4590,In_16,In_1559);
nor U4591 (N_4591,In_828,In_1345);
or U4592 (N_4592,In_558,In_305);
or U4593 (N_4593,In_1826,In_417);
and U4594 (N_4594,In_1460,In_461);
or U4595 (N_4595,In_84,In_309);
and U4596 (N_4596,In_545,In_871);
and U4597 (N_4597,In_1481,In_1101);
and U4598 (N_4598,In_474,In_1854);
nand U4599 (N_4599,In_878,In_1981);
and U4600 (N_4600,In_1709,In_796);
nand U4601 (N_4601,In_1796,In_1608);
and U4602 (N_4602,In_267,In_1441);
or U4603 (N_4603,In_1688,In_390);
or U4604 (N_4604,In_1003,In_1782);
xor U4605 (N_4605,In_1453,In_1034);
and U4606 (N_4606,In_787,In_1116);
or U4607 (N_4607,In_811,In_1729);
or U4608 (N_4608,In_1164,In_1133);
xor U4609 (N_4609,In_1570,In_540);
and U4610 (N_4610,In_510,In_1309);
nor U4611 (N_4611,In_534,In_1801);
or U4612 (N_4612,In_1957,In_1220);
and U4613 (N_4613,In_1814,In_1724);
or U4614 (N_4614,In_1426,In_384);
nor U4615 (N_4615,In_592,In_1444);
or U4616 (N_4616,In_876,In_850);
and U4617 (N_4617,In_133,In_1155);
nor U4618 (N_4618,In_456,In_1090);
nand U4619 (N_4619,In_276,In_1465);
nor U4620 (N_4620,In_1500,In_1448);
nor U4621 (N_4621,In_732,In_1719);
nand U4622 (N_4622,In_1333,In_53);
nand U4623 (N_4623,In_303,In_26);
nor U4624 (N_4624,In_534,In_127);
nor U4625 (N_4625,In_1681,In_1461);
and U4626 (N_4626,In_376,In_510);
and U4627 (N_4627,In_975,In_440);
nor U4628 (N_4628,In_1162,In_1727);
or U4629 (N_4629,In_503,In_1007);
and U4630 (N_4630,In_1676,In_904);
and U4631 (N_4631,In_382,In_1170);
nand U4632 (N_4632,In_353,In_850);
or U4633 (N_4633,In_451,In_1984);
xnor U4634 (N_4634,In_711,In_360);
and U4635 (N_4635,In_1562,In_986);
or U4636 (N_4636,In_251,In_761);
and U4637 (N_4637,In_1274,In_893);
nand U4638 (N_4638,In_1937,In_203);
nor U4639 (N_4639,In_104,In_145);
nor U4640 (N_4640,In_827,In_1741);
nand U4641 (N_4641,In_1025,In_682);
nand U4642 (N_4642,In_355,In_402);
or U4643 (N_4643,In_1734,In_395);
nor U4644 (N_4644,In_1195,In_1241);
or U4645 (N_4645,In_1053,In_472);
xnor U4646 (N_4646,In_1907,In_879);
or U4647 (N_4647,In_1493,In_214);
nand U4648 (N_4648,In_1496,In_628);
or U4649 (N_4649,In_565,In_1725);
and U4650 (N_4650,In_967,In_983);
xor U4651 (N_4651,In_1487,In_94);
nor U4652 (N_4652,In_1232,In_920);
and U4653 (N_4653,In_123,In_1236);
and U4654 (N_4654,In_1113,In_10);
nor U4655 (N_4655,In_1707,In_357);
nand U4656 (N_4656,In_1822,In_1871);
nor U4657 (N_4657,In_1214,In_1444);
or U4658 (N_4658,In_963,In_258);
xor U4659 (N_4659,In_1996,In_510);
or U4660 (N_4660,In_292,In_1321);
and U4661 (N_4661,In_1575,In_179);
nand U4662 (N_4662,In_1583,In_424);
nor U4663 (N_4663,In_28,In_1818);
xnor U4664 (N_4664,In_1068,In_698);
nand U4665 (N_4665,In_1331,In_689);
nor U4666 (N_4666,In_447,In_1013);
xnor U4667 (N_4667,In_591,In_444);
nor U4668 (N_4668,In_6,In_1342);
nor U4669 (N_4669,In_60,In_596);
xor U4670 (N_4670,In_785,In_1227);
xnor U4671 (N_4671,In_1806,In_1552);
and U4672 (N_4672,In_1634,In_436);
and U4673 (N_4673,In_400,In_1851);
or U4674 (N_4674,In_1080,In_1347);
or U4675 (N_4675,In_654,In_394);
and U4676 (N_4676,In_1267,In_657);
nand U4677 (N_4677,In_1909,In_1797);
nand U4678 (N_4678,In_1509,In_582);
and U4679 (N_4679,In_973,In_509);
or U4680 (N_4680,In_759,In_1380);
xor U4681 (N_4681,In_1299,In_57);
or U4682 (N_4682,In_1762,In_1943);
or U4683 (N_4683,In_1251,In_924);
or U4684 (N_4684,In_1051,In_449);
and U4685 (N_4685,In_1952,In_564);
nor U4686 (N_4686,In_1584,In_1885);
and U4687 (N_4687,In_398,In_1533);
nand U4688 (N_4688,In_48,In_329);
and U4689 (N_4689,In_1400,In_1540);
or U4690 (N_4690,In_964,In_1352);
or U4691 (N_4691,In_23,In_1258);
or U4692 (N_4692,In_1034,In_587);
nor U4693 (N_4693,In_1404,In_1248);
xnor U4694 (N_4694,In_107,In_1021);
and U4695 (N_4695,In_1428,In_296);
and U4696 (N_4696,In_879,In_1478);
or U4697 (N_4697,In_475,In_1425);
nand U4698 (N_4698,In_178,In_1910);
nand U4699 (N_4699,In_678,In_1823);
or U4700 (N_4700,In_609,In_504);
or U4701 (N_4701,In_1799,In_492);
xor U4702 (N_4702,In_1054,In_855);
and U4703 (N_4703,In_1499,In_1654);
or U4704 (N_4704,In_1362,In_1755);
and U4705 (N_4705,In_1472,In_1720);
nor U4706 (N_4706,In_1635,In_48);
or U4707 (N_4707,In_601,In_1831);
or U4708 (N_4708,In_1696,In_293);
and U4709 (N_4709,In_520,In_1738);
nor U4710 (N_4710,In_445,In_1149);
nand U4711 (N_4711,In_1768,In_709);
or U4712 (N_4712,In_888,In_375);
nand U4713 (N_4713,In_1255,In_1076);
or U4714 (N_4714,In_479,In_1339);
nand U4715 (N_4715,In_235,In_1854);
or U4716 (N_4716,In_1497,In_1136);
or U4717 (N_4717,In_1585,In_81);
nand U4718 (N_4718,In_442,In_956);
nand U4719 (N_4719,In_500,In_189);
or U4720 (N_4720,In_1792,In_1823);
nand U4721 (N_4721,In_533,In_272);
xnor U4722 (N_4722,In_1779,In_1310);
nand U4723 (N_4723,In_599,In_860);
or U4724 (N_4724,In_444,In_100);
nand U4725 (N_4725,In_2,In_671);
xor U4726 (N_4726,In_1963,In_846);
or U4727 (N_4727,In_909,In_24);
or U4728 (N_4728,In_469,In_1300);
nand U4729 (N_4729,In_1862,In_1787);
xor U4730 (N_4730,In_1242,In_1308);
nor U4731 (N_4731,In_907,In_732);
or U4732 (N_4732,In_461,In_647);
xnor U4733 (N_4733,In_596,In_528);
nor U4734 (N_4734,In_257,In_869);
xnor U4735 (N_4735,In_0,In_84);
or U4736 (N_4736,In_496,In_676);
or U4737 (N_4737,In_265,In_718);
nand U4738 (N_4738,In_1088,In_1796);
or U4739 (N_4739,In_279,In_601);
nand U4740 (N_4740,In_1447,In_1943);
nor U4741 (N_4741,In_677,In_1405);
or U4742 (N_4742,In_1056,In_464);
or U4743 (N_4743,In_1170,In_787);
or U4744 (N_4744,In_1609,In_1556);
and U4745 (N_4745,In_359,In_1562);
nand U4746 (N_4746,In_967,In_1281);
nand U4747 (N_4747,In_115,In_1357);
nor U4748 (N_4748,In_800,In_1282);
nor U4749 (N_4749,In_1084,In_1385);
or U4750 (N_4750,In_921,In_543);
nand U4751 (N_4751,In_347,In_446);
and U4752 (N_4752,In_539,In_348);
or U4753 (N_4753,In_1850,In_530);
xnor U4754 (N_4754,In_1476,In_1003);
nand U4755 (N_4755,In_1464,In_609);
and U4756 (N_4756,In_1640,In_630);
nor U4757 (N_4757,In_337,In_1505);
or U4758 (N_4758,In_1530,In_881);
or U4759 (N_4759,In_695,In_1948);
xnor U4760 (N_4760,In_1989,In_1702);
nor U4761 (N_4761,In_1348,In_972);
nor U4762 (N_4762,In_500,In_898);
nor U4763 (N_4763,In_1072,In_1306);
nor U4764 (N_4764,In_1520,In_1221);
nor U4765 (N_4765,In_1070,In_169);
and U4766 (N_4766,In_1451,In_1926);
nor U4767 (N_4767,In_101,In_1165);
nand U4768 (N_4768,In_452,In_1264);
nor U4769 (N_4769,In_1827,In_878);
xnor U4770 (N_4770,In_674,In_1865);
nor U4771 (N_4771,In_282,In_132);
nor U4772 (N_4772,In_1108,In_1454);
nor U4773 (N_4773,In_1493,In_1622);
nor U4774 (N_4774,In_664,In_882);
nand U4775 (N_4775,In_820,In_14);
or U4776 (N_4776,In_1611,In_129);
nand U4777 (N_4777,In_141,In_652);
and U4778 (N_4778,In_470,In_1623);
or U4779 (N_4779,In_1375,In_1941);
xor U4780 (N_4780,In_1853,In_1144);
nor U4781 (N_4781,In_1480,In_468);
and U4782 (N_4782,In_1491,In_1705);
and U4783 (N_4783,In_436,In_550);
xnor U4784 (N_4784,In_1781,In_659);
or U4785 (N_4785,In_395,In_2);
or U4786 (N_4786,In_1546,In_302);
or U4787 (N_4787,In_383,In_133);
nor U4788 (N_4788,In_186,In_615);
and U4789 (N_4789,In_87,In_660);
or U4790 (N_4790,In_239,In_997);
nor U4791 (N_4791,In_330,In_1047);
or U4792 (N_4792,In_962,In_859);
nand U4793 (N_4793,In_1414,In_1004);
nand U4794 (N_4794,In_734,In_1101);
nand U4795 (N_4795,In_462,In_404);
nand U4796 (N_4796,In_1534,In_1782);
and U4797 (N_4797,In_1653,In_421);
xnor U4798 (N_4798,In_628,In_323);
or U4799 (N_4799,In_1407,In_1006);
xor U4800 (N_4800,In_971,In_1192);
nor U4801 (N_4801,In_1781,In_79);
nor U4802 (N_4802,In_1693,In_1739);
or U4803 (N_4803,In_1418,In_531);
nor U4804 (N_4804,In_228,In_1156);
or U4805 (N_4805,In_1591,In_1707);
nand U4806 (N_4806,In_85,In_315);
nand U4807 (N_4807,In_1257,In_997);
or U4808 (N_4808,In_1890,In_670);
nor U4809 (N_4809,In_442,In_486);
nor U4810 (N_4810,In_621,In_365);
xnor U4811 (N_4811,In_1089,In_1176);
and U4812 (N_4812,In_1024,In_317);
and U4813 (N_4813,In_1054,In_35);
or U4814 (N_4814,In_317,In_1036);
and U4815 (N_4815,In_1862,In_1142);
and U4816 (N_4816,In_1252,In_1375);
nand U4817 (N_4817,In_1898,In_660);
and U4818 (N_4818,In_1058,In_1700);
or U4819 (N_4819,In_93,In_306);
xor U4820 (N_4820,In_1355,In_1959);
and U4821 (N_4821,In_1467,In_1209);
or U4822 (N_4822,In_712,In_1844);
nor U4823 (N_4823,In_1065,In_1374);
and U4824 (N_4824,In_376,In_961);
nor U4825 (N_4825,In_1509,In_1658);
and U4826 (N_4826,In_669,In_103);
and U4827 (N_4827,In_1509,In_1152);
and U4828 (N_4828,In_1001,In_1689);
or U4829 (N_4829,In_160,In_1184);
nor U4830 (N_4830,In_1968,In_1963);
or U4831 (N_4831,In_1266,In_1937);
nor U4832 (N_4832,In_427,In_42);
nor U4833 (N_4833,In_1646,In_1660);
or U4834 (N_4834,In_1436,In_1973);
xnor U4835 (N_4835,In_410,In_1746);
nor U4836 (N_4836,In_199,In_778);
or U4837 (N_4837,In_706,In_1852);
and U4838 (N_4838,In_1807,In_1539);
nor U4839 (N_4839,In_617,In_1185);
and U4840 (N_4840,In_1672,In_966);
or U4841 (N_4841,In_796,In_1791);
or U4842 (N_4842,In_1165,In_1504);
or U4843 (N_4843,In_1814,In_1135);
nand U4844 (N_4844,In_1192,In_785);
or U4845 (N_4845,In_111,In_1048);
nor U4846 (N_4846,In_1882,In_1881);
nor U4847 (N_4847,In_497,In_157);
or U4848 (N_4848,In_1180,In_208);
or U4849 (N_4849,In_1028,In_581);
nand U4850 (N_4850,In_1980,In_1183);
and U4851 (N_4851,In_1444,In_703);
nor U4852 (N_4852,In_867,In_1856);
and U4853 (N_4853,In_392,In_830);
and U4854 (N_4854,In_1942,In_241);
nor U4855 (N_4855,In_868,In_1145);
nand U4856 (N_4856,In_60,In_380);
and U4857 (N_4857,In_974,In_219);
nor U4858 (N_4858,In_245,In_1664);
or U4859 (N_4859,In_1349,In_174);
nand U4860 (N_4860,In_926,In_1653);
nor U4861 (N_4861,In_1256,In_24);
xnor U4862 (N_4862,In_1446,In_1857);
and U4863 (N_4863,In_1279,In_683);
or U4864 (N_4864,In_1254,In_1482);
or U4865 (N_4865,In_1549,In_1629);
and U4866 (N_4866,In_72,In_804);
or U4867 (N_4867,In_1640,In_1581);
and U4868 (N_4868,In_190,In_1404);
and U4869 (N_4869,In_1592,In_1058);
nor U4870 (N_4870,In_102,In_1740);
and U4871 (N_4871,In_1479,In_1565);
and U4872 (N_4872,In_1773,In_94);
nand U4873 (N_4873,In_839,In_56);
nor U4874 (N_4874,In_1489,In_1132);
and U4875 (N_4875,In_861,In_418);
or U4876 (N_4876,In_1285,In_1167);
nor U4877 (N_4877,In_677,In_1611);
nor U4878 (N_4878,In_1222,In_1403);
nand U4879 (N_4879,In_1303,In_1604);
nor U4880 (N_4880,In_1437,In_1059);
nor U4881 (N_4881,In_1557,In_1320);
or U4882 (N_4882,In_121,In_1261);
or U4883 (N_4883,In_1177,In_1859);
nor U4884 (N_4884,In_1197,In_78);
nand U4885 (N_4885,In_1119,In_925);
or U4886 (N_4886,In_1501,In_1190);
xor U4887 (N_4887,In_869,In_1842);
nand U4888 (N_4888,In_845,In_1789);
nor U4889 (N_4889,In_508,In_1536);
nor U4890 (N_4890,In_739,In_323);
and U4891 (N_4891,In_1473,In_333);
nand U4892 (N_4892,In_471,In_454);
or U4893 (N_4893,In_73,In_545);
nor U4894 (N_4894,In_941,In_1168);
and U4895 (N_4895,In_1014,In_611);
nand U4896 (N_4896,In_288,In_1242);
or U4897 (N_4897,In_1514,In_66);
nor U4898 (N_4898,In_934,In_1808);
nand U4899 (N_4899,In_899,In_1478);
nor U4900 (N_4900,In_1932,In_1097);
nor U4901 (N_4901,In_357,In_1795);
nor U4902 (N_4902,In_1311,In_117);
nor U4903 (N_4903,In_1564,In_1515);
nor U4904 (N_4904,In_1094,In_1540);
and U4905 (N_4905,In_822,In_735);
xnor U4906 (N_4906,In_658,In_1540);
nand U4907 (N_4907,In_849,In_1406);
xor U4908 (N_4908,In_641,In_1203);
xor U4909 (N_4909,In_308,In_1974);
xnor U4910 (N_4910,In_550,In_474);
nand U4911 (N_4911,In_473,In_747);
nor U4912 (N_4912,In_461,In_1582);
nand U4913 (N_4913,In_712,In_1578);
nor U4914 (N_4914,In_263,In_623);
nand U4915 (N_4915,In_255,In_658);
nor U4916 (N_4916,In_1844,In_338);
nor U4917 (N_4917,In_1271,In_39);
and U4918 (N_4918,In_121,In_1730);
or U4919 (N_4919,In_1019,In_1710);
nor U4920 (N_4920,In_2,In_637);
nor U4921 (N_4921,In_1232,In_272);
nand U4922 (N_4922,In_1814,In_1808);
nand U4923 (N_4923,In_1792,In_1733);
and U4924 (N_4924,In_1038,In_346);
and U4925 (N_4925,In_388,In_1464);
xor U4926 (N_4926,In_63,In_1141);
and U4927 (N_4927,In_156,In_1978);
and U4928 (N_4928,In_332,In_1132);
or U4929 (N_4929,In_440,In_1343);
and U4930 (N_4930,In_878,In_211);
or U4931 (N_4931,In_1395,In_1034);
xor U4932 (N_4932,In_536,In_1860);
nor U4933 (N_4933,In_1797,In_544);
nor U4934 (N_4934,In_1716,In_222);
nor U4935 (N_4935,In_599,In_192);
nor U4936 (N_4936,In_38,In_656);
and U4937 (N_4937,In_1739,In_84);
nand U4938 (N_4938,In_1556,In_41);
xnor U4939 (N_4939,In_244,In_1788);
and U4940 (N_4940,In_662,In_1787);
nand U4941 (N_4941,In_947,In_1935);
and U4942 (N_4942,In_1560,In_1945);
and U4943 (N_4943,In_1168,In_1274);
nor U4944 (N_4944,In_1029,In_1371);
nor U4945 (N_4945,In_404,In_992);
xor U4946 (N_4946,In_1000,In_207);
nand U4947 (N_4947,In_1812,In_11);
nor U4948 (N_4948,In_981,In_626);
nand U4949 (N_4949,In_974,In_1224);
nand U4950 (N_4950,In_1627,In_386);
or U4951 (N_4951,In_292,In_1837);
nor U4952 (N_4952,In_24,In_356);
nor U4953 (N_4953,In_544,In_1360);
nand U4954 (N_4954,In_866,In_1814);
or U4955 (N_4955,In_644,In_400);
xor U4956 (N_4956,In_729,In_47);
and U4957 (N_4957,In_1211,In_51);
xnor U4958 (N_4958,In_1082,In_342);
nand U4959 (N_4959,In_57,In_1749);
nor U4960 (N_4960,In_535,In_1246);
and U4961 (N_4961,In_1717,In_1543);
or U4962 (N_4962,In_1494,In_157);
nor U4963 (N_4963,In_98,In_538);
nand U4964 (N_4964,In_565,In_353);
or U4965 (N_4965,In_1747,In_1488);
nor U4966 (N_4966,In_1314,In_101);
or U4967 (N_4967,In_1956,In_938);
and U4968 (N_4968,In_348,In_1511);
nand U4969 (N_4969,In_437,In_1547);
and U4970 (N_4970,In_1058,In_1622);
nand U4971 (N_4971,In_739,In_506);
xor U4972 (N_4972,In_292,In_576);
nor U4973 (N_4973,In_589,In_416);
and U4974 (N_4974,In_48,In_1387);
and U4975 (N_4975,In_1118,In_164);
or U4976 (N_4976,In_575,In_338);
or U4977 (N_4977,In_980,In_129);
nand U4978 (N_4978,In_390,In_220);
nor U4979 (N_4979,In_327,In_88);
or U4980 (N_4980,In_1134,In_230);
nor U4981 (N_4981,In_1997,In_1981);
and U4982 (N_4982,In_837,In_1263);
and U4983 (N_4983,In_826,In_1505);
nand U4984 (N_4984,In_1064,In_789);
and U4985 (N_4985,In_1846,In_1468);
or U4986 (N_4986,In_443,In_1169);
xnor U4987 (N_4987,In_768,In_258);
and U4988 (N_4988,In_1028,In_1523);
and U4989 (N_4989,In_398,In_1955);
or U4990 (N_4990,In_417,In_293);
and U4991 (N_4991,In_215,In_1753);
nand U4992 (N_4992,In_909,In_348);
or U4993 (N_4993,In_92,In_889);
or U4994 (N_4994,In_1681,In_484);
xor U4995 (N_4995,In_354,In_1663);
xor U4996 (N_4996,In_1947,In_1784);
xor U4997 (N_4997,In_1000,In_316);
and U4998 (N_4998,In_1053,In_499);
and U4999 (N_4999,In_431,In_880);
and U5000 (N_5000,N_2309,N_600);
nand U5001 (N_5001,N_3173,N_4297);
nand U5002 (N_5002,N_4326,N_3848);
nor U5003 (N_5003,N_2214,N_595);
nor U5004 (N_5004,N_2956,N_4278);
nor U5005 (N_5005,N_2538,N_4758);
or U5006 (N_5006,N_4345,N_3245);
nand U5007 (N_5007,N_2328,N_3316);
nand U5008 (N_5008,N_1617,N_4130);
and U5009 (N_5009,N_1951,N_4997);
and U5010 (N_5010,N_4347,N_2926);
and U5011 (N_5011,N_4514,N_4795);
nand U5012 (N_5012,N_4917,N_1297);
nor U5013 (N_5013,N_4127,N_399);
nand U5014 (N_5014,N_739,N_4006);
or U5015 (N_5015,N_4384,N_307);
or U5016 (N_5016,N_129,N_930);
xor U5017 (N_5017,N_3044,N_3124);
or U5018 (N_5018,N_4872,N_1314);
and U5019 (N_5019,N_3365,N_4283);
and U5020 (N_5020,N_2356,N_151);
nor U5021 (N_5021,N_508,N_3298);
nand U5022 (N_5022,N_1807,N_2868);
nor U5023 (N_5023,N_4670,N_2667);
nand U5024 (N_5024,N_191,N_3233);
or U5025 (N_5025,N_80,N_3780);
nor U5026 (N_5026,N_3289,N_4901);
and U5027 (N_5027,N_1776,N_758);
nor U5028 (N_5028,N_1852,N_2860);
nor U5029 (N_5029,N_3211,N_1840);
or U5030 (N_5030,N_4094,N_4449);
nor U5031 (N_5031,N_4859,N_4215);
nor U5032 (N_5032,N_2879,N_4823);
or U5033 (N_5033,N_3686,N_1964);
nor U5034 (N_5034,N_4181,N_2326);
xnor U5035 (N_5035,N_784,N_3128);
or U5036 (N_5036,N_2741,N_3244);
and U5037 (N_5037,N_4827,N_4579);
nand U5038 (N_5038,N_2774,N_3236);
and U5039 (N_5039,N_4694,N_1935);
nand U5040 (N_5040,N_1699,N_1121);
or U5041 (N_5041,N_966,N_3599);
and U5042 (N_5042,N_3088,N_3162);
nand U5043 (N_5043,N_2047,N_131);
nor U5044 (N_5044,N_4397,N_2573);
nor U5045 (N_5045,N_807,N_4117);
and U5046 (N_5046,N_1100,N_3594);
nor U5047 (N_5047,N_16,N_4342);
and U5048 (N_5048,N_3020,N_3426);
nand U5049 (N_5049,N_3308,N_1465);
and U5050 (N_5050,N_1226,N_71);
and U5051 (N_5051,N_4647,N_4325);
or U5052 (N_5052,N_4580,N_1391);
xnor U5053 (N_5053,N_4003,N_2599);
or U5054 (N_5054,N_1167,N_1948);
nor U5055 (N_5055,N_4222,N_1546);
nand U5056 (N_5056,N_1480,N_2636);
nor U5057 (N_5057,N_4780,N_4777);
nand U5058 (N_5058,N_368,N_4979);
nand U5059 (N_5059,N_2255,N_3938);
or U5060 (N_5060,N_23,N_2761);
or U5061 (N_5061,N_2021,N_3579);
nor U5062 (N_5062,N_3732,N_3635);
nand U5063 (N_5063,N_3603,N_3620);
and U5064 (N_5064,N_4096,N_3906);
and U5065 (N_5065,N_3272,N_1111);
nand U5066 (N_5066,N_513,N_589);
or U5067 (N_5067,N_2086,N_1108);
and U5068 (N_5068,N_2011,N_4816);
nor U5069 (N_5069,N_3184,N_701);
or U5070 (N_5070,N_1675,N_4078);
xnor U5071 (N_5071,N_2253,N_4155);
nand U5072 (N_5072,N_99,N_4961);
and U5073 (N_5073,N_1061,N_2828);
nor U5074 (N_5074,N_3217,N_1640);
or U5075 (N_5075,N_4951,N_887);
or U5076 (N_5076,N_4674,N_4451);
and U5077 (N_5077,N_2503,N_2690);
or U5078 (N_5078,N_2885,N_216);
and U5079 (N_5079,N_4160,N_4019);
nand U5080 (N_5080,N_2587,N_3553);
nor U5081 (N_5081,N_2040,N_123);
or U5082 (N_5082,N_2839,N_3076);
or U5083 (N_5083,N_3019,N_926);
and U5084 (N_5084,N_2207,N_1097);
or U5085 (N_5085,N_1728,N_156);
or U5086 (N_5086,N_1043,N_232);
xor U5087 (N_5087,N_1444,N_1901);
and U5088 (N_5088,N_1451,N_4730);
or U5089 (N_5089,N_4771,N_4878);
nor U5090 (N_5090,N_2299,N_3089);
nor U5091 (N_5091,N_1014,N_2558);
and U5092 (N_5092,N_3218,N_4529);
nand U5093 (N_5093,N_3182,N_4273);
nand U5094 (N_5094,N_4282,N_803);
xnor U5095 (N_5095,N_2897,N_2089);
or U5096 (N_5096,N_956,N_3597);
xnor U5097 (N_5097,N_2576,N_1742);
nor U5098 (N_5098,N_722,N_712);
nand U5099 (N_5099,N_1495,N_1659);
and U5100 (N_5100,N_3480,N_1323);
and U5101 (N_5101,N_4124,N_119);
nand U5102 (N_5102,N_1357,N_155);
and U5103 (N_5103,N_138,N_4533);
and U5104 (N_5104,N_1073,N_19);
nor U5105 (N_5105,N_2051,N_321);
and U5106 (N_5106,N_3009,N_3045);
nand U5107 (N_5107,N_348,N_4088);
nand U5108 (N_5108,N_295,N_3264);
nor U5109 (N_5109,N_2130,N_2683);
nand U5110 (N_5110,N_1739,N_1668);
and U5111 (N_5111,N_1956,N_3057);
nand U5112 (N_5112,N_2807,N_4501);
xnor U5113 (N_5113,N_3969,N_3136);
xnor U5114 (N_5114,N_2606,N_3622);
nor U5115 (N_5115,N_943,N_3806);
xnor U5116 (N_5116,N_4252,N_4906);
nor U5117 (N_5117,N_1228,N_4836);
or U5118 (N_5118,N_685,N_3572);
and U5119 (N_5119,N_1512,N_4043);
nor U5120 (N_5120,N_329,N_337);
and U5121 (N_5121,N_4865,N_2111);
nand U5122 (N_5122,N_3214,N_4148);
nand U5123 (N_5123,N_2343,N_3836);
nand U5124 (N_5124,N_4195,N_3667);
or U5125 (N_5125,N_945,N_4495);
and U5126 (N_5126,N_1486,N_148);
nor U5127 (N_5127,N_1131,N_3285);
nand U5128 (N_5128,N_3766,N_2507);
nor U5129 (N_5129,N_4534,N_3249);
nand U5130 (N_5130,N_1576,N_147);
and U5131 (N_5131,N_1696,N_2793);
nor U5132 (N_5132,N_2217,N_2);
nor U5133 (N_5133,N_3976,N_362);
nor U5134 (N_5134,N_3576,N_1849);
and U5135 (N_5135,N_2300,N_648);
or U5136 (N_5136,N_573,N_3439);
and U5137 (N_5137,N_455,N_1508);
nand U5138 (N_5138,N_2026,N_3159);
nand U5139 (N_5139,N_890,N_4556);
nand U5140 (N_5140,N_2668,N_1063);
xor U5141 (N_5141,N_4938,N_1866);
nand U5142 (N_5142,N_965,N_1406);
nor U5143 (N_5143,N_1544,N_1745);
nor U5144 (N_5144,N_2733,N_1494);
or U5145 (N_5145,N_4856,N_139);
and U5146 (N_5146,N_3802,N_3811);
nand U5147 (N_5147,N_4058,N_892);
nor U5148 (N_5148,N_1672,N_4469);
nand U5149 (N_5149,N_4757,N_950);
nor U5150 (N_5150,N_4732,N_4850);
and U5151 (N_5151,N_838,N_2732);
and U5152 (N_5152,N_4335,N_1091);
or U5153 (N_5153,N_4753,N_1527);
and U5154 (N_5154,N_3307,N_227);
nand U5155 (N_5155,N_1263,N_651);
and U5156 (N_5156,N_4327,N_1693);
xor U5157 (N_5157,N_4625,N_1504);
nand U5158 (N_5158,N_1254,N_1239);
nand U5159 (N_5159,N_2240,N_1242);
or U5160 (N_5160,N_3041,N_2292);
nand U5161 (N_5161,N_2940,N_235);
nor U5162 (N_5162,N_2184,N_4992);
nor U5163 (N_5163,N_1196,N_1836);
or U5164 (N_5164,N_4959,N_1031);
nand U5165 (N_5165,N_539,N_3452);
nor U5166 (N_5166,N_2059,N_2035);
and U5167 (N_5167,N_2015,N_3016);
nor U5168 (N_5168,N_3784,N_4634);
or U5169 (N_5169,N_3427,N_4035);
and U5170 (N_5170,N_3065,N_3582);
and U5171 (N_5171,N_336,N_3751);
or U5172 (N_5172,N_2395,N_2904);
or U5173 (N_5173,N_1846,N_3372);
nand U5174 (N_5174,N_4635,N_2675);
or U5175 (N_5175,N_2983,N_2321);
nand U5176 (N_5176,N_1850,N_2799);
or U5177 (N_5177,N_4624,N_1268);
or U5178 (N_5178,N_4955,N_4974);
nor U5179 (N_5179,N_3261,N_578);
nand U5180 (N_5180,N_2482,N_2486);
and U5181 (N_5181,N_3359,N_4266);
and U5182 (N_5182,N_4542,N_1454);
or U5183 (N_5183,N_3896,N_4401);
or U5184 (N_5184,N_4973,N_2781);
or U5185 (N_5185,N_3329,N_538);
nor U5186 (N_5186,N_3197,N_4191);
or U5187 (N_5187,N_176,N_1394);
and U5188 (N_5188,N_1908,N_4940);
nand U5189 (N_5189,N_204,N_2596);
nand U5190 (N_5190,N_396,N_2866);
nand U5191 (N_5191,N_891,N_1806);
or U5192 (N_5192,N_4581,N_3335);
nand U5193 (N_5193,N_4792,N_440);
nand U5194 (N_5194,N_1980,N_39);
and U5195 (N_5195,N_1190,N_1855);
nand U5196 (N_5196,N_4456,N_2802);
and U5197 (N_5197,N_3604,N_4369);
and U5198 (N_5198,N_2995,N_2716);
and U5199 (N_5199,N_1760,N_1626);
or U5200 (N_5200,N_4560,N_883);
nor U5201 (N_5201,N_3042,N_2544);
nand U5202 (N_5202,N_2796,N_361);
xnor U5203 (N_5203,N_2391,N_2303);
nor U5204 (N_5204,N_671,N_2663);
nor U5205 (N_5205,N_563,N_3734);
nand U5206 (N_5206,N_1689,N_4781);
xor U5207 (N_5207,N_639,N_2138);
and U5208 (N_5208,N_2669,N_757);
nor U5209 (N_5209,N_3823,N_4405);
nor U5210 (N_5210,N_3382,N_2585);
nor U5211 (N_5211,N_593,N_3440);
or U5212 (N_5212,N_798,N_4180);
and U5213 (N_5213,N_2363,N_2920);
or U5214 (N_5214,N_4292,N_2247);
nand U5215 (N_5215,N_1040,N_3477);
and U5216 (N_5216,N_4047,N_1525);
nor U5217 (N_5217,N_3060,N_17);
xnor U5218 (N_5218,N_1079,N_2360);
or U5219 (N_5219,N_3221,N_2088);
nand U5220 (N_5220,N_4386,N_679);
nor U5221 (N_5221,N_2156,N_385);
nor U5222 (N_5222,N_3761,N_1996);
nand U5223 (N_5223,N_692,N_2944);
nand U5224 (N_5224,N_2730,N_1518);
and U5225 (N_5225,N_4804,N_2206);
or U5226 (N_5226,N_1028,N_4843);
or U5227 (N_5227,N_4923,N_4935);
and U5228 (N_5228,N_468,N_4614);
and U5229 (N_5229,N_4887,N_4566);
nor U5230 (N_5230,N_1348,N_3101);
nor U5231 (N_5231,N_942,N_1255);
nor U5232 (N_5232,N_1788,N_1191);
or U5233 (N_5233,N_2313,N_3633);
xnor U5234 (N_5234,N_4165,N_3792);
or U5235 (N_5235,N_3405,N_4832);
and U5236 (N_5236,N_163,N_4174);
nor U5237 (N_5237,N_3430,N_4914);
nand U5238 (N_5238,N_3425,N_4380);
nand U5239 (N_5239,N_1984,N_1256);
xor U5240 (N_5240,N_4686,N_3420);
xnor U5241 (N_5241,N_542,N_3978);
nor U5242 (N_5242,N_3879,N_1827);
xor U5243 (N_5243,N_2264,N_4368);
or U5244 (N_5244,N_3283,N_364);
nand U5245 (N_5245,N_3276,N_844);
nor U5246 (N_5246,N_1030,N_4038);
nand U5247 (N_5247,N_932,N_878);
and U5248 (N_5248,N_630,N_2621);
and U5249 (N_5249,N_3115,N_2519);
or U5250 (N_5250,N_283,N_1000);
nand U5251 (N_5251,N_1279,N_4442);
nand U5252 (N_5252,N_3393,N_3563);
or U5253 (N_5253,N_2358,N_497);
nor U5254 (N_5254,N_528,N_958);
or U5255 (N_5255,N_192,N_1733);
or U5256 (N_5256,N_1194,N_3254);
xnor U5257 (N_5257,N_2268,N_535);
nor U5258 (N_5258,N_3110,N_3927);
or U5259 (N_5259,N_1053,N_3485);
nor U5260 (N_5260,N_4661,N_771);
nor U5261 (N_5261,N_4659,N_2511);
nand U5262 (N_5262,N_4595,N_806);
and U5263 (N_5263,N_1823,N_318);
and U5264 (N_5264,N_2662,N_2929);
nor U5265 (N_5265,N_986,N_2000);
nor U5266 (N_5266,N_817,N_1140);
nand U5267 (N_5267,N_1708,N_1877);
nor U5268 (N_5268,N_531,N_561);
and U5269 (N_5269,N_1630,N_3137);
nor U5270 (N_5270,N_3967,N_4217);
and U5271 (N_5271,N_1312,N_3215);
nand U5272 (N_5272,N_1857,N_3656);
nor U5273 (N_5273,N_4285,N_3730);
and U5274 (N_5274,N_3237,N_2136);
xnor U5275 (N_5275,N_697,N_3388);
or U5276 (N_5276,N_4607,N_1257);
xnor U5277 (N_5277,N_1511,N_1738);
and U5278 (N_5278,N_3345,N_4313);
nand U5279 (N_5279,N_2372,N_580);
nand U5280 (N_5280,N_634,N_4485);
xor U5281 (N_5281,N_2842,N_3188);
and U5282 (N_5282,N_4178,N_68);
nor U5283 (N_5283,N_1241,N_4101);
nor U5284 (N_5284,N_611,N_1155);
nand U5285 (N_5285,N_3573,N_657);
nor U5286 (N_5286,N_2124,N_3257);
and U5287 (N_5287,N_4837,N_1673);
or U5288 (N_5288,N_4762,N_1897);
nor U5289 (N_5289,N_1808,N_4724);
nand U5290 (N_5290,N_2525,N_4765);
xor U5291 (N_5291,N_3996,N_1260);
or U5292 (N_5292,N_2362,N_824);
or U5293 (N_5293,N_1747,N_3346);
xnor U5294 (N_5294,N_1661,N_158);
and U5295 (N_5295,N_3856,N_1837);
and U5296 (N_5296,N_2581,N_1744);
and U5297 (N_5297,N_767,N_3474);
xnor U5298 (N_5298,N_4681,N_4122);
or U5299 (N_5299,N_287,N_105);
xor U5300 (N_5300,N_84,N_1178);
nand U5301 (N_5301,N_1386,N_4689);
nand U5302 (N_5302,N_3096,N_2421);
nor U5303 (N_5303,N_2789,N_1423);
nand U5304 (N_5304,N_1695,N_3810);
or U5305 (N_5305,N_2521,N_3581);
nand U5306 (N_5306,N_202,N_1915);
nand U5307 (N_5307,N_3093,N_1607);
and U5308 (N_5308,N_2711,N_924);
xnor U5309 (N_5309,N_818,N_2458);
nor U5310 (N_5310,N_490,N_4862);
xor U5311 (N_5311,N_1482,N_4507);
nor U5312 (N_5312,N_1906,N_4294);
or U5313 (N_5313,N_1200,N_3659);
nand U5314 (N_5314,N_4551,N_1685);
nand U5315 (N_5315,N_334,N_2344);
nor U5316 (N_5316,N_1970,N_34);
nor U5317 (N_5317,N_1417,N_1118);
xor U5318 (N_5318,N_4840,N_2477);
xor U5319 (N_5319,N_3523,N_30);
nand U5320 (N_5320,N_212,N_523);
nand U5321 (N_5321,N_1973,N_3947);
and U5322 (N_5322,N_587,N_1151);
or U5323 (N_5323,N_917,N_2226);
nor U5324 (N_5324,N_1765,N_2151);
and U5325 (N_5325,N_3818,N_206);
nor U5326 (N_5326,N_4939,N_494);
or U5327 (N_5327,N_832,N_322);
or U5328 (N_5328,N_3959,N_1321);
nor U5329 (N_5329,N_1360,N_239);
nand U5330 (N_5330,N_4336,N_1054);
nand U5331 (N_5331,N_2960,N_3488);
nand U5332 (N_5332,N_444,N_2735);
and U5333 (N_5333,N_940,N_4735);
nor U5334 (N_5334,N_4594,N_354);
nor U5335 (N_5335,N_1815,N_4791);
nand U5336 (N_5336,N_3478,N_3641);
and U5337 (N_5337,N_2227,N_4298);
nor U5338 (N_5338,N_3479,N_584);
and U5339 (N_5339,N_4240,N_3195);
and U5340 (N_5340,N_1313,N_3164);
and U5341 (N_5341,N_1130,N_3491);
or U5342 (N_5342,N_3074,N_4963);
nand U5343 (N_5343,N_4158,N_4597);
nand U5344 (N_5344,N_540,N_2348);
and U5345 (N_5345,N_568,N_2623);
nor U5346 (N_5346,N_1233,N_4864);
and U5347 (N_5347,N_2847,N_4330);
nand U5348 (N_5348,N_3031,N_1210);
and U5349 (N_5349,N_387,N_853);
nand U5350 (N_5350,N_2301,N_209);
or U5351 (N_5351,N_2287,N_2512);
and U5352 (N_5352,N_137,N_2390);
or U5353 (N_5353,N_873,N_3299);
nand U5354 (N_5354,N_2575,N_2568);
nor U5355 (N_5355,N_3246,N_303);
nor U5356 (N_5356,N_1707,N_747);
nand U5357 (N_5357,N_552,N_1109);
nand U5358 (N_5358,N_2579,N_505);
and U5359 (N_5359,N_4225,N_470);
nor U5360 (N_5360,N_2405,N_4902);
or U5361 (N_5361,N_833,N_677);
nand U5362 (N_5362,N_2834,N_4880);
nor U5363 (N_5363,N_243,N_4817);
nand U5364 (N_5364,N_211,N_3116);
nor U5365 (N_5365,N_1520,N_1794);
or U5366 (N_5366,N_4554,N_3004);
nand U5367 (N_5367,N_1577,N_4544);
nor U5368 (N_5368,N_782,N_1496);
nor U5369 (N_5369,N_426,N_35);
nor U5370 (N_5370,N_915,N_1472);
nor U5371 (N_5371,N_2996,N_1272);
nor U5372 (N_5372,N_4164,N_1998);
or U5373 (N_5373,N_2819,N_2312);
or U5374 (N_5374,N_4565,N_3629);
and U5375 (N_5375,N_4466,N_3681);
or U5376 (N_5376,N_352,N_826);
nand U5377 (N_5377,N_3022,N_2892);
or U5378 (N_5378,N_876,N_2204);
or U5379 (N_5379,N_2531,N_2355);
nand U5380 (N_5380,N_4219,N_1952);
or U5381 (N_5381,N_4848,N_2141);
and U5382 (N_5382,N_2058,N_3274);
nor U5383 (N_5383,N_668,N_1663);
or U5384 (N_5384,N_1466,N_1162);
and U5385 (N_5385,N_1221,N_646);
and U5386 (N_5386,N_3558,N_3841);
or U5387 (N_5387,N_3112,N_4839);
nor U5388 (N_5388,N_1845,N_617);
nor U5389 (N_5389,N_3339,N_3153);
xor U5390 (N_5390,N_1428,N_2024);
nor U5391 (N_5391,N_2656,N_2388);
xnor U5392 (N_5392,N_1336,N_2549);
and U5393 (N_5393,N_1538,N_2384);
nor U5394 (N_5394,N_4896,N_710);
nand U5395 (N_5395,N_1563,N_2784);
xor U5396 (N_5396,N_2378,N_1289);
nor U5397 (N_5397,N_1521,N_4455);
and U5398 (N_5398,N_3338,N_1045);
nand U5399 (N_5399,N_4739,N_4747);
nor U5400 (N_5400,N_2112,N_1631);
or U5401 (N_5401,N_529,N_213);
and U5402 (N_5402,N_721,N_2065);
nand U5403 (N_5403,N_4564,N_4348);
or U5404 (N_5404,N_3490,N_2472);
nor U5405 (N_5405,N_4526,N_3929);
and U5406 (N_5406,N_1570,N_909);
nand U5407 (N_5407,N_4211,N_2666);
or U5408 (N_5408,N_4582,N_1723);
xor U5409 (N_5409,N_3500,N_3658);
nand U5410 (N_5410,N_558,N_1035);
nor U5411 (N_5411,N_4891,N_2517);
xor U5412 (N_5412,N_823,N_2710);
or U5413 (N_5413,N_4632,N_2106);
nor U5414 (N_5414,N_330,N_3105);
or U5415 (N_5415,N_2137,N_3349);
and U5416 (N_5416,N_3034,N_2870);
and U5417 (N_5417,N_2044,N_4616);
and U5418 (N_5418,N_2357,N_1821);
xnor U5419 (N_5419,N_240,N_2972);
and U5420 (N_5420,N_2645,N_4194);
and U5421 (N_5421,N_4382,N_4677);
or U5422 (N_5422,N_4408,N_1800);
or U5423 (N_5423,N_4941,N_4262);
nor U5424 (N_5424,N_4633,N_2790);
nor U5425 (N_5425,N_3753,N_4621);
xor U5426 (N_5426,N_1421,N_1900);
or U5427 (N_5427,N_755,N_1802);
nor U5428 (N_5428,N_3931,N_1614);
or U5429 (N_5429,N_44,N_2444);
and U5430 (N_5430,N_4143,N_2166);
nor U5431 (N_5431,N_2397,N_2967);
nand U5432 (N_5432,N_245,N_2977);
or U5433 (N_5433,N_3552,N_370);
nor U5434 (N_5434,N_929,N_3600);
nor U5435 (N_5435,N_2561,N_4705);
nor U5436 (N_5436,N_4729,N_4908);
nand U5437 (N_5437,N_2708,N_1912);
and U5438 (N_5438,N_2496,N_4053);
nor U5439 (N_5439,N_3156,N_1934);
and U5440 (N_5440,N_1785,N_691);
xnor U5441 (N_5441,N_1771,N_2750);
nand U5442 (N_5442,N_643,N_3417);
or U5443 (N_5443,N_2428,N_4310);
and U5444 (N_5444,N_948,N_3690);
or U5445 (N_5445,N_1379,N_4928);
or U5446 (N_5446,N_1224,N_2552);
or U5447 (N_5447,N_2896,N_3917);
nand U5448 (N_5448,N_2365,N_2332);
or U5449 (N_5449,N_4018,N_604);
and U5450 (N_5450,N_406,N_4700);
nand U5451 (N_5451,N_1600,N_2696);
or U5452 (N_5452,N_4617,N_4587);
xor U5453 (N_5453,N_3281,N_2043);
or U5454 (N_5454,N_3240,N_3389);
nor U5455 (N_5455,N_955,N_4321);
nand U5456 (N_5456,N_74,N_3470);
and U5457 (N_5457,N_1368,N_2942);
or U5458 (N_5458,N_3235,N_4135);
or U5459 (N_5459,N_2122,N_3348);
nor U5460 (N_5460,N_484,N_3733);
nor U5461 (N_5461,N_3125,N_38);
nor U5462 (N_5462,N_78,N_3185);
nor U5463 (N_5463,N_1058,N_193);
nor U5464 (N_5464,N_702,N_4322);
nand U5465 (N_5465,N_1896,N_1356);
nor U5466 (N_5466,N_2975,N_1981);
or U5467 (N_5467,N_3984,N_4858);
or U5468 (N_5468,N_2808,N_2671);
and U5469 (N_5469,N_3271,N_907);
or U5470 (N_5470,N_506,N_3242);
nor U5471 (N_5471,N_4479,N_2233);
nor U5472 (N_5472,N_3707,N_445);
nand U5473 (N_5473,N_1294,N_4084);
and U5474 (N_5474,N_2695,N_2113);
nand U5475 (N_5475,N_3243,N_162);
nor U5476 (N_5476,N_1519,N_3516);
and U5477 (N_5477,N_4618,N_3058);
nand U5478 (N_5478,N_4190,N_740);
or U5479 (N_5479,N_1502,N_1326);
nand U5480 (N_5480,N_4026,N_4360);
xnor U5481 (N_5481,N_1070,N_609);
and U5482 (N_5482,N_1916,N_4697);
and U5483 (N_5483,N_495,N_3496);
nand U5484 (N_5484,N_2578,N_4299);
and U5485 (N_5485,N_3035,N_4966);
nand U5486 (N_5486,N_1447,N_811);
nand U5487 (N_5487,N_2811,N_1752);
and U5488 (N_5488,N_316,N_973);
xnor U5489 (N_5489,N_2293,N_2075);
and U5490 (N_5490,N_2545,N_2825);
nor U5491 (N_5491,N_3054,N_3351);
and U5492 (N_5492,N_900,N_2354);
and U5493 (N_5493,N_3857,N_292);
nor U5494 (N_5494,N_3229,N_867);
or U5495 (N_5495,N_1266,N_4344);
and U5496 (N_5496,N_1625,N_4432);
and U5497 (N_5497,N_3864,N_3828);
nand U5498 (N_5498,N_3962,N_3071);
or U5499 (N_5499,N_3369,N_473);
or U5500 (N_5500,N_2001,N_82);
nand U5501 (N_5501,N_884,N_1829);
nand U5502 (N_5502,N_4125,N_4287);
nor U5503 (N_5503,N_1475,N_4524);
and U5504 (N_5504,N_4583,N_1875);
nand U5505 (N_5505,N_500,N_4482);
nor U5506 (N_5506,N_1461,N_3158);
or U5507 (N_5507,N_1619,N_550);
nand U5508 (N_5508,N_4573,N_1243);
and U5509 (N_5509,N_1522,N_1982);
nor U5510 (N_5510,N_1277,N_4413);
and U5511 (N_5511,N_3404,N_2569);
and U5512 (N_5512,N_4079,N_3596);
nand U5513 (N_5513,N_1290,N_751);
and U5514 (N_5514,N_3903,N_1950);
nand U5515 (N_5515,N_3080,N_486);
nand U5516 (N_5516,N_3981,N_2199);
xor U5517 (N_5517,N_4365,N_2943);
nor U5518 (N_5518,N_1531,N_4000);
and U5519 (N_5519,N_143,N_1703);
nand U5520 (N_5520,N_4210,N_10);
or U5521 (N_5521,N_4609,N_3670);
nor U5522 (N_5522,N_2245,N_4809);
nor U5523 (N_5523,N_400,N_866);
nand U5524 (N_5524,N_4366,N_2631);
or U5525 (N_5525,N_310,N_3181);
nor U5526 (N_5526,N_2403,N_4358);
nor U5527 (N_5527,N_3370,N_413);
nand U5528 (N_5528,N_4188,N_3796);
and U5529 (N_5529,N_2702,N_3831);
nor U5530 (N_5530,N_4340,N_1753);
nor U5531 (N_5531,N_1425,N_2154);
or U5532 (N_5532,N_4831,N_4289);
nor U5533 (N_5533,N_4076,N_1832);
nand U5534 (N_5534,N_4846,N_3736);
nand U5535 (N_5535,N_4478,N_4286);
and U5536 (N_5536,N_298,N_1083);
and U5537 (N_5537,N_636,N_605);
nor U5538 (N_5538,N_972,N_4776);
and U5539 (N_5539,N_4688,N_3321);
nand U5540 (N_5540,N_4907,N_971);
xor U5541 (N_5541,N_1944,N_4978);
xnor U5542 (N_5542,N_4658,N_1138);
nor U5543 (N_5543,N_1868,N_4568);
or U5544 (N_5544,N_2768,N_2805);
nor U5545 (N_5545,N_4717,N_2485);
or U5546 (N_5546,N_4768,N_4712);
and U5547 (N_5547,N_4610,N_1732);
nor U5548 (N_5548,N_2175,N_1334);
xor U5549 (N_5549,N_3531,N_1358);
or U5550 (N_5550,N_2727,N_4701);
nor U5551 (N_5551,N_773,N_2817);
nor U5552 (N_5552,N_3548,N_678);
nand U5553 (N_5553,N_2165,N_1678);
nor U5554 (N_5554,N_2908,N_4539);
nor U5555 (N_5555,N_3443,N_2193);
xor U5556 (N_5556,N_2862,N_168);
nand U5557 (N_5557,N_190,N_391);
or U5558 (N_5558,N_1680,N_4049);
or U5559 (N_5559,N_4468,N_2700);
and U5560 (N_5560,N_1917,N_111);
or U5561 (N_5561,N_2346,N_479);
xnor U5562 (N_5562,N_2787,N_2627);
and U5563 (N_5563,N_4206,N_3875);
nand U5564 (N_5564,N_3511,N_3398);
nor U5565 (N_5565,N_2964,N_4280);
and U5566 (N_5566,N_1104,N_896);
xnor U5567 (N_5567,N_3460,N_4502);
or U5568 (N_5568,N_1959,N_3627);
nand U5569 (N_5569,N_3987,N_1572);
nand U5570 (N_5570,N_4664,N_4116);
and U5571 (N_5571,N_2597,N_3654);
xnor U5572 (N_5572,N_1187,N_3560);
nand U5573 (N_5573,N_3555,N_3433);
nor U5574 (N_5574,N_1966,N_556);
nand U5575 (N_5575,N_4142,N_3677);
nand U5576 (N_5576,N_353,N_4435);
or U5577 (N_5577,N_1139,N_637);
nand U5578 (N_5578,N_1468,N_1422);
and U5579 (N_5579,N_1276,N_4668);
xnor U5580 (N_5580,N_459,N_642);
or U5581 (N_5581,N_4975,N_1351);
nor U5582 (N_5582,N_3256,N_1185);
nand U5583 (N_5583,N_4748,N_207);
and U5584 (N_5584,N_1628,N_1904);
nor U5585 (N_5585,N_2046,N_793);
and U5586 (N_5586,N_1925,N_91);
or U5587 (N_5587,N_3739,N_3935);
nor U5588 (N_5588,N_3203,N_1976);
or U5589 (N_5589,N_69,N_3362);
and U5590 (N_5590,N_2595,N_4259);
or U5591 (N_5591,N_1426,N_2563);
and U5592 (N_5592,N_4013,N_2469);
nand U5593 (N_5593,N_544,N_2102);
nand U5594 (N_5594,N_536,N_4028);
or U5595 (N_5595,N_3375,N_1936);
or U5596 (N_5596,N_1974,N_1350);
xor U5597 (N_5597,N_2854,N_1892);
nor U5598 (N_5598,N_3717,N_4139);
and U5599 (N_5599,N_2389,N_901);
and U5600 (N_5600,N_3133,N_619);
nand U5601 (N_5601,N_1259,N_4231);
or U5602 (N_5602,N_1005,N_4806);
nor U5603 (N_5603,N_3637,N_2949);
or U5604 (N_5604,N_3591,N_3092);
or U5605 (N_5605,N_98,N_1088);
xnor U5606 (N_5606,N_3771,N_408);
nand U5607 (N_5607,N_3401,N_3788);
and U5608 (N_5608,N_402,N_4773);
nand U5609 (N_5609,N_968,N_2013);
nand U5610 (N_5610,N_1036,N_3201);
nand U5611 (N_5611,N_1193,N_3565);
or U5612 (N_5612,N_1355,N_1069);
nor U5613 (N_5613,N_746,N_2653);
or U5614 (N_5614,N_1437,N_4745);
or U5615 (N_5615,N_1361,N_4156);
nor U5616 (N_5616,N_1669,N_2160);
nor U5617 (N_5617,N_2100,N_1181);
xnor U5618 (N_5618,N_2280,N_2213);
nand U5619 (N_5619,N_1978,N_83);
and U5620 (N_5620,N_4829,N_4108);
nor U5621 (N_5621,N_4707,N_3748);
and U5622 (N_5622,N_1711,N_2955);
and U5623 (N_5623,N_4987,N_1180);
or U5624 (N_5624,N_4982,N_3412);
or U5625 (N_5625,N_1624,N_4027);
and U5626 (N_5626,N_4835,N_4430);
nand U5627 (N_5627,N_768,N_331);
or U5628 (N_5628,N_4037,N_3252);
xnor U5629 (N_5629,N_4176,N_2331);
and U5630 (N_5630,N_1335,N_1886);
and U5631 (N_5631,N_3813,N_3048);
nor U5632 (N_5632,N_4371,N_3795);
nor U5633 (N_5633,N_2535,N_2383);
and U5634 (N_5634,N_4815,N_1551);
xor U5635 (N_5635,N_2800,N_456);
or U5636 (N_5636,N_1433,N_32);
and U5637 (N_5637,N_2707,N_582);
and U5638 (N_5638,N_4640,N_462);
and U5639 (N_5639,N_3328,N_2368);
and U5640 (N_5640,N_885,N_2715);
and U5641 (N_5641,N_586,N_666);
nor U5642 (N_5642,N_418,N_2682);
or U5643 (N_5643,N_2342,N_3205);
nor U5644 (N_5644,N_2639,N_4615);
and U5645 (N_5645,N_1142,N_1748);
nand U5646 (N_5646,N_4441,N_441);
or U5647 (N_5647,N_1267,N_2728);
and U5648 (N_5648,N_374,N_165);
nor U5649 (N_5649,N_911,N_4458);
nand U5650 (N_5650,N_1281,N_1464);
nand U5651 (N_5651,N_1914,N_3535);
nand U5652 (N_5652,N_3010,N_1777);
xor U5653 (N_5653,N_1397,N_4471);
nor U5654 (N_5654,N_4574,N_794);
nor U5655 (N_5655,N_839,N_121);
and U5656 (N_5656,N_5,N_3225);
or U5657 (N_5657,N_1347,N_1743);
or U5658 (N_5658,N_2577,N_1933);
or U5659 (N_5659,N_4489,N_1467);
and U5660 (N_5660,N_1602,N_2982);
or U5661 (N_5661,N_1367,N_507);
nor U5662 (N_5662,N_530,N_4121);
nor U5663 (N_5663,N_4611,N_3317);
nand U5664 (N_5664,N_333,N_1939);
or U5665 (N_5665,N_263,N_748);
or U5666 (N_5666,N_1405,N_951);
nor U5667 (N_5667,N_607,N_2537);
or U5668 (N_5668,N_1330,N_450);
nand U5669 (N_5669,N_4883,N_1158);
nor U5670 (N_5670,N_2744,N_4650);
or U5671 (N_5671,N_1238,N_3920);
nor U5672 (N_5672,N_4508,N_4518);
nand U5673 (N_5673,N_4304,N_3923);
and U5674 (N_5674,N_4461,N_3719);
xor U5675 (N_5675,N_2352,N_4249);
xnor U5676 (N_5676,N_2275,N_1930);
and U5677 (N_5677,N_1288,N_4725);
nor U5678 (N_5678,N_534,N_2501);
or U5679 (N_5679,N_291,N_1214);
nor U5680 (N_5680,N_1033,N_2891);
and U5681 (N_5681,N_1006,N_2294);
and U5682 (N_5682,N_1213,N_754);
and U5683 (N_5683,N_4722,N_1793);
xnor U5684 (N_5684,N_4584,N_635);
nor U5685 (N_5685,N_1016,N_1702);
nand U5686 (N_5686,N_3194,N_1887);
nor U5687 (N_5687,N_102,N_3687);
xor U5688 (N_5688,N_3294,N_1609);
nand U5689 (N_5689,N_4893,N_4281);
nor U5690 (N_5690,N_4089,N_3954);
nor U5691 (N_5691,N_4642,N_2818);
or U5692 (N_5692,N_4488,N_3157);
nand U5693 (N_5693,N_1215,N_1389);
and U5694 (N_5694,N_1574,N_644);
or U5695 (N_5695,N_2607,N_3822);
or U5696 (N_5696,N_3539,N_2235);
xor U5697 (N_5697,N_3107,N_3406);
and U5698 (N_5698,N_4513,N_113);
nand U5699 (N_5699,N_4980,N_2670);
or U5700 (N_5700,N_511,N_548);
and U5701 (N_5701,N_2797,N_918);
and U5702 (N_5702,N_4460,N_3988);
nand U5703 (N_5703,N_2640,N_274);
xor U5704 (N_5704,N_2502,N_1579);
nor U5705 (N_5705,N_3638,N_1160);
or U5706 (N_5706,N_1816,N_2269);
or U5707 (N_5707,N_4177,N_846);
and U5708 (N_5708,N_1457,N_1220);
or U5709 (N_5709,N_3320,N_3169);
nand U5710 (N_5710,N_3196,N_2895);
nor U5711 (N_5711,N_4059,N_3778);
nor U5712 (N_5712,N_4072,N_1573);
nand U5713 (N_5713,N_4570,N_4504);
or U5714 (N_5714,N_2042,N_4789);
nor U5715 (N_5715,N_4794,N_1273);
nand U5716 (N_5716,N_94,N_628);
and U5717 (N_5717,N_923,N_3459);
or U5718 (N_5718,N_2329,N_1720);
or U5719 (N_5719,N_1957,N_3323);
nand U5720 (N_5720,N_1611,N_2243);
or U5721 (N_5721,N_1754,N_2330);
nor U5722 (N_5722,N_1910,N_3982);
nand U5723 (N_5723,N_2449,N_2145);
or U5724 (N_5724,N_1448,N_1924);
nor U5725 (N_5725,N_1919,N_3561);
nor U5726 (N_5726,N_3008,N_2688);
nor U5727 (N_5727,N_4372,N_4074);
nand U5728 (N_5728,N_1946,N_1963);
or U5729 (N_5729,N_1549,N_4763);
and U5730 (N_5730,N_1462,N_1789);
nor U5731 (N_5731,N_132,N_925);
nor U5732 (N_5732,N_1046,N_1796);
and U5733 (N_5733,N_4433,N_1558);
xnor U5734 (N_5734,N_2878,N_750);
and U5735 (N_5735,N_0,N_4097);
or U5736 (N_5736,N_1880,N_3537);
nand U5737 (N_5737,N_3248,N_2276);
and U5738 (N_5738,N_3361,N_921);
nand U5739 (N_5739,N_128,N_4797);
nor U5740 (N_5740,N_4258,N_3662);
nor U5741 (N_5741,N_3880,N_4415);
nor U5742 (N_5742,N_2029,N_419);
nor U5743 (N_5743,N_857,N_4434);
and U5744 (N_5744,N_4667,N_3534);
and U5745 (N_5745,N_1384,N_2133);
nor U5746 (N_5746,N_3311,N_2867);
or U5747 (N_5747,N_964,N_2463);
nor U5748 (N_5748,N_1025,N_2215);
nor U5749 (N_5749,N_141,N_4306);
nand U5750 (N_5750,N_4359,N_3765);
or U5751 (N_5751,N_2832,N_2677);
nand U5752 (N_5752,N_3508,N_2387);
or U5753 (N_5753,N_3147,N_4301);
nand U5754 (N_5754,N_1209,N_2016);
or U5755 (N_5755,N_1670,N_42);
and U5756 (N_5756,N_1271,N_2641);
or U5757 (N_5757,N_3394,N_4844);
nor U5758 (N_5758,N_1082,N_2144);
nand U5759 (N_5759,N_4239,N_89);
nor U5760 (N_5760,N_499,N_2146);
and U5761 (N_5761,N_359,N_871);
nor U5762 (N_5762,N_4948,N_4131);
or U5763 (N_5763,N_4221,N_4509);
nand U5764 (N_5764,N_4492,N_1353);
or U5765 (N_5765,N_2270,N_2055);
and U5766 (N_5766,N_2978,N_1644);
or U5767 (N_5767,N_343,N_4119);
nand U5768 (N_5768,N_2123,N_1884);
nor U5769 (N_5769,N_1874,N_110);
nor U5770 (N_5770,N_2686,N_166);
nand U5771 (N_5771,N_3610,N_753);
and U5772 (N_5772,N_2212,N_3557);
and U5773 (N_5773,N_2453,N_4698);
nand U5774 (N_5774,N_4713,N_4530);
or U5775 (N_5775,N_3867,N_3919);
and U5776 (N_5776,N_2087,N_2803);
or U5777 (N_5777,N_724,N_1413);
nand U5778 (N_5778,N_1550,N_152);
nor U5779 (N_5779,N_814,N_1470);
and U5780 (N_5780,N_410,N_4100);
or U5781 (N_5781,N_2763,N_2109);
and U5782 (N_5782,N_4162,N_234);
and U5783 (N_5783,N_1764,N_2174);
nor U5784 (N_5784,N_3313,N_728);
xnor U5785 (N_5785,N_3538,N_3100);
xnor U5786 (N_5786,N_4167,N_1197);
or U5787 (N_5787,N_830,N_3253);
xor U5788 (N_5788,N_2177,N_4873);
nand U5789 (N_5789,N_2810,N_4740);
and U5790 (N_5790,N_2692,N_851);
xnor U5791 (N_5791,N_1048,N_2260);
and U5792 (N_5792,N_3693,N_3583);
and U5793 (N_5793,N_4702,N_1123);
xor U5794 (N_5794,N_90,N_2717);
nor U5795 (N_5795,N_2238,N_4062);
or U5796 (N_5796,N_2062,N_4989);
or U5797 (N_5797,N_1251,N_3493);
nor U5798 (N_5798,N_698,N_2161);
and U5799 (N_5799,N_1023,N_255);
xor U5800 (N_5800,N_2965,N_2907);
and U5801 (N_5801,N_3288,N_4709);
xor U5802 (N_5802,N_3783,N_45);
nor U5803 (N_5803,N_3505,N_3332);
or U5804 (N_5804,N_4860,N_3942);
nand U5805 (N_5805,N_1055,N_4419);
nand U5806 (N_5806,N_2722,N_547);
nor U5807 (N_5807,N_2143,N_2527);
xnor U5808 (N_5808,N_140,N_2020);
nor U5809 (N_5809,N_3680,N_2918);
nor U5810 (N_5810,N_373,N_3015);
nor U5811 (N_5811,N_3273,N_1019);
or U5812 (N_5812,N_2007,N_2082);
xor U5813 (N_5813,N_3609,N_4387);
and U5814 (N_5814,N_1715,N_543);
or U5815 (N_5815,N_938,N_1431);
and U5816 (N_5816,N_3575,N_1092);
nor U5817 (N_5817,N_388,N_2037);
or U5818 (N_5818,N_3860,N_4044);
nand U5819 (N_5819,N_3714,N_1740);
and U5820 (N_5820,N_2376,N_4903);
nor U5821 (N_5821,N_3395,N_4684);
or U5822 (N_5822,N_447,N_2990);
xor U5823 (N_5823,N_4510,N_1432);
and U5824 (N_5824,N_1757,N_2090);
nand U5825 (N_5825,N_1841,N_4402);
or U5826 (N_5826,N_575,N_1926);
nand U5827 (N_5827,N_1047,N_564);
or U5828 (N_5828,N_4971,N_3868);
nor U5829 (N_5829,N_993,N_1488);
and U5830 (N_5830,N_1867,N_4427);
or U5831 (N_5831,N_3758,N_55);
or U5832 (N_5832,N_2608,N_514);
xnor U5833 (N_5833,N_3522,N_2452);
and U5834 (N_5834,N_1727,N_2858);
nand U5835 (N_5835,N_1208,N_1681);
xnor U5836 (N_5836,N_4586,N_2959);
xor U5837 (N_5837,N_357,N_3843);
nor U5838 (N_5838,N_2250,N_4912);
nor U5839 (N_5839,N_546,N_4242);
or U5840 (N_5840,N_2635,N_2963);
or U5841 (N_5841,N_2288,N_827);
and U5842 (N_5842,N_656,N_116);
nor U5843 (N_5843,N_1649,N_3737);
and U5844 (N_5844,N_4814,N_2077);
nor U5845 (N_5845,N_4798,N_2905);
xnor U5846 (N_5846,N_3944,N_183);
or U5847 (N_5847,N_1618,N_3373);
nand U5848 (N_5848,N_3222,N_4726);
nor U5849 (N_5849,N_420,N_3053);
nor U5850 (N_5850,N_302,N_1059);
nor U5851 (N_5851,N_663,N_4422);
nand U5852 (N_5852,N_2375,N_3624);
and U5853 (N_5853,N_4613,N_4603);
or U5854 (N_5854,N_1074,N_3353);
or U5855 (N_5855,N_394,N_282);
or U5856 (N_5856,N_761,N_4708);
xnor U5857 (N_5857,N_4720,N_424);
nand U5858 (N_5858,N_4654,N_1291);
or U5859 (N_5859,N_2191,N_1322);
nand U5860 (N_5860,N_2261,N_2523);
xor U5861 (N_5861,N_2986,N_1556);
or U5862 (N_5862,N_4438,N_4522);
nand U5863 (N_5863,N_4233,N_4699);
xnor U5864 (N_5864,N_3742,N_1986);
nand U5865 (N_5865,N_4063,N_3892);
or U5866 (N_5866,N_959,N_2497);
or U5867 (N_5867,N_4106,N_1888);
nand U5868 (N_5868,N_1385,N_660);
or U5869 (N_5869,N_865,N_3259);
nand U5870 (N_5870,N_417,N_849);
nand U5871 (N_5871,N_1768,N_1749);
or U5872 (N_5872,N_2655,N_284);
and U5873 (N_5873,N_2347,N_3779);
nand U5874 (N_5874,N_3608,N_3180);
or U5875 (N_5875,N_4404,N_3718);
nor U5876 (N_5876,N_218,N_267);
and U5877 (N_5877,N_2927,N_652);
xnor U5878 (N_5878,N_3012,N_4378);
and U5879 (N_5879,N_4030,N_2869);
or U5880 (N_5880,N_992,N_300);
nor U5881 (N_5881,N_745,N_11);
nand U5882 (N_5882,N_2381,N_3595);
and U5883 (N_5883,N_1275,N_3356);
nor U5884 (N_5884,N_2468,N_2127);
nand U5885 (N_5885,N_430,N_3396);
and U5886 (N_5886,N_1507,N_114);
nand U5887 (N_5887,N_734,N_4927);
and U5888 (N_5888,N_2684,N_3432);
or U5889 (N_5889,N_1026,N_2396);
nor U5890 (N_5890,N_1137,N_4041);
and U5891 (N_5891,N_3556,N_4900);
nor U5892 (N_5892,N_1126,N_3106);
and U5893 (N_5893,N_401,N_365);
nand U5894 (N_5894,N_4017,N_1369);
nor U5895 (N_5895,N_1168,N_2720);
nand U5896 (N_5896,N_825,N_185);
nand U5897 (N_5897,N_1265,N_4678);
nand U5898 (N_5898,N_2718,N_1721);
and U5899 (N_5899,N_3883,N_501);
nor U5900 (N_5900,N_1854,N_1893);
nor U5901 (N_5901,N_2070,N_3666);
nand U5902 (N_5902,N_802,N_524);
nand U5903 (N_5903,N_4436,N_4414);
and U5904 (N_5904,N_3363,N_808);
xor U5905 (N_5905,N_4352,N_1756);
nand U5906 (N_5906,N_3464,N_1022);
and U5907 (N_5907,N_449,N_3852);
xor U5908 (N_5908,N_1420,N_77);
nand U5909 (N_5909,N_1879,N_1762);
or U5910 (N_5910,N_975,N_2795);
nand U5911 (N_5911,N_2582,N_3728);
and U5912 (N_5912,N_1145,N_4852);
nor U5913 (N_5913,N_3151,N_1419);
xor U5914 (N_5914,N_2751,N_1247);
nor U5915 (N_5915,N_1004,N_2719);
and U5916 (N_5916,N_2182,N_1424);
nand U5917 (N_5917,N_3530,N_4457);
nand U5918 (N_5918,N_3333,N_574);
xor U5919 (N_5919,N_693,N_2064);
xnor U5920 (N_5920,N_4810,N_1763);
and U5921 (N_5921,N_912,N_1530);
and U5922 (N_5922,N_1922,N_2361);
nor U5923 (N_5923,N_4090,N_2945);
or U5924 (N_5924,N_4187,N_4150);
or U5925 (N_5925,N_1440,N_2230);
or U5926 (N_5926,N_569,N_2382);
or U5927 (N_5927,N_4412,N_344);
and U5928 (N_5928,N_3145,N_4367);
nor U5929 (N_5929,N_4916,N_1819);
or U5930 (N_5930,N_4663,N_623);
or U5931 (N_5931,N_4552,N_1090);
and U5932 (N_5932,N_2454,N_1333);
and U5933 (N_5933,N_1805,N_403);
or U5934 (N_5934,N_4105,N_2284);
nor U5935 (N_5935,N_277,N_2804);
nand U5936 (N_5936,N_428,N_2216);
and U5937 (N_5937,N_4424,N_312);
and U5938 (N_5938,N_2129,N_2371);
nand U5939 (N_5939,N_3546,N_4170);
or U5940 (N_5940,N_2902,N_3835);
nor U5941 (N_5941,N_358,N_1913);
nand U5942 (N_5942,N_872,N_4443);
xnor U5943 (N_5943,N_820,N_4571);
or U5944 (N_5944,N_1834,N_1791);
nand U5945 (N_5945,N_1814,N_2826);
nand U5946 (N_5946,N_647,N_1182);
and U5947 (N_5947,N_880,N_1403);
or U5948 (N_5948,N_2052,N_4452);
nor U5949 (N_5949,N_4550,N_2786);
nand U5950 (N_5950,N_2638,N_1582);
or U5951 (N_5951,N_3447,N_3756);
nand U5952 (N_5952,N_144,N_1020);
nand U5953 (N_5953,N_860,N_3391);
nor U5954 (N_5954,N_2370,N_910);
or U5955 (N_5955,N_1456,N_1730);
nor U5956 (N_5956,N_1766,N_43);
xnor U5957 (N_5957,N_4656,N_1141);
nor U5958 (N_5958,N_1,N_1216);
xnor U5959 (N_5959,N_2262,N_3774);
nand U5960 (N_5960,N_1250,N_4186);
nand U5961 (N_5961,N_49,N_2282);
or U5962 (N_5962,N_2499,N_3726);
and U5963 (N_5963,N_2505,N_2461);
nand U5964 (N_5964,N_3204,N_922);
and U5965 (N_5965,N_4937,N_1717);
nand U5966 (N_5966,N_3187,N_2925);
and U5967 (N_5967,N_3782,N_3451);
or U5968 (N_5968,N_2822,N_2006);
nor U5969 (N_5969,N_4356,N_4040);
nand U5970 (N_5970,N_2734,N_4786);
xor U5971 (N_5971,N_4132,N_1057);
nor U5972 (N_5972,N_196,N_1452);
or U5973 (N_5973,N_1152,N_3958);
nor U5974 (N_5974,N_3642,N_86);
and U5975 (N_5975,N_59,N_2465);
nand U5976 (N_5976,N_3025,N_301);
and U5977 (N_5977,N_4014,N_3081);
nand U5978 (N_5978,N_998,N_4834);
xor U5979 (N_5979,N_2069,N_730);
or U5980 (N_5980,N_1665,N_52);
nor U5981 (N_5981,N_3940,N_2056);
and U5982 (N_5982,N_2756,N_601);
or U5983 (N_5983,N_4318,N_2456);
nand U5984 (N_5984,N_1490,N_645);
or U5985 (N_5985,N_4820,N_3611);
nor U5986 (N_5986,N_2672,N_649);
xnor U5987 (N_5987,N_3897,N_4228);
or U5988 (N_5988,N_2296,N_888);
xor U5989 (N_5989,N_2224,N_1891);
and U5990 (N_5990,N_4871,N_2455);
and U5991 (N_5991,N_1371,N_4970);
nand U5992 (N_5992,N_4464,N_1635);
and U5993 (N_5993,N_2252,N_3397);
xnor U5994 (N_5994,N_2023,N_363);
xor U5995 (N_5995,N_3378,N_870);
nand U5996 (N_5996,N_3854,N_2764);
nor U5997 (N_5997,N_3231,N_429);
or U5998 (N_5998,N_4716,N_594);
nand U5999 (N_5999,N_1853,N_3794);
and U6000 (N_6000,N_2876,N_2833);
nand U6001 (N_6001,N_3414,N_3722);
or U6002 (N_6002,N_4894,N_3077);
or U6003 (N_6003,N_485,N_2633);
or U6004 (N_6004,N_2674,N_4525);
nand U6005 (N_6005,N_4398,N_1905);
or U6006 (N_6006,N_4651,N_3489);
nand U6007 (N_6007,N_442,N_3513);
and U6008 (N_6008,N_4328,N_1694);
nand U6009 (N_6009,N_725,N_3371);
xnor U6010 (N_6010,N_3979,N_1284);
nand U6011 (N_6011,N_276,N_228);
or U6012 (N_6012,N_4021,N_4099);
and U6013 (N_6013,N_1317,N_837);
and U6014 (N_6014,N_641,N_4711);
nor U6015 (N_6015,N_4045,N_4750);
or U6016 (N_6016,N_4481,N_2121);
and U6017 (N_6017,N_205,N_1491);
or U6018 (N_6018,N_3789,N_2420);
nor U6019 (N_6019,N_270,N_1688);
nand U6020 (N_6020,N_895,N_2814);
nor U6021 (N_6021,N_2950,N_2612);
and U6022 (N_6022,N_4734,N_467);
or U6023 (N_6023,N_3099,N_4854);
and U6024 (N_6024,N_2757,N_3267);
nand U6025 (N_6025,N_4976,N_2731);
nor U6026 (N_6026,N_4913,N_4769);
nand U6027 (N_6027,N_705,N_4954);
nand U6028 (N_6028,N_1627,N_3613);
nor U6029 (N_6029,N_1229,N_1842);
and U6030 (N_6030,N_4775,N_62);
and U6031 (N_6031,N_1050,N_3862);
and U6032 (N_6032,N_2080,N_1146);
or U6033 (N_6033,N_482,N_4056);
xnor U6034 (N_6034,N_1993,N_1755);
or U6035 (N_6035,N_4218,N_63);
nand U6036 (N_6036,N_3429,N_4737);
and U6037 (N_6037,N_1099,N_3937);
nor U6038 (N_6038,N_1205,N_3354);
nand U6039 (N_6039,N_3193,N_1010);
or U6040 (N_6040,N_3082,N_439);
nor U6041 (N_6041,N_453,N_483);
or U6042 (N_6042,N_4715,N_3300);
or U6043 (N_6043,N_898,N_257);
xnor U6044 (N_6044,N_392,N_1775);
and U6045 (N_6045,N_4212,N_478);
xor U6046 (N_6046,N_970,N_4983);
nand U6047 (N_6047,N_2208,N_145);
nor U6048 (N_6048,N_650,N_1298);
nand U6049 (N_6049,N_4171,N_2572);
nor U6050 (N_6050,N_1818,N_2526);
or U6051 (N_6051,N_4754,N_3885);
nor U6052 (N_6052,N_2745,N_498);
nor U6053 (N_6053,N_2911,N_3683);
or U6054 (N_6054,N_3094,N_1176);
and U6055 (N_6055,N_3781,N_2410);
or U6056 (N_6056,N_842,N_324);
nand U6057 (N_6057,N_2436,N_1234);
or U6058 (N_6058,N_3498,N_1784);
nand U6059 (N_6059,N_3529,N_2541);
nor U6060 (N_6060,N_3098,N_603);
or U6061 (N_6061,N_2097,N_3708);
nand U6062 (N_6062,N_4549,N_1093);
nor U6063 (N_6063,N_2748,N_3902);
or U6064 (N_6064,N_4107,N_2017);
or U6065 (N_6065,N_3946,N_3991);
and U6066 (N_6066,N_250,N_3669);
nor U6067 (N_6067,N_1072,N_1856);
or U6068 (N_6068,N_4085,N_3415);
and U6069 (N_6069,N_2237,N_3032);
nor U6070 (N_6070,N_4051,N_2167);
or U6071 (N_6071,N_2437,N_4996);
and U6072 (N_6072,N_4392,N_493);
or U6073 (N_6073,N_4399,N_3230);
nor U6074 (N_6074,N_4691,N_4759);
or U6075 (N_6075,N_1340,N_3786);
nor U6076 (N_6076,N_4755,N_244);
or U6077 (N_6077,N_3011,N_696);
xnor U6078 (N_6078,N_4824,N_2706);
and U6079 (N_6079,N_366,N_2882);
nand U6080 (N_6080,N_309,N_491);
or U6081 (N_6081,N_1300,N_4123);
nor U6082 (N_6082,N_3083,N_4467);
nor U6083 (N_6083,N_4183,N_1811);
nor U6084 (N_6084,N_1958,N_4007);
and U6085 (N_6085,N_3154,N_939);
nor U6086 (N_6086,N_1545,N_4364);
or U6087 (N_6087,N_3972,N_126);
and U6088 (N_6088,N_2571,N_4224);
or U6089 (N_6089,N_4911,N_2628);
nor U6090 (N_6090,N_1174,N_3501);
and U6091 (N_6091,N_2584,N_4001);
nor U6092 (N_6092,N_1870,N_3007);
xnor U6093 (N_6093,N_1643,N_1383);
or U6094 (N_6094,N_1065,N_863);
xor U6095 (N_6095,N_4995,N_2289);
or U6096 (N_6096,N_2324,N_2438);
xnor U6097 (N_6097,N_3507,N_4115);
and U6098 (N_6098,N_606,N_233);
xor U6099 (N_6099,N_226,N_706);
and U6100 (N_6100,N_381,N_4114);
nand U6101 (N_6101,N_4054,N_4676);
nor U6102 (N_6102,N_2654,N_4665);
nand U6103 (N_6103,N_3564,N_3206);
nand U6104 (N_6104,N_3518,N_3804);
nor U6105 (N_6105,N_3091,N_3303);
nor U6106 (N_6106,N_3520,N_3287);
and U6107 (N_6107,N_1127,N_3840);
nor U6108 (N_6108,N_266,N_3033);
or U6109 (N_6109,N_3072,N_1697);
xor U6110 (N_6110,N_1780,N_989);
nand U6111 (N_6111,N_1478,N_395);
and U6112 (N_6112,N_4350,N_2266);
nand U6113 (N_6113,N_251,N_1484);
and U6114 (N_6114,N_1566,N_437);
xnor U6115 (N_6115,N_659,N_2594);
nand U6116 (N_6116,N_1262,N_3698);
nand U6117 (N_6117,N_2780,N_2012);
and U6118 (N_6118,N_2951,N_4134);
nor U6119 (N_6119,N_2279,N_1593);
nand U6120 (N_6120,N_3241,N_4619);
and U6121 (N_6121,N_1953,N_412);
or U6122 (N_6122,N_805,N_4141);
or U6123 (N_6123,N_433,N_4562);
nand U6124 (N_6124,N_4445,N_4144);
nor U6125 (N_6125,N_3980,N_4943);
nand U6126 (N_6126,N_1248,N_1622);
nor U6127 (N_6127,N_2460,N_61);
nor U6128 (N_6128,N_598,N_4519);
nand U6129 (N_6129,N_4137,N_592);
or U6130 (N_6130,N_1096,N_60);
nand U6131 (N_6131,N_142,N_1726);
nor U6132 (N_6132,N_3027,N_1441);
and U6133 (N_6133,N_3955,N_3700);
and U6134 (N_6134,N_854,N_4338);
nand U6135 (N_6135,N_4695,N_3970);
nor U6136 (N_6136,N_4048,N_576);
or U6137 (N_6137,N_2098,N_4189);
nand U6138 (N_6138,N_4881,N_1513);
or U6139 (N_6139,N_2327,N_1725);
nor U6140 (N_6140,N_2337,N_1489);
and U6141 (N_6141,N_315,N_1231);
nor U6142 (N_6142,N_1532,N_3585);
nand U6143 (N_6143,N_2248,N_1927);
and U6144 (N_6144,N_3652,N_451);
xnor U6145 (N_6145,N_2546,N_3149);
nand U6146 (N_6146,N_4207,N_4349);
xnor U6147 (N_6147,N_1438,N_2412);
or U6148 (N_6148,N_3648,N_1132);
nor U6149 (N_6149,N_2490,N_3472);
nor U6150 (N_6150,N_1129,N_1529);
or U6151 (N_6151,N_1166,N_2588);
or U6152 (N_6152,N_1679,N_3992);
xor U6153 (N_6153,N_3445,N_4547);
or U6154 (N_6154,N_1169,N_1479);
nor U6155 (N_6155,N_2530,N_4802);
nor U6156 (N_6156,N_252,N_4474);
nand U6157 (N_6157,N_2693,N_2551);
nand U6158 (N_6158,N_3586,N_4738);
and U6159 (N_6159,N_4933,N_3292);
or U6160 (N_6160,N_733,N_699);
and U6161 (N_6161,N_1712,N_2393);
or U6162 (N_6162,N_1992,N_1646);
xor U6163 (N_6163,N_4673,N_1645);
or U6164 (N_6164,N_4830,N_2419);
or U6165 (N_6165,N_1171,N_4377);
and U6166 (N_6166,N_4361,N_2139);
or U6167 (N_6167,N_4203,N_3703);
and U6168 (N_6168,N_3280,N_1586);
and U6169 (N_6169,N_2574,N_2322);
nand U6170 (N_6170,N_1972,N_2772);
nand U6171 (N_6171,N_3260,N_4145);
or U6172 (N_6172,N_3830,N_1458);
nand U6173 (N_6173,N_3383,N_4113);
nor U6174 (N_6174,N_2619,N_3038);
or U6175 (N_6175,N_3704,N_1772);
nand U6176 (N_6176,N_3842,N_411);
and U6177 (N_6177,N_3350,N_4354);
nand U6178 (N_6178,N_3615,N_2831);
nor U6179 (N_6179,N_4480,N_181);
nand U6180 (N_6180,N_2316,N_4052);
nor U6181 (N_6181,N_777,N_760);
nor U6182 (N_6182,N_843,N_3882);
and U6183 (N_6183,N_3598,N_1117);
and U6184 (N_6184,N_4949,N_960);
and U6185 (N_6185,N_4608,N_3284);
nor U6186 (N_6186,N_4324,N_3893);
and U6187 (N_6187,N_350,N_781);
and U6188 (N_6188,N_3441,N_1967);
or U6189 (N_6189,N_4080,N_2310);
nor U6190 (N_6190,N_4406,N_3798);
nor U6191 (N_6191,N_4291,N_3894);
and U6192 (N_6192,N_1098,N_2893);
nand U6193 (N_6193,N_1561,N_53);
and U6194 (N_6194,N_769,N_2532);
nor U6195 (N_6195,N_3960,N_1382);
and U6196 (N_6196,N_4209,N_2081);
or U6197 (N_6197,N_1184,N_2922);
nand U6198 (N_6198,N_108,N_1575);
nor U6199 (N_6199,N_4965,N_703);
nand U6200 (N_6200,N_2820,N_551);
or U6201 (N_6201,N_3661,N_1287);
or U6202 (N_6202,N_1991,N_2286);
nor U6203 (N_6203,N_4577,N_3747);
nand U6204 (N_6204,N_1352,N_446);
or U6205 (N_6205,N_1081,N_2379);
nor U6206 (N_6206,N_4921,N_4511);
or U6207 (N_6207,N_1009,N_3495);
and U6208 (N_6208,N_3884,N_2225);
or U6209 (N_6209,N_2071,N_3924);
or U6210 (N_6210,N_908,N_3189);
nor U6211 (N_6211,N_3234,N_3913);
nor U6212 (N_6212,N_2613,N_2039);
and U6213 (N_6213,N_713,N_4885);
nor U6214 (N_6214,N_2152,N_796);
or U6215 (N_6215,N_2738,N_4950);
nor U6216 (N_6216,N_4323,N_1085);
xor U6217 (N_6217,N_952,N_590);
nand U6218 (N_6218,N_4346,N_4543);
nor U6219 (N_6219,N_3023,N_799);
and U6220 (N_6220,N_4154,N_1001);
nand U6221 (N_6221,N_4036,N_2168);
or U6222 (N_6222,N_2837,N_572);
xor U6223 (N_6223,N_2473,N_4483);
and U6224 (N_6224,N_2915,N_2072);
nor U6225 (N_6225,N_4521,N_518);
xor U6226 (N_6226,N_946,N_3995);
and U6227 (N_6227,N_3407,N_3536);
nor U6228 (N_6228,N_1400,N_4420);
nor U6229 (N_6229,N_223,N_375);
and U6230 (N_6230,N_2032,N_999);
nor U6231 (N_6231,N_4869,N_160);
or U6232 (N_6232,N_1154,N_2560);
or U6233 (N_6233,N_3735,N_3519);
and U6234 (N_6234,N_2267,N_2457);
or U6235 (N_6235,N_150,N_2514);
nor U6236 (N_6236,N_4015,N_1683);
nand U6237 (N_6237,N_3061,N_2611);
and U6238 (N_6238,N_4591,N_272);
nor U6239 (N_6239,N_894,N_3814);
xnor U6240 (N_6240,N_2104,N_475);
nand U6241 (N_6241,N_1007,N_3863);
and U6242 (N_6242,N_1056,N_103);
nor U6243 (N_6243,N_3422,N_788);
xor U6244 (N_6244,N_2994,N_81);
and U6245 (N_6245,N_3837,N_4800);
nor U6246 (N_6246,N_3497,N_2219);
and U6247 (N_6247,N_448,N_4638);
and U6248 (N_6248,N_1439,N_625);
xnor U6249 (N_6249,N_1863,N_3904);
xnor U6250 (N_6250,N_1409,N_1285);
nor U6251 (N_6251,N_3912,N_3509);
nand U6252 (N_6252,N_2536,N_360);
and U6253 (N_6253,N_3660,N_474);
and U6254 (N_6254,N_4256,N_3653);
xnor U6255 (N_6255,N_801,N_1078);
nand U6256 (N_6256,N_3279,N_3876);
and U6257 (N_6257,N_2500,N_899);
nand U6258 (N_6258,N_201,N_1598);
and U6259 (N_6259,N_4271,N_3068);
and U6260 (N_6260,N_4394,N_3657);
xnor U6261 (N_6261,N_763,N_1202);
and U6262 (N_6262,N_3952,N_1037);
xor U6263 (N_6263,N_1153,N_3918);
nor U6264 (N_6264,N_661,N_2249);
or U6265 (N_6265,N_3793,N_4895);
nor U6266 (N_6266,N_2721,N_3172);
and U6267 (N_6267,N_2755,N_2431);
nand U6268 (N_6268,N_3334,N_1990);
or U6269 (N_6269,N_2019,N_1787);
nor U6270 (N_6270,N_957,N_4390);
nand U6271 (N_6271,N_4333,N_4589);
and U6272 (N_6272,N_4523,N_2119);
and U6273 (N_6273,N_1249,N_711);
nand U6274 (N_6274,N_727,N_1560);
and U6275 (N_6275,N_4193,N_3132);
xnor U6276 (N_6276,N_3431,N_367);
xnor U6277 (N_6277,N_2958,N_2259);
and U6278 (N_6278,N_1562,N_1264);
or U6279 (N_6279,N_714,N_2462);
nand U6280 (N_6280,N_583,N_4572);
or U6281 (N_6281,N_3347,N_1851);
and U6282 (N_6282,N_882,N_2147);
or U6283 (N_6283,N_4453,N_2027);
nand U6284 (N_6284,N_3562,N_2678);
or U6285 (N_6285,N_2424,N_3668);
or U6286 (N_6286,N_2791,N_2778);
or U6287 (N_6287,N_520,N_791);
and U6288 (N_6288,N_2989,N_3741);
and U6289 (N_6289,N_4491,N_780);
and U6290 (N_6290,N_3998,N_2953);
nand U6291 (N_6291,N_1373,N_4253);
nor U6292 (N_6292,N_3908,N_3762);
nand U6293 (N_6293,N_3834,N_1921);
or U6294 (N_6294,N_70,N_488);
nor U6295 (N_6295,N_341,N_1103);
and U6296 (N_6296,N_3319,N_1667);
and U6297 (N_6297,N_3097,N_602);
nor U6298 (N_6298,N_342,N_3777);
or U6299 (N_6299,N_46,N_1434);
nand U6300 (N_6300,N_4868,N_2103);
and U6301 (N_6301,N_4714,N_1013);
nor U6302 (N_6302,N_2776,N_2852);
xnor U6303 (N_6303,N_1770,N_2353);
nor U6304 (N_6304,N_3725,N_2697);
xnor U6305 (N_6305,N_3983,N_976);
nor U6306 (N_6306,N_299,N_1839);
nor U6307 (N_6307,N_2443,N_4499);
and U6308 (N_6308,N_3715,N_3616);
or U6309 (N_6309,N_3997,N_613);
and U6310 (N_6310,N_2318,N_4826);
nand U6311 (N_6311,N_2705,N_744);
nor U6312 (N_6312,N_2244,N_3251);
nor U6313 (N_6313,N_3481,N_4303);
or U6314 (N_6314,N_3721,N_436);
nor U6315 (N_6315,N_297,N_279);
or U6316 (N_6316,N_1395,N_3746);
nand U6317 (N_6317,N_2779,N_1309);
nand U6318 (N_6318,N_1817,N_2078);
and U6319 (N_6319,N_2031,N_2467);
or U6320 (N_6320,N_219,N_2242);
and U6321 (N_6321,N_3933,N_1949);
or U6322 (N_6322,N_517,N_4853);
and U6323 (N_6323,N_662,N_3829);
nor U6324 (N_6324,N_3421,N_4537);
nand U6325 (N_6325,N_4962,N_674);
and U6326 (N_6326,N_4274,N_770);
xnor U6327 (N_6327,N_304,N_3387);
xnor U6328 (N_6328,N_4046,N_4244);
xor U6329 (N_6329,N_3593,N_308);
nand U6330 (N_6330,N_3699,N_1223);
or U6331 (N_6331,N_2162,N_2851);
xor U6332 (N_6332,N_1962,N_2843);
and U6333 (N_6333,N_3113,N_1450);
nand U6334 (N_6334,N_1310,N_3446);
and U6335 (N_6335,N_3528,N_4652);
or U6336 (N_6336,N_3148,N_4683);
nor U6337 (N_6337,N_3621,N_1399);
nor U6338 (N_6338,N_620,N_4986);
nand U6339 (N_6339,N_3226,N_4793);
nand U6340 (N_6340,N_93,N_1843);
or U6341 (N_6341,N_1542,N_4159);
nand U6342 (N_6342,N_1810,N_1364);
nand U6343 (N_6343,N_3410,N_4515);
or U6344 (N_6344,N_463,N_1741);
and U6345 (N_6345,N_1388,N_622);
nor U6346 (N_6346,N_3368,N_3018);
nor U6347 (N_6347,N_1404,N_3821);
or U6348 (N_6348,N_2935,N_541);
xnor U6349 (N_6349,N_979,N_1858);
xor U6350 (N_6350,N_1307,N_476);
and U6351 (N_6351,N_3851,N_1402);
and U6352 (N_6352,N_3064,N_4849);
xor U6353 (N_6353,N_4855,N_1412);
xor U6354 (N_6354,N_1524,N_3731);
nand U6355 (N_6355,N_1920,N_1638);
xnor U6356 (N_6356,N_3494,N_88);
and U6357 (N_6357,N_978,N_4863);
nor U6358 (N_6358,N_3209,N_2910);
or U6359 (N_6359,N_4284,N_1345);
or U6360 (N_6360,N_87,N_3701);
nor U6361 (N_6361,N_2923,N_57);
nor U6362 (N_6362,N_4744,N_4690);
nand U6363 (N_6363,N_2591,N_624);
and U6364 (N_6364,N_2232,N_2466);
xor U6365 (N_6365,N_1608,N_2493);
and U6366 (N_6366,N_1869,N_3186);
and U6367 (N_6367,N_1407,N_3754);
nand U6368 (N_6368,N_4355,N_3989);
or U6369 (N_6369,N_4828,N_2556);
and U6370 (N_6370,N_3037,N_4528);
nor U6371 (N_6371,N_3506,N_2083);
or U6372 (N_6372,N_2271,N_3914);
nand U6373 (N_6373,N_1320,N_2736);
and U6374 (N_6374,N_4011,N_1541);
xor U6375 (N_6375,N_199,N_1476);
or U6376 (N_6376,N_383,N_253);
nand U6377 (N_6377,N_1199,N_3296);
and U6378 (N_6378,N_4476,N_3679);
and U6379 (N_6379,N_4490,N_4487);
nand U6380 (N_6380,N_380,N_3475);
or U6381 (N_6381,N_2518,N_4920);
and U6382 (N_6382,N_1961,N_4779);
or U6383 (N_6383,N_4075,N_819);
and U6384 (N_6384,N_3131,N_585);
and U6385 (N_6385,N_3866,N_2345);
nor U6386 (N_6386,N_3381,N_686);
nand U6387 (N_6387,N_2061,N_3846);
and U6388 (N_6388,N_2906,N_3966);
nand U6389 (N_6389,N_36,N_2196);
or U6390 (N_6390,N_3672,N_1492);
xnor U6391 (N_6391,N_285,N_4315);
and U6392 (N_6392,N_3664,N_2898);
xnor U6393 (N_6393,N_3644,N_2947);
nor U6394 (N_6394,N_3974,N_3712);
nor U6395 (N_6395,N_242,N_741);
or U6396 (N_6396,N_560,N_96);
nor U6397 (N_6397,N_22,N_1283);
and U6398 (N_6398,N_3824,N_1596);
and U6399 (N_6399,N_1555,N_3805);
nand U6400 (N_6400,N_4919,N_1116);
and U6401 (N_6401,N_1316,N_2492);
nor U6402 (N_6402,N_3342,N_2849);
or U6403 (N_6403,N_4721,N_1883);
and U6404 (N_6404,N_3800,N_2614);
or U6405 (N_6405,N_1983,N_1170);
or U6406 (N_6406,N_452,N_3729);
and U6407 (N_6407,N_2589,N_4669);
nand U6408 (N_6408,N_2760,N_3078);
nand U6409 (N_6409,N_4752,N_3678);
nor U6410 (N_6410,N_4593,N_3930);
nand U6411 (N_6411,N_2338,N_3129);
nand U6412 (N_6412,N_1435,N_3916);
nand U6413 (N_6413,N_4357,N_4944);
and U6414 (N_6414,N_3402,N_4110);
nor U6415 (N_6415,N_3002,N_2899);
nor U6416 (N_6416,N_774,N_56);
nand U6417 (N_6417,N_2794,N_2010);
or U6418 (N_6418,N_743,N_3079);
xor U6419 (N_6419,N_614,N_153);
nand U6420 (N_6420,N_169,N_2340);
and U6421 (N_6421,N_4770,N_2647);
nor U6422 (N_6422,N_4229,N_3744);
and U6423 (N_6423,N_4706,N_3130);
nor U6424 (N_6424,N_1526,N_1516);
xnor U6425 (N_6425,N_2542,N_2036);
and U6426 (N_6426,N_1592,N_1620);
xor U6427 (N_6427,N_626,N_1410);
nor U6428 (N_6428,N_3605,N_1114);
or U6429 (N_6429,N_3062,N_4727);
nand U6430 (N_6430,N_1094,N_3250);
nor U6431 (N_6431,N_3957,N_1354);
nand U6432 (N_6432,N_4307,N_3216);
and U6433 (N_6433,N_3628,N_2190);
and U6434 (N_6434,N_2857,N_2566);
nand U6435 (N_6435,N_2297,N_4599);
or U6436 (N_6436,N_3499,N_2314);
or U6437 (N_6437,N_4555,N_723);
nor U6438 (N_6438,N_1246,N_4329);
nand U6439 (N_6439,N_3977,N_3461);
nor U6440 (N_6440,N_1398,N_4216);
nor U6441 (N_6441,N_2481,N_3764);
nor U6442 (N_6442,N_1274,N_2491);
xor U6443 (N_6443,N_2305,N_700);
and U6444 (N_6444,N_4120,N_2176);
nand U6445 (N_6445,N_4248,N_1865);
nor U6446 (N_6446,N_1370,N_2180);
or U6447 (N_6447,N_3457,N_3239);
and U6448 (N_6448,N_664,N_718);
xor U6449 (N_6449,N_2274,N_2149);
xnor U6450 (N_6450,N_1535,N_2850);
and U6451 (N_6451,N_969,N_1282);
xnor U6452 (N_6452,N_4351,N_4149);
and U6453 (N_6453,N_1706,N_2652);
xnor U6454 (N_6454,N_2630,N_58);
nand U6455 (N_6455,N_2914,N_1164);
xnor U6456 (N_6456,N_3797,N_1017);
nand U6457 (N_6457,N_2725,N_902);
or U6458 (N_6458,N_3673,N_3975);
nor U6459 (N_6459,N_2509,N_2422);
and U6460 (N_6460,N_4151,N_1318);
nor U6461 (N_6461,N_2447,N_3026);
and U6462 (N_6462,N_812,N_2003);
nor U6463 (N_6463,N_627,N_306);
nor U6464 (N_6464,N_3602,N_4066);
or U6465 (N_6465,N_328,N_1809);
nand U6466 (N_6466,N_2350,N_3922);
or U6467 (N_6467,N_3543,N_4641);
nor U6468 (N_6468,N_4439,N_2970);
or U6469 (N_6469,N_170,N_1718);
nand U6470 (N_6470,N_762,N_3247);
nand U6471 (N_6471,N_4264,N_2844);
or U6472 (N_6472,N_12,N_1937);
nand U6473 (N_6473,N_658,N_729);
nor U6474 (N_6474,N_687,N_2565);
or U6475 (N_6475,N_3567,N_2665);
nor U6476 (N_6476,N_1449,N_384);
nand U6477 (N_6477,N_868,N_3763);
or U6478 (N_6478,N_742,N_4002);
nand U6479 (N_6479,N_3379,N_3521);
or U6480 (N_6480,N_3208,N_4403);
nor U6481 (N_6481,N_3619,N_3297);
nand U6482 (N_6482,N_1311,N_349);
and U6483 (N_6483,N_3993,N_3671);
nand U6484 (N_6484,N_1258,N_3238);
nand U6485 (N_6485,N_3694,N_1942);
or U6486 (N_6486,N_2096,N_1985);
or U6487 (N_6487,N_4396,N_338);
or U6488 (N_6488,N_2369,N_4268);
nor U6489 (N_6489,N_4277,N_1613);
or U6490 (N_6490,N_4267,N_371);
and U6491 (N_6491,N_2813,N_4825);
nor U6492 (N_6492,N_2698,N_3676);
and U6493 (N_6493,N_208,N_4111);
or U6494 (N_6494,N_280,N_1929);
or U6495 (N_6495,N_612,N_2221);
nor U6496 (N_6496,N_120,N_1537);
nor U6497 (N_6497,N_4060,N_1195);
nand U6498 (N_6498,N_709,N_906);
or U6499 (N_6499,N_1860,N_1331);
nand U6500 (N_6500,N_3291,N_532);
nor U6501 (N_6501,N_3874,N_3890);
xnor U6502 (N_6502,N_2685,N_2974);
nor U6503 (N_6503,N_472,N_4818);
nor U6504 (N_6504,N_1583,N_4649);
nand U6505 (N_6505,N_3374,N_457);
nor U6506 (N_6506,N_1895,N_4205);
nand U6507 (N_6507,N_4857,N_1401);
nor U6508 (N_6508,N_3815,N_778);
nand U6509 (N_6509,N_186,N_1533);
nor U6510 (N_6510,N_1528,N_1700);
or U6511 (N_6511,N_4269,N_4157);
or U6512 (N_6512,N_4838,N_4751);
or U6513 (N_6513,N_355,N_3134);
xnor U6514 (N_6514,N_3524,N_2099);
nand U6515 (N_6515,N_3767,N_1087);
nor U6516 (N_6516,N_4602,N_4103);
nor U6517 (N_6517,N_3337,N_1641);
or U6518 (N_6518,N_3651,N_3844);
nand U6519 (N_6519,N_1089,N_4473);
xor U6520 (N_6520,N_1671,N_2030);
nand U6521 (N_6521,N_3438,N_2434);
or U6522 (N_6522,N_3326,N_3850);
xnor U6523 (N_6523,N_3462,N_4985);
nor U6524 (N_6524,N_3588,N_3785);
nor U6525 (N_6525,N_1150,N_4411);
nor U6526 (N_6526,N_1734,N_4450);
nand U6527 (N_6527,N_2916,N_3973);
or U6528 (N_6528,N_3227,N_987);
xor U6529 (N_6529,N_995,N_2873);
or U6530 (N_6530,N_3881,N_2701);
or U6531 (N_6531,N_2131,N_2409);
or U6532 (N_6532,N_4288,N_4749);
or U6533 (N_6533,N_3544,N_4538);
nor U6534 (N_6534,N_4767,N_4548);
nor U6535 (N_6535,N_994,N_719);
nor U6536 (N_6536,N_1786,N_3269);
xor U6537 (N_6537,N_4703,N_259);
or U6538 (N_6538,N_2973,N_3278);
xnor U6539 (N_6539,N_327,N_2120);
and U6540 (N_6540,N_1106,N_2186);
xnor U6541 (N_6541,N_3075,N_4208);
or U6542 (N_6542,N_549,N_2516);
and U6543 (N_6543,N_934,N_2610);
nor U6544 (N_6544,N_3845,N_897);
nand U6545 (N_6545,N_4426,N_665);
nand U6546 (N_6546,N_2754,N_4093);
and U6547 (N_6547,N_100,N_822);
and U6548 (N_6548,N_1201,N_3455);
and U6549 (N_6549,N_1125,N_4875);
nor U6550 (N_6550,N_236,N_1102);
nor U6551 (N_6551,N_2723,N_2179);
nand U6552 (N_6552,N_1684,N_2140);
or U6553 (N_6553,N_1296,N_2470);
nand U6554 (N_6554,N_1797,N_3052);
xnor U6555 (N_6555,N_4146,N_4061);
and U6556 (N_6556,N_673,N_4172);
xnor U6557 (N_6557,N_1585,N_3198);
or U6558 (N_6558,N_3849,N_1204);
nand U6559 (N_6559,N_2335,N_716);
or U6560 (N_6560,N_3385,N_4173);
or U6561 (N_6561,N_3144,N_1135);
and U6562 (N_6562,N_2239,N_3322);
nor U6563 (N_6563,N_2257,N_2164);
and U6564 (N_6564,N_4416,N_2411);
and U6565 (N_6565,N_290,N_2999);
or U6566 (N_6566,N_1844,N_2687);
and U6567 (N_6567,N_4034,N_4337);
and U6568 (N_6568,N_616,N_1783);
nor U6569 (N_6569,N_2366,N_4601);
nand U6570 (N_6570,N_3416,N_26);
and U6571 (N_6571,N_1245,N_815);
or U6572 (N_6572,N_3087,N_2562);
or U6573 (N_6573,N_736,N_4185);
xnor U6574 (N_6574,N_787,N_4421);
and U6575 (N_6575,N_351,N_988);
nand U6576 (N_6576,N_2084,N_2425);
nor U6577 (N_6577,N_2689,N_1606);
nor U6578 (N_6578,N_2642,N_2992);
or U6579 (N_6579,N_3456,N_2615);
or U6580 (N_6580,N_4029,N_792);
nand U6581 (N_6581,N_2806,N_2617);
nor U6582 (N_6582,N_4653,N_2737);
and U6583 (N_6583,N_3014,N_785);
and U6584 (N_6584,N_615,N_4516);
and U6585 (N_6585,N_1062,N_2583);
and U6586 (N_6586,N_2406,N_4645);
nor U6587 (N_6587,N_1473,N_4425);
nor U6588 (N_6588,N_320,N_2661);
nand U6589 (N_6589,N_3448,N_766);
and U6590 (N_6590,N_1095,N_4385);
or U6591 (N_6591,N_3047,N_2278);
nor U6592 (N_6592,N_3121,N_4050);
and U6593 (N_6593,N_1411,N_2234);
nand U6594 (N_6594,N_1804,N_4463);
nand U6595 (N_6595,N_3040,N_3161);
or U6596 (N_6596,N_1503,N_2901);
nand U6597 (N_6597,N_2092,N_237);
nand U6598 (N_6598,N_195,N_1588);
and U6599 (N_6599,N_2827,N_1653);
and U6600 (N_6600,N_2427,N_707);
xnor U6601 (N_6601,N_776,N_2676);
and U6602 (N_6602,N_1987,N_980);
nor U6603 (N_6603,N_2446,N_1034);
and U6604 (N_6604,N_3776,N_425);
or U6605 (N_6605,N_1477,N_2609);
xor U6606 (N_6606,N_260,N_4822);
xor U6607 (N_6607,N_3170,N_4073);
nor U6608 (N_6608,N_3926,N_783);
nand U6609 (N_6609,N_1833,N_4687);
or U6610 (N_6610,N_522,N_3423);
xor U6611 (N_6611,N_4977,N_3436);
nand U6612 (N_6612,N_4503,N_3486);
nor U6613 (N_6613,N_2178,N_1655);
and U6614 (N_6614,N_1232,N_3341);
and U6615 (N_6615,N_903,N_2050);
nand U6616 (N_6616,N_389,N_864);
or U6617 (N_6617,N_738,N_1559);
and U6618 (N_6618,N_4742,N_4214);
nand U6619 (N_6619,N_4785,N_519);
nand U6620 (N_6620,N_4005,N_4606);
and U6621 (N_6621,N_4276,N_4605);
xor U6622 (N_6622,N_2471,N_1124);
or U6623 (N_6623,N_3895,N_2320);
or U6624 (N_6624,N_397,N_4945);
and U6625 (N_6625,N_1736,N_1514);
or U6626 (N_6626,N_3525,N_875);
xor U6627 (N_6627,N_2533,N_2835);
and U6628 (N_6628,N_752,N_256);
nor U6629 (N_6629,N_4255,N_3314);
nand U6630 (N_6630,N_1303,N_670);
nand U6631 (N_6631,N_941,N_2317);
xor U6632 (N_6632,N_4316,N_3111);
or U6633 (N_6633,N_772,N_481);
nand U6634 (N_6634,N_4196,N_2290);
nand U6635 (N_6635,N_1820,N_1128);
and U6636 (N_6636,N_241,N_1342);
and U6637 (N_6637,N_4363,N_2210);
xor U6638 (N_6638,N_3367,N_4870);
or U6639 (N_6639,N_4373,N_1722);
nor U6640 (N_6640,N_4138,N_4942);
xnor U6641 (N_6641,N_1188,N_2644);
and U6642 (N_6642,N_4559,N_347);
nand U6643 (N_6643,N_2246,N_3454);
nor U6644 (N_6644,N_4343,N_431);
or U6645 (N_6645,N_1003,N_3357);
xor U6646 (N_6646,N_2014,N_4275);
nand U6647 (N_6647,N_3965,N_4314);
nand U6648 (N_6648,N_913,N_1315);
nand U6649 (N_6649,N_2333,N_1442);
nor U6650 (N_6650,N_2254,N_3706);
nand U6651 (N_6651,N_4733,N_3617);
or U6652 (N_6652,N_2889,N_2846);
xor U6653 (N_6653,N_4493,N_2351);
and U6654 (N_6654,N_795,N_2529);
or U6655 (N_6655,N_4477,N_1143);
xnor U6656 (N_6656,N_4250,N_2564);
nor U6657 (N_6657,N_146,N_3069);
nor U6658 (N_6658,N_1838,N_4563);
or U6659 (N_6659,N_3355,N_4886);
and U6660 (N_6660,N_3120,N_852);
and U6661 (N_6661,N_3891,N_4672);
nand U6662 (N_6662,N_4305,N_1278);
nor U6663 (N_6663,N_1682,N_4918);
nand U6664 (N_6664,N_732,N_3554);
and U6665 (N_6665,N_599,N_1505);
and U6666 (N_6666,N_2539,N_2859);
or U6667 (N_6667,N_3587,N_489);
xor U6668 (N_6668,N_4922,N_1885);
nand U6669 (N_6669,N_2865,N_264);
nor U6670 (N_6670,N_4161,N_305);
nor U6671 (N_6671,N_66,N_4535);
nand U6672 (N_6672,N_3791,N_3139);
and U6673 (N_6673,N_3517,N_3095);
and U6674 (N_6674,N_3945,N_4102);
and U6675 (N_6675,N_3601,N_4375);
and U6676 (N_6676,N_840,N_4578);
xor U6677 (N_6677,N_3709,N_4520);
nand U6678 (N_6678,N_4235,N_4067);
or U6679 (N_6679,N_1207,N_2399);
nand U6680 (N_6680,N_2931,N_3290);
xor U6681 (N_6681,N_2554,N_4077);
or U6682 (N_6682,N_1523,N_4575);
and U6683 (N_6683,N_2066,N_3847);
nand U6684 (N_6684,N_1878,N_1416);
or U6685 (N_6685,N_4639,N_3017);
and U6686 (N_6686,N_3386,N_254);
nand U6687 (N_6687,N_2163,N_246);
or U6688 (N_6688,N_3178,N_3086);
nand U6689 (N_6689,N_3710,N_2277);
nand U6690 (N_6690,N_3000,N_2426);
and U6691 (N_6691,N_4008,N_1795);
nor U6692 (N_6692,N_2590,N_2919);
and U6693 (N_6693,N_3986,N_2624);
and U6694 (N_6694,N_4813,N_3887);
and U6695 (N_6695,N_372,N_314);
nor U6696 (N_6696,N_3312,N_4472);
and U6697 (N_6697,N_869,N_2074);
and U6698 (N_6698,N_1107,N_215);
and U6699 (N_6699,N_3167,N_2998);
nand U6700 (N_6700,N_3366,N_847);
nand U6701 (N_6701,N_4199,N_4604);
nand U6702 (N_6702,N_3713,N_845);
and U6703 (N_6703,N_3921,N_526);
nor U6704 (N_6704,N_3634,N_4567);
nand U6705 (N_6705,N_1835,N_4662);
or U6706 (N_6706,N_2306,N_1509);
nor U6707 (N_6707,N_1731,N_3909);
or U6708 (N_6708,N_67,N_1329);
nand U6709 (N_6709,N_1547,N_1824);
and U6710 (N_6710,N_2478,N_2747);
or U6711 (N_6711,N_3630,N_1332);
nor U6712 (N_6712,N_3199,N_4087);
and U6713 (N_6713,N_1021,N_4851);
nor U6714 (N_6714,N_2134,N_248);
nand U6715 (N_6715,N_2506,N_3905);
and U6716 (N_6716,N_73,N_2022);
nand U6717 (N_6717,N_14,N_2480);
and U6718 (N_6718,N_570,N_1705);
xnor U6719 (N_6719,N_2172,N_1443);
nor U6720 (N_6720,N_1161,N_3213);
or U6721 (N_6721,N_4540,N_1446);
nand U6722 (N_6722,N_3275,N_3743);
and U6723 (N_6723,N_3142,N_4969);
nand U6724 (N_6724,N_1252,N_3409);
xnor U6725 (N_6725,N_4320,N_3752);
and U6726 (N_6726,N_4756,N_2432);
or U6727 (N_6727,N_1219,N_4251);
or U6728 (N_6728,N_27,N_1691);
and U6729 (N_6729,N_4821,N_2009);
xor U6730 (N_6730,N_2900,N_1601);
nor U6731 (N_6731,N_2629,N_1767);
xor U6732 (N_6732,N_4630,N_2202);
and U6733 (N_6733,N_1292,N_4391);
or U6734 (N_6734,N_2769,N_2115);
nand U6735 (N_6735,N_1156,N_471);
nor U6736 (N_6736,N_1928,N_3853);
or U6737 (N_6737,N_1186,N_3769);
and U6738 (N_6738,N_2952,N_765);
nand U6739 (N_6739,N_1902,N_1429);
or U6740 (N_6740,N_919,N_2553);
nor U6741 (N_6741,N_1828,N_1534);
nor U6742 (N_6742,N_3030,N_1710);
or U6743 (N_6743,N_3968,N_393);
nand U6744 (N_6744,N_3114,N_4991);
and U6745 (N_6745,N_2108,N_2928);
nor U6746 (N_6746,N_117,N_1859);
and U6747 (N_6747,N_2875,N_4261);
nand U6748 (N_6748,N_1954,N_4236);
or U6749 (N_6749,N_172,N_2785);
xnor U6750 (N_6750,N_848,N_1510);
nand U6751 (N_6751,N_997,N_2004);
nand U6752 (N_6752,N_759,N_2765);
or U6753 (N_6753,N_4446,N_559);
and U6754 (N_6754,N_877,N_4104);
and U6755 (N_6755,N_3138,N_1280);
and U6756 (N_6756,N_618,N_177);
nand U6757 (N_6757,N_1890,N_675);
and U6758 (N_6758,N_1218,N_949);
nor U6759 (N_6759,N_1483,N_1286);
nand U6760 (N_6760,N_3858,N_3309);
nor U6761 (N_6761,N_4990,N_326);
nand U6762 (N_6762,N_2605,N_2341);
nand U6763 (N_6763,N_1414,N_4409);
and U6764 (N_6764,N_3809,N_3655);
and U6765 (N_6765,N_4561,N_2984);
nor U6766 (N_6766,N_4500,N_164);
xor U6767 (N_6767,N_4968,N_296);
or U6768 (N_6768,N_1632,N_2660);
nor U6769 (N_6769,N_2209,N_2401);
or U6770 (N_6770,N_1105,N_4783);
nor U6771 (N_6771,N_1968,N_2985);
or U6772 (N_6772,N_1941,N_4071);
or U6773 (N_6773,N_1076,N_2228);
nand U6774 (N_6774,N_779,N_1889);
nor U6775 (N_6775,N_3787,N_1071);
or U6776 (N_6776,N_3790,N_4782);
xor U6777 (N_6777,N_125,N_1459);
nor U6778 (N_6778,N_3310,N_3344);
nor U6779 (N_6779,N_2187,N_4447);
nor U6780 (N_6780,N_4807,N_311);
and U6781 (N_6781,N_2729,N_2439);
and U6782 (N_6782,N_4994,N_230);
or U6783 (N_6783,N_1616,N_4761);
or U6784 (N_6784,N_2445,N_933);
nand U6785 (N_6785,N_1876,N_1657);
nor U6786 (N_6786,N_2855,N_1633);
nor U6787 (N_6787,N_2759,N_914);
nor U6788 (N_6788,N_4666,N_101);
nor U6789 (N_6789,N_2185,N_3886);
xor U6790 (N_6790,N_1911,N_217);
or U6791 (N_6791,N_3705,N_3418);
or U6792 (N_6792,N_1605,N_3559);
nor U6793 (N_6793,N_4925,N_4905);
or U6794 (N_6794,N_2433,N_2838);
nor U6795 (N_6795,N_1595,N_502);
or U6796 (N_6796,N_3390,N_1677);
nor U6797 (N_6797,N_1206,N_3304);
or U6798 (N_6798,N_3990,N_4070);
xnor U6799 (N_6799,N_3364,N_2694);
or U6800 (N_6800,N_1068,N_134);
nor U6801 (N_6801,N_1341,N_2740);
nand U6802 (N_6802,N_1363,N_2302);
or U6803 (N_6803,N_3685,N_828);
or U6804 (N_6804,N_4295,N_632);
or U6805 (N_6805,N_4801,N_1032);
or U6806 (N_6806,N_97,N_1295);
xnor U6807 (N_6807,N_95,N_3643);
and U6808 (N_6808,N_789,N_874);
or U6809 (N_6809,N_4505,N_4109);
xnor U6810 (N_6810,N_492,N_4897);
and U6811 (N_6811,N_2118,N_545);
and U6812 (N_6812,N_1052,N_3377);
nand U6813 (N_6813,N_3750,N_2125);
or U6814 (N_6814,N_4201,N_3085);
xor U6815 (N_6815,N_2981,N_920);
nand U6816 (N_6816,N_1366,N_229);
nand U6817 (N_6817,N_2775,N_4024);
and U6818 (N_6818,N_3614,N_510);
and U6819 (N_6819,N_112,N_2991);
nand U6820 (N_6820,N_4541,N_1378);
or U6821 (N_6821,N_1110,N_1704);
and U6822 (N_6822,N_608,N_422);
nand U6823 (N_6823,N_1293,N_2386);
nand U6824 (N_6824,N_136,N_862);
nand U6825 (N_6825,N_2961,N_2417);
nand U6826 (N_6826,N_813,N_4636);
nor U6827 (N_6827,N_4444,N_4031);
xor U6828 (N_6828,N_1305,N_1539);
or U6829 (N_6829,N_2085,N_737);
and U6830 (N_6830,N_2128,N_3571);
or U6831 (N_6831,N_28,N_1894);
or U6832 (N_6832,N_15,N_3502);
nor U6833 (N_6833,N_695,N_936);
nor U6834 (N_6834,N_24,N_4257);
and U6835 (N_6835,N_3941,N_3483);
or U6836 (N_6836,N_3632,N_1177);
xor U6837 (N_6837,N_1134,N_2880);
or U6838 (N_6838,N_1995,N_1709);
nor U6839 (N_6839,N_1938,N_4932);
or U6840 (N_6840,N_2201,N_271);
nand U6841 (N_6841,N_916,N_1060);
or U6842 (N_6842,N_3675,N_2547);
or U6843 (N_6843,N_2380,N_3119);
nand U6844 (N_6844,N_1080,N_2913);
and U6845 (N_6845,N_2872,N_3570);
xor U6846 (N_6846,N_4998,N_1172);
xnor U6847 (N_6847,N_3900,N_3302);
or U6848 (N_6848,N_1301,N_1049);
or U6849 (N_6849,N_2709,N_1830);
xor U6850 (N_6850,N_2567,N_1376);
xor U6851 (N_6851,N_3191,N_2997);
and U6852 (N_6852,N_2117,N_2815);
nor U6853 (N_6853,N_3487,N_2198);
nand U6854 (N_6854,N_931,N_3258);
nor U6855 (N_6855,N_3861,N_1792);
and U6856 (N_6856,N_4163,N_3090);
nor U6857 (N_6857,N_2976,N_4972);
xor U6858 (N_6858,N_262,N_2550);
or U6859 (N_6859,N_3803,N_2620);
nor U6860 (N_6860,N_749,N_2703);
and U6861 (N_6861,N_4475,N_3899);
nor U6862 (N_6862,N_3469,N_2934);
or U6863 (N_6863,N_480,N_2451);
nand U6864 (N_6864,N_3512,N_3612);
xnor U6865 (N_6865,N_6,N_438);
nor U6866 (N_6866,N_2195,N_3578);
nand U6867 (N_6867,N_4039,N_996);
and U6868 (N_6868,N_3697,N_2430);
and U6869 (N_6869,N_1029,N_1327);
or U6870 (N_6870,N_4845,N_708);
nand U6871 (N_6871,N_1861,N_512);
or U6872 (N_6872,N_3155,N_180);
nand U6873 (N_6873,N_2746,N_3055);
xnor U6874 (N_6874,N_3265,N_2921);
and U6875 (N_6875,N_435,N_4265);
and U6876 (N_6876,N_278,N_1603);
nor U6877 (N_6877,N_1660,N_2743);
nor U6878 (N_6878,N_3636,N_127);
nor U6879 (N_6879,N_2586,N_1543);
and U6880 (N_6880,N_3428,N_4339);
xor U6881 (N_6881,N_423,N_407);
nand U6882 (N_6882,N_161,N_3569);
nand U6883 (N_6883,N_167,N_3360);
and U6884 (N_6884,N_786,N_3141);
or U6885 (N_6885,N_173,N_4936);
nor U6886 (N_6886,N_157,N_2418);
nor U6887 (N_6887,N_2464,N_947);
nor U6888 (N_6888,N_124,N_2489);
and U6889 (N_6889,N_1418,N_2076);
xor U6890 (N_6890,N_2291,N_107);
nand U6891 (N_6891,N_1338,N_3463);
or U6892 (N_6892,N_2107,N_4332);
and U6893 (N_6893,N_4622,N_3859);
or U6894 (N_6894,N_1498,N_4334);
nor U6895 (N_6895,N_4245,N_346);
or U6896 (N_6896,N_2159,N_4879);
nor U6897 (N_6897,N_1396,N_2909);
and U6898 (N_6898,N_2966,N_1192);
xnor U6899 (N_6899,N_1761,N_2181);
nand U6900 (N_6900,N_13,N_3146);
or U6901 (N_6901,N_1041,N_4042);
nor U6902 (N_6902,N_4628,N_4437);
or U6903 (N_6903,N_2742,N_688);
xor U6904 (N_6904,N_1719,N_2265);
and U6905 (N_6905,N_655,N_3331);
nand U6906 (N_6906,N_133,N_2753);
nand U6907 (N_6907,N_3807,N_1716);
xor U6908 (N_6908,N_1650,N_3542);
and U6909 (N_6909,N_3663,N_4202);
nor U6910 (N_6910,N_633,N_2513);
xor U6911 (N_6911,N_2273,N_2930);
nand U6912 (N_6912,N_2339,N_571);
and U6913 (N_6913,N_1390,N_2408);
or U6914 (N_6914,N_4778,N_1591);
nand U6915 (N_6915,N_954,N_4898);
and U6916 (N_6916,N_690,N_2649);
or U6917 (N_6917,N_4682,N_2158);
or U6918 (N_6918,N_3190,N_2413);
or U6919 (N_6919,N_974,N_555);
nand U6920 (N_6920,N_4746,N_184);
nand U6921 (N_6921,N_3228,N_2494);
or U6922 (N_6922,N_1737,N_1515);
nor U6923 (N_6923,N_2203,N_2679);
xnor U6924 (N_6924,N_1994,N_2241);
nor U6925 (N_6925,N_4592,N_3545);
or U6926 (N_6926,N_2980,N_2222);
or U6927 (N_6927,N_3400,N_515);
nor U6928 (N_6928,N_3577,N_2773);
and U6929 (N_6929,N_3816,N_1328);
and U6930 (N_6930,N_2936,N_1359);
xor U6931 (N_6931,N_1113,N_4410);
and U6932 (N_6932,N_4506,N_2968);
nor U6933 (N_6933,N_4981,N_4128);
and U6934 (N_6934,N_4175,N_4924);
nor U6935 (N_6935,N_1365,N_3994);
nor U6936 (N_6936,N_1778,N_2604);
or U6937 (N_6937,N_3325,N_4147);
and U6938 (N_6938,N_2598,N_2155);
nand U6939 (N_6939,N_4081,N_390);
nor U6940 (N_6940,N_398,N_2887);
nand U6941 (N_6941,N_3224,N_4796);
or U6942 (N_6942,N_2877,N_405);
or U6943 (N_6943,N_1831,N_4083);
or U6944 (N_6944,N_629,N_2830);
nor U6945 (N_6945,N_2871,N_3870);
or U6946 (N_6946,N_3639,N_1997);
xor U6947 (N_6947,N_79,N_179);
or U6948 (N_6948,N_2528,N_967);
and U6949 (N_6949,N_3174,N_2038);
nor U6950 (N_6950,N_2848,N_4428);
nand U6951 (N_6951,N_504,N_1862);
xnor U6952 (N_6952,N_4423,N_2504);
xor U6953 (N_6953,N_1578,N_2157);
nor U6954 (N_6954,N_4395,N_1907);
or U6955 (N_6955,N_3165,N_1571);
nor U6956 (N_6956,N_340,N_2555);
nor U6957 (N_6957,N_3948,N_1687);
xnor U6958 (N_6958,N_4279,N_1493);
or U6959 (N_6959,N_2625,N_3102);
nand U6960 (N_6960,N_3492,N_1871);
nor U6961 (N_6961,N_4736,N_3738);
nand U6962 (N_6962,N_416,N_681);
or U6963 (N_6963,N_1230,N_4379);
nand U6964 (N_6964,N_3408,N_1517);
or U6965 (N_6965,N_2435,N_904);
or U6966 (N_6966,N_3005,N_1415);
and U6967 (N_6967,N_4842,N_3006);
or U6968 (N_6968,N_4136,N_2766);
nor U6969 (N_6969,N_1463,N_4226);
xor U6970 (N_6970,N_1339,N_174);
or U6971 (N_6971,N_720,N_4704);
nand U6972 (N_6972,N_4407,N_680);
xor U6973 (N_6973,N_694,N_1554);
and U6974 (N_6974,N_2646,N_4065);
nor U6975 (N_6975,N_621,N_4317);
nand U6976 (N_6976,N_4888,N_3869);
nor U6977 (N_6977,N_3934,N_4680);
or U6978 (N_6978,N_591,N_3759);
or U6979 (N_6979,N_4929,N_2334);
or U6980 (N_6980,N_3674,N_3838);
nand U6981 (N_6981,N_64,N_3515);
nand U6982 (N_6982,N_335,N_3999);
nand U6983 (N_6983,N_3380,N_2673);
and U6984 (N_6984,N_4660,N_1587);
nand U6985 (N_6985,N_2704,N_3476);
or U6986 (N_6986,N_1136,N_858);
or U6987 (N_6987,N_203,N_2394);
and U6988 (N_6988,N_2192,N_2823);
nand U6989 (N_6989,N_1898,N_669);
nand U6990 (N_6990,N_4787,N_1299);
nor U6991 (N_6991,N_4531,N_4741);
nor U6992 (N_6992,N_182,N_1629);
nor U6993 (N_6993,N_2101,N_4260);
or U6994 (N_6994,N_41,N_893);
xor U6995 (N_6995,N_317,N_3770);
nand U6996 (N_6996,N_3684,N_1149);
nor U6997 (N_6997,N_2487,N_4637);
and U6998 (N_6998,N_261,N_225);
and U6999 (N_6999,N_4882,N_2488);
nand U7000 (N_7000,N_982,N_667);
and U7001 (N_7001,N_2114,N_3143);
or U7002 (N_7002,N_1506,N_928);
nor U7003 (N_7003,N_4192,N_1826);
or U7004 (N_7004,N_983,N_1955);
and U7005 (N_7005,N_1977,N_1122);
nand U7006 (N_7006,N_3618,N_1701);
or U7007 (N_7007,N_3442,N_1306);
or U7008 (N_7008,N_1304,N_3568);
or U7009 (N_7009,N_2197,N_92);
nor U7010 (N_7010,N_3063,N_2057);
nand U7011 (N_7011,N_790,N_1086);
or U7012 (N_7012,N_1798,N_4246);
nor U7013 (N_7013,N_3692,N_3695);
xnor U7014 (N_7014,N_325,N_2510);
or U7015 (N_7015,N_1565,N_1790);
and U7016 (N_7016,N_2298,N_4588);
and U7017 (N_7017,N_2603,N_3282);
nand U7018 (N_7018,N_1375,N_432);
or U7019 (N_7019,N_4220,N_4867);
or U7020 (N_7020,N_4988,N_1674);
nor U7021 (N_7021,N_3046,N_3839);
and U7022 (N_7022,N_3262,N_3403);
nor U7023 (N_7023,N_1923,N_2053);
nor U7024 (N_7024,N_4200,N_1581);
and U7025 (N_7025,N_3036,N_3901);
nand U7026 (N_7026,N_577,N_1064);
xor U7027 (N_7027,N_927,N_2520);
or U7028 (N_7028,N_2726,N_610);
nand U7029 (N_7029,N_1801,N_2853);
nor U7030 (N_7030,N_2045,N_4847);
xnor U7031 (N_7031,N_2752,N_2200);
and U7032 (N_7032,N_1500,N_4238);
and U7033 (N_7033,N_1120,N_836);
or U7034 (N_7034,N_2739,N_3503);
and U7035 (N_7035,N_4400,N_2148);
nand U7036 (N_7036,N_1848,N_4930);
nor U7037 (N_7037,N_810,N_4241);
xnor U7038 (N_7038,N_2256,N_1002);
and U7039 (N_7039,N_2924,N_3315);
and U7040 (N_7040,N_3108,N_4300);
or U7041 (N_7041,N_3324,N_4032);
or U7042 (N_7042,N_3336,N_85);
or U7043 (N_7043,N_1337,N_1779);
or U7044 (N_7044,N_3953,N_2863);
or U7045 (N_7045,N_2548,N_1940);
or U7046 (N_7046,N_944,N_1408);
and U7047 (N_7047,N_4129,N_962);
and U7048 (N_7048,N_3551,N_3140);
nand U7049 (N_7049,N_4470,N_1308);
and U7050 (N_7050,N_379,N_3122);
nor U7051 (N_7051,N_4788,N_427);
xnor U7052 (N_7052,N_2570,N_676);
nand U7053 (N_7053,N_4910,N_477);
nor U7054 (N_7054,N_3971,N_3878);
nor U7055 (N_7055,N_516,N_1481);
nand U7056 (N_7056,N_3723,N_1008);
xor U7057 (N_7057,N_2957,N_3270);
or U7058 (N_7058,N_200,N_1899);
xor U7059 (N_7059,N_1658,N_3716);
xor U7060 (N_7060,N_1610,N_4884);
xnor U7061 (N_7061,N_1686,N_247);
nor U7062 (N_7062,N_4627,N_3566);
nor U7063 (N_7063,N_2856,N_3434);
and U7064 (N_7064,N_1039,N_4557);
or U7065 (N_7065,N_2658,N_2543);
nor U7066 (N_7066,N_1666,N_3911);
xor U7067 (N_7067,N_1751,N_1381);
nand U7068 (N_7068,N_683,N_3943);
nor U7069 (N_7069,N_4388,N_2377);
nor U7070 (N_7070,N_4204,N_4693);
nor U7071 (N_7071,N_3049,N_2188);
nand U7072 (N_7072,N_122,N_1067);
xnor U7073 (N_7073,N_4648,N_3855);
and U7074 (N_7074,N_377,N_3135);
nor U7075 (N_7075,N_29,N_3305);
nor U7076 (N_7076,N_1261,N_640);
and U7077 (N_7077,N_2223,N_4309);
xor U7078 (N_7078,N_4784,N_434);
nand U7079 (N_7079,N_2681,N_2398);
and U7080 (N_7080,N_3024,N_3724);
nor U7081 (N_7081,N_1474,N_2864);
xnor U7082 (N_7082,N_1636,N_4999);
and U7083 (N_7083,N_1782,N_4819);
nor U7084 (N_7084,N_1225,N_4964);
and U7085 (N_7085,N_1427,N_831);
nand U7086 (N_7086,N_3915,N_2861);
nand U7087 (N_7087,N_461,N_465);
nor U7088 (N_7088,N_294,N_2325);
nand U7089 (N_7089,N_4234,N_4448);
nand U7090 (N_7090,N_4496,N_554);
or U7091 (N_7091,N_3649,N_3727);
nand U7092 (N_7092,N_684,N_1664);
nand U7093 (N_7093,N_3812,N_797);
or U7094 (N_7094,N_1639,N_2771);
nor U7095 (N_7095,N_2600,N_3223);
and U7096 (N_7096,N_1217,N_3872);
nand U7097 (N_7097,N_1567,N_861);
nand U7098 (N_7098,N_3533,N_1568);
or U7099 (N_7099,N_4153,N_3956);
and U7100 (N_7100,N_454,N_1075);
nor U7101 (N_7101,N_268,N_2767);
nor U7102 (N_7102,N_2295,N_2824);
and U7103 (N_7103,N_4517,N_3833);
or U7104 (N_7104,N_3889,N_4383);
and U7105 (N_7105,N_3580,N_2105);
or U7106 (N_7106,N_2194,N_3749);
nand U7107 (N_7107,N_4558,N_3001);
or U7108 (N_7108,N_2713,N_597);
nor U7109 (N_7109,N_1236,N_2788);
and U7110 (N_7110,N_1729,N_1430);
xnor U7111 (N_7111,N_3471,N_3939);
or U7112 (N_7112,N_1244,N_3003);
nor U7113 (N_7113,N_3392,N_3192);
and U7114 (N_7114,N_3117,N_51);
or U7115 (N_7115,N_4227,N_3877);
nor U7116 (N_7116,N_2068,N_1564);
and U7117 (N_7117,N_4465,N_2304);
and U7118 (N_7118,N_2258,N_4655);
nor U7119 (N_7119,N_672,N_1872);
nand U7120 (N_7120,N_2263,N_1198);
nor U7121 (N_7121,N_2475,N_2749);
or U7122 (N_7122,N_2315,N_3817);
nor U7123 (N_7123,N_2349,N_2416);
nor U7124 (N_7124,N_4719,N_1769);
nand U7125 (N_7125,N_4376,N_3453);
nand U7126 (N_7126,N_3711,N_4926);
and U7127 (N_7127,N_4016,N_9);
xnor U7128 (N_7128,N_2005,N_756);
or U7129 (N_7129,N_378,N_3263);
nor U7130 (N_7130,N_829,N_4626);
or U7131 (N_7131,N_1599,N_2792);
and U7132 (N_7132,N_4532,N_4892);
or U7133 (N_7133,N_3589,N_4429);
or U7134 (N_7134,N_985,N_3286);
nand U7135 (N_7135,N_3070,N_1909);
nand U7136 (N_7136,N_3449,N_4068);
xor U7137 (N_7137,N_3210,N_2699);
or U7138 (N_7138,N_1024,N_118);
and U7139 (N_7139,N_834,N_109);
or U7140 (N_7140,N_2407,N_1594);
or U7141 (N_7141,N_1746,N_889);
nor U7142 (N_7142,N_4569,N_3466);
nor U7143 (N_7143,N_115,N_171);
xnor U7144 (N_7144,N_4576,N_4497);
nand U7145 (N_7145,N_4841,N_1750);
or U7146 (N_7146,N_2632,N_188);
or U7147 (N_7147,N_3757,N_1077);
and U7148 (N_7148,N_4486,N_2251);
and U7149 (N_7149,N_4213,N_977);
or U7150 (N_7150,N_2971,N_4459);
and U7151 (N_7151,N_2323,N_1960);
and U7152 (N_7152,N_3888,N_3951);
xor U7153 (N_7153,N_3760,N_3682);
nand U7154 (N_7154,N_3691,N_537);
nor U7155 (N_7155,N_197,N_1989);
and U7156 (N_7156,N_2616,N_3827);
and U7157 (N_7157,N_404,N_3590);
or U7158 (N_7158,N_4389,N_4899);
nand U7159 (N_7159,N_1436,N_2008);
and U7160 (N_7160,N_4182,N_4484);
xor U7161 (N_7161,N_2659,N_4197);
and U7162 (N_7162,N_4179,N_3720);
and U7163 (N_7163,N_4952,N_2067);
nand U7164 (N_7164,N_1584,N_4418);
and U7165 (N_7165,N_4166,N_981);
nor U7166 (N_7166,N_4811,N_4232);
nand U7167 (N_7167,N_2601,N_4915);
and U7168 (N_7168,N_4631,N_2048);
and U7169 (N_7169,N_566,N_2657);
or U7170 (N_7170,N_2912,N_2903);
and U7171 (N_7171,N_3631,N_4696);
or U7172 (N_7172,N_20,N_339);
and U7173 (N_7173,N_1799,N_3826);
or U7174 (N_7174,N_1548,N_2954);
or U7175 (N_7175,N_4909,N_2073);
or U7176 (N_7176,N_4023,N_7);
xor U7177 (N_7177,N_4022,N_3527);
or U7178 (N_7178,N_1642,N_72);
or U7179 (N_7179,N_881,N_4931);
nor U7180 (N_7180,N_3419,N_466);
nand U7181 (N_7181,N_2441,N_2034);
xnor U7182 (N_7182,N_269,N_2402);
nand U7183 (N_7183,N_198,N_3220);
xnor U7184 (N_7184,N_2592,N_3103);
or U7185 (N_7185,N_654,N_2415);
or U7186 (N_7186,N_4140,N_4064);
or U7187 (N_7187,N_286,N_4370);
and U7188 (N_7188,N_1637,N_2622);
and U7189 (N_7189,N_187,N_3963);
nor U7190 (N_7190,N_4184,N_841);
or U7191 (N_7191,N_689,N_2883);
or U7192 (N_7192,N_963,N_3623);
or U7193 (N_7193,N_726,N_319);
nand U7194 (N_7194,N_984,N_4657);
nand U7195 (N_7195,N_293,N_3775);
and U7196 (N_7196,N_4092,N_2593);
nor U7197 (N_7197,N_1144,N_1374);
nor U7198 (N_7198,N_2308,N_1652);
nor U7199 (N_7199,N_579,N_3437);
or U7200 (N_7200,N_224,N_859);
or U7201 (N_7201,N_2515,N_1735);
nand U7202 (N_7202,N_1847,N_2359);
xnor U7203 (N_7203,N_804,N_4833);
and U7204 (N_7204,N_2189,N_4866);
or U7205 (N_7205,N_1460,N_565);
nand U7206 (N_7206,N_1945,N_443);
or U7207 (N_7207,N_1455,N_1179);
or U7208 (N_7208,N_4805,N_1724);
nor U7209 (N_7209,N_3330,N_3177);
nand U7210 (N_7210,N_3768,N_3413);
nand U7211 (N_7211,N_2770,N_2423);
nor U7212 (N_7212,N_1759,N_1038);
xor U7213 (N_7213,N_3510,N_2364);
and U7214 (N_7214,N_1119,N_47);
nand U7215 (N_7215,N_2841,N_2557);
and U7216 (N_7216,N_1557,N_2962);
nand U7217 (N_7217,N_1881,N_1066);
and U7218 (N_7218,N_835,N_2888);
and U7219 (N_7219,N_2809,N_1781);
nor U7220 (N_7220,N_3985,N_991);
xnor U7221 (N_7221,N_3465,N_2758);
and U7222 (N_7222,N_3013,N_4766);
xor U7223 (N_7223,N_4247,N_3152);
or U7224 (N_7224,N_1999,N_135);
xnor U7225 (N_7225,N_4876,N_281);
or U7226 (N_7226,N_3202,N_4381);
or U7227 (N_7227,N_3825,N_313);
or U7228 (N_7228,N_1044,N_178);
or U7229 (N_7229,N_905,N_104);
nor U7230 (N_7230,N_3327,N_210);
xor U7231 (N_7231,N_1580,N_4967);
nor U7232 (N_7232,N_3650,N_1147);
or U7233 (N_7233,N_4808,N_1011);
and U7234 (N_7234,N_2283,N_1237);
or U7235 (N_7235,N_3928,N_4393);
and U7236 (N_7236,N_2018,N_4743);
nand U7237 (N_7237,N_4112,N_2311);
nor U7238 (N_7238,N_2440,N_3);
or U7239 (N_7239,N_856,N_4033);
nand U7240 (N_7240,N_3043,N_4957);
or U7241 (N_7241,N_1302,N_3640);
xor U7242 (N_7242,N_265,N_3073);
xnor U7243 (N_7243,N_4082,N_2205);
nor U7244 (N_7244,N_3932,N_1758);
xnor U7245 (N_7245,N_3504,N_503);
nor U7246 (N_7246,N_1873,N_369);
or U7247 (N_7247,N_588,N_4598);
xnor U7248 (N_7248,N_3171,N_2483);
nor U7249 (N_7249,N_1569,N_3175);
and U7250 (N_7250,N_2459,N_2664);
or U7251 (N_7251,N_3646,N_1499);
nand U7252 (N_7252,N_2777,N_1018);
nor U7253 (N_7253,N_3150,N_21);
nor U7254 (N_7254,N_3358,N_1932);
nor U7255 (N_7255,N_1344,N_3056);
or U7256 (N_7256,N_2890,N_1392);
nand U7257 (N_7257,N_2524,N_4512);
nand U7258 (N_7258,N_2110,N_4889);
nor U7259 (N_7259,N_1372,N_4374);
nand U7260 (N_7260,N_1183,N_2534);
nor U7261 (N_7261,N_2126,N_4009);
or U7262 (N_7262,N_1471,N_521);
or U7263 (N_7263,N_2648,N_2948);
xnor U7264 (N_7264,N_1175,N_1165);
nor U7265 (N_7265,N_4431,N_1979);
nor U7266 (N_7266,N_1621,N_1212);
and U7267 (N_7267,N_275,N_1346);
or U7268 (N_7268,N_2392,N_4956);
nand U7269 (N_7269,N_715,N_3268);
and U7270 (N_7270,N_3295,N_3219);
and U7271 (N_7271,N_2637,N_3318);
nor U7272 (N_7272,N_4620,N_4454);
or U7273 (N_7273,N_1654,N_3212);
or U7274 (N_7274,N_4272,N_3301);
nor U7275 (N_7275,N_1864,N_4675);
nand U7276 (N_7276,N_3532,N_2714);
and U7277 (N_7277,N_4237,N_4760);
and U7278 (N_7278,N_935,N_4958);
nor U7279 (N_7279,N_3910,N_1319);
xor U7280 (N_7280,N_2580,N_2319);
nor U7281 (N_7281,N_376,N_3066);
and U7282 (N_7282,N_4629,N_2367);
nand U7283 (N_7283,N_3773,N_2894);
nand U7284 (N_7284,N_4946,N_382);
nor U7285 (N_7285,N_3352,N_2448);
xor U7286 (N_7286,N_4590,N_3745);
and U7287 (N_7287,N_4679,N_76);
nor U7288 (N_7288,N_2724,N_2091);
nand U7289 (N_7289,N_2063,N_2783);
nor U7290 (N_7290,N_2028,N_596);
nor U7291 (N_7291,N_3755,N_4710);
nand U7292 (N_7292,N_289,N_4877);
nand U7293 (N_7293,N_1148,N_421);
nor U7294 (N_7294,N_4091,N_3625);
or U7295 (N_7295,N_1803,N_1343);
or U7296 (N_7296,N_458,N_3424);
and U7297 (N_7297,N_1713,N_3688);
nand U7298 (N_7298,N_1971,N_3293);
or U7299 (N_7299,N_3084,N_4960);
and U7300 (N_7300,N_4440,N_4308);
and U7301 (N_7301,N_2933,N_3574);
nor U7302 (N_7302,N_2522,N_2476);
or U7303 (N_7303,N_4126,N_2218);
nor U7304 (N_7304,N_1485,N_1813);
and U7305 (N_7305,N_194,N_855);
nor U7306 (N_7306,N_4133,N_4934);
nor U7307 (N_7307,N_2049,N_1662);
nor U7308 (N_7308,N_3467,N_1203);
and U7309 (N_7309,N_2979,N_4168);
or U7310 (N_7310,N_509,N_2285);
nand U7311 (N_7311,N_50,N_1387);
or U7312 (N_7312,N_937,N_1487);
or U7313 (N_7313,N_2041,N_3160);
nor U7314 (N_7314,N_2969,N_1623);
and U7315 (N_7315,N_2414,N_3873);
nand U7316 (N_7316,N_1015,N_1133);
and U7317 (N_7317,N_3801,N_953);
or U7318 (N_7318,N_3176,N_1042);
nand U7319 (N_7319,N_3028,N_4596);
or U7320 (N_7320,N_3808,N_3702);
nor U7321 (N_7321,N_2374,N_2634);
nor U7322 (N_7322,N_4536,N_2993);
and U7323 (N_7323,N_3936,N_2142);
or U7324 (N_7324,N_1159,N_4290);
or U7325 (N_7325,N_1698,N_2798);
and U7326 (N_7326,N_2712,N_4545);
nor U7327 (N_7327,N_258,N_2937);
nand U7328 (N_7328,N_4293,N_3799);
nor U7329 (N_7329,N_1349,N_3647);
nand U7330 (N_7330,N_4861,N_40);
nand U7331 (N_7331,N_3832,N_3819);
and U7332 (N_7332,N_533,N_1536);
or U7333 (N_7333,N_1975,N_1325);
and U7334 (N_7334,N_356,N_4086);
nand U7335 (N_7335,N_33,N_2429);
xnor U7336 (N_7336,N_4152,N_2183);
xor U7337 (N_7337,N_2559,N_3444);
nand U7338 (N_7338,N_4230,N_2618);
nor U7339 (N_7339,N_527,N_2132);
or U7340 (N_7340,N_4612,N_704);
xor U7341 (N_7341,N_3232,N_2932);
and U7342 (N_7342,N_4012,N_222);
and U7343 (N_7343,N_1969,N_37);
nor U7344 (N_7344,N_4055,N_631);
and U7345 (N_7345,N_2988,N_2821);
nand U7346 (N_7346,N_1393,N_4353);
nand U7347 (N_7347,N_2495,N_48);
or U7348 (N_7348,N_1269,N_821);
xor U7349 (N_7349,N_238,N_1101);
and U7350 (N_7350,N_3964,N_1773);
nand U7351 (N_7351,N_3050,N_2135);
and U7352 (N_7352,N_3865,N_3645);
and U7353 (N_7353,N_3696,N_1324);
and U7354 (N_7354,N_2946,N_1227);
and U7355 (N_7355,N_4270,N_3514);
or U7356 (N_7356,N_1211,N_496);
and U7357 (N_7357,N_4243,N_2281);
and U7358 (N_7358,N_2150,N_2829);
nor U7359 (N_7359,N_4020,N_2307);
or U7360 (N_7360,N_1235,N_2229);
or U7361 (N_7361,N_2231,N_557);
nor U7362 (N_7362,N_3526,N_1362);
nor U7363 (N_7363,N_4169,N_4790);
xor U7364 (N_7364,N_2153,N_159);
nor U7365 (N_7365,N_961,N_3109);
nand U7366 (N_7366,N_1825,N_154);
or U7367 (N_7367,N_1597,N_4718);
nor U7368 (N_7368,N_4993,N_2060);
nand U7369 (N_7369,N_2033,N_3450);
or U7370 (N_7370,N_4311,N_4692);
nor U7371 (N_7371,N_2602,N_3468);
or U7372 (N_7372,N_1903,N_4585);
and U7373 (N_7373,N_2220,N_4643);
nand U7374 (N_7374,N_3021,N_1157);
nor U7375 (N_7375,N_4010,N_2479);
nand U7376 (N_7376,N_4546,N_562);
and U7377 (N_7377,N_1453,N_2801);
and U7378 (N_7378,N_8,N_3689);
nor U7379 (N_7379,N_1604,N_1714);
or U7380 (N_7380,N_1676,N_3166);
and U7381 (N_7381,N_3123,N_4312);
or U7382 (N_7382,N_4417,N_4341);
or U7383 (N_7383,N_3104,N_2211);
or U7384 (N_7384,N_65,N_1377);
nand U7385 (N_7385,N_2782,N_249);
and U7386 (N_7386,N_4772,N_1012);
nor U7387 (N_7387,N_2484,N_3584);
and U7388 (N_7388,N_735,N_3266);
or U7389 (N_7389,N_4057,N_3540);
and U7390 (N_7390,N_345,N_3411);
or U7391 (N_7391,N_464,N_54);
or U7392 (N_7392,N_2498,N_2917);
nand U7393 (N_7393,N_3626,N_3482);
and U7394 (N_7394,N_3067,N_2680);
nand U7395 (N_7395,N_1189,N_816);
and U7396 (N_7396,N_4953,N_4644);
xor U7397 (N_7397,N_4623,N_2836);
or U7398 (N_7398,N_469,N_2540);
nand U7399 (N_7399,N_775,N_3772);
nor U7400 (N_7400,N_214,N_4764);
nand U7401 (N_7401,N_2874,N_2651);
nand U7402 (N_7402,N_4498,N_2938);
nor U7403 (N_7403,N_2173,N_2236);
or U7404 (N_7404,N_1163,N_4331);
nand U7405 (N_7405,N_3592,N_553);
nand U7406 (N_7406,N_189,N_220);
xor U7407 (N_7407,N_1553,N_1692);
xnor U7408 (N_7408,N_175,N_3059);
nor U7409 (N_7409,N_4799,N_4319);
or U7410 (N_7410,N_764,N_638);
and U7411 (N_7411,N_106,N_4671);
nand U7412 (N_7412,N_1647,N_3126);
and U7413 (N_7413,N_3907,N_879);
nand U7414 (N_7414,N_2762,N_4462);
or U7415 (N_7415,N_1589,N_2025);
nand U7416 (N_7416,N_231,N_1173);
nand U7417 (N_7417,N_4731,N_3949);
and U7418 (N_7418,N_2404,N_4198);
xor U7419 (N_7419,N_1918,N_3340);
and U7420 (N_7420,N_31,N_3961);
nand U7421 (N_7421,N_2508,N_415);
nand U7422 (N_7422,N_460,N_2626);
nor U7423 (N_7423,N_2939,N_3127);
and U7424 (N_7424,N_1445,N_4685);
and U7425 (N_7425,N_1615,N_2691);
xnor U7426 (N_7426,N_75,N_567);
nand U7427 (N_7427,N_3484,N_653);
and U7428 (N_7428,N_3399,N_4);
nor U7429 (N_7429,N_3458,N_3183);
nor U7430 (N_7430,N_1253,N_1931);
nor U7431 (N_7431,N_886,N_682);
nand U7432 (N_7432,N_2400,N_1552);
and U7433 (N_7433,N_809,N_2840);
and U7434 (N_7434,N_3039,N_2385);
or U7435 (N_7435,N_4600,N_3820);
xnor U7436 (N_7436,N_4812,N_2373);
or U7437 (N_7437,N_332,N_2079);
nor U7438 (N_7438,N_2886,N_25);
nor U7439 (N_7439,N_2093,N_4095);
and U7440 (N_7440,N_1112,N_3168);
nor U7441 (N_7441,N_4004,N_4646);
nor U7442 (N_7442,N_1943,N_4803);
and U7443 (N_7443,N_2884,N_3871);
or U7444 (N_7444,N_221,N_2845);
nand U7445 (N_7445,N_3207,N_3200);
and U7446 (N_7446,N_3118,N_2812);
and U7447 (N_7447,N_717,N_2987);
nand U7448 (N_7448,N_3541,N_1965);
or U7449 (N_7449,N_3547,N_2116);
nand U7450 (N_7450,N_4874,N_1822);
or U7451 (N_7451,N_1027,N_3435);
or U7452 (N_7452,N_1648,N_1084);
or U7453 (N_7453,N_1634,N_2054);
or U7454 (N_7454,N_1690,N_1222);
nor U7455 (N_7455,N_1947,N_2816);
and U7456 (N_7456,N_4527,N_3163);
or U7457 (N_7457,N_1882,N_4069);
and U7458 (N_7458,N_3925,N_1988);
or U7459 (N_7459,N_2650,N_2171);
xnor U7460 (N_7460,N_4296,N_525);
xnor U7461 (N_7461,N_409,N_3277);
and U7462 (N_7462,N_414,N_1497);
nor U7463 (N_7463,N_2881,N_2450);
or U7464 (N_7464,N_3665,N_731);
and U7465 (N_7465,N_4890,N_3549);
nor U7466 (N_7466,N_4494,N_3376);
and U7467 (N_7467,N_2941,N_3898);
xnor U7468 (N_7468,N_3051,N_1115);
nand U7469 (N_7469,N_4302,N_4984);
nor U7470 (N_7470,N_2474,N_273);
and U7471 (N_7471,N_386,N_3179);
nor U7472 (N_7472,N_990,N_3606);
and U7473 (N_7473,N_2095,N_1774);
or U7474 (N_7474,N_4254,N_1651);
and U7475 (N_7475,N_3255,N_4098);
or U7476 (N_7476,N_800,N_1469);
nor U7477 (N_7477,N_1380,N_4223);
or U7478 (N_7478,N_850,N_323);
and U7479 (N_7479,N_3343,N_130);
nor U7480 (N_7480,N_3607,N_2272);
nand U7481 (N_7481,N_2336,N_3473);
nand U7482 (N_7482,N_1656,N_4362);
or U7483 (N_7483,N_581,N_2169);
and U7484 (N_7484,N_3306,N_4728);
or U7485 (N_7485,N_2002,N_3550);
nor U7486 (N_7486,N_1270,N_4774);
and U7487 (N_7487,N_4118,N_288);
or U7488 (N_7488,N_2442,N_4025);
nand U7489 (N_7489,N_149,N_18);
or U7490 (N_7490,N_1612,N_2643);
and U7491 (N_7491,N_4904,N_1540);
and U7492 (N_7492,N_3950,N_4263);
and U7493 (N_7493,N_3029,N_1501);
xnor U7494 (N_7494,N_4947,N_1240);
nor U7495 (N_7495,N_2094,N_1590);
nand U7496 (N_7496,N_3740,N_1812);
or U7497 (N_7497,N_487,N_1051);
or U7498 (N_7498,N_4723,N_2170);
nor U7499 (N_7499,N_4553,N_3384);
nor U7500 (N_7500,N_4656,N_4311);
and U7501 (N_7501,N_1174,N_1680);
or U7502 (N_7502,N_1978,N_4868);
nor U7503 (N_7503,N_856,N_2506);
nand U7504 (N_7504,N_329,N_2776);
or U7505 (N_7505,N_1507,N_748);
and U7506 (N_7506,N_4854,N_4481);
xnor U7507 (N_7507,N_3539,N_56);
or U7508 (N_7508,N_3815,N_3176);
nand U7509 (N_7509,N_3565,N_211);
and U7510 (N_7510,N_3631,N_4515);
and U7511 (N_7511,N_4452,N_3472);
nor U7512 (N_7512,N_312,N_2160);
xnor U7513 (N_7513,N_4073,N_4617);
nand U7514 (N_7514,N_3051,N_3109);
nand U7515 (N_7515,N_2959,N_1860);
nor U7516 (N_7516,N_1002,N_1221);
nand U7517 (N_7517,N_2053,N_2009);
nand U7518 (N_7518,N_384,N_23);
nand U7519 (N_7519,N_3498,N_2830);
nor U7520 (N_7520,N_4674,N_1952);
nand U7521 (N_7521,N_2078,N_2086);
and U7522 (N_7522,N_1884,N_3239);
or U7523 (N_7523,N_1313,N_1430);
and U7524 (N_7524,N_4076,N_1025);
nor U7525 (N_7525,N_2802,N_4195);
xor U7526 (N_7526,N_445,N_2418);
nor U7527 (N_7527,N_2833,N_1617);
nor U7528 (N_7528,N_2222,N_838);
and U7529 (N_7529,N_2051,N_505);
and U7530 (N_7530,N_149,N_4270);
nor U7531 (N_7531,N_1838,N_544);
nand U7532 (N_7532,N_193,N_1343);
nand U7533 (N_7533,N_147,N_1622);
xnor U7534 (N_7534,N_276,N_1883);
and U7535 (N_7535,N_688,N_4885);
xor U7536 (N_7536,N_1372,N_3230);
and U7537 (N_7537,N_1297,N_1200);
and U7538 (N_7538,N_1773,N_1942);
or U7539 (N_7539,N_254,N_1627);
and U7540 (N_7540,N_2309,N_2612);
nand U7541 (N_7541,N_4759,N_996);
nor U7542 (N_7542,N_3891,N_941);
xor U7543 (N_7543,N_3482,N_3828);
xnor U7544 (N_7544,N_1183,N_2430);
and U7545 (N_7545,N_1725,N_1733);
and U7546 (N_7546,N_2495,N_1275);
xor U7547 (N_7547,N_4876,N_2967);
nand U7548 (N_7548,N_4409,N_3902);
or U7549 (N_7549,N_1986,N_4302);
nor U7550 (N_7550,N_3173,N_1554);
nor U7551 (N_7551,N_166,N_657);
or U7552 (N_7552,N_2257,N_2602);
or U7553 (N_7553,N_3541,N_544);
xor U7554 (N_7554,N_4953,N_4845);
or U7555 (N_7555,N_4440,N_1461);
or U7556 (N_7556,N_2278,N_3555);
and U7557 (N_7557,N_3574,N_1722);
nor U7558 (N_7558,N_2543,N_811);
nor U7559 (N_7559,N_2181,N_475);
nor U7560 (N_7560,N_456,N_3345);
and U7561 (N_7561,N_1184,N_4377);
and U7562 (N_7562,N_1663,N_316);
nand U7563 (N_7563,N_1153,N_3049);
nor U7564 (N_7564,N_1157,N_3214);
and U7565 (N_7565,N_159,N_1644);
and U7566 (N_7566,N_4043,N_133);
or U7567 (N_7567,N_1322,N_388);
or U7568 (N_7568,N_613,N_72);
nor U7569 (N_7569,N_524,N_1621);
xor U7570 (N_7570,N_3485,N_1055);
nand U7571 (N_7571,N_4420,N_1345);
or U7572 (N_7572,N_2569,N_3572);
nor U7573 (N_7573,N_2099,N_1589);
nand U7574 (N_7574,N_4300,N_942);
nor U7575 (N_7575,N_643,N_1615);
xor U7576 (N_7576,N_4428,N_4013);
nand U7577 (N_7577,N_1228,N_4802);
nand U7578 (N_7578,N_579,N_4010);
xor U7579 (N_7579,N_537,N_884);
or U7580 (N_7580,N_4219,N_74);
and U7581 (N_7581,N_2993,N_2842);
or U7582 (N_7582,N_532,N_558);
nand U7583 (N_7583,N_3571,N_811);
xor U7584 (N_7584,N_2670,N_2410);
nand U7585 (N_7585,N_3446,N_2937);
nor U7586 (N_7586,N_484,N_3026);
or U7587 (N_7587,N_4788,N_4572);
nor U7588 (N_7588,N_2959,N_2643);
and U7589 (N_7589,N_370,N_3096);
and U7590 (N_7590,N_1298,N_3388);
nand U7591 (N_7591,N_1768,N_1559);
nor U7592 (N_7592,N_2326,N_135);
or U7593 (N_7593,N_3201,N_4233);
nand U7594 (N_7594,N_2604,N_3418);
or U7595 (N_7595,N_79,N_3575);
or U7596 (N_7596,N_1547,N_2059);
and U7597 (N_7597,N_353,N_4710);
or U7598 (N_7598,N_3817,N_1037);
nor U7599 (N_7599,N_3897,N_3007);
nor U7600 (N_7600,N_1534,N_2565);
nor U7601 (N_7601,N_2227,N_2945);
nand U7602 (N_7602,N_3701,N_3153);
nor U7603 (N_7603,N_2085,N_3481);
nor U7604 (N_7604,N_667,N_4812);
xnor U7605 (N_7605,N_1510,N_295);
nor U7606 (N_7606,N_464,N_4597);
or U7607 (N_7607,N_222,N_1380);
xor U7608 (N_7608,N_2073,N_191);
or U7609 (N_7609,N_2915,N_876);
nor U7610 (N_7610,N_2855,N_3662);
or U7611 (N_7611,N_278,N_2954);
nand U7612 (N_7612,N_3186,N_2844);
xor U7613 (N_7613,N_4075,N_2666);
or U7614 (N_7614,N_591,N_2576);
and U7615 (N_7615,N_3029,N_1296);
nor U7616 (N_7616,N_3362,N_4564);
and U7617 (N_7617,N_4817,N_3304);
nand U7618 (N_7618,N_185,N_4469);
or U7619 (N_7619,N_4999,N_529);
xnor U7620 (N_7620,N_3444,N_3081);
xnor U7621 (N_7621,N_338,N_2807);
xor U7622 (N_7622,N_1083,N_1676);
nand U7623 (N_7623,N_3026,N_4242);
nand U7624 (N_7624,N_3442,N_494);
and U7625 (N_7625,N_1355,N_4046);
xor U7626 (N_7626,N_2519,N_3309);
nand U7627 (N_7627,N_1584,N_3361);
nor U7628 (N_7628,N_4765,N_1597);
or U7629 (N_7629,N_1043,N_2152);
nor U7630 (N_7630,N_3378,N_4224);
and U7631 (N_7631,N_1348,N_3171);
nand U7632 (N_7632,N_4108,N_1665);
nand U7633 (N_7633,N_1028,N_3875);
xor U7634 (N_7634,N_4186,N_2083);
or U7635 (N_7635,N_1467,N_3273);
nand U7636 (N_7636,N_2955,N_343);
nand U7637 (N_7637,N_2974,N_1432);
xnor U7638 (N_7638,N_1016,N_4031);
nor U7639 (N_7639,N_689,N_475);
and U7640 (N_7640,N_3070,N_1846);
and U7641 (N_7641,N_3930,N_2429);
and U7642 (N_7642,N_2693,N_2570);
or U7643 (N_7643,N_2089,N_424);
and U7644 (N_7644,N_729,N_2789);
nor U7645 (N_7645,N_4532,N_4827);
or U7646 (N_7646,N_1716,N_3536);
and U7647 (N_7647,N_881,N_206);
or U7648 (N_7648,N_4688,N_4661);
or U7649 (N_7649,N_4160,N_4980);
or U7650 (N_7650,N_3503,N_1209);
nand U7651 (N_7651,N_181,N_3449);
and U7652 (N_7652,N_1237,N_3689);
nand U7653 (N_7653,N_1081,N_1969);
nand U7654 (N_7654,N_1462,N_233);
and U7655 (N_7655,N_348,N_2508);
or U7656 (N_7656,N_4261,N_2917);
or U7657 (N_7657,N_1381,N_4045);
or U7658 (N_7658,N_3247,N_2038);
and U7659 (N_7659,N_650,N_3852);
or U7660 (N_7660,N_1001,N_552);
and U7661 (N_7661,N_2412,N_4777);
or U7662 (N_7662,N_487,N_1107);
nand U7663 (N_7663,N_837,N_1705);
and U7664 (N_7664,N_2386,N_949);
nand U7665 (N_7665,N_2163,N_2016);
nand U7666 (N_7666,N_787,N_888);
nor U7667 (N_7667,N_2174,N_1853);
nor U7668 (N_7668,N_1396,N_2268);
nand U7669 (N_7669,N_1724,N_3001);
nand U7670 (N_7670,N_2564,N_4450);
nor U7671 (N_7671,N_812,N_4404);
nand U7672 (N_7672,N_4873,N_4510);
or U7673 (N_7673,N_4483,N_3304);
and U7674 (N_7674,N_1360,N_874);
or U7675 (N_7675,N_3045,N_2330);
and U7676 (N_7676,N_2548,N_3016);
or U7677 (N_7677,N_2574,N_170);
nor U7678 (N_7678,N_4695,N_4174);
or U7679 (N_7679,N_3145,N_4181);
nand U7680 (N_7680,N_2589,N_1940);
nor U7681 (N_7681,N_3729,N_715);
nand U7682 (N_7682,N_179,N_363);
nand U7683 (N_7683,N_1955,N_1478);
xor U7684 (N_7684,N_4533,N_4311);
and U7685 (N_7685,N_3752,N_4431);
nand U7686 (N_7686,N_2536,N_770);
and U7687 (N_7687,N_210,N_1388);
or U7688 (N_7688,N_1430,N_2289);
nand U7689 (N_7689,N_204,N_2767);
or U7690 (N_7690,N_2173,N_1650);
nor U7691 (N_7691,N_3541,N_2974);
xor U7692 (N_7692,N_1951,N_2812);
or U7693 (N_7693,N_1900,N_3382);
or U7694 (N_7694,N_1463,N_4963);
nor U7695 (N_7695,N_1582,N_174);
nor U7696 (N_7696,N_2242,N_3902);
or U7697 (N_7697,N_3043,N_3926);
or U7698 (N_7698,N_2736,N_4264);
or U7699 (N_7699,N_2016,N_1607);
nand U7700 (N_7700,N_2131,N_884);
xor U7701 (N_7701,N_430,N_2018);
nor U7702 (N_7702,N_491,N_2198);
and U7703 (N_7703,N_2410,N_3405);
and U7704 (N_7704,N_3221,N_1276);
and U7705 (N_7705,N_3852,N_1421);
and U7706 (N_7706,N_318,N_4924);
and U7707 (N_7707,N_3555,N_3944);
nor U7708 (N_7708,N_1363,N_1016);
and U7709 (N_7709,N_1170,N_4356);
nor U7710 (N_7710,N_4412,N_1531);
xnor U7711 (N_7711,N_553,N_4870);
and U7712 (N_7712,N_3803,N_4456);
and U7713 (N_7713,N_919,N_1431);
nor U7714 (N_7714,N_3451,N_1103);
nand U7715 (N_7715,N_4455,N_836);
or U7716 (N_7716,N_920,N_1354);
nor U7717 (N_7717,N_439,N_1845);
and U7718 (N_7718,N_3806,N_2800);
and U7719 (N_7719,N_4447,N_385);
xor U7720 (N_7720,N_1452,N_4330);
or U7721 (N_7721,N_3634,N_2139);
nor U7722 (N_7722,N_4858,N_4730);
nor U7723 (N_7723,N_4944,N_915);
or U7724 (N_7724,N_4347,N_3755);
and U7725 (N_7725,N_1869,N_4448);
xor U7726 (N_7726,N_4906,N_2045);
xor U7727 (N_7727,N_1605,N_3060);
or U7728 (N_7728,N_4395,N_4415);
or U7729 (N_7729,N_4472,N_2830);
xor U7730 (N_7730,N_3471,N_3293);
nor U7731 (N_7731,N_4538,N_4913);
nand U7732 (N_7732,N_1455,N_3261);
and U7733 (N_7733,N_2381,N_1225);
xor U7734 (N_7734,N_2070,N_1017);
nor U7735 (N_7735,N_3270,N_3935);
nand U7736 (N_7736,N_4325,N_3401);
nor U7737 (N_7737,N_4690,N_3960);
nor U7738 (N_7738,N_2476,N_4274);
or U7739 (N_7739,N_2388,N_1637);
nor U7740 (N_7740,N_459,N_1684);
nor U7741 (N_7741,N_1542,N_3804);
nor U7742 (N_7742,N_1936,N_2010);
and U7743 (N_7743,N_1697,N_2335);
or U7744 (N_7744,N_1494,N_1797);
nand U7745 (N_7745,N_3492,N_4244);
xor U7746 (N_7746,N_1007,N_2387);
and U7747 (N_7747,N_2997,N_478);
nor U7748 (N_7748,N_920,N_3985);
nand U7749 (N_7749,N_1090,N_555);
and U7750 (N_7750,N_3718,N_2943);
and U7751 (N_7751,N_4148,N_3632);
or U7752 (N_7752,N_70,N_4503);
nor U7753 (N_7753,N_641,N_3415);
and U7754 (N_7754,N_1375,N_588);
nor U7755 (N_7755,N_4343,N_2591);
or U7756 (N_7756,N_4555,N_794);
nand U7757 (N_7757,N_2958,N_1912);
nand U7758 (N_7758,N_3808,N_1735);
xnor U7759 (N_7759,N_4790,N_46);
nor U7760 (N_7760,N_4668,N_3048);
xnor U7761 (N_7761,N_3458,N_4040);
or U7762 (N_7762,N_1287,N_3976);
and U7763 (N_7763,N_1530,N_1180);
or U7764 (N_7764,N_3873,N_1050);
nor U7765 (N_7765,N_1086,N_2998);
or U7766 (N_7766,N_2146,N_1654);
nand U7767 (N_7767,N_1368,N_1413);
and U7768 (N_7768,N_3657,N_563);
and U7769 (N_7769,N_123,N_4341);
nand U7770 (N_7770,N_3010,N_4193);
nor U7771 (N_7771,N_226,N_2340);
nand U7772 (N_7772,N_4961,N_4675);
nand U7773 (N_7773,N_1812,N_4468);
xnor U7774 (N_7774,N_3974,N_3434);
nor U7775 (N_7775,N_4929,N_1554);
or U7776 (N_7776,N_2276,N_3596);
and U7777 (N_7777,N_2648,N_3649);
nand U7778 (N_7778,N_3601,N_4433);
and U7779 (N_7779,N_4641,N_4718);
xor U7780 (N_7780,N_24,N_2802);
nor U7781 (N_7781,N_1067,N_1540);
and U7782 (N_7782,N_29,N_346);
and U7783 (N_7783,N_1005,N_3446);
or U7784 (N_7784,N_504,N_3824);
nand U7785 (N_7785,N_2504,N_3519);
and U7786 (N_7786,N_3406,N_2668);
nor U7787 (N_7787,N_11,N_3807);
and U7788 (N_7788,N_2574,N_2629);
nand U7789 (N_7789,N_4486,N_1757);
and U7790 (N_7790,N_4099,N_2192);
or U7791 (N_7791,N_2169,N_1270);
nor U7792 (N_7792,N_1853,N_4042);
and U7793 (N_7793,N_4346,N_409);
xnor U7794 (N_7794,N_1437,N_630);
or U7795 (N_7795,N_9,N_949);
nor U7796 (N_7796,N_4787,N_792);
nand U7797 (N_7797,N_608,N_3642);
or U7798 (N_7798,N_1972,N_444);
and U7799 (N_7799,N_561,N_3639);
and U7800 (N_7800,N_287,N_1117);
nand U7801 (N_7801,N_1363,N_2365);
and U7802 (N_7802,N_3396,N_1946);
nor U7803 (N_7803,N_3252,N_3247);
nand U7804 (N_7804,N_2556,N_598);
or U7805 (N_7805,N_2817,N_501);
and U7806 (N_7806,N_2537,N_1981);
xor U7807 (N_7807,N_4103,N_4917);
nor U7808 (N_7808,N_2837,N_4822);
or U7809 (N_7809,N_564,N_3219);
xnor U7810 (N_7810,N_2660,N_4063);
or U7811 (N_7811,N_893,N_385);
nor U7812 (N_7812,N_4955,N_2677);
nor U7813 (N_7813,N_2698,N_12);
nand U7814 (N_7814,N_2835,N_4510);
nor U7815 (N_7815,N_1458,N_3347);
nand U7816 (N_7816,N_3515,N_2963);
nand U7817 (N_7817,N_782,N_2239);
or U7818 (N_7818,N_1596,N_775);
xnor U7819 (N_7819,N_3399,N_4223);
or U7820 (N_7820,N_2178,N_2458);
nor U7821 (N_7821,N_2598,N_1902);
nor U7822 (N_7822,N_3704,N_667);
xor U7823 (N_7823,N_3930,N_1304);
or U7824 (N_7824,N_2763,N_4094);
nand U7825 (N_7825,N_418,N_4568);
or U7826 (N_7826,N_767,N_3432);
nand U7827 (N_7827,N_1649,N_843);
nand U7828 (N_7828,N_921,N_1776);
nor U7829 (N_7829,N_4258,N_1240);
or U7830 (N_7830,N_2821,N_4709);
nor U7831 (N_7831,N_317,N_2514);
nor U7832 (N_7832,N_1928,N_4819);
nand U7833 (N_7833,N_30,N_1924);
nor U7834 (N_7834,N_3470,N_1287);
nor U7835 (N_7835,N_4831,N_1696);
nor U7836 (N_7836,N_1099,N_2838);
nor U7837 (N_7837,N_2011,N_4291);
xor U7838 (N_7838,N_1213,N_4273);
and U7839 (N_7839,N_381,N_4388);
nor U7840 (N_7840,N_2991,N_2559);
or U7841 (N_7841,N_874,N_2531);
nor U7842 (N_7842,N_1326,N_906);
nor U7843 (N_7843,N_266,N_2673);
nand U7844 (N_7844,N_547,N_3383);
and U7845 (N_7845,N_1482,N_977);
or U7846 (N_7846,N_2404,N_1812);
or U7847 (N_7847,N_2284,N_2829);
nand U7848 (N_7848,N_3046,N_1385);
and U7849 (N_7849,N_2955,N_582);
and U7850 (N_7850,N_2903,N_2264);
or U7851 (N_7851,N_4196,N_2901);
and U7852 (N_7852,N_747,N_3247);
and U7853 (N_7853,N_2062,N_0);
nor U7854 (N_7854,N_3346,N_1640);
nand U7855 (N_7855,N_4895,N_2161);
or U7856 (N_7856,N_3682,N_4276);
nor U7857 (N_7857,N_3224,N_4907);
and U7858 (N_7858,N_4939,N_3589);
xor U7859 (N_7859,N_2681,N_3732);
xnor U7860 (N_7860,N_4777,N_3243);
and U7861 (N_7861,N_357,N_4662);
nor U7862 (N_7862,N_1152,N_42);
xor U7863 (N_7863,N_1788,N_3975);
or U7864 (N_7864,N_1925,N_4806);
nor U7865 (N_7865,N_1417,N_4050);
nand U7866 (N_7866,N_4658,N_3440);
and U7867 (N_7867,N_4289,N_2778);
and U7868 (N_7868,N_883,N_1451);
and U7869 (N_7869,N_1998,N_97);
nand U7870 (N_7870,N_720,N_2716);
nor U7871 (N_7871,N_345,N_698);
or U7872 (N_7872,N_4802,N_3596);
or U7873 (N_7873,N_46,N_2151);
or U7874 (N_7874,N_1170,N_2074);
or U7875 (N_7875,N_3469,N_3524);
or U7876 (N_7876,N_3891,N_959);
or U7877 (N_7877,N_2195,N_1339);
nor U7878 (N_7878,N_1940,N_3358);
xor U7879 (N_7879,N_1649,N_188);
xnor U7880 (N_7880,N_3321,N_714);
nand U7881 (N_7881,N_656,N_1599);
nor U7882 (N_7882,N_4572,N_1581);
nor U7883 (N_7883,N_242,N_2777);
nand U7884 (N_7884,N_1282,N_1746);
xor U7885 (N_7885,N_414,N_1118);
and U7886 (N_7886,N_2551,N_2445);
and U7887 (N_7887,N_4480,N_616);
nand U7888 (N_7888,N_1348,N_2361);
nand U7889 (N_7889,N_2686,N_4544);
nor U7890 (N_7890,N_3947,N_4415);
and U7891 (N_7891,N_435,N_4471);
nand U7892 (N_7892,N_3767,N_4600);
nor U7893 (N_7893,N_1000,N_2138);
and U7894 (N_7894,N_4827,N_4416);
nand U7895 (N_7895,N_1500,N_1672);
nor U7896 (N_7896,N_334,N_3545);
nor U7897 (N_7897,N_561,N_3918);
nand U7898 (N_7898,N_4759,N_4133);
nand U7899 (N_7899,N_4924,N_2674);
and U7900 (N_7900,N_360,N_285);
nor U7901 (N_7901,N_1019,N_4542);
nand U7902 (N_7902,N_565,N_3810);
and U7903 (N_7903,N_1907,N_1861);
or U7904 (N_7904,N_1898,N_193);
and U7905 (N_7905,N_3104,N_4113);
and U7906 (N_7906,N_1608,N_3371);
or U7907 (N_7907,N_4559,N_4928);
or U7908 (N_7908,N_1022,N_2749);
nand U7909 (N_7909,N_958,N_4574);
and U7910 (N_7910,N_3985,N_4503);
nor U7911 (N_7911,N_3887,N_2854);
nor U7912 (N_7912,N_2923,N_4182);
xor U7913 (N_7913,N_3159,N_3785);
nor U7914 (N_7914,N_1014,N_4854);
nand U7915 (N_7915,N_3633,N_1218);
nor U7916 (N_7916,N_4986,N_3760);
or U7917 (N_7917,N_3882,N_2906);
xnor U7918 (N_7918,N_3498,N_203);
and U7919 (N_7919,N_803,N_881);
and U7920 (N_7920,N_4723,N_653);
nor U7921 (N_7921,N_4261,N_1742);
and U7922 (N_7922,N_3323,N_3470);
xnor U7923 (N_7923,N_215,N_741);
nor U7924 (N_7924,N_2143,N_4789);
and U7925 (N_7925,N_2473,N_1929);
or U7926 (N_7926,N_3339,N_2470);
nand U7927 (N_7927,N_4874,N_2495);
or U7928 (N_7928,N_2595,N_1418);
and U7929 (N_7929,N_2598,N_233);
or U7930 (N_7930,N_2520,N_4695);
nor U7931 (N_7931,N_3061,N_1275);
or U7932 (N_7932,N_3129,N_4479);
nand U7933 (N_7933,N_4815,N_2981);
nand U7934 (N_7934,N_1838,N_3255);
nand U7935 (N_7935,N_2208,N_2477);
or U7936 (N_7936,N_1024,N_2770);
nor U7937 (N_7937,N_194,N_4535);
or U7938 (N_7938,N_4381,N_413);
nand U7939 (N_7939,N_287,N_2749);
and U7940 (N_7940,N_1494,N_531);
nor U7941 (N_7941,N_314,N_3261);
nand U7942 (N_7942,N_1360,N_131);
or U7943 (N_7943,N_2649,N_1511);
and U7944 (N_7944,N_2087,N_228);
nor U7945 (N_7945,N_1316,N_1734);
or U7946 (N_7946,N_2430,N_4379);
and U7947 (N_7947,N_3817,N_4622);
and U7948 (N_7948,N_3949,N_4103);
and U7949 (N_7949,N_1573,N_2626);
and U7950 (N_7950,N_2850,N_2581);
nand U7951 (N_7951,N_2719,N_4107);
xnor U7952 (N_7952,N_2825,N_1843);
xor U7953 (N_7953,N_3592,N_4603);
nor U7954 (N_7954,N_3746,N_2927);
or U7955 (N_7955,N_2498,N_1536);
or U7956 (N_7956,N_2452,N_1033);
or U7957 (N_7957,N_224,N_3532);
or U7958 (N_7958,N_2115,N_2631);
nor U7959 (N_7959,N_3615,N_140);
and U7960 (N_7960,N_2869,N_4539);
nor U7961 (N_7961,N_2508,N_3449);
and U7962 (N_7962,N_876,N_3475);
xor U7963 (N_7963,N_956,N_4713);
or U7964 (N_7964,N_3182,N_533);
nand U7965 (N_7965,N_1656,N_2825);
nor U7966 (N_7966,N_330,N_1975);
and U7967 (N_7967,N_1202,N_158);
nand U7968 (N_7968,N_4130,N_3134);
nor U7969 (N_7969,N_1576,N_2622);
nor U7970 (N_7970,N_3500,N_1822);
or U7971 (N_7971,N_4232,N_4502);
nor U7972 (N_7972,N_4431,N_1057);
and U7973 (N_7973,N_3214,N_1780);
nand U7974 (N_7974,N_1756,N_4110);
nand U7975 (N_7975,N_4057,N_1320);
and U7976 (N_7976,N_4447,N_4842);
nor U7977 (N_7977,N_1114,N_560);
nand U7978 (N_7978,N_2595,N_709);
nand U7979 (N_7979,N_2428,N_1887);
nor U7980 (N_7980,N_4007,N_415);
and U7981 (N_7981,N_762,N_1568);
or U7982 (N_7982,N_4752,N_3396);
nand U7983 (N_7983,N_2631,N_1211);
xor U7984 (N_7984,N_540,N_1390);
nand U7985 (N_7985,N_4941,N_1018);
nand U7986 (N_7986,N_2784,N_2644);
or U7987 (N_7987,N_3565,N_4462);
or U7988 (N_7988,N_815,N_73);
nand U7989 (N_7989,N_3195,N_4008);
nand U7990 (N_7990,N_105,N_2516);
nand U7991 (N_7991,N_2800,N_2658);
nor U7992 (N_7992,N_1295,N_4197);
and U7993 (N_7993,N_3838,N_834);
xor U7994 (N_7994,N_3633,N_3563);
nor U7995 (N_7995,N_2534,N_481);
and U7996 (N_7996,N_1320,N_3636);
or U7997 (N_7997,N_2752,N_3936);
nand U7998 (N_7998,N_1941,N_968);
nor U7999 (N_7999,N_822,N_170);
nand U8000 (N_8000,N_4617,N_406);
nand U8001 (N_8001,N_4344,N_2358);
or U8002 (N_8002,N_1526,N_4315);
nand U8003 (N_8003,N_4085,N_2591);
nand U8004 (N_8004,N_465,N_428);
nor U8005 (N_8005,N_2024,N_4201);
and U8006 (N_8006,N_1716,N_4924);
xnor U8007 (N_8007,N_4285,N_3863);
nand U8008 (N_8008,N_2371,N_4608);
nor U8009 (N_8009,N_3576,N_2704);
and U8010 (N_8010,N_4298,N_27);
and U8011 (N_8011,N_3944,N_2895);
nor U8012 (N_8012,N_4198,N_2942);
nor U8013 (N_8013,N_2470,N_2279);
nor U8014 (N_8014,N_2157,N_389);
or U8015 (N_8015,N_2461,N_216);
nor U8016 (N_8016,N_2695,N_1002);
nand U8017 (N_8017,N_4198,N_4784);
or U8018 (N_8018,N_4374,N_1136);
xor U8019 (N_8019,N_4243,N_3548);
and U8020 (N_8020,N_1972,N_3096);
and U8021 (N_8021,N_3016,N_500);
or U8022 (N_8022,N_2173,N_4608);
and U8023 (N_8023,N_4119,N_441);
nand U8024 (N_8024,N_1871,N_582);
and U8025 (N_8025,N_4684,N_3644);
and U8026 (N_8026,N_1333,N_3621);
nand U8027 (N_8027,N_3912,N_2513);
and U8028 (N_8028,N_3212,N_2846);
xor U8029 (N_8029,N_3499,N_2914);
nor U8030 (N_8030,N_2404,N_639);
nand U8031 (N_8031,N_4925,N_2411);
nor U8032 (N_8032,N_3788,N_15);
nor U8033 (N_8033,N_340,N_837);
nand U8034 (N_8034,N_3137,N_2349);
nor U8035 (N_8035,N_4144,N_3691);
nor U8036 (N_8036,N_4499,N_290);
and U8037 (N_8037,N_4439,N_596);
nand U8038 (N_8038,N_1296,N_1196);
nand U8039 (N_8039,N_2406,N_1165);
and U8040 (N_8040,N_1842,N_3487);
nand U8041 (N_8041,N_489,N_1804);
and U8042 (N_8042,N_9,N_1623);
nand U8043 (N_8043,N_1196,N_2484);
or U8044 (N_8044,N_1878,N_4733);
nor U8045 (N_8045,N_2756,N_4514);
nand U8046 (N_8046,N_4148,N_4309);
or U8047 (N_8047,N_3685,N_3623);
and U8048 (N_8048,N_1824,N_2049);
nand U8049 (N_8049,N_1249,N_4078);
or U8050 (N_8050,N_3165,N_4677);
nor U8051 (N_8051,N_1430,N_3808);
nor U8052 (N_8052,N_1124,N_899);
and U8053 (N_8053,N_4089,N_181);
nor U8054 (N_8054,N_2400,N_3158);
nor U8055 (N_8055,N_3113,N_83);
and U8056 (N_8056,N_2100,N_2488);
or U8057 (N_8057,N_1308,N_4389);
and U8058 (N_8058,N_2148,N_2500);
nor U8059 (N_8059,N_2116,N_209);
nor U8060 (N_8060,N_2642,N_1148);
nor U8061 (N_8061,N_1982,N_41);
nor U8062 (N_8062,N_3778,N_2981);
nand U8063 (N_8063,N_1023,N_247);
or U8064 (N_8064,N_3456,N_4073);
or U8065 (N_8065,N_2209,N_652);
or U8066 (N_8066,N_1250,N_3385);
nand U8067 (N_8067,N_2166,N_2250);
nor U8068 (N_8068,N_3797,N_3034);
nand U8069 (N_8069,N_3089,N_980);
or U8070 (N_8070,N_2785,N_2575);
nand U8071 (N_8071,N_3366,N_2831);
nor U8072 (N_8072,N_2186,N_548);
xnor U8073 (N_8073,N_782,N_4576);
nor U8074 (N_8074,N_2643,N_3143);
and U8075 (N_8075,N_3255,N_3037);
nand U8076 (N_8076,N_3513,N_3188);
nor U8077 (N_8077,N_3733,N_4397);
xor U8078 (N_8078,N_2145,N_651);
or U8079 (N_8079,N_3884,N_3623);
or U8080 (N_8080,N_4080,N_987);
or U8081 (N_8081,N_2342,N_1054);
xnor U8082 (N_8082,N_547,N_1160);
and U8083 (N_8083,N_300,N_1616);
xor U8084 (N_8084,N_3113,N_3714);
nor U8085 (N_8085,N_4575,N_2769);
or U8086 (N_8086,N_4196,N_1870);
nor U8087 (N_8087,N_2039,N_4250);
nand U8088 (N_8088,N_1340,N_2635);
nor U8089 (N_8089,N_3834,N_4538);
nand U8090 (N_8090,N_220,N_1418);
and U8091 (N_8091,N_2132,N_2679);
nand U8092 (N_8092,N_3814,N_1620);
nand U8093 (N_8093,N_4128,N_368);
and U8094 (N_8094,N_2297,N_2281);
and U8095 (N_8095,N_2826,N_3721);
nor U8096 (N_8096,N_11,N_441);
nand U8097 (N_8097,N_4574,N_1619);
and U8098 (N_8098,N_1827,N_2483);
and U8099 (N_8099,N_1210,N_2979);
or U8100 (N_8100,N_3317,N_1013);
and U8101 (N_8101,N_4501,N_393);
nor U8102 (N_8102,N_4976,N_4245);
or U8103 (N_8103,N_4567,N_68);
and U8104 (N_8104,N_4028,N_2199);
and U8105 (N_8105,N_2714,N_3328);
or U8106 (N_8106,N_646,N_2222);
nand U8107 (N_8107,N_2271,N_779);
nor U8108 (N_8108,N_2997,N_1372);
nand U8109 (N_8109,N_3022,N_1471);
or U8110 (N_8110,N_3421,N_953);
nor U8111 (N_8111,N_2512,N_2183);
and U8112 (N_8112,N_718,N_3182);
nand U8113 (N_8113,N_2819,N_2364);
and U8114 (N_8114,N_1254,N_1939);
xnor U8115 (N_8115,N_3016,N_933);
nor U8116 (N_8116,N_1626,N_883);
nand U8117 (N_8117,N_348,N_3291);
nor U8118 (N_8118,N_2257,N_3932);
nand U8119 (N_8119,N_4289,N_2345);
and U8120 (N_8120,N_1389,N_968);
nor U8121 (N_8121,N_1008,N_4382);
nand U8122 (N_8122,N_248,N_4116);
or U8123 (N_8123,N_3792,N_2673);
nand U8124 (N_8124,N_2957,N_1350);
xor U8125 (N_8125,N_1280,N_2906);
or U8126 (N_8126,N_11,N_782);
or U8127 (N_8127,N_2226,N_3866);
nor U8128 (N_8128,N_4032,N_2065);
nand U8129 (N_8129,N_2721,N_2293);
nand U8130 (N_8130,N_859,N_3499);
nand U8131 (N_8131,N_4486,N_3520);
nand U8132 (N_8132,N_3663,N_4455);
nand U8133 (N_8133,N_1670,N_1072);
and U8134 (N_8134,N_4657,N_1992);
and U8135 (N_8135,N_3174,N_884);
nor U8136 (N_8136,N_119,N_4920);
xor U8137 (N_8137,N_4104,N_2245);
or U8138 (N_8138,N_1028,N_2982);
nand U8139 (N_8139,N_906,N_3650);
and U8140 (N_8140,N_4659,N_3250);
and U8141 (N_8141,N_89,N_3096);
xor U8142 (N_8142,N_2104,N_4960);
nor U8143 (N_8143,N_968,N_4944);
or U8144 (N_8144,N_2964,N_1136);
and U8145 (N_8145,N_2941,N_1456);
nor U8146 (N_8146,N_2224,N_4600);
and U8147 (N_8147,N_3780,N_2240);
xnor U8148 (N_8148,N_4353,N_4955);
or U8149 (N_8149,N_4437,N_1596);
nor U8150 (N_8150,N_562,N_3486);
or U8151 (N_8151,N_3912,N_2719);
or U8152 (N_8152,N_4969,N_4781);
xor U8153 (N_8153,N_3747,N_4894);
and U8154 (N_8154,N_4431,N_4215);
nor U8155 (N_8155,N_1163,N_2985);
nor U8156 (N_8156,N_125,N_3050);
and U8157 (N_8157,N_4398,N_3533);
nand U8158 (N_8158,N_3134,N_2283);
and U8159 (N_8159,N_3873,N_654);
or U8160 (N_8160,N_1047,N_3992);
or U8161 (N_8161,N_486,N_1925);
or U8162 (N_8162,N_3915,N_3838);
and U8163 (N_8163,N_3389,N_4636);
xor U8164 (N_8164,N_263,N_1482);
or U8165 (N_8165,N_4578,N_1956);
and U8166 (N_8166,N_3048,N_1186);
or U8167 (N_8167,N_415,N_4935);
and U8168 (N_8168,N_4509,N_2205);
xor U8169 (N_8169,N_2319,N_1076);
nor U8170 (N_8170,N_1643,N_3647);
or U8171 (N_8171,N_1367,N_111);
nand U8172 (N_8172,N_223,N_1560);
or U8173 (N_8173,N_4738,N_2590);
nor U8174 (N_8174,N_1984,N_217);
nand U8175 (N_8175,N_16,N_211);
nand U8176 (N_8176,N_2668,N_3220);
or U8177 (N_8177,N_4619,N_2120);
nand U8178 (N_8178,N_2782,N_3838);
or U8179 (N_8179,N_4674,N_3388);
and U8180 (N_8180,N_1072,N_2537);
xor U8181 (N_8181,N_4388,N_691);
nand U8182 (N_8182,N_3269,N_4773);
nand U8183 (N_8183,N_1481,N_345);
nor U8184 (N_8184,N_4909,N_4797);
or U8185 (N_8185,N_3710,N_3691);
nand U8186 (N_8186,N_3045,N_3504);
nand U8187 (N_8187,N_4193,N_3941);
nor U8188 (N_8188,N_3615,N_633);
or U8189 (N_8189,N_1856,N_1553);
and U8190 (N_8190,N_33,N_1584);
or U8191 (N_8191,N_3382,N_4730);
and U8192 (N_8192,N_2266,N_3667);
or U8193 (N_8193,N_2836,N_990);
nor U8194 (N_8194,N_4077,N_110);
xor U8195 (N_8195,N_3800,N_4137);
or U8196 (N_8196,N_500,N_985);
or U8197 (N_8197,N_4797,N_4934);
nand U8198 (N_8198,N_3001,N_2510);
or U8199 (N_8199,N_4773,N_1053);
xor U8200 (N_8200,N_3635,N_3965);
or U8201 (N_8201,N_3402,N_2554);
and U8202 (N_8202,N_2931,N_1291);
or U8203 (N_8203,N_3776,N_2819);
xnor U8204 (N_8204,N_1862,N_2460);
nor U8205 (N_8205,N_823,N_225);
nand U8206 (N_8206,N_49,N_989);
or U8207 (N_8207,N_462,N_3371);
nand U8208 (N_8208,N_524,N_680);
nor U8209 (N_8209,N_1258,N_1097);
or U8210 (N_8210,N_2909,N_615);
nand U8211 (N_8211,N_4502,N_310);
nand U8212 (N_8212,N_2476,N_3754);
and U8213 (N_8213,N_1,N_2032);
nor U8214 (N_8214,N_2713,N_4077);
and U8215 (N_8215,N_1035,N_3346);
nor U8216 (N_8216,N_1626,N_664);
and U8217 (N_8217,N_790,N_281);
nand U8218 (N_8218,N_2345,N_1307);
and U8219 (N_8219,N_3718,N_4062);
nand U8220 (N_8220,N_2925,N_2870);
nor U8221 (N_8221,N_387,N_3848);
nand U8222 (N_8222,N_1957,N_1602);
or U8223 (N_8223,N_1602,N_1433);
nor U8224 (N_8224,N_158,N_922);
nand U8225 (N_8225,N_1365,N_3924);
nand U8226 (N_8226,N_2082,N_4687);
or U8227 (N_8227,N_2464,N_2299);
xnor U8228 (N_8228,N_1202,N_2847);
and U8229 (N_8229,N_1649,N_704);
nand U8230 (N_8230,N_1541,N_3278);
and U8231 (N_8231,N_4247,N_2353);
nor U8232 (N_8232,N_2104,N_3534);
xnor U8233 (N_8233,N_1852,N_1883);
xor U8234 (N_8234,N_4539,N_111);
and U8235 (N_8235,N_4940,N_4590);
and U8236 (N_8236,N_4899,N_4801);
nand U8237 (N_8237,N_3552,N_2819);
or U8238 (N_8238,N_2023,N_1727);
and U8239 (N_8239,N_1048,N_4093);
or U8240 (N_8240,N_422,N_105);
and U8241 (N_8241,N_1344,N_2705);
nand U8242 (N_8242,N_2717,N_2864);
nand U8243 (N_8243,N_1654,N_4662);
and U8244 (N_8244,N_2192,N_2897);
or U8245 (N_8245,N_2826,N_3208);
nor U8246 (N_8246,N_4463,N_3662);
or U8247 (N_8247,N_4298,N_161);
and U8248 (N_8248,N_1636,N_2072);
and U8249 (N_8249,N_1801,N_1060);
nor U8250 (N_8250,N_4002,N_1767);
nor U8251 (N_8251,N_424,N_1002);
nor U8252 (N_8252,N_2864,N_4139);
nand U8253 (N_8253,N_255,N_90);
or U8254 (N_8254,N_4001,N_4646);
nand U8255 (N_8255,N_3463,N_1009);
or U8256 (N_8256,N_2681,N_2397);
nor U8257 (N_8257,N_455,N_530);
xnor U8258 (N_8258,N_4316,N_123);
nor U8259 (N_8259,N_1938,N_4245);
or U8260 (N_8260,N_832,N_1319);
and U8261 (N_8261,N_3057,N_3008);
or U8262 (N_8262,N_3453,N_2095);
or U8263 (N_8263,N_4576,N_2717);
xnor U8264 (N_8264,N_4592,N_540);
and U8265 (N_8265,N_4404,N_960);
nor U8266 (N_8266,N_168,N_3320);
or U8267 (N_8267,N_1774,N_2808);
nand U8268 (N_8268,N_115,N_1940);
and U8269 (N_8269,N_1065,N_4924);
nand U8270 (N_8270,N_2298,N_4288);
or U8271 (N_8271,N_4070,N_820);
nor U8272 (N_8272,N_2351,N_2140);
nand U8273 (N_8273,N_2340,N_4791);
nor U8274 (N_8274,N_2482,N_290);
and U8275 (N_8275,N_4344,N_2755);
and U8276 (N_8276,N_4281,N_3110);
and U8277 (N_8277,N_2194,N_4155);
or U8278 (N_8278,N_3846,N_1098);
nand U8279 (N_8279,N_2703,N_1877);
nor U8280 (N_8280,N_2121,N_3737);
and U8281 (N_8281,N_524,N_1062);
and U8282 (N_8282,N_3956,N_3536);
or U8283 (N_8283,N_849,N_1635);
nand U8284 (N_8284,N_2734,N_1923);
nand U8285 (N_8285,N_692,N_3311);
and U8286 (N_8286,N_4597,N_140);
and U8287 (N_8287,N_633,N_2281);
nor U8288 (N_8288,N_2941,N_3425);
nand U8289 (N_8289,N_415,N_398);
xnor U8290 (N_8290,N_3180,N_721);
xnor U8291 (N_8291,N_4585,N_850);
or U8292 (N_8292,N_4371,N_2170);
or U8293 (N_8293,N_3126,N_4930);
nor U8294 (N_8294,N_140,N_3766);
or U8295 (N_8295,N_1273,N_4987);
and U8296 (N_8296,N_35,N_1473);
and U8297 (N_8297,N_1616,N_2736);
or U8298 (N_8298,N_2798,N_3890);
xor U8299 (N_8299,N_3100,N_1791);
or U8300 (N_8300,N_524,N_3796);
or U8301 (N_8301,N_916,N_4931);
xnor U8302 (N_8302,N_4193,N_2132);
nand U8303 (N_8303,N_576,N_2575);
and U8304 (N_8304,N_3822,N_3194);
or U8305 (N_8305,N_2731,N_201);
nor U8306 (N_8306,N_1665,N_3807);
xor U8307 (N_8307,N_3679,N_1141);
xor U8308 (N_8308,N_4159,N_1240);
nor U8309 (N_8309,N_94,N_2966);
or U8310 (N_8310,N_2268,N_1885);
or U8311 (N_8311,N_2846,N_3935);
and U8312 (N_8312,N_2237,N_2602);
nor U8313 (N_8313,N_1898,N_3786);
nor U8314 (N_8314,N_4694,N_2571);
nand U8315 (N_8315,N_2598,N_3178);
nor U8316 (N_8316,N_4738,N_1217);
and U8317 (N_8317,N_2099,N_2678);
nand U8318 (N_8318,N_4117,N_537);
nor U8319 (N_8319,N_4003,N_953);
nor U8320 (N_8320,N_4594,N_638);
or U8321 (N_8321,N_1552,N_3321);
nor U8322 (N_8322,N_4386,N_284);
nand U8323 (N_8323,N_776,N_4110);
and U8324 (N_8324,N_1008,N_3400);
nor U8325 (N_8325,N_597,N_1072);
nor U8326 (N_8326,N_4236,N_3235);
or U8327 (N_8327,N_752,N_2533);
or U8328 (N_8328,N_3776,N_4817);
nand U8329 (N_8329,N_2528,N_888);
nand U8330 (N_8330,N_2245,N_1299);
xor U8331 (N_8331,N_3227,N_4781);
nand U8332 (N_8332,N_4948,N_4672);
nand U8333 (N_8333,N_2207,N_3194);
or U8334 (N_8334,N_762,N_4361);
or U8335 (N_8335,N_47,N_2446);
or U8336 (N_8336,N_85,N_1278);
xor U8337 (N_8337,N_4579,N_4541);
xor U8338 (N_8338,N_252,N_3973);
nor U8339 (N_8339,N_1977,N_3042);
nand U8340 (N_8340,N_1102,N_4482);
nand U8341 (N_8341,N_2739,N_4682);
xor U8342 (N_8342,N_4348,N_3193);
and U8343 (N_8343,N_3467,N_3775);
and U8344 (N_8344,N_398,N_3705);
and U8345 (N_8345,N_2294,N_819);
nand U8346 (N_8346,N_4449,N_2985);
xnor U8347 (N_8347,N_2165,N_4523);
xnor U8348 (N_8348,N_2029,N_1248);
and U8349 (N_8349,N_3303,N_4072);
nor U8350 (N_8350,N_3331,N_2388);
nor U8351 (N_8351,N_369,N_2452);
and U8352 (N_8352,N_2423,N_2473);
nand U8353 (N_8353,N_3613,N_1503);
and U8354 (N_8354,N_2654,N_4295);
nor U8355 (N_8355,N_235,N_2044);
nor U8356 (N_8356,N_21,N_2347);
or U8357 (N_8357,N_2965,N_235);
nor U8358 (N_8358,N_2733,N_4229);
nor U8359 (N_8359,N_291,N_4926);
nand U8360 (N_8360,N_4131,N_73);
nand U8361 (N_8361,N_1499,N_4833);
and U8362 (N_8362,N_3391,N_4402);
nand U8363 (N_8363,N_4984,N_1418);
nand U8364 (N_8364,N_1177,N_3889);
xor U8365 (N_8365,N_3567,N_3672);
and U8366 (N_8366,N_3272,N_2128);
or U8367 (N_8367,N_2841,N_1469);
or U8368 (N_8368,N_287,N_2624);
nor U8369 (N_8369,N_3796,N_4236);
or U8370 (N_8370,N_786,N_747);
nand U8371 (N_8371,N_1211,N_2870);
nand U8372 (N_8372,N_4207,N_1907);
nor U8373 (N_8373,N_858,N_1910);
and U8374 (N_8374,N_1287,N_619);
and U8375 (N_8375,N_2417,N_951);
and U8376 (N_8376,N_3686,N_4386);
nand U8377 (N_8377,N_2915,N_1924);
nand U8378 (N_8378,N_394,N_4007);
nand U8379 (N_8379,N_3214,N_3844);
or U8380 (N_8380,N_4214,N_228);
and U8381 (N_8381,N_3351,N_2629);
nor U8382 (N_8382,N_26,N_4922);
nand U8383 (N_8383,N_72,N_1900);
or U8384 (N_8384,N_1619,N_3977);
nor U8385 (N_8385,N_1697,N_252);
nor U8386 (N_8386,N_1551,N_4044);
nor U8387 (N_8387,N_3341,N_3913);
and U8388 (N_8388,N_4796,N_3890);
nor U8389 (N_8389,N_1196,N_491);
nor U8390 (N_8390,N_703,N_2028);
and U8391 (N_8391,N_2624,N_4256);
and U8392 (N_8392,N_1130,N_1940);
nand U8393 (N_8393,N_4048,N_547);
nor U8394 (N_8394,N_269,N_2562);
nor U8395 (N_8395,N_3,N_4572);
xor U8396 (N_8396,N_1562,N_2390);
nor U8397 (N_8397,N_3146,N_652);
nor U8398 (N_8398,N_2255,N_2632);
nor U8399 (N_8399,N_392,N_2276);
xnor U8400 (N_8400,N_4866,N_2541);
and U8401 (N_8401,N_2113,N_3712);
nand U8402 (N_8402,N_1249,N_4505);
nand U8403 (N_8403,N_1050,N_2594);
and U8404 (N_8404,N_1304,N_4936);
xor U8405 (N_8405,N_4335,N_109);
or U8406 (N_8406,N_595,N_3578);
xor U8407 (N_8407,N_4065,N_1433);
or U8408 (N_8408,N_3548,N_1742);
and U8409 (N_8409,N_1439,N_2689);
nor U8410 (N_8410,N_4249,N_1671);
nor U8411 (N_8411,N_2883,N_4664);
nand U8412 (N_8412,N_2957,N_925);
or U8413 (N_8413,N_2701,N_2250);
nand U8414 (N_8414,N_1009,N_2421);
nand U8415 (N_8415,N_969,N_1441);
nor U8416 (N_8416,N_180,N_3720);
xor U8417 (N_8417,N_2251,N_1510);
or U8418 (N_8418,N_4809,N_2331);
and U8419 (N_8419,N_3636,N_369);
or U8420 (N_8420,N_2468,N_4791);
and U8421 (N_8421,N_3899,N_3248);
nand U8422 (N_8422,N_4410,N_4034);
or U8423 (N_8423,N_4742,N_4026);
or U8424 (N_8424,N_274,N_2607);
nand U8425 (N_8425,N_3972,N_2619);
nand U8426 (N_8426,N_3609,N_1221);
nand U8427 (N_8427,N_3790,N_3950);
and U8428 (N_8428,N_564,N_4972);
nand U8429 (N_8429,N_3622,N_2711);
nand U8430 (N_8430,N_3826,N_3449);
and U8431 (N_8431,N_660,N_656);
and U8432 (N_8432,N_1057,N_4256);
and U8433 (N_8433,N_1892,N_3570);
or U8434 (N_8434,N_2496,N_831);
or U8435 (N_8435,N_3000,N_786);
nand U8436 (N_8436,N_1,N_3636);
nand U8437 (N_8437,N_1632,N_2134);
and U8438 (N_8438,N_945,N_1078);
nand U8439 (N_8439,N_4467,N_3623);
nand U8440 (N_8440,N_3111,N_2212);
and U8441 (N_8441,N_3015,N_582);
nand U8442 (N_8442,N_1788,N_4514);
or U8443 (N_8443,N_3836,N_3152);
nand U8444 (N_8444,N_4076,N_4220);
and U8445 (N_8445,N_2104,N_3425);
nand U8446 (N_8446,N_2865,N_3316);
or U8447 (N_8447,N_3942,N_2677);
or U8448 (N_8448,N_4877,N_4225);
nand U8449 (N_8449,N_1079,N_2380);
and U8450 (N_8450,N_1251,N_1198);
nand U8451 (N_8451,N_1918,N_4681);
nor U8452 (N_8452,N_3931,N_247);
nor U8453 (N_8453,N_1374,N_770);
and U8454 (N_8454,N_4386,N_348);
nand U8455 (N_8455,N_340,N_3594);
nand U8456 (N_8456,N_2274,N_1697);
or U8457 (N_8457,N_2848,N_2977);
xor U8458 (N_8458,N_4472,N_2092);
nand U8459 (N_8459,N_1256,N_3068);
and U8460 (N_8460,N_692,N_288);
nand U8461 (N_8461,N_2203,N_3615);
xnor U8462 (N_8462,N_887,N_4267);
nor U8463 (N_8463,N_783,N_491);
or U8464 (N_8464,N_1321,N_663);
nand U8465 (N_8465,N_3989,N_1434);
nor U8466 (N_8466,N_2954,N_2992);
nand U8467 (N_8467,N_2578,N_2988);
or U8468 (N_8468,N_4194,N_1422);
nor U8469 (N_8469,N_4998,N_2062);
xnor U8470 (N_8470,N_1897,N_3399);
or U8471 (N_8471,N_3567,N_1711);
nor U8472 (N_8472,N_1713,N_1945);
nand U8473 (N_8473,N_4226,N_1822);
nand U8474 (N_8474,N_1909,N_2855);
or U8475 (N_8475,N_866,N_773);
or U8476 (N_8476,N_4732,N_1657);
or U8477 (N_8477,N_603,N_2324);
nand U8478 (N_8478,N_3363,N_1430);
and U8479 (N_8479,N_3223,N_4394);
nor U8480 (N_8480,N_1489,N_1875);
and U8481 (N_8481,N_349,N_3237);
and U8482 (N_8482,N_1895,N_3796);
xnor U8483 (N_8483,N_2853,N_2589);
nand U8484 (N_8484,N_4283,N_1488);
nor U8485 (N_8485,N_2102,N_997);
and U8486 (N_8486,N_3462,N_553);
or U8487 (N_8487,N_2469,N_1425);
and U8488 (N_8488,N_3542,N_3004);
nor U8489 (N_8489,N_332,N_3837);
nor U8490 (N_8490,N_4728,N_4437);
nand U8491 (N_8491,N_4846,N_2354);
xor U8492 (N_8492,N_3441,N_3821);
nand U8493 (N_8493,N_3378,N_1135);
nor U8494 (N_8494,N_3444,N_1091);
and U8495 (N_8495,N_3545,N_970);
or U8496 (N_8496,N_4111,N_3319);
or U8497 (N_8497,N_1571,N_3548);
nand U8498 (N_8498,N_197,N_1941);
xnor U8499 (N_8499,N_3982,N_4395);
nor U8500 (N_8500,N_4634,N_3727);
and U8501 (N_8501,N_465,N_4934);
nor U8502 (N_8502,N_1093,N_3177);
or U8503 (N_8503,N_3212,N_4241);
or U8504 (N_8504,N_4101,N_3116);
xnor U8505 (N_8505,N_2934,N_2834);
or U8506 (N_8506,N_3759,N_1226);
and U8507 (N_8507,N_379,N_4760);
xnor U8508 (N_8508,N_1686,N_1472);
xnor U8509 (N_8509,N_2138,N_2101);
or U8510 (N_8510,N_86,N_821);
or U8511 (N_8511,N_1448,N_3589);
and U8512 (N_8512,N_3576,N_3755);
and U8513 (N_8513,N_2400,N_4270);
nor U8514 (N_8514,N_3360,N_1114);
nor U8515 (N_8515,N_318,N_364);
nor U8516 (N_8516,N_1737,N_3439);
xnor U8517 (N_8517,N_862,N_354);
or U8518 (N_8518,N_3196,N_1108);
or U8519 (N_8519,N_1525,N_1810);
nand U8520 (N_8520,N_3649,N_854);
nor U8521 (N_8521,N_3271,N_4868);
or U8522 (N_8522,N_4623,N_259);
or U8523 (N_8523,N_4860,N_4300);
or U8524 (N_8524,N_1460,N_312);
and U8525 (N_8525,N_2304,N_2954);
and U8526 (N_8526,N_3266,N_1221);
nor U8527 (N_8527,N_3562,N_1486);
or U8528 (N_8528,N_2075,N_1780);
nor U8529 (N_8529,N_1068,N_629);
xor U8530 (N_8530,N_128,N_1251);
and U8531 (N_8531,N_158,N_4605);
nand U8532 (N_8532,N_3456,N_432);
or U8533 (N_8533,N_1601,N_2578);
xnor U8534 (N_8534,N_3955,N_3162);
and U8535 (N_8535,N_4877,N_4132);
and U8536 (N_8536,N_3528,N_3746);
xor U8537 (N_8537,N_4224,N_782);
or U8538 (N_8538,N_2510,N_115);
and U8539 (N_8539,N_41,N_921);
or U8540 (N_8540,N_3765,N_4850);
nand U8541 (N_8541,N_4399,N_809);
nor U8542 (N_8542,N_453,N_1547);
nand U8543 (N_8543,N_4081,N_1403);
or U8544 (N_8544,N_4323,N_4929);
xnor U8545 (N_8545,N_4805,N_1288);
or U8546 (N_8546,N_2400,N_4828);
nor U8547 (N_8547,N_4618,N_1772);
and U8548 (N_8548,N_4050,N_4268);
and U8549 (N_8549,N_3849,N_522);
or U8550 (N_8550,N_2357,N_4657);
xor U8551 (N_8551,N_786,N_592);
nand U8552 (N_8552,N_564,N_1368);
and U8553 (N_8553,N_2867,N_2577);
and U8554 (N_8554,N_4911,N_1549);
nand U8555 (N_8555,N_2099,N_4586);
xnor U8556 (N_8556,N_1532,N_210);
or U8557 (N_8557,N_2161,N_1360);
or U8558 (N_8558,N_1409,N_4795);
nor U8559 (N_8559,N_3553,N_1632);
and U8560 (N_8560,N_1566,N_1932);
or U8561 (N_8561,N_3396,N_2738);
and U8562 (N_8562,N_2072,N_270);
and U8563 (N_8563,N_3000,N_168);
nand U8564 (N_8564,N_188,N_4513);
xnor U8565 (N_8565,N_602,N_4213);
nand U8566 (N_8566,N_1828,N_3447);
or U8567 (N_8567,N_3371,N_2503);
or U8568 (N_8568,N_3703,N_4298);
and U8569 (N_8569,N_2819,N_632);
nor U8570 (N_8570,N_4365,N_1296);
xor U8571 (N_8571,N_786,N_4451);
xnor U8572 (N_8572,N_2645,N_3978);
or U8573 (N_8573,N_4140,N_866);
nand U8574 (N_8574,N_3469,N_583);
or U8575 (N_8575,N_605,N_4740);
nand U8576 (N_8576,N_14,N_3389);
or U8577 (N_8577,N_3339,N_3976);
nor U8578 (N_8578,N_2828,N_3742);
or U8579 (N_8579,N_1405,N_1565);
nand U8580 (N_8580,N_2528,N_1256);
and U8581 (N_8581,N_4511,N_3377);
nor U8582 (N_8582,N_3617,N_835);
nand U8583 (N_8583,N_1247,N_598);
and U8584 (N_8584,N_4544,N_1645);
nor U8585 (N_8585,N_149,N_488);
nand U8586 (N_8586,N_4053,N_1209);
nand U8587 (N_8587,N_2779,N_173);
nand U8588 (N_8588,N_2630,N_4349);
nand U8589 (N_8589,N_2735,N_110);
nor U8590 (N_8590,N_93,N_3790);
nor U8591 (N_8591,N_3870,N_1962);
nor U8592 (N_8592,N_301,N_2833);
nand U8593 (N_8593,N_4429,N_212);
or U8594 (N_8594,N_1443,N_4351);
nor U8595 (N_8595,N_994,N_3005);
nor U8596 (N_8596,N_355,N_3913);
xnor U8597 (N_8597,N_597,N_4457);
and U8598 (N_8598,N_2519,N_4688);
xor U8599 (N_8599,N_182,N_790);
or U8600 (N_8600,N_2303,N_1435);
nand U8601 (N_8601,N_3617,N_1580);
nor U8602 (N_8602,N_2445,N_3941);
and U8603 (N_8603,N_560,N_4270);
nor U8604 (N_8604,N_3034,N_312);
or U8605 (N_8605,N_4665,N_4082);
or U8606 (N_8606,N_2558,N_4622);
and U8607 (N_8607,N_1038,N_2850);
nor U8608 (N_8608,N_4973,N_2518);
and U8609 (N_8609,N_2772,N_2876);
nand U8610 (N_8610,N_3067,N_2626);
nand U8611 (N_8611,N_4245,N_1286);
nand U8612 (N_8612,N_4040,N_3053);
and U8613 (N_8613,N_4765,N_4658);
nor U8614 (N_8614,N_1676,N_3187);
or U8615 (N_8615,N_527,N_3869);
and U8616 (N_8616,N_2000,N_2411);
or U8617 (N_8617,N_1886,N_4373);
nand U8618 (N_8618,N_2064,N_4807);
or U8619 (N_8619,N_1744,N_3830);
and U8620 (N_8620,N_1990,N_2616);
or U8621 (N_8621,N_1957,N_1355);
and U8622 (N_8622,N_1844,N_445);
and U8623 (N_8623,N_3867,N_2230);
and U8624 (N_8624,N_2820,N_4650);
and U8625 (N_8625,N_991,N_658);
xnor U8626 (N_8626,N_1551,N_1194);
and U8627 (N_8627,N_1287,N_4669);
nand U8628 (N_8628,N_1298,N_252);
nand U8629 (N_8629,N_917,N_3145);
nand U8630 (N_8630,N_1910,N_3126);
nand U8631 (N_8631,N_3108,N_4836);
nand U8632 (N_8632,N_789,N_558);
nor U8633 (N_8633,N_3003,N_3431);
and U8634 (N_8634,N_129,N_1447);
nor U8635 (N_8635,N_3232,N_1201);
xnor U8636 (N_8636,N_4045,N_383);
nor U8637 (N_8637,N_3991,N_835);
or U8638 (N_8638,N_2361,N_737);
and U8639 (N_8639,N_4228,N_3040);
and U8640 (N_8640,N_2799,N_238);
or U8641 (N_8641,N_4195,N_245);
and U8642 (N_8642,N_4652,N_1879);
xnor U8643 (N_8643,N_3036,N_4913);
or U8644 (N_8644,N_4116,N_634);
or U8645 (N_8645,N_2480,N_3149);
nand U8646 (N_8646,N_199,N_561);
nor U8647 (N_8647,N_4782,N_3376);
xnor U8648 (N_8648,N_44,N_1761);
nand U8649 (N_8649,N_99,N_1931);
and U8650 (N_8650,N_4358,N_1466);
or U8651 (N_8651,N_255,N_14);
nand U8652 (N_8652,N_271,N_4167);
nand U8653 (N_8653,N_2361,N_4871);
or U8654 (N_8654,N_1605,N_623);
and U8655 (N_8655,N_4379,N_4213);
nor U8656 (N_8656,N_648,N_3570);
nor U8657 (N_8657,N_3403,N_4599);
and U8658 (N_8658,N_1509,N_2552);
nand U8659 (N_8659,N_2491,N_2050);
nor U8660 (N_8660,N_3547,N_2686);
xor U8661 (N_8661,N_2673,N_2183);
nand U8662 (N_8662,N_4298,N_2340);
and U8663 (N_8663,N_2020,N_3108);
nor U8664 (N_8664,N_680,N_1060);
and U8665 (N_8665,N_3230,N_4680);
nand U8666 (N_8666,N_4480,N_1512);
and U8667 (N_8667,N_3198,N_2898);
nor U8668 (N_8668,N_1332,N_1101);
or U8669 (N_8669,N_3294,N_3269);
nand U8670 (N_8670,N_26,N_2710);
xor U8671 (N_8671,N_1630,N_4842);
or U8672 (N_8672,N_1549,N_3765);
xnor U8673 (N_8673,N_4426,N_2386);
nor U8674 (N_8674,N_4610,N_214);
or U8675 (N_8675,N_335,N_2095);
and U8676 (N_8676,N_4347,N_2083);
or U8677 (N_8677,N_1125,N_4112);
or U8678 (N_8678,N_1835,N_2149);
nor U8679 (N_8679,N_3065,N_2994);
xor U8680 (N_8680,N_4613,N_4063);
nand U8681 (N_8681,N_3163,N_1848);
nor U8682 (N_8682,N_298,N_1415);
or U8683 (N_8683,N_4459,N_1857);
or U8684 (N_8684,N_717,N_4645);
nand U8685 (N_8685,N_2592,N_439);
nor U8686 (N_8686,N_4550,N_4720);
and U8687 (N_8687,N_4582,N_3731);
nand U8688 (N_8688,N_1297,N_4852);
or U8689 (N_8689,N_2785,N_1497);
and U8690 (N_8690,N_3903,N_2658);
and U8691 (N_8691,N_4262,N_2547);
nand U8692 (N_8692,N_4924,N_106);
nor U8693 (N_8693,N_344,N_2785);
or U8694 (N_8694,N_4124,N_4221);
or U8695 (N_8695,N_1239,N_1270);
nand U8696 (N_8696,N_1923,N_2671);
nand U8697 (N_8697,N_3500,N_1697);
or U8698 (N_8698,N_2248,N_2707);
nor U8699 (N_8699,N_4081,N_885);
or U8700 (N_8700,N_4844,N_2873);
and U8701 (N_8701,N_1929,N_3563);
and U8702 (N_8702,N_4552,N_985);
or U8703 (N_8703,N_4882,N_3377);
nand U8704 (N_8704,N_2334,N_56);
nand U8705 (N_8705,N_4826,N_4779);
or U8706 (N_8706,N_4390,N_2293);
nor U8707 (N_8707,N_4832,N_499);
and U8708 (N_8708,N_4751,N_3258);
nor U8709 (N_8709,N_4100,N_1583);
xor U8710 (N_8710,N_3980,N_1262);
and U8711 (N_8711,N_1507,N_190);
nand U8712 (N_8712,N_3930,N_3596);
nor U8713 (N_8713,N_3281,N_3230);
nor U8714 (N_8714,N_1377,N_4040);
or U8715 (N_8715,N_3412,N_1693);
nor U8716 (N_8716,N_1796,N_234);
nand U8717 (N_8717,N_1409,N_4502);
nor U8718 (N_8718,N_4772,N_2913);
or U8719 (N_8719,N_3985,N_1181);
and U8720 (N_8720,N_1852,N_1091);
nand U8721 (N_8721,N_2109,N_4335);
nor U8722 (N_8722,N_4535,N_1572);
nand U8723 (N_8723,N_2668,N_2200);
and U8724 (N_8724,N_3947,N_4441);
nor U8725 (N_8725,N_2444,N_1032);
nand U8726 (N_8726,N_65,N_2270);
and U8727 (N_8727,N_2608,N_3615);
nand U8728 (N_8728,N_3261,N_2195);
nand U8729 (N_8729,N_2247,N_2715);
nand U8730 (N_8730,N_3820,N_943);
or U8731 (N_8731,N_2332,N_3434);
nor U8732 (N_8732,N_4905,N_4812);
and U8733 (N_8733,N_3088,N_348);
or U8734 (N_8734,N_3532,N_437);
or U8735 (N_8735,N_4146,N_2440);
or U8736 (N_8736,N_4040,N_4274);
xor U8737 (N_8737,N_2060,N_2683);
and U8738 (N_8738,N_1450,N_3842);
or U8739 (N_8739,N_2119,N_1067);
xor U8740 (N_8740,N_3555,N_687);
xor U8741 (N_8741,N_112,N_1499);
nand U8742 (N_8742,N_720,N_627);
and U8743 (N_8743,N_2119,N_4482);
nor U8744 (N_8744,N_4060,N_2135);
nand U8745 (N_8745,N_3336,N_3825);
or U8746 (N_8746,N_1049,N_2454);
or U8747 (N_8747,N_1142,N_969);
or U8748 (N_8748,N_682,N_626);
or U8749 (N_8749,N_2997,N_2683);
nor U8750 (N_8750,N_1000,N_3123);
nand U8751 (N_8751,N_4791,N_1828);
nand U8752 (N_8752,N_4351,N_2534);
nand U8753 (N_8753,N_362,N_2411);
and U8754 (N_8754,N_3288,N_4678);
and U8755 (N_8755,N_1942,N_4796);
or U8756 (N_8756,N_478,N_4236);
or U8757 (N_8757,N_3885,N_3201);
and U8758 (N_8758,N_1864,N_2401);
or U8759 (N_8759,N_1282,N_1797);
or U8760 (N_8760,N_81,N_4015);
nor U8761 (N_8761,N_1611,N_2612);
nand U8762 (N_8762,N_1630,N_1234);
and U8763 (N_8763,N_798,N_1421);
and U8764 (N_8764,N_1430,N_2617);
xor U8765 (N_8765,N_1030,N_856);
nand U8766 (N_8766,N_2572,N_1976);
nor U8767 (N_8767,N_4442,N_2736);
or U8768 (N_8768,N_501,N_3425);
or U8769 (N_8769,N_3028,N_4471);
nor U8770 (N_8770,N_1608,N_49);
nand U8771 (N_8771,N_813,N_2179);
xor U8772 (N_8772,N_4068,N_2431);
nand U8773 (N_8773,N_748,N_1066);
xor U8774 (N_8774,N_4900,N_3021);
xor U8775 (N_8775,N_2472,N_1923);
or U8776 (N_8776,N_180,N_913);
nand U8777 (N_8777,N_1125,N_1120);
nor U8778 (N_8778,N_3659,N_1799);
xnor U8779 (N_8779,N_2897,N_3259);
nand U8780 (N_8780,N_3826,N_4895);
or U8781 (N_8781,N_3422,N_4578);
or U8782 (N_8782,N_3504,N_3096);
nand U8783 (N_8783,N_2632,N_1613);
xor U8784 (N_8784,N_81,N_3323);
nor U8785 (N_8785,N_4283,N_4471);
nand U8786 (N_8786,N_1389,N_2454);
nand U8787 (N_8787,N_1710,N_1003);
xor U8788 (N_8788,N_4243,N_1587);
nor U8789 (N_8789,N_4660,N_3960);
nor U8790 (N_8790,N_2126,N_336);
or U8791 (N_8791,N_1194,N_3041);
and U8792 (N_8792,N_1531,N_1157);
or U8793 (N_8793,N_4112,N_2572);
nand U8794 (N_8794,N_2108,N_3121);
or U8795 (N_8795,N_1197,N_2659);
or U8796 (N_8796,N_2229,N_2690);
and U8797 (N_8797,N_3423,N_3993);
nor U8798 (N_8798,N_4891,N_120);
nand U8799 (N_8799,N_2766,N_4831);
nand U8800 (N_8800,N_2370,N_1601);
nand U8801 (N_8801,N_3871,N_3282);
nor U8802 (N_8802,N_3711,N_872);
nor U8803 (N_8803,N_192,N_1624);
or U8804 (N_8804,N_2584,N_4208);
or U8805 (N_8805,N_758,N_2999);
nor U8806 (N_8806,N_2604,N_1126);
or U8807 (N_8807,N_2881,N_2104);
nand U8808 (N_8808,N_2327,N_3217);
or U8809 (N_8809,N_1439,N_3082);
xor U8810 (N_8810,N_2341,N_4847);
and U8811 (N_8811,N_3347,N_3454);
or U8812 (N_8812,N_2525,N_1137);
and U8813 (N_8813,N_2415,N_2244);
and U8814 (N_8814,N_4972,N_1081);
or U8815 (N_8815,N_4573,N_2812);
nand U8816 (N_8816,N_2488,N_1570);
xor U8817 (N_8817,N_1075,N_3521);
nor U8818 (N_8818,N_2597,N_4249);
xor U8819 (N_8819,N_2888,N_3904);
or U8820 (N_8820,N_3673,N_145);
and U8821 (N_8821,N_3154,N_3614);
and U8822 (N_8822,N_3090,N_4386);
and U8823 (N_8823,N_874,N_1490);
nand U8824 (N_8824,N_3826,N_2066);
nor U8825 (N_8825,N_4930,N_4295);
nor U8826 (N_8826,N_4220,N_1777);
and U8827 (N_8827,N_212,N_4621);
or U8828 (N_8828,N_3438,N_4856);
or U8829 (N_8829,N_1165,N_2800);
nor U8830 (N_8830,N_3035,N_3481);
or U8831 (N_8831,N_1507,N_2113);
and U8832 (N_8832,N_2960,N_2321);
and U8833 (N_8833,N_3675,N_628);
and U8834 (N_8834,N_3774,N_551);
nand U8835 (N_8835,N_4010,N_4932);
nor U8836 (N_8836,N_593,N_2898);
nand U8837 (N_8837,N_2835,N_2729);
or U8838 (N_8838,N_2666,N_895);
or U8839 (N_8839,N_2955,N_484);
nor U8840 (N_8840,N_3826,N_1279);
nand U8841 (N_8841,N_1985,N_1023);
and U8842 (N_8842,N_411,N_4995);
or U8843 (N_8843,N_3944,N_2581);
or U8844 (N_8844,N_575,N_2927);
nand U8845 (N_8845,N_1282,N_711);
or U8846 (N_8846,N_2759,N_1697);
or U8847 (N_8847,N_3101,N_2813);
nand U8848 (N_8848,N_2824,N_1087);
xor U8849 (N_8849,N_2245,N_257);
and U8850 (N_8850,N_3082,N_1608);
and U8851 (N_8851,N_3082,N_1972);
and U8852 (N_8852,N_1264,N_4366);
nor U8853 (N_8853,N_3241,N_160);
nor U8854 (N_8854,N_3005,N_4861);
or U8855 (N_8855,N_2685,N_1506);
nand U8856 (N_8856,N_1572,N_1183);
and U8857 (N_8857,N_2862,N_332);
xnor U8858 (N_8858,N_267,N_3664);
xor U8859 (N_8859,N_1697,N_2293);
nor U8860 (N_8860,N_1553,N_2397);
and U8861 (N_8861,N_4703,N_1947);
nand U8862 (N_8862,N_2964,N_2655);
and U8863 (N_8863,N_1640,N_1564);
and U8864 (N_8864,N_3641,N_3491);
nand U8865 (N_8865,N_9,N_3358);
nand U8866 (N_8866,N_678,N_3669);
and U8867 (N_8867,N_3681,N_143);
and U8868 (N_8868,N_2124,N_1874);
and U8869 (N_8869,N_3798,N_2617);
or U8870 (N_8870,N_1255,N_4027);
nand U8871 (N_8871,N_1343,N_674);
nand U8872 (N_8872,N_2183,N_2010);
nor U8873 (N_8873,N_3731,N_3953);
nand U8874 (N_8874,N_3983,N_2945);
nand U8875 (N_8875,N_4458,N_2376);
or U8876 (N_8876,N_4324,N_3620);
nor U8877 (N_8877,N_1489,N_2724);
nor U8878 (N_8878,N_4362,N_862);
or U8879 (N_8879,N_3757,N_1127);
and U8880 (N_8880,N_2204,N_2807);
nor U8881 (N_8881,N_963,N_2867);
nand U8882 (N_8882,N_446,N_4898);
or U8883 (N_8883,N_3025,N_4995);
nor U8884 (N_8884,N_1425,N_2528);
and U8885 (N_8885,N_3825,N_2021);
or U8886 (N_8886,N_1012,N_2771);
nand U8887 (N_8887,N_1202,N_2941);
nor U8888 (N_8888,N_2730,N_1435);
and U8889 (N_8889,N_3552,N_4727);
and U8890 (N_8890,N_2135,N_4452);
or U8891 (N_8891,N_1361,N_1510);
or U8892 (N_8892,N_632,N_4094);
and U8893 (N_8893,N_4332,N_3545);
nor U8894 (N_8894,N_1365,N_4187);
nor U8895 (N_8895,N_3457,N_3394);
xnor U8896 (N_8896,N_3455,N_3884);
nor U8897 (N_8897,N_3221,N_1779);
and U8898 (N_8898,N_3324,N_1423);
xnor U8899 (N_8899,N_799,N_317);
and U8900 (N_8900,N_4188,N_1825);
nand U8901 (N_8901,N_4667,N_4529);
nor U8902 (N_8902,N_2416,N_2935);
nand U8903 (N_8903,N_2969,N_4639);
nor U8904 (N_8904,N_1623,N_2450);
or U8905 (N_8905,N_1589,N_2735);
or U8906 (N_8906,N_3515,N_958);
nand U8907 (N_8907,N_1816,N_919);
and U8908 (N_8908,N_4766,N_1309);
and U8909 (N_8909,N_2072,N_4242);
nand U8910 (N_8910,N_2196,N_1300);
nor U8911 (N_8911,N_916,N_4159);
or U8912 (N_8912,N_1825,N_4916);
and U8913 (N_8913,N_585,N_2266);
and U8914 (N_8914,N_1066,N_2979);
and U8915 (N_8915,N_3540,N_1529);
nor U8916 (N_8916,N_2668,N_3751);
nand U8917 (N_8917,N_553,N_3994);
or U8918 (N_8918,N_2078,N_3768);
nand U8919 (N_8919,N_4935,N_3336);
and U8920 (N_8920,N_1593,N_3570);
and U8921 (N_8921,N_3841,N_3735);
or U8922 (N_8922,N_1678,N_2599);
xnor U8923 (N_8923,N_4226,N_4119);
nor U8924 (N_8924,N_277,N_4623);
nand U8925 (N_8925,N_4622,N_1693);
and U8926 (N_8926,N_224,N_1694);
and U8927 (N_8927,N_3421,N_4760);
xnor U8928 (N_8928,N_4168,N_2785);
and U8929 (N_8929,N_2160,N_3538);
xnor U8930 (N_8930,N_2137,N_1826);
nor U8931 (N_8931,N_740,N_44);
and U8932 (N_8932,N_1096,N_4843);
or U8933 (N_8933,N_4710,N_4199);
nand U8934 (N_8934,N_724,N_2767);
or U8935 (N_8935,N_1950,N_4591);
nand U8936 (N_8936,N_4846,N_214);
nor U8937 (N_8937,N_3757,N_4340);
nor U8938 (N_8938,N_3221,N_3667);
or U8939 (N_8939,N_10,N_170);
and U8940 (N_8940,N_3842,N_3844);
nor U8941 (N_8941,N_2514,N_4430);
and U8942 (N_8942,N_3155,N_2594);
or U8943 (N_8943,N_3673,N_4362);
nor U8944 (N_8944,N_2807,N_661);
and U8945 (N_8945,N_454,N_1854);
nand U8946 (N_8946,N_4239,N_1707);
nand U8947 (N_8947,N_3026,N_1934);
xnor U8948 (N_8948,N_337,N_2689);
nand U8949 (N_8949,N_3168,N_4541);
or U8950 (N_8950,N_4396,N_999);
and U8951 (N_8951,N_1794,N_222);
nand U8952 (N_8952,N_1127,N_1133);
nor U8953 (N_8953,N_4295,N_4332);
or U8954 (N_8954,N_4944,N_3039);
and U8955 (N_8955,N_3406,N_543);
nand U8956 (N_8956,N_1589,N_596);
nor U8957 (N_8957,N_1533,N_1200);
or U8958 (N_8958,N_277,N_2107);
nor U8959 (N_8959,N_4175,N_1334);
nand U8960 (N_8960,N_1517,N_1478);
nor U8961 (N_8961,N_2442,N_1644);
and U8962 (N_8962,N_3863,N_2621);
and U8963 (N_8963,N_4422,N_3218);
or U8964 (N_8964,N_284,N_2904);
nor U8965 (N_8965,N_3017,N_3817);
nor U8966 (N_8966,N_4854,N_3729);
or U8967 (N_8967,N_904,N_4096);
nand U8968 (N_8968,N_417,N_88);
nor U8969 (N_8969,N_1298,N_2921);
and U8970 (N_8970,N_2489,N_4828);
and U8971 (N_8971,N_540,N_2364);
xnor U8972 (N_8972,N_2732,N_4179);
xor U8973 (N_8973,N_2772,N_4806);
or U8974 (N_8974,N_3330,N_1780);
nor U8975 (N_8975,N_3583,N_1019);
nor U8976 (N_8976,N_222,N_3639);
and U8977 (N_8977,N_337,N_937);
nand U8978 (N_8978,N_369,N_2389);
and U8979 (N_8979,N_3179,N_4940);
and U8980 (N_8980,N_159,N_4216);
xnor U8981 (N_8981,N_674,N_4725);
or U8982 (N_8982,N_492,N_3721);
nand U8983 (N_8983,N_3185,N_2502);
or U8984 (N_8984,N_1859,N_2674);
or U8985 (N_8985,N_4691,N_4197);
nor U8986 (N_8986,N_3074,N_1312);
nor U8987 (N_8987,N_909,N_3612);
nor U8988 (N_8988,N_4587,N_3785);
or U8989 (N_8989,N_3169,N_2085);
or U8990 (N_8990,N_3353,N_4443);
xnor U8991 (N_8991,N_1037,N_4628);
nand U8992 (N_8992,N_4008,N_3640);
or U8993 (N_8993,N_513,N_2989);
or U8994 (N_8994,N_3050,N_2542);
or U8995 (N_8995,N_3121,N_3634);
nor U8996 (N_8996,N_3291,N_4349);
nand U8997 (N_8997,N_1359,N_3754);
nand U8998 (N_8998,N_2667,N_2056);
or U8999 (N_8999,N_2398,N_3049);
nor U9000 (N_9000,N_3521,N_71);
or U9001 (N_9001,N_43,N_2343);
or U9002 (N_9002,N_842,N_1456);
and U9003 (N_9003,N_1604,N_2696);
and U9004 (N_9004,N_673,N_2243);
nand U9005 (N_9005,N_808,N_4148);
nand U9006 (N_9006,N_1102,N_4582);
nand U9007 (N_9007,N_3304,N_2897);
nor U9008 (N_9008,N_4323,N_726);
nand U9009 (N_9009,N_1684,N_3983);
nand U9010 (N_9010,N_2339,N_1939);
nand U9011 (N_9011,N_3613,N_763);
nor U9012 (N_9012,N_2696,N_1784);
nand U9013 (N_9013,N_2565,N_2305);
nor U9014 (N_9014,N_4626,N_4029);
nand U9015 (N_9015,N_596,N_2008);
or U9016 (N_9016,N_203,N_1241);
nand U9017 (N_9017,N_1321,N_1205);
or U9018 (N_9018,N_2508,N_1334);
and U9019 (N_9019,N_3604,N_3814);
or U9020 (N_9020,N_2034,N_1019);
xnor U9021 (N_9021,N_3181,N_3188);
and U9022 (N_9022,N_4553,N_2088);
nand U9023 (N_9023,N_4768,N_4818);
or U9024 (N_9024,N_745,N_3111);
nor U9025 (N_9025,N_3410,N_115);
or U9026 (N_9026,N_3603,N_2793);
nand U9027 (N_9027,N_3615,N_215);
nand U9028 (N_9028,N_2703,N_4889);
and U9029 (N_9029,N_4564,N_4672);
nand U9030 (N_9030,N_3005,N_2531);
nand U9031 (N_9031,N_4340,N_2837);
and U9032 (N_9032,N_2707,N_4741);
and U9033 (N_9033,N_762,N_2067);
nand U9034 (N_9034,N_2249,N_1358);
nor U9035 (N_9035,N_1519,N_1728);
and U9036 (N_9036,N_3290,N_3680);
nor U9037 (N_9037,N_310,N_4685);
nor U9038 (N_9038,N_4384,N_1160);
and U9039 (N_9039,N_4096,N_1258);
and U9040 (N_9040,N_2002,N_3996);
nor U9041 (N_9041,N_1270,N_2079);
and U9042 (N_9042,N_1017,N_4411);
and U9043 (N_9043,N_1967,N_674);
nor U9044 (N_9044,N_1415,N_4682);
xnor U9045 (N_9045,N_1195,N_4615);
and U9046 (N_9046,N_3934,N_609);
and U9047 (N_9047,N_3166,N_2127);
nor U9048 (N_9048,N_1343,N_4109);
nand U9049 (N_9049,N_4170,N_558);
and U9050 (N_9050,N_2593,N_4406);
nand U9051 (N_9051,N_3878,N_2102);
or U9052 (N_9052,N_866,N_108);
nor U9053 (N_9053,N_2561,N_587);
or U9054 (N_9054,N_3220,N_1464);
nand U9055 (N_9055,N_2913,N_3521);
nor U9056 (N_9056,N_1897,N_2380);
or U9057 (N_9057,N_1951,N_1136);
nand U9058 (N_9058,N_4327,N_3615);
nand U9059 (N_9059,N_4254,N_420);
and U9060 (N_9060,N_4364,N_2537);
and U9061 (N_9061,N_2610,N_2343);
nand U9062 (N_9062,N_290,N_4329);
nor U9063 (N_9063,N_3113,N_3234);
and U9064 (N_9064,N_1683,N_503);
or U9065 (N_9065,N_3939,N_4076);
nand U9066 (N_9066,N_3747,N_3024);
or U9067 (N_9067,N_51,N_3396);
nand U9068 (N_9068,N_2590,N_4467);
and U9069 (N_9069,N_2144,N_4259);
nand U9070 (N_9070,N_546,N_3728);
and U9071 (N_9071,N_386,N_3944);
nand U9072 (N_9072,N_375,N_2636);
or U9073 (N_9073,N_796,N_1200);
nor U9074 (N_9074,N_4864,N_2418);
nor U9075 (N_9075,N_3206,N_4152);
nor U9076 (N_9076,N_4083,N_2527);
or U9077 (N_9077,N_4821,N_3984);
or U9078 (N_9078,N_2499,N_4039);
xor U9079 (N_9079,N_4229,N_4749);
xor U9080 (N_9080,N_1925,N_914);
and U9081 (N_9081,N_1635,N_1747);
nor U9082 (N_9082,N_10,N_770);
nor U9083 (N_9083,N_3825,N_260);
and U9084 (N_9084,N_932,N_3833);
xor U9085 (N_9085,N_888,N_3434);
or U9086 (N_9086,N_2571,N_1974);
nand U9087 (N_9087,N_1427,N_4159);
nor U9088 (N_9088,N_345,N_522);
xor U9089 (N_9089,N_309,N_3970);
or U9090 (N_9090,N_1274,N_1645);
nand U9091 (N_9091,N_4014,N_4107);
or U9092 (N_9092,N_3601,N_680);
and U9093 (N_9093,N_1661,N_3734);
or U9094 (N_9094,N_4424,N_4643);
nand U9095 (N_9095,N_3713,N_2733);
or U9096 (N_9096,N_4768,N_2808);
or U9097 (N_9097,N_2343,N_1965);
nand U9098 (N_9098,N_502,N_1118);
and U9099 (N_9099,N_4912,N_1775);
nor U9100 (N_9100,N_1938,N_4791);
and U9101 (N_9101,N_2487,N_2869);
nand U9102 (N_9102,N_995,N_3638);
nor U9103 (N_9103,N_4279,N_3874);
nand U9104 (N_9104,N_1185,N_1105);
or U9105 (N_9105,N_3582,N_1410);
and U9106 (N_9106,N_34,N_3832);
nand U9107 (N_9107,N_350,N_3109);
and U9108 (N_9108,N_1951,N_3270);
nor U9109 (N_9109,N_4252,N_3619);
nand U9110 (N_9110,N_4925,N_1383);
or U9111 (N_9111,N_2606,N_4943);
nand U9112 (N_9112,N_3804,N_3510);
nor U9113 (N_9113,N_659,N_2383);
nand U9114 (N_9114,N_373,N_3423);
or U9115 (N_9115,N_4236,N_3834);
or U9116 (N_9116,N_4402,N_3876);
or U9117 (N_9117,N_2469,N_1850);
and U9118 (N_9118,N_890,N_3186);
nor U9119 (N_9119,N_4224,N_734);
or U9120 (N_9120,N_1481,N_4753);
and U9121 (N_9121,N_2952,N_1455);
and U9122 (N_9122,N_3144,N_3050);
and U9123 (N_9123,N_4102,N_4378);
nand U9124 (N_9124,N_485,N_2072);
or U9125 (N_9125,N_4375,N_2995);
or U9126 (N_9126,N_1584,N_4441);
and U9127 (N_9127,N_1950,N_36);
nand U9128 (N_9128,N_3480,N_4237);
nor U9129 (N_9129,N_3295,N_4643);
nand U9130 (N_9130,N_423,N_3782);
nand U9131 (N_9131,N_3538,N_831);
and U9132 (N_9132,N_224,N_1510);
nand U9133 (N_9133,N_4964,N_2200);
nand U9134 (N_9134,N_2345,N_4108);
or U9135 (N_9135,N_2248,N_653);
and U9136 (N_9136,N_2378,N_949);
or U9137 (N_9137,N_119,N_4209);
nand U9138 (N_9138,N_766,N_866);
or U9139 (N_9139,N_382,N_4090);
xor U9140 (N_9140,N_1817,N_862);
nand U9141 (N_9141,N_4018,N_734);
nand U9142 (N_9142,N_4646,N_1124);
nand U9143 (N_9143,N_636,N_4334);
nand U9144 (N_9144,N_4081,N_3859);
nor U9145 (N_9145,N_4496,N_1315);
nand U9146 (N_9146,N_2464,N_477);
and U9147 (N_9147,N_483,N_4417);
nor U9148 (N_9148,N_4446,N_4656);
xor U9149 (N_9149,N_3901,N_4460);
nor U9150 (N_9150,N_998,N_2519);
nand U9151 (N_9151,N_2662,N_3099);
nor U9152 (N_9152,N_1238,N_3392);
nor U9153 (N_9153,N_2094,N_4446);
nand U9154 (N_9154,N_3654,N_4873);
nor U9155 (N_9155,N_3060,N_4018);
and U9156 (N_9156,N_1186,N_773);
nand U9157 (N_9157,N_4413,N_720);
xnor U9158 (N_9158,N_2198,N_2418);
nor U9159 (N_9159,N_2813,N_3331);
or U9160 (N_9160,N_589,N_3259);
nor U9161 (N_9161,N_2712,N_3995);
xor U9162 (N_9162,N_1100,N_467);
nor U9163 (N_9163,N_2789,N_4362);
nor U9164 (N_9164,N_1477,N_4562);
nor U9165 (N_9165,N_1305,N_2726);
and U9166 (N_9166,N_2349,N_299);
or U9167 (N_9167,N_3555,N_883);
or U9168 (N_9168,N_4789,N_2479);
nor U9169 (N_9169,N_369,N_3944);
or U9170 (N_9170,N_405,N_461);
or U9171 (N_9171,N_4835,N_3001);
or U9172 (N_9172,N_1615,N_43);
nor U9173 (N_9173,N_2213,N_868);
xnor U9174 (N_9174,N_2300,N_2959);
and U9175 (N_9175,N_889,N_1478);
nand U9176 (N_9176,N_4482,N_896);
or U9177 (N_9177,N_1904,N_3614);
xor U9178 (N_9178,N_4017,N_1943);
nor U9179 (N_9179,N_1395,N_4646);
nand U9180 (N_9180,N_2769,N_1510);
nor U9181 (N_9181,N_4997,N_120);
nor U9182 (N_9182,N_3687,N_2284);
or U9183 (N_9183,N_2063,N_1917);
xor U9184 (N_9184,N_3760,N_3972);
or U9185 (N_9185,N_434,N_1325);
or U9186 (N_9186,N_1045,N_1023);
nand U9187 (N_9187,N_4986,N_2571);
or U9188 (N_9188,N_1154,N_4997);
or U9189 (N_9189,N_2243,N_2822);
or U9190 (N_9190,N_352,N_3957);
nor U9191 (N_9191,N_2951,N_235);
xnor U9192 (N_9192,N_1353,N_410);
and U9193 (N_9193,N_4360,N_2867);
and U9194 (N_9194,N_4983,N_179);
nand U9195 (N_9195,N_3967,N_4824);
and U9196 (N_9196,N_2701,N_4709);
nand U9197 (N_9197,N_4710,N_3837);
nand U9198 (N_9198,N_4432,N_4225);
nor U9199 (N_9199,N_4234,N_4630);
nor U9200 (N_9200,N_1276,N_1409);
and U9201 (N_9201,N_4070,N_2213);
nand U9202 (N_9202,N_1633,N_3865);
nand U9203 (N_9203,N_1694,N_28);
nand U9204 (N_9204,N_2474,N_1718);
nand U9205 (N_9205,N_2440,N_4735);
and U9206 (N_9206,N_3062,N_3479);
nand U9207 (N_9207,N_2676,N_1264);
and U9208 (N_9208,N_4235,N_4975);
nor U9209 (N_9209,N_2380,N_1160);
nor U9210 (N_9210,N_4382,N_2145);
or U9211 (N_9211,N_3071,N_2842);
xor U9212 (N_9212,N_1136,N_1970);
or U9213 (N_9213,N_3998,N_2903);
and U9214 (N_9214,N_4188,N_2697);
nand U9215 (N_9215,N_4627,N_4917);
nor U9216 (N_9216,N_2115,N_1172);
and U9217 (N_9217,N_3715,N_426);
nand U9218 (N_9218,N_2028,N_1776);
nand U9219 (N_9219,N_2700,N_3355);
or U9220 (N_9220,N_3982,N_3055);
and U9221 (N_9221,N_3102,N_797);
and U9222 (N_9222,N_3562,N_266);
and U9223 (N_9223,N_628,N_4265);
nor U9224 (N_9224,N_322,N_2580);
or U9225 (N_9225,N_1222,N_148);
or U9226 (N_9226,N_4076,N_446);
xnor U9227 (N_9227,N_3409,N_1543);
or U9228 (N_9228,N_3081,N_4954);
or U9229 (N_9229,N_1130,N_763);
and U9230 (N_9230,N_3299,N_4884);
and U9231 (N_9231,N_1338,N_4579);
or U9232 (N_9232,N_2328,N_653);
nor U9233 (N_9233,N_1656,N_2631);
and U9234 (N_9234,N_4249,N_118);
nor U9235 (N_9235,N_3509,N_1723);
or U9236 (N_9236,N_428,N_1234);
or U9237 (N_9237,N_725,N_654);
or U9238 (N_9238,N_4676,N_1037);
xor U9239 (N_9239,N_2611,N_4521);
xnor U9240 (N_9240,N_1902,N_867);
and U9241 (N_9241,N_1388,N_1210);
xnor U9242 (N_9242,N_117,N_4973);
and U9243 (N_9243,N_3605,N_4848);
nand U9244 (N_9244,N_1649,N_416);
nand U9245 (N_9245,N_4237,N_3784);
nand U9246 (N_9246,N_2304,N_473);
xnor U9247 (N_9247,N_832,N_687);
nand U9248 (N_9248,N_2178,N_4183);
or U9249 (N_9249,N_3852,N_3272);
and U9250 (N_9250,N_413,N_2434);
and U9251 (N_9251,N_2701,N_2644);
nand U9252 (N_9252,N_4444,N_3227);
nor U9253 (N_9253,N_1864,N_4723);
and U9254 (N_9254,N_3928,N_3245);
nor U9255 (N_9255,N_2552,N_3718);
nor U9256 (N_9256,N_4825,N_1989);
nand U9257 (N_9257,N_3408,N_1962);
and U9258 (N_9258,N_2616,N_3674);
nand U9259 (N_9259,N_2337,N_3932);
or U9260 (N_9260,N_4468,N_4958);
or U9261 (N_9261,N_1659,N_2572);
nor U9262 (N_9262,N_4584,N_1882);
nor U9263 (N_9263,N_4785,N_4294);
nand U9264 (N_9264,N_739,N_854);
xnor U9265 (N_9265,N_1247,N_4635);
nor U9266 (N_9266,N_3261,N_4846);
and U9267 (N_9267,N_2074,N_4628);
or U9268 (N_9268,N_995,N_3476);
and U9269 (N_9269,N_3489,N_389);
nor U9270 (N_9270,N_4306,N_90);
nor U9271 (N_9271,N_2811,N_1670);
and U9272 (N_9272,N_2954,N_2330);
nand U9273 (N_9273,N_1102,N_1898);
nor U9274 (N_9274,N_1449,N_4207);
nand U9275 (N_9275,N_469,N_3302);
and U9276 (N_9276,N_2684,N_968);
or U9277 (N_9277,N_454,N_4167);
and U9278 (N_9278,N_21,N_2195);
xnor U9279 (N_9279,N_904,N_3023);
xor U9280 (N_9280,N_1474,N_743);
and U9281 (N_9281,N_4328,N_3341);
or U9282 (N_9282,N_2794,N_2235);
or U9283 (N_9283,N_3854,N_543);
nand U9284 (N_9284,N_2281,N_1851);
and U9285 (N_9285,N_4357,N_304);
nor U9286 (N_9286,N_3239,N_1011);
nor U9287 (N_9287,N_586,N_4113);
nor U9288 (N_9288,N_4619,N_4293);
nand U9289 (N_9289,N_807,N_33);
and U9290 (N_9290,N_2212,N_1172);
or U9291 (N_9291,N_2828,N_676);
xor U9292 (N_9292,N_1489,N_514);
and U9293 (N_9293,N_4074,N_2533);
and U9294 (N_9294,N_1086,N_3166);
or U9295 (N_9295,N_2915,N_1005);
xor U9296 (N_9296,N_113,N_3954);
and U9297 (N_9297,N_4391,N_2123);
nand U9298 (N_9298,N_4051,N_161);
xor U9299 (N_9299,N_457,N_392);
nand U9300 (N_9300,N_856,N_4697);
nor U9301 (N_9301,N_1317,N_824);
and U9302 (N_9302,N_3782,N_2887);
nand U9303 (N_9303,N_1370,N_2010);
nand U9304 (N_9304,N_4872,N_2947);
nand U9305 (N_9305,N_939,N_2361);
nor U9306 (N_9306,N_1439,N_1040);
and U9307 (N_9307,N_2118,N_4970);
or U9308 (N_9308,N_529,N_72);
nor U9309 (N_9309,N_2270,N_260);
and U9310 (N_9310,N_670,N_3221);
xnor U9311 (N_9311,N_4973,N_562);
and U9312 (N_9312,N_1480,N_1949);
nor U9313 (N_9313,N_835,N_2165);
or U9314 (N_9314,N_857,N_4990);
or U9315 (N_9315,N_3495,N_4773);
nor U9316 (N_9316,N_1068,N_665);
nand U9317 (N_9317,N_421,N_4336);
and U9318 (N_9318,N_2010,N_4028);
or U9319 (N_9319,N_3964,N_4964);
or U9320 (N_9320,N_1558,N_2552);
or U9321 (N_9321,N_2383,N_1560);
and U9322 (N_9322,N_4351,N_535);
xor U9323 (N_9323,N_2050,N_175);
and U9324 (N_9324,N_184,N_3850);
and U9325 (N_9325,N_680,N_1289);
and U9326 (N_9326,N_2784,N_4793);
nor U9327 (N_9327,N_3690,N_3573);
nand U9328 (N_9328,N_505,N_1375);
nand U9329 (N_9329,N_4158,N_529);
nor U9330 (N_9330,N_4420,N_3441);
and U9331 (N_9331,N_2594,N_44);
and U9332 (N_9332,N_1939,N_1723);
nand U9333 (N_9333,N_3921,N_2762);
nand U9334 (N_9334,N_3655,N_4750);
nor U9335 (N_9335,N_4739,N_4236);
and U9336 (N_9336,N_1758,N_1812);
nand U9337 (N_9337,N_4018,N_3241);
xnor U9338 (N_9338,N_154,N_4181);
or U9339 (N_9339,N_1327,N_3123);
or U9340 (N_9340,N_4558,N_619);
or U9341 (N_9341,N_29,N_862);
nand U9342 (N_9342,N_3654,N_3861);
nand U9343 (N_9343,N_4840,N_3931);
or U9344 (N_9344,N_2974,N_3391);
nor U9345 (N_9345,N_2392,N_2200);
nand U9346 (N_9346,N_2875,N_1648);
nand U9347 (N_9347,N_3188,N_3068);
or U9348 (N_9348,N_1348,N_2703);
or U9349 (N_9349,N_722,N_3269);
and U9350 (N_9350,N_2196,N_3646);
nand U9351 (N_9351,N_848,N_3466);
nand U9352 (N_9352,N_450,N_961);
nor U9353 (N_9353,N_3779,N_4843);
nand U9354 (N_9354,N_1867,N_1884);
and U9355 (N_9355,N_894,N_344);
nand U9356 (N_9356,N_1912,N_4035);
xor U9357 (N_9357,N_4285,N_2599);
and U9358 (N_9358,N_3594,N_758);
and U9359 (N_9359,N_1236,N_2394);
nor U9360 (N_9360,N_1537,N_473);
nor U9361 (N_9361,N_4211,N_1051);
nand U9362 (N_9362,N_1926,N_3077);
or U9363 (N_9363,N_186,N_4794);
nand U9364 (N_9364,N_424,N_2324);
or U9365 (N_9365,N_4244,N_1388);
and U9366 (N_9366,N_3118,N_4925);
or U9367 (N_9367,N_4104,N_4749);
xor U9368 (N_9368,N_1528,N_4977);
nor U9369 (N_9369,N_1392,N_4383);
nor U9370 (N_9370,N_185,N_256);
nor U9371 (N_9371,N_4719,N_397);
nand U9372 (N_9372,N_1473,N_805);
nor U9373 (N_9373,N_4531,N_3892);
nor U9374 (N_9374,N_2530,N_3926);
and U9375 (N_9375,N_985,N_2242);
nand U9376 (N_9376,N_762,N_1469);
nor U9377 (N_9377,N_4631,N_4064);
nand U9378 (N_9378,N_4898,N_2956);
nand U9379 (N_9379,N_1726,N_4751);
nor U9380 (N_9380,N_1319,N_1359);
and U9381 (N_9381,N_3271,N_3837);
nor U9382 (N_9382,N_3294,N_4925);
or U9383 (N_9383,N_4005,N_3949);
and U9384 (N_9384,N_1977,N_193);
nand U9385 (N_9385,N_3775,N_850);
nand U9386 (N_9386,N_3947,N_4788);
nand U9387 (N_9387,N_4275,N_4129);
nor U9388 (N_9388,N_3521,N_4080);
nand U9389 (N_9389,N_2927,N_3648);
or U9390 (N_9390,N_305,N_3155);
and U9391 (N_9391,N_1439,N_2492);
or U9392 (N_9392,N_4566,N_841);
nand U9393 (N_9393,N_4842,N_4514);
nand U9394 (N_9394,N_796,N_3630);
nand U9395 (N_9395,N_202,N_3023);
or U9396 (N_9396,N_1550,N_3341);
and U9397 (N_9397,N_443,N_1774);
xor U9398 (N_9398,N_2065,N_3314);
and U9399 (N_9399,N_457,N_1679);
or U9400 (N_9400,N_2273,N_4654);
or U9401 (N_9401,N_4267,N_2335);
or U9402 (N_9402,N_1955,N_1594);
or U9403 (N_9403,N_935,N_3871);
nor U9404 (N_9404,N_1986,N_1774);
nand U9405 (N_9405,N_2602,N_2529);
nor U9406 (N_9406,N_1550,N_3294);
nand U9407 (N_9407,N_2368,N_652);
or U9408 (N_9408,N_2293,N_1235);
or U9409 (N_9409,N_606,N_1065);
nor U9410 (N_9410,N_554,N_704);
nor U9411 (N_9411,N_2291,N_202);
nor U9412 (N_9412,N_1175,N_1143);
xor U9413 (N_9413,N_278,N_3377);
or U9414 (N_9414,N_4093,N_626);
nor U9415 (N_9415,N_2910,N_530);
xor U9416 (N_9416,N_3365,N_4539);
and U9417 (N_9417,N_2408,N_268);
nand U9418 (N_9418,N_1608,N_877);
nand U9419 (N_9419,N_1812,N_3770);
nor U9420 (N_9420,N_2771,N_766);
and U9421 (N_9421,N_1676,N_954);
nand U9422 (N_9422,N_2960,N_3278);
xnor U9423 (N_9423,N_665,N_3458);
or U9424 (N_9424,N_3916,N_2024);
nor U9425 (N_9425,N_4303,N_239);
nor U9426 (N_9426,N_941,N_1923);
and U9427 (N_9427,N_3627,N_2116);
xnor U9428 (N_9428,N_1351,N_3787);
or U9429 (N_9429,N_3651,N_379);
nand U9430 (N_9430,N_2951,N_1194);
nand U9431 (N_9431,N_2182,N_306);
nor U9432 (N_9432,N_4696,N_1826);
or U9433 (N_9433,N_33,N_330);
nor U9434 (N_9434,N_3386,N_3692);
or U9435 (N_9435,N_3491,N_1901);
nand U9436 (N_9436,N_1391,N_2285);
nor U9437 (N_9437,N_267,N_649);
nor U9438 (N_9438,N_781,N_2190);
nor U9439 (N_9439,N_1604,N_1593);
and U9440 (N_9440,N_3372,N_3055);
xnor U9441 (N_9441,N_2022,N_3832);
nand U9442 (N_9442,N_4731,N_2224);
and U9443 (N_9443,N_871,N_2528);
or U9444 (N_9444,N_3481,N_4070);
nor U9445 (N_9445,N_168,N_2256);
nand U9446 (N_9446,N_816,N_2851);
and U9447 (N_9447,N_1146,N_1055);
or U9448 (N_9448,N_1617,N_3189);
or U9449 (N_9449,N_4784,N_422);
or U9450 (N_9450,N_1303,N_4152);
and U9451 (N_9451,N_1054,N_4897);
nor U9452 (N_9452,N_1144,N_2012);
nor U9453 (N_9453,N_2246,N_753);
xor U9454 (N_9454,N_3759,N_3711);
nor U9455 (N_9455,N_3327,N_4853);
and U9456 (N_9456,N_606,N_2420);
and U9457 (N_9457,N_758,N_2817);
or U9458 (N_9458,N_3881,N_2596);
and U9459 (N_9459,N_441,N_517);
or U9460 (N_9460,N_4585,N_3162);
nor U9461 (N_9461,N_2668,N_2570);
nor U9462 (N_9462,N_2358,N_1896);
and U9463 (N_9463,N_3875,N_4997);
nor U9464 (N_9464,N_244,N_414);
or U9465 (N_9465,N_2987,N_2035);
nor U9466 (N_9466,N_1808,N_42);
nand U9467 (N_9467,N_4576,N_2297);
and U9468 (N_9468,N_264,N_3724);
and U9469 (N_9469,N_1085,N_4449);
and U9470 (N_9470,N_1380,N_608);
nor U9471 (N_9471,N_304,N_1456);
xor U9472 (N_9472,N_1771,N_1623);
or U9473 (N_9473,N_1721,N_2870);
nor U9474 (N_9474,N_3339,N_387);
or U9475 (N_9475,N_2147,N_4876);
and U9476 (N_9476,N_3144,N_4799);
xnor U9477 (N_9477,N_3011,N_442);
and U9478 (N_9478,N_1243,N_606);
or U9479 (N_9479,N_3422,N_2411);
nand U9480 (N_9480,N_4740,N_1995);
xor U9481 (N_9481,N_3514,N_3175);
nand U9482 (N_9482,N_846,N_4423);
and U9483 (N_9483,N_523,N_851);
nor U9484 (N_9484,N_789,N_2406);
nand U9485 (N_9485,N_68,N_770);
nand U9486 (N_9486,N_3637,N_2435);
and U9487 (N_9487,N_4555,N_164);
or U9488 (N_9488,N_2019,N_4021);
nand U9489 (N_9489,N_3168,N_197);
or U9490 (N_9490,N_2917,N_2938);
or U9491 (N_9491,N_1375,N_198);
and U9492 (N_9492,N_3069,N_4328);
or U9493 (N_9493,N_4001,N_252);
and U9494 (N_9494,N_3398,N_2233);
xnor U9495 (N_9495,N_1798,N_9);
or U9496 (N_9496,N_2575,N_591);
and U9497 (N_9497,N_3228,N_2044);
xor U9498 (N_9498,N_44,N_1805);
and U9499 (N_9499,N_11,N_104);
nand U9500 (N_9500,N_3531,N_1936);
and U9501 (N_9501,N_1633,N_612);
and U9502 (N_9502,N_2596,N_3969);
nand U9503 (N_9503,N_2816,N_2419);
nand U9504 (N_9504,N_3614,N_3263);
nand U9505 (N_9505,N_1402,N_2928);
nand U9506 (N_9506,N_1559,N_1252);
nand U9507 (N_9507,N_188,N_2533);
or U9508 (N_9508,N_79,N_4932);
or U9509 (N_9509,N_2212,N_4757);
and U9510 (N_9510,N_3890,N_3146);
nor U9511 (N_9511,N_806,N_2457);
nand U9512 (N_9512,N_563,N_2908);
or U9513 (N_9513,N_4544,N_2336);
nand U9514 (N_9514,N_606,N_2094);
nor U9515 (N_9515,N_1291,N_4210);
and U9516 (N_9516,N_418,N_1326);
or U9517 (N_9517,N_3511,N_2319);
and U9518 (N_9518,N_4971,N_617);
and U9519 (N_9519,N_4732,N_3265);
or U9520 (N_9520,N_3140,N_2517);
xnor U9521 (N_9521,N_1397,N_2791);
nor U9522 (N_9522,N_3814,N_948);
nor U9523 (N_9523,N_1085,N_4524);
xnor U9524 (N_9524,N_2513,N_4476);
nand U9525 (N_9525,N_3864,N_1147);
nand U9526 (N_9526,N_3913,N_4082);
xor U9527 (N_9527,N_85,N_1941);
and U9528 (N_9528,N_4650,N_3587);
and U9529 (N_9529,N_50,N_4518);
nor U9530 (N_9530,N_1893,N_4888);
nand U9531 (N_9531,N_3432,N_4543);
or U9532 (N_9532,N_4888,N_1315);
or U9533 (N_9533,N_4466,N_3402);
nor U9534 (N_9534,N_4499,N_2091);
or U9535 (N_9535,N_1732,N_2613);
xor U9536 (N_9536,N_2668,N_2387);
or U9537 (N_9537,N_59,N_3905);
nand U9538 (N_9538,N_4175,N_143);
nor U9539 (N_9539,N_1186,N_3216);
nand U9540 (N_9540,N_420,N_4193);
nor U9541 (N_9541,N_4422,N_781);
nand U9542 (N_9542,N_2431,N_1992);
nand U9543 (N_9543,N_2657,N_4367);
nor U9544 (N_9544,N_4583,N_1281);
nand U9545 (N_9545,N_2442,N_1539);
nor U9546 (N_9546,N_1925,N_4805);
or U9547 (N_9547,N_3061,N_650);
nand U9548 (N_9548,N_770,N_2890);
nor U9549 (N_9549,N_2919,N_473);
nor U9550 (N_9550,N_1038,N_4578);
nand U9551 (N_9551,N_1278,N_2205);
and U9552 (N_9552,N_3043,N_3908);
or U9553 (N_9553,N_3557,N_4240);
xnor U9554 (N_9554,N_711,N_508);
nor U9555 (N_9555,N_2264,N_2504);
and U9556 (N_9556,N_1681,N_1617);
nand U9557 (N_9557,N_2607,N_4601);
and U9558 (N_9558,N_2404,N_4117);
nor U9559 (N_9559,N_3992,N_2575);
xnor U9560 (N_9560,N_526,N_2085);
and U9561 (N_9561,N_3839,N_2474);
nand U9562 (N_9562,N_4718,N_50);
xor U9563 (N_9563,N_151,N_2395);
or U9564 (N_9564,N_3700,N_4711);
or U9565 (N_9565,N_527,N_3269);
or U9566 (N_9566,N_4310,N_1622);
and U9567 (N_9567,N_594,N_1710);
xnor U9568 (N_9568,N_770,N_2300);
or U9569 (N_9569,N_1687,N_2493);
nand U9570 (N_9570,N_4603,N_3848);
nand U9571 (N_9571,N_3918,N_1449);
or U9572 (N_9572,N_4599,N_3970);
xor U9573 (N_9573,N_4389,N_2326);
nand U9574 (N_9574,N_2932,N_2651);
or U9575 (N_9575,N_4188,N_338);
nand U9576 (N_9576,N_165,N_2174);
nand U9577 (N_9577,N_901,N_449);
nor U9578 (N_9578,N_533,N_4289);
and U9579 (N_9579,N_4176,N_4159);
and U9580 (N_9580,N_2402,N_4759);
nor U9581 (N_9581,N_4076,N_3448);
nand U9582 (N_9582,N_1556,N_360);
and U9583 (N_9583,N_4457,N_238);
nand U9584 (N_9584,N_1554,N_532);
nor U9585 (N_9585,N_2280,N_3309);
or U9586 (N_9586,N_3934,N_4387);
and U9587 (N_9587,N_1796,N_473);
or U9588 (N_9588,N_3654,N_2022);
nand U9589 (N_9589,N_2760,N_2059);
nor U9590 (N_9590,N_2961,N_1379);
nor U9591 (N_9591,N_3237,N_1725);
and U9592 (N_9592,N_4824,N_3239);
or U9593 (N_9593,N_1190,N_400);
and U9594 (N_9594,N_43,N_68);
nand U9595 (N_9595,N_944,N_4607);
and U9596 (N_9596,N_4345,N_4589);
nand U9597 (N_9597,N_1362,N_2295);
nor U9598 (N_9598,N_3271,N_3637);
nor U9599 (N_9599,N_2125,N_40);
or U9600 (N_9600,N_3238,N_586);
nor U9601 (N_9601,N_3537,N_4843);
and U9602 (N_9602,N_695,N_532);
nor U9603 (N_9603,N_3294,N_830);
nand U9604 (N_9604,N_4431,N_2101);
or U9605 (N_9605,N_813,N_2066);
nor U9606 (N_9606,N_1772,N_243);
xnor U9607 (N_9607,N_427,N_4690);
nor U9608 (N_9608,N_1157,N_2609);
nor U9609 (N_9609,N_4063,N_3959);
nor U9610 (N_9610,N_1802,N_3036);
and U9611 (N_9611,N_577,N_1940);
xnor U9612 (N_9612,N_4100,N_4988);
and U9613 (N_9613,N_2809,N_4716);
nor U9614 (N_9614,N_2251,N_561);
and U9615 (N_9615,N_1128,N_2408);
or U9616 (N_9616,N_570,N_4068);
or U9617 (N_9617,N_2709,N_4325);
nor U9618 (N_9618,N_3730,N_4360);
nand U9619 (N_9619,N_2326,N_1687);
nor U9620 (N_9620,N_3005,N_2078);
nor U9621 (N_9621,N_3077,N_2340);
xnor U9622 (N_9622,N_4342,N_1863);
nand U9623 (N_9623,N_2951,N_1828);
and U9624 (N_9624,N_2828,N_829);
xnor U9625 (N_9625,N_73,N_3433);
and U9626 (N_9626,N_3815,N_4350);
and U9627 (N_9627,N_1058,N_1570);
or U9628 (N_9628,N_3662,N_4115);
nand U9629 (N_9629,N_61,N_365);
nor U9630 (N_9630,N_3995,N_4449);
and U9631 (N_9631,N_2831,N_113);
and U9632 (N_9632,N_2013,N_4854);
and U9633 (N_9633,N_2698,N_603);
and U9634 (N_9634,N_3304,N_20);
or U9635 (N_9635,N_825,N_3954);
and U9636 (N_9636,N_1874,N_4963);
nand U9637 (N_9637,N_4886,N_2742);
or U9638 (N_9638,N_1388,N_1567);
or U9639 (N_9639,N_3588,N_3308);
nor U9640 (N_9640,N_4999,N_2966);
xor U9641 (N_9641,N_3247,N_1436);
xor U9642 (N_9642,N_1791,N_3764);
xnor U9643 (N_9643,N_1581,N_1500);
or U9644 (N_9644,N_3940,N_997);
nor U9645 (N_9645,N_1355,N_2927);
xor U9646 (N_9646,N_3722,N_2840);
nand U9647 (N_9647,N_987,N_1483);
or U9648 (N_9648,N_1583,N_206);
nand U9649 (N_9649,N_2174,N_3390);
nor U9650 (N_9650,N_1585,N_3225);
xnor U9651 (N_9651,N_1261,N_1416);
or U9652 (N_9652,N_4455,N_504);
nor U9653 (N_9653,N_1481,N_1800);
and U9654 (N_9654,N_1093,N_2170);
xor U9655 (N_9655,N_754,N_1703);
xnor U9656 (N_9656,N_1470,N_238);
and U9657 (N_9657,N_1807,N_3927);
nand U9658 (N_9658,N_3033,N_2885);
or U9659 (N_9659,N_1679,N_4571);
and U9660 (N_9660,N_974,N_963);
xor U9661 (N_9661,N_4455,N_3534);
xnor U9662 (N_9662,N_4433,N_751);
nand U9663 (N_9663,N_4188,N_1749);
nor U9664 (N_9664,N_711,N_741);
nand U9665 (N_9665,N_3534,N_1292);
or U9666 (N_9666,N_2911,N_4205);
or U9667 (N_9667,N_4940,N_1095);
or U9668 (N_9668,N_2476,N_4289);
and U9669 (N_9669,N_1688,N_4529);
or U9670 (N_9670,N_1779,N_1200);
and U9671 (N_9671,N_1288,N_1135);
xnor U9672 (N_9672,N_2423,N_1134);
and U9673 (N_9673,N_3482,N_2449);
nor U9674 (N_9674,N_213,N_4265);
and U9675 (N_9675,N_483,N_1666);
nand U9676 (N_9676,N_679,N_2152);
nor U9677 (N_9677,N_2180,N_3449);
xor U9678 (N_9678,N_1404,N_3536);
and U9679 (N_9679,N_2739,N_4953);
nor U9680 (N_9680,N_4022,N_2799);
or U9681 (N_9681,N_4881,N_4783);
nor U9682 (N_9682,N_3829,N_395);
xor U9683 (N_9683,N_4329,N_2448);
nand U9684 (N_9684,N_1457,N_1846);
nor U9685 (N_9685,N_1757,N_4131);
or U9686 (N_9686,N_4115,N_1579);
and U9687 (N_9687,N_4363,N_334);
and U9688 (N_9688,N_1950,N_662);
and U9689 (N_9689,N_1950,N_2700);
xnor U9690 (N_9690,N_4277,N_1245);
xnor U9691 (N_9691,N_391,N_323);
xnor U9692 (N_9692,N_3517,N_3057);
nor U9693 (N_9693,N_1856,N_391);
and U9694 (N_9694,N_228,N_210);
or U9695 (N_9695,N_3108,N_4388);
nor U9696 (N_9696,N_2616,N_3110);
and U9697 (N_9697,N_4755,N_2517);
nand U9698 (N_9698,N_4265,N_3466);
nor U9699 (N_9699,N_3289,N_2072);
nor U9700 (N_9700,N_3644,N_1887);
nand U9701 (N_9701,N_1390,N_4827);
and U9702 (N_9702,N_3324,N_2158);
nor U9703 (N_9703,N_2282,N_4932);
or U9704 (N_9704,N_4376,N_4327);
nand U9705 (N_9705,N_495,N_864);
nand U9706 (N_9706,N_2858,N_1959);
nand U9707 (N_9707,N_4017,N_2242);
and U9708 (N_9708,N_1560,N_1586);
and U9709 (N_9709,N_1046,N_800);
or U9710 (N_9710,N_3276,N_1444);
nor U9711 (N_9711,N_2513,N_4766);
nand U9712 (N_9712,N_355,N_367);
or U9713 (N_9713,N_182,N_746);
nor U9714 (N_9714,N_3581,N_4633);
and U9715 (N_9715,N_4779,N_2948);
nor U9716 (N_9716,N_3192,N_2240);
or U9717 (N_9717,N_1174,N_2377);
nor U9718 (N_9718,N_4396,N_4884);
or U9719 (N_9719,N_3025,N_2394);
nand U9720 (N_9720,N_3646,N_2089);
or U9721 (N_9721,N_2727,N_3113);
nand U9722 (N_9722,N_3868,N_2533);
and U9723 (N_9723,N_371,N_4637);
or U9724 (N_9724,N_2769,N_4526);
and U9725 (N_9725,N_3053,N_3906);
or U9726 (N_9726,N_2317,N_1408);
and U9727 (N_9727,N_2816,N_3517);
nand U9728 (N_9728,N_3767,N_2140);
or U9729 (N_9729,N_2114,N_4616);
nor U9730 (N_9730,N_1088,N_3816);
nor U9731 (N_9731,N_1702,N_3713);
nor U9732 (N_9732,N_4095,N_2301);
xnor U9733 (N_9733,N_329,N_2865);
and U9734 (N_9734,N_3023,N_4879);
xor U9735 (N_9735,N_2171,N_3543);
and U9736 (N_9736,N_4079,N_1879);
or U9737 (N_9737,N_1793,N_1497);
or U9738 (N_9738,N_4866,N_3228);
and U9739 (N_9739,N_3830,N_4942);
or U9740 (N_9740,N_4353,N_2637);
nor U9741 (N_9741,N_1446,N_4885);
and U9742 (N_9742,N_2111,N_748);
nor U9743 (N_9743,N_1841,N_195);
nand U9744 (N_9744,N_654,N_2681);
or U9745 (N_9745,N_4664,N_1028);
nand U9746 (N_9746,N_779,N_3290);
nand U9747 (N_9747,N_180,N_2517);
or U9748 (N_9748,N_1906,N_3847);
and U9749 (N_9749,N_3333,N_465);
and U9750 (N_9750,N_4564,N_3140);
nor U9751 (N_9751,N_1942,N_1171);
nand U9752 (N_9752,N_3527,N_191);
and U9753 (N_9753,N_2966,N_547);
and U9754 (N_9754,N_3108,N_589);
or U9755 (N_9755,N_3243,N_230);
nand U9756 (N_9756,N_3719,N_4210);
or U9757 (N_9757,N_755,N_4183);
xnor U9758 (N_9758,N_1226,N_2196);
and U9759 (N_9759,N_1863,N_1759);
nand U9760 (N_9760,N_3712,N_3106);
or U9761 (N_9761,N_3351,N_2985);
nor U9762 (N_9762,N_2687,N_68);
nand U9763 (N_9763,N_1571,N_2306);
xnor U9764 (N_9764,N_2466,N_605);
nor U9765 (N_9765,N_4223,N_688);
nor U9766 (N_9766,N_84,N_4437);
nand U9767 (N_9767,N_4588,N_4405);
or U9768 (N_9768,N_4784,N_4664);
or U9769 (N_9769,N_2848,N_3094);
nand U9770 (N_9770,N_4724,N_914);
and U9771 (N_9771,N_2143,N_1804);
or U9772 (N_9772,N_3661,N_4040);
nor U9773 (N_9773,N_3239,N_1029);
and U9774 (N_9774,N_2067,N_2305);
and U9775 (N_9775,N_1830,N_972);
and U9776 (N_9776,N_446,N_851);
xor U9777 (N_9777,N_783,N_3913);
nor U9778 (N_9778,N_3481,N_2610);
or U9779 (N_9779,N_2169,N_4462);
nand U9780 (N_9780,N_3272,N_1252);
nor U9781 (N_9781,N_3098,N_734);
and U9782 (N_9782,N_2200,N_210);
nand U9783 (N_9783,N_4210,N_3437);
nor U9784 (N_9784,N_2033,N_1531);
and U9785 (N_9785,N_587,N_4239);
or U9786 (N_9786,N_613,N_3611);
nor U9787 (N_9787,N_1493,N_1734);
nor U9788 (N_9788,N_2777,N_2059);
nand U9789 (N_9789,N_3742,N_2940);
nand U9790 (N_9790,N_277,N_3867);
xnor U9791 (N_9791,N_1767,N_2051);
xnor U9792 (N_9792,N_4140,N_383);
xor U9793 (N_9793,N_4432,N_2256);
and U9794 (N_9794,N_153,N_1889);
nand U9795 (N_9795,N_4481,N_1545);
or U9796 (N_9796,N_3292,N_4198);
nor U9797 (N_9797,N_2571,N_3461);
nor U9798 (N_9798,N_1468,N_41);
nor U9799 (N_9799,N_3923,N_425);
xnor U9800 (N_9800,N_4753,N_1376);
nor U9801 (N_9801,N_1819,N_3798);
nand U9802 (N_9802,N_1530,N_2854);
or U9803 (N_9803,N_2969,N_3229);
nand U9804 (N_9804,N_3984,N_4415);
or U9805 (N_9805,N_3394,N_2204);
nor U9806 (N_9806,N_898,N_4368);
and U9807 (N_9807,N_3807,N_2887);
and U9808 (N_9808,N_2911,N_2181);
and U9809 (N_9809,N_1633,N_4260);
nor U9810 (N_9810,N_2880,N_1553);
or U9811 (N_9811,N_2540,N_2292);
nand U9812 (N_9812,N_2284,N_3777);
and U9813 (N_9813,N_3140,N_4441);
nor U9814 (N_9814,N_2122,N_145);
nand U9815 (N_9815,N_335,N_1036);
and U9816 (N_9816,N_629,N_3173);
or U9817 (N_9817,N_2043,N_3384);
and U9818 (N_9818,N_3524,N_2412);
nor U9819 (N_9819,N_1597,N_3241);
nand U9820 (N_9820,N_2704,N_2625);
or U9821 (N_9821,N_2350,N_1433);
nand U9822 (N_9822,N_1250,N_2341);
and U9823 (N_9823,N_3723,N_4286);
or U9824 (N_9824,N_4075,N_3849);
or U9825 (N_9825,N_2805,N_2882);
nor U9826 (N_9826,N_4878,N_643);
or U9827 (N_9827,N_1671,N_4123);
or U9828 (N_9828,N_1808,N_2852);
nand U9829 (N_9829,N_1020,N_3589);
or U9830 (N_9830,N_3665,N_3438);
nor U9831 (N_9831,N_281,N_3234);
nor U9832 (N_9832,N_2773,N_1464);
nor U9833 (N_9833,N_4124,N_3461);
or U9834 (N_9834,N_2356,N_3966);
nand U9835 (N_9835,N_3051,N_548);
nand U9836 (N_9836,N_3095,N_4775);
xnor U9837 (N_9837,N_3084,N_4006);
nor U9838 (N_9838,N_2239,N_2669);
nand U9839 (N_9839,N_3366,N_2791);
xnor U9840 (N_9840,N_3160,N_416);
nand U9841 (N_9841,N_3680,N_2632);
xor U9842 (N_9842,N_4370,N_4145);
nor U9843 (N_9843,N_3953,N_3264);
nor U9844 (N_9844,N_3134,N_3490);
nand U9845 (N_9845,N_2218,N_1061);
and U9846 (N_9846,N_4313,N_1719);
or U9847 (N_9847,N_4510,N_1414);
and U9848 (N_9848,N_3342,N_1804);
xnor U9849 (N_9849,N_2370,N_216);
nand U9850 (N_9850,N_1433,N_1586);
nand U9851 (N_9851,N_1471,N_4713);
or U9852 (N_9852,N_4507,N_641);
and U9853 (N_9853,N_3631,N_257);
and U9854 (N_9854,N_4518,N_1312);
nor U9855 (N_9855,N_261,N_3249);
nor U9856 (N_9856,N_3706,N_3513);
or U9857 (N_9857,N_2875,N_4691);
and U9858 (N_9858,N_1343,N_1620);
and U9859 (N_9859,N_1713,N_4117);
nor U9860 (N_9860,N_2903,N_1814);
nor U9861 (N_9861,N_4165,N_2955);
nand U9862 (N_9862,N_2050,N_1948);
nor U9863 (N_9863,N_1275,N_3638);
or U9864 (N_9864,N_4592,N_1769);
nor U9865 (N_9865,N_2692,N_4367);
xor U9866 (N_9866,N_1941,N_4817);
and U9867 (N_9867,N_833,N_2931);
nand U9868 (N_9868,N_3721,N_2446);
nor U9869 (N_9869,N_2433,N_3816);
or U9870 (N_9870,N_4292,N_3759);
and U9871 (N_9871,N_1292,N_256);
nor U9872 (N_9872,N_1680,N_4666);
or U9873 (N_9873,N_2821,N_3995);
nand U9874 (N_9874,N_4585,N_695);
nand U9875 (N_9875,N_4403,N_218);
nand U9876 (N_9876,N_3565,N_3980);
and U9877 (N_9877,N_630,N_4226);
nor U9878 (N_9878,N_2268,N_1042);
nand U9879 (N_9879,N_3544,N_1658);
xor U9880 (N_9880,N_2374,N_2529);
or U9881 (N_9881,N_2692,N_1333);
or U9882 (N_9882,N_684,N_3538);
or U9883 (N_9883,N_4455,N_1654);
nand U9884 (N_9884,N_4663,N_1792);
and U9885 (N_9885,N_2541,N_3955);
nor U9886 (N_9886,N_141,N_520);
and U9887 (N_9887,N_2258,N_989);
and U9888 (N_9888,N_770,N_2771);
nand U9889 (N_9889,N_3656,N_2595);
xor U9890 (N_9890,N_1685,N_1457);
or U9891 (N_9891,N_555,N_4085);
nand U9892 (N_9892,N_156,N_3879);
nand U9893 (N_9893,N_455,N_3348);
or U9894 (N_9894,N_2233,N_2534);
nand U9895 (N_9895,N_3030,N_4601);
or U9896 (N_9896,N_471,N_3060);
and U9897 (N_9897,N_336,N_287);
and U9898 (N_9898,N_3557,N_1569);
nor U9899 (N_9899,N_4647,N_3223);
xnor U9900 (N_9900,N_4778,N_3208);
xnor U9901 (N_9901,N_1209,N_1171);
nand U9902 (N_9902,N_1376,N_2221);
nand U9903 (N_9903,N_1715,N_385);
nor U9904 (N_9904,N_1189,N_207);
and U9905 (N_9905,N_2946,N_4882);
nand U9906 (N_9906,N_4614,N_3066);
or U9907 (N_9907,N_3713,N_722);
nand U9908 (N_9908,N_2462,N_237);
nor U9909 (N_9909,N_655,N_4898);
and U9910 (N_9910,N_3708,N_3112);
xor U9911 (N_9911,N_1358,N_3088);
nor U9912 (N_9912,N_1533,N_1347);
or U9913 (N_9913,N_1792,N_936);
xor U9914 (N_9914,N_4395,N_3085);
nand U9915 (N_9915,N_582,N_564);
nand U9916 (N_9916,N_1724,N_2169);
or U9917 (N_9917,N_4254,N_3881);
and U9918 (N_9918,N_3163,N_4235);
and U9919 (N_9919,N_943,N_2806);
or U9920 (N_9920,N_336,N_1176);
nor U9921 (N_9921,N_857,N_4503);
and U9922 (N_9922,N_4855,N_199);
nand U9923 (N_9923,N_231,N_3758);
nand U9924 (N_9924,N_2334,N_2913);
or U9925 (N_9925,N_4742,N_2612);
or U9926 (N_9926,N_110,N_3333);
or U9927 (N_9927,N_4802,N_937);
nor U9928 (N_9928,N_228,N_4432);
nand U9929 (N_9929,N_1691,N_4604);
nand U9930 (N_9930,N_1767,N_1183);
xnor U9931 (N_9931,N_4517,N_3689);
xor U9932 (N_9932,N_2317,N_210);
and U9933 (N_9933,N_3447,N_4958);
and U9934 (N_9934,N_697,N_3656);
or U9935 (N_9935,N_1681,N_1132);
nor U9936 (N_9936,N_1753,N_3876);
and U9937 (N_9937,N_131,N_1154);
nor U9938 (N_9938,N_618,N_541);
nand U9939 (N_9939,N_467,N_4402);
nand U9940 (N_9940,N_4641,N_1480);
nor U9941 (N_9941,N_1223,N_2197);
nand U9942 (N_9942,N_1298,N_3991);
nand U9943 (N_9943,N_496,N_1612);
nor U9944 (N_9944,N_392,N_4890);
xnor U9945 (N_9945,N_4187,N_576);
and U9946 (N_9946,N_3742,N_780);
or U9947 (N_9947,N_3514,N_296);
nor U9948 (N_9948,N_4423,N_3096);
or U9949 (N_9949,N_3750,N_3486);
and U9950 (N_9950,N_154,N_543);
nor U9951 (N_9951,N_195,N_1281);
nor U9952 (N_9952,N_3784,N_208);
nand U9953 (N_9953,N_2506,N_3054);
nor U9954 (N_9954,N_4280,N_2283);
nor U9955 (N_9955,N_464,N_2608);
nand U9956 (N_9956,N_3396,N_4160);
nor U9957 (N_9957,N_4788,N_1615);
or U9958 (N_9958,N_1312,N_1372);
or U9959 (N_9959,N_3436,N_182);
or U9960 (N_9960,N_1743,N_3572);
and U9961 (N_9961,N_2302,N_4789);
and U9962 (N_9962,N_2446,N_529);
and U9963 (N_9963,N_3060,N_693);
and U9964 (N_9964,N_2163,N_4598);
nor U9965 (N_9965,N_2019,N_4971);
xnor U9966 (N_9966,N_489,N_1567);
or U9967 (N_9967,N_4525,N_1482);
nor U9968 (N_9968,N_4817,N_3699);
xnor U9969 (N_9969,N_454,N_570);
xnor U9970 (N_9970,N_3264,N_4750);
or U9971 (N_9971,N_4284,N_1088);
and U9972 (N_9972,N_1562,N_2241);
and U9973 (N_9973,N_4670,N_4811);
and U9974 (N_9974,N_282,N_3991);
and U9975 (N_9975,N_851,N_4831);
nand U9976 (N_9976,N_2033,N_3495);
nand U9977 (N_9977,N_4616,N_3208);
and U9978 (N_9978,N_4687,N_3332);
nor U9979 (N_9979,N_2599,N_1433);
and U9980 (N_9980,N_3811,N_77);
xnor U9981 (N_9981,N_4638,N_2454);
nand U9982 (N_9982,N_936,N_4901);
or U9983 (N_9983,N_813,N_1749);
nor U9984 (N_9984,N_495,N_1771);
or U9985 (N_9985,N_1163,N_4303);
nand U9986 (N_9986,N_485,N_4861);
and U9987 (N_9987,N_2223,N_1082);
or U9988 (N_9988,N_1521,N_391);
nand U9989 (N_9989,N_1131,N_4012);
or U9990 (N_9990,N_4567,N_3471);
xor U9991 (N_9991,N_228,N_3540);
xor U9992 (N_9992,N_4739,N_2906);
or U9993 (N_9993,N_2776,N_1796);
nor U9994 (N_9994,N_2935,N_267);
and U9995 (N_9995,N_1878,N_1508);
nor U9996 (N_9996,N_2773,N_4031);
nand U9997 (N_9997,N_1160,N_1162);
nand U9998 (N_9998,N_1846,N_4839);
nand U9999 (N_9999,N_4247,N_3899);
and U10000 (N_10000,N_5988,N_7931);
or U10001 (N_10001,N_5860,N_7510);
nand U10002 (N_10002,N_9189,N_9891);
nor U10003 (N_10003,N_9581,N_6375);
or U10004 (N_10004,N_8444,N_7649);
nand U10005 (N_10005,N_5947,N_5001);
nor U10006 (N_10006,N_8719,N_6699);
and U10007 (N_10007,N_9706,N_9553);
nor U10008 (N_10008,N_7841,N_8833);
and U10009 (N_10009,N_5191,N_6051);
and U10010 (N_10010,N_5351,N_5362);
nand U10011 (N_10011,N_6752,N_6255);
nand U10012 (N_10012,N_6425,N_5037);
and U10013 (N_10013,N_7724,N_6118);
nand U10014 (N_10014,N_9556,N_8159);
xor U10015 (N_10015,N_8795,N_9000);
nor U10016 (N_10016,N_8506,N_5332);
and U10017 (N_10017,N_7028,N_9435);
nand U10018 (N_10018,N_8805,N_9676);
or U10019 (N_10019,N_7234,N_7680);
xnor U10020 (N_10020,N_7088,N_8151);
xor U10021 (N_10021,N_6065,N_7795);
xor U10022 (N_10022,N_8778,N_9145);
and U10023 (N_10023,N_7302,N_7557);
and U10024 (N_10024,N_6626,N_5182);
or U10025 (N_10025,N_5698,N_5903);
and U10026 (N_10026,N_8145,N_5284);
and U10027 (N_10027,N_5190,N_5591);
and U10028 (N_10028,N_8561,N_5868);
and U10029 (N_10029,N_5401,N_9601);
and U10030 (N_10030,N_9453,N_9052);
or U10031 (N_10031,N_7970,N_6088);
nand U10032 (N_10032,N_5295,N_5376);
xnor U10033 (N_10033,N_8403,N_6237);
nor U10034 (N_10034,N_5747,N_9301);
and U10035 (N_10035,N_6863,N_7683);
nor U10036 (N_10036,N_6976,N_6713);
nor U10037 (N_10037,N_6350,N_7330);
and U10038 (N_10038,N_7732,N_7698);
or U10039 (N_10039,N_9386,N_6321);
nand U10040 (N_10040,N_9436,N_9076);
nand U10041 (N_10041,N_6407,N_8324);
nor U10042 (N_10042,N_7417,N_8238);
nand U10043 (N_10043,N_7639,N_7231);
nor U10044 (N_10044,N_9982,N_9126);
nand U10045 (N_10045,N_7863,N_7191);
xor U10046 (N_10046,N_9294,N_5861);
nand U10047 (N_10047,N_7118,N_5631);
or U10048 (N_10048,N_5467,N_6023);
and U10049 (N_10049,N_7364,N_9127);
or U10050 (N_10050,N_7291,N_8697);
nand U10051 (N_10051,N_8943,N_5677);
nand U10052 (N_10052,N_7225,N_5403);
nand U10053 (N_10053,N_8550,N_7584);
or U10054 (N_10054,N_8015,N_7937);
and U10055 (N_10055,N_7445,N_6226);
xnor U10056 (N_10056,N_9783,N_5466);
nor U10057 (N_10057,N_5349,N_6929);
xnor U10058 (N_10058,N_9230,N_8141);
or U10059 (N_10059,N_5079,N_6074);
nand U10060 (N_10060,N_7611,N_7399);
nand U10061 (N_10061,N_7890,N_6664);
and U10062 (N_10062,N_6563,N_6076);
nor U10063 (N_10063,N_9867,N_5850);
and U10064 (N_10064,N_7507,N_5587);
nor U10065 (N_10065,N_6768,N_6735);
nor U10066 (N_10066,N_6609,N_5487);
nand U10067 (N_10067,N_9139,N_8144);
and U10068 (N_10068,N_8856,N_8659);
nand U10069 (N_10069,N_8094,N_8733);
nor U10070 (N_10070,N_9485,N_8575);
xor U10071 (N_10071,N_7927,N_6759);
nand U10072 (N_10072,N_6603,N_7664);
nor U10073 (N_10073,N_6693,N_7098);
nor U10074 (N_10074,N_5302,N_9447);
or U10075 (N_10075,N_7532,N_7884);
or U10076 (N_10076,N_5086,N_7735);
nor U10077 (N_10077,N_8158,N_5519);
nor U10078 (N_10078,N_5525,N_9961);
nand U10079 (N_10079,N_7423,N_9379);
nand U10080 (N_10080,N_8361,N_9307);
nand U10081 (N_10081,N_8537,N_6339);
or U10082 (N_10082,N_5453,N_6641);
and U10083 (N_10083,N_7027,N_6048);
or U10084 (N_10084,N_8173,N_5489);
or U10085 (N_10085,N_9659,N_9773);
xor U10086 (N_10086,N_8655,N_8801);
xnor U10087 (N_10087,N_7778,N_5815);
or U10088 (N_10088,N_9749,N_5112);
nand U10089 (N_10089,N_9089,N_6689);
nand U10090 (N_10090,N_9158,N_9930);
and U10091 (N_10091,N_7530,N_7121);
or U10092 (N_10092,N_9480,N_6814);
nand U10093 (N_10093,N_6963,N_7934);
nor U10094 (N_10094,N_6148,N_5473);
and U10095 (N_10095,N_7730,N_8237);
and U10096 (N_10096,N_6110,N_7387);
nand U10097 (N_10097,N_7046,N_9980);
or U10098 (N_10098,N_5755,N_5609);
nand U10099 (N_10099,N_6409,N_6960);
and U10100 (N_10100,N_6182,N_5049);
nand U10101 (N_10101,N_8342,N_7908);
nand U10102 (N_10102,N_7564,N_6097);
nor U10103 (N_10103,N_5343,N_6083);
nor U10104 (N_10104,N_7705,N_9279);
nand U10105 (N_10105,N_5347,N_7774);
nand U10106 (N_10106,N_8335,N_6945);
and U10107 (N_10107,N_9907,N_6000);
and U10108 (N_10108,N_8024,N_8551);
nand U10109 (N_10109,N_9310,N_5433);
nand U10110 (N_10110,N_7430,N_8842);
nor U10111 (N_10111,N_9190,N_7701);
nor U10112 (N_10112,N_9092,N_8382);
nand U10113 (N_10113,N_5895,N_8080);
or U10114 (N_10114,N_9639,N_7287);
and U10115 (N_10115,N_5047,N_8200);
nor U10116 (N_10116,N_5278,N_6211);
xnor U10117 (N_10117,N_8855,N_5382);
or U10118 (N_10118,N_8681,N_8534);
and U10119 (N_10119,N_6515,N_6253);
nand U10120 (N_10120,N_5948,N_7961);
xor U10121 (N_10121,N_9734,N_9314);
and U10122 (N_10122,N_8139,N_9586);
nand U10123 (N_10123,N_7853,N_5003);
and U10124 (N_10124,N_9383,N_8826);
nor U10125 (N_10125,N_7099,N_5134);
xnor U10126 (N_10126,N_9454,N_8288);
nand U10127 (N_10127,N_6840,N_6050);
or U10128 (N_10128,N_7630,N_5375);
nand U10129 (N_10129,N_6346,N_7646);
xor U10130 (N_10130,N_7901,N_7294);
and U10131 (N_10131,N_8230,N_5844);
and U10132 (N_10132,N_8973,N_9547);
nor U10133 (N_10133,N_9575,N_8735);
nor U10134 (N_10134,N_8220,N_5304);
nand U10135 (N_10135,N_8884,N_5042);
xnor U10136 (N_10136,N_5230,N_8279);
and U10137 (N_10137,N_5852,N_5331);
or U10138 (N_10138,N_8022,N_8677);
nand U10139 (N_10139,N_5156,N_9959);
nor U10140 (N_10140,N_8194,N_7142);
or U10141 (N_10141,N_7616,N_9585);
and U10142 (N_10142,N_6964,N_8251);
and U10143 (N_10143,N_8385,N_6614);
nor U10144 (N_10144,N_5069,N_5132);
nand U10145 (N_10145,N_7017,N_5618);
nor U10146 (N_10146,N_8766,N_6465);
xor U10147 (N_10147,N_9596,N_9433);
or U10148 (N_10148,N_9122,N_7095);
nor U10149 (N_10149,N_9362,N_6442);
nor U10150 (N_10150,N_7957,N_5380);
and U10151 (N_10151,N_7904,N_9934);
and U10152 (N_10152,N_5701,N_7916);
and U10153 (N_10153,N_9572,N_5252);
nor U10154 (N_10154,N_5143,N_6127);
xnor U10155 (N_10155,N_7561,N_7779);
and U10156 (N_10156,N_8001,N_8223);
nand U10157 (N_10157,N_9239,N_9155);
or U10158 (N_10158,N_8789,N_7137);
or U10159 (N_10159,N_6286,N_7565);
and U10160 (N_10160,N_8713,N_8982);
nand U10161 (N_10161,N_8028,N_6259);
and U10162 (N_10162,N_6128,N_9945);
and U10163 (N_10163,N_5658,N_8295);
or U10164 (N_10164,N_6739,N_7866);
nand U10165 (N_10165,N_7899,N_7501);
and U10166 (N_10166,N_9681,N_7588);
nor U10167 (N_10167,N_6108,N_6970);
nor U10168 (N_10168,N_7110,N_5825);
nand U10169 (N_10169,N_7216,N_7462);
xnor U10170 (N_10170,N_6933,N_7435);
or U10171 (N_10171,N_8396,N_7335);
nand U10172 (N_10172,N_9180,N_6272);
or U10173 (N_10173,N_6293,N_6303);
nor U10174 (N_10174,N_6469,N_9025);
or U10175 (N_10175,N_7247,N_6058);
nand U10176 (N_10176,N_7105,N_6310);
nand U10177 (N_10177,N_5711,N_8176);
nor U10178 (N_10178,N_6135,N_5665);
nand U10179 (N_10179,N_5002,N_9367);
and U10180 (N_10180,N_6763,N_5247);
xor U10181 (N_10181,N_8377,N_6341);
and U10182 (N_10182,N_8228,N_9120);
nand U10183 (N_10183,N_9428,N_6969);
and U10184 (N_10184,N_9763,N_8800);
nand U10185 (N_10185,N_5961,N_6480);
and U10186 (N_10186,N_7875,N_7062);
nand U10187 (N_10187,N_8863,N_7472);
or U10188 (N_10188,N_6112,N_6142);
or U10189 (N_10189,N_8702,N_8014);
nand U10190 (N_10190,N_9444,N_9911);
xor U10191 (N_10191,N_8399,N_6646);
and U10192 (N_10192,N_8480,N_8057);
and U10193 (N_10193,N_7114,N_6500);
and U10194 (N_10194,N_9072,N_6367);
or U10195 (N_10195,N_5041,N_9932);
nand U10196 (N_10196,N_5790,N_9516);
nor U10197 (N_10197,N_6477,N_5785);
nand U10198 (N_10198,N_6361,N_9908);
nor U10199 (N_10199,N_9873,N_7091);
or U10200 (N_10200,N_5862,N_7032);
nand U10201 (N_10201,N_9974,N_6443);
and U10202 (N_10202,N_5651,N_6610);
nand U10203 (N_10203,N_7535,N_7080);
and U10204 (N_10204,N_5240,N_5583);
or U10205 (N_10205,N_6144,N_5006);
or U10206 (N_10206,N_7877,N_7828);
and U10207 (N_10207,N_5779,N_8454);
or U10208 (N_10208,N_5219,N_7835);
and U10209 (N_10209,N_8972,N_9758);
and U10210 (N_10210,N_8054,N_5067);
and U10211 (N_10211,N_6206,N_5611);
nor U10212 (N_10212,N_5938,N_5022);
nor U10213 (N_10213,N_6014,N_5916);
nand U10214 (N_10214,N_5661,N_6439);
and U10215 (N_10215,N_7684,N_9097);
nand U10216 (N_10216,N_9549,N_6714);
nor U10217 (N_10217,N_7892,N_5404);
and U10218 (N_10218,N_9465,N_7311);
or U10219 (N_10219,N_9309,N_7550);
nor U10220 (N_10220,N_7458,N_8665);
xor U10221 (N_10221,N_9935,N_6604);
and U10222 (N_10222,N_8513,N_8021);
nand U10223 (N_10223,N_6619,N_7883);
and U10224 (N_10224,N_8264,N_8287);
nor U10225 (N_10225,N_7713,N_6851);
nand U10226 (N_10226,N_6354,N_5432);
nand U10227 (N_10227,N_9674,N_7181);
and U10228 (N_10228,N_9537,N_7796);
nand U10229 (N_10229,N_7051,N_8065);
nor U10230 (N_10230,N_5847,N_5570);
or U10231 (N_10231,N_7707,N_7289);
nor U10232 (N_10232,N_8540,N_6337);
and U10233 (N_10233,N_6841,N_8607);
nand U10234 (N_10234,N_7002,N_6416);
and U10235 (N_10235,N_6218,N_9457);
nand U10236 (N_10236,N_6878,N_5964);
xor U10237 (N_10237,N_5004,N_6165);
nor U10238 (N_10238,N_8286,N_7825);
nor U10239 (N_10239,N_7048,N_6162);
xor U10240 (N_10240,N_6663,N_9999);
nor U10241 (N_10241,N_9916,N_7756);
xnor U10242 (N_10242,N_6791,N_5799);
nand U10243 (N_10243,N_7372,N_7809);
or U10244 (N_10244,N_9176,N_5249);
nand U10245 (N_10245,N_6308,N_5142);
or U10246 (N_10246,N_7852,N_9501);
nor U10247 (N_10247,N_9430,N_8612);
and U10248 (N_10248,N_6141,N_7477);
or U10249 (N_10249,N_7188,N_5336);
nor U10250 (N_10250,N_6181,N_7743);
nor U10251 (N_10251,N_5501,N_5526);
or U10252 (N_10252,N_7856,N_7422);
nor U10253 (N_10253,N_7227,N_6180);
nor U10254 (N_10254,N_8868,N_7545);
nand U10255 (N_10255,N_7769,N_6157);
and U10256 (N_10256,N_9303,N_8323);
or U10257 (N_10257,N_5930,N_8351);
nand U10258 (N_10258,N_8373,N_6015);
and U10259 (N_10259,N_7751,N_6616);
nand U10260 (N_10260,N_8572,N_7156);
xnor U10261 (N_10261,N_8860,N_5664);
or U10262 (N_10262,N_8661,N_6309);
and U10263 (N_10263,N_5911,N_5700);
nand U10264 (N_10264,N_7541,N_5605);
or U10265 (N_10265,N_6622,N_8316);
nand U10266 (N_10266,N_6234,N_6612);
nand U10267 (N_10267,N_8913,N_7251);
and U10268 (N_10268,N_7327,N_5321);
nor U10269 (N_10269,N_6795,N_5722);
nor U10270 (N_10270,N_5090,N_7714);
nor U10271 (N_10271,N_6456,N_8168);
and U10272 (N_10272,N_6244,N_5222);
xnor U10273 (N_10273,N_8031,N_6736);
nor U10274 (N_10274,N_5133,N_7633);
nand U10275 (N_10275,N_8870,N_9166);
nor U10276 (N_10276,N_6574,N_8343);
nand U10277 (N_10277,N_7393,N_8588);
nor U10278 (N_10278,N_9746,N_5293);
xor U10279 (N_10279,N_6230,N_8050);
nor U10280 (N_10280,N_9712,N_9020);
and U10281 (N_10281,N_9250,N_8005);
nand U10282 (N_10282,N_8664,N_8099);
and U10283 (N_10283,N_8011,N_7911);
or U10284 (N_10284,N_9757,N_5276);
xor U10285 (N_10285,N_8874,N_7447);
nand U10286 (N_10286,N_6915,N_5465);
and U10287 (N_10287,N_8197,N_5460);
or U10288 (N_10288,N_5091,N_9210);
nor U10289 (N_10289,N_7451,N_7233);
nor U10290 (N_10290,N_7093,N_8346);
and U10291 (N_10291,N_5866,N_5810);
or U10292 (N_10292,N_9918,N_8755);
nand U10293 (N_10293,N_9896,N_8147);
nand U10294 (N_10294,N_8381,N_8522);
xnor U10295 (N_10295,N_9741,N_5491);
nor U10296 (N_10296,N_6860,N_5007);
nand U10297 (N_10297,N_5084,N_9743);
or U10298 (N_10298,N_7413,N_8265);
or U10299 (N_10299,N_6815,N_8420);
nand U10300 (N_10300,N_6401,N_8306);
nor U10301 (N_10301,N_9762,N_5474);
or U10302 (N_10302,N_8450,N_6973);
nor U10303 (N_10303,N_7845,N_6966);
nor U10304 (N_10304,N_5572,N_8921);
xnor U10305 (N_10305,N_7305,N_9081);
or U10306 (N_10306,N_8280,N_9850);
nand U10307 (N_10307,N_6913,N_5288);
nand U10308 (N_10308,N_9288,N_7326);
and U10309 (N_10309,N_6314,N_9859);
nand U10310 (N_10310,N_6468,N_6712);
nor U10311 (N_10311,N_7461,N_9002);
or U10312 (N_10312,N_9728,N_9666);
nand U10313 (N_10313,N_9701,N_5741);
or U10314 (N_10314,N_8552,N_7591);
nand U10315 (N_10315,N_8658,N_8797);
nor U10316 (N_10316,N_9869,N_5103);
and U10317 (N_10317,N_9616,N_5652);
and U10318 (N_10318,N_5914,N_8148);
xnor U10319 (N_10319,N_7404,N_8625);
nor U10320 (N_10320,N_9544,N_5859);
nor U10321 (N_10321,N_9730,N_7590);
nand U10322 (N_10322,N_5193,N_8121);
or U10323 (N_10323,N_6734,N_8850);
nand U10324 (N_10324,N_6508,N_7479);
nor U10325 (N_10325,N_6613,N_8662);
and U10326 (N_10326,N_6555,N_6406);
or U10327 (N_10327,N_7199,N_7960);
xnor U10328 (N_10328,N_9012,N_8394);
or U10329 (N_10329,N_6249,N_7349);
nand U10330 (N_10330,N_8566,N_6971);
xnor U10331 (N_10331,N_9231,N_5726);
nand U10332 (N_10332,N_9017,N_9764);
or U10333 (N_10333,N_8689,N_6078);
nor U10334 (N_10334,N_5452,N_7256);
and U10335 (N_10335,N_5176,N_6570);
or U10336 (N_10336,N_6880,N_9446);
nor U10337 (N_10337,N_9868,N_9084);
nor U10338 (N_10338,N_8901,N_6844);
nand U10339 (N_10339,N_7965,N_8362);
and U10340 (N_10340,N_9156,N_7694);
or U10341 (N_10341,N_8811,N_7949);
or U10342 (N_10342,N_7159,N_7872);
and U10343 (N_10343,N_9577,N_9904);
or U10344 (N_10344,N_9320,N_5280);
nand U10345 (N_10345,N_9490,N_5910);
and U10346 (N_10346,N_8613,N_9341);
or U10347 (N_10347,N_8975,N_5115);
or U10348 (N_10348,N_6022,N_9654);
nor U10349 (N_10349,N_9579,N_7755);
xor U10350 (N_10350,N_6411,N_5532);
or U10351 (N_10351,N_6030,N_9455);
or U10352 (N_10352,N_6886,N_6576);
or U10353 (N_10353,N_9500,N_5077);
nor U10354 (N_10354,N_5034,N_9543);
and U10355 (N_10355,N_6273,N_7147);
nor U10356 (N_10356,N_9766,N_9075);
and U10357 (N_10357,N_6849,N_7448);
nand U10358 (N_10358,N_9829,N_8933);
or U10359 (N_10359,N_5628,N_8196);
and U10360 (N_10360,N_7351,N_7165);
nor U10361 (N_10361,N_9368,N_7946);
xnor U10362 (N_10362,N_5326,N_9791);
nand U10363 (N_10363,N_7084,N_5013);
nand U10364 (N_10364,N_6615,N_6997);
and U10365 (N_10365,N_8807,N_8949);
nand U10366 (N_10366,N_7208,N_7651);
nor U10367 (N_10367,N_9302,N_5148);
or U10368 (N_10368,N_9021,N_7983);
xnor U10369 (N_10369,N_7466,N_5420);
xnor U10370 (N_10370,N_7858,N_5345);
nor U10371 (N_10371,N_5913,N_7782);
nor U10372 (N_10372,N_7534,N_9315);
nor U10373 (N_10373,N_6605,N_7553);
and U10374 (N_10374,N_7258,N_7166);
nand U10375 (N_10375,N_8268,N_8932);
nor U10376 (N_10376,N_6084,N_6954);
xnor U10377 (N_10377,N_8471,N_9078);
nand U10378 (N_10378,N_5337,N_7500);
and U10379 (N_10379,N_8744,N_5738);
nor U10380 (N_10380,N_9761,N_8181);
or U10381 (N_10381,N_7986,N_8847);
nor U10382 (N_10382,N_8649,N_8259);
or U10383 (N_10383,N_9469,N_8441);
and U10384 (N_10384,N_6787,N_8869);
and U10385 (N_10385,N_6214,N_9598);
and U10386 (N_10386,N_6530,N_5752);
and U10387 (N_10387,N_9718,N_6430);
and U10388 (N_10388,N_6398,N_5399);
nor U10389 (N_10389,N_8329,N_8986);
nor U10390 (N_10390,N_7797,N_9562);
nor U10391 (N_10391,N_8963,N_5596);
nand U10392 (N_10392,N_5025,N_9173);
and U10393 (N_10393,N_5997,N_5610);
nand U10394 (N_10394,N_7280,N_6898);
or U10395 (N_10395,N_5707,N_9476);
xnor U10396 (N_10396,N_5068,N_9193);
or U10397 (N_10397,N_8871,N_7855);
nand U10398 (N_10398,N_9318,N_8563);
nor U10399 (N_10399,N_9118,N_8055);
nand U10400 (N_10400,N_9160,N_5482);
and U10401 (N_10401,N_7265,N_6326);
and U10402 (N_10402,N_6043,N_7576);
and U10403 (N_10403,N_5621,N_5975);
nand U10404 (N_10404,N_9576,N_8872);
nand U10405 (N_10405,N_9838,N_6564);
and U10406 (N_10406,N_9280,N_9382);
nor U10407 (N_10407,N_5392,N_6947);
and U10408 (N_10408,N_6085,N_8107);
nand U10409 (N_10409,N_5051,N_9846);
nor U10410 (N_10410,N_8020,N_7001);
and U10411 (N_10411,N_7641,N_8352);
or U10412 (N_10412,N_6634,N_8751);
xor U10413 (N_10413,N_5490,N_9287);
or U10414 (N_10414,N_5987,N_9834);
or U10415 (N_10415,N_9881,N_6396);
and U10416 (N_10416,N_9950,N_8971);
or U10417 (N_10417,N_9074,N_6593);
xnor U10418 (N_10418,N_6119,N_7711);
nor U10419 (N_10419,N_7094,N_7631);
nand U10420 (N_10420,N_8939,N_5286);
and U10421 (N_10421,N_6818,N_5232);
nor U10422 (N_10422,N_7090,N_6392);
xnor U10423 (N_10423,N_9107,N_7921);
or U10424 (N_10424,N_9936,N_6202);
xnor U10425 (N_10425,N_9512,N_8070);
xnor U10426 (N_10426,N_7082,N_9413);
xnor U10427 (N_10427,N_6645,N_8447);
nor U10428 (N_10428,N_5437,N_5147);
xor U10429 (N_10429,N_6064,N_6158);
nor U10430 (N_10430,N_5704,N_5434);
nor U10431 (N_10431,N_7948,N_7804);
nor U10432 (N_10432,N_5687,N_9731);
nor U10433 (N_10433,N_5499,N_8473);
nand U10434 (N_10434,N_7967,N_8698);
or U10435 (N_10435,N_7681,N_9487);
nand U10436 (N_10436,N_9886,N_9550);
or U10437 (N_10437,N_5902,N_7108);
nand U10438 (N_10438,N_6283,N_7973);
and U10439 (N_10439,N_5165,N_8046);
nand U10440 (N_10440,N_7475,N_5045);
xnor U10441 (N_10441,N_9608,N_8296);
nor U10442 (N_10442,N_6212,N_6934);
or U10443 (N_10443,N_8559,N_9632);
and U10444 (N_10444,N_7169,N_8711);
nor U10445 (N_10445,N_6654,N_5909);
nand U10446 (N_10446,N_7982,N_5679);
or U10447 (N_10447,N_7932,N_9135);
nor U10448 (N_10448,N_6728,N_9340);
or U10449 (N_10449,N_8814,N_5052);
nand U10450 (N_10450,N_7602,N_5794);
or U10451 (N_10451,N_5188,N_6059);
or U10452 (N_10452,N_9124,N_8045);
nand U10453 (N_10453,N_5019,N_6952);
and U10454 (N_10454,N_9528,N_9778);
nand U10455 (N_10455,N_5248,N_8684);
or U10456 (N_10456,N_5443,N_7918);
nand U10457 (N_10457,N_5297,N_6608);
and U10458 (N_10458,N_5877,N_8954);
or U10459 (N_10459,N_9635,N_6792);
nor U10460 (N_10460,N_9634,N_9324);
nor U10461 (N_10461,N_7253,N_9806);
nand U10462 (N_10462,N_5942,N_7329);
nand U10463 (N_10463,N_8166,N_6424);
nor U10464 (N_10464,N_9004,N_6513);
xnor U10465 (N_10465,N_5598,N_8812);
or U10466 (N_10466,N_7943,N_6669);
and U10467 (N_10467,N_5926,N_6385);
or U10468 (N_10468,N_5130,N_7994);
or U10469 (N_10469,N_8034,N_9989);
nor U10470 (N_10470,N_8904,N_9964);
nand U10471 (N_10471,N_5509,N_5279);
or U10472 (N_10472,N_6154,N_7800);
nor U10473 (N_10473,N_5363,N_5372);
nor U10474 (N_10474,N_8968,N_7385);
nand U10475 (N_10475,N_8603,N_5254);
nor U10476 (N_10476,N_7146,N_6188);
and U10477 (N_10477,N_8648,N_6368);
and U10478 (N_10478,N_6575,N_7211);
nor U10479 (N_10479,N_5770,N_6276);
xnor U10480 (N_10480,N_8978,N_7220);
nor U10481 (N_10481,N_9364,N_9938);
or U10482 (N_10482,N_8400,N_5105);
xnor U10483 (N_10483,N_7650,N_9187);
and U10484 (N_10484,N_9841,N_6884);
or U10485 (N_10485,N_8359,N_9931);
nand U10486 (N_10486,N_6107,N_6100);
nor U10487 (N_10487,N_6070,N_8602);
or U10488 (N_10488,N_5692,N_8995);
nand U10489 (N_10489,N_8866,N_8452);
or U10490 (N_10490,N_5873,N_7636);
and U10491 (N_10491,N_5114,N_8113);
xnor U10492 (N_10492,N_5348,N_6241);
nor U10493 (N_10493,N_8327,N_7594);
or U10494 (N_10494,N_6010,N_6675);
nand U10495 (N_10495,N_9801,N_7944);
or U10496 (N_10496,N_5344,N_5080);
and U10497 (N_10497,N_5455,N_6149);
nor U10498 (N_10498,N_7881,N_9401);
or U10499 (N_10499,N_7533,N_7629);
and U10500 (N_10500,N_7012,N_5458);
xnor U10501 (N_10501,N_5070,N_5020);
nand U10502 (N_10502,N_7910,N_5875);
nor U10503 (N_10503,N_7008,N_5361);
nand U10504 (N_10504,N_7543,N_5093);
and U10505 (N_10505,N_8774,N_5542);
nand U10506 (N_10506,N_9702,N_6129);
or U10507 (N_10507,N_9726,N_6926);
nand U10508 (N_10508,N_9745,N_7940);
nor U10509 (N_10509,N_7540,N_5980);
nor U10510 (N_10510,N_9880,N_6071);
or U10511 (N_10511,N_5179,N_7242);
nand U10512 (N_10512,N_8406,N_9966);
and U10513 (N_10513,N_8409,N_8301);
and U10514 (N_10514,N_9445,N_9864);
nand U10515 (N_10515,N_9810,N_8297);
xor U10516 (N_10516,N_7959,N_6986);
nor U10517 (N_10517,N_8078,N_9857);
xor U10518 (N_10518,N_5116,N_8970);
nor U10519 (N_10519,N_5921,N_7504);
xor U10520 (N_10520,N_9957,N_8348);
xnor U10521 (N_10521,N_7695,N_5146);
nand U10522 (N_10522,N_7366,N_9797);
nor U10523 (N_10523,N_6873,N_9399);
nand U10524 (N_10524,N_9612,N_5874);
or U10525 (N_10525,N_8790,N_5480);
and U10526 (N_10526,N_9613,N_8077);
nor U10527 (N_10527,N_9767,N_8535);
nor U10528 (N_10528,N_5322,N_8114);
and U10529 (N_10529,N_5220,N_6967);
and U10530 (N_10530,N_9233,N_9607);
and U10531 (N_10531,N_9879,N_6243);
nand U10532 (N_10532,N_7509,N_9359);
nand U10533 (N_10533,N_7026,N_6270);
nor U10534 (N_10534,N_8467,N_8300);
xnor U10535 (N_10535,N_9019,N_6994);
nand U10536 (N_10536,N_5205,N_9722);
and U10537 (N_10537,N_5060,N_7131);
xnor U10538 (N_10538,N_8235,N_8333);
nand U10539 (N_10539,N_7862,N_8977);
nor U10540 (N_10540,N_8752,N_9924);
and U10541 (N_10541,N_9069,N_8516);
nor U10542 (N_10542,N_9776,N_8341);
and U10543 (N_10543,N_6105,N_5567);
xnor U10544 (N_10544,N_7260,N_5026);
or U10545 (N_10545,N_8309,N_6855);
nand U10546 (N_10546,N_7930,N_9686);
xnor U10547 (N_10547,N_7757,N_5816);
xor U10548 (N_10548,N_6049,N_6598);
nor U10549 (N_10549,N_8782,N_6062);
nor U10550 (N_10550,N_5812,N_7341);
or U10551 (N_10551,N_9129,N_9584);
nor U10552 (N_10552,N_6541,N_8788);
and U10553 (N_10553,N_5035,N_6932);
nand U10554 (N_10554,N_6205,N_5038);
or U10555 (N_10555,N_7784,N_9199);
xnor U10556 (N_10556,N_9725,N_8787);
and U10557 (N_10557,N_9204,N_6447);
nand U10558 (N_10558,N_6327,N_8414);
or U10559 (N_10559,N_9224,N_8209);
nand U10560 (N_10560,N_7975,N_8347);
or U10561 (N_10561,N_6280,N_9708);
and U10562 (N_10562,N_5291,N_8395);
nand U10563 (N_10563,N_6707,N_7136);
and U10564 (N_10564,N_6090,N_8435);
and U10565 (N_10565,N_7492,N_5168);
nor U10566 (N_10566,N_9787,N_8085);
nand U10567 (N_10567,N_5531,N_6377);
and U10568 (N_10568,N_8564,N_7537);
nor U10569 (N_10569,N_5937,N_9484);
or U10570 (N_10570,N_9903,N_6196);
and U10571 (N_10571,N_9086,N_5479);
and U10572 (N_10572,N_7928,N_6706);
and U10573 (N_10573,N_9132,N_7869);
nand U10574 (N_10574,N_8095,N_8412);
and U10575 (N_10575,N_6463,N_5608);
nand U10576 (N_10576,N_6037,N_6004);
and U10577 (N_10577,N_5040,N_9098);
xnor U10578 (N_10578,N_6727,N_8118);
nand U10579 (N_10579,N_7058,N_5588);
xor U10580 (N_10580,N_5686,N_7360);
or U10581 (N_10581,N_6749,N_9472);
and U10582 (N_10582,N_6271,N_8991);
xor U10583 (N_10583,N_5538,N_5659);
nand U10584 (N_10584,N_6872,N_5733);
nand U10585 (N_10585,N_8549,N_9358);
nor U10586 (N_10586,N_6066,N_7328);
or U10587 (N_10587,N_7497,N_6340);
and U10588 (N_10588,N_6708,N_6024);
and U10589 (N_10589,N_5149,N_9704);
xor U10590 (N_10590,N_6720,N_5884);
nand U10591 (N_10591,N_5296,N_9700);
and U10592 (N_10592,N_9717,N_5318);
nand U10593 (N_10593,N_5124,N_8289);
or U10594 (N_10594,N_6784,N_6025);
and U10595 (N_10595,N_5208,N_5811);
nor U10596 (N_10596,N_5207,N_7061);
and U10597 (N_10597,N_8482,N_9848);
nor U10598 (N_10598,N_6091,N_7151);
or U10599 (N_10599,N_5768,N_8569);
nand U10600 (N_10600,N_6171,N_7980);
nand U10601 (N_10601,N_8088,N_6774);
nand U10602 (N_10602,N_5824,N_7463);
nand U10603 (N_10603,N_7392,N_6850);
and U10604 (N_10604,N_5511,N_9511);
nor U10605 (N_10605,N_8270,N_5865);
nor U10606 (N_10606,N_6962,N_6876);
nand U10607 (N_10607,N_8000,N_8715);
xnor U10608 (N_10608,N_5855,N_6016);
and U10609 (N_10609,N_9981,N_7568);
nor U10610 (N_10610,N_6571,N_5268);
and U10611 (N_10611,N_6861,N_5919);
nor U10612 (N_10612,N_9450,N_7459);
or U10613 (N_10613,N_9297,N_7605);
nor U10614 (N_10614,N_9893,N_9317);
nor U10615 (N_10615,N_9010,N_6591);
nand U10616 (N_10616,N_5521,N_7338);
or U10617 (N_10617,N_8241,N_5756);
or U10618 (N_10618,N_5981,N_6155);
and U10619 (N_10619,N_7712,N_7288);
nand U10620 (N_10620,N_8092,N_5275);
nor U10621 (N_10621,N_8438,N_6242);
xor U10622 (N_10622,N_9094,N_6265);
xnor U10623 (N_10623,N_5424,N_8006);
or U10624 (N_10624,N_8858,N_5690);
nand U10625 (N_10625,N_6039,N_9254);
nand U10626 (N_10626,N_6800,N_8928);
or U10627 (N_10627,N_7812,N_9994);
nand U10628 (N_10628,N_5887,N_6569);
nor U10629 (N_10629,N_9887,N_5260);
or U10630 (N_10630,N_8468,N_8802);
nand U10631 (N_10631,N_5929,N_6291);
and U10632 (N_10632,N_9304,N_9710);
nor U10633 (N_10633,N_9526,N_7127);
and U10634 (N_10634,N_6737,N_6067);
and U10635 (N_10635,N_6109,N_8248);
nand U10636 (N_10636,N_9611,N_6560);
and U10637 (N_10637,N_5012,N_6289);
nor U10638 (N_10638,N_9590,N_8526);
or U10639 (N_10639,N_5616,N_8007);
nor U10640 (N_10640,N_9404,N_6238);
nor U10641 (N_10641,N_8650,N_8762);
and U10642 (N_10642,N_8630,N_7212);
or U10643 (N_10643,N_6003,N_5294);
nor U10644 (N_10644,N_6421,N_9240);
nand U10645 (N_10645,N_9571,N_6586);
and U10646 (N_10646,N_9853,N_7968);
or U10647 (N_10647,N_5451,N_9988);
nor U10648 (N_10648,N_8063,N_5739);
xor U10649 (N_10649,N_8272,N_7438);
and U10650 (N_10650,N_8616,N_6438);
and U10651 (N_10651,N_9672,N_6018);
nor U10652 (N_10652,N_7138,N_9014);
nand U10653 (N_10653,N_6903,N_9419);
and U10654 (N_10654,N_5303,N_5640);
nand U10655 (N_10655,N_9733,N_8882);
and U10656 (N_10656,N_6600,N_8753);
nor U10657 (N_10657,N_7054,N_6429);
nor U10658 (N_10658,N_6179,N_7599);
nor U10659 (N_10659,N_8250,N_5500);
nor U10660 (N_10660,N_9604,N_5680);
nand U10661 (N_10661,N_5829,N_9372);
or U10662 (N_10662,N_6801,N_7607);
or U10663 (N_10663,N_5579,N_9407);
nor U10664 (N_10664,N_7271,N_5655);
nand U10665 (N_10665,N_9685,N_9817);
nand U10666 (N_10666,N_7635,N_9154);
or U10667 (N_10667,N_9920,N_8937);
nand U10668 (N_10668,N_7257,N_8221);
or U10669 (N_10669,N_8691,N_6342);
and U10670 (N_10670,N_5406,N_7333);
and U10671 (N_10671,N_6503,N_9330);
nor U10672 (N_10672,N_7988,N_9535);
and U10673 (N_10673,N_5617,N_5830);
nor U10674 (N_10674,N_5101,N_6019);
nand U10675 (N_10675,N_7457,N_5582);
and U10676 (N_10676,N_7867,N_6833);
nor U10677 (N_10677,N_9525,N_5777);
xnor U10678 (N_10678,N_8199,N_9387);
nor U10679 (N_10679,N_7483,N_5261);
xor U10680 (N_10680,N_7401,N_6909);
or U10681 (N_10681,N_9177,N_7966);
nand U10682 (N_10682,N_6949,N_6546);
nand U10683 (N_10683,N_6741,N_6215);
or U10684 (N_10684,N_7525,N_6684);
or U10685 (N_10685,N_5214,N_7347);
xnor U10686 (N_10686,N_6279,N_5078);
or U10687 (N_10687,N_5064,N_6134);
or U10688 (N_10688,N_6836,N_6470);
nand U10689 (N_10689,N_5708,N_7494);
and U10690 (N_10690,N_9420,N_7951);
and U10691 (N_10691,N_6290,N_5057);
and U10692 (N_10692,N_9007,N_7692);
or U10693 (N_10693,N_5120,N_7186);
and U10694 (N_10694,N_5580,N_8459);
nor U10695 (N_10695,N_7659,N_9312);
nand U10696 (N_10696,N_9583,N_9405);
or U10697 (N_10697,N_8101,N_6905);
or U10698 (N_10698,N_6151,N_5387);
nand U10699 (N_10699,N_7130,N_7697);
and U10700 (N_10700,N_8672,N_5059);
or U10701 (N_10701,N_5228,N_8910);
or U10702 (N_10702,N_5414,N_9271);
and U10703 (N_10703,N_6582,N_8922);
or U10704 (N_10704,N_9792,N_6553);
and U10705 (N_10705,N_9357,N_5513);
nor U10706 (N_10706,N_7781,N_7941);
nor U10707 (N_10707,N_9198,N_7601);
or U10708 (N_10708,N_8429,N_7597);
nand U10709 (N_10709,N_7063,N_8003);
and U10710 (N_10710,N_9133,N_6081);
nor U10711 (N_10711,N_8758,N_6123);
or U10712 (N_10712,N_7874,N_8777);
nor U10713 (N_10713,N_9805,N_7361);
and U10714 (N_10714,N_9660,N_7604);
and U10715 (N_10715,N_9281,N_9520);
or U10716 (N_10716,N_8831,N_6137);
nand U10717 (N_10717,N_8740,N_6579);
xor U10718 (N_10718,N_7645,N_5027);
and U10719 (N_10719,N_9178,N_6332);
nor U10720 (N_10720,N_8053,N_8893);
nor U10721 (N_10721,N_8336,N_5181);
and U10722 (N_10722,N_5102,N_7945);
nand U10723 (N_10723,N_7808,N_6435);
nand U10724 (N_10724,N_5312,N_8133);
or U10725 (N_10725,N_5867,N_7558);
nand U10726 (N_10726,N_6902,N_5602);
nand U10727 (N_10727,N_5076,N_8675);
or U10728 (N_10728,N_7298,N_8123);
and U10729 (N_10729,N_5428,N_7811);
nor U10730 (N_10730,N_8531,N_6894);
xnor U10731 (N_10731,N_7240,N_8694);
or U10732 (N_10732,N_8164,N_7603);
nor U10733 (N_10733,N_7015,N_6998);
nand U10734 (N_10734,N_5018,N_6912);
and U10735 (N_10735,N_6153,N_5478);
nor U10736 (N_10736,N_8266,N_6458);
or U10737 (N_10737,N_9148,N_6369);
or U10738 (N_10738,N_8844,N_5368);
or U10739 (N_10739,N_6121,N_9852);
and U10740 (N_10740,N_9416,N_6676);
nor U10741 (N_10741,N_9671,N_9560);
and U10742 (N_10742,N_7065,N_6606);
or U10743 (N_10743,N_5435,N_7820);
or U10744 (N_10744,N_5940,N_8974);
nand U10745 (N_10745,N_7304,N_6979);
nand U10746 (N_10746,N_8463,N_6349);
or U10747 (N_10747,N_5872,N_8062);
nand U10748 (N_10748,N_7572,N_8584);
nor U10749 (N_10749,N_6370,N_7920);
nand U10750 (N_10750,N_7956,N_6681);
nor U10751 (N_10751,N_6315,N_6487);
nor U10752 (N_10752,N_7997,N_5849);
and U10753 (N_10753,N_9971,N_6620);
xnor U10754 (N_10754,N_8518,N_9910);
or U10755 (N_10755,N_7158,N_6034);
and U10756 (N_10756,N_9265,N_7758);
and U10757 (N_10757,N_6195,N_6403);
xnor U10758 (N_10758,N_6665,N_9975);
and U10759 (N_10759,N_5524,N_9862);
and U10760 (N_10760,N_7049,N_9181);
nor U10761 (N_10761,N_6136,N_5954);
and U10762 (N_10762,N_7370,N_8927);
nand U10763 (N_10763,N_8775,N_7144);
or U10764 (N_10764,N_8226,N_8332);
nand U10765 (N_10765,N_5140,N_5215);
nor U10766 (N_10766,N_6687,N_6796);
and U10767 (N_10767,N_6285,N_7337);
or U10768 (N_10768,N_8985,N_5204);
nand U10769 (N_10769,N_8487,N_5669);
and U10770 (N_10770,N_5535,N_8838);
and U10771 (N_10771,N_7174,N_7919);
and U10772 (N_10772,N_9927,N_8619);
nor U10773 (N_10773,N_8829,N_7503);
nand U10774 (N_10774,N_8281,N_5750);
nor U10775 (N_10775,N_6147,N_9532);
and U10776 (N_10776,N_7880,N_9594);
or U10777 (N_10777,N_7860,N_7373);
xnor U10778 (N_10778,N_5157,N_7412);
nand U10779 (N_10779,N_9184,N_9227);
nor U10780 (N_10780,N_8208,N_7133);
xor U10781 (N_10781,N_5163,N_8803);
or U10782 (N_10782,N_6866,N_6192);
nor U10783 (N_10783,N_7505,N_7762);
nor U10784 (N_10784,N_7079,N_5314);
nor U10785 (N_10785,N_7848,N_5088);
nand U10786 (N_10786,N_8679,N_7571);
nor U10787 (N_10787,N_8565,N_8345);
or U10788 (N_10788,N_8889,N_6817);
or U10789 (N_10789,N_6618,N_9360);
nand U10790 (N_10790,N_8523,N_9698);
or U10791 (N_10791,N_6983,N_6779);
nor U10792 (N_10792,N_7391,N_9036);
nor U10793 (N_10793,N_9277,N_7499);
nand U10794 (N_10794,N_7021,N_5654);
and U10795 (N_10795,N_7575,N_7276);
nor U10796 (N_10796,N_8380,N_7837);
nand U10797 (N_10797,N_8489,N_9900);
or U10798 (N_10798,N_5472,N_8948);
nand U10799 (N_10799,N_7278,N_7086);
or U10800 (N_10800,N_9006,N_9219);
nor U10801 (N_10801,N_6719,N_7316);
nand U10802 (N_10802,N_6343,N_9032);
nor U10803 (N_10803,N_6418,N_5355);
or U10804 (N_10804,N_7296,N_8894);
or U10805 (N_10805,N_7308,N_8712);
and U10806 (N_10806,N_6816,N_8374);
nor U10807 (N_10807,N_8247,N_9095);
nand U10808 (N_10808,N_6652,N_7440);
or U10809 (N_10809,N_9216,N_5890);
and U10810 (N_10810,N_8834,N_8791);
nand U10811 (N_10811,N_9649,N_5468);
and U10812 (N_10812,N_8779,N_7903);
or U10813 (N_10813,N_7777,N_6750);
and U10814 (N_10814,N_5740,N_7320);
nand U10815 (N_10815,N_7716,N_5095);
or U10816 (N_10816,N_8839,N_6138);
or U10817 (N_10817,N_6700,N_5774);
and U10818 (N_10818,N_7718,N_5673);
nand U10819 (N_10819,N_9237,N_7357);
or U10820 (N_10820,N_8903,N_9735);
or U10821 (N_10821,N_8424,N_8792);
and U10822 (N_10822,N_8401,N_9906);
nand U10823 (N_10823,N_5742,N_7823);
nand U10824 (N_10824,N_6742,N_6671);
and U10825 (N_10825,N_9521,N_9588);
or U10826 (N_10826,N_6987,N_5772);
or U10827 (N_10827,N_5650,N_5725);
nor U10828 (N_10828,N_8180,N_7160);
nor U10829 (N_10829,N_5446,N_9788);
nand U10830 (N_10830,N_5670,N_6258);
and U10831 (N_10831,N_8946,N_8182);
xor U10832 (N_10832,N_7345,N_9332);
or U10833 (N_10833,N_8783,N_8384);
and U10834 (N_10834,N_8895,N_5226);
and U10835 (N_10835,N_5544,N_5566);
and U10836 (N_10836,N_6756,N_7925);
or U10837 (N_10837,N_5904,N_7020);
nor U10838 (N_10838,N_6585,N_8402);
and U10839 (N_10839,N_5340,N_9922);
and U10840 (N_10840,N_6688,N_5292);
nor U10841 (N_10841,N_8198,N_6937);
nand U10842 (N_10842,N_9353,N_6941);
and U10843 (N_10843,N_5171,N_9821);
xnor U10844 (N_10844,N_9533,N_7678);
or U10845 (N_10845,N_9432,N_9343);
nor U10846 (N_10846,N_7431,N_8290);
or U10847 (N_10847,N_9040,N_9901);
and U10848 (N_10848,N_7878,N_6655);
xor U10849 (N_10849,N_6492,N_7068);
nand U10850 (N_10850,N_5560,N_7325);
and U10851 (N_10851,N_6644,N_8645);
or U10852 (N_10852,N_5806,N_7523);
nand U10853 (N_10853,N_7059,N_8186);
or U10854 (N_10854,N_7621,N_7914);
or U10855 (N_10855,N_7773,N_8038);
or U10856 (N_10856,N_6012,N_5668);
nand U10857 (N_10857,N_8263,N_9819);
nor U10858 (N_10858,N_7444,N_5601);
nor U10859 (N_10859,N_7517,N_6991);
xnor U10860 (N_10860,N_9496,N_8304);
nor U10861 (N_10861,N_6723,N_5557);
and U10862 (N_10862,N_7245,N_5029);
nand U10863 (N_10863,N_9053,N_7421);
nor U10864 (N_10864,N_5217,N_6239);
and U10865 (N_10865,N_7419,N_8245);
and U10866 (N_10866,N_6278,N_7014);
or U10867 (N_10867,N_5696,N_5761);
and U10868 (N_10868,N_6928,N_5405);
and U10869 (N_10869,N_6405,N_7388);
and U10870 (N_10870,N_7839,N_6547);
nor U10871 (N_10871,N_5836,N_5174);
or U10872 (N_10872,N_7162,N_8586);
and U10873 (N_10873,N_5957,N_9243);
xnor U10874 (N_10874,N_7213,N_5104);
nor U10875 (N_10875,N_9840,N_8996);
xor U10876 (N_10876,N_7627,N_5754);
nor U10877 (N_10877,N_7292,N_8069);
or U10878 (N_10878,N_9695,N_7827);
nand U10879 (N_10879,N_8623,N_8079);
nor U10880 (N_10880,N_9822,N_7785);
nand U10881 (N_10881,N_9593,N_9782);
nand U10882 (N_10882,N_9742,N_9890);
nor U10883 (N_10883,N_8660,N_8721);
and U10884 (N_10884,N_6701,N_5121);
nor U10885 (N_10885,N_8232,N_7512);
xor U10886 (N_10886,N_7549,N_7053);
nand U10887 (N_10887,N_7460,N_5237);
nor U10888 (N_10888,N_8538,N_5416);
and U10889 (N_10889,N_9477,N_5447);
nand U10890 (N_10890,N_9952,N_8582);
and U10891 (N_10891,N_7585,N_5854);
nand U10892 (N_10892,N_8275,N_8609);
or U10893 (N_10893,N_9874,N_9721);
and U10894 (N_10894,N_9046,N_5736);
or U10895 (N_10895,N_6204,N_6462);
nor U10896 (N_10896,N_8597,N_5398);
nor U10897 (N_10897,N_9709,N_8484);
nand U10898 (N_10898,N_8883,N_6578);
or U10899 (N_10899,N_7310,N_9389);
and U10900 (N_10900,N_8578,N_9467);
and U10901 (N_10901,N_6968,N_9417);
or U10902 (N_10902,N_8029,N_5507);
or U10903 (N_10903,N_5211,N_8727);
or U10904 (N_10904,N_9755,N_8162);
or U10905 (N_10905,N_8240,N_8378);
and U10906 (N_10906,N_9397,N_6725);
or U10907 (N_10907,N_8068,N_6379);
and U10908 (N_10908,N_5831,N_8369);
or U10909 (N_10909,N_5118,N_9917);
nor U10910 (N_10910,N_5169,N_6160);
nand U10911 (N_10911,N_7269,N_7476);
or U10912 (N_10912,N_7464,N_6395);
and U10913 (N_10913,N_5979,N_9941);
nor U10914 (N_10914,N_8126,N_9955);
nand U10915 (N_10915,N_7969,N_6099);
nand U10916 (N_10916,N_6120,N_8189);
and U10917 (N_10917,N_6302,N_8417);
nand U10918 (N_10918,N_7096,N_7623);
or U10919 (N_10919,N_6027,N_9104);
nor U10920 (N_10920,N_7788,N_7661);
and U10921 (N_10921,N_6057,N_5719);
or U10922 (N_10922,N_5265,N_6222);
or U10923 (N_10923,N_7764,N_9615);
or U10924 (N_10924,N_9424,N_6764);
xor U10925 (N_10925,N_8951,N_7439);
nor U10926 (N_10926,N_5505,N_8035);
or U10927 (N_10927,N_8512,N_8600);
or U10928 (N_10928,N_9754,N_8849);
and U10929 (N_10929,N_6746,N_8363);
nor U10930 (N_10930,N_8084,N_5912);
or U10931 (N_10931,N_7350,N_9462);
nand U10932 (N_10932,N_5697,N_6717);
or U10933 (N_10933,N_5857,N_9488);
nand U10934 (N_10934,N_6358,N_8195);
or U10935 (N_10935,N_6907,N_6449);
xor U10936 (N_10936,N_5469,N_9677);
nand U10937 (N_10937,N_9926,N_5967);
xnor U10938 (N_10938,N_6296,N_8914);
nor U10939 (N_10939,N_5154,N_6721);
nand U10940 (N_10940,N_8170,N_7671);
nor U10941 (N_10941,N_8642,N_6532);
nand U10942 (N_10942,N_6247,N_8353);
nand U10943 (N_10943,N_9513,N_9298);
or U10944 (N_10944,N_7667,N_7155);
nor U10945 (N_10945,N_8016,N_5032);
and U10946 (N_10946,N_9474,N_7076);
nand U10947 (N_10947,N_9564,N_5200);
and U10948 (N_10948,N_7589,N_7840);
and U10949 (N_10949,N_6931,N_8638);
or U10950 (N_10950,N_9739,N_5923);
nand U10951 (N_10951,N_7274,N_9679);
or U10952 (N_10952,N_9851,N_6729);
and U10953 (N_10953,N_6374,N_9825);
and U10954 (N_10954,N_7414,N_5634);
or U10955 (N_10955,N_7761,N_9262);
nand U10956 (N_10956,N_7924,N_7936);
nand U10957 (N_10957,N_6250,N_5048);
nand U10958 (N_10958,N_7487,N_8628);
nor U10959 (N_10959,N_6115,N_5563);
nor U10960 (N_10960,N_8960,N_6075);
nor U10961 (N_10961,N_6517,N_5061);
xnor U10962 (N_10962,N_8108,N_9391);
and U10963 (N_10963,N_7995,N_8366);
nor U10964 (N_10964,N_6724,N_8585);
xor U10965 (N_10965,N_6832,N_8994);
or U10966 (N_10966,N_6999,N_8009);
or U10967 (N_10967,N_9680,N_9131);
nand U10968 (N_10968,N_7369,N_7569);
and U10969 (N_10969,N_7362,N_5444);
nand U10970 (N_10970,N_5769,N_8190);
nand U10971 (N_10971,N_7989,N_6366);
or U10972 (N_10972,N_7844,N_6830);
and U10973 (N_10973,N_8483,N_6589);
and U10974 (N_10974,N_7728,N_8364);
nor U10975 (N_10975,N_8111,N_6328);
nand U10976 (N_10976,N_5075,N_6233);
xnor U10977 (N_10977,N_7116,N_9714);
or U10978 (N_10978,N_7453,N_9650);
nand U10979 (N_10979,N_9174,N_8117);
and U10980 (N_10980,N_9724,N_8455);
nand U10981 (N_10981,N_5993,N_5881);
nor U10982 (N_10982,N_8076,N_7230);
and U10983 (N_10983,N_8710,N_6990);
nand U10984 (N_10984,N_5941,N_7991);
nor U10985 (N_10985,N_7145,N_8514);
and U10986 (N_10986,N_8817,N_8581);
nand U10987 (N_10987,N_6213,N_7729);
and U10988 (N_10988,N_8036,N_7672);
xor U10989 (N_10989,N_7905,N_5083);
and U10990 (N_10990,N_9134,N_9136);
xnor U10991 (N_10991,N_5164,N_9411);
or U10992 (N_10992,N_6520,N_5978);
nor U10993 (N_10993,N_8056,N_8433);
and U10994 (N_10994,N_5883,N_7803);
nor U10995 (N_10995,N_9418,N_6164);
or U10996 (N_10996,N_8415,N_8555);
and U10997 (N_10997,N_9523,N_5571);
nand U10998 (N_10998,N_6026,N_9090);
or U10999 (N_10999,N_8897,N_6510);
nor U11000 (N_11000,N_5629,N_5360);
or U11001 (N_11001,N_6868,N_5427);
or U11002 (N_11002,N_7261,N_5520);
nor U11003 (N_11003,N_6890,N_6643);
and U11004 (N_11004,N_5888,N_8207);
nand U11005 (N_11005,N_7041,N_8896);
and U11006 (N_11006,N_7273,N_5944);
nor U11007 (N_11007,N_8548,N_8218);
nor U11008 (N_11008,N_9688,N_6177);
nor U11009 (N_11009,N_6544,N_5053);
or U11010 (N_11010,N_8980,N_8568);
nand U11011 (N_11011,N_6838,N_6474);
nor U11012 (N_11012,N_5626,N_5197);
nor U11013 (N_11013,N_9414,N_6197);
and U11014 (N_11014,N_8785,N_9845);
nor U11015 (N_11015,N_8161,N_9033);
nand U11016 (N_11016,N_8437,N_8656);
or U11017 (N_11017,N_7963,N_5951);
or U11018 (N_11018,N_5365,N_5800);
nor U11019 (N_11019,N_7277,N_5170);
and U11020 (N_11020,N_9486,N_9259);
or U11021 (N_11021,N_6683,N_8541);
and U11022 (N_11022,N_6082,N_9928);
nor U11023 (N_11023,N_7871,N_5724);
or U11024 (N_11024,N_9558,N_8171);
and U11025 (N_11025,N_7998,N_5390);
nor U11026 (N_11026,N_7207,N_6131);
nor U11027 (N_11027,N_6762,N_7551);
nand U11028 (N_11028,N_9167,N_9682);
or U11029 (N_11029,N_9494,N_9034);
xnor U11030 (N_11030,N_6965,N_6047);
nand U11031 (N_11031,N_5407,N_8204);
nor U11032 (N_11032,N_9497,N_5581);
xor U11033 (N_11033,N_6194,N_7567);
nor U11034 (N_11034,N_6946,N_5549);
and U11035 (N_11035,N_9038,N_5989);
nor U11036 (N_11036,N_7420,N_8666);
or U11037 (N_11037,N_6776,N_5339);
nor U11038 (N_11038,N_8730,N_6461);
and U11039 (N_11039,N_5684,N_6633);
or U11040 (N_11040,N_8310,N_8678);
nand U11041 (N_11041,N_9956,N_7189);
nand U11042 (N_11042,N_9260,N_6351);
or U11043 (N_11043,N_6953,N_8061);
nand U11044 (N_11044,N_8554,N_8692);
or U11045 (N_11045,N_6479,N_8669);
nor U11046 (N_11046,N_7654,N_6925);
or U11047 (N_11047,N_7733,N_9800);
nand U11048 (N_11048,N_8357,N_7715);
nor U11049 (N_11049,N_5328,N_8673);
nand U11050 (N_11050,N_7942,N_6344);
nand U11051 (N_11051,N_9983,N_7238);
nor U11052 (N_11052,N_8325,N_5558);
and U11053 (N_11053,N_8491,N_8128);
and U11054 (N_11054,N_9354,N_6942);
and U11055 (N_11055,N_5787,N_7215);
nand U11056 (N_11056,N_8539,N_9545);
nor U11057 (N_11057,N_9214,N_8019);
or U11058 (N_11058,N_5250,N_9508);
and U11059 (N_11059,N_9464,N_5442);
or U11060 (N_11060,N_9657,N_5846);
or U11061 (N_11061,N_6821,N_7592);
nand U11062 (N_11062,N_9153,N_8469);
and U11063 (N_11063,N_7666,N_9400);
nand U11064 (N_11064,N_5589,N_5073);
and U11065 (N_11065,N_7148,N_8075);
or U11066 (N_11066,N_7011,N_8416);
nor U11067 (N_11067,N_6790,N_5636);
nand U11068 (N_11068,N_5381,N_5906);
nor U11069 (N_11069,N_6268,N_9823);
nor U11070 (N_11070,N_5123,N_8862);
and U11071 (N_11071,N_6301,N_9765);
nand U11072 (N_11072,N_6512,N_9258);
nand U11073 (N_11073,N_5714,N_5695);
or U11074 (N_11074,N_7617,N_8611);
nand U11075 (N_11075,N_9770,N_6400);
or U11076 (N_11076,N_6595,N_5841);
nand U11077 (N_11077,N_6989,N_8668);
nand U11078 (N_11078,N_8912,N_5573);
nand U11079 (N_11079,N_7129,N_6748);
nor U11080 (N_11080,N_9816,N_5412);
or U11081 (N_11081,N_8379,N_6529);
or U11082 (N_11082,N_6095,N_9620);
nand U11083 (N_11083,N_8709,N_5771);
nor U11084 (N_11084,N_9252,N_6751);
and U11085 (N_11085,N_6130,N_7038);
or U11086 (N_11086,N_7524,N_8328);
nand U11087 (N_11087,N_9188,N_8929);
nand U11088 (N_11088,N_6333,N_8081);
nor U11089 (N_11089,N_9169,N_5529);
or U11090 (N_11090,N_5238,N_6471);
nand U11091 (N_11091,N_6364,N_7010);
and U11092 (N_11092,N_8651,N_9439);
and U11093 (N_11093,N_8641,N_9202);
or U11094 (N_11094,N_8685,N_9316);
nor U11095 (N_11095,N_8940,N_8073);
nand U11096 (N_11096,N_5984,N_8966);
nor U11097 (N_11097,N_7085,N_9171);
and U11098 (N_11098,N_6434,N_9561);
nor U11099 (N_11099,N_9539,N_7656);
nand U11100 (N_11100,N_7172,N_6331);
xor U11101 (N_11101,N_8308,N_5054);
and U11102 (N_11102,N_6311,N_6581);
nand U11103 (N_11103,N_7449,N_6698);
nand U11104 (N_11104,N_8594,N_7224);
or U11105 (N_11105,N_8479,N_6601);
and U11106 (N_11106,N_7815,N_9889);
xor U11107 (N_11107,N_6845,N_8271);
or U11108 (N_11108,N_8370,N_7838);
nand U11109 (N_11109,N_5965,N_8703);
nand U11110 (N_11110,N_9820,N_8018);
nand U11111 (N_11111,N_5267,N_6299);
nor U11112 (N_11112,N_8481,N_8432);
xor U11113 (N_11113,N_6041,N_6320);
nand U11114 (N_11114,N_5106,N_7275);
or U11115 (N_11115,N_5475,N_7752);
nand U11116 (N_11116,N_9055,N_7473);
or U11117 (N_11117,N_6640,N_9468);
nor U11118 (N_11118,N_9610,N_7953);
or U11119 (N_11119,N_9614,N_9831);
nand U11120 (N_11120,N_7861,N_6911);
nand U11121 (N_11121,N_9716,N_6747);
or U11122 (N_11122,N_6857,N_7175);
nand U11123 (N_11123,N_7248,N_9863);
nor U11124 (N_11124,N_9723,N_9812);
and U11125 (N_11125,N_6402,N_9824);
nand U11126 (N_11126,N_7832,N_5796);
nor U11127 (N_11127,N_6098,N_9538);
or U11128 (N_11128,N_6260,N_6252);
nor U11129 (N_11129,N_6495,N_6505);
and U11130 (N_11130,N_5385,N_8337);
nor U11131 (N_11131,N_5388,N_8756);
nand U11132 (N_11132,N_8130,N_7185);
and U11133 (N_11133,N_8935,N_5410);
nor U11134 (N_11134,N_7354,N_6908);
and U11135 (N_11135,N_9146,N_8916);
and U11136 (N_11136,N_9152,N_9909);
and U11137 (N_11137,N_6548,N_9648);
xor U11138 (N_11138,N_5633,N_9452);
or U11139 (N_11139,N_6208,N_8816);
nand U11140 (N_11140,N_6426,N_7005);
nand U11141 (N_11141,N_7829,N_9073);
xnor U11142 (N_11142,N_9703,N_8472);
or U11143 (N_11143,N_7025,N_9684);
nor U11144 (N_11144,N_7993,N_9209);
and U11145 (N_11145,N_8558,N_7425);
xnor U11146 (N_11146,N_9996,N_5198);
nor U11147 (N_11147,N_8154,N_5528);
nor U11148 (N_11148,N_9466,N_9035);
nor U11149 (N_11149,N_5795,N_5166);
nand U11150 (N_11150,N_5717,N_7072);
or U11151 (N_11151,N_8880,N_6891);
or U11152 (N_11152,N_8821,N_6936);
or U11153 (N_11153,N_6347,N_8302);
nand U11154 (N_11154,N_8474,N_8179);
or U11155 (N_11155,N_6506,N_6335);
and U11156 (N_11156,N_7394,N_6334);
or U11157 (N_11157,N_6009,N_6420);
or U11158 (N_11158,N_6781,N_9830);
nor U11159 (N_11159,N_7443,N_6338);
and U11160 (N_11160,N_5421,N_7622);
nand U11161 (N_11161,N_9276,N_9337);
xnor U11162 (N_11162,N_6770,N_6454);
and U11163 (N_11163,N_6256,N_7000);
and U11164 (N_11164,N_7690,N_9987);
nor U11165 (N_11165,N_8244,N_7300);
or U11166 (N_11166,N_9505,N_7821);
and U11167 (N_11167,N_8234,N_9839);
nand U11168 (N_11168,N_7632,N_9603);
xor U11169 (N_11169,N_6352,N_9244);
xor U11170 (N_11170,N_5820,N_6446);
nand U11171 (N_11171,N_7170,N_9774);
or U11172 (N_11172,N_5244,N_8653);
or U11173 (N_11173,N_6526,N_8105);
nor U11174 (N_11174,N_7322,N_9888);
nand U11175 (N_11175,N_9223,N_6478);
or U11176 (N_11176,N_5614,N_9768);
and U11177 (N_11177,N_6772,N_9995);
and U11178 (N_11178,N_8515,N_9067);
or U11179 (N_11179,N_5788,N_5422);
or U11180 (N_11180,N_7198,N_6679);
and U11181 (N_11181,N_5269,N_6704);
xnor U11182 (N_11182,N_6562,N_8203);
xnor U11183 (N_11183,N_5891,N_8873);
nor U11184 (N_11184,N_6635,N_8276);
nor U11185 (N_11185,N_9548,N_7400);
or U11186 (N_11186,N_8945,N_6697);
xnor U11187 (N_11187,N_8533,N_9977);
nor U11188 (N_11188,N_5781,N_6584);
nor U11189 (N_11189,N_8553,N_8590);
nor U11190 (N_11190,N_7849,N_8303);
or U11191 (N_11191,N_5408,N_9238);
or U11192 (N_11192,N_8989,N_8285);
xor U11193 (N_11193,N_9946,N_6629);
nor U11194 (N_11194,N_5389,N_9715);
xor U11195 (N_11195,N_5746,N_8291);
nor U11196 (N_11196,N_9321,N_5643);
and U11197 (N_11197,N_7418,N_7677);
nand U11198 (N_11198,N_5556,N_8714);
nand U11199 (N_11199,N_9573,N_9162);
and U11200 (N_11200,N_5612,N_6567);
and U11201 (N_11201,N_5982,N_9412);
or U11202 (N_11202,N_7511,N_5737);
nor U11203 (N_11203,N_7241,N_9719);
and U11204 (N_11204,N_7353,N_5445);
nand U11205 (N_11205,N_6744,N_6885);
nand U11206 (N_11206,N_9013,N_6918);
and U11207 (N_11207,N_6843,N_6481);
xor U11208 (N_11208,N_5956,N_9088);
or U11209 (N_11209,N_7488,N_7267);
nand U11210 (N_11210,N_6703,N_8367);
nor U11211 (N_11211,N_5417,N_6178);
xnor U11212 (N_11212,N_5793,N_5189);
and U11213 (N_11213,N_5177,N_5024);
nor U11214 (N_11214,N_5845,N_8532);
or U11215 (N_11215,N_5813,N_6220);
xor U11216 (N_11216,N_9781,N_5258);
or U11217 (N_11217,N_9351,N_8132);
nand U11218 (N_11218,N_8837,N_6103);
nand U11219 (N_11219,N_8720,N_6094);
or U11220 (N_11220,N_5597,N_8686);
and U11221 (N_11221,N_5663,N_9344);
nor U11222 (N_11222,N_6384,N_8261);
or U11223 (N_11223,N_6269,N_7745);
nor U11224 (N_11224,N_5313,N_6722);
nor U11225 (N_11225,N_5464,N_8449);
nor U11226 (N_11226,N_9667,N_8907);
or U11227 (N_11227,N_8340,N_6122);
or U11228 (N_11228,N_7907,N_8905);
and U11229 (N_11229,N_5537,N_8967);
and U11230 (N_11230,N_5194,N_9186);
or U11231 (N_11231,N_8987,N_6415);
nand U11232 (N_11232,N_8722,N_8654);
xor U11233 (N_11233,N_8906,N_9644);
or U11234 (N_11234,N_9103,N_5681);
nand U11235 (N_11235,N_7819,N_5578);
or U11236 (N_11236,N_7070,N_8443);
nand U11237 (N_11237,N_8748,N_6771);
xor U11238 (N_11238,N_9849,N_5792);
and U11239 (N_11239,N_9415,N_8184);
nor U11240 (N_11240,N_6190,N_8030);
xor U11241 (N_11241,N_5959,N_5352);
nor U11242 (N_11242,N_9308,N_9168);
and U11243 (N_11243,N_5023,N_8707);
xor U11244 (N_11244,N_8930,N_7237);
xor U11245 (N_11245,N_7888,N_6383);
nand U11246 (N_11246,N_8644,N_5333);
or U11247 (N_11247,N_5858,N_8521);
nor U11248 (N_11248,N_9756,N_9226);
nand U11249 (N_11249,N_9619,N_9047);
nand U11250 (N_11250,N_6572,N_5235);
xnor U11251 (N_11251,N_7870,N_8269);
nand U11252 (N_11252,N_9595,N_9645);
xnor U11253 (N_11253,N_5409,N_6422);
nand U11254 (N_11254,N_8606,N_9119);
or U11255 (N_11255,N_6988,N_6306);
xnor U11256 (N_11256,N_7263,N_6355);
nor U11257 (N_11257,N_7381,N_6621);
nand U11258 (N_11258,N_7608,N_9589);
nor U11259 (N_11259,N_8864,N_5162);
nor U11260 (N_11260,N_9876,N_9182);
or U11261 (N_11261,N_6777,N_8093);
xnor U11262 (N_11262,N_9356,N_8225);
xor U11263 (N_11263,N_9205,N_9093);
xor U11264 (N_11264,N_9272,N_6874);
and U11265 (N_11265,N_7560,N_7977);
or U11266 (N_11266,N_9574,N_5233);
or U11267 (N_11267,N_8219,N_5000);
and U11268 (N_11268,N_5758,N_5097);
xor U11269 (N_11269,N_8059,N_7471);
or U11270 (N_11270,N_6642,N_6901);
nor U11271 (N_11271,N_7578,N_8827);
nor U11272 (N_11272,N_5449,N_9266);
nor U11273 (N_11273,N_9937,N_7219);
xor U11274 (N_11274,N_7056,N_8626);
nand U11275 (N_11275,N_5011,N_9263);
nor U11276 (N_11276,N_5439,N_6236);
nor U11277 (N_11277,N_9437,N_6036);
and U11278 (N_11278,N_9738,N_5839);
nand U11279 (N_11279,N_7675,N_7895);
nor U11280 (N_11280,N_7933,N_5675);
nor U11281 (N_11281,N_5028,N_7873);
and U11282 (N_11282,N_6087,N_7386);
nand U11283 (N_11283,N_9208,N_5778);
and U11284 (N_11284,N_9295,N_8690);
and U11285 (N_11285,N_7252,N_6951);
and U11286 (N_11286,N_7009,N_6831);
or U11287 (N_11287,N_5441,N_8008);
nor U11288 (N_11288,N_9196,N_6668);
or U11289 (N_11289,N_7375,N_5595);
or U11290 (N_11290,N_6673,N_5055);
and U11291 (N_11291,N_7490,N_9837);
or U11292 (N_11292,N_9440,N_5734);
nor U11293 (N_11293,N_8504,N_7614);
and U11294 (N_11294,N_6557,N_8693);
or U11295 (N_11295,N_9406,N_9048);
or U11296 (N_11296,N_5809,N_5705);
and U11297 (N_11297,N_7268,N_9495);
and U11298 (N_11298,N_5089,N_6113);
and U11299 (N_11299,N_9394,N_8683);
nor U11300 (N_11300,N_7772,N_5763);
nand U11301 (N_11301,N_6282,N_8636);
nor U11302 (N_11302,N_5050,N_8205);
nand U11303 (N_11303,N_7452,N_9925);
or U11304 (N_11304,N_5277,N_7749);
nor U11305 (N_11305,N_5972,N_6246);
and U11306 (N_11306,N_5346,N_6802);
nor U11307 (N_11307,N_6086,N_7529);
and U11308 (N_11308,N_7210,N_5255);
and U11309 (N_11309,N_6982,N_5735);
nand U11310 (N_11310,N_7050,N_9913);
or U11311 (N_11311,N_6726,N_5933);
and U11312 (N_11312,N_8598,N_7824);
nand U11313 (N_11313,N_6068,N_9775);
nand U11314 (N_11314,N_7674,N_5559);
or U11315 (N_11315,N_6893,N_7384);
or U11316 (N_11316,N_8041,N_8979);
or U11317 (N_11317,N_8843,N_6323);
or U11318 (N_11318,N_6682,N_8887);
nand U11319 (N_11319,N_6955,N_8411);
xor U11320 (N_11320,N_9016,N_8004);
and U11321 (N_11321,N_9070,N_8614);
and U11322 (N_11322,N_5335,N_6054);
or U11323 (N_11323,N_9313,N_7243);
or U11324 (N_11324,N_6266,N_9828);
nor U11325 (N_11325,N_9519,N_8757);
or U11326 (N_11326,N_6718,N_6758);
and U11327 (N_11327,N_5324,N_6780);
nand U11328 (N_11328,N_5689,N_7217);
or U11329 (N_11329,N_9100,N_9629);
or U11330 (N_11330,N_5273,N_8891);
nor U11331 (N_11331,N_8298,N_5728);
nor U11332 (N_11332,N_5008,N_7736);
nor U11333 (N_11333,N_9352,N_8595);
nand U11334 (N_11334,N_7628,N_6145);
nor U11335 (N_11335,N_6658,N_5718);
or U11336 (N_11336,N_9663,N_8969);
nand U11337 (N_11337,N_9292,N_6417);
nand U11338 (N_11338,N_6628,N_9319);
nand U11339 (N_11339,N_7506,N_6497);
xor U11340 (N_11340,N_6978,N_6900);
nor U11341 (N_11341,N_7434,N_7854);
xnor U11342 (N_11342,N_8027,N_5221);
or U11343 (N_11343,N_8859,N_7746);
and U11344 (N_11344,N_9037,N_7087);
nor U11345 (N_11345,N_9507,N_9459);
and U11346 (N_11346,N_8499,N_5383);
nor U11347 (N_11347,N_9692,N_5970);
nand U11348 (N_11348,N_8319,N_8140);
nor U11349 (N_11349,N_7204,N_8737);
or U11350 (N_11350,N_5014,N_5371);
and U11351 (N_11351,N_7134,N_8498);
nor U11352 (N_11352,N_5851,N_7132);
and U11353 (N_11353,N_9915,N_8520);
nor U11354 (N_11354,N_9191,N_5309);
or U11355 (N_11355,N_8254,N_7876);
nor U11356 (N_11356,N_9375,N_9066);
nor U11357 (N_11357,N_8993,N_8824);
and U11358 (N_11358,N_8574,N_5682);
and U11359 (N_11359,N_8355,N_5299);
nand U11360 (N_11360,N_7972,N_8836);
and U11361 (N_11361,N_9105,N_6531);
or U11362 (N_11362,N_5184,N_9687);
or U11363 (N_11363,N_8627,N_8457);
nand U11364 (N_11364,N_7339,N_5721);
nand U11365 (N_11365,N_9245,N_8938);
nand U11366 (N_11366,N_5122,N_7682);
or U11367 (N_11367,N_7744,N_5848);
and U11368 (N_11368,N_5627,N_5637);
or U11369 (N_11369,N_8178,N_7115);
and U11370 (N_11370,N_6317,N_6175);
nor U11371 (N_11371,N_7753,N_6459);
nand U11372 (N_11372,N_6412,N_9689);
or U11373 (N_11373,N_5354,N_7754);
and U11374 (N_11374,N_7480,N_5834);
nor U11375 (N_11375,N_6556,N_5329);
and U11376 (N_11376,N_5161,N_7882);
and U11377 (N_11377,N_7315,N_7520);
or U11378 (N_11378,N_6298,N_5720);
and U11379 (N_11379,N_8430,N_9636);
or U11380 (N_11380,N_8761,N_7486);
nor U11381 (N_11381,N_7579,N_9137);
xor U11382 (N_11382,N_7613,N_9625);
nand U11383 (N_11383,N_5864,N_9963);
xor U11384 (N_11384,N_9844,N_5564);
nor U11385 (N_11385,N_9628,N_8704);
nand U11386 (N_11386,N_6464,N_5126);
nor U11387 (N_11387,N_6881,N_8127);
xnor U11388 (N_11388,N_5256,N_5212);
xnor U11389 (N_11389,N_5550,N_9786);
nor U11390 (N_11390,N_7580,N_6552);
nor U11391 (N_11391,N_9808,N_6797);
and U11392 (N_11392,N_7390,N_7022);
or U11393 (N_11393,N_5766,N_8599);
xor U11394 (N_11394,N_7112,N_6496);
or U11395 (N_11395,N_6111,N_8579);
nand U11396 (N_11396,N_9366,N_7408);
nand U11397 (N_11397,N_7100,N_6391);
xnor U11398 (N_11398,N_7552,N_5394);
nor U11399 (N_11399,N_7868,N_9541);
or U11400 (N_11400,N_8135,N_9121);
and U11401 (N_11401,N_9970,N_6408);
and U11402 (N_11402,N_8466,N_6972);
nor U11403 (N_11403,N_9029,N_6549);
nand U11404 (N_11404,N_9335,N_7563);
nor U11405 (N_11405,N_7182,N_8852);
or U11406 (N_11406,N_9499,N_7723);
nor U11407 (N_11407,N_8201,N_7526);
xor U11408 (N_11408,N_6691,N_6126);
nor U11409 (N_11409,N_8249,N_5234);
or U11410 (N_11410,N_9515,N_9195);
nand U11411 (N_11411,N_9965,N_9943);
nor U11412 (N_11412,N_6484,N_5271);
and U11413 (N_11413,N_8311,N_9056);
or U11414 (N_11414,N_8900,N_6159);
or U11415 (N_11415,N_7092,N_5030);
xnor U11416 (N_11416,N_7974,N_8643);
nand U11417 (N_11417,N_6692,N_8277);
or U11418 (N_11418,N_9207,N_6482);
or U11419 (N_11419,N_9396,N_5900);
nor U11420 (N_11420,N_6485,N_8796);
or U11421 (N_11421,N_7259,N_8637);
nand U11422 (N_11422,N_5044,N_9602);
and U11423 (N_11423,N_9431,N_6587);
nor U11424 (N_11424,N_7710,N_9144);
nand U11425 (N_11425,N_8759,N_5922);
xor U11426 (N_11426,N_5694,N_7498);
nor U11427 (N_11427,N_6167,N_8155);
nor U11428 (N_11428,N_7833,N_7813);
nor U11429 (N_11429,N_9854,N_8460);
nor U11430 (N_11430,N_9165,N_5649);
and U11431 (N_11431,N_5843,N_5730);
nand U11432 (N_11432,N_7285,N_9883);
and U11433 (N_11433,N_6826,N_9099);
xnor U11434 (N_11434,N_5641,N_8840);
and U11435 (N_11435,N_9479,N_5015);
and U11436 (N_11436,N_5065,N_5353);
nand U11437 (N_11437,N_9422,N_5648);
nand U11438 (N_11438,N_7371,N_7057);
or U11439 (N_11439,N_9711,N_7455);
or U11440 (N_11440,N_9531,N_9150);
and U11441 (N_11441,N_8798,N_6189);
nor U11442 (N_11442,N_7029,N_6005);
or U11443 (N_11443,N_5159,N_6060);
and U11444 (N_11444,N_7979,N_8390);
nor U11445 (N_11445,N_7411,N_9393);
or U11446 (N_11446,N_7805,N_5223);
nor U11447 (N_11447,N_9410,N_7696);
nor U11448 (N_11448,N_7652,N_5918);
nor U11449 (N_11449,N_6666,N_6069);
and U11450 (N_11450,N_5359,N_5391);
or U11451 (N_11451,N_7660,N_9678);
nand U11452 (N_11452,N_8830,N_6824);
and U11453 (N_11453,N_9551,N_6499);
or U11454 (N_11454,N_9892,N_8419);
nor U11455 (N_11455,N_7826,N_5977);
or U11456 (N_11456,N_7765,N_7107);
and U11457 (N_11457,N_7232,N_7902);
nor U11458 (N_11458,N_7060,N_7200);
or U11459 (N_11459,N_6017,N_9470);
nand U11460 (N_11460,N_8815,N_6388);
or U11461 (N_11461,N_8486,N_5882);
xor U11462 (N_11462,N_5647,N_6329);
or U11463 (N_11463,N_7668,N_7378);
nor U11464 (N_11464,N_9385,N_7178);
and U11465 (N_11465,N_7798,N_8734);
xnor U11466 (N_11466,N_9027,N_6445);
xnor U11467 (N_11467,N_5470,N_8911);
or U11468 (N_11468,N_9967,N_6920);
nor U11469 (N_11469,N_9408,N_9234);
or U11470 (N_11470,N_9771,N_9269);
nor U11471 (N_11471,N_9976,N_5553);
and U11472 (N_11472,N_5958,N_6172);
or U11473 (N_11473,N_8725,N_7075);
nand U11474 (N_11474,N_8167,N_6169);
nor U11475 (N_11475,N_8315,N_7206);
and U11476 (N_11476,N_5300,N_6143);
and U11477 (N_11477,N_9524,N_7141);
or U11478 (N_11478,N_7912,N_6173);
nand U11479 (N_11479,N_5110,N_9051);
and U11480 (N_11480,N_7104,N_5046);
or U11481 (N_11481,N_7179,N_5869);
and U11482 (N_11482,N_6466,N_5876);
and U11483 (N_11483,N_5671,N_6199);
nand U11484 (N_11484,N_6089,N_9071);
nor U11485 (N_11485,N_6783,N_7317);
nor U11486 (N_11486,N_6916,N_5554);
and U11487 (N_11487,N_7437,N_8408);
and U11488 (N_11488,N_6288,N_5183);
or U11489 (N_11489,N_7321,N_6808);
nand U11490 (N_11490,N_7428,N_5539);
or U11491 (N_11491,N_5245,N_7140);
or U11492 (N_11492,N_8392,N_8784);
nand U11493 (N_11493,N_5495,N_5397);
nor U11494 (N_11494,N_7493,N_6507);
nand U11495 (N_11495,N_6021,N_7365);
and U11496 (N_11496,N_8322,N_5100);
and U11497 (N_11497,N_6690,N_5751);
nor U11498 (N_11498,N_8376,N_9110);
and U11499 (N_11499,N_9478,N_9807);
and U11500 (N_11500,N_5832,N_5630);
xor U11501 (N_11501,N_9855,N_9606);
nand U11502 (N_11502,N_8492,N_6072);
and U11503 (N_11503,N_9861,N_5782);
nand U11504 (N_11504,N_9990,N_6869);
nor U11505 (N_11505,N_6139,N_5229);
or U11506 (N_11506,N_7067,N_7264);
nand U11507 (N_11507,N_8407,N_9426);
nand U11508 (N_11508,N_5266,N_6313);
nor U11509 (N_11509,N_5378,N_8048);
xor U11510 (N_11510,N_8657,N_6325);
and U11511 (N_11511,N_7004,N_6275);
or U11512 (N_11512,N_7562,N_8502);
nor U11513 (N_11513,N_8743,N_8239);
and U11514 (N_11514,N_7717,N_6561);
xnor U11515 (N_11515,N_7229,N_7266);
nand U11516 (N_11516,N_6028,N_9921);
nor U11517 (N_11517,N_6985,N_8577);
and U11518 (N_11518,N_6674,N_6380);
or U11519 (N_11519,N_8146,N_9605);
nor U11520 (N_11520,N_9713,N_8456);
and U11521 (N_11521,N_5743,N_8500);
or U11522 (N_11522,N_6887,N_9370);
nand U11523 (N_11523,N_5213,N_8440);
xnor U11524 (N_11524,N_8557,N_8211);
and U11525 (N_11525,N_7023,N_8040);
nand U11526 (N_11526,N_5209,N_6133);
or U11527 (N_11527,N_5153,N_8461);
and U11528 (N_11528,N_5672,N_5225);
or U11529 (N_11529,N_9102,N_9759);
nand U11530 (N_11530,N_8242,N_7760);
nand U11531 (N_11531,N_6504,N_7693);
nor U11532 (N_11532,N_9109,N_6922);
nand U11533 (N_11533,N_6046,N_9933);
or U11534 (N_11534,N_7518,N_7024);
xnor U11535 (N_11535,N_9877,N_8314);
or U11536 (N_11536,N_9065,N_7139);
nor U11537 (N_11537,N_6678,N_8580);
or U11538 (N_11538,N_9510,N_9274);
and U11539 (N_11539,N_5160,N_7700);
and U11540 (N_11540,N_6413,N_6740);
and U11541 (N_11541,N_8439,N_9255);
nor U11542 (N_11542,N_8428,N_7748);
and U11543 (N_11543,N_7950,N_6847);
or U11544 (N_11544,N_5486,N_8090);
or U11545 (N_11545,N_5727,N_7078);
and U11546 (N_11546,N_5807,N_6217);
nand U11547 (N_11547,N_7319,N_7045);
nor U11548 (N_11548,N_9653,N_9130);
nor U11549 (N_11549,N_5311,N_7546);
and U11550 (N_11550,N_5369,N_7708);
nand U11551 (N_11551,N_5606,N_7624);
nand U11552 (N_11552,N_6914,N_6006);
and U11553 (N_11553,N_8478,N_9647);
nand U11554 (N_11554,N_8724,N_5483);
nor U11555 (N_11555,N_9997,N_8344);
nor U11556 (N_11556,N_6755,N_5262);
or U11557 (N_11557,N_6104,N_9815);
nand U11558 (N_11558,N_9506,N_9691);
nand U11559 (N_11559,N_7042,N_9005);
nor U11560 (N_11560,N_6187,N_9958);
nand U11561 (N_11561,N_6011,N_7859);
nand U11562 (N_11562,N_9059,N_7019);
xor U11563 (N_11563,N_7314,N_7801);
or U11564 (N_11564,N_7954,N_9149);
nand U11565 (N_11565,N_7513,N_8273);
and U11566 (N_11566,N_5819,N_7767);
or U11567 (N_11567,N_6828,N_7343);
or U11568 (N_11568,N_5243,N_5457);
nor U11569 (N_11569,N_5536,N_9322);
nand U11570 (N_11570,N_6102,N_6371);
and U11571 (N_11571,N_5949,N_5508);
nor U11572 (N_11572,N_9972,N_5236);
nand U11573 (N_11573,N_6889,N_6980);
nand U11574 (N_11574,N_6106,N_7040);
or U11575 (N_11575,N_8025,N_9261);
nand U11576 (N_11576,N_6568,N_6757);
and U11577 (N_11577,N_7817,N_8936);
nor U11578 (N_11578,N_7309,N_5619);
or U11579 (N_11579,N_8695,N_6033);
and U11580 (N_11580,N_9257,N_6494);
nor U11581 (N_11581,N_5016,N_8465);
nor U11582 (N_11582,N_9878,N_7737);
nand U11583 (N_11583,N_5357,N_8143);
or U11584 (N_11584,N_7117,N_8592);
and U11585 (N_11585,N_7405,N_9557);
and U11586 (N_11586,N_5950,N_9200);
nor U11587 (N_11587,N_6489,N_7235);
or U11588 (N_11588,N_9658,N_7077);
nand U11589 (N_11589,N_8509,N_5765);
and U11590 (N_11590,N_7239,N_7679);
or U11591 (N_11591,N_6811,N_5801);
nor U11592 (N_11592,N_8576,N_7120);
nand U11593 (N_11593,N_9115,N_9201);
nand U11594 (N_11594,N_7615,N_9656);
xnor U11595 (N_11595,N_6854,N_5454);
nand U11596 (N_11596,N_8742,N_8002);
or U11597 (N_11597,N_5574,N_8210);
xnor U11598 (N_11598,N_6812,N_9345);
or U11599 (N_11599,N_9157,N_5603);
or U11600 (N_11600,N_9842,N_9836);
and U11601 (N_11601,N_5492,N_7255);
and U11602 (N_11602,N_6451,N_9623);
nand U11603 (N_11603,N_7374,N_8191);
or U11604 (N_11604,N_5879,N_5562);
or U11605 (N_11605,N_7583,N_7706);
or U11606 (N_11606,N_7363,N_5117);
nor U11607 (N_11607,N_5272,N_9675);
nor U11608 (N_11608,N_9473,N_6397);
nor U11609 (N_11609,N_8183,N_8010);
and U11610 (N_11610,N_6229,N_5108);
or U11611 (N_11611,N_8350,N_6923);
xnor U11612 (N_11612,N_7843,N_5342);
nor U11613 (N_11613,N_6428,N_5731);
and U11614 (N_11614,N_8542,N_9599);
nor U11615 (N_11615,N_5203,N_5135);
nand U11616 (N_11616,N_7581,N_6316);
nor U11617 (N_11617,N_6709,N_9621);
or U11618 (N_11618,N_9669,N_6231);
nand U11619 (N_11619,N_5264,N_8187);
or U11620 (N_11620,N_9030,N_9172);
and U11621 (N_11621,N_6330,N_8556);
nor U11622 (N_11622,N_6944,N_9609);
and U11623 (N_11623,N_9395,N_6785);
nor U11624 (N_11624,N_9793,N_8699);
or U11625 (N_11625,N_8865,N_9179);
nor U11626 (N_11626,N_7454,N_6363);
and U11627 (N_11627,N_7964,N_7787);
xnor U11628 (N_11628,N_9870,N_8620);
or U11629 (N_11629,N_8527,N_6879);
nand U11630 (N_11630,N_7606,N_9300);
nand U11631 (N_11631,N_5775,N_5512);
or U11632 (N_11632,N_8120,N_5878);
or U11633 (N_11633,N_9438,N_7721);
or U11634 (N_11634,N_8902,N_9498);
xnor U11635 (N_11635,N_9592,N_6399);
and U11636 (N_11636,N_7984,N_9534);
and U11637 (N_11637,N_5729,N_7618);
nand U11638 (N_11638,N_6140,N_9123);
nand U11639 (N_11639,N_7064,N_5939);
nand U11640 (N_11640,N_5773,N_9954);
and U11641 (N_11641,N_8258,N_8941);
and U11642 (N_11642,N_9286,N_9111);
nor U11643 (N_11643,N_8772,N_9493);
or U11644 (N_11644,N_7850,N_8216);
xor U11645 (N_11645,N_7468,N_8156);
and U11646 (N_11646,N_8877,N_8624);
and U11647 (N_11647,N_8511,N_8947);
or U11648 (N_11648,N_5992,N_5986);
and U11649 (N_11649,N_8925,N_8043);
or U11650 (N_11650,N_7427,N_5518);
xor U11651 (N_11651,N_8047,N_9514);
nor U11652 (N_11652,N_6927,N_9241);
or U11653 (N_11653,N_8646,N_8206);
or U11654 (N_11654,N_9872,N_5281);
and U11655 (N_11655,N_8605,N_6819);
xnor U11656 (N_11656,N_7307,N_7894);
or U11657 (N_11657,N_5604,N_6490);
nor U11658 (N_11658,N_5702,N_6825);
and U11659 (N_11659,N_7647,N_5285);
nor U11660 (N_11660,N_9331,N_6389);
and U11661 (N_11661,N_5259,N_5568);
nor U11662 (N_11662,N_7864,N_5893);
nand U11663 (N_11663,N_5653,N_6055);
and U11664 (N_11664,N_7018,N_8129);
nor U11665 (N_11665,N_7896,N_7482);
nand U11666 (N_11666,N_7625,N_7857);
nand U11667 (N_11667,N_9388,N_7396);
nor U11668 (N_11668,N_8663,N_8086);
and U11669 (N_11669,N_6754,N_7658);
and U11670 (N_11670,N_9328,N_9655);
and U11671 (N_11671,N_8705,N_9138);
or U11672 (N_11672,N_5131,N_6117);
nand U11673 (N_11673,N_8175,N_5657);
nand U11674 (N_11674,N_6093,N_5092);
or U11675 (N_11675,N_7971,N_5081);
nor U11676 (N_11676,N_8017,N_9737);
nand U11677 (N_11677,N_7135,N_9565);
xnor U11678 (N_11678,N_8371,N_5366);
nand U11679 (N_11679,N_8470,N_7906);
nand U11680 (N_11680,N_6410,N_8992);
nand U11681 (N_11681,N_6052,N_6534);
nor U11682 (N_11682,N_8252,N_7152);
nand U11683 (N_11683,N_7407,N_5377);
nand U11684 (N_11684,N_5969,N_7776);
or U11685 (N_11685,N_7495,N_6650);
nor U11686 (N_11686,N_8898,N_5327);
nor U11687 (N_11687,N_6373,N_9897);
nor U11688 (N_11688,N_9213,N_6166);
or U11689 (N_11689,N_5119,N_9536);
nand U11690 (N_11690,N_5430,N_8546);
nor U11691 (N_11691,N_6200,N_7295);
and U11692 (N_11692,N_8458,N_7409);
xor U11693 (N_11693,N_8137,N_6261);
nand U11694 (N_11694,N_8879,N_8888);
nand U11695 (N_11695,N_9338,N_5315);
xor U11696 (N_11696,N_9381,N_8942);
nor U11697 (N_11697,N_8934,N_6450);
nor U11698 (N_11698,N_5527,N_6381);
nand U11699 (N_11699,N_8749,N_6453);
and U11700 (N_11700,N_5907,N_5607);
xor U11701 (N_11701,N_9633,N_6766);
nor U11702 (N_11702,N_9833,N_9998);
or U11703 (N_11703,N_7865,N_5575);
or U11704 (N_11704,N_9696,N_5569);
or U11705 (N_11705,N_9253,N_7446);
or U11706 (N_11706,N_8999,N_7467);
xnor U11707 (N_11707,N_5129,N_7184);
or U11708 (N_11708,N_7368,N_5966);
and U11709 (N_11709,N_5167,N_8153);
or U11710 (N_11710,N_6542,N_8547);
or U11711 (N_11711,N_9640,N_9600);
xor U11712 (N_11712,N_5411,N_7089);
nor U11713 (N_11713,N_8560,N_9947);
and U11714 (N_11714,N_6959,N_8109);
and U11715 (N_11715,N_7097,N_7312);
and U11716 (N_11716,N_5925,N_8841);
and U11717 (N_11717,N_8519,N_8358);
nand U11718 (N_11718,N_8631,N_5953);
nor U11719 (N_11719,N_7102,N_6829);
nand U11720 (N_11720,N_9744,N_7889);
or U11721 (N_11721,N_6156,N_9641);
nand U11722 (N_11722,N_7780,N_8082);
nor U11723 (N_11723,N_5780,N_6491);
or U11724 (N_11724,N_5175,N_7344);
or U11725 (N_11725,N_7432,N_8152);
and U11726 (N_11726,N_8857,N_9282);
and U11727 (N_11727,N_6823,N_6822);
or U11728 (N_11728,N_7124,N_9348);
xnor U11729 (N_11729,N_9175,N_8562);
or U11730 (N_11730,N_6948,N_6472);
nand U11731 (N_11731,N_6186,N_6696);
or U11732 (N_11732,N_7818,N_5764);
or U11733 (N_11733,N_5199,N_5996);
or U11734 (N_11734,N_7055,N_5693);
nand U11735 (N_11735,N_7270,N_5425);
nor U11736 (N_11736,N_6519,N_5367);
xor U11737 (N_11737,N_7709,N_7149);
and U11738 (N_11738,N_5485,N_5426);
xor U11739 (N_11739,N_6318,N_6799);
or U11740 (N_11740,N_7886,N_8294);
and U11741 (N_11741,N_9264,N_5514);
and U11742 (N_11742,N_8214,N_7990);
or U11743 (N_11743,N_7587,N_9015);
or U11744 (N_11744,N_6080,N_6096);
and U11745 (N_11745,N_7469,N_9108);
nand U11746 (N_11746,N_9802,N_8959);
nand U11747 (N_11747,N_8202,N_6858);
nor U11748 (N_11748,N_5565,N_8591);
nand U11749 (N_11749,N_5306,N_9361);
xor U11750 (N_11750,N_8767,N_7397);
or U11751 (N_11751,N_5305,N_9736);
xor U11752 (N_11752,N_6264,N_8256);
or U11753 (N_11753,N_8368,N_7544);
or U11754 (N_11754,N_7922,N_7379);
or U11755 (N_11755,N_8962,N_9811);
or U11756 (N_11756,N_6502,N_5749);
nor U11757 (N_11757,N_5943,N_7069);
nand U11758 (N_11758,N_6661,N_7547);
and U11759 (N_11759,N_9798,N_6300);
xor U11760 (N_11760,N_7741,N_6883);
nand U11761 (N_11761,N_5128,N_5438);
nand U11762 (N_11762,N_7006,N_9502);
or U11763 (N_11763,N_8773,N_5936);
nor U11764 (N_11764,N_9206,N_9378);
or U11765 (N_11765,N_7548,N_8997);
or U11766 (N_11766,N_8794,N_5010);
or U11767 (N_11767,N_9662,N_8422);
nand U11768 (N_11768,N_5892,N_7297);
nand U11769 (N_11769,N_6125,N_5138);
and U11770 (N_11770,N_6225,N_9923);
or U11771 (N_11771,N_9217,N_7822);
nand U11772 (N_11772,N_5172,N_8283);
xor U11773 (N_11773,N_5952,N_9329);
and U11774 (N_11774,N_7433,N_6993);
or U11775 (N_11775,N_6694,N_6958);
nand U11776 (N_11776,N_6657,N_5983);
or U11777 (N_11777,N_9530,N_9096);
nor U11778 (N_11778,N_5837,N_8243);
nor U11779 (N_11779,N_7441,N_9899);
or U11780 (N_11780,N_9799,N_6710);
nand U11781 (N_11781,N_9642,N_7938);
nor U11782 (N_11782,N_8464,N_8639);
nor U11783 (N_11783,N_9212,N_6738);
nor U11784 (N_11784,N_6813,N_6695);
nor U11785 (N_11785,N_5477,N_9804);
or U11786 (N_11786,N_8536,N_6730);
nor U11787 (N_11787,N_8853,N_6862);
xor U11788 (N_11788,N_8640,N_5543);
or U11789 (N_11789,N_6662,N_9346);
and U11790 (N_11790,N_7836,N_9894);
nor U11791 (N_11791,N_9569,N_8851);
xor U11792 (N_11792,N_6842,N_7657);
and U11793 (N_11793,N_7726,N_8097);
xnor U11794 (N_11794,N_8490,N_6509);
and U11795 (N_11795,N_7847,N_9461);
xnor U11796 (N_11796,N_6577,N_6853);
nor U11797 (N_11797,N_9085,N_8634);
nor U11798 (N_11798,N_5395,N_7176);
or U11799 (N_11799,N_5915,N_8953);
and U11800 (N_11800,N_7074,N_8507);
and U11801 (N_11801,N_7403,N_7786);
nor U11802 (N_11802,N_6773,N_7508);
and U11803 (N_11803,N_8372,N_5036);
and U11804 (N_11804,N_9142,N_5323);
or U11805 (N_11805,N_6917,N_6035);
or U11806 (N_11806,N_7346,N_7047);
and U11807 (N_11807,N_7052,N_9856);
or U11808 (N_11808,N_8593,N_7719);
and U11809 (N_11809,N_8845,N_7926);
or U11810 (N_11810,N_6267,N_8629);
or U11811 (N_11811,N_6262,N_7226);
nand U11812 (N_11812,N_8885,N_7484);
nand U11813 (N_11813,N_7196,N_5356);
or U11814 (N_11814,N_6209,N_6715);
and U11815 (N_11815,N_6743,N_6667);
or U11816 (N_11816,N_5960,N_5071);
nor U11817 (N_11817,N_7528,N_8317);
xor U11818 (N_11818,N_7013,N_8193);
nor U11819 (N_11819,N_8224,N_7720);
nand U11820 (N_11820,N_6956,N_7691);
or U11821 (N_11821,N_8058,N_8955);
nor U11822 (N_11822,N_5031,N_9060);
nand U11823 (N_11823,N_7673,N_8957);
nor U11824 (N_11824,N_9185,N_8313);
xor U11825 (N_11825,N_8809,N_7197);
nor U11826 (N_11826,N_9591,N_5541);
xnor U11827 (N_11827,N_6008,N_9747);
nor U11828 (N_11828,N_9939,N_7619);
nand U11829 (N_11829,N_7214,N_5257);
xor U11830 (N_11830,N_6386,N_5753);
and U11831 (N_11831,N_9568,N_6761);
nor U11832 (N_11832,N_7791,N_9390);
nor U11833 (N_11833,N_8886,N_6798);
nor U11834 (N_11834,N_6977,N_9347);
and U11835 (N_11835,N_9236,N_6254);
nor U11836 (N_11836,N_8339,N_7790);
nor U11837 (N_11837,N_6382,N_7171);
nand U11838 (N_11838,N_5087,N_8861);
and U11839 (N_11839,N_9905,N_8545);
or U11840 (N_11840,N_5418,N_6558);
xnor U11841 (N_11841,N_6174,N_7637);
xor U11842 (N_11842,N_9858,N_8670);
nor U11843 (N_11843,N_9732,N_9228);
and U11844 (N_11844,N_7262,N_9369);
or U11845 (N_11845,N_5289,N_6805);
nor U11846 (N_11846,N_7323,N_8104);
or U11847 (N_11847,N_9960,N_5341);
or U11848 (N_11848,N_5590,N_8674);
nor U11849 (N_11849,N_9559,N_5316);
and U11850 (N_11850,N_8825,N_9384);
and U11851 (N_11851,N_8823,N_5635);
and U11852 (N_11852,N_8293,N_5908);
or U11853 (N_11853,N_7456,N_6324);
nand U11854 (N_11854,N_6518,N_5263);
or U11855 (N_11855,N_7367,N_6210);
xnor U11856 (N_11856,N_7595,N_8032);
or U11857 (N_11857,N_5415,N_9284);
xor U11858 (N_11858,N_9567,N_6336);
xnor U11859 (N_11859,N_7436,N_5870);
xor U11860 (N_11860,N_5043,N_5561);
nand U11861 (N_11861,N_8122,N_7626);
and U11862 (N_11862,N_9114,N_6219);
nor U11863 (N_11863,N_7806,N_7952);
or U11864 (N_11864,N_7037,N_5760);
nor U11865 (N_11865,N_8365,N_7193);
xnor U11866 (N_11866,N_7039,N_8621);
xor U11867 (N_11867,N_7034,N_7324);
xnor U11868 (N_11868,N_6376,N_7398);
and U11869 (N_11869,N_5822,N_6827);
and U11870 (N_11870,N_9827,N_8119);
xnor U11871 (N_11871,N_8890,N_6788);
nor U11872 (N_11872,N_5494,N_9627);
and U11873 (N_11873,N_9349,N_9062);
nor U11874 (N_11874,N_9866,N_6864);
and U11875 (N_11875,N_6867,N_9748);
nor U11876 (N_11876,N_6390,N_8848);
or U11877 (N_11877,N_7609,N_6596);
or U11878 (N_11878,N_5757,N_9159);
and U11879 (N_11879,N_8768,N_6378);
nor U11880 (N_11880,N_7887,N_7531);
or U11881 (N_11881,N_5555,N_9529);
and U11882 (N_11882,N_8356,N_9342);
or U11883 (N_11883,N_5545,N_9011);
and U11884 (N_11884,N_6297,N_7106);
nor U11885 (N_11885,N_6834,N_8185);
nor U11886 (N_11886,N_8023,N_8318);
nand U11887 (N_11887,N_6295,N_5533);
or U11888 (N_11888,N_7228,N_7699);
and U11889 (N_11889,N_5173,N_9045);
nand U11890 (N_11890,N_8622,N_6685);
nor U11891 (N_11891,N_6001,N_8958);
or U11892 (N_11892,N_8503,N_9540);
or U11893 (N_11893,N_6896,N_8398);
or U11894 (N_11894,N_6486,N_7103);
nor U11895 (N_11895,N_7879,N_5586);
nor U11896 (N_11896,N_6251,N_8174);
nor U11897 (N_11897,N_7279,N_6040);
nand U11898 (N_11898,N_5413,N_7750);
nor U11899 (N_11899,N_6974,N_9232);
or U11900 (N_11900,N_8051,N_6516);
or U11901 (N_11901,N_7167,N_9481);
or U11902 (N_11902,N_5894,N_7377);
nand U11903 (N_11903,N_7066,N_7775);
nand U11904 (N_11904,N_5685,N_5481);
nand U11905 (N_11905,N_8875,N_5310);
and U11906 (N_11906,N_5307,N_7642);
nor U11907 (N_11907,N_8071,N_9458);
nor U11908 (N_11908,N_9221,N_9546);
nand U11909 (N_11909,N_9009,N_8781);
nor U11910 (N_11910,N_8098,N_8033);
nand U11911 (N_11911,N_6550,N_5709);
and U11912 (N_11912,N_8508,N_8103);
nor U11913 (N_11913,N_7122,N_5828);
and U11914 (N_11914,N_6670,N_8632);
nor U11915 (N_11915,N_7939,N_9694);
and U11916 (N_11916,N_5622,N_8100);
or U11917 (N_11917,N_8321,N_7759);
and U11918 (N_11918,N_6536,N_7893);
or U11919 (N_11919,N_9256,N_9456);
nand U11920 (N_11920,N_8387,N_8708);
nand U11921 (N_11921,N_9460,N_7282);
nand U11922 (N_11922,N_7202,N_7634);
nand U11923 (N_11923,N_9063,N_6029);
nand U11924 (N_11924,N_8596,N_6031);
nand U11925 (N_11925,N_5370,N_7383);
nand U11926 (N_11926,N_8881,N_7559);
nor U11927 (N_11927,N_6493,N_6716);
and U11928 (N_11928,N_5317,N_9402);
or U11929 (N_11929,N_5808,N_5374);
xnor U11930 (N_11930,N_8716,N_9215);
xor U11931 (N_11931,N_6523,N_7987);
and U11932 (N_11932,N_9705,N_6680);
nand U11933 (N_11933,N_6705,N_9080);
xor U11934 (N_11934,N_5534,N_9809);
nor U11935 (N_11935,N_6427,N_6935);
nor U11936 (N_11936,N_9670,N_9760);
nand U11937 (N_11937,N_8822,N_5551);
and U11938 (N_11938,N_9847,N_5840);
nor U11939 (N_11939,N_9043,N_6423);
nand U11940 (N_11940,N_5516,N_9229);
nand U11941 (N_11941,N_7663,N_6852);
nand U11942 (N_11942,N_6624,N_8115);
and U11943 (N_11943,N_7272,N_8013);
nand U11944 (N_11944,N_8764,N_5660);
and U11945 (N_11945,N_9339,N_7909);
and U11946 (N_11946,N_9772,N_6859);
or U11947 (N_11947,N_5144,N_6457);
or U11948 (N_11948,N_5546,N_9727);
or U11949 (N_11949,N_5998,N_9163);
nor U11950 (N_11950,N_6592,N_7996);
nand U11951 (N_11951,N_5522,N_7340);
nor U11952 (N_11952,N_8089,N_6630);
nand U11953 (N_11953,N_6775,N_9164);
or U11954 (N_11954,N_5136,N_8421);
or U11955 (N_11955,N_9365,N_5158);
or U11956 (N_11956,N_8635,N_9194);
or U11957 (N_11957,N_8418,N_7429);
xor U11958 (N_11958,N_9183,N_9289);
xnor U11959 (N_11959,N_6414,N_5419);
and U11960 (N_11960,N_5210,N_5201);
nand U11961 (N_11961,N_6875,N_5180);
and U11962 (N_11962,N_9832,N_8835);
nor U11963 (N_11963,N_6877,N_7702);
or U11964 (N_11964,N_7450,N_7030);
nand U11965 (N_11965,N_8981,N_7725);
and U11966 (N_11966,N_8044,N_7083);
and U11967 (N_11967,N_5459,N_8320);
and U11968 (N_11968,N_5584,N_8233);
nand U11969 (N_11969,N_5074,N_9570);
or U11970 (N_11970,N_6950,N_9871);
and U11971 (N_11971,N_6533,N_9986);
or U11972 (N_11972,N_6207,N_8984);
nor U11973 (N_11973,N_7689,N_5113);
nand U11974 (N_11974,N_9079,N_7281);
nor U11975 (N_11975,N_9638,N_5488);
nand U11976 (N_11976,N_8813,N_9141);
and U11977 (N_11977,N_9022,N_7125);
nor U11978 (N_11978,N_5552,N_5674);
xor U11979 (N_11979,N_9042,N_5835);
or U11980 (N_11980,N_9409,N_7789);
and U11981 (N_11981,N_8453,N_6185);
xnor U11982 (N_11982,N_8160,N_7610);
xor U11983 (N_11983,N_6356,N_6359);
nand U11984 (N_11984,N_5762,N_5827);
nand U11985 (N_11985,N_5576,N_6996);
nor U11986 (N_11986,N_5440,N_6778);
xnor U11987 (N_11987,N_6294,N_8066);
and U11988 (N_11988,N_6056,N_9091);
nand U11989 (N_11989,N_7739,N_7516);
or U11990 (N_11990,N_5889,N_6865);
and U11991 (N_11991,N_5298,N_8052);
xor U11992 (N_11992,N_5185,N_6525);
xnor U11993 (N_11993,N_5928,N_9969);
nand U11994 (N_11994,N_5594,N_5955);
or U11995 (N_11995,N_9061,N_7514);
and U11996 (N_11996,N_6848,N_8528);
or U11997 (N_11997,N_5985,N_8236);
and U11998 (N_11998,N_9491,N_7638);
xnor U11999 (N_11999,N_5107,N_6161);
nor U12000 (N_12000,N_5759,N_5968);
and U12001 (N_12001,N_5817,N_6353);
or U12002 (N_12002,N_8282,N_8426);
and U12003 (N_12003,N_9796,N_7209);
or U12004 (N_12004,N_8142,N_5699);
nand U12005 (N_12005,N_9814,N_7897);
and U12006 (N_12006,N_8615,N_5946);
nor U12007 (N_12007,N_5833,N_6038);
nand U12008 (N_12008,N_6871,N_8793);
and U12009 (N_12009,N_9492,N_5821);
and U12010 (N_12010,N_6537,N_9374);
or U12011 (N_12011,N_7236,N_6277);
or U12012 (N_12012,N_7570,N_6789);
and U12013 (N_12013,N_9283,N_8388);
and U12014 (N_12014,N_9326,N_6539);
and U12015 (N_12015,N_5517,N_8476);
nor U12016 (N_12016,N_5373,N_5274);
and U12017 (N_12017,N_8307,N_5632);
and U12018 (N_12018,N_7539,N_7958);
and U12019 (N_12019,N_8680,N_7173);
nand U12020 (N_12020,N_6580,N_7502);
nor U12021 (N_12021,N_6992,N_5145);
and U12022 (N_12022,N_5150,N_6731);
nand U12023 (N_12023,N_8750,N_8375);
and U12024 (N_12024,N_8136,N_6224);
and U12025 (N_12025,N_6540,N_8998);
or U12026 (N_12026,N_7742,N_5227);
xor U12027 (N_12027,N_6702,N_5384);
nand U12028 (N_12028,N_8765,N_5216);
and U12029 (N_12029,N_9517,N_6216);
nor U12030 (N_12030,N_9542,N_6514);
nor U12031 (N_12031,N_5776,N_6245);
nor U12032 (N_12032,N_9441,N_5678);
nor U12033 (N_12033,N_8604,N_6767);
or U12034 (N_12034,N_7620,N_9377);
or U12035 (N_12035,N_5853,N_5503);
nor U12036 (N_12036,N_5688,N_7600);
and U12037 (N_12037,N_5710,N_5623);
and U12038 (N_12038,N_8920,N_8124);
and U12039 (N_12039,N_7731,N_9246);
nor U12040 (N_12040,N_7161,N_5703);
or U12041 (N_12041,N_8923,N_9249);
nor U12042 (N_12042,N_5784,N_9449);
or U12043 (N_12043,N_6184,N_9489);
nor U12044 (N_12044,N_6432,N_7293);
nand U12045 (N_12045,N_5715,N_6452);
nand U12046 (N_12046,N_6176,N_6287);
nand U12047 (N_12047,N_6511,N_8618);
and U12048 (N_12048,N_9617,N_9993);
nand U12049 (N_12049,N_7380,N_9125);
and U12050 (N_12050,N_9041,N_6623);
or U12051 (N_12051,N_5599,N_8488);
nand U12052 (N_12052,N_5990,N_5282);
nand U12053 (N_12053,N_7222,N_9769);
nand U12054 (N_12054,N_8134,N_9355);
nand U12055 (N_12055,N_5239,N_8213);
and U12056 (N_12056,N_5251,N_8462);
nand U12057 (N_12057,N_8485,N_5017);
or U12058 (N_12058,N_6940,N_8701);
nor U12059 (N_12059,N_7164,N_8723);
or U12060 (N_12060,N_8212,N_8530);
nor U12061 (N_12061,N_9363,N_5805);
nor U12062 (N_12062,N_7128,N_7555);
nor U12063 (N_12063,N_6617,N_7342);
or U12064 (N_12064,N_7831,N_6938);
nand U12065 (N_12065,N_6483,N_7035);
nand U12066 (N_12066,N_6436,N_8961);
nor U12067 (N_12067,N_8349,N_8828);
nor U12068 (N_12068,N_9587,N_6433);
or U12069 (N_12069,N_7205,N_6648);
and U12070 (N_12070,N_7947,N_5496);
nor U12071 (N_12071,N_5706,N_9949);
nor U12072 (N_12072,N_8964,N_7218);
and U12073 (N_12073,N_6686,N_7402);
nand U12074 (N_12074,N_5082,N_7426);
nor U12075 (N_12075,N_5615,N_7573);
and U12076 (N_12076,N_8846,N_5099);
nand U12077 (N_12077,N_8517,N_9197);
nand U12078 (N_12078,N_9563,N_9299);
nand U12079 (N_12079,N_8215,N_8477);
and U12080 (N_12080,N_9398,N_7814);
nor U12081 (N_12081,N_6611,N_8818);
or U12082 (N_12082,N_9803,N_9777);
nor U12083 (N_12083,N_6810,N_5585);
nor U12084 (N_12084,N_8177,N_7898);
xnor U12085 (N_12085,N_7442,N_9860);
nor U12086 (N_12086,N_7643,N_5364);
nor U12087 (N_12087,N_5732,N_9423);
nand U12088 (N_12088,N_6809,N_7043);
and U12089 (N_12089,N_9003,N_7109);
and U12090 (N_12090,N_8257,N_5141);
nor U12091 (N_12091,N_7740,N_7923);
nor U12092 (N_12092,N_5350,N_9273);
nand U12093 (N_12093,N_8601,N_5995);
nor U12094 (N_12094,N_7415,N_8222);
nor U12095 (N_12095,N_7071,N_9028);
and U12096 (N_12096,N_9101,N_9509);
xnor U12097 (N_12097,N_9327,N_6221);
nor U12098 (N_12098,N_6227,N_7470);
and U12099 (N_12099,N_6522,N_8741);
and U12100 (N_12100,N_7648,N_8529);
nor U12101 (N_12101,N_8983,N_7527);
nor U12102 (N_12102,N_7810,N_5178);
nor U12103 (N_12103,N_6460,N_7766);
and U12104 (N_12104,N_9929,N_8899);
nand U12105 (N_12105,N_7424,N_6594);
nor U12106 (N_12106,N_7722,N_5218);
and U12107 (N_12107,N_5901,N_9373);
and U12108 (N_12108,N_9376,N_9248);
xnor U12109 (N_12109,N_7119,N_6372);
and U12110 (N_12110,N_6042,N_9668);
and U12111 (N_12111,N_6360,N_9794);
nand U12112 (N_12112,N_7955,N_8867);
and U12113 (N_12113,N_7842,N_6235);
xnor U12114 (N_12114,N_7406,N_8312);
and U12115 (N_12115,N_9978,N_6981);
nand U12116 (N_12116,N_5137,N_5393);
xor U12117 (N_12117,N_5802,N_9789);
or U12118 (N_12118,N_7522,N_7665);
or U12119 (N_12119,N_7830,N_8729);
nand U12120 (N_12120,N_8102,N_5471);
xor U12121 (N_12121,N_6146,N_8383);
and U12122 (N_12122,N_8965,N_8067);
nor U12123 (N_12123,N_9058,N_9504);
or U12124 (N_12124,N_8587,N_5638);
xor U12125 (N_12125,N_6292,N_7221);
or U12126 (N_12126,N_7126,N_5644);
or U12127 (N_12127,N_9618,N_7359);
nand U12128 (N_12128,N_5899,N_8393);
nand U12129 (N_12129,N_9720,N_6583);
nor U12130 (N_12130,N_6248,N_5974);
nor U12131 (N_12131,N_5920,N_8832);
nor U12132 (N_12132,N_8738,N_8138);
and U12133 (N_12133,N_8326,N_6892);
nand U12134 (N_12134,N_9242,N_9443);
nor U12135 (N_12135,N_5358,N_8163);
nor U12136 (N_12136,N_7985,N_8731);
xnor U12137 (N_12137,N_9117,N_6807);
nand U12138 (N_12138,N_6882,N_7566);
nor U12139 (N_12139,N_6032,N_9665);
xnor U12140 (N_12140,N_9522,N_6554);
and U12141 (N_12141,N_6651,N_9942);
nand U12142 (N_12142,N_5656,N_8072);
and U12143 (N_12143,N_8917,N_7192);
nor U12144 (N_12144,N_7978,N_8804);
nand U12145 (N_12145,N_6475,N_7771);
or U12146 (N_12146,N_7474,N_5593);
nor U12147 (N_12147,N_6163,N_6794);
nor U12148 (N_12148,N_8652,N_5396);
and U12149 (N_12149,N_7355,N_5429);
or U12150 (N_12150,N_5880,N_9475);
xnor U12151 (N_12151,N_5379,N_9429);
nor U12152 (N_12152,N_5797,N_8188);
or U12153 (N_12153,N_7313,N_9140);
or U12154 (N_12154,N_6995,N_8746);
nor U12155 (N_12155,N_6820,N_5523);
nand U12156 (N_12156,N_5111,N_7168);
nor U12157 (N_12157,N_6345,N_5971);
and U12158 (N_12158,N_8667,N_7538);
or U12159 (N_12159,N_8260,N_9270);
and U12160 (N_12160,N_5994,N_9451);
xnor U12161 (N_12161,N_8012,N_5056);
and U12162 (N_12162,N_7703,N_5402);
xnor U12163 (N_12163,N_7688,N_9054);
nand U12164 (N_12164,N_8255,N_7783);
nor U12165 (N_12165,N_9323,N_7802);
nand U12166 (N_12166,N_5613,N_8676);
nand U12167 (N_12167,N_8231,N_9001);
and U12168 (N_12168,N_8876,N_6904);
or U12169 (N_12169,N_6856,N_6910);
nor U12170 (N_12170,N_9083,N_6527);
and U12171 (N_12171,N_5476,N_9630);
or U12172 (N_12172,N_5058,N_5066);
nor U12173 (N_12173,N_7153,N_9044);
or U12174 (N_12174,N_8918,N_8915);
and U12175 (N_12175,N_7478,N_6639);
and U12176 (N_12176,N_9651,N_6191);
nor U12177 (N_12177,N_7653,N_6124);
nand U12178 (N_12178,N_8771,N_8042);
nand U12179 (N_12179,N_8131,N_9463);
and U12180 (N_12180,N_9235,N_6975);
nand U12181 (N_12181,N_8074,N_5935);
and U12182 (N_12182,N_5814,N_6672);
nor U12183 (N_12183,N_9780,N_7157);
nor U12184 (N_12184,N_8524,N_8397);
nand U12185 (N_12185,N_7249,N_6930);
nor U12186 (N_12186,N_7303,N_9087);
or U12187 (N_12187,N_5826,N_6152);
or U12188 (N_12188,N_8405,N_8106);
nor U12189 (N_12189,N_7356,N_7799);
and U12190 (N_12190,N_6455,N_9350);
or U12191 (N_12191,N_8386,N_8278);
and U12192 (N_12192,N_8718,N_9483);
and U12193 (N_12193,N_6782,N_6625);
and U12194 (N_12194,N_8494,N_8745);
nor U12195 (N_12195,N_7574,N_8988);
nand U12196 (N_12196,N_7143,N_6240);
xor U12197 (N_12197,N_9637,N_5504);
xor U12198 (N_12198,N_8976,N_9392);
xor U12199 (N_12199,N_7807,N_9031);
or U12200 (N_12200,N_5231,N_9740);
or U12201 (N_12201,N_8331,N_5206);
nand U12202 (N_12202,N_8769,N_9984);
or U12203 (N_12203,N_7244,N_5667);
nor U12204 (N_12204,N_6919,N_7596);
or U12205 (N_12205,N_8434,N_8544);
and U12206 (N_12206,N_8700,N_5963);
and U12207 (N_12207,N_7885,N_8696);
or U12208 (N_12208,N_9578,N_6232);
or U12209 (N_12209,N_6092,N_6431);
and U12210 (N_12210,N_5098,N_6647);
nor U12211 (N_12211,N_8475,N_5639);
or U12212 (N_12212,N_5818,N_6627);
and U12213 (N_12213,N_6079,N_8217);
nor U12214 (N_12214,N_6559,N_9646);
and U12215 (N_12215,N_7250,N_6304);
xnor U12216 (N_12216,N_8776,N_9425);
nor U12217 (N_12217,N_6257,N_6899);
nand U12218 (N_12218,N_9434,N_5085);
nand U12219 (N_12219,N_9979,N_9882);
nor U12220 (N_12220,N_6437,N_9057);
or U12221 (N_12221,N_8510,N_6441);
or U12222 (N_12222,N_7929,N_6895);
nand U12223 (N_12223,N_9018,N_9049);
xnor U12224 (N_12224,N_6203,N_6839);
nand U12225 (N_12225,N_7073,N_9626);
xor U12226 (N_12226,N_9580,N_7685);
nand U12227 (N_12227,N_7016,N_6193);
nor U12228 (N_12228,N_7382,N_6307);
nand U12229 (N_12229,N_9785,N_5662);
nor U12230 (N_12230,N_8445,N_6602);
nor U12231 (N_12231,N_8227,N_8806);
nand U12232 (N_12232,N_5886,N_6733);
nor U12233 (N_12233,N_5991,N_9527);
nand U12234 (N_12234,N_7180,N_5400);
nor U12235 (N_12235,N_9895,N_7491);
nand U12236 (N_12236,N_9884,N_9661);
or U12237 (N_12237,N_7542,N_5152);
nor U12238 (N_12238,N_6573,N_7669);
xnor U12239 (N_12239,N_9296,N_9752);
or U12240 (N_12240,N_8267,N_8169);
nor U12241 (N_12241,N_7003,N_6943);
nand U12242 (N_12242,N_7348,N_5187);
or U12243 (N_12243,N_5325,N_7593);
and U12244 (N_12244,N_5976,N_8799);
xor U12245 (N_12245,N_6590,N_5683);
nand U12246 (N_12246,N_6632,N_9225);
and U12247 (N_12247,N_9336,N_8754);
nand U12248 (N_12248,N_6804,N_6806);
nor U12249 (N_12249,N_9552,N_8633);
and U12250 (N_12250,N_8360,N_7976);
and U12251 (N_12251,N_9865,N_5241);
or U12252 (N_12252,N_5999,N_5461);
or U12253 (N_12253,N_9885,N_5927);
nand U12254 (N_12254,N_9707,N_6677);
or U12255 (N_12255,N_8944,N_5547);
and U12256 (N_12256,N_7113,N_9278);
and U12257 (N_12257,N_8493,N_9940);
or U12258 (N_12258,N_8165,N_8410);
and U12259 (N_12259,N_5917,N_9039);
nand U12260 (N_12260,N_6053,N_6551);
and U12261 (N_12261,N_5195,N_6404);
and U12262 (N_12262,N_7187,N_5155);
and U12263 (N_12263,N_7301,N_8391);
and U12264 (N_12264,N_9023,N_7389);
nand U12265 (N_12265,N_5246,N_7770);
or U12266 (N_12266,N_7336,N_6921);
nand U12267 (N_12267,N_6362,N_8413);
or U12268 (N_12268,N_7150,N_9147);
nand U12269 (N_12269,N_8305,N_5021);
nor U12270 (N_12270,N_8253,N_7290);
nor U12271 (N_12271,N_9843,N_5186);
nor U12272 (N_12272,N_8292,N_6656);
xor U12273 (N_12273,N_8404,N_5723);
or U12274 (N_12274,N_9750,N_9991);
or U12275 (N_12275,N_5139,N_8110);
nand U12276 (N_12276,N_8717,N_5502);
nor U12277 (N_12277,N_9790,N_9729);
and U12278 (N_12278,N_9826,N_7846);
nor U12279 (N_12279,N_7190,N_8037);
or U12280 (N_12280,N_9919,N_7687);
or U12281 (N_12281,N_6007,N_8125);
or U12282 (N_12282,N_7981,N_9597);
or U12283 (N_12283,N_7670,N_6274);
nor U12284 (N_12284,N_9008,N_8064);
nor U12285 (N_12285,N_9403,N_9582);
nand U12286 (N_12286,N_9334,N_8525);
nand U12287 (N_12287,N_8854,N_6312);
nand U12288 (N_12288,N_5885,N_8919);
nor U12289 (N_12289,N_9077,N_6077);
nand U12290 (N_12290,N_5548,N_7465);
and U12291 (N_12291,N_6476,N_7763);
or U12292 (N_12292,N_7612,N_5863);
and U12293 (N_12293,N_8543,N_8820);
or U12294 (N_12294,N_7284,N_8610);
or U12295 (N_12295,N_6803,N_6357);
xnor U12296 (N_12296,N_6101,N_9306);
and U12297 (N_12297,N_9693,N_9203);
nand U12298 (N_12298,N_6659,N_8687);
nand U12299 (N_12299,N_5009,N_5510);
nand U12300 (N_12300,N_7111,N_9293);
nand U12301 (N_12301,N_7515,N_9912);
xor U12302 (N_12302,N_8501,N_9222);
or U12303 (N_12303,N_9448,N_9170);
nand U12304 (N_12304,N_7915,N_6002);
nand U12305 (N_12305,N_5973,N_6846);
nor U12306 (N_12306,N_9290,N_9471);
or U12307 (N_12307,N_7081,N_6228);
and U12308 (N_12308,N_7900,N_5620);
or U12309 (N_12309,N_5823,N_5934);
or U12310 (N_12310,N_7007,N_8819);
nor U12311 (N_12311,N_6281,N_9116);
and U12312 (N_12312,N_7917,N_8571);
nand U12313 (N_12313,N_6957,N_5666);
nor U12314 (N_12314,N_7485,N_9624);
nor U12315 (N_12315,N_9631,N_9664);
or U12316 (N_12316,N_6223,N_5842);
nor U12317 (N_12317,N_9690,N_9380);
and U12318 (N_12318,N_5062,N_8338);
and U12319 (N_12319,N_9161,N_5871);
and U12320 (N_12320,N_7521,N_9951);
xor U12321 (N_12321,N_5803,N_9064);
nor U12322 (N_12322,N_6732,N_7704);
or U12323 (N_12323,N_8908,N_8083);
nor U12324 (N_12324,N_6870,N_5767);
nand U12325 (N_12325,N_5932,N_8112);
or U12326 (N_12326,N_6765,N_6150);
nor U12327 (N_12327,N_7299,N_8497);
xor U12328 (N_12328,N_8567,N_7644);
nor U12329 (N_12329,N_9220,N_7655);
and U12330 (N_12330,N_5196,N_8330);
xnor U12331 (N_12331,N_8760,N_6631);
nor U12332 (N_12332,N_5334,N_7044);
nor U12333 (N_12333,N_8436,N_5386);
xnor U12334 (N_12334,N_9697,N_5676);
nor U12335 (N_12335,N_8780,N_6538);
nand U12336 (N_12336,N_6116,N_9325);
and U12337 (N_12337,N_5745,N_8909);
xnor U12338 (N_12338,N_5498,N_8172);
xor U12339 (N_12339,N_5798,N_5897);
nand U12340 (N_12340,N_6263,N_9026);
nor U12341 (N_12341,N_5896,N_5450);
nor U12342 (N_12342,N_7201,N_6387);
xnor U12343 (N_12343,N_7033,N_5319);
and U12344 (N_12344,N_8786,N_7123);
nand U12345 (N_12345,N_6448,N_8570);
nand U12346 (N_12346,N_9652,N_9795);
or U12347 (N_12347,N_9973,N_5270);
and U12348 (N_12348,N_7962,N_9503);
nand U12349 (N_12349,N_5202,N_9948);
xor U12350 (N_12350,N_7793,N_8950);
nor U12351 (N_12351,N_7734,N_6653);
and U12352 (N_12352,N_5905,N_9106);
xnor U12353 (N_12353,N_9962,N_8728);
xor U12354 (N_12354,N_9751,N_9128);
or U12355 (N_12355,N_5625,N_8150);
nand U12356 (N_12356,N_7031,N_5804);
nand U12357 (N_12357,N_5151,N_9112);
and U12358 (N_12358,N_7101,N_9113);
nand U12359 (N_12359,N_8091,N_9555);
or U12360 (N_12360,N_6020,N_5497);
or U12361 (N_12361,N_6501,N_9914);
xnor U12362 (N_12362,N_8726,N_9902);
and U12363 (N_12363,N_6419,N_8682);
and U12364 (N_12364,N_8990,N_6597);
and U12365 (N_12365,N_5783,N_7331);
nor U12366 (N_12366,N_8423,N_5713);
nand U12367 (N_12367,N_8284,N_6198);
or U12368 (N_12368,N_8956,N_8706);
nor U12369 (N_12369,N_9898,N_7410);
xor U12370 (N_12370,N_7358,N_6488);
xnor U12371 (N_12371,N_9371,N_8442);
and U12372 (N_12372,N_6365,N_7519);
or U12373 (N_12373,N_5072,N_5646);
nand U12374 (N_12374,N_6636,N_8039);
nor U12375 (N_12375,N_7223,N_9554);
nor U12376 (N_12376,N_7577,N_6786);
nor U12377 (N_12377,N_6888,N_8952);
or U12378 (N_12378,N_5540,N_5838);
or U12379 (N_12379,N_9673,N_8425);
and U12380 (N_12380,N_9427,N_7792);
or U12381 (N_12381,N_8732,N_8589);
or U12382 (N_12382,N_8431,N_7286);
or U12383 (N_12383,N_9985,N_9753);
and U12384 (N_12384,N_8878,N_5506);
xnor U12385 (N_12385,N_9218,N_6897);
nor U12386 (N_12386,N_7794,N_9835);
nand U12387 (N_12387,N_8617,N_6543);
nand U12388 (N_12388,N_9944,N_5431);
nor U12389 (N_12389,N_7306,N_6170);
or U12390 (N_12390,N_6837,N_6467);
nor U12391 (N_12391,N_9143,N_8573);
or U12392 (N_12392,N_6183,N_5592);
xor U12393 (N_12393,N_5224,N_9082);
nand U12394 (N_12394,N_5301,N_5456);
nand U12395 (N_12395,N_5192,N_8770);
and U12396 (N_12396,N_6045,N_8451);
nand U12397 (N_12397,N_9992,N_8747);
or U12398 (N_12398,N_8810,N_9643);
or U12399 (N_12399,N_9024,N_9784);
and U12400 (N_12400,N_6521,N_6607);
or U12401 (N_12401,N_8892,N_5962);
nand U12402 (N_12402,N_7676,N_7992);
nand U12403 (N_12403,N_7036,N_7163);
or U12404 (N_12404,N_7747,N_7416);
nor U12405 (N_12405,N_6637,N_9151);
nor U12406 (N_12406,N_5463,N_5931);
and U12407 (N_12407,N_5744,N_6649);
nor U12408 (N_12408,N_6769,N_6566);
and U12409 (N_12409,N_7154,N_6013);
nor U12410 (N_12410,N_9268,N_8736);
xor U12411 (N_12411,N_5748,N_5462);
or U12412 (N_12412,N_5716,N_5645);
and U12413 (N_12413,N_8583,N_9875);
and U12414 (N_12414,N_8924,N_9421);
nand U12415 (N_12415,N_7554,N_7395);
and U12416 (N_12416,N_9050,N_8049);
nor U12417 (N_12417,N_5109,N_6348);
xnor U12418 (N_12418,N_7183,N_6835);
xor U12419 (N_12419,N_6535,N_5530);
or U12420 (N_12420,N_7640,N_8229);
nor U12421 (N_12421,N_7332,N_5242);
or U12422 (N_12422,N_8739,N_7586);
nor U12423 (N_12423,N_9566,N_6444);
and U12424 (N_12424,N_9482,N_5786);
nor U12425 (N_12425,N_9311,N_7496);
nor U12426 (N_12426,N_6201,N_5330);
nor U12427 (N_12427,N_5791,N_7194);
and U12428 (N_12428,N_6393,N_6924);
or U12429 (N_12429,N_6168,N_5691);
or U12430 (N_12430,N_6528,N_8446);
xnor U12431 (N_12431,N_6305,N_9622);
nor U12432 (N_12432,N_7376,N_7582);
nand U12433 (N_12433,N_6599,N_7738);
or U12434 (N_12434,N_9247,N_9291);
or U12435 (N_12435,N_6498,N_5924);
nor U12436 (N_12436,N_8299,N_8671);
and U12437 (N_12437,N_6711,N_6114);
xnor U12438 (N_12438,N_5094,N_8087);
nand U12439 (N_12439,N_6473,N_5600);
and U12440 (N_12440,N_9305,N_8808);
nand U12441 (N_12441,N_6132,N_9518);
or U12442 (N_12442,N_6588,N_5127);
nand U12443 (N_12443,N_9068,N_5945);
nor U12444 (N_12444,N_6044,N_8647);
xor U12445 (N_12445,N_5423,N_8060);
xnor U12446 (N_12446,N_9953,N_7203);
and U12447 (N_12447,N_5856,N_8246);
nand U12448 (N_12448,N_5063,N_5283);
or U12449 (N_12449,N_7816,N_7489);
or U12450 (N_12450,N_5624,N_5493);
nand U12451 (N_12451,N_7891,N_8763);
nand U12452 (N_12452,N_6961,N_6063);
xor U12453 (N_12453,N_7254,N_7177);
nand U12454 (N_12454,N_5789,N_9683);
or U12455 (N_12455,N_5436,N_5125);
nand U12456 (N_12456,N_9267,N_5287);
nor U12457 (N_12457,N_5005,N_5033);
nand U12458 (N_12458,N_6745,N_7851);
xnor U12459 (N_12459,N_9251,N_9211);
nand U12460 (N_12460,N_8262,N_5712);
nor U12461 (N_12461,N_6906,N_8505);
or U12462 (N_12462,N_7662,N_7935);
nor U12463 (N_12463,N_5484,N_9779);
and U12464 (N_12464,N_6394,N_5290);
nand U12465 (N_12465,N_5338,N_8096);
or U12466 (N_12466,N_5096,N_8274);
nor U12467 (N_12467,N_7999,N_9333);
nor U12468 (N_12468,N_6793,N_5308);
nand U12469 (N_12469,N_6660,N_7352);
and U12470 (N_12470,N_8448,N_8026);
nor U12471 (N_12471,N_6322,N_9442);
nand U12472 (N_12472,N_6284,N_8688);
xnor U12473 (N_12473,N_6524,N_6565);
xnor U12474 (N_12474,N_9813,N_6939);
nand U12475 (N_12475,N_8149,N_9818);
nor U12476 (N_12476,N_7246,N_7913);
nor U12477 (N_12477,N_8354,N_5577);
nand U12478 (N_12478,N_8116,N_7195);
or U12479 (N_12479,N_5898,N_5448);
nand U12480 (N_12480,N_6753,N_6440);
or U12481 (N_12481,N_7334,N_8926);
nor U12482 (N_12482,N_7283,N_8496);
nand U12483 (N_12483,N_9968,N_8389);
and U12484 (N_12484,N_8427,N_6319);
or U12485 (N_12485,N_7536,N_9699);
nand U12486 (N_12486,N_9285,N_5320);
or U12487 (N_12487,N_7556,N_6638);
nand U12488 (N_12488,N_5253,N_5039);
nor U12489 (N_12489,N_7481,N_6545);
nor U12490 (N_12490,N_8334,N_7318);
nor U12491 (N_12491,N_9192,N_9275);
nor U12492 (N_12492,N_7727,N_7768);
nand U12493 (N_12493,N_7686,N_5642);
nor U12494 (N_12494,N_8495,N_8157);
or U12495 (N_12495,N_8608,N_6061);
or U12496 (N_12496,N_6984,N_7834);
and U12497 (N_12497,N_7598,N_5515);
and U12498 (N_12498,N_8192,N_6760);
or U12499 (N_12499,N_6073,N_8931);
and U12500 (N_12500,N_6552,N_9795);
or U12501 (N_12501,N_8312,N_9733);
and U12502 (N_12502,N_6360,N_5845);
or U12503 (N_12503,N_8505,N_8314);
nor U12504 (N_12504,N_9682,N_7578);
nor U12505 (N_12505,N_7721,N_9448);
and U12506 (N_12506,N_7746,N_8092);
nand U12507 (N_12507,N_8395,N_5744);
nand U12508 (N_12508,N_8738,N_8772);
nand U12509 (N_12509,N_5852,N_8135);
nand U12510 (N_12510,N_9025,N_7663);
nor U12511 (N_12511,N_5149,N_8043);
nor U12512 (N_12512,N_9092,N_8125);
nor U12513 (N_12513,N_8906,N_5398);
nor U12514 (N_12514,N_6379,N_5349);
or U12515 (N_12515,N_9873,N_6319);
nand U12516 (N_12516,N_5982,N_8334);
xor U12517 (N_12517,N_5598,N_7478);
and U12518 (N_12518,N_7797,N_7025);
and U12519 (N_12519,N_7307,N_8292);
xor U12520 (N_12520,N_6216,N_5915);
or U12521 (N_12521,N_8043,N_6326);
or U12522 (N_12522,N_9288,N_5033);
or U12523 (N_12523,N_7668,N_9110);
or U12524 (N_12524,N_6443,N_7893);
and U12525 (N_12525,N_8440,N_7029);
nor U12526 (N_12526,N_9612,N_6953);
nand U12527 (N_12527,N_7449,N_9277);
nand U12528 (N_12528,N_5585,N_5482);
xnor U12529 (N_12529,N_6689,N_9659);
nand U12530 (N_12530,N_8940,N_5206);
and U12531 (N_12531,N_7103,N_8181);
and U12532 (N_12532,N_5890,N_7657);
and U12533 (N_12533,N_9623,N_9646);
xnor U12534 (N_12534,N_9768,N_8207);
nand U12535 (N_12535,N_7092,N_7447);
nand U12536 (N_12536,N_9416,N_7866);
and U12537 (N_12537,N_6340,N_9896);
or U12538 (N_12538,N_7183,N_5182);
nor U12539 (N_12539,N_7258,N_7816);
or U12540 (N_12540,N_6396,N_7243);
or U12541 (N_12541,N_5038,N_5510);
or U12542 (N_12542,N_5985,N_7179);
or U12543 (N_12543,N_8507,N_7633);
or U12544 (N_12544,N_5647,N_8306);
nand U12545 (N_12545,N_5801,N_6789);
xnor U12546 (N_12546,N_7500,N_8595);
and U12547 (N_12547,N_6892,N_5862);
or U12548 (N_12548,N_8217,N_6773);
xnor U12549 (N_12549,N_9127,N_9826);
or U12550 (N_12550,N_9084,N_6831);
nand U12551 (N_12551,N_8043,N_6909);
nor U12552 (N_12552,N_7047,N_6294);
and U12553 (N_12553,N_5929,N_5449);
nor U12554 (N_12554,N_9824,N_7573);
and U12555 (N_12555,N_6491,N_7381);
and U12556 (N_12556,N_9536,N_7850);
nor U12557 (N_12557,N_8991,N_7780);
nand U12558 (N_12558,N_6675,N_5992);
nor U12559 (N_12559,N_9872,N_9397);
and U12560 (N_12560,N_9552,N_8201);
xnor U12561 (N_12561,N_6149,N_6721);
xnor U12562 (N_12562,N_7551,N_5738);
nor U12563 (N_12563,N_9299,N_7537);
nor U12564 (N_12564,N_6006,N_5587);
or U12565 (N_12565,N_6922,N_5276);
nand U12566 (N_12566,N_7814,N_5502);
nand U12567 (N_12567,N_7717,N_6353);
or U12568 (N_12568,N_5290,N_8985);
nand U12569 (N_12569,N_7681,N_5765);
or U12570 (N_12570,N_7414,N_5893);
or U12571 (N_12571,N_7965,N_7061);
nor U12572 (N_12572,N_5404,N_8689);
or U12573 (N_12573,N_7875,N_9727);
nand U12574 (N_12574,N_8407,N_7134);
xnor U12575 (N_12575,N_7098,N_6469);
or U12576 (N_12576,N_5073,N_7829);
nor U12577 (N_12577,N_9735,N_5240);
and U12578 (N_12578,N_6900,N_6828);
nand U12579 (N_12579,N_7937,N_6258);
nor U12580 (N_12580,N_7570,N_9425);
nand U12581 (N_12581,N_5936,N_7351);
or U12582 (N_12582,N_5799,N_8468);
nor U12583 (N_12583,N_9018,N_8826);
nand U12584 (N_12584,N_8163,N_9083);
nor U12585 (N_12585,N_9480,N_8413);
nand U12586 (N_12586,N_9303,N_7284);
nor U12587 (N_12587,N_6515,N_5238);
and U12588 (N_12588,N_8851,N_6499);
nor U12589 (N_12589,N_7612,N_5436);
xor U12590 (N_12590,N_6747,N_9439);
nor U12591 (N_12591,N_5149,N_8746);
or U12592 (N_12592,N_9460,N_9609);
nand U12593 (N_12593,N_8743,N_8354);
nor U12594 (N_12594,N_8191,N_6184);
and U12595 (N_12595,N_6650,N_9242);
nor U12596 (N_12596,N_9776,N_6264);
nand U12597 (N_12597,N_5246,N_6726);
or U12598 (N_12598,N_9308,N_5407);
and U12599 (N_12599,N_7236,N_6098);
nor U12600 (N_12600,N_9415,N_8263);
and U12601 (N_12601,N_5484,N_6585);
nor U12602 (N_12602,N_5970,N_7568);
nor U12603 (N_12603,N_6606,N_7213);
nand U12604 (N_12604,N_5495,N_7128);
nand U12605 (N_12605,N_5102,N_6477);
xnor U12606 (N_12606,N_5668,N_5918);
or U12607 (N_12607,N_5805,N_7928);
nor U12608 (N_12608,N_8401,N_7617);
and U12609 (N_12609,N_5735,N_8746);
and U12610 (N_12610,N_7308,N_9601);
nor U12611 (N_12611,N_6282,N_8952);
nor U12612 (N_12612,N_5590,N_5739);
or U12613 (N_12613,N_8658,N_7821);
nand U12614 (N_12614,N_6207,N_8893);
nand U12615 (N_12615,N_8002,N_9438);
xor U12616 (N_12616,N_7906,N_7750);
nand U12617 (N_12617,N_8035,N_7700);
nand U12618 (N_12618,N_6586,N_5068);
or U12619 (N_12619,N_7043,N_8019);
or U12620 (N_12620,N_7665,N_8852);
nand U12621 (N_12621,N_8231,N_9314);
or U12622 (N_12622,N_5476,N_7011);
xnor U12623 (N_12623,N_7129,N_9909);
and U12624 (N_12624,N_7832,N_9725);
and U12625 (N_12625,N_6182,N_6843);
or U12626 (N_12626,N_8744,N_8147);
nor U12627 (N_12627,N_8595,N_8949);
nand U12628 (N_12628,N_6568,N_5569);
nand U12629 (N_12629,N_7936,N_6783);
and U12630 (N_12630,N_5064,N_7464);
nor U12631 (N_12631,N_9178,N_7145);
and U12632 (N_12632,N_9973,N_9992);
or U12633 (N_12633,N_7752,N_7081);
nor U12634 (N_12634,N_7640,N_5954);
or U12635 (N_12635,N_7603,N_6496);
nor U12636 (N_12636,N_8202,N_5853);
nand U12637 (N_12637,N_6457,N_9167);
nor U12638 (N_12638,N_9242,N_6074);
nor U12639 (N_12639,N_7127,N_8031);
and U12640 (N_12640,N_9294,N_5028);
nand U12641 (N_12641,N_8283,N_5472);
xor U12642 (N_12642,N_8678,N_8538);
and U12643 (N_12643,N_9266,N_5121);
or U12644 (N_12644,N_6103,N_9012);
xnor U12645 (N_12645,N_6242,N_6860);
nor U12646 (N_12646,N_5206,N_8043);
and U12647 (N_12647,N_9305,N_8121);
or U12648 (N_12648,N_9535,N_6940);
and U12649 (N_12649,N_5032,N_7051);
and U12650 (N_12650,N_7356,N_9841);
nor U12651 (N_12651,N_5580,N_9294);
nand U12652 (N_12652,N_5222,N_6340);
and U12653 (N_12653,N_5330,N_9138);
nand U12654 (N_12654,N_5614,N_9012);
nand U12655 (N_12655,N_9882,N_8411);
nand U12656 (N_12656,N_8969,N_5684);
and U12657 (N_12657,N_9273,N_6390);
nand U12658 (N_12658,N_9487,N_7242);
and U12659 (N_12659,N_7798,N_8530);
and U12660 (N_12660,N_9323,N_8680);
or U12661 (N_12661,N_6955,N_6397);
and U12662 (N_12662,N_5207,N_5333);
or U12663 (N_12663,N_9772,N_6644);
nor U12664 (N_12664,N_5700,N_8598);
and U12665 (N_12665,N_9127,N_9397);
or U12666 (N_12666,N_8748,N_7661);
and U12667 (N_12667,N_5305,N_6713);
and U12668 (N_12668,N_9503,N_9143);
nand U12669 (N_12669,N_9600,N_6163);
and U12670 (N_12670,N_5654,N_6864);
nor U12671 (N_12671,N_5827,N_8761);
nand U12672 (N_12672,N_5553,N_7474);
nor U12673 (N_12673,N_9313,N_6340);
nor U12674 (N_12674,N_5159,N_5615);
or U12675 (N_12675,N_6658,N_6293);
nor U12676 (N_12676,N_9890,N_7184);
and U12677 (N_12677,N_5246,N_6497);
or U12678 (N_12678,N_8341,N_6006);
or U12679 (N_12679,N_5769,N_9748);
xor U12680 (N_12680,N_7545,N_6518);
nand U12681 (N_12681,N_8389,N_6275);
and U12682 (N_12682,N_8781,N_5179);
nand U12683 (N_12683,N_5550,N_6174);
nand U12684 (N_12684,N_9018,N_8769);
nand U12685 (N_12685,N_7399,N_5135);
nor U12686 (N_12686,N_9946,N_5382);
xor U12687 (N_12687,N_9451,N_8342);
nand U12688 (N_12688,N_7452,N_6401);
and U12689 (N_12689,N_6491,N_8786);
nand U12690 (N_12690,N_9997,N_5362);
or U12691 (N_12691,N_6082,N_9267);
or U12692 (N_12692,N_5193,N_6131);
or U12693 (N_12693,N_8885,N_7702);
or U12694 (N_12694,N_6546,N_5585);
nand U12695 (N_12695,N_5029,N_8895);
nand U12696 (N_12696,N_5347,N_8830);
or U12697 (N_12697,N_6378,N_6874);
nand U12698 (N_12698,N_7246,N_8181);
or U12699 (N_12699,N_5765,N_5605);
and U12700 (N_12700,N_8381,N_5430);
xnor U12701 (N_12701,N_6781,N_5773);
xnor U12702 (N_12702,N_6471,N_8414);
or U12703 (N_12703,N_9469,N_9651);
nor U12704 (N_12704,N_5944,N_6837);
xor U12705 (N_12705,N_6352,N_7484);
nor U12706 (N_12706,N_8188,N_8633);
nand U12707 (N_12707,N_9738,N_6836);
nand U12708 (N_12708,N_6780,N_8302);
or U12709 (N_12709,N_6120,N_7353);
and U12710 (N_12710,N_6229,N_5746);
nand U12711 (N_12711,N_5795,N_6858);
nor U12712 (N_12712,N_7873,N_6095);
and U12713 (N_12713,N_5795,N_5015);
xor U12714 (N_12714,N_6022,N_6016);
and U12715 (N_12715,N_6950,N_6596);
nor U12716 (N_12716,N_7850,N_9721);
xnor U12717 (N_12717,N_5575,N_7150);
nor U12718 (N_12718,N_6909,N_6749);
and U12719 (N_12719,N_8540,N_7422);
and U12720 (N_12720,N_9443,N_9822);
nor U12721 (N_12721,N_7217,N_6085);
or U12722 (N_12722,N_7784,N_6953);
nor U12723 (N_12723,N_9352,N_9122);
nor U12724 (N_12724,N_6229,N_9287);
xnor U12725 (N_12725,N_6817,N_5937);
nor U12726 (N_12726,N_8024,N_5410);
nor U12727 (N_12727,N_7053,N_6299);
or U12728 (N_12728,N_7354,N_9824);
nor U12729 (N_12729,N_5913,N_7284);
and U12730 (N_12730,N_9975,N_9394);
nand U12731 (N_12731,N_8383,N_7500);
nor U12732 (N_12732,N_7496,N_5520);
nor U12733 (N_12733,N_8380,N_5092);
or U12734 (N_12734,N_9046,N_9820);
and U12735 (N_12735,N_5247,N_6143);
xor U12736 (N_12736,N_9156,N_5112);
and U12737 (N_12737,N_6111,N_6971);
or U12738 (N_12738,N_5768,N_7720);
xor U12739 (N_12739,N_5360,N_6960);
nor U12740 (N_12740,N_9432,N_7165);
and U12741 (N_12741,N_9462,N_6393);
nor U12742 (N_12742,N_6984,N_8516);
nand U12743 (N_12743,N_8736,N_8857);
nor U12744 (N_12744,N_5329,N_5401);
nand U12745 (N_12745,N_5004,N_9879);
and U12746 (N_12746,N_5332,N_7577);
nor U12747 (N_12747,N_5918,N_8515);
and U12748 (N_12748,N_7700,N_6441);
nand U12749 (N_12749,N_8933,N_8891);
or U12750 (N_12750,N_9062,N_7073);
nand U12751 (N_12751,N_6606,N_7475);
or U12752 (N_12752,N_8117,N_5741);
nor U12753 (N_12753,N_7405,N_6614);
or U12754 (N_12754,N_6580,N_7281);
or U12755 (N_12755,N_7204,N_6170);
xnor U12756 (N_12756,N_8211,N_8646);
and U12757 (N_12757,N_5923,N_7205);
and U12758 (N_12758,N_5459,N_8552);
and U12759 (N_12759,N_7652,N_9769);
and U12760 (N_12760,N_6051,N_9736);
and U12761 (N_12761,N_5528,N_7836);
or U12762 (N_12762,N_7134,N_6537);
and U12763 (N_12763,N_8625,N_5957);
or U12764 (N_12764,N_8792,N_6724);
and U12765 (N_12765,N_6711,N_6485);
and U12766 (N_12766,N_7295,N_9464);
or U12767 (N_12767,N_6685,N_5273);
nand U12768 (N_12768,N_8467,N_6402);
xnor U12769 (N_12769,N_8526,N_9033);
and U12770 (N_12770,N_5210,N_5256);
and U12771 (N_12771,N_6058,N_9864);
nor U12772 (N_12772,N_9785,N_7214);
and U12773 (N_12773,N_5398,N_6097);
nand U12774 (N_12774,N_5726,N_9187);
or U12775 (N_12775,N_6627,N_6384);
xnor U12776 (N_12776,N_8942,N_7325);
xor U12777 (N_12777,N_6280,N_7157);
nand U12778 (N_12778,N_7173,N_9195);
or U12779 (N_12779,N_9768,N_7055);
and U12780 (N_12780,N_5570,N_6825);
nor U12781 (N_12781,N_9223,N_8404);
xor U12782 (N_12782,N_8218,N_5589);
and U12783 (N_12783,N_9562,N_7280);
and U12784 (N_12784,N_8896,N_6967);
xor U12785 (N_12785,N_5881,N_8261);
and U12786 (N_12786,N_9893,N_5316);
or U12787 (N_12787,N_6462,N_5974);
and U12788 (N_12788,N_8922,N_6368);
xor U12789 (N_12789,N_5826,N_7029);
xor U12790 (N_12790,N_5602,N_9952);
or U12791 (N_12791,N_6166,N_6939);
or U12792 (N_12792,N_9287,N_9540);
nor U12793 (N_12793,N_7639,N_8401);
and U12794 (N_12794,N_5342,N_7150);
nor U12795 (N_12795,N_6358,N_6047);
nand U12796 (N_12796,N_5893,N_7901);
nand U12797 (N_12797,N_5677,N_8295);
nand U12798 (N_12798,N_8962,N_9550);
nor U12799 (N_12799,N_7192,N_5334);
nor U12800 (N_12800,N_9288,N_9075);
nor U12801 (N_12801,N_9831,N_5434);
nand U12802 (N_12802,N_6658,N_6488);
and U12803 (N_12803,N_8261,N_7283);
nor U12804 (N_12804,N_6740,N_9538);
xor U12805 (N_12805,N_7956,N_7707);
and U12806 (N_12806,N_8385,N_6242);
or U12807 (N_12807,N_9662,N_8450);
or U12808 (N_12808,N_9991,N_5007);
or U12809 (N_12809,N_8957,N_9831);
nand U12810 (N_12810,N_9956,N_7941);
or U12811 (N_12811,N_6790,N_7323);
nand U12812 (N_12812,N_5173,N_8756);
nand U12813 (N_12813,N_6831,N_8508);
or U12814 (N_12814,N_6930,N_7337);
nor U12815 (N_12815,N_5675,N_9392);
nor U12816 (N_12816,N_6550,N_9267);
nand U12817 (N_12817,N_5050,N_5364);
or U12818 (N_12818,N_5249,N_6698);
and U12819 (N_12819,N_9785,N_9171);
xor U12820 (N_12820,N_8609,N_6416);
nand U12821 (N_12821,N_9733,N_7764);
and U12822 (N_12822,N_7285,N_7932);
or U12823 (N_12823,N_7337,N_8492);
or U12824 (N_12824,N_9599,N_6134);
and U12825 (N_12825,N_7917,N_6879);
nand U12826 (N_12826,N_7847,N_8679);
and U12827 (N_12827,N_5713,N_7536);
nor U12828 (N_12828,N_7669,N_8901);
or U12829 (N_12829,N_9116,N_8649);
nand U12830 (N_12830,N_9264,N_9776);
and U12831 (N_12831,N_8150,N_5199);
or U12832 (N_12832,N_7367,N_9697);
xnor U12833 (N_12833,N_7306,N_5702);
nor U12834 (N_12834,N_5721,N_9829);
xor U12835 (N_12835,N_9469,N_6217);
and U12836 (N_12836,N_6393,N_6422);
and U12837 (N_12837,N_5118,N_9519);
and U12838 (N_12838,N_5040,N_7099);
nor U12839 (N_12839,N_8959,N_6353);
or U12840 (N_12840,N_8214,N_6484);
and U12841 (N_12841,N_8642,N_6493);
xnor U12842 (N_12842,N_8069,N_5068);
nor U12843 (N_12843,N_5858,N_6855);
or U12844 (N_12844,N_8830,N_8409);
nor U12845 (N_12845,N_9971,N_6456);
and U12846 (N_12846,N_7438,N_7340);
nor U12847 (N_12847,N_6919,N_8433);
nand U12848 (N_12848,N_9798,N_9744);
nand U12849 (N_12849,N_7330,N_6500);
and U12850 (N_12850,N_9166,N_7439);
or U12851 (N_12851,N_6400,N_8987);
or U12852 (N_12852,N_6945,N_9703);
and U12853 (N_12853,N_9766,N_6539);
or U12854 (N_12854,N_8605,N_5503);
and U12855 (N_12855,N_6082,N_5504);
nand U12856 (N_12856,N_6997,N_5715);
nand U12857 (N_12857,N_8479,N_9819);
or U12858 (N_12858,N_9553,N_5629);
nand U12859 (N_12859,N_5904,N_5219);
nand U12860 (N_12860,N_9062,N_8793);
or U12861 (N_12861,N_5878,N_7512);
nand U12862 (N_12862,N_5276,N_7002);
nand U12863 (N_12863,N_5581,N_7373);
and U12864 (N_12864,N_6989,N_9062);
and U12865 (N_12865,N_8826,N_8484);
nand U12866 (N_12866,N_9848,N_6614);
and U12867 (N_12867,N_6142,N_8842);
nand U12868 (N_12868,N_6912,N_9591);
nand U12869 (N_12869,N_8177,N_9049);
xor U12870 (N_12870,N_7423,N_9768);
and U12871 (N_12871,N_8867,N_5249);
and U12872 (N_12872,N_8615,N_9436);
and U12873 (N_12873,N_7629,N_6305);
xnor U12874 (N_12874,N_6994,N_8588);
and U12875 (N_12875,N_5173,N_9294);
nand U12876 (N_12876,N_9783,N_6645);
and U12877 (N_12877,N_6799,N_6591);
nand U12878 (N_12878,N_9444,N_5385);
nand U12879 (N_12879,N_9951,N_7450);
nand U12880 (N_12880,N_8362,N_9207);
or U12881 (N_12881,N_5346,N_5955);
nor U12882 (N_12882,N_8084,N_9502);
or U12883 (N_12883,N_7339,N_7197);
nor U12884 (N_12884,N_5422,N_7543);
xor U12885 (N_12885,N_8368,N_8301);
nor U12886 (N_12886,N_7525,N_8678);
nor U12887 (N_12887,N_6129,N_5497);
and U12888 (N_12888,N_6578,N_5647);
and U12889 (N_12889,N_9379,N_5335);
nand U12890 (N_12890,N_5866,N_8860);
or U12891 (N_12891,N_7168,N_6532);
nand U12892 (N_12892,N_8929,N_8077);
or U12893 (N_12893,N_8156,N_7867);
or U12894 (N_12894,N_6423,N_5066);
and U12895 (N_12895,N_5472,N_8745);
nand U12896 (N_12896,N_7517,N_9094);
and U12897 (N_12897,N_5381,N_6065);
nand U12898 (N_12898,N_9614,N_9391);
or U12899 (N_12899,N_5710,N_9711);
nand U12900 (N_12900,N_9137,N_7517);
nand U12901 (N_12901,N_9844,N_6491);
and U12902 (N_12902,N_5286,N_7624);
nor U12903 (N_12903,N_6099,N_9770);
and U12904 (N_12904,N_6767,N_5191);
nand U12905 (N_12905,N_8177,N_6726);
nand U12906 (N_12906,N_6855,N_6996);
and U12907 (N_12907,N_6197,N_6864);
nand U12908 (N_12908,N_6608,N_6229);
nor U12909 (N_12909,N_7939,N_8320);
or U12910 (N_12910,N_9969,N_9773);
nor U12911 (N_12911,N_5726,N_8316);
nand U12912 (N_12912,N_8373,N_5404);
and U12913 (N_12913,N_9837,N_8992);
and U12914 (N_12914,N_9118,N_9526);
or U12915 (N_12915,N_5700,N_9329);
nand U12916 (N_12916,N_9090,N_5686);
or U12917 (N_12917,N_8928,N_9402);
xnor U12918 (N_12918,N_6783,N_9806);
nor U12919 (N_12919,N_5487,N_7309);
nand U12920 (N_12920,N_9145,N_7856);
nand U12921 (N_12921,N_5667,N_9089);
nor U12922 (N_12922,N_6908,N_5824);
or U12923 (N_12923,N_5764,N_6739);
nand U12924 (N_12924,N_7378,N_7879);
nor U12925 (N_12925,N_6814,N_6143);
nand U12926 (N_12926,N_6160,N_8679);
nor U12927 (N_12927,N_8124,N_8778);
nor U12928 (N_12928,N_9217,N_7829);
nand U12929 (N_12929,N_5187,N_8901);
nor U12930 (N_12930,N_9435,N_7071);
and U12931 (N_12931,N_6699,N_8181);
xor U12932 (N_12932,N_7673,N_9778);
nor U12933 (N_12933,N_9214,N_5658);
nor U12934 (N_12934,N_5437,N_5133);
nand U12935 (N_12935,N_8531,N_9846);
xor U12936 (N_12936,N_9276,N_5042);
or U12937 (N_12937,N_5449,N_9739);
nand U12938 (N_12938,N_6328,N_9474);
nor U12939 (N_12939,N_8122,N_6418);
xor U12940 (N_12940,N_9390,N_8395);
nand U12941 (N_12941,N_9623,N_9849);
and U12942 (N_12942,N_5854,N_9549);
nand U12943 (N_12943,N_5756,N_5376);
or U12944 (N_12944,N_9724,N_8296);
xnor U12945 (N_12945,N_8413,N_6454);
nand U12946 (N_12946,N_6269,N_7089);
xor U12947 (N_12947,N_9402,N_7244);
and U12948 (N_12948,N_7663,N_7936);
and U12949 (N_12949,N_5468,N_5032);
xor U12950 (N_12950,N_8081,N_9724);
and U12951 (N_12951,N_9352,N_6337);
and U12952 (N_12952,N_7013,N_8379);
or U12953 (N_12953,N_6228,N_8180);
or U12954 (N_12954,N_6422,N_5363);
or U12955 (N_12955,N_8082,N_8178);
or U12956 (N_12956,N_9871,N_5892);
or U12957 (N_12957,N_9365,N_9980);
nand U12958 (N_12958,N_6247,N_5688);
nor U12959 (N_12959,N_6739,N_9538);
or U12960 (N_12960,N_5515,N_9811);
and U12961 (N_12961,N_9209,N_5769);
and U12962 (N_12962,N_8491,N_8381);
or U12963 (N_12963,N_7402,N_9082);
nand U12964 (N_12964,N_8923,N_5291);
nor U12965 (N_12965,N_6323,N_8312);
xnor U12966 (N_12966,N_8350,N_8134);
nor U12967 (N_12967,N_7729,N_6762);
nand U12968 (N_12968,N_6153,N_9079);
and U12969 (N_12969,N_5008,N_8562);
or U12970 (N_12970,N_7255,N_8753);
and U12971 (N_12971,N_8557,N_6011);
nor U12972 (N_12972,N_7066,N_8540);
nand U12973 (N_12973,N_5430,N_8488);
and U12974 (N_12974,N_9585,N_5704);
nand U12975 (N_12975,N_8998,N_8030);
nor U12976 (N_12976,N_5503,N_6943);
and U12977 (N_12977,N_5385,N_5468);
nand U12978 (N_12978,N_7690,N_9250);
or U12979 (N_12979,N_6830,N_7653);
nand U12980 (N_12980,N_6526,N_5954);
xnor U12981 (N_12981,N_8734,N_5084);
or U12982 (N_12982,N_5408,N_9120);
nand U12983 (N_12983,N_8421,N_6540);
or U12984 (N_12984,N_8019,N_6001);
nand U12985 (N_12985,N_8566,N_9734);
nand U12986 (N_12986,N_8941,N_6433);
nand U12987 (N_12987,N_9025,N_5360);
nand U12988 (N_12988,N_6729,N_8644);
nor U12989 (N_12989,N_8571,N_7821);
and U12990 (N_12990,N_8374,N_6624);
nor U12991 (N_12991,N_8251,N_9957);
or U12992 (N_12992,N_6580,N_7882);
nor U12993 (N_12993,N_5288,N_7727);
or U12994 (N_12994,N_9194,N_5580);
or U12995 (N_12995,N_5399,N_8713);
and U12996 (N_12996,N_8564,N_9215);
nand U12997 (N_12997,N_8517,N_8393);
xor U12998 (N_12998,N_5402,N_8321);
nor U12999 (N_12999,N_8965,N_5370);
and U13000 (N_13000,N_5531,N_8781);
or U13001 (N_13001,N_6222,N_9493);
and U13002 (N_13002,N_7401,N_6350);
and U13003 (N_13003,N_5579,N_5562);
or U13004 (N_13004,N_5261,N_7011);
nand U13005 (N_13005,N_7392,N_8016);
and U13006 (N_13006,N_9403,N_9650);
nand U13007 (N_13007,N_5271,N_9871);
xnor U13008 (N_13008,N_5018,N_7045);
nand U13009 (N_13009,N_8747,N_7161);
nand U13010 (N_13010,N_9815,N_8057);
or U13011 (N_13011,N_9996,N_7457);
and U13012 (N_13012,N_7636,N_5988);
nor U13013 (N_13013,N_9288,N_9838);
xnor U13014 (N_13014,N_9866,N_9135);
nor U13015 (N_13015,N_6853,N_8154);
nor U13016 (N_13016,N_5652,N_6125);
nor U13017 (N_13017,N_7329,N_6651);
nor U13018 (N_13018,N_6850,N_6062);
or U13019 (N_13019,N_7899,N_8457);
or U13020 (N_13020,N_5849,N_5874);
or U13021 (N_13021,N_6509,N_8939);
nand U13022 (N_13022,N_6184,N_5323);
nand U13023 (N_13023,N_7053,N_7843);
nor U13024 (N_13024,N_5252,N_9972);
or U13025 (N_13025,N_9796,N_9031);
and U13026 (N_13026,N_9450,N_8803);
or U13027 (N_13027,N_8353,N_8918);
nor U13028 (N_13028,N_9517,N_8786);
or U13029 (N_13029,N_9163,N_5152);
and U13030 (N_13030,N_9946,N_6757);
nor U13031 (N_13031,N_5382,N_6322);
and U13032 (N_13032,N_6082,N_5301);
nor U13033 (N_13033,N_8498,N_8661);
or U13034 (N_13034,N_9372,N_6469);
nor U13035 (N_13035,N_7962,N_9652);
nand U13036 (N_13036,N_7256,N_9710);
nand U13037 (N_13037,N_5016,N_5384);
and U13038 (N_13038,N_9982,N_9759);
nor U13039 (N_13039,N_6797,N_6199);
nor U13040 (N_13040,N_7332,N_7973);
xor U13041 (N_13041,N_5430,N_6895);
nand U13042 (N_13042,N_9282,N_7034);
nor U13043 (N_13043,N_9884,N_8949);
or U13044 (N_13044,N_7575,N_6494);
and U13045 (N_13045,N_6825,N_6729);
nand U13046 (N_13046,N_7226,N_7072);
nand U13047 (N_13047,N_9305,N_7922);
nor U13048 (N_13048,N_5960,N_5871);
nor U13049 (N_13049,N_5101,N_8928);
and U13050 (N_13050,N_6840,N_8439);
nor U13051 (N_13051,N_7986,N_9582);
or U13052 (N_13052,N_6045,N_7657);
xor U13053 (N_13053,N_7930,N_9498);
nor U13054 (N_13054,N_9420,N_6684);
and U13055 (N_13055,N_9916,N_6792);
xor U13056 (N_13056,N_9975,N_8581);
nor U13057 (N_13057,N_7383,N_5467);
or U13058 (N_13058,N_7011,N_5904);
xor U13059 (N_13059,N_9149,N_6379);
nor U13060 (N_13060,N_6052,N_7913);
or U13061 (N_13061,N_8846,N_6284);
and U13062 (N_13062,N_9042,N_6361);
nor U13063 (N_13063,N_5668,N_9157);
nor U13064 (N_13064,N_7142,N_5188);
nor U13065 (N_13065,N_7716,N_5472);
or U13066 (N_13066,N_7347,N_7403);
xnor U13067 (N_13067,N_6275,N_9814);
nand U13068 (N_13068,N_6242,N_8994);
or U13069 (N_13069,N_5881,N_8919);
nand U13070 (N_13070,N_9335,N_9706);
nor U13071 (N_13071,N_6856,N_5447);
nand U13072 (N_13072,N_6472,N_8736);
nand U13073 (N_13073,N_9690,N_6083);
and U13074 (N_13074,N_8214,N_5180);
or U13075 (N_13075,N_8547,N_9686);
and U13076 (N_13076,N_5145,N_6497);
and U13077 (N_13077,N_8174,N_5679);
nand U13078 (N_13078,N_9252,N_8642);
and U13079 (N_13079,N_9996,N_9898);
nand U13080 (N_13080,N_8828,N_6383);
nand U13081 (N_13081,N_9799,N_7803);
xnor U13082 (N_13082,N_8788,N_6259);
or U13083 (N_13083,N_9543,N_9882);
nand U13084 (N_13084,N_5397,N_8507);
nand U13085 (N_13085,N_9934,N_8402);
or U13086 (N_13086,N_9100,N_9046);
or U13087 (N_13087,N_6853,N_5793);
or U13088 (N_13088,N_7247,N_7658);
nand U13089 (N_13089,N_6458,N_9079);
or U13090 (N_13090,N_9679,N_7836);
or U13091 (N_13091,N_5614,N_7526);
and U13092 (N_13092,N_7531,N_8479);
nand U13093 (N_13093,N_5408,N_7224);
and U13094 (N_13094,N_8325,N_6657);
or U13095 (N_13095,N_7823,N_9851);
and U13096 (N_13096,N_9298,N_9756);
or U13097 (N_13097,N_7529,N_9483);
nand U13098 (N_13098,N_8390,N_8547);
nand U13099 (N_13099,N_6000,N_6351);
nand U13100 (N_13100,N_5556,N_7882);
and U13101 (N_13101,N_8749,N_8311);
nor U13102 (N_13102,N_6716,N_5036);
or U13103 (N_13103,N_7319,N_8118);
nor U13104 (N_13104,N_5399,N_6322);
and U13105 (N_13105,N_9114,N_9587);
nor U13106 (N_13106,N_8442,N_5682);
nor U13107 (N_13107,N_6755,N_8515);
xnor U13108 (N_13108,N_5054,N_7099);
and U13109 (N_13109,N_9234,N_7847);
nand U13110 (N_13110,N_7406,N_8297);
nand U13111 (N_13111,N_5782,N_5765);
nor U13112 (N_13112,N_6024,N_7428);
nor U13113 (N_13113,N_5080,N_5688);
and U13114 (N_13114,N_5321,N_7357);
and U13115 (N_13115,N_7205,N_8053);
nor U13116 (N_13116,N_8101,N_7705);
nand U13117 (N_13117,N_7702,N_8146);
nor U13118 (N_13118,N_6874,N_6421);
and U13119 (N_13119,N_5686,N_5460);
or U13120 (N_13120,N_5152,N_8064);
and U13121 (N_13121,N_9755,N_5939);
and U13122 (N_13122,N_8614,N_6674);
nand U13123 (N_13123,N_5671,N_9166);
nor U13124 (N_13124,N_9883,N_5966);
and U13125 (N_13125,N_9186,N_6648);
or U13126 (N_13126,N_6052,N_7821);
nor U13127 (N_13127,N_8285,N_7139);
or U13128 (N_13128,N_8426,N_5213);
and U13129 (N_13129,N_9520,N_5312);
nor U13130 (N_13130,N_6593,N_6280);
nor U13131 (N_13131,N_7178,N_8025);
nand U13132 (N_13132,N_6268,N_5920);
and U13133 (N_13133,N_9522,N_7458);
nand U13134 (N_13134,N_7654,N_6124);
and U13135 (N_13135,N_5392,N_5610);
nor U13136 (N_13136,N_9424,N_7454);
nor U13137 (N_13137,N_5890,N_8797);
and U13138 (N_13138,N_7215,N_9954);
nor U13139 (N_13139,N_8955,N_5614);
and U13140 (N_13140,N_9818,N_9505);
nand U13141 (N_13141,N_5178,N_7978);
or U13142 (N_13142,N_6737,N_7347);
nor U13143 (N_13143,N_7916,N_9111);
nand U13144 (N_13144,N_9304,N_9712);
and U13145 (N_13145,N_8306,N_7488);
and U13146 (N_13146,N_8481,N_9103);
or U13147 (N_13147,N_6569,N_8088);
and U13148 (N_13148,N_9236,N_7495);
nand U13149 (N_13149,N_8413,N_8017);
nand U13150 (N_13150,N_7321,N_7370);
nand U13151 (N_13151,N_8494,N_9764);
nor U13152 (N_13152,N_9945,N_8842);
and U13153 (N_13153,N_9851,N_7883);
or U13154 (N_13154,N_7978,N_8620);
and U13155 (N_13155,N_7021,N_6132);
nor U13156 (N_13156,N_6425,N_7998);
nand U13157 (N_13157,N_9234,N_7790);
or U13158 (N_13158,N_7782,N_6780);
or U13159 (N_13159,N_9278,N_7806);
or U13160 (N_13160,N_9713,N_6349);
or U13161 (N_13161,N_9989,N_9786);
and U13162 (N_13162,N_7175,N_9089);
and U13163 (N_13163,N_9372,N_9666);
or U13164 (N_13164,N_8812,N_9734);
nor U13165 (N_13165,N_8025,N_9410);
nor U13166 (N_13166,N_8279,N_5045);
xor U13167 (N_13167,N_8913,N_9997);
nand U13168 (N_13168,N_8990,N_7458);
nand U13169 (N_13169,N_9616,N_7888);
and U13170 (N_13170,N_8949,N_5839);
nand U13171 (N_13171,N_6289,N_6398);
nand U13172 (N_13172,N_7797,N_7472);
nor U13173 (N_13173,N_6473,N_7545);
nor U13174 (N_13174,N_7437,N_5357);
and U13175 (N_13175,N_6881,N_9634);
or U13176 (N_13176,N_8185,N_9081);
nor U13177 (N_13177,N_7230,N_8186);
and U13178 (N_13178,N_6096,N_9506);
or U13179 (N_13179,N_8736,N_5537);
nand U13180 (N_13180,N_8313,N_8957);
nor U13181 (N_13181,N_9909,N_8504);
nor U13182 (N_13182,N_6059,N_7486);
or U13183 (N_13183,N_8126,N_6088);
nand U13184 (N_13184,N_9516,N_6125);
or U13185 (N_13185,N_5430,N_6125);
nand U13186 (N_13186,N_8630,N_6065);
nor U13187 (N_13187,N_6768,N_6187);
and U13188 (N_13188,N_8648,N_5295);
and U13189 (N_13189,N_7792,N_5710);
and U13190 (N_13190,N_5999,N_6804);
nor U13191 (N_13191,N_5528,N_8059);
or U13192 (N_13192,N_7134,N_6001);
and U13193 (N_13193,N_6726,N_7670);
nor U13194 (N_13194,N_9920,N_8635);
nand U13195 (N_13195,N_7806,N_8532);
nand U13196 (N_13196,N_8053,N_6949);
and U13197 (N_13197,N_9176,N_7291);
nor U13198 (N_13198,N_9047,N_8641);
or U13199 (N_13199,N_6944,N_7285);
and U13200 (N_13200,N_8100,N_6672);
or U13201 (N_13201,N_7080,N_8568);
or U13202 (N_13202,N_6559,N_6337);
and U13203 (N_13203,N_6250,N_7503);
and U13204 (N_13204,N_8492,N_7390);
or U13205 (N_13205,N_7905,N_7727);
nor U13206 (N_13206,N_7064,N_7472);
and U13207 (N_13207,N_6664,N_8047);
nor U13208 (N_13208,N_6898,N_7409);
nand U13209 (N_13209,N_8025,N_5522);
nand U13210 (N_13210,N_5326,N_8669);
or U13211 (N_13211,N_6257,N_8773);
nor U13212 (N_13212,N_5540,N_7859);
nand U13213 (N_13213,N_8637,N_9081);
and U13214 (N_13214,N_8103,N_8502);
xor U13215 (N_13215,N_5376,N_6313);
or U13216 (N_13216,N_6112,N_6126);
and U13217 (N_13217,N_9219,N_8364);
xor U13218 (N_13218,N_8410,N_6288);
nor U13219 (N_13219,N_7811,N_7055);
or U13220 (N_13220,N_8812,N_7756);
xor U13221 (N_13221,N_9535,N_5583);
xor U13222 (N_13222,N_7327,N_8993);
nor U13223 (N_13223,N_5971,N_6078);
nand U13224 (N_13224,N_7930,N_8939);
and U13225 (N_13225,N_7304,N_8323);
nand U13226 (N_13226,N_6431,N_9722);
and U13227 (N_13227,N_7841,N_6738);
nand U13228 (N_13228,N_7575,N_5318);
or U13229 (N_13229,N_7376,N_6270);
nand U13230 (N_13230,N_5482,N_7024);
nor U13231 (N_13231,N_9153,N_7970);
or U13232 (N_13232,N_8581,N_8248);
and U13233 (N_13233,N_9813,N_7338);
or U13234 (N_13234,N_6973,N_6648);
nor U13235 (N_13235,N_7419,N_7061);
nor U13236 (N_13236,N_5291,N_7757);
nor U13237 (N_13237,N_8596,N_6939);
or U13238 (N_13238,N_7726,N_7614);
nand U13239 (N_13239,N_6894,N_9347);
or U13240 (N_13240,N_7390,N_6304);
and U13241 (N_13241,N_8495,N_6433);
nand U13242 (N_13242,N_7850,N_5928);
and U13243 (N_13243,N_7579,N_5019);
nor U13244 (N_13244,N_7978,N_5274);
nand U13245 (N_13245,N_9301,N_9340);
nor U13246 (N_13246,N_5167,N_6983);
xor U13247 (N_13247,N_8533,N_5727);
nor U13248 (N_13248,N_6183,N_9816);
or U13249 (N_13249,N_9587,N_6430);
or U13250 (N_13250,N_5107,N_8855);
xnor U13251 (N_13251,N_8834,N_9109);
nor U13252 (N_13252,N_5856,N_5003);
nor U13253 (N_13253,N_5606,N_9365);
and U13254 (N_13254,N_8784,N_8733);
nand U13255 (N_13255,N_8884,N_5754);
and U13256 (N_13256,N_7233,N_6655);
nor U13257 (N_13257,N_7621,N_6081);
xor U13258 (N_13258,N_9793,N_9315);
and U13259 (N_13259,N_6077,N_5728);
or U13260 (N_13260,N_8067,N_6658);
and U13261 (N_13261,N_7987,N_8500);
or U13262 (N_13262,N_6513,N_9868);
nand U13263 (N_13263,N_7883,N_7322);
or U13264 (N_13264,N_5177,N_6472);
nand U13265 (N_13265,N_6011,N_8787);
nor U13266 (N_13266,N_7815,N_6381);
and U13267 (N_13267,N_6506,N_5948);
and U13268 (N_13268,N_9855,N_7893);
and U13269 (N_13269,N_5004,N_9500);
xor U13270 (N_13270,N_7908,N_5088);
and U13271 (N_13271,N_8229,N_5218);
and U13272 (N_13272,N_5940,N_7302);
nor U13273 (N_13273,N_9801,N_5255);
and U13274 (N_13274,N_8460,N_5560);
or U13275 (N_13275,N_5225,N_7559);
xnor U13276 (N_13276,N_7603,N_9307);
nor U13277 (N_13277,N_5856,N_7569);
and U13278 (N_13278,N_6208,N_9654);
and U13279 (N_13279,N_5498,N_5935);
and U13280 (N_13280,N_5842,N_5094);
nand U13281 (N_13281,N_5237,N_5495);
or U13282 (N_13282,N_7318,N_9644);
nor U13283 (N_13283,N_8253,N_5489);
nand U13284 (N_13284,N_8062,N_8484);
xor U13285 (N_13285,N_9996,N_7301);
nand U13286 (N_13286,N_9740,N_7453);
nor U13287 (N_13287,N_7059,N_8585);
nand U13288 (N_13288,N_9791,N_9103);
nor U13289 (N_13289,N_5567,N_8180);
nor U13290 (N_13290,N_5634,N_5710);
and U13291 (N_13291,N_6370,N_8970);
and U13292 (N_13292,N_7221,N_9918);
nor U13293 (N_13293,N_5300,N_7729);
nand U13294 (N_13294,N_9415,N_8487);
nor U13295 (N_13295,N_6915,N_7236);
nor U13296 (N_13296,N_7820,N_6645);
nand U13297 (N_13297,N_6808,N_8899);
nor U13298 (N_13298,N_6929,N_6353);
or U13299 (N_13299,N_9192,N_7005);
nand U13300 (N_13300,N_6630,N_6131);
or U13301 (N_13301,N_5859,N_7834);
nand U13302 (N_13302,N_5728,N_7243);
nor U13303 (N_13303,N_6925,N_8381);
nand U13304 (N_13304,N_8946,N_8695);
nor U13305 (N_13305,N_7798,N_7097);
nand U13306 (N_13306,N_7413,N_6295);
or U13307 (N_13307,N_9743,N_7283);
or U13308 (N_13308,N_6472,N_9642);
or U13309 (N_13309,N_8302,N_8614);
nand U13310 (N_13310,N_8630,N_7056);
or U13311 (N_13311,N_7729,N_6293);
xor U13312 (N_13312,N_7753,N_8688);
nor U13313 (N_13313,N_9736,N_6687);
nand U13314 (N_13314,N_7070,N_9343);
nand U13315 (N_13315,N_5489,N_6129);
and U13316 (N_13316,N_7332,N_7263);
or U13317 (N_13317,N_9037,N_7156);
xor U13318 (N_13318,N_8750,N_5189);
or U13319 (N_13319,N_7806,N_9180);
or U13320 (N_13320,N_5433,N_5430);
or U13321 (N_13321,N_8169,N_6486);
nand U13322 (N_13322,N_5521,N_6246);
nand U13323 (N_13323,N_9605,N_8280);
nand U13324 (N_13324,N_6560,N_6948);
or U13325 (N_13325,N_5784,N_6704);
nor U13326 (N_13326,N_5035,N_8840);
nor U13327 (N_13327,N_9126,N_7221);
nand U13328 (N_13328,N_5059,N_7409);
nand U13329 (N_13329,N_5072,N_9788);
xor U13330 (N_13330,N_7482,N_7968);
nand U13331 (N_13331,N_5844,N_9231);
and U13332 (N_13332,N_7775,N_5444);
and U13333 (N_13333,N_7697,N_9708);
and U13334 (N_13334,N_7273,N_5230);
and U13335 (N_13335,N_5855,N_5164);
nor U13336 (N_13336,N_8985,N_6249);
nand U13337 (N_13337,N_6017,N_8941);
nand U13338 (N_13338,N_6313,N_5273);
and U13339 (N_13339,N_5520,N_8238);
nand U13340 (N_13340,N_6619,N_6321);
nand U13341 (N_13341,N_6824,N_8871);
nand U13342 (N_13342,N_9325,N_5559);
nand U13343 (N_13343,N_9698,N_6716);
nand U13344 (N_13344,N_8339,N_9816);
or U13345 (N_13345,N_5293,N_6797);
nor U13346 (N_13346,N_5077,N_9542);
or U13347 (N_13347,N_8969,N_6838);
and U13348 (N_13348,N_9208,N_7698);
and U13349 (N_13349,N_6173,N_8201);
or U13350 (N_13350,N_5712,N_8231);
and U13351 (N_13351,N_8013,N_6696);
nor U13352 (N_13352,N_9861,N_7239);
nand U13353 (N_13353,N_5249,N_7250);
nand U13354 (N_13354,N_8967,N_8225);
nor U13355 (N_13355,N_7735,N_8851);
nor U13356 (N_13356,N_7761,N_5540);
and U13357 (N_13357,N_6888,N_8436);
nand U13358 (N_13358,N_7477,N_6033);
nand U13359 (N_13359,N_6559,N_6593);
xnor U13360 (N_13360,N_9725,N_7027);
nand U13361 (N_13361,N_9527,N_6660);
or U13362 (N_13362,N_9817,N_7218);
xor U13363 (N_13363,N_5578,N_6504);
or U13364 (N_13364,N_8772,N_8581);
nand U13365 (N_13365,N_5096,N_7397);
nand U13366 (N_13366,N_5100,N_8513);
or U13367 (N_13367,N_9882,N_5680);
or U13368 (N_13368,N_5287,N_8015);
nor U13369 (N_13369,N_9860,N_8404);
nor U13370 (N_13370,N_8118,N_6230);
nand U13371 (N_13371,N_6044,N_9652);
nor U13372 (N_13372,N_6752,N_8816);
and U13373 (N_13373,N_9240,N_5139);
and U13374 (N_13374,N_6118,N_8884);
or U13375 (N_13375,N_9921,N_7408);
nand U13376 (N_13376,N_6081,N_5100);
or U13377 (N_13377,N_6198,N_9392);
or U13378 (N_13378,N_9856,N_8594);
nand U13379 (N_13379,N_9499,N_6006);
nand U13380 (N_13380,N_9367,N_6229);
and U13381 (N_13381,N_7237,N_7321);
or U13382 (N_13382,N_9646,N_5607);
and U13383 (N_13383,N_6787,N_8610);
nand U13384 (N_13384,N_8403,N_8018);
nor U13385 (N_13385,N_7734,N_9378);
nor U13386 (N_13386,N_5385,N_7158);
and U13387 (N_13387,N_9919,N_9583);
nand U13388 (N_13388,N_5135,N_8862);
and U13389 (N_13389,N_7536,N_5541);
or U13390 (N_13390,N_5684,N_9819);
and U13391 (N_13391,N_6078,N_5885);
or U13392 (N_13392,N_6438,N_9100);
and U13393 (N_13393,N_6474,N_8227);
or U13394 (N_13394,N_6207,N_9762);
or U13395 (N_13395,N_9366,N_6256);
or U13396 (N_13396,N_8702,N_6611);
nand U13397 (N_13397,N_9385,N_7377);
or U13398 (N_13398,N_9797,N_7598);
or U13399 (N_13399,N_5583,N_8720);
nor U13400 (N_13400,N_5151,N_8217);
and U13401 (N_13401,N_8188,N_7958);
nor U13402 (N_13402,N_6258,N_5362);
or U13403 (N_13403,N_7941,N_7033);
and U13404 (N_13404,N_9109,N_9930);
nand U13405 (N_13405,N_6534,N_6600);
xor U13406 (N_13406,N_7250,N_6416);
or U13407 (N_13407,N_5389,N_9743);
nor U13408 (N_13408,N_5125,N_9408);
or U13409 (N_13409,N_8398,N_5996);
or U13410 (N_13410,N_7138,N_5928);
nand U13411 (N_13411,N_6311,N_5377);
or U13412 (N_13412,N_9138,N_7292);
nand U13413 (N_13413,N_7145,N_9697);
nor U13414 (N_13414,N_5973,N_8733);
nor U13415 (N_13415,N_8039,N_6372);
or U13416 (N_13416,N_8235,N_7650);
and U13417 (N_13417,N_7029,N_8588);
nor U13418 (N_13418,N_6919,N_7282);
nand U13419 (N_13419,N_7992,N_6808);
nor U13420 (N_13420,N_8535,N_9394);
nor U13421 (N_13421,N_6331,N_6517);
nor U13422 (N_13422,N_7536,N_7292);
nand U13423 (N_13423,N_5707,N_6257);
nand U13424 (N_13424,N_8796,N_9397);
or U13425 (N_13425,N_5632,N_7719);
or U13426 (N_13426,N_5019,N_5362);
nand U13427 (N_13427,N_6356,N_6037);
nor U13428 (N_13428,N_8568,N_7612);
and U13429 (N_13429,N_8057,N_7806);
nor U13430 (N_13430,N_7113,N_8883);
nand U13431 (N_13431,N_7415,N_5548);
or U13432 (N_13432,N_9446,N_6356);
nand U13433 (N_13433,N_5959,N_8341);
nand U13434 (N_13434,N_9479,N_5507);
nand U13435 (N_13435,N_7884,N_7339);
or U13436 (N_13436,N_5762,N_6616);
nand U13437 (N_13437,N_8950,N_7678);
nand U13438 (N_13438,N_5502,N_6896);
nor U13439 (N_13439,N_5384,N_7867);
nor U13440 (N_13440,N_9116,N_6089);
xor U13441 (N_13441,N_7202,N_9817);
xor U13442 (N_13442,N_5517,N_9631);
nand U13443 (N_13443,N_5207,N_7540);
nor U13444 (N_13444,N_7275,N_7394);
nand U13445 (N_13445,N_8218,N_6944);
nand U13446 (N_13446,N_7665,N_5080);
nor U13447 (N_13447,N_6186,N_9032);
or U13448 (N_13448,N_7700,N_5833);
xor U13449 (N_13449,N_9411,N_6075);
nor U13450 (N_13450,N_7170,N_9886);
or U13451 (N_13451,N_7138,N_9688);
xnor U13452 (N_13452,N_7931,N_9578);
and U13453 (N_13453,N_9813,N_8168);
nor U13454 (N_13454,N_5885,N_8185);
nand U13455 (N_13455,N_6607,N_5143);
nand U13456 (N_13456,N_5208,N_9634);
xor U13457 (N_13457,N_5079,N_6497);
or U13458 (N_13458,N_9930,N_9546);
or U13459 (N_13459,N_7146,N_5152);
or U13460 (N_13460,N_9175,N_9550);
nand U13461 (N_13461,N_8342,N_8298);
nor U13462 (N_13462,N_9520,N_9172);
nand U13463 (N_13463,N_9942,N_9080);
xnor U13464 (N_13464,N_6689,N_7497);
xnor U13465 (N_13465,N_9497,N_8105);
and U13466 (N_13466,N_8744,N_9081);
xnor U13467 (N_13467,N_5115,N_6844);
and U13468 (N_13468,N_9807,N_5712);
and U13469 (N_13469,N_9191,N_6666);
nand U13470 (N_13470,N_8192,N_7648);
and U13471 (N_13471,N_8493,N_7185);
xor U13472 (N_13472,N_9052,N_8105);
or U13473 (N_13473,N_9486,N_5444);
and U13474 (N_13474,N_6840,N_9326);
nand U13475 (N_13475,N_6628,N_5712);
or U13476 (N_13476,N_6624,N_5460);
nor U13477 (N_13477,N_8756,N_6021);
or U13478 (N_13478,N_7415,N_6140);
and U13479 (N_13479,N_8386,N_6641);
and U13480 (N_13480,N_9662,N_8321);
and U13481 (N_13481,N_8341,N_6346);
and U13482 (N_13482,N_5445,N_5218);
xnor U13483 (N_13483,N_8177,N_8362);
xnor U13484 (N_13484,N_7789,N_9847);
xor U13485 (N_13485,N_9662,N_6725);
and U13486 (N_13486,N_6625,N_5364);
or U13487 (N_13487,N_5080,N_9497);
or U13488 (N_13488,N_8754,N_6797);
nor U13489 (N_13489,N_7107,N_5396);
and U13490 (N_13490,N_6520,N_6149);
and U13491 (N_13491,N_7382,N_5679);
or U13492 (N_13492,N_6465,N_5153);
nor U13493 (N_13493,N_9863,N_9642);
and U13494 (N_13494,N_6058,N_8229);
nor U13495 (N_13495,N_8903,N_5524);
nor U13496 (N_13496,N_7189,N_7066);
nor U13497 (N_13497,N_6767,N_7023);
nand U13498 (N_13498,N_9254,N_5249);
nand U13499 (N_13499,N_9833,N_6510);
nand U13500 (N_13500,N_7208,N_8248);
nand U13501 (N_13501,N_7832,N_8864);
nor U13502 (N_13502,N_6741,N_8128);
and U13503 (N_13503,N_9156,N_9853);
nand U13504 (N_13504,N_8248,N_9041);
and U13505 (N_13505,N_6804,N_7902);
and U13506 (N_13506,N_7638,N_5514);
nand U13507 (N_13507,N_8541,N_8023);
nor U13508 (N_13508,N_7364,N_5336);
or U13509 (N_13509,N_6712,N_9346);
nand U13510 (N_13510,N_7849,N_6059);
nand U13511 (N_13511,N_7805,N_7209);
xnor U13512 (N_13512,N_8978,N_6814);
or U13513 (N_13513,N_7200,N_8326);
and U13514 (N_13514,N_5432,N_9808);
and U13515 (N_13515,N_9009,N_6702);
and U13516 (N_13516,N_8548,N_8729);
or U13517 (N_13517,N_7444,N_7356);
and U13518 (N_13518,N_6590,N_9948);
or U13519 (N_13519,N_6701,N_7826);
xnor U13520 (N_13520,N_5459,N_6903);
and U13521 (N_13521,N_7075,N_8249);
and U13522 (N_13522,N_7698,N_5365);
nand U13523 (N_13523,N_9490,N_8697);
and U13524 (N_13524,N_5831,N_6572);
nand U13525 (N_13525,N_8243,N_5496);
nor U13526 (N_13526,N_5943,N_5442);
xor U13527 (N_13527,N_8043,N_9775);
and U13528 (N_13528,N_8726,N_5340);
nor U13529 (N_13529,N_5951,N_8236);
or U13530 (N_13530,N_9861,N_8441);
nor U13531 (N_13531,N_5383,N_7872);
and U13532 (N_13532,N_6654,N_8985);
nor U13533 (N_13533,N_5001,N_5747);
nor U13534 (N_13534,N_8563,N_6670);
nor U13535 (N_13535,N_7063,N_8095);
xor U13536 (N_13536,N_9849,N_7767);
nor U13537 (N_13537,N_6611,N_7574);
nor U13538 (N_13538,N_7157,N_6494);
or U13539 (N_13539,N_7109,N_6513);
nand U13540 (N_13540,N_8843,N_7181);
and U13541 (N_13541,N_5204,N_7945);
or U13542 (N_13542,N_5949,N_6808);
and U13543 (N_13543,N_7574,N_7349);
nand U13544 (N_13544,N_9954,N_5078);
and U13545 (N_13545,N_6588,N_9084);
nand U13546 (N_13546,N_8214,N_7277);
nand U13547 (N_13547,N_8954,N_7986);
nor U13548 (N_13548,N_8958,N_8763);
xor U13549 (N_13549,N_8322,N_7826);
and U13550 (N_13550,N_9697,N_8882);
nand U13551 (N_13551,N_8408,N_8178);
and U13552 (N_13552,N_9700,N_5020);
nand U13553 (N_13553,N_9370,N_6423);
xnor U13554 (N_13554,N_5127,N_6190);
or U13555 (N_13555,N_9364,N_6796);
nand U13556 (N_13556,N_9465,N_7083);
nor U13557 (N_13557,N_7027,N_7263);
and U13558 (N_13558,N_7684,N_8003);
nor U13559 (N_13559,N_8788,N_5638);
and U13560 (N_13560,N_8465,N_5573);
xnor U13561 (N_13561,N_8181,N_8188);
nand U13562 (N_13562,N_5629,N_7707);
or U13563 (N_13563,N_7575,N_7693);
nor U13564 (N_13564,N_6510,N_9655);
nor U13565 (N_13565,N_6341,N_5408);
or U13566 (N_13566,N_9203,N_7294);
xnor U13567 (N_13567,N_8790,N_8144);
and U13568 (N_13568,N_9365,N_5426);
xor U13569 (N_13569,N_6692,N_7048);
and U13570 (N_13570,N_6756,N_6293);
nor U13571 (N_13571,N_5047,N_8020);
and U13572 (N_13572,N_5570,N_6911);
nor U13573 (N_13573,N_5748,N_5514);
nand U13574 (N_13574,N_5410,N_5086);
or U13575 (N_13575,N_6862,N_8154);
nand U13576 (N_13576,N_6040,N_9324);
nand U13577 (N_13577,N_7531,N_9443);
nor U13578 (N_13578,N_5369,N_7782);
nand U13579 (N_13579,N_9803,N_6857);
or U13580 (N_13580,N_5011,N_6546);
nand U13581 (N_13581,N_8022,N_8649);
nor U13582 (N_13582,N_6849,N_7605);
nor U13583 (N_13583,N_5768,N_7264);
or U13584 (N_13584,N_6718,N_8351);
and U13585 (N_13585,N_9031,N_8830);
nand U13586 (N_13586,N_9519,N_5174);
nor U13587 (N_13587,N_8479,N_9895);
and U13588 (N_13588,N_7627,N_9263);
nand U13589 (N_13589,N_8639,N_6751);
nand U13590 (N_13590,N_8611,N_8687);
nand U13591 (N_13591,N_8523,N_7746);
xnor U13592 (N_13592,N_5647,N_8838);
nor U13593 (N_13593,N_8664,N_6244);
nor U13594 (N_13594,N_9653,N_5014);
and U13595 (N_13595,N_8892,N_5820);
or U13596 (N_13596,N_5629,N_9713);
nand U13597 (N_13597,N_6745,N_5891);
nand U13598 (N_13598,N_6822,N_5533);
nand U13599 (N_13599,N_9996,N_7371);
nand U13600 (N_13600,N_6557,N_7718);
or U13601 (N_13601,N_7202,N_8383);
and U13602 (N_13602,N_8813,N_5768);
or U13603 (N_13603,N_6079,N_9381);
nor U13604 (N_13604,N_6751,N_9629);
nand U13605 (N_13605,N_6511,N_8558);
and U13606 (N_13606,N_8466,N_5796);
or U13607 (N_13607,N_8693,N_9168);
nand U13608 (N_13608,N_5978,N_8015);
or U13609 (N_13609,N_5725,N_7521);
or U13610 (N_13610,N_7283,N_5565);
and U13611 (N_13611,N_6736,N_7756);
or U13612 (N_13612,N_7607,N_7704);
or U13613 (N_13613,N_5683,N_8201);
xnor U13614 (N_13614,N_8787,N_8304);
and U13615 (N_13615,N_7357,N_9263);
xnor U13616 (N_13616,N_9621,N_7485);
and U13617 (N_13617,N_7614,N_8635);
nand U13618 (N_13618,N_8371,N_7158);
nor U13619 (N_13619,N_5361,N_6616);
nor U13620 (N_13620,N_6148,N_8577);
and U13621 (N_13621,N_5357,N_8931);
nand U13622 (N_13622,N_7832,N_9038);
nor U13623 (N_13623,N_5638,N_9956);
nor U13624 (N_13624,N_6758,N_8234);
and U13625 (N_13625,N_6238,N_7049);
nand U13626 (N_13626,N_5287,N_8227);
or U13627 (N_13627,N_7402,N_6926);
xnor U13628 (N_13628,N_9486,N_9821);
nand U13629 (N_13629,N_9456,N_5921);
and U13630 (N_13630,N_7179,N_5696);
nand U13631 (N_13631,N_7115,N_8600);
or U13632 (N_13632,N_9549,N_6995);
and U13633 (N_13633,N_8949,N_6178);
xnor U13634 (N_13634,N_5892,N_7657);
and U13635 (N_13635,N_9871,N_5121);
and U13636 (N_13636,N_7509,N_8853);
nor U13637 (N_13637,N_8202,N_6524);
or U13638 (N_13638,N_9098,N_6463);
or U13639 (N_13639,N_7409,N_7279);
nor U13640 (N_13640,N_7799,N_7183);
and U13641 (N_13641,N_5837,N_9428);
nor U13642 (N_13642,N_8107,N_7904);
xor U13643 (N_13643,N_9610,N_8918);
nand U13644 (N_13644,N_9895,N_6715);
nor U13645 (N_13645,N_7934,N_8824);
xnor U13646 (N_13646,N_8090,N_7612);
or U13647 (N_13647,N_8252,N_9090);
nand U13648 (N_13648,N_5757,N_8406);
nand U13649 (N_13649,N_5166,N_7608);
and U13650 (N_13650,N_6081,N_5664);
or U13651 (N_13651,N_9955,N_6749);
nor U13652 (N_13652,N_9689,N_9747);
nor U13653 (N_13653,N_5608,N_7953);
or U13654 (N_13654,N_7433,N_9804);
and U13655 (N_13655,N_5056,N_8063);
and U13656 (N_13656,N_7633,N_5389);
or U13657 (N_13657,N_6218,N_5576);
nor U13658 (N_13658,N_9349,N_7574);
xor U13659 (N_13659,N_9934,N_5263);
and U13660 (N_13660,N_6237,N_9879);
and U13661 (N_13661,N_6729,N_9740);
or U13662 (N_13662,N_7036,N_9128);
and U13663 (N_13663,N_8403,N_6762);
nor U13664 (N_13664,N_7754,N_5750);
or U13665 (N_13665,N_5219,N_6847);
or U13666 (N_13666,N_5779,N_6954);
or U13667 (N_13667,N_5034,N_8711);
nand U13668 (N_13668,N_5117,N_6464);
nand U13669 (N_13669,N_8901,N_7647);
or U13670 (N_13670,N_7238,N_9006);
or U13671 (N_13671,N_5779,N_6624);
or U13672 (N_13672,N_8862,N_9401);
and U13673 (N_13673,N_9877,N_5304);
nor U13674 (N_13674,N_8938,N_7457);
or U13675 (N_13675,N_6496,N_6799);
nor U13676 (N_13676,N_6599,N_5824);
or U13677 (N_13677,N_7679,N_7583);
nand U13678 (N_13678,N_5888,N_8519);
and U13679 (N_13679,N_9924,N_7230);
xnor U13680 (N_13680,N_6237,N_8625);
nand U13681 (N_13681,N_5824,N_5595);
nand U13682 (N_13682,N_9258,N_9676);
nand U13683 (N_13683,N_7889,N_9705);
or U13684 (N_13684,N_7635,N_7392);
or U13685 (N_13685,N_8619,N_9848);
nor U13686 (N_13686,N_7504,N_6991);
nand U13687 (N_13687,N_6873,N_9723);
xnor U13688 (N_13688,N_9250,N_9866);
and U13689 (N_13689,N_9086,N_8236);
and U13690 (N_13690,N_9867,N_5952);
or U13691 (N_13691,N_8459,N_8936);
or U13692 (N_13692,N_8221,N_5030);
and U13693 (N_13693,N_5066,N_8672);
or U13694 (N_13694,N_6360,N_8193);
nand U13695 (N_13695,N_7750,N_9645);
or U13696 (N_13696,N_5262,N_8876);
and U13697 (N_13697,N_8001,N_5962);
and U13698 (N_13698,N_8984,N_8205);
or U13699 (N_13699,N_6245,N_6769);
nor U13700 (N_13700,N_6451,N_8807);
nand U13701 (N_13701,N_5294,N_5055);
or U13702 (N_13702,N_6039,N_7300);
and U13703 (N_13703,N_7152,N_6861);
or U13704 (N_13704,N_5228,N_8012);
nor U13705 (N_13705,N_9597,N_9544);
and U13706 (N_13706,N_5166,N_9195);
and U13707 (N_13707,N_8722,N_7326);
or U13708 (N_13708,N_6685,N_8299);
nand U13709 (N_13709,N_5544,N_6926);
nand U13710 (N_13710,N_7534,N_8065);
or U13711 (N_13711,N_8860,N_7214);
and U13712 (N_13712,N_6325,N_6019);
nor U13713 (N_13713,N_5267,N_6969);
nand U13714 (N_13714,N_7670,N_9832);
or U13715 (N_13715,N_6903,N_6890);
nand U13716 (N_13716,N_7621,N_9394);
nor U13717 (N_13717,N_7512,N_6885);
or U13718 (N_13718,N_7149,N_5249);
and U13719 (N_13719,N_6379,N_9317);
nor U13720 (N_13720,N_7271,N_9447);
or U13721 (N_13721,N_6874,N_7096);
nand U13722 (N_13722,N_8946,N_8645);
and U13723 (N_13723,N_9381,N_9837);
xor U13724 (N_13724,N_7745,N_8014);
nand U13725 (N_13725,N_7834,N_6174);
xnor U13726 (N_13726,N_8807,N_8055);
and U13727 (N_13727,N_9810,N_9280);
nor U13728 (N_13728,N_5593,N_8433);
xor U13729 (N_13729,N_9302,N_7655);
xnor U13730 (N_13730,N_6060,N_7623);
and U13731 (N_13731,N_6596,N_6283);
nand U13732 (N_13732,N_5730,N_6912);
or U13733 (N_13733,N_8833,N_7976);
or U13734 (N_13734,N_6002,N_9539);
or U13735 (N_13735,N_9709,N_9456);
or U13736 (N_13736,N_9247,N_6777);
or U13737 (N_13737,N_9030,N_7945);
nand U13738 (N_13738,N_5638,N_6230);
xor U13739 (N_13739,N_7629,N_6429);
and U13740 (N_13740,N_5912,N_6629);
nand U13741 (N_13741,N_5815,N_7534);
xor U13742 (N_13742,N_9391,N_9813);
xor U13743 (N_13743,N_6143,N_7186);
nand U13744 (N_13744,N_8602,N_5927);
nor U13745 (N_13745,N_8745,N_7529);
nor U13746 (N_13746,N_8851,N_6897);
nor U13747 (N_13747,N_8596,N_8972);
xor U13748 (N_13748,N_8171,N_8497);
and U13749 (N_13749,N_7818,N_6396);
nand U13750 (N_13750,N_7684,N_6622);
and U13751 (N_13751,N_5402,N_8129);
and U13752 (N_13752,N_6829,N_7151);
or U13753 (N_13753,N_5478,N_9845);
or U13754 (N_13754,N_5887,N_5473);
nand U13755 (N_13755,N_7073,N_9598);
xnor U13756 (N_13756,N_6912,N_7595);
and U13757 (N_13757,N_7671,N_6219);
or U13758 (N_13758,N_7368,N_6488);
nand U13759 (N_13759,N_8192,N_9165);
nand U13760 (N_13760,N_9527,N_9430);
nor U13761 (N_13761,N_7261,N_6406);
nand U13762 (N_13762,N_7990,N_6248);
or U13763 (N_13763,N_5822,N_6281);
nand U13764 (N_13764,N_6526,N_7006);
nand U13765 (N_13765,N_9318,N_8365);
and U13766 (N_13766,N_9790,N_9401);
nand U13767 (N_13767,N_9499,N_9104);
nor U13768 (N_13768,N_7146,N_7174);
and U13769 (N_13769,N_9371,N_9681);
nand U13770 (N_13770,N_6392,N_7822);
and U13771 (N_13771,N_7168,N_7905);
nor U13772 (N_13772,N_7456,N_8622);
or U13773 (N_13773,N_8299,N_9389);
nand U13774 (N_13774,N_6141,N_8431);
and U13775 (N_13775,N_5225,N_5232);
nor U13776 (N_13776,N_9084,N_9487);
nor U13777 (N_13777,N_9126,N_6016);
nor U13778 (N_13778,N_8195,N_8012);
or U13779 (N_13779,N_6060,N_6202);
and U13780 (N_13780,N_8250,N_6601);
and U13781 (N_13781,N_6091,N_6212);
or U13782 (N_13782,N_8935,N_6893);
and U13783 (N_13783,N_9069,N_7043);
or U13784 (N_13784,N_8942,N_7250);
and U13785 (N_13785,N_5521,N_5280);
xnor U13786 (N_13786,N_8556,N_9787);
nand U13787 (N_13787,N_8129,N_7443);
nand U13788 (N_13788,N_5490,N_8223);
or U13789 (N_13789,N_7626,N_5732);
nand U13790 (N_13790,N_5416,N_7892);
xnor U13791 (N_13791,N_5475,N_9543);
xnor U13792 (N_13792,N_6665,N_7149);
nor U13793 (N_13793,N_8343,N_6151);
nor U13794 (N_13794,N_7470,N_5861);
nor U13795 (N_13795,N_8901,N_7296);
nor U13796 (N_13796,N_6271,N_8277);
nand U13797 (N_13797,N_5799,N_9191);
or U13798 (N_13798,N_6170,N_6341);
nor U13799 (N_13799,N_6633,N_5118);
nor U13800 (N_13800,N_8309,N_7949);
nand U13801 (N_13801,N_9508,N_7599);
nor U13802 (N_13802,N_5207,N_6316);
nand U13803 (N_13803,N_6382,N_5977);
or U13804 (N_13804,N_5280,N_5625);
or U13805 (N_13805,N_6697,N_7365);
nor U13806 (N_13806,N_8222,N_5478);
or U13807 (N_13807,N_7393,N_6536);
nand U13808 (N_13808,N_9137,N_8053);
and U13809 (N_13809,N_6167,N_7386);
and U13810 (N_13810,N_5715,N_9157);
nor U13811 (N_13811,N_6657,N_5309);
nor U13812 (N_13812,N_9681,N_5565);
and U13813 (N_13813,N_6554,N_9894);
nor U13814 (N_13814,N_8259,N_9288);
or U13815 (N_13815,N_7554,N_5850);
nor U13816 (N_13816,N_5521,N_5245);
nand U13817 (N_13817,N_5392,N_6269);
nand U13818 (N_13818,N_9954,N_5192);
nor U13819 (N_13819,N_7967,N_8340);
xor U13820 (N_13820,N_9145,N_9556);
or U13821 (N_13821,N_6608,N_7612);
and U13822 (N_13822,N_6124,N_7284);
or U13823 (N_13823,N_8401,N_5856);
nand U13824 (N_13824,N_6001,N_5889);
nand U13825 (N_13825,N_6295,N_8851);
nor U13826 (N_13826,N_9281,N_5812);
or U13827 (N_13827,N_5307,N_9308);
or U13828 (N_13828,N_7330,N_7832);
and U13829 (N_13829,N_5650,N_9408);
xnor U13830 (N_13830,N_8323,N_8664);
xnor U13831 (N_13831,N_5931,N_6923);
or U13832 (N_13832,N_7416,N_6170);
and U13833 (N_13833,N_7977,N_7653);
or U13834 (N_13834,N_7488,N_5433);
nand U13835 (N_13835,N_8766,N_8419);
or U13836 (N_13836,N_6724,N_6040);
or U13837 (N_13837,N_6318,N_8011);
nand U13838 (N_13838,N_7729,N_6380);
and U13839 (N_13839,N_7477,N_7074);
and U13840 (N_13840,N_5310,N_7267);
xor U13841 (N_13841,N_9999,N_5220);
nand U13842 (N_13842,N_7167,N_6000);
nand U13843 (N_13843,N_9849,N_7166);
or U13844 (N_13844,N_9993,N_6910);
nor U13845 (N_13845,N_8410,N_6571);
and U13846 (N_13846,N_6899,N_9226);
nor U13847 (N_13847,N_6501,N_6493);
or U13848 (N_13848,N_6307,N_6184);
nand U13849 (N_13849,N_5672,N_8072);
or U13850 (N_13850,N_6245,N_9938);
nor U13851 (N_13851,N_6258,N_9341);
and U13852 (N_13852,N_6570,N_8550);
nand U13853 (N_13853,N_9118,N_5535);
nand U13854 (N_13854,N_6452,N_9761);
and U13855 (N_13855,N_8535,N_7830);
and U13856 (N_13856,N_5892,N_9643);
xor U13857 (N_13857,N_8723,N_8798);
nor U13858 (N_13858,N_6649,N_5004);
xnor U13859 (N_13859,N_7765,N_6861);
nor U13860 (N_13860,N_9339,N_5876);
nor U13861 (N_13861,N_5006,N_5474);
nor U13862 (N_13862,N_9228,N_7481);
or U13863 (N_13863,N_8041,N_6588);
or U13864 (N_13864,N_6616,N_5566);
or U13865 (N_13865,N_9648,N_6877);
nor U13866 (N_13866,N_7561,N_9109);
nor U13867 (N_13867,N_5307,N_7919);
and U13868 (N_13868,N_5112,N_6929);
nor U13869 (N_13869,N_9492,N_8569);
or U13870 (N_13870,N_9943,N_5102);
nand U13871 (N_13871,N_9089,N_5422);
and U13872 (N_13872,N_7844,N_6249);
or U13873 (N_13873,N_8052,N_8511);
nor U13874 (N_13874,N_7914,N_5175);
xor U13875 (N_13875,N_7139,N_8392);
nand U13876 (N_13876,N_6615,N_8173);
and U13877 (N_13877,N_7830,N_7938);
xnor U13878 (N_13878,N_8829,N_8212);
nor U13879 (N_13879,N_5268,N_7529);
and U13880 (N_13880,N_5436,N_9009);
nand U13881 (N_13881,N_7471,N_7107);
nand U13882 (N_13882,N_5843,N_5299);
or U13883 (N_13883,N_7553,N_8235);
or U13884 (N_13884,N_7199,N_7450);
nand U13885 (N_13885,N_6687,N_6682);
or U13886 (N_13886,N_5693,N_8660);
and U13887 (N_13887,N_6028,N_6667);
xnor U13888 (N_13888,N_6205,N_7233);
or U13889 (N_13889,N_6192,N_5405);
or U13890 (N_13890,N_5784,N_9110);
or U13891 (N_13891,N_8147,N_9905);
xor U13892 (N_13892,N_7809,N_8540);
and U13893 (N_13893,N_6867,N_8459);
nor U13894 (N_13894,N_9967,N_7174);
xnor U13895 (N_13895,N_6503,N_9015);
nand U13896 (N_13896,N_7667,N_6778);
nor U13897 (N_13897,N_6011,N_7115);
nor U13898 (N_13898,N_6797,N_6470);
nand U13899 (N_13899,N_8426,N_7732);
and U13900 (N_13900,N_5178,N_5132);
nand U13901 (N_13901,N_6049,N_6681);
nor U13902 (N_13902,N_8765,N_9521);
nand U13903 (N_13903,N_7318,N_6142);
or U13904 (N_13904,N_8442,N_5009);
and U13905 (N_13905,N_8884,N_5919);
nor U13906 (N_13906,N_7660,N_8420);
and U13907 (N_13907,N_8355,N_5333);
and U13908 (N_13908,N_9271,N_6534);
nor U13909 (N_13909,N_5238,N_9316);
or U13910 (N_13910,N_5046,N_6728);
xor U13911 (N_13911,N_9488,N_5249);
and U13912 (N_13912,N_5895,N_9403);
xor U13913 (N_13913,N_8447,N_8522);
nand U13914 (N_13914,N_5986,N_6554);
or U13915 (N_13915,N_8390,N_7475);
nor U13916 (N_13916,N_7685,N_7895);
nor U13917 (N_13917,N_8733,N_9893);
or U13918 (N_13918,N_8015,N_9401);
nor U13919 (N_13919,N_5396,N_7049);
nand U13920 (N_13920,N_9460,N_8387);
xnor U13921 (N_13921,N_5338,N_5488);
and U13922 (N_13922,N_8225,N_7259);
or U13923 (N_13923,N_5947,N_7417);
nand U13924 (N_13924,N_9176,N_6327);
or U13925 (N_13925,N_7185,N_5825);
and U13926 (N_13926,N_9937,N_8398);
xnor U13927 (N_13927,N_7329,N_9505);
nor U13928 (N_13928,N_6054,N_5616);
nand U13929 (N_13929,N_7616,N_5433);
nand U13930 (N_13930,N_8227,N_6969);
nand U13931 (N_13931,N_9877,N_6535);
nand U13932 (N_13932,N_8432,N_8365);
nor U13933 (N_13933,N_6853,N_8733);
xor U13934 (N_13934,N_7334,N_6367);
or U13935 (N_13935,N_6746,N_9911);
nand U13936 (N_13936,N_6760,N_5221);
and U13937 (N_13937,N_5305,N_5960);
nand U13938 (N_13938,N_9581,N_7268);
and U13939 (N_13939,N_6938,N_9856);
nor U13940 (N_13940,N_9932,N_9180);
and U13941 (N_13941,N_5269,N_5526);
nor U13942 (N_13942,N_8239,N_6653);
xor U13943 (N_13943,N_6873,N_6025);
nand U13944 (N_13944,N_9875,N_7569);
nor U13945 (N_13945,N_6462,N_9570);
and U13946 (N_13946,N_5380,N_9750);
and U13947 (N_13947,N_5245,N_9984);
xor U13948 (N_13948,N_7189,N_7325);
nand U13949 (N_13949,N_6167,N_7638);
or U13950 (N_13950,N_8400,N_7732);
nand U13951 (N_13951,N_9221,N_6628);
and U13952 (N_13952,N_9983,N_7176);
and U13953 (N_13953,N_5409,N_8539);
and U13954 (N_13954,N_7703,N_9344);
nor U13955 (N_13955,N_8461,N_5333);
nand U13956 (N_13956,N_9285,N_5508);
nor U13957 (N_13957,N_7215,N_6870);
and U13958 (N_13958,N_7730,N_5087);
nor U13959 (N_13959,N_8599,N_5427);
or U13960 (N_13960,N_7868,N_8502);
and U13961 (N_13961,N_7646,N_8787);
nor U13962 (N_13962,N_8356,N_8800);
or U13963 (N_13963,N_6738,N_5352);
or U13964 (N_13964,N_5763,N_9909);
or U13965 (N_13965,N_8616,N_6182);
nor U13966 (N_13966,N_9961,N_9604);
and U13967 (N_13967,N_6097,N_8625);
nor U13968 (N_13968,N_5263,N_8388);
nor U13969 (N_13969,N_9934,N_9076);
and U13970 (N_13970,N_8054,N_6695);
nand U13971 (N_13971,N_7395,N_7782);
xor U13972 (N_13972,N_5228,N_8949);
or U13973 (N_13973,N_9167,N_8958);
and U13974 (N_13974,N_9545,N_6132);
and U13975 (N_13975,N_8912,N_7958);
or U13976 (N_13976,N_7845,N_6399);
or U13977 (N_13977,N_8792,N_8995);
nor U13978 (N_13978,N_5217,N_8444);
and U13979 (N_13979,N_8189,N_5063);
or U13980 (N_13980,N_9669,N_6287);
and U13981 (N_13981,N_8108,N_9894);
nand U13982 (N_13982,N_7002,N_9588);
xor U13983 (N_13983,N_8100,N_9827);
nor U13984 (N_13984,N_7743,N_7523);
or U13985 (N_13985,N_8775,N_5405);
nor U13986 (N_13986,N_8096,N_9391);
xnor U13987 (N_13987,N_8164,N_5869);
or U13988 (N_13988,N_8177,N_8809);
and U13989 (N_13989,N_6286,N_9027);
and U13990 (N_13990,N_5420,N_8319);
and U13991 (N_13991,N_6750,N_7504);
and U13992 (N_13992,N_5624,N_9061);
nand U13993 (N_13993,N_6072,N_9755);
and U13994 (N_13994,N_7817,N_8301);
xor U13995 (N_13995,N_6289,N_7605);
nor U13996 (N_13996,N_7441,N_9978);
and U13997 (N_13997,N_6873,N_7105);
and U13998 (N_13998,N_5239,N_5725);
nand U13999 (N_13999,N_8460,N_5177);
nor U14000 (N_14000,N_5122,N_5869);
and U14001 (N_14001,N_8363,N_5325);
or U14002 (N_14002,N_6427,N_5540);
nand U14003 (N_14003,N_9846,N_9226);
or U14004 (N_14004,N_6230,N_8501);
nand U14005 (N_14005,N_6759,N_9077);
and U14006 (N_14006,N_9602,N_5465);
and U14007 (N_14007,N_7749,N_7095);
xnor U14008 (N_14008,N_8889,N_6556);
xnor U14009 (N_14009,N_8924,N_9254);
or U14010 (N_14010,N_8738,N_9479);
nor U14011 (N_14011,N_9750,N_6955);
nor U14012 (N_14012,N_9838,N_6676);
and U14013 (N_14013,N_7796,N_8263);
nor U14014 (N_14014,N_6876,N_5694);
nand U14015 (N_14015,N_6254,N_6461);
nand U14016 (N_14016,N_6446,N_5484);
nor U14017 (N_14017,N_7706,N_5474);
and U14018 (N_14018,N_6816,N_6261);
and U14019 (N_14019,N_5392,N_8410);
or U14020 (N_14020,N_6528,N_6465);
and U14021 (N_14021,N_8491,N_9245);
nor U14022 (N_14022,N_8939,N_5083);
xor U14023 (N_14023,N_5282,N_9936);
xnor U14024 (N_14024,N_5405,N_8277);
nand U14025 (N_14025,N_5617,N_5737);
nand U14026 (N_14026,N_5042,N_5212);
nand U14027 (N_14027,N_7101,N_9386);
and U14028 (N_14028,N_9568,N_9131);
and U14029 (N_14029,N_7201,N_5541);
nor U14030 (N_14030,N_8843,N_6017);
nor U14031 (N_14031,N_6218,N_8656);
and U14032 (N_14032,N_5097,N_5445);
nand U14033 (N_14033,N_5340,N_8043);
and U14034 (N_14034,N_6349,N_7709);
nand U14035 (N_14035,N_8890,N_5462);
nand U14036 (N_14036,N_6858,N_9124);
xor U14037 (N_14037,N_9642,N_5540);
or U14038 (N_14038,N_6831,N_5378);
or U14039 (N_14039,N_5487,N_8214);
xor U14040 (N_14040,N_8486,N_6710);
or U14041 (N_14041,N_6211,N_6764);
nand U14042 (N_14042,N_6617,N_6352);
and U14043 (N_14043,N_5392,N_8385);
xnor U14044 (N_14044,N_6990,N_6119);
or U14045 (N_14045,N_8894,N_9085);
nand U14046 (N_14046,N_6777,N_5238);
and U14047 (N_14047,N_9466,N_9874);
nand U14048 (N_14048,N_7484,N_5431);
or U14049 (N_14049,N_6946,N_7342);
nand U14050 (N_14050,N_7983,N_9425);
nor U14051 (N_14051,N_9033,N_6741);
and U14052 (N_14052,N_7026,N_8235);
nand U14053 (N_14053,N_9292,N_5755);
nor U14054 (N_14054,N_8883,N_7276);
nor U14055 (N_14055,N_6175,N_5779);
nand U14056 (N_14056,N_9939,N_9401);
and U14057 (N_14057,N_6435,N_7493);
xnor U14058 (N_14058,N_7436,N_9963);
xnor U14059 (N_14059,N_5224,N_8056);
or U14060 (N_14060,N_9429,N_9657);
nor U14061 (N_14061,N_6603,N_5995);
xor U14062 (N_14062,N_5704,N_9533);
nor U14063 (N_14063,N_5459,N_6699);
or U14064 (N_14064,N_8625,N_6415);
nand U14065 (N_14065,N_9755,N_7639);
and U14066 (N_14066,N_7771,N_8403);
nand U14067 (N_14067,N_6942,N_9645);
nor U14068 (N_14068,N_8442,N_7750);
or U14069 (N_14069,N_6188,N_6348);
nand U14070 (N_14070,N_9356,N_8327);
or U14071 (N_14071,N_5052,N_7135);
nand U14072 (N_14072,N_7514,N_9402);
xnor U14073 (N_14073,N_5099,N_7585);
or U14074 (N_14074,N_7253,N_5951);
nor U14075 (N_14075,N_6963,N_6478);
and U14076 (N_14076,N_6772,N_8701);
nand U14077 (N_14077,N_6732,N_6562);
or U14078 (N_14078,N_7917,N_6408);
nor U14079 (N_14079,N_7218,N_8917);
or U14080 (N_14080,N_5932,N_6712);
or U14081 (N_14081,N_9240,N_7806);
nand U14082 (N_14082,N_9250,N_9289);
nand U14083 (N_14083,N_7107,N_5679);
or U14084 (N_14084,N_6881,N_7508);
nand U14085 (N_14085,N_7034,N_9671);
nor U14086 (N_14086,N_8578,N_9442);
xor U14087 (N_14087,N_9777,N_6345);
or U14088 (N_14088,N_7958,N_9602);
nor U14089 (N_14089,N_6978,N_5507);
nand U14090 (N_14090,N_9914,N_8060);
or U14091 (N_14091,N_9968,N_7339);
or U14092 (N_14092,N_8996,N_8682);
nor U14093 (N_14093,N_7160,N_8321);
and U14094 (N_14094,N_7316,N_8664);
or U14095 (N_14095,N_8618,N_6915);
nand U14096 (N_14096,N_9731,N_9052);
nor U14097 (N_14097,N_9958,N_9750);
and U14098 (N_14098,N_9599,N_6477);
and U14099 (N_14099,N_5528,N_5643);
and U14100 (N_14100,N_5151,N_8732);
or U14101 (N_14101,N_5783,N_8711);
nor U14102 (N_14102,N_8139,N_9422);
or U14103 (N_14103,N_7816,N_9852);
nand U14104 (N_14104,N_7757,N_7776);
nand U14105 (N_14105,N_8137,N_6976);
nand U14106 (N_14106,N_7356,N_6864);
and U14107 (N_14107,N_6286,N_7442);
nand U14108 (N_14108,N_7362,N_6986);
nor U14109 (N_14109,N_9919,N_6481);
xnor U14110 (N_14110,N_7728,N_8138);
nor U14111 (N_14111,N_7558,N_5044);
and U14112 (N_14112,N_8863,N_8977);
and U14113 (N_14113,N_5774,N_8912);
or U14114 (N_14114,N_6613,N_7575);
nand U14115 (N_14115,N_7685,N_7571);
nand U14116 (N_14116,N_8763,N_9633);
and U14117 (N_14117,N_5419,N_7159);
nand U14118 (N_14118,N_9676,N_9661);
xnor U14119 (N_14119,N_9853,N_9467);
nor U14120 (N_14120,N_5068,N_9707);
xnor U14121 (N_14121,N_5348,N_8849);
nand U14122 (N_14122,N_6571,N_7685);
nor U14123 (N_14123,N_9955,N_7842);
nor U14124 (N_14124,N_6388,N_8110);
or U14125 (N_14125,N_6932,N_9664);
or U14126 (N_14126,N_8962,N_5973);
or U14127 (N_14127,N_9404,N_6674);
and U14128 (N_14128,N_7379,N_5186);
and U14129 (N_14129,N_7362,N_8535);
or U14130 (N_14130,N_8058,N_6792);
xor U14131 (N_14131,N_7465,N_6010);
nand U14132 (N_14132,N_9614,N_8761);
nand U14133 (N_14133,N_8794,N_7151);
nor U14134 (N_14134,N_7651,N_9098);
nand U14135 (N_14135,N_5525,N_5500);
or U14136 (N_14136,N_8980,N_7481);
nand U14137 (N_14137,N_9649,N_6125);
nor U14138 (N_14138,N_6713,N_9877);
nor U14139 (N_14139,N_6432,N_6881);
or U14140 (N_14140,N_8925,N_6303);
nor U14141 (N_14141,N_8477,N_8540);
and U14142 (N_14142,N_8162,N_8755);
or U14143 (N_14143,N_8190,N_5308);
or U14144 (N_14144,N_9872,N_6358);
nor U14145 (N_14145,N_9938,N_6083);
and U14146 (N_14146,N_5076,N_8135);
and U14147 (N_14147,N_6831,N_7466);
xor U14148 (N_14148,N_6240,N_7667);
nor U14149 (N_14149,N_8114,N_7034);
and U14150 (N_14150,N_6684,N_7800);
nand U14151 (N_14151,N_6394,N_8726);
xor U14152 (N_14152,N_8025,N_7659);
or U14153 (N_14153,N_8892,N_9706);
nor U14154 (N_14154,N_7088,N_6859);
xnor U14155 (N_14155,N_5517,N_9741);
nor U14156 (N_14156,N_6954,N_7605);
nor U14157 (N_14157,N_6149,N_8076);
or U14158 (N_14158,N_5531,N_5024);
nand U14159 (N_14159,N_7932,N_8720);
and U14160 (N_14160,N_7705,N_7926);
and U14161 (N_14161,N_9519,N_8724);
nor U14162 (N_14162,N_8000,N_5214);
or U14163 (N_14163,N_7772,N_7750);
or U14164 (N_14164,N_6466,N_9788);
nand U14165 (N_14165,N_9833,N_5056);
or U14166 (N_14166,N_6739,N_7159);
and U14167 (N_14167,N_7217,N_7319);
xnor U14168 (N_14168,N_6319,N_8329);
nor U14169 (N_14169,N_6946,N_5244);
nor U14170 (N_14170,N_6895,N_8555);
and U14171 (N_14171,N_7648,N_9372);
nor U14172 (N_14172,N_7970,N_9978);
or U14173 (N_14173,N_7460,N_5779);
or U14174 (N_14174,N_8514,N_8517);
nor U14175 (N_14175,N_6411,N_6946);
xnor U14176 (N_14176,N_8940,N_6032);
and U14177 (N_14177,N_6068,N_6407);
or U14178 (N_14178,N_8322,N_5458);
or U14179 (N_14179,N_9170,N_9370);
and U14180 (N_14180,N_7705,N_6674);
or U14181 (N_14181,N_7783,N_8789);
nand U14182 (N_14182,N_7831,N_8764);
nand U14183 (N_14183,N_7653,N_5222);
nand U14184 (N_14184,N_5872,N_7099);
nand U14185 (N_14185,N_5478,N_5711);
nand U14186 (N_14186,N_8903,N_6914);
or U14187 (N_14187,N_5241,N_7905);
or U14188 (N_14188,N_8011,N_6340);
and U14189 (N_14189,N_9480,N_6493);
nand U14190 (N_14190,N_7765,N_8306);
nand U14191 (N_14191,N_9734,N_9223);
nand U14192 (N_14192,N_6768,N_8459);
or U14193 (N_14193,N_8532,N_9939);
nor U14194 (N_14194,N_8990,N_8816);
nor U14195 (N_14195,N_6740,N_5278);
and U14196 (N_14196,N_9633,N_6753);
nand U14197 (N_14197,N_9569,N_6321);
nand U14198 (N_14198,N_9873,N_7627);
nand U14199 (N_14199,N_5406,N_5288);
nor U14200 (N_14200,N_8513,N_9412);
or U14201 (N_14201,N_6723,N_6289);
xor U14202 (N_14202,N_7914,N_5436);
nor U14203 (N_14203,N_9144,N_7396);
xnor U14204 (N_14204,N_8194,N_9443);
and U14205 (N_14205,N_6600,N_8494);
and U14206 (N_14206,N_7156,N_5288);
and U14207 (N_14207,N_5681,N_5703);
or U14208 (N_14208,N_6706,N_8750);
xor U14209 (N_14209,N_9866,N_9414);
or U14210 (N_14210,N_5757,N_6898);
and U14211 (N_14211,N_8616,N_7094);
nand U14212 (N_14212,N_7306,N_9045);
nand U14213 (N_14213,N_5665,N_6895);
and U14214 (N_14214,N_9120,N_5786);
and U14215 (N_14215,N_8420,N_8937);
nand U14216 (N_14216,N_6200,N_8539);
nor U14217 (N_14217,N_6643,N_8716);
nor U14218 (N_14218,N_7384,N_5256);
nor U14219 (N_14219,N_7189,N_6504);
xnor U14220 (N_14220,N_9770,N_5014);
or U14221 (N_14221,N_9252,N_6065);
nand U14222 (N_14222,N_6596,N_8313);
or U14223 (N_14223,N_5351,N_9524);
nor U14224 (N_14224,N_8750,N_7880);
nor U14225 (N_14225,N_6814,N_6526);
or U14226 (N_14226,N_7756,N_7976);
nor U14227 (N_14227,N_6954,N_8557);
nor U14228 (N_14228,N_8368,N_9393);
or U14229 (N_14229,N_8664,N_5000);
nand U14230 (N_14230,N_8664,N_6748);
and U14231 (N_14231,N_5542,N_6076);
nand U14232 (N_14232,N_5221,N_6530);
or U14233 (N_14233,N_9440,N_6595);
nand U14234 (N_14234,N_9692,N_5258);
and U14235 (N_14235,N_8735,N_7857);
and U14236 (N_14236,N_6891,N_6523);
nor U14237 (N_14237,N_8468,N_6612);
and U14238 (N_14238,N_5572,N_9217);
or U14239 (N_14239,N_8736,N_8751);
and U14240 (N_14240,N_5763,N_9788);
nor U14241 (N_14241,N_7900,N_8446);
nor U14242 (N_14242,N_5137,N_9045);
nor U14243 (N_14243,N_9190,N_6123);
or U14244 (N_14244,N_7730,N_8090);
or U14245 (N_14245,N_6769,N_6573);
and U14246 (N_14246,N_7750,N_7020);
or U14247 (N_14247,N_5792,N_7753);
nor U14248 (N_14248,N_7228,N_5734);
nor U14249 (N_14249,N_9170,N_9130);
nor U14250 (N_14250,N_8493,N_6047);
nor U14251 (N_14251,N_7091,N_9591);
or U14252 (N_14252,N_5396,N_7738);
or U14253 (N_14253,N_6601,N_7406);
and U14254 (N_14254,N_8415,N_9788);
nor U14255 (N_14255,N_7575,N_8292);
xnor U14256 (N_14256,N_6575,N_5496);
nor U14257 (N_14257,N_8759,N_7839);
and U14258 (N_14258,N_5764,N_5299);
or U14259 (N_14259,N_7782,N_9949);
and U14260 (N_14260,N_5500,N_9389);
nor U14261 (N_14261,N_8830,N_7576);
xnor U14262 (N_14262,N_8913,N_8215);
or U14263 (N_14263,N_8588,N_6437);
and U14264 (N_14264,N_7404,N_7915);
and U14265 (N_14265,N_9382,N_5629);
or U14266 (N_14266,N_8069,N_7943);
xor U14267 (N_14267,N_8637,N_9135);
xor U14268 (N_14268,N_5376,N_8312);
or U14269 (N_14269,N_6342,N_6542);
nand U14270 (N_14270,N_9189,N_8677);
xnor U14271 (N_14271,N_7851,N_5309);
and U14272 (N_14272,N_9432,N_8177);
xor U14273 (N_14273,N_7543,N_8235);
nand U14274 (N_14274,N_5978,N_7209);
and U14275 (N_14275,N_7314,N_6354);
nand U14276 (N_14276,N_8606,N_5897);
nand U14277 (N_14277,N_6244,N_9534);
or U14278 (N_14278,N_6206,N_8555);
nand U14279 (N_14279,N_6923,N_7919);
xor U14280 (N_14280,N_6647,N_8945);
nand U14281 (N_14281,N_8807,N_5065);
nor U14282 (N_14282,N_5676,N_6948);
or U14283 (N_14283,N_8322,N_7485);
and U14284 (N_14284,N_5578,N_5175);
and U14285 (N_14285,N_5952,N_5928);
nor U14286 (N_14286,N_7699,N_8946);
or U14287 (N_14287,N_6994,N_8330);
and U14288 (N_14288,N_7965,N_9053);
or U14289 (N_14289,N_5938,N_9088);
nand U14290 (N_14290,N_8494,N_6826);
or U14291 (N_14291,N_5137,N_8719);
or U14292 (N_14292,N_6642,N_7699);
nand U14293 (N_14293,N_9303,N_8533);
nor U14294 (N_14294,N_7694,N_9267);
or U14295 (N_14295,N_7432,N_7943);
nor U14296 (N_14296,N_6166,N_7541);
nor U14297 (N_14297,N_5075,N_6662);
or U14298 (N_14298,N_9441,N_9889);
xnor U14299 (N_14299,N_6922,N_7161);
xnor U14300 (N_14300,N_9371,N_9292);
nand U14301 (N_14301,N_5340,N_5592);
or U14302 (N_14302,N_8517,N_5101);
nand U14303 (N_14303,N_7625,N_8614);
and U14304 (N_14304,N_8957,N_9233);
and U14305 (N_14305,N_7650,N_9510);
nor U14306 (N_14306,N_8418,N_9922);
and U14307 (N_14307,N_7742,N_6001);
and U14308 (N_14308,N_5451,N_8766);
xor U14309 (N_14309,N_8884,N_5982);
and U14310 (N_14310,N_9923,N_9236);
and U14311 (N_14311,N_5811,N_7836);
and U14312 (N_14312,N_8546,N_6318);
nand U14313 (N_14313,N_6832,N_5260);
or U14314 (N_14314,N_7348,N_7887);
nor U14315 (N_14315,N_8053,N_8389);
nand U14316 (N_14316,N_6547,N_6418);
or U14317 (N_14317,N_7930,N_8984);
or U14318 (N_14318,N_8069,N_6809);
nand U14319 (N_14319,N_7048,N_5935);
nand U14320 (N_14320,N_9791,N_9305);
nor U14321 (N_14321,N_6526,N_8237);
nor U14322 (N_14322,N_6651,N_5551);
or U14323 (N_14323,N_6719,N_6531);
and U14324 (N_14324,N_7376,N_6630);
or U14325 (N_14325,N_6058,N_5512);
or U14326 (N_14326,N_6955,N_5141);
and U14327 (N_14327,N_7910,N_8801);
and U14328 (N_14328,N_8187,N_5224);
nand U14329 (N_14329,N_9000,N_9691);
or U14330 (N_14330,N_8768,N_9944);
nand U14331 (N_14331,N_8565,N_5322);
nand U14332 (N_14332,N_9001,N_9046);
and U14333 (N_14333,N_5958,N_5206);
nand U14334 (N_14334,N_8752,N_9315);
nand U14335 (N_14335,N_6293,N_6480);
or U14336 (N_14336,N_9192,N_8368);
xor U14337 (N_14337,N_8260,N_7270);
or U14338 (N_14338,N_8750,N_9667);
and U14339 (N_14339,N_7477,N_8392);
and U14340 (N_14340,N_9902,N_8669);
nand U14341 (N_14341,N_5903,N_9284);
or U14342 (N_14342,N_6124,N_7315);
nor U14343 (N_14343,N_5036,N_9588);
and U14344 (N_14344,N_5397,N_9701);
nor U14345 (N_14345,N_7831,N_6006);
nand U14346 (N_14346,N_9109,N_5108);
xor U14347 (N_14347,N_5788,N_5933);
and U14348 (N_14348,N_5364,N_9338);
or U14349 (N_14349,N_8364,N_9186);
or U14350 (N_14350,N_7284,N_6989);
nand U14351 (N_14351,N_8856,N_5751);
nor U14352 (N_14352,N_9068,N_6619);
and U14353 (N_14353,N_6392,N_9704);
and U14354 (N_14354,N_9832,N_9651);
nand U14355 (N_14355,N_9049,N_5494);
and U14356 (N_14356,N_8068,N_7997);
or U14357 (N_14357,N_8818,N_8252);
or U14358 (N_14358,N_5718,N_6431);
or U14359 (N_14359,N_7665,N_9099);
nor U14360 (N_14360,N_5624,N_6386);
nor U14361 (N_14361,N_8355,N_5214);
nor U14362 (N_14362,N_8395,N_9461);
nor U14363 (N_14363,N_5905,N_5177);
or U14364 (N_14364,N_8734,N_7491);
xnor U14365 (N_14365,N_8394,N_6205);
nand U14366 (N_14366,N_7093,N_8151);
and U14367 (N_14367,N_6401,N_6756);
nor U14368 (N_14368,N_9200,N_9708);
xor U14369 (N_14369,N_8632,N_5026);
nor U14370 (N_14370,N_6203,N_7244);
nand U14371 (N_14371,N_5130,N_8773);
xor U14372 (N_14372,N_9639,N_6115);
nor U14373 (N_14373,N_7824,N_6697);
xor U14374 (N_14374,N_8690,N_9081);
nand U14375 (N_14375,N_5514,N_8768);
and U14376 (N_14376,N_7363,N_8752);
nand U14377 (N_14377,N_6399,N_5064);
or U14378 (N_14378,N_5663,N_7344);
nand U14379 (N_14379,N_6977,N_8105);
and U14380 (N_14380,N_8602,N_6862);
or U14381 (N_14381,N_8411,N_9400);
or U14382 (N_14382,N_6433,N_5738);
or U14383 (N_14383,N_7681,N_9266);
nor U14384 (N_14384,N_6219,N_5306);
or U14385 (N_14385,N_7627,N_9700);
or U14386 (N_14386,N_5610,N_6222);
xor U14387 (N_14387,N_5317,N_9157);
and U14388 (N_14388,N_6058,N_8916);
xor U14389 (N_14389,N_7956,N_9816);
nor U14390 (N_14390,N_5496,N_9956);
nor U14391 (N_14391,N_7344,N_8850);
or U14392 (N_14392,N_6835,N_9442);
or U14393 (N_14393,N_6827,N_8054);
and U14394 (N_14394,N_9907,N_5058);
nand U14395 (N_14395,N_8899,N_9014);
nor U14396 (N_14396,N_8995,N_5269);
and U14397 (N_14397,N_9205,N_9295);
or U14398 (N_14398,N_5248,N_5332);
nand U14399 (N_14399,N_7252,N_9097);
and U14400 (N_14400,N_5796,N_9802);
nor U14401 (N_14401,N_9432,N_6501);
nor U14402 (N_14402,N_9382,N_5631);
nand U14403 (N_14403,N_8753,N_6384);
nand U14404 (N_14404,N_8268,N_7245);
nand U14405 (N_14405,N_6486,N_9977);
nand U14406 (N_14406,N_9379,N_8116);
or U14407 (N_14407,N_5658,N_6686);
nor U14408 (N_14408,N_6191,N_7783);
nor U14409 (N_14409,N_6551,N_7417);
nand U14410 (N_14410,N_9783,N_6034);
or U14411 (N_14411,N_5350,N_8292);
and U14412 (N_14412,N_6516,N_5089);
nor U14413 (N_14413,N_6333,N_9697);
or U14414 (N_14414,N_5652,N_7799);
or U14415 (N_14415,N_5439,N_6870);
nor U14416 (N_14416,N_9175,N_7597);
nor U14417 (N_14417,N_7735,N_7719);
nor U14418 (N_14418,N_9755,N_5550);
or U14419 (N_14419,N_8938,N_5003);
or U14420 (N_14420,N_5524,N_8084);
nand U14421 (N_14421,N_6355,N_9043);
and U14422 (N_14422,N_6532,N_5597);
nand U14423 (N_14423,N_8929,N_7856);
nand U14424 (N_14424,N_6868,N_5916);
or U14425 (N_14425,N_6812,N_9142);
nand U14426 (N_14426,N_9456,N_8222);
or U14427 (N_14427,N_5480,N_8882);
and U14428 (N_14428,N_9606,N_8238);
xor U14429 (N_14429,N_7351,N_7706);
nor U14430 (N_14430,N_8252,N_6435);
nand U14431 (N_14431,N_9705,N_7211);
nand U14432 (N_14432,N_9321,N_8401);
nand U14433 (N_14433,N_8347,N_5741);
xor U14434 (N_14434,N_7508,N_9836);
and U14435 (N_14435,N_6120,N_7596);
nor U14436 (N_14436,N_9168,N_9814);
or U14437 (N_14437,N_8956,N_9351);
or U14438 (N_14438,N_9037,N_5179);
nand U14439 (N_14439,N_5196,N_8099);
xor U14440 (N_14440,N_6111,N_7725);
and U14441 (N_14441,N_8358,N_5092);
or U14442 (N_14442,N_5934,N_5396);
nand U14443 (N_14443,N_5775,N_6902);
nor U14444 (N_14444,N_8270,N_6567);
nand U14445 (N_14445,N_5772,N_7071);
xor U14446 (N_14446,N_7569,N_7860);
or U14447 (N_14447,N_6628,N_6272);
nand U14448 (N_14448,N_8141,N_7677);
nand U14449 (N_14449,N_5187,N_8722);
nand U14450 (N_14450,N_5508,N_6005);
or U14451 (N_14451,N_5077,N_5504);
or U14452 (N_14452,N_5600,N_5655);
nand U14453 (N_14453,N_8872,N_5250);
or U14454 (N_14454,N_8720,N_7766);
and U14455 (N_14455,N_9707,N_9415);
nor U14456 (N_14456,N_9190,N_9537);
or U14457 (N_14457,N_8438,N_9544);
xor U14458 (N_14458,N_9308,N_7701);
xnor U14459 (N_14459,N_9663,N_7810);
or U14460 (N_14460,N_8209,N_5050);
or U14461 (N_14461,N_7537,N_5637);
or U14462 (N_14462,N_6639,N_9381);
or U14463 (N_14463,N_7348,N_5923);
nor U14464 (N_14464,N_7620,N_5039);
nand U14465 (N_14465,N_5262,N_8887);
or U14466 (N_14466,N_5261,N_9834);
and U14467 (N_14467,N_7189,N_8246);
xnor U14468 (N_14468,N_6695,N_6787);
nand U14469 (N_14469,N_8628,N_7639);
and U14470 (N_14470,N_9232,N_7171);
or U14471 (N_14471,N_6414,N_5229);
and U14472 (N_14472,N_8881,N_5549);
nand U14473 (N_14473,N_6652,N_8356);
and U14474 (N_14474,N_9606,N_5016);
xor U14475 (N_14475,N_9513,N_8730);
and U14476 (N_14476,N_8088,N_9861);
or U14477 (N_14477,N_9276,N_6250);
or U14478 (N_14478,N_5442,N_5250);
or U14479 (N_14479,N_9140,N_7846);
and U14480 (N_14480,N_8870,N_7003);
nand U14481 (N_14481,N_8925,N_8358);
and U14482 (N_14482,N_6241,N_9081);
xnor U14483 (N_14483,N_6693,N_6365);
nor U14484 (N_14484,N_9486,N_8369);
or U14485 (N_14485,N_5187,N_7436);
or U14486 (N_14486,N_7262,N_9289);
or U14487 (N_14487,N_5651,N_8425);
or U14488 (N_14488,N_6960,N_7196);
or U14489 (N_14489,N_9700,N_8386);
nand U14490 (N_14490,N_8429,N_7374);
and U14491 (N_14491,N_6156,N_8632);
nand U14492 (N_14492,N_6110,N_5024);
or U14493 (N_14493,N_7385,N_5174);
or U14494 (N_14494,N_5883,N_9582);
or U14495 (N_14495,N_9734,N_7667);
and U14496 (N_14496,N_8683,N_9221);
nor U14497 (N_14497,N_5102,N_7037);
nor U14498 (N_14498,N_8930,N_6694);
and U14499 (N_14499,N_9428,N_7858);
and U14500 (N_14500,N_7669,N_7487);
xor U14501 (N_14501,N_6600,N_8706);
or U14502 (N_14502,N_9587,N_9537);
nand U14503 (N_14503,N_7321,N_8856);
nand U14504 (N_14504,N_6370,N_9057);
nand U14505 (N_14505,N_8219,N_9732);
or U14506 (N_14506,N_9224,N_8067);
or U14507 (N_14507,N_9080,N_6417);
nor U14508 (N_14508,N_8423,N_9186);
and U14509 (N_14509,N_8609,N_5107);
nand U14510 (N_14510,N_9431,N_5764);
and U14511 (N_14511,N_9998,N_5636);
nand U14512 (N_14512,N_6322,N_8655);
or U14513 (N_14513,N_7007,N_7614);
xor U14514 (N_14514,N_5809,N_6056);
nand U14515 (N_14515,N_9399,N_5800);
or U14516 (N_14516,N_7349,N_9410);
and U14517 (N_14517,N_7490,N_8789);
nor U14518 (N_14518,N_9432,N_7685);
nor U14519 (N_14519,N_8568,N_7013);
or U14520 (N_14520,N_8551,N_9887);
and U14521 (N_14521,N_8833,N_8198);
or U14522 (N_14522,N_6048,N_6165);
or U14523 (N_14523,N_6690,N_8183);
nand U14524 (N_14524,N_7996,N_6528);
nor U14525 (N_14525,N_6784,N_8374);
nor U14526 (N_14526,N_8299,N_6128);
nor U14527 (N_14527,N_8084,N_8790);
or U14528 (N_14528,N_5721,N_7833);
or U14529 (N_14529,N_8145,N_6761);
or U14530 (N_14530,N_8086,N_5433);
nand U14531 (N_14531,N_8661,N_5512);
or U14532 (N_14532,N_8170,N_5551);
or U14533 (N_14533,N_9680,N_5170);
nor U14534 (N_14534,N_9639,N_7647);
xnor U14535 (N_14535,N_5504,N_9286);
and U14536 (N_14536,N_6560,N_8009);
and U14537 (N_14537,N_6449,N_5944);
or U14538 (N_14538,N_8239,N_6166);
or U14539 (N_14539,N_6336,N_6920);
nor U14540 (N_14540,N_7311,N_9616);
nor U14541 (N_14541,N_8966,N_5920);
nand U14542 (N_14542,N_9780,N_9777);
xor U14543 (N_14543,N_9477,N_9366);
nand U14544 (N_14544,N_5448,N_7228);
and U14545 (N_14545,N_7659,N_6467);
nand U14546 (N_14546,N_5742,N_9935);
xor U14547 (N_14547,N_9491,N_6908);
nand U14548 (N_14548,N_8397,N_8886);
or U14549 (N_14549,N_5278,N_7229);
and U14550 (N_14550,N_6791,N_6698);
nand U14551 (N_14551,N_9078,N_7164);
xor U14552 (N_14552,N_6858,N_9519);
and U14553 (N_14553,N_8679,N_8439);
or U14554 (N_14554,N_9793,N_7310);
xor U14555 (N_14555,N_5379,N_5554);
nor U14556 (N_14556,N_7294,N_6717);
nand U14557 (N_14557,N_6212,N_8175);
nand U14558 (N_14558,N_7885,N_5248);
nor U14559 (N_14559,N_9162,N_5169);
or U14560 (N_14560,N_9596,N_7474);
or U14561 (N_14561,N_9197,N_7037);
or U14562 (N_14562,N_9338,N_8563);
and U14563 (N_14563,N_8303,N_5429);
xor U14564 (N_14564,N_9029,N_5603);
nor U14565 (N_14565,N_6479,N_5125);
nand U14566 (N_14566,N_5369,N_7056);
xnor U14567 (N_14567,N_5755,N_9395);
and U14568 (N_14568,N_6805,N_8304);
and U14569 (N_14569,N_9467,N_5813);
or U14570 (N_14570,N_5902,N_5727);
or U14571 (N_14571,N_9426,N_8880);
and U14572 (N_14572,N_7160,N_9012);
nand U14573 (N_14573,N_9873,N_5842);
or U14574 (N_14574,N_8569,N_6819);
nand U14575 (N_14575,N_7287,N_5270);
and U14576 (N_14576,N_7206,N_8263);
or U14577 (N_14577,N_8228,N_8353);
xor U14578 (N_14578,N_8524,N_7753);
nor U14579 (N_14579,N_6818,N_7823);
nand U14580 (N_14580,N_7941,N_9512);
nand U14581 (N_14581,N_9408,N_9215);
xor U14582 (N_14582,N_7309,N_9575);
and U14583 (N_14583,N_8171,N_8503);
or U14584 (N_14584,N_6270,N_5350);
nand U14585 (N_14585,N_8987,N_8285);
or U14586 (N_14586,N_8865,N_7673);
and U14587 (N_14587,N_6053,N_5158);
and U14588 (N_14588,N_8338,N_8290);
nand U14589 (N_14589,N_5700,N_7113);
or U14590 (N_14590,N_7445,N_9782);
nor U14591 (N_14591,N_5890,N_8457);
and U14592 (N_14592,N_8523,N_9784);
and U14593 (N_14593,N_5889,N_5908);
nor U14594 (N_14594,N_5461,N_9030);
nand U14595 (N_14595,N_9935,N_5532);
xnor U14596 (N_14596,N_8207,N_7703);
or U14597 (N_14597,N_5099,N_7752);
and U14598 (N_14598,N_8920,N_6041);
or U14599 (N_14599,N_6913,N_8052);
nand U14600 (N_14600,N_5612,N_8274);
or U14601 (N_14601,N_8628,N_9215);
or U14602 (N_14602,N_6436,N_9002);
nand U14603 (N_14603,N_9262,N_5982);
and U14604 (N_14604,N_9204,N_8245);
xor U14605 (N_14605,N_7937,N_5803);
nand U14606 (N_14606,N_8167,N_8931);
nor U14607 (N_14607,N_8431,N_9733);
nand U14608 (N_14608,N_7242,N_9960);
nand U14609 (N_14609,N_7861,N_5338);
xor U14610 (N_14610,N_6874,N_8321);
nand U14611 (N_14611,N_7034,N_5020);
or U14612 (N_14612,N_9262,N_8740);
and U14613 (N_14613,N_6138,N_9930);
nand U14614 (N_14614,N_5780,N_6409);
or U14615 (N_14615,N_9320,N_5907);
nor U14616 (N_14616,N_9586,N_9133);
and U14617 (N_14617,N_5523,N_8330);
nand U14618 (N_14618,N_5646,N_9595);
and U14619 (N_14619,N_7313,N_6540);
nand U14620 (N_14620,N_9521,N_9101);
and U14621 (N_14621,N_8493,N_7062);
nand U14622 (N_14622,N_5903,N_7429);
xnor U14623 (N_14623,N_7251,N_8873);
nor U14624 (N_14624,N_8012,N_5503);
or U14625 (N_14625,N_6465,N_5270);
and U14626 (N_14626,N_5789,N_6568);
nor U14627 (N_14627,N_8179,N_9885);
nand U14628 (N_14628,N_8805,N_5976);
or U14629 (N_14629,N_9156,N_8811);
or U14630 (N_14630,N_6554,N_6847);
or U14631 (N_14631,N_8343,N_8518);
nor U14632 (N_14632,N_6778,N_7940);
and U14633 (N_14633,N_9393,N_7346);
or U14634 (N_14634,N_9087,N_5007);
nor U14635 (N_14635,N_8292,N_9819);
or U14636 (N_14636,N_7085,N_9280);
nor U14637 (N_14637,N_9873,N_7072);
and U14638 (N_14638,N_8832,N_5319);
or U14639 (N_14639,N_9004,N_8565);
nor U14640 (N_14640,N_6717,N_9014);
nor U14641 (N_14641,N_6532,N_7998);
nand U14642 (N_14642,N_9057,N_7093);
and U14643 (N_14643,N_9518,N_7049);
or U14644 (N_14644,N_8076,N_6733);
and U14645 (N_14645,N_8862,N_6298);
nand U14646 (N_14646,N_6179,N_9833);
nor U14647 (N_14647,N_6987,N_9987);
and U14648 (N_14648,N_8783,N_5042);
and U14649 (N_14649,N_8906,N_6343);
nand U14650 (N_14650,N_7643,N_5618);
nor U14651 (N_14651,N_9778,N_8896);
nor U14652 (N_14652,N_7359,N_5835);
xor U14653 (N_14653,N_9895,N_5275);
nand U14654 (N_14654,N_6808,N_6447);
or U14655 (N_14655,N_7241,N_9338);
nand U14656 (N_14656,N_9443,N_5169);
or U14657 (N_14657,N_6041,N_5441);
and U14658 (N_14658,N_9625,N_6105);
nand U14659 (N_14659,N_6983,N_9533);
nand U14660 (N_14660,N_8128,N_6127);
xor U14661 (N_14661,N_7839,N_8345);
and U14662 (N_14662,N_5504,N_8431);
nor U14663 (N_14663,N_6758,N_5588);
nor U14664 (N_14664,N_9993,N_8362);
nand U14665 (N_14665,N_5161,N_7714);
nand U14666 (N_14666,N_7659,N_6388);
xor U14667 (N_14667,N_6727,N_5249);
and U14668 (N_14668,N_5255,N_5721);
xor U14669 (N_14669,N_8470,N_5182);
or U14670 (N_14670,N_9288,N_6232);
or U14671 (N_14671,N_6259,N_8985);
xor U14672 (N_14672,N_5885,N_5841);
nor U14673 (N_14673,N_7966,N_9147);
and U14674 (N_14674,N_6024,N_6758);
and U14675 (N_14675,N_7891,N_6733);
xor U14676 (N_14676,N_7997,N_8386);
nor U14677 (N_14677,N_6973,N_5553);
and U14678 (N_14678,N_5223,N_7712);
or U14679 (N_14679,N_9503,N_5644);
or U14680 (N_14680,N_8327,N_9776);
nand U14681 (N_14681,N_7251,N_8285);
nand U14682 (N_14682,N_9324,N_9974);
nor U14683 (N_14683,N_8362,N_8200);
nor U14684 (N_14684,N_6375,N_6286);
or U14685 (N_14685,N_8632,N_6263);
nor U14686 (N_14686,N_7640,N_5181);
nor U14687 (N_14687,N_8478,N_5872);
and U14688 (N_14688,N_7757,N_8361);
nor U14689 (N_14689,N_5807,N_6149);
and U14690 (N_14690,N_7544,N_6489);
and U14691 (N_14691,N_5075,N_6023);
and U14692 (N_14692,N_8074,N_6986);
nand U14693 (N_14693,N_8569,N_6017);
and U14694 (N_14694,N_7497,N_8504);
xor U14695 (N_14695,N_8144,N_6400);
and U14696 (N_14696,N_8822,N_5548);
or U14697 (N_14697,N_6954,N_6105);
nand U14698 (N_14698,N_8452,N_9488);
nor U14699 (N_14699,N_5783,N_6676);
nor U14700 (N_14700,N_7765,N_9407);
or U14701 (N_14701,N_7506,N_5320);
or U14702 (N_14702,N_8022,N_8095);
nor U14703 (N_14703,N_7450,N_9692);
and U14704 (N_14704,N_8007,N_9974);
nor U14705 (N_14705,N_8821,N_8866);
or U14706 (N_14706,N_6069,N_8505);
nor U14707 (N_14707,N_7022,N_5203);
nand U14708 (N_14708,N_9149,N_5781);
and U14709 (N_14709,N_8598,N_6002);
nor U14710 (N_14710,N_6309,N_5110);
nor U14711 (N_14711,N_7853,N_9904);
or U14712 (N_14712,N_6523,N_8445);
xnor U14713 (N_14713,N_7766,N_5831);
nand U14714 (N_14714,N_8521,N_7185);
nand U14715 (N_14715,N_7688,N_5279);
or U14716 (N_14716,N_5208,N_7222);
and U14717 (N_14717,N_8773,N_9725);
and U14718 (N_14718,N_5637,N_5693);
xor U14719 (N_14719,N_5045,N_7526);
nor U14720 (N_14720,N_6402,N_8448);
and U14721 (N_14721,N_8772,N_7505);
xor U14722 (N_14722,N_9418,N_9012);
nor U14723 (N_14723,N_5315,N_5057);
nand U14724 (N_14724,N_6186,N_9137);
or U14725 (N_14725,N_7720,N_9386);
or U14726 (N_14726,N_7576,N_7323);
nand U14727 (N_14727,N_6345,N_7531);
or U14728 (N_14728,N_7359,N_6033);
and U14729 (N_14729,N_6663,N_7863);
or U14730 (N_14730,N_5911,N_6736);
and U14731 (N_14731,N_7671,N_7046);
nor U14732 (N_14732,N_5431,N_7841);
nor U14733 (N_14733,N_6083,N_9804);
nor U14734 (N_14734,N_7242,N_5651);
and U14735 (N_14735,N_6592,N_7958);
and U14736 (N_14736,N_9484,N_9637);
and U14737 (N_14737,N_5111,N_8549);
and U14738 (N_14738,N_5777,N_7668);
or U14739 (N_14739,N_7566,N_6414);
nor U14740 (N_14740,N_8296,N_5621);
or U14741 (N_14741,N_9909,N_7227);
or U14742 (N_14742,N_7370,N_8337);
and U14743 (N_14743,N_6746,N_5783);
and U14744 (N_14744,N_7277,N_7454);
nor U14745 (N_14745,N_8992,N_6545);
and U14746 (N_14746,N_7443,N_8911);
or U14747 (N_14747,N_7846,N_8358);
or U14748 (N_14748,N_5761,N_7084);
and U14749 (N_14749,N_5332,N_5976);
nor U14750 (N_14750,N_6748,N_5768);
and U14751 (N_14751,N_7113,N_8486);
nand U14752 (N_14752,N_8204,N_5836);
or U14753 (N_14753,N_8492,N_6562);
and U14754 (N_14754,N_8842,N_9403);
nor U14755 (N_14755,N_9421,N_5818);
or U14756 (N_14756,N_6591,N_5001);
and U14757 (N_14757,N_9080,N_6154);
nand U14758 (N_14758,N_5931,N_8265);
nor U14759 (N_14759,N_8665,N_6491);
and U14760 (N_14760,N_7887,N_8734);
and U14761 (N_14761,N_7019,N_9705);
or U14762 (N_14762,N_8123,N_6456);
or U14763 (N_14763,N_5793,N_6834);
nand U14764 (N_14764,N_7575,N_8252);
and U14765 (N_14765,N_6866,N_5757);
nand U14766 (N_14766,N_8507,N_7576);
or U14767 (N_14767,N_8785,N_9681);
nand U14768 (N_14768,N_9309,N_8251);
or U14769 (N_14769,N_5811,N_6777);
nand U14770 (N_14770,N_9765,N_5548);
or U14771 (N_14771,N_8805,N_5671);
and U14772 (N_14772,N_5037,N_7507);
xnor U14773 (N_14773,N_7029,N_9065);
or U14774 (N_14774,N_7961,N_7787);
or U14775 (N_14775,N_8181,N_7703);
and U14776 (N_14776,N_6204,N_9078);
and U14777 (N_14777,N_7180,N_8212);
or U14778 (N_14778,N_5463,N_7270);
nor U14779 (N_14779,N_6770,N_8100);
and U14780 (N_14780,N_7572,N_5730);
or U14781 (N_14781,N_7916,N_9690);
or U14782 (N_14782,N_6884,N_5448);
or U14783 (N_14783,N_7906,N_9159);
nor U14784 (N_14784,N_6115,N_5099);
nor U14785 (N_14785,N_8071,N_7996);
xnor U14786 (N_14786,N_6696,N_7260);
and U14787 (N_14787,N_8603,N_6807);
or U14788 (N_14788,N_8826,N_5829);
nand U14789 (N_14789,N_7050,N_6803);
nand U14790 (N_14790,N_5340,N_9252);
nor U14791 (N_14791,N_9490,N_6151);
and U14792 (N_14792,N_9643,N_5171);
nand U14793 (N_14793,N_5932,N_5007);
nand U14794 (N_14794,N_8908,N_8647);
nor U14795 (N_14795,N_9778,N_9519);
nor U14796 (N_14796,N_6164,N_7473);
nor U14797 (N_14797,N_5347,N_5850);
nand U14798 (N_14798,N_9797,N_6855);
nand U14799 (N_14799,N_6794,N_6338);
or U14800 (N_14800,N_7928,N_6764);
nand U14801 (N_14801,N_5749,N_9144);
and U14802 (N_14802,N_7281,N_9358);
nand U14803 (N_14803,N_7480,N_6342);
nand U14804 (N_14804,N_7003,N_8096);
nand U14805 (N_14805,N_8302,N_6755);
or U14806 (N_14806,N_9664,N_9860);
or U14807 (N_14807,N_6206,N_8720);
nand U14808 (N_14808,N_9152,N_8620);
and U14809 (N_14809,N_5456,N_9235);
xor U14810 (N_14810,N_5456,N_7501);
or U14811 (N_14811,N_5154,N_5514);
and U14812 (N_14812,N_6212,N_6110);
nand U14813 (N_14813,N_8579,N_7216);
xnor U14814 (N_14814,N_5288,N_7849);
xor U14815 (N_14815,N_7162,N_9116);
nor U14816 (N_14816,N_7010,N_5513);
or U14817 (N_14817,N_5079,N_9719);
nand U14818 (N_14818,N_9451,N_6552);
and U14819 (N_14819,N_5321,N_9919);
nor U14820 (N_14820,N_9368,N_8251);
nor U14821 (N_14821,N_5151,N_6959);
and U14822 (N_14822,N_6568,N_5445);
and U14823 (N_14823,N_7523,N_5936);
nor U14824 (N_14824,N_8677,N_8627);
and U14825 (N_14825,N_9406,N_5240);
xor U14826 (N_14826,N_9377,N_8994);
and U14827 (N_14827,N_8644,N_5587);
nand U14828 (N_14828,N_6202,N_7755);
nand U14829 (N_14829,N_5604,N_7844);
xor U14830 (N_14830,N_8307,N_7541);
nor U14831 (N_14831,N_9042,N_6933);
nor U14832 (N_14832,N_5356,N_5982);
or U14833 (N_14833,N_6829,N_7106);
nor U14834 (N_14834,N_5208,N_8300);
nor U14835 (N_14835,N_7573,N_9782);
and U14836 (N_14836,N_8877,N_5063);
nand U14837 (N_14837,N_7555,N_7761);
or U14838 (N_14838,N_9707,N_6438);
nor U14839 (N_14839,N_8089,N_5200);
nand U14840 (N_14840,N_8922,N_9453);
and U14841 (N_14841,N_9409,N_5272);
and U14842 (N_14842,N_8821,N_5810);
and U14843 (N_14843,N_7260,N_5785);
or U14844 (N_14844,N_9554,N_5679);
or U14845 (N_14845,N_9483,N_9397);
nand U14846 (N_14846,N_6429,N_9878);
nand U14847 (N_14847,N_7902,N_9213);
nor U14848 (N_14848,N_7041,N_8941);
nand U14849 (N_14849,N_8818,N_9377);
nand U14850 (N_14850,N_7240,N_9762);
nor U14851 (N_14851,N_6274,N_6386);
and U14852 (N_14852,N_8443,N_8048);
or U14853 (N_14853,N_5886,N_5902);
and U14854 (N_14854,N_8287,N_9970);
xnor U14855 (N_14855,N_7613,N_5414);
nor U14856 (N_14856,N_9190,N_5847);
xor U14857 (N_14857,N_8019,N_7617);
or U14858 (N_14858,N_9298,N_9952);
and U14859 (N_14859,N_7152,N_6796);
nor U14860 (N_14860,N_8388,N_5191);
and U14861 (N_14861,N_8509,N_6000);
nor U14862 (N_14862,N_5878,N_9535);
nand U14863 (N_14863,N_9805,N_7301);
xnor U14864 (N_14864,N_7205,N_7951);
nand U14865 (N_14865,N_9304,N_9727);
xor U14866 (N_14866,N_7710,N_5447);
nand U14867 (N_14867,N_6990,N_5350);
nand U14868 (N_14868,N_6192,N_6954);
xnor U14869 (N_14869,N_6277,N_5564);
nor U14870 (N_14870,N_6822,N_5312);
xnor U14871 (N_14871,N_7164,N_9874);
or U14872 (N_14872,N_5968,N_8527);
and U14873 (N_14873,N_7415,N_5958);
or U14874 (N_14874,N_9474,N_6194);
xnor U14875 (N_14875,N_5707,N_7871);
nor U14876 (N_14876,N_9326,N_8125);
or U14877 (N_14877,N_7077,N_7044);
nand U14878 (N_14878,N_9096,N_7478);
nor U14879 (N_14879,N_5077,N_7909);
nand U14880 (N_14880,N_8352,N_7667);
nand U14881 (N_14881,N_5926,N_9586);
nor U14882 (N_14882,N_8121,N_7472);
nand U14883 (N_14883,N_8884,N_9034);
or U14884 (N_14884,N_9254,N_6729);
and U14885 (N_14885,N_9139,N_6993);
nand U14886 (N_14886,N_9812,N_8146);
or U14887 (N_14887,N_7162,N_5706);
xnor U14888 (N_14888,N_6081,N_8463);
or U14889 (N_14889,N_6846,N_6026);
and U14890 (N_14890,N_8350,N_8102);
nor U14891 (N_14891,N_8022,N_9140);
nand U14892 (N_14892,N_9725,N_5329);
or U14893 (N_14893,N_5729,N_9402);
nand U14894 (N_14894,N_6002,N_6316);
nor U14895 (N_14895,N_8340,N_7451);
or U14896 (N_14896,N_9527,N_5747);
nor U14897 (N_14897,N_8600,N_5246);
and U14898 (N_14898,N_7853,N_7493);
and U14899 (N_14899,N_5145,N_5887);
or U14900 (N_14900,N_7936,N_8970);
nor U14901 (N_14901,N_7733,N_6955);
or U14902 (N_14902,N_6620,N_6942);
nor U14903 (N_14903,N_9076,N_5499);
xor U14904 (N_14904,N_9675,N_9455);
or U14905 (N_14905,N_5987,N_6875);
and U14906 (N_14906,N_9631,N_6223);
and U14907 (N_14907,N_8172,N_6883);
and U14908 (N_14908,N_8431,N_8290);
nand U14909 (N_14909,N_9232,N_6871);
or U14910 (N_14910,N_6704,N_7594);
or U14911 (N_14911,N_7791,N_9265);
or U14912 (N_14912,N_8531,N_8030);
nor U14913 (N_14913,N_5275,N_9492);
or U14914 (N_14914,N_9141,N_7032);
and U14915 (N_14915,N_6221,N_7204);
xor U14916 (N_14916,N_9848,N_7996);
nor U14917 (N_14917,N_7967,N_8210);
and U14918 (N_14918,N_7172,N_8221);
and U14919 (N_14919,N_7434,N_7926);
nor U14920 (N_14920,N_7161,N_7575);
or U14921 (N_14921,N_8508,N_9331);
and U14922 (N_14922,N_9557,N_9703);
and U14923 (N_14923,N_6809,N_5296);
nand U14924 (N_14924,N_7150,N_9871);
xnor U14925 (N_14925,N_6795,N_7306);
nand U14926 (N_14926,N_7399,N_8983);
nand U14927 (N_14927,N_5185,N_5885);
or U14928 (N_14928,N_8405,N_5604);
nand U14929 (N_14929,N_6929,N_5131);
or U14930 (N_14930,N_9916,N_5008);
or U14931 (N_14931,N_8933,N_8475);
nand U14932 (N_14932,N_8024,N_6062);
xnor U14933 (N_14933,N_5048,N_8961);
xnor U14934 (N_14934,N_8550,N_7064);
nor U14935 (N_14935,N_7355,N_9810);
or U14936 (N_14936,N_7619,N_6014);
and U14937 (N_14937,N_7905,N_9928);
nand U14938 (N_14938,N_7458,N_7659);
or U14939 (N_14939,N_9502,N_6744);
xnor U14940 (N_14940,N_6516,N_6507);
nand U14941 (N_14941,N_7002,N_9898);
or U14942 (N_14942,N_8188,N_8177);
nor U14943 (N_14943,N_8696,N_8530);
nand U14944 (N_14944,N_8208,N_5170);
or U14945 (N_14945,N_5614,N_9061);
nand U14946 (N_14946,N_9728,N_6853);
xor U14947 (N_14947,N_8377,N_7305);
or U14948 (N_14948,N_8105,N_7184);
or U14949 (N_14949,N_6554,N_5260);
nor U14950 (N_14950,N_5806,N_6056);
xor U14951 (N_14951,N_9340,N_5228);
nor U14952 (N_14952,N_8451,N_7386);
nor U14953 (N_14953,N_9831,N_8812);
nand U14954 (N_14954,N_9036,N_9114);
nand U14955 (N_14955,N_8407,N_8324);
or U14956 (N_14956,N_7950,N_5256);
and U14957 (N_14957,N_9451,N_6522);
and U14958 (N_14958,N_7885,N_7799);
nand U14959 (N_14959,N_7725,N_5446);
and U14960 (N_14960,N_8699,N_9231);
nand U14961 (N_14961,N_5164,N_6824);
and U14962 (N_14962,N_7451,N_5146);
or U14963 (N_14963,N_9681,N_6382);
nor U14964 (N_14964,N_7352,N_6719);
nor U14965 (N_14965,N_8199,N_6876);
xnor U14966 (N_14966,N_9320,N_8494);
nor U14967 (N_14967,N_8443,N_8308);
xor U14968 (N_14968,N_5744,N_7778);
nor U14969 (N_14969,N_9726,N_7281);
nand U14970 (N_14970,N_8048,N_9428);
or U14971 (N_14971,N_8010,N_6357);
nor U14972 (N_14972,N_7158,N_7442);
xor U14973 (N_14973,N_6262,N_8931);
or U14974 (N_14974,N_5655,N_8938);
nor U14975 (N_14975,N_6574,N_6371);
or U14976 (N_14976,N_7558,N_5883);
nand U14977 (N_14977,N_5539,N_9119);
and U14978 (N_14978,N_7299,N_9577);
or U14979 (N_14979,N_9127,N_9689);
or U14980 (N_14980,N_8206,N_9750);
nand U14981 (N_14981,N_9323,N_8918);
nor U14982 (N_14982,N_6695,N_6924);
nor U14983 (N_14983,N_9830,N_5223);
and U14984 (N_14984,N_6932,N_6791);
or U14985 (N_14985,N_5592,N_7401);
xor U14986 (N_14986,N_8522,N_6496);
xnor U14987 (N_14987,N_9349,N_7976);
nand U14988 (N_14988,N_9562,N_8487);
and U14989 (N_14989,N_9763,N_7878);
nor U14990 (N_14990,N_9605,N_6880);
and U14991 (N_14991,N_9108,N_9365);
or U14992 (N_14992,N_8676,N_8075);
nand U14993 (N_14993,N_9936,N_8859);
and U14994 (N_14994,N_6611,N_8913);
xor U14995 (N_14995,N_8825,N_5637);
nor U14996 (N_14996,N_6573,N_6863);
and U14997 (N_14997,N_8183,N_8971);
and U14998 (N_14998,N_7458,N_9557);
xnor U14999 (N_14999,N_7304,N_5922);
or U15000 (N_15000,N_14598,N_13154);
nand U15001 (N_15001,N_13566,N_14576);
or U15002 (N_15002,N_13415,N_12187);
nor U15003 (N_15003,N_13427,N_14532);
nor U15004 (N_15004,N_11629,N_13753);
and U15005 (N_15005,N_13056,N_14872);
nor U15006 (N_15006,N_14294,N_10399);
or U15007 (N_15007,N_11514,N_14408);
nor U15008 (N_15008,N_11607,N_13145);
xor U15009 (N_15009,N_10348,N_10760);
nor U15010 (N_15010,N_13240,N_11770);
nand U15011 (N_15011,N_13182,N_12370);
and U15012 (N_15012,N_10004,N_14934);
or U15013 (N_15013,N_14647,N_14825);
nor U15014 (N_15014,N_12545,N_10613);
or U15015 (N_15015,N_12269,N_13435);
and U15016 (N_15016,N_14811,N_14416);
xnor U15017 (N_15017,N_11823,N_12121);
nor U15018 (N_15018,N_11047,N_12407);
nand U15019 (N_15019,N_13982,N_14435);
and U15020 (N_15020,N_11013,N_11413);
nand U15021 (N_15021,N_11791,N_12787);
nor U15022 (N_15022,N_12989,N_10293);
and U15023 (N_15023,N_12045,N_14241);
and U15024 (N_15024,N_10472,N_12313);
xor U15025 (N_15025,N_14649,N_11621);
nand U15026 (N_15026,N_14267,N_11160);
nor U15027 (N_15027,N_10061,N_12247);
or U15028 (N_15028,N_13530,N_14918);
nand U15029 (N_15029,N_10618,N_13223);
nand U15030 (N_15030,N_11051,N_13459);
xnor U15031 (N_15031,N_12780,N_14575);
or U15032 (N_15032,N_14310,N_13541);
nor U15033 (N_15033,N_12261,N_13087);
and U15034 (N_15034,N_11281,N_10540);
and U15035 (N_15035,N_10351,N_10683);
or U15036 (N_15036,N_14105,N_11066);
and U15037 (N_15037,N_13014,N_13705);
nand U15038 (N_15038,N_10296,N_11605);
and U15039 (N_15039,N_13698,N_11023);
nand U15040 (N_15040,N_10135,N_12974);
nand U15041 (N_15041,N_11722,N_11469);
or U15042 (N_15042,N_10038,N_14172);
or U15043 (N_15043,N_13318,N_12636);
xnor U15044 (N_15044,N_13481,N_10762);
nor U15045 (N_15045,N_12795,N_10813);
nor U15046 (N_15046,N_13767,N_11911);
nand U15047 (N_15047,N_13516,N_14523);
or U15048 (N_15048,N_14827,N_10938);
nor U15049 (N_15049,N_12430,N_12620);
nor U15050 (N_15050,N_14099,N_11069);
and U15051 (N_15051,N_13099,N_12087);
nand U15052 (N_15052,N_13444,N_10854);
nand U15053 (N_15053,N_11463,N_11252);
or U15054 (N_15054,N_11902,N_14029);
nor U15055 (N_15055,N_14577,N_14604);
nand U15056 (N_15056,N_12466,N_14380);
and U15057 (N_15057,N_10736,N_14363);
and U15058 (N_15058,N_14221,N_11601);
nor U15059 (N_15059,N_10263,N_13887);
and U15060 (N_15060,N_14291,N_10478);
nand U15061 (N_15061,N_11624,N_13022);
or U15062 (N_15062,N_11080,N_11753);
or U15063 (N_15063,N_13817,N_10984);
nor U15064 (N_15064,N_14656,N_11206);
and U15065 (N_15065,N_11454,N_12808);
nor U15066 (N_15066,N_14373,N_10109);
xor U15067 (N_15067,N_11239,N_11232);
nand U15068 (N_15068,N_14789,N_14238);
or U15069 (N_15069,N_12576,N_13072);
or U15070 (N_15070,N_11082,N_10810);
nor U15071 (N_15071,N_12608,N_14591);
or U15072 (N_15072,N_13218,N_10918);
nand U15073 (N_15073,N_14754,N_10531);
nand U15074 (N_15074,N_11555,N_12901);
nor U15075 (N_15075,N_14637,N_10616);
and U15076 (N_15076,N_13302,N_11338);
or U15077 (N_15077,N_10852,N_12020);
or U15078 (N_15078,N_14376,N_12625);
and U15079 (N_15079,N_12423,N_13197);
and U15080 (N_15080,N_12053,N_10922);
nand U15081 (N_15081,N_13569,N_10331);
or U15082 (N_15082,N_13059,N_13143);
xor U15083 (N_15083,N_12554,N_10889);
and U15084 (N_15084,N_13659,N_12497);
nand U15085 (N_15085,N_12951,N_13667);
xnor U15086 (N_15086,N_11456,N_11848);
nor U15087 (N_15087,N_12299,N_13579);
nor U15088 (N_15088,N_10771,N_13251);
nand U15089 (N_15089,N_11966,N_13019);
or U15090 (N_15090,N_14243,N_13121);
nor U15091 (N_15091,N_12415,N_14348);
and U15092 (N_15092,N_10416,N_10907);
nand U15093 (N_15093,N_14962,N_14981);
and U15094 (N_15094,N_14201,N_12238);
or U15095 (N_15095,N_12578,N_13872);
or U15096 (N_15096,N_12022,N_14834);
nand U15097 (N_15097,N_10214,N_10601);
nand U15098 (N_15098,N_12420,N_10875);
nand U15099 (N_15099,N_14928,N_10180);
and U15100 (N_15100,N_13965,N_10971);
or U15101 (N_15101,N_13419,N_11937);
nor U15102 (N_15102,N_11596,N_12995);
and U15103 (N_15103,N_11512,N_10735);
xor U15104 (N_15104,N_12535,N_10697);
xor U15105 (N_15105,N_13720,N_12230);
or U15106 (N_15106,N_14704,N_14430);
or U15107 (N_15107,N_13763,N_10352);
and U15108 (N_15108,N_11914,N_10315);
or U15109 (N_15109,N_12517,N_14228);
or U15110 (N_15110,N_12820,N_14236);
and U15111 (N_15111,N_14566,N_12809);
and U15112 (N_15112,N_12613,N_11659);
nand U15113 (N_15113,N_12573,N_10928);
and U15114 (N_15114,N_10402,N_10693);
and U15115 (N_15115,N_10093,N_13142);
nand U15116 (N_15116,N_11059,N_12461);
nor U15117 (N_15117,N_14075,N_10503);
or U15118 (N_15118,N_14164,N_14752);
nor U15119 (N_15119,N_13139,N_10120);
or U15120 (N_15120,N_13396,N_12871);
nor U15121 (N_15121,N_14061,N_14046);
nor U15122 (N_15122,N_12255,N_12579);
or U15123 (N_15123,N_12450,N_14003);
nand U15124 (N_15124,N_13583,N_13126);
or U15125 (N_15125,N_14020,N_13421);
and U15126 (N_15126,N_14545,N_10749);
and U15127 (N_15127,N_14657,N_11813);
nand U15128 (N_15128,N_14472,N_13880);
nand U15129 (N_15129,N_13050,N_10040);
nor U15130 (N_15130,N_12043,N_13008);
nor U15131 (N_15131,N_14091,N_14452);
nor U15132 (N_15132,N_14331,N_12274);
nand U15133 (N_15133,N_14793,N_12742);
or U15134 (N_15134,N_10567,N_10539);
and U15135 (N_15135,N_12357,N_11092);
nand U15136 (N_15136,N_14546,N_12186);
nor U15137 (N_15137,N_11064,N_13348);
or U15138 (N_15138,N_10519,N_13450);
nand U15139 (N_15139,N_13621,N_13160);
and U15140 (N_15140,N_13372,N_12102);
nor U15141 (N_15141,N_10378,N_11274);
xnor U15142 (N_15142,N_11570,N_10667);
and U15143 (N_15143,N_14551,N_14964);
xnor U15144 (N_15144,N_10328,N_10238);
nand U15145 (N_15145,N_12325,N_14326);
and U15146 (N_15146,N_14305,N_14448);
nand U15147 (N_15147,N_13106,N_13242);
nor U15148 (N_15148,N_11270,N_10851);
xor U15149 (N_15149,N_13342,N_13109);
and U15150 (N_15150,N_10610,N_12124);
or U15151 (N_15151,N_13407,N_10264);
and U15152 (N_15152,N_10013,N_10888);
or U15153 (N_15153,N_12271,N_11974);
nor U15154 (N_15154,N_11331,N_13624);
and U15155 (N_15155,N_13849,N_10273);
and U15156 (N_15156,N_13007,N_14512);
or U15157 (N_15157,N_12418,N_10964);
nor U15158 (N_15158,N_14322,N_14403);
or U15159 (N_15159,N_11612,N_13042);
or U15160 (N_15160,N_14325,N_12318);
nand U15161 (N_15161,N_13046,N_14854);
and U15162 (N_15162,N_10972,N_11461);
nor U15163 (N_15163,N_10747,N_10921);
and U15164 (N_15164,N_11280,N_10623);
and U15165 (N_15165,N_10757,N_13426);
nor U15166 (N_15166,N_10552,N_13997);
xnor U15167 (N_15167,N_14304,N_10802);
or U15168 (N_15168,N_11345,N_12036);
and U15169 (N_15169,N_13264,N_12574);
xnor U15170 (N_15170,N_14968,N_10104);
nand U15171 (N_15171,N_10193,N_11482);
nor U15172 (N_15172,N_11958,N_10565);
nand U15173 (N_15173,N_13319,N_11585);
and U15174 (N_15174,N_13171,N_10787);
nor U15175 (N_15175,N_14599,N_11645);
nand U15176 (N_15176,N_13577,N_11674);
nor U15177 (N_15177,N_12954,N_10189);
nor U15178 (N_15178,N_14278,N_12847);
nand U15179 (N_15179,N_12559,N_14174);
or U15180 (N_15180,N_10224,N_11265);
nand U15181 (N_15181,N_12289,N_10817);
and U15182 (N_15182,N_11116,N_10829);
nor U15183 (N_15183,N_10827,N_14952);
and U15184 (N_15184,N_10611,N_13995);
nor U15185 (N_15185,N_14824,N_10671);
and U15186 (N_15186,N_12499,N_13905);
xnor U15187 (N_15187,N_12642,N_12646);
nand U15188 (N_15188,N_12540,N_14786);
nand U15189 (N_15189,N_12500,N_10421);
or U15190 (N_15190,N_12745,N_11863);
xnor U15191 (N_15191,N_11943,N_11316);
nand U15192 (N_15192,N_13322,N_12414);
nor U15193 (N_15193,N_14026,N_13876);
nor U15194 (N_15194,N_10592,N_13495);
nor U15195 (N_15195,N_13216,N_12394);
nand U15196 (N_15196,N_11936,N_11362);
nor U15197 (N_15197,N_12052,N_10807);
nand U15198 (N_15198,N_14372,N_13846);
nand U15199 (N_15199,N_13703,N_14763);
nor U15200 (N_15200,N_11704,N_14117);
nor U15201 (N_15201,N_12235,N_14313);
or U15202 (N_15202,N_13693,N_14818);
and U15203 (N_15203,N_13815,N_14541);
and U15204 (N_15204,N_12383,N_11844);
xor U15205 (N_15205,N_11416,N_13899);
nor U15206 (N_15206,N_10513,N_13339);
or U15207 (N_15207,N_10857,N_11654);
and U15208 (N_15208,N_13490,N_12301);
and U15209 (N_15209,N_10115,N_14944);
nor U15210 (N_15210,N_14664,N_10275);
or U15211 (N_15211,N_11490,N_11054);
nand U15212 (N_15212,N_13534,N_12718);
or U15213 (N_15213,N_11616,N_11201);
and U15214 (N_15214,N_11420,N_11320);
nand U15215 (N_15215,N_14254,N_11744);
and U15216 (N_15216,N_12722,N_11003);
nand U15217 (N_15217,N_13984,N_12976);
nand U15218 (N_15218,N_12577,N_13232);
nand U15219 (N_15219,N_14764,N_12580);
and U15220 (N_15220,N_11878,N_12980);
nand U15221 (N_15221,N_11314,N_14893);
or U15222 (N_15222,N_12009,N_11646);
and U15223 (N_15223,N_13290,N_11904);
or U15224 (N_15224,N_13727,N_12338);
nor U15225 (N_15225,N_14625,N_12899);
or U15226 (N_15226,N_13128,N_13431);
or U15227 (N_15227,N_11325,N_10725);
or U15228 (N_15228,N_12404,N_12647);
nand U15229 (N_15229,N_12427,N_14734);
or U15230 (N_15230,N_13871,N_12199);
nor U15231 (N_15231,N_10590,N_13535);
xor U15232 (N_15232,N_10433,N_10242);
nor U15233 (N_15233,N_14891,N_13889);
and U15234 (N_15234,N_13119,N_13906);
nand U15235 (N_15235,N_14629,N_14317);
nand U15236 (N_15236,N_13980,N_13606);
and U15237 (N_15237,N_12965,N_10199);
nand U15238 (N_15238,N_14205,N_14343);
nor U15239 (N_15239,N_10170,N_13432);
nor U15240 (N_15240,N_10371,N_11954);
or U15241 (N_15241,N_10772,N_12277);
xor U15242 (N_15242,N_10222,N_11130);
nor U15243 (N_15243,N_12323,N_13797);
and U15244 (N_15244,N_10420,N_10368);
nor U15245 (N_15245,N_13992,N_12228);
or U15246 (N_15246,N_14052,N_10290);
nand U15247 (N_15247,N_14642,N_14908);
and U15248 (N_15248,N_13902,N_11705);
and U15249 (N_15249,N_13069,N_14162);
nor U15250 (N_15250,N_12754,N_10377);
xnor U15251 (N_15251,N_14300,N_10660);
xor U15252 (N_15252,N_10720,N_12772);
xnor U15253 (N_15253,N_14142,N_12986);
nor U15254 (N_15254,N_12963,N_13248);
xnor U15255 (N_15255,N_11896,N_14220);
nor U15256 (N_15256,N_13466,N_12463);
and U15257 (N_15257,N_12555,N_14086);
nor U15258 (N_15258,N_13863,N_14947);
or U15259 (N_15259,N_11979,N_14777);
and U15260 (N_15260,N_10094,N_13532);
and U15261 (N_15261,N_14415,N_12770);
nor U15262 (N_15262,N_12978,N_11366);
xnor U15263 (N_15263,N_14101,N_13035);
nand U15264 (N_15264,N_12674,N_14769);
xnor U15265 (N_15265,N_14796,N_13161);
and U15266 (N_15266,N_12640,N_11226);
or U15267 (N_15267,N_10396,N_11683);
and U15268 (N_15268,N_12098,N_10309);
nor U15269 (N_15269,N_11496,N_13528);
or U15270 (N_15270,N_13546,N_13036);
nor U15271 (N_15271,N_14048,N_13335);
or U15272 (N_15272,N_14986,N_11711);
or U15273 (N_15273,N_10544,N_11984);
nor U15274 (N_15274,N_13941,N_12833);
nand U15275 (N_15275,N_10583,N_10225);
and U15276 (N_15276,N_14862,N_14203);
nand U15277 (N_15277,N_11712,N_12694);
and U15278 (N_15278,N_12119,N_12519);
xor U15279 (N_15279,N_10249,N_12107);
nor U15280 (N_15280,N_13857,N_10450);
nand U15281 (N_15281,N_13102,N_13328);
nand U15282 (N_15282,N_11488,N_13475);
nor U15283 (N_15283,N_13295,N_11223);
nor U15284 (N_15284,N_14804,N_12032);
and U15285 (N_15285,N_12455,N_10607);
nor U15286 (N_15286,N_11898,N_14723);
or U15287 (N_15287,N_14992,N_14732);
and U15288 (N_15288,N_14128,N_12624);
nor U15289 (N_15289,N_14840,N_11495);
nor U15290 (N_15290,N_10471,N_14065);
and U15291 (N_15291,N_12035,N_11908);
or U15292 (N_15292,N_11737,N_12944);
nor U15293 (N_15293,N_14386,N_14590);
or U15294 (N_15294,N_11244,N_14096);
xnor U15295 (N_15295,N_12641,N_11525);
or U15296 (N_15296,N_11784,N_13162);
xnor U15297 (N_15297,N_11963,N_10107);
or U15298 (N_15298,N_14250,N_14171);
nor U15299 (N_15299,N_14716,N_14062);
and U15300 (N_15300,N_12309,N_10241);
xnor U15301 (N_15301,N_14730,N_14593);
nor U15302 (N_15302,N_12633,N_13356);
nor U15303 (N_15303,N_14829,N_12200);
and U15304 (N_15304,N_11897,N_11732);
xnor U15305 (N_15305,N_13023,N_11716);
and U15306 (N_15306,N_11661,N_14700);
or U15307 (N_15307,N_14258,N_14850);
and U15308 (N_15308,N_13101,N_10205);
nor U15309 (N_15309,N_11222,N_13428);
or U15310 (N_15310,N_11090,N_13167);
nor U15311 (N_15311,N_11589,N_11321);
nor U15312 (N_15312,N_13491,N_12308);
nand U15313 (N_15313,N_12769,N_10404);
nor U15314 (N_15314,N_12533,N_13608);
nand U15315 (N_15315,N_12223,N_11934);
nand U15316 (N_15316,N_12538,N_13951);
and U15317 (N_15317,N_14078,N_13647);
nand U15318 (N_15318,N_10323,N_12807);
nand U15319 (N_15319,N_12214,N_11335);
xnor U15320 (N_15320,N_11472,N_13325);
and U15321 (N_15321,N_14869,N_14297);
nand U15322 (N_15322,N_11796,N_12355);
nor U15323 (N_15323,N_11558,N_13550);
nand U15324 (N_15324,N_10215,N_13658);
xor U15325 (N_15325,N_12347,N_14342);
xnor U15326 (N_15326,N_10380,N_11079);
and U15327 (N_15327,N_10367,N_13685);
and U15328 (N_15328,N_10538,N_10021);
and U15329 (N_15329,N_10555,N_10451);
and U15330 (N_15330,N_13637,N_10291);
xnor U15331 (N_15331,N_10071,N_12703);
and U15332 (N_15332,N_12331,N_12557);
xor U15333 (N_15333,N_12652,N_12391);
and U15334 (N_15334,N_13144,N_12680);
and U15335 (N_15335,N_10561,N_11219);
nor U15336 (N_15336,N_11052,N_14059);
and U15337 (N_15337,N_11916,N_14442);
nor U15338 (N_15338,N_10432,N_13988);
or U15339 (N_15339,N_11688,N_13417);
nand U15340 (N_15340,N_11011,N_10288);
nor U15341 (N_15341,N_11238,N_14196);
or U15342 (N_15342,N_10882,N_14368);
and U15343 (N_15343,N_12921,N_11697);
or U15344 (N_15344,N_14803,N_13524);
nor U15345 (N_15345,N_11019,N_13645);
or U15346 (N_15346,N_14311,N_12791);
nor U15347 (N_15347,N_10550,N_11967);
nor U15348 (N_15348,N_13808,N_14856);
nand U15349 (N_15349,N_14023,N_14182);
nor U15350 (N_15350,N_12846,N_11377);
or U15351 (N_15351,N_14034,N_11418);
or U15352 (N_15352,N_14272,N_12182);
nand U15353 (N_15353,N_12526,N_10808);
nand U15354 (N_15354,N_14815,N_13153);
or U15355 (N_15355,N_14580,N_13411);
nor U15356 (N_15356,N_12425,N_12167);
or U15357 (N_15357,N_14633,N_11992);
and U15358 (N_15358,N_14244,N_13085);
nand U15359 (N_15359,N_10691,N_10409);
nor U15360 (N_15360,N_13410,N_14123);
or U15361 (N_15361,N_10248,N_11421);
or U15362 (N_15362,N_14838,N_10437);
or U15363 (N_15363,N_13304,N_10558);
or U15364 (N_15364,N_12419,N_13299);
and U15365 (N_15365,N_11409,N_13355);
and U15366 (N_15366,N_10981,N_14788);
nand U15367 (N_15367,N_11040,N_12948);
nand U15368 (N_15368,N_10463,N_12815);
xnor U15369 (N_15369,N_12992,N_11257);
nand U15370 (N_15370,N_11315,N_14044);
and U15371 (N_15371,N_12145,N_14939);
and U15372 (N_15372,N_11759,N_12918);
nand U15373 (N_15373,N_13627,N_14334);
and U15374 (N_15374,N_13639,N_11837);
or U15375 (N_15375,N_11946,N_13843);
or U15376 (N_15376,N_11277,N_14858);
xor U15377 (N_15377,N_10418,N_12074);
or U15378 (N_15378,N_11286,N_10111);
or U15379 (N_15379,N_13329,N_12738);
nand U15380 (N_15380,N_13231,N_12249);
nor U15381 (N_15381,N_14747,N_11288);
or U15382 (N_15382,N_10486,N_14043);
xnor U15383 (N_15383,N_10721,N_10443);
or U15384 (N_15384,N_12628,N_10985);
or U15385 (N_15385,N_11459,N_12066);
and U15386 (N_15386,N_12439,N_14961);
xnor U15387 (N_15387,N_10308,N_10920);
nor U15388 (N_15388,N_14279,N_13386);
or U15389 (N_15389,N_13560,N_14722);
and U15390 (N_15390,N_14190,N_12507);
and U15391 (N_15391,N_12821,N_11522);
or U15392 (N_15392,N_13625,N_13125);
and U15393 (N_15393,N_10904,N_13931);
nand U15394 (N_15394,N_10496,N_13116);
nor U15395 (N_15395,N_11284,N_14214);
nand U15396 (N_15396,N_12159,N_12155);
or U15397 (N_15397,N_12909,N_11031);
or U15398 (N_15398,N_11969,N_11489);
nand U15399 (N_15399,N_12089,N_11307);
nand U15400 (N_15400,N_13467,N_12822);
nor U15401 (N_15401,N_11207,N_12049);
nor U15402 (N_15402,N_13100,N_14892);
and U15403 (N_15403,N_14366,N_13391);
or U15404 (N_15404,N_14296,N_10456);
nand U15405 (N_15405,N_10259,N_12568);
nand U15406 (N_15406,N_11457,N_13986);
and U15407 (N_15407,N_11107,N_12710);
nor U15408 (N_15408,N_12851,N_12057);
nand U15409 (N_15409,N_10332,N_10726);
nor U15410 (N_15410,N_14424,N_14739);
xor U15411 (N_15411,N_12164,N_10588);
and U15412 (N_15412,N_10303,N_12867);
xor U15413 (N_15413,N_14674,N_11725);
or U15414 (N_15414,N_11910,N_10289);
nand U15415 (N_15415,N_14570,N_10568);
nor U15416 (N_15416,N_11012,N_11115);
nand U15417 (N_15417,N_12442,N_14271);
or U15418 (N_15418,N_14725,N_14581);
or U15419 (N_15419,N_11310,N_12071);
or U15420 (N_15420,N_13373,N_12334);
and U15421 (N_15421,N_14170,N_10000);
and U15422 (N_15422,N_10641,N_12597);
and U15423 (N_15423,N_10564,N_13312);
nor U15424 (N_15424,N_12964,N_13499);
nand U15425 (N_15425,N_10390,N_11780);
nand U15426 (N_15426,N_12571,N_10006);
nor U15427 (N_15427,N_14379,N_14400);
or U15428 (N_15428,N_14684,N_12421);
or U15429 (N_15429,N_11691,N_11939);
nand U15430 (N_15430,N_14618,N_13034);
nand U15431 (N_15431,N_10255,N_10270);
and U15432 (N_15432,N_10043,N_12881);
nand U15433 (N_15433,N_10980,N_11842);
nand U15434 (N_15434,N_11535,N_11774);
nand U15435 (N_15435,N_10614,N_14165);
nand U15436 (N_15436,N_11041,N_12708);
nor U15437 (N_15437,N_11886,N_14724);
or U15438 (N_15438,N_13193,N_11533);
and U15439 (N_15439,N_11743,N_10152);
or U15440 (N_15440,N_12008,N_13283);
or U15441 (N_15441,N_14149,N_12493);
nand U15442 (N_15442,N_14897,N_10258);
nand U15443 (N_15443,N_10990,N_10133);
nand U15444 (N_15444,N_14371,N_14421);
or U15445 (N_15445,N_14257,N_13096);
and U15446 (N_15446,N_14554,N_14066);
or U15447 (N_15447,N_11145,N_14444);
or U15448 (N_15448,N_11700,N_14436);
and U15449 (N_15449,N_13226,N_12161);
nor U15450 (N_15450,N_10350,N_10156);
or U15451 (N_15451,N_12868,N_13227);
and U15452 (N_15452,N_14175,N_14330);
nor U15453 (N_15453,N_10364,N_13664);
nand U15454 (N_15454,N_14359,N_11768);
or U15455 (N_15455,N_10487,N_13548);
or U15456 (N_15456,N_12514,N_14974);
nor U15457 (N_15457,N_10202,N_10317);
or U15458 (N_15458,N_14073,N_13826);
nor U15459 (N_15459,N_14639,N_10479);
and U15460 (N_15460,N_13307,N_10412);
nand U15461 (N_15461,N_11049,N_13555);
and U15462 (N_15462,N_10385,N_10843);
nand U15463 (N_15463,N_10183,N_10912);
and U15464 (N_15464,N_11398,N_12885);
or U15465 (N_15465,N_13385,N_14832);
nor U15466 (N_15466,N_14127,N_13853);
nand U15467 (N_15467,N_11800,N_12835);
nand U15468 (N_15468,N_12490,N_14636);
or U15469 (N_15469,N_11304,N_11322);
and U15470 (N_15470,N_11074,N_10692);
and U15471 (N_15471,N_10655,N_14828);
and U15472 (N_15472,N_10481,N_10455);
nor U15473 (N_15473,N_10041,N_11499);
nand U15474 (N_15474,N_13107,N_13520);
nand U15475 (N_15475,N_12586,N_10698);
nor U15476 (N_15476,N_14107,N_10831);
nand U15477 (N_15477,N_13200,N_11430);
and U15478 (N_15478,N_14841,N_14874);
nand U15479 (N_15479,N_14204,N_13253);
and U15480 (N_15480,N_10830,N_14081);
or U15481 (N_15481,N_11828,N_14536);
nor U15482 (N_15482,N_14660,N_12563);
and U15483 (N_15483,N_13246,N_11524);
and U15484 (N_15484,N_11617,N_12521);
and U15485 (N_15485,N_11113,N_14845);
and U15486 (N_15486,N_11255,N_13090);
xor U15487 (N_15487,N_11452,N_11870);
or U15488 (N_15488,N_14530,N_11932);
nand U15489 (N_15489,N_11851,N_11433);
nand U15490 (N_15490,N_11808,N_14457);
and U15491 (N_15491,N_13949,N_13781);
and U15492 (N_15492,N_14715,N_12184);
nor U15493 (N_15493,N_14277,N_10163);
nand U15494 (N_15494,N_14925,N_11258);
nor U15495 (N_15495,N_11050,N_12111);
nand U15496 (N_15496,N_11819,N_10457);
xnor U15497 (N_15497,N_10936,N_13701);
or U15498 (N_15498,N_13821,N_14574);
and U15499 (N_15499,N_10379,N_13613);
nor U15500 (N_15500,N_13237,N_10983);
nor U15501 (N_15501,N_13665,N_13829);
and U15502 (N_15502,N_14863,N_10805);
or U15503 (N_15503,N_14115,N_11531);
and U15504 (N_15504,N_13836,N_10870);
nand U15505 (N_15505,N_14596,N_14375);
or U15506 (N_15506,N_14222,N_14899);
nand U15507 (N_15507,N_14669,N_12943);
xnor U15508 (N_15508,N_12038,N_10458);
and U15509 (N_15509,N_11152,N_13732);
nand U15510 (N_15510,N_12542,N_10203);
and U15511 (N_15511,N_12583,N_14388);
or U15512 (N_15512,N_12934,N_13867);
nand U15513 (N_15513,N_10247,N_13183);
nand U15514 (N_15514,N_14791,N_13883);
nand U15515 (N_15515,N_14767,N_13651);
and U15516 (N_15516,N_13215,N_12166);
nand U15517 (N_15517,N_12859,N_11169);
nor U15518 (N_15518,N_12737,N_11384);
nand U15519 (N_15519,N_14844,N_13558);
or U15520 (N_15520,N_12375,N_13083);
and U15521 (N_15521,N_12106,N_14447);
or U15522 (N_15522,N_11833,N_14640);
nor U15523 (N_15523,N_11260,N_11141);
xor U15524 (N_15524,N_10220,N_11503);
or U15525 (N_15525,N_10557,N_10063);
and U15526 (N_15526,N_13212,N_11336);
nor U15527 (N_15527,N_14058,N_12409);
nor U15528 (N_15528,N_13765,N_13999);
nand U15529 (N_15529,N_13314,N_14833);
or U15530 (N_15530,N_11541,N_13810);
or U15531 (N_15531,N_12013,N_14905);
and U15532 (N_15532,N_13881,N_11408);
or U15533 (N_15533,N_13626,N_13205);
or U15534 (N_15534,N_12330,N_11824);
or U15535 (N_15535,N_12093,N_13075);
nor U15536 (N_15536,N_11872,N_10929);
and U15537 (N_15537,N_12887,N_10838);
and U15538 (N_15538,N_13172,N_14439);
nand U15539 (N_15539,N_11730,N_13848);
xnor U15540 (N_15540,N_10105,N_13683);
nor U15541 (N_15541,N_14682,N_10039);
and U15542 (N_15542,N_13222,N_11276);
or U15543 (N_15543,N_13729,N_12385);
or U15544 (N_15544,N_10598,N_14987);
or U15545 (N_15545,N_11960,N_11578);
or U15546 (N_15546,N_10609,N_11648);
xnor U15547 (N_15547,N_10911,N_13204);
or U15548 (N_15548,N_13184,N_13500);
nor U15549 (N_15549,N_12103,N_13320);
nor U15550 (N_15550,N_13054,N_12589);
and U15551 (N_15551,N_10201,N_12569);
nand U15552 (N_15552,N_14216,N_11002);
nand U15553 (N_15553,N_12544,N_11637);
nor U15554 (N_15554,N_12458,N_10410);
or U15555 (N_15555,N_11020,N_13855);
or U15556 (N_15556,N_13958,N_11926);
xor U15557 (N_15557,N_13582,N_11104);
nor U15558 (N_15558,N_11727,N_13492);
nand U15559 (N_15559,N_13671,N_12252);
or U15560 (N_15560,N_10318,N_12411);
nand U15561 (N_15561,N_12687,N_10355);
and U15562 (N_15562,N_11644,N_11234);
nand U15563 (N_15563,N_14487,N_10821);
xnor U15564 (N_15564,N_12340,N_11640);
nand U15565 (N_15565,N_11752,N_14045);
and U15566 (N_15566,N_10153,N_13779);
nor U15567 (N_15567,N_12185,N_14644);
and U15568 (N_15568,N_14514,N_10666);
or U15569 (N_15569,N_10718,N_11538);
nor U15570 (N_15570,N_14434,N_13839);
nand U15571 (N_15571,N_11361,N_10635);
nand U15572 (N_15572,N_12373,N_14180);
and U15573 (N_15573,N_13833,N_14412);
or U15574 (N_15574,N_10257,N_14332);
nor U15575 (N_15575,N_11584,N_11740);
nor U15576 (N_15576,N_13470,N_13148);
or U15577 (N_15577,N_11950,N_14426);
or U15578 (N_15578,N_14270,N_14904);
nor U15579 (N_15579,N_10297,N_13878);
and U15580 (N_15580,N_10855,N_12688);
and U15581 (N_15581,N_14999,N_10982);
or U15582 (N_15582,N_13504,N_11396);
or U15583 (N_15583,N_14208,N_13201);
and U15584 (N_15584,N_11952,N_13137);
and U15585 (N_15585,N_11738,N_10621);
or U15586 (N_15586,N_14607,N_14197);
nand U15587 (N_15587,N_12192,N_13830);
xnor U15588 (N_15588,N_14624,N_14836);
nand U15589 (N_15589,N_11532,N_10512);
nor U15590 (N_15590,N_11838,N_10335);
nand U15591 (N_15591,N_13165,N_10100);
and U15592 (N_15592,N_14153,N_11526);
nand U15593 (N_15593,N_13480,N_10322);
xor U15594 (N_15594,N_13398,N_10642);
and U15595 (N_15595,N_11745,N_14861);
nand U15596 (N_15596,N_12587,N_13323);
nand U15597 (N_15597,N_10998,N_13985);
xor U15598 (N_15598,N_12505,N_13864);
nand U15599 (N_15599,N_13272,N_10434);
nor U15600 (N_15600,N_12716,N_10663);
and U15601 (N_15601,N_11509,N_10498);
nand U15602 (N_15602,N_13488,N_12863);
nor U15603 (N_15603,N_11576,N_13818);
and U15604 (N_15604,N_10708,N_10979);
and U15605 (N_15605,N_12367,N_13131);
xor U15606 (N_15606,N_14612,N_12548);
nor U15607 (N_15607,N_14184,N_14347);
or U15608 (N_15608,N_12403,N_14678);
nand U15609 (N_15609,N_14568,N_12151);
and U15610 (N_15610,N_10036,N_12734);
or U15611 (N_15611,N_11028,N_10865);
or U15612 (N_15612,N_11504,N_11015);
or U15613 (N_15613,N_11455,N_11655);
nand U15614 (N_15614,N_10957,N_11138);
and U15615 (N_15615,N_11410,N_12004);
nor U15616 (N_15616,N_14980,N_10902);
and U15617 (N_15617,N_12024,N_11678);
nand U15618 (N_15618,N_12031,N_13702);
or U15619 (N_15619,N_14028,N_12824);
nand U15620 (N_15620,N_14499,N_13694);
xnor U15621 (N_15621,N_12695,N_11694);
nand U15622 (N_15622,N_10284,N_12643);
and U15623 (N_15623,N_12621,N_11442);
and U15624 (N_15624,N_10685,N_13037);
nor U15625 (N_15625,N_12552,N_10413);
nor U15626 (N_15626,N_13894,N_14748);
nand U15627 (N_15627,N_10700,N_10764);
nand U15628 (N_15628,N_10411,N_10744);
nand U15629 (N_15629,N_14776,N_13633);
and U15630 (N_15630,N_12696,N_10669);
nor U15631 (N_15631,N_11042,N_14606);
and U15632 (N_15632,N_11798,N_10160);
or U15633 (N_15633,N_12831,N_12528);
nor U15634 (N_15634,N_14775,N_11208);
and U15635 (N_15635,N_13601,N_14641);
and U15636 (N_15636,N_11048,N_12495);
nor U15637 (N_15637,N_11350,N_10643);
nand U15638 (N_15638,N_12698,N_13819);
nor U15639 (N_15639,N_14476,N_10231);
nor U15640 (N_15640,N_13374,N_11468);
or U15641 (N_15641,N_11633,N_12139);
xor U15642 (N_15642,N_11548,N_13277);
or U15643 (N_15643,N_10415,N_11435);
nor U15644 (N_15644,N_13884,N_13932);
and U15645 (N_15645,N_14198,N_14813);
nand U15646 (N_15646,N_11183,N_11033);
or U15647 (N_15647,N_10712,N_10340);
or U15648 (N_15648,N_13230,N_10417);
nand U15649 (N_15649,N_14605,N_14920);
nand U15650 (N_15650,N_12910,N_10474);
and U15651 (N_15651,N_14309,N_14146);
and U15652 (N_15652,N_14790,N_13789);
nor U15653 (N_15653,N_11211,N_12491);
or U15654 (N_15654,N_10723,N_11484);
xor U15655 (N_15655,N_12715,N_10239);
xnor U15656 (N_15656,N_12058,N_13898);
and U15657 (N_15657,N_14705,N_14179);
or U15658 (N_15658,N_14785,N_10049);
nand U15659 (N_15659,N_14805,N_10065);
nand U15660 (N_15660,N_10345,N_11632);
and U15661 (N_15661,N_13185,N_11856);
or U15662 (N_15662,N_11200,N_12484);
nor U15663 (N_15663,N_10579,N_12610);
nand U15664 (N_15664,N_14665,N_13369);
nand U15665 (N_15665,N_13948,N_11864);
and U15666 (N_15666,N_13287,N_12241);
nand U15667 (N_15667,N_13414,N_11279);
or U15668 (N_15668,N_12651,N_10140);
or U15669 (N_15669,N_12862,N_10612);
or U15670 (N_15670,N_12509,N_11811);
or U15671 (N_15671,N_10863,N_10502);
nor U15672 (N_15672,N_12667,N_14626);
xor U15673 (N_15673,N_11831,N_10182);
nor U15674 (N_15674,N_14923,N_11976);
nand U15675 (N_15675,N_12923,N_13938);
and U15676 (N_15676,N_10816,N_10068);
nor U15677 (N_15677,N_14798,N_14124);
nor U15678 (N_15678,N_10110,N_13164);
and U15679 (N_15679,N_10581,N_14274);
xor U15680 (N_15680,N_10150,N_13443);
or U15681 (N_15681,N_10750,N_13623);
nand U15682 (N_15682,N_13286,N_14007);
or U15683 (N_15683,N_12762,N_12915);
or U15684 (N_15684,N_14542,N_10253);
nand U15685 (N_15685,N_13801,N_14427);
nor U15686 (N_15686,N_10398,N_13759);
xnor U15687 (N_15687,N_10791,N_12279);
or U15688 (N_15688,N_12344,N_11177);
or U15689 (N_15689,N_11562,N_11093);
nand U15690 (N_15690,N_13788,N_10690);
nand U15691 (N_15691,N_11782,N_12209);
or U15692 (N_15692,N_14289,N_12496);
and U15693 (N_15693,N_12176,N_14004);
xnor U15694 (N_15694,N_11144,N_14886);
nor U15695 (N_15695,N_12190,N_14391);
or U15696 (N_15696,N_13213,N_11294);
nor U15697 (N_15697,N_11907,N_14087);
nand U15698 (N_15698,N_12854,N_11581);
nor U15699 (N_15699,N_11108,N_12889);
nand U15700 (N_15700,N_11034,N_13129);
nand U15701 (N_15701,N_11679,N_10790);
or U15702 (N_15702,N_14389,N_12068);
and U15703 (N_15703,N_14823,N_10946);
nor U15704 (N_15704,N_11205,N_14207);
and U15705 (N_15705,N_12005,N_13440);
nor U15706 (N_15706,N_14273,N_13547);
and U15707 (N_15707,N_13211,N_14240);
or U15708 (N_15708,N_10730,N_13795);
and U15709 (N_15709,N_13512,N_11259);
and U15710 (N_15710,N_11874,N_11806);
nor U15711 (N_15711,N_13522,N_10316);
nand U15712 (N_15712,N_12848,N_12281);
or U15713 (N_15713,N_10837,N_10260);
or U15714 (N_15714,N_10953,N_11431);
and U15715 (N_15715,N_13820,N_10951);
or U15716 (N_15716,N_12101,N_11502);
and U15717 (N_15717,N_10098,N_14510);
xor U15718 (N_15718,N_10277,N_12361);
xor U15719 (N_15719,N_13405,N_12666);
and U15720 (N_15720,N_14314,N_14687);
nand U15721 (N_15721,N_11728,N_12838);
nor U15722 (N_15722,N_11295,N_14337);
nand U15723 (N_15723,N_13349,N_13576);
or U15724 (N_15724,N_14917,N_12839);
nor U15725 (N_15725,N_11411,N_12388);
and U15726 (N_15726,N_12805,N_14852);
and U15727 (N_15727,N_12118,N_11906);
nand U15728 (N_15728,N_11805,N_14496);
and U15729 (N_15729,N_11696,N_11359);
nand U15730 (N_15730,N_13219,N_11133);
and U15731 (N_15731,N_14946,N_10741);
or U15732 (N_15732,N_10738,N_11383);
xor U15733 (N_15733,N_10861,N_13244);
nor U15734 (N_15734,N_10619,N_12094);
nand U15735 (N_15735,N_10795,N_11826);
nor U15736 (N_15736,N_13382,N_11603);
nor U15737 (N_15737,N_14242,N_13486);
nand U15738 (N_15738,N_14055,N_13599);
xor U15739 (N_15739,N_14323,N_10536);
or U15740 (N_15740,N_10595,N_14193);
nor U15741 (N_15741,N_13828,N_14983);
and U15742 (N_15742,N_14396,N_13058);
nor U15743 (N_15743,N_13433,N_13635);
nand U15744 (N_15744,N_12320,N_14619);
and U15745 (N_15745,N_13760,N_11763);
nand U15746 (N_15746,N_10034,N_13769);
xor U15747 (N_15747,N_13631,N_12702);
nor U15748 (N_15748,N_10064,N_13811);
or U15749 (N_15749,N_13224,N_14901);
and U15750 (N_15750,N_12471,N_10715);
nand U15751 (N_15751,N_11550,N_13690);
and U15752 (N_15752,N_10114,N_10525);
xnor U15753 (N_15753,N_11735,N_11583);
or U15754 (N_15754,N_14037,N_14896);
nor U15755 (N_15755,N_12669,N_11311);
xor U15756 (N_15756,N_13429,N_11240);
and U15757 (N_15757,N_11053,N_13586);
nor U15758 (N_15758,N_12069,N_10950);
and U15759 (N_15759,N_10765,N_13838);
nand U15760 (N_15760,N_10706,N_12358);
and U15761 (N_15761,N_14875,N_13930);
and U15762 (N_15762,N_14188,N_13439);
xor U15763 (N_15763,N_13575,N_14772);
or U15764 (N_15764,N_12352,N_13451);
and U15765 (N_15765,N_10129,N_10828);
and U15766 (N_15766,N_10495,N_12488);
xnor U15767 (N_15767,N_11861,N_11235);
and U15768 (N_15768,N_13353,N_14491);
or U15769 (N_15769,N_12939,N_12756);
nand U15770 (N_15770,N_14136,N_11256);
nand U15771 (N_15771,N_14039,N_14745);
nor U15772 (N_15772,N_10710,N_14770);
or U15773 (N_15773,N_14143,N_12254);
or U15774 (N_15774,N_14275,N_13713);
nor U15775 (N_15775,N_11360,N_13735);
nor U15776 (N_15776,N_11604,N_12931);
xnor U15777 (N_15777,N_13750,N_10535);
nand U15778 (N_15778,N_14534,N_10009);
xnor U15779 (N_15779,N_10704,N_12021);
and U15780 (N_15780,N_10245,N_13343);
nand U15781 (N_15781,N_10716,N_11096);
nand U15782 (N_15782,N_12212,N_12971);
and U15783 (N_15783,N_14392,N_10121);
nand U15784 (N_15784,N_12077,N_10839);
nand U15785 (N_15785,N_10559,N_12172);
nor U15786 (N_15786,N_10906,N_13267);
or U15787 (N_15787,N_14638,N_14390);
and U15788 (N_15788,N_12543,N_13799);
or U15789 (N_15789,N_10459,N_11810);
nor U15790 (N_15790,N_11736,N_12880);
nand U15791 (N_15791,N_14288,N_10200);
nor U15792 (N_15792,N_10869,N_14063);
and U15793 (N_15793,N_13649,N_11120);
or U15794 (N_15794,N_14589,N_11572);
xor U15795 (N_15795,N_12171,N_14129);
or U15796 (N_15796,N_13910,N_10369);
and U15797 (N_15797,N_12136,N_11528);
or U15798 (N_15798,N_13517,N_14148);
nor U15799 (N_15799,N_12541,N_11018);
and U15800 (N_15800,N_13020,N_12852);
nor U15801 (N_15801,N_13105,N_14147);
xor U15802 (N_15802,N_10626,N_10798);
xnor U15803 (N_15803,N_13961,N_14398);
and U15804 (N_15804,N_11893,N_11626);
xnor U15805 (N_15805,N_12627,N_14361);
and U15806 (N_15806,N_13340,N_14474);
nor U15807 (N_15807,N_13055,N_11180);
nor U15808 (N_15808,N_12799,N_12494);
nand U15809 (N_15809,N_10186,N_13942);
and U15810 (N_15810,N_14726,N_10354);
or U15811 (N_15811,N_10896,N_12360);
nor U15812 (N_15812,N_12257,N_10794);
or U15813 (N_15813,N_12549,N_12969);
nor U15814 (N_15814,N_12447,N_11063);
nor U15815 (N_15815,N_10349,N_14602);
nor U15816 (N_15816,N_11176,N_11005);
nand U15817 (N_15817,N_13040,N_14533);
and U15818 (N_15818,N_10518,N_11827);
nand U15819 (N_15819,N_13552,N_10890);
and U15820 (N_15820,N_14806,N_11742);
nor U15821 (N_15821,N_14378,N_11450);
or U15822 (N_15822,N_12489,N_12104);
and U15823 (N_15823,N_12844,N_10464);
nand U15824 (N_15824,N_13854,N_10211);
and U15825 (N_15825,N_13392,N_10499);
nand U15826 (N_15826,N_11720,N_10822);
or U15827 (N_15827,N_14318,N_12202);
nor U15828 (N_15828,N_12713,N_10136);
nand U15829 (N_15829,N_12814,N_13937);
and U15830 (N_15830,N_12786,N_12692);
or U15831 (N_15831,N_13888,N_10370);
or U15832 (N_15832,N_14132,N_10394);
and U15833 (N_15833,N_14927,N_11246);
nor U15834 (N_15834,N_11915,N_10207);
nand U15835 (N_15835,N_13156,N_12766);
nor U15836 (N_15836,N_11961,N_12566);
or U15837 (N_15837,N_12983,N_10312);
or U15838 (N_15838,N_10966,N_14341);
and U15839 (N_15839,N_14616,N_12001);
nor U15840 (N_15840,N_11227,N_13371);
and U15841 (N_15841,N_14915,N_11167);
nor U15842 (N_15842,N_11717,N_10566);
xnor U15843 (N_15843,N_13892,N_11766);
or U15844 (N_15844,N_12283,N_10756);
and U15845 (N_15845,N_12356,N_10969);
nor U15846 (N_15846,N_11602,N_12565);
and U15847 (N_15847,N_14733,N_10157);
and U15848 (N_15848,N_13933,N_14324);
nand U15849 (N_15849,N_10388,N_14260);
nand U15850 (N_15850,N_14527,N_13513);
or U15851 (N_15851,N_12029,N_13990);
nand U15852 (N_15852,N_12828,N_11203);
or U15853 (N_15853,N_12152,N_13983);
xnor U15854 (N_15854,N_10509,N_12462);
nor U15855 (N_15855,N_14907,N_12018);
xnor U15856 (N_15856,N_10326,N_13141);
and U15857 (N_15857,N_12843,N_12693);
nand U15858 (N_15858,N_13502,N_14402);
nand U15859 (N_15859,N_10493,N_11195);
nand U15860 (N_15860,N_14224,N_11021);
or U15861 (N_15861,N_12861,N_10751);
nand U15862 (N_15862,N_14729,N_10346);
or U15863 (N_15863,N_14819,N_12429);
and U15864 (N_15864,N_13478,N_11598);
nor U15865 (N_15865,N_12894,N_12353);
nor U15866 (N_15866,N_10302,N_14652);
and U15867 (N_15867,N_13717,N_13173);
or U15868 (N_15868,N_12717,N_14761);
or U15869 (N_15869,N_13798,N_12206);
nor U15870 (N_15870,N_10597,N_14406);
or U15871 (N_15871,N_11401,N_14900);
or U15872 (N_15872,N_10940,N_11989);
or U15873 (N_15873,N_13704,N_14394);
nand U15874 (N_15874,N_14140,N_13954);
nor U15875 (N_15875,N_10130,N_12433);
nor U15876 (N_15876,N_14673,N_12975);
and U15877 (N_15877,N_11143,N_14269);
or U15878 (N_15878,N_12990,N_13650);
or U15879 (N_15879,N_10321,N_11639);
nand U15880 (N_15880,N_13743,N_13057);
xor U15881 (N_15881,N_12173,N_13861);
or U15882 (N_15882,N_10256,N_10871);
or U15883 (N_15883,N_12721,N_11731);
xor U15884 (N_15884,N_10719,N_14490);
nor U15885 (N_15885,N_10789,N_13776);
nor U15886 (N_15886,N_12314,N_13458);
nand U15887 (N_15887,N_14183,N_10002);
nand U15888 (N_15888,N_12925,N_12048);
nor U15889 (N_15889,N_11067,N_10124);
and U15890 (N_15890,N_13768,N_14585);
nand U15891 (N_15891,N_13317,N_11600);
nand U15892 (N_15892,N_10733,N_12413);
nor U15893 (N_15893,N_14991,N_11123);
or U15894 (N_15894,N_11941,N_11865);
or U15895 (N_15895,N_10470,N_10761);
and U15896 (N_15896,N_14470,N_13383);
xor U15897 (N_15897,N_12947,N_14564);
or U15898 (N_15898,N_12075,N_12537);
nand U15899 (N_15899,N_12759,N_10887);
xor U15900 (N_15900,N_11014,N_11078);
nor U15901 (N_15901,N_11832,N_13070);
nand U15902 (N_15902,N_13858,N_10800);
or U15903 (N_15903,N_11101,N_11458);
or U15904 (N_15904,N_11741,N_11075);
or U15905 (N_15905,N_13337,N_11122);
nor U15906 (N_15906,N_12100,N_13536);
xnor U15907 (N_15907,N_13744,N_13368);
and U15908 (N_15908,N_13393,N_14989);
nor U15909 (N_15909,N_12988,N_14360);
and U15910 (N_15910,N_11000,N_10073);
nor U15911 (N_15911,N_12449,N_14615);
or U15912 (N_15912,N_12406,N_10766);
or U15913 (N_15913,N_11841,N_10276);
nand U15914 (N_15914,N_14882,N_11085);
nor U15915 (N_15915,N_13778,N_12665);
nor U15916 (N_15916,N_14108,N_12476);
or U15917 (N_15917,N_12294,N_12645);
xnor U15918 (N_15918,N_14762,N_12293);
xor U15919 (N_15919,N_13764,N_10868);
xnor U15920 (N_15920,N_13669,N_13113);
or U15921 (N_15921,N_13514,N_13178);
or U15922 (N_15922,N_14022,N_13457);
xnor U15923 (N_15923,N_11747,N_11557);
nor U15924 (N_15924,N_11756,N_10746);
nand U15925 (N_15925,N_10881,N_10188);
nor U15926 (N_15926,N_14731,N_12801);
nand U15927 (N_15927,N_14888,N_11118);
nand U15928 (N_15928,N_14467,N_11788);
and U15929 (N_15929,N_13924,N_10679);
xor U15930 (N_15930,N_10461,N_12768);
nor U15931 (N_15931,N_12900,N_12561);
or U15932 (N_15932,N_10571,N_10573);
and U15933 (N_15933,N_11783,N_12285);
or U15934 (N_15934,N_14455,N_10684);
nor U15935 (N_15935,N_13775,N_12113);
nor U15936 (N_15936,N_14209,N_10931);
nand U15937 (N_15937,N_13278,N_10075);
nand U15938 (N_15938,N_13807,N_12751);
or U15939 (N_15939,N_14680,N_13198);
nand U15940 (N_15940,N_10426,N_12460);
nor U15941 (N_15941,N_12984,N_14157);
nand U15942 (N_15942,N_10507,N_13194);
nor U15943 (N_15943,N_14038,N_12513);
and U15944 (N_15944,N_14975,N_13300);
xnor U15945 (N_15945,N_14150,N_12363);
and U15946 (N_15946,N_10804,N_14595);
nand U15947 (N_15947,N_11666,N_13330);
or U15948 (N_15948,N_12752,N_10029);
nand U15949 (N_15949,N_12236,N_14758);
nor U15950 (N_15950,N_13845,N_14531);
or U15951 (N_15951,N_14808,N_12883);
nor U15952 (N_15952,N_13563,N_10729);
or U15953 (N_15953,N_10914,N_11840);
and U15954 (N_15954,N_10395,N_10763);
xor U15955 (N_15955,N_10419,N_10342);
nand U15956 (N_15956,N_10194,N_10537);
nand U15957 (N_15957,N_12767,N_12431);
nand U15958 (N_15958,N_14126,N_14969);
nand U15959 (N_15959,N_14812,N_11942);
xnor U15960 (N_15960,N_13220,N_11352);
and U15961 (N_15961,N_12523,N_12396);
xnor U15962 (N_15962,N_11767,N_13001);
xor U15963 (N_15963,N_11534,N_12650);
or U15964 (N_15964,N_11977,N_11347);
nor U15965 (N_15965,N_14486,N_14248);
nand U15966 (N_15966,N_11198,N_13243);
and U15967 (N_15967,N_10134,N_14556);
and U15968 (N_15968,N_11537,N_11970);
nor U15969 (N_15969,N_12127,N_12371);
nor U15970 (N_15970,N_13043,N_11777);
and U15971 (N_15971,N_13981,N_13134);
nor U15972 (N_15972,N_11845,N_10563);
nand U15973 (N_15973,N_11894,N_14346);
and U15974 (N_15974,N_14050,N_11475);
xnor U15975 (N_15975,N_10089,N_10047);
or U15976 (N_15976,N_10362,N_12611);
nor U15977 (N_15977,N_10532,N_14956);
or U15978 (N_15978,N_10630,N_13851);
or U15979 (N_15979,N_10734,N_12668);
nor U15980 (N_15980,N_13168,N_13233);
nor U15981 (N_15981,N_12999,N_11044);
nor U15982 (N_15982,N_12506,N_12599);
or U15983 (N_15983,N_12876,N_11429);
nor U15984 (N_15984,N_12584,N_14387);
and U15985 (N_15985,N_10196,N_11949);
or U15986 (N_15986,N_14645,N_12193);
nand U15987 (N_15987,N_14592,N_12333);
and U15988 (N_15988,N_12448,N_12864);
nand U15989 (N_15989,N_12928,N_13925);
and U15990 (N_15990,N_14440,N_11680);
nand U15991 (N_15991,N_14941,N_11673);
nand U15992 (N_15992,N_11529,N_12201);
or U15993 (N_15993,N_11554,N_11663);
nor U15994 (N_15994,N_14912,N_13806);
nand U15995 (N_15995,N_13928,N_13420);
xor U15996 (N_15996,N_14251,N_10070);
xor U15997 (N_15997,N_11723,N_14794);
and U15998 (N_15998,N_10659,N_11924);
nor U15999 (N_15999,N_14997,N_14988);
and U16000 (N_16000,N_12467,N_12775);
nor U16001 (N_16001,N_11835,N_11631);
or U16002 (N_16002,N_13206,N_10894);
or U16003 (N_16003,N_10825,N_13505);
or U16004 (N_16004,N_10793,N_12108);
nand U16005 (N_16005,N_10106,N_12134);
nand U16006 (N_16006,N_12595,N_12996);
nand U16007 (N_16007,N_10862,N_13362);
or U16008 (N_16008,N_11380,N_11955);
and U16009 (N_16009,N_13065,N_11393);
nand U16010 (N_16010,N_10801,N_13687);
xor U16011 (N_16011,N_10942,N_13027);
or U16012 (N_16012,N_10283,N_14609);
and U16013 (N_16013,N_14951,N_13973);
and U16014 (N_16014,N_12962,N_14083);
and U16015 (N_16015,N_13108,N_11521);
nand U16016 (N_16016,N_11425,N_13048);
nor U16017 (N_16017,N_12656,N_11566);
nand U16018 (N_16018,N_13152,N_11592);
nor U16019 (N_16019,N_10647,N_11718);
and U16020 (N_16020,N_14320,N_10265);
and U16021 (N_16021,N_11724,N_11676);
xnor U16022 (N_16022,N_12234,N_10923);
nand U16023 (N_16023,N_13571,N_14885);
xor U16024 (N_16024,N_13255,N_14133);
and U16025 (N_16025,N_11846,N_14218);
nor U16026 (N_16026,N_10711,N_12012);
nor U16027 (N_16027,N_13891,N_14878);
xnor U16028 (N_16028,N_10430,N_14848);
or U16029 (N_16029,N_10082,N_12585);
and U16030 (N_16030,N_14653,N_12487);
nand U16031 (N_16031,N_13180,N_14031);
nor U16032 (N_16032,N_14759,N_13235);
and U16033 (N_16033,N_13772,N_11923);
nand U16034 (N_16034,N_13654,N_14077);
and U16035 (N_16035,N_13442,N_10527);
nand U16036 (N_16036,N_11303,N_14493);
nand U16037 (N_16037,N_13568,N_11754);
xor U16038 (N_16038,N_11436,N_14914);
and U16039 (N_16039,N_14092,N_14870);
nand U16040 (N_16040,N_10483,N_14417);
nor U16041 (N_16041,N_10492,N_11611);
nor U16042 (N_16042,N_13822,N_10467);
and U16043 (N_16043,N_11985,N_13611);
nor U16044 (N_16044,N_13422,N_13610);
or U16045 (N_16045,N_14049,N_10924);
nand U16046 (N_16046,N_11587,N_12618);
nand U16047 (N_16047,N_12451,N_10674);
nor U16048 (N_16048,N_10240,N_13666);
nand U16049 (N_16049,N_13408,N_10545);
and U16050 (N_16050,N_14385,N_13503);
or U16051 (N_16051,N_11057,N_14284);
or U16052 (N_16052,N_11690,N_12437);
nor U16053 (N_16053,N_13617,N_14356);
nand U16054 (N_16054,N_14329,N_10171);
xnor U16055 (N_16055,N_14929,N_13423);
nor U16056 (N_16056,N_12654,N_14367);
and U16057 (N_16057,N_10101,N_12677);
xnor U16058 (N_16058,N_10359,N_12480);
nor U16059 (N_16059,N_11511,N_11427);
and U16060 (N_16060,N_14890,N_11282);
xnor U16061 (N_16061,N_13214,N_11820);
or U16062 (N_16062,N_11196,N_14741);
nor U16063 (N_16063,N_12564,N_12345);
nand U16064 (N_16064,N_11312,N_14110);
nand U16065 (N_16065,N_10678,N_10523);
or U16066 (N_16066,N_12858,N_11625);
and U16067 (N_16067,N_11588,N_14998);
and U16068 (N_16068,N_13190,N_13841);
nor U16069 (N_16069,N_14357,N_11990);
xnor U16070 (N_16070,N_14627,N_10206);
and U16071 (N_16071,N_14212,N_11699);
nand U16072 (N_16072,N_11477,N_13409);
nor U16073 (N_16073,N_10195,N_10758);
or U16074 (N_16074,N_14141,N_14792);
nor U16075 (N_16075,N_12841,N_12845);
nand U16076 (N_16076,N_12141,N_13076);
nor U16077 (N_16077,N_11278,N_10305);
and U16078 (N_16078,N_12304,N_12034);
and U16079 (N_16079,N_13354,N_10576);
xor U16080 (N_16080,N_10548,N_11220);
and U16081 (N_16081,N_14600,N_12379);
nand U16082 (N_16082,N_12359,N_11778);
and U16083 (N_16083,N_10313,N_14630);
nor U16084 (N_16084,N_14100,N_14340);
nor U16085 (N_16085,N_14569,N_12711);
xor U16086 (N_16086,N_11035,N_10934);
and U16087 (N_16087,N_10099,N_10594);
nor U16088 (N_16088,N_14816,N_14902);
nand U16089 (N_16089,N_13590,N_12114);
and U16090 (N_16090,N_11171,N_12207);
nor U16091 (N_16091,N_11772,N_10858);
nand U16092 (N_16092,N_12556,N_13358);
nor U16093 (N_16093,N_12761,N_12478);
or U16094 (N_16094,N_11174,N_14102);
and U16095 (N_16095,N_11614,N_13783);
and U16096 (N_16096,N_13465,N_11447);
xnor U16097 (N_16097,N_13309,N_10397);
or U16098 (N_16098,N_14355,N_10740);
or U16099 (N_16099,N_13699,N_12792);
nand U16100 (N_16100,N_14782,N_14578);
and U16101 (N_16101,N_12503,N_14338);
and U16102 (N_16102,N_10165,N_12602);
or U16103 (N_16103,N_11577,N_13430);
nand U16104 (N_16104,N_14458,N_11216);
nand U16105 (N_16105,N_12306,N_12648);
nor U16106 (N_16106,N_11933,N_13496);
nand U16107 (N_16107,N_13979,N_14707);
or U16108 (N_16108,N_10060,N_12225);
and U16109 (N_16109,N_10947,N_11586);
nor U16110 (N_16110,N_11501,N_13691);
nand U16111 (N_16111,N_11868,N_13315);
nand U16112 (N_16112,N_13199,N_12504);
nand U16113 (N_16113,N_13953,N_13551);
nand U16114 (N_16114,N_13934,N_12724);
or U16115 (N_16115,N_13091,N_10147);
and U16116 (N_16116,N_12473,N_13539);
nor U16117 (N_16117,N_10727,N_11309);
xnor U16118 (N_16118,N_14744,N_12365);
nor U16119 (N_16119,N_11221,N_10688);
or U16120 (N_16120,N_11641,N_14405);
nor U16121 (N_16121,N_10491,N_11913);
nor U16122 (N_16122,N_10123,N_12501);
or U16123 (N_16123,N_10176,N_13276);
nand U16124 (N_16124,N_14736,N_10005);
nor U16125 (N_16125,N_13094,N_12350);
nand U16126 (N_16126,N_14779,N_12982);
and U16127 (N_16127,N_14737,N_12935);
nand U16128 (N_16128,N_14719,N_12816);
nand U16129 (N_16129,N_12920,N_12138);
and U16130 (N_16130,N_13574,N_14299);
nor U16131 (N_16131,N_13195,N_10185);
or U16132 (N_16132,N_13380,N_13998);
nor U16133 (N_16133,N_14079,N_11406);
nor U16134 (N_16134,N_12605,N_13441);
and U16135 (N_16135,N_14588,N_12492);
nand U16136 (N_16136,N_12047,N_11859);
nand U16137 (N_16137,N_12945,N_14335);
nor U16138 (N_16138,N_10879,N_12966);
nand U16139 (N_16139,N_14211,N_11262);
and U16140 (N_16140,N_11407,N_13132);
and U16141 (N_16141,N_13943,N_13081);
nor U16142 (N_16142,N_11965,N_10577);
and U16143 (N_16143,N_12758,N_11790);
or U16144 (N_16144,N_13870,N_10438);
or U16145 (N_16145,N_11986,N_14765);
nor U16146 (N_16146,N_13436,N_13485);
nand U16147 (N_16147,N_12727,N_12998);
or U16148 (N_16148,N_13700,N_11793);
or U16149 (N_16149,N_13510,N_13964);
and U16150 (N_16150,N_14352,N_13929);
nor U16151 (N_16151,N_11702,N_11812);
and U16152 (N_16152,N_13281,N_10383);
nand U16153 (N_16153,N_11225,N_10670);
and U16154 (N_16154,N_14894,N_11186);
or U16155 (N_16155,N_13874,N_13086);
xor U16156 (N_16156,N_11334,N_10637);
xor U16157 (N_16157,N_11857,N_10236);
nand U16158 (N_16158,N_14670,N_14933);
nor U16159 (N_16159,N_11638,N_14206);
nand U16160 (N_16160,N_13399,N_11400);
nand U16161 (N_16161,N_10617,N_11185);
nor U16162 (N_16162,N_12993,N_12307);
nand U16163 (N_16163,N_10504,N_10977);
and U16164 (N_16164,N_12592,N_10439);
and U16165 (N_16165,N_13572,N_13561);
or U16166 (N_16166,N_12091,N_13802);
nand U16167 (N_16167,N_14027,N_12797);
nand U16168 (N_16168,N_11154,N_11804);
nand U16169 (N_16169,N_11156,N_10596);
and U16170 (N_16170,N_11665,N_11001);
nand U16171 (N_16171,N_11797,N_10809);
and U16172 (N_16172,N_12678,N_13316);
and U16173 (N_16173,N_13010,N_12081);
and U16174 (N_16174,N_11371,N_10127);
or U16175 (N_16175,N_11230,N_10445);
nand U16176 (N_16176,N_10069,N_11591);
nand U16177 (N_16177,N_10190,N_10948);
nor U16178 (N_16178,N_11088,N_12593);
nand U16179 (N_16179,N_10913,N_12936);
or U16180 (N_16180,N_11905,N_11373);
or U16181 (N_16181,N_12177,N_12558);
xnor U16182 (N_16182,N_14281,N_11520);
and U16183 (N_16183,N_11672,N_12158);
and U16184 (N_16184,N_13360,N_13875);
or U16185 (N_16185,N_14345,N_13424);
xor U16186 (N_16186,N_11385,N_14507);
nor U16187 (N_16187,N_13519,N_13636);
nor U16188 (N_16188,N_10970,N_11776);
and U16189 (N_16189,N_10722,N_12511);
nor U16190 (N_16190,N_10125,N_12679);
nor U16191 (N_16191,N_11058,N_13533);
nand U16192 (N_16192,N_11191,N_11444);
xnor U16193 (N_16193,N_12188,N_14252);
nor U16194 (N_16194,N_13413,N_12025);
nor U16195 (N_16195,N_14677,N_12781);
nand U16196 (N_16196,N_14173,N_12486);
or U16197 (N_16197,N_12596,N_12664);
nand U16198 (N_16198,N_12110,N_11686);
xnor U16199 (N_16199,N_12256,N_14810);
or U16200 (N_16200,N_14696,N_11698);
nor U16201 (N_16201,N_14014,N_13785);
and U16202 (N_16202,N_13553,N_13766);
and U16203 (N_16203,N_10836,N_14967);
nand U16204 (N_16204,N_10285,N_10158);
or U16205 (N_16205,N_14795,N_10651);
nor U16206 (N_16206,N_12922,N_14781);
nor U16207 (N_16207,N_11168,N_12263);
and U16208 (N_16208,N_10219,N_10533);
or U16209 (N_16209,N_12707,N_12381);
or U16210 (N_16210,N_13039,N_12788);
nor U16211 (N_16211,N_11830,N_11378);
xnor U16212 (N_16212,N_14691,N_14423);
xor U16213 (N_16213,N_14985,N_10883);
or U16214 (N_16214,N_11158,N_11987);
nand U16215 (N_16215,N_14488,N_11119);
nor U16216 (N_16216,N_13250,N_13991);
nand U16217 (N_16217,N_10392,N_11382);
and U16218 (N_16218,N_13347,N_11332);
or U16219 (N_16219,N_11151,N_14067);
xnor U16220 (N_16220,N_14181,N_12961);
or U16221 (N_16221,N_14202,N_10728);
xor U16222 (N_16222,N_13578,N_10585);
nor U16223 (N_16223,N_14689,N_10142);
nand U16224 (N_16224,N_14328,N_12837);
nor U16225 (N_16225,N_11419,N_14714);
nand U16226 (N_16226,N_12906,N_14701);
nand U16227 (N_16227,N_13384,N_13163);
nand U16228 (N_16228,N_14930,N_13721);
and U16229 (N_16229,N_13740,N_13919);
nand U16230 (N_16230,N_10664,N_10932);
and U16231 (N_16231,N_14966,N_11300);
or U16232 (N_16232,N_13404,N_13730);
nor U16233 (N_16233,N_11026,N_14333);
nor U16234 (N_16234,N_14071,N_12477);
nor U16235 (N_16235,N_11348,N_10223);
or U16236 (N_16236,N_12878,N_10962);
or U16237 (N_16237,N_13885,N_13974);
nand U16238 (N_16238,N_13570,N_11329);
or U16239 (N_16239,N_11649,N_12875);
nor U16240 (N_16240,N_12870,N_12615);
xnor U16241 (N_16241,N_13900,N_13098);
or U16242 (N_16242,N_13712,N_14094);
and U16243 (N_16243,N_13676,N_13207);
and U16244 (N_16244,N_12719,N_12850);
and U16245 (N_16245,N_10234,N_13976);
nand U16246 (N_16246,N_14276,N_11710);
nor U16247 (N_16247,N_14990,N_11978);
nand U16248 (N_16248,N_10252,N_13718);
nor U16249 (N_16249,N_10051,N_14268);
xor U16250 (N_16250,N_10677,N_12659);
nor U16251 (N_16251,N_11386,N_11871);
nor U16252 (N_16252,N_12213,N_13603);
and U16253 (N_16253,N_12970,N_10485);
or U16254 (N_16254,N_13030,N_10785);
nand U16255 (N_16255,N_11497,N_13588);
or U16256 (N_16256,N_10574,N_10676);
nand U16257 (N_16257,N_13209,N_14057);
nand U16258 (N_16258,N_13282,N_14685);
or U16259 (N_16259,N_14404,N_12440);
nor U16260 (N_16260,N_13688,N_10524);
nor U16261 (N_16261,N_14287,N_10226);
xor U16262 (N_16262,N_10033,N_11166);
nand U16263 (N_16263,N_14321,N_12525);
nand U16264 (N_16264,N_12116,N_11822);
nand U16265 (N_16265,N_12575,N_11445);
or U16266 (N_16266,N_10282,N_12417);
and U16267 (N_16267,N_14821,N_12003);
nand U16268 (N_16268,N_10449,N_13969);
nor U16269 (N_16269,N_13711,N_12051);
nand U16270 (N_16270,N_14122,N_10973);
xnor U16271 (N_16271,N_12903,N_10910);
or U16272 (N_16272,N_10141,N_11068);
or U16273 (N_16273,N_11643,N_12725);
nand U16274 (N_16274,N_14911,N_14970);
and U16275 (N_16275,N_12882,N_13893);
nor U16276 (N_16276,N_10373,N_10824);
nor U16277 (N_16277,N_14672,N_14538);
or U16278 (N_16278,N_11709,N_13288);
xnor U16279 (N_16279,N_14613,N_11179);
nor U16280 (N_16280,N_12547,N_13527);
nand U16281 (N_16281,N_13782,N_10799);
nand U16282 (N_16282,N_14558,N_13259);
nor U16283 (N_16283,N_12096,N_10657);
nor U16284 (N_16284,N_11781,N_11917);
and U16285 (N_16285,N_10849,N_11008);
nand U16286 (N_16286,N_10958,N_12662);
or U16287 (N_16287,N_13455,N_12146);
and U16288 (N_16288,N_14365,N_11899);
nor U16289 (N_16289,N_12532,N_14634);
and U16290 (N_16290,N_12465,N_12253);
nor U16291 (N_16291,N_10916,N_10386);
xnor U16292 (N_16292,N_14187,N_14483);
and U16293 (N_16293,N_13112,N_12348);
or U16294 (N_16294,N_13728,N_13935);
nand U16295 (N_16295,N_11953,N_12829);
and U16296 (N_16296,N_11392,N_11236);
and U16297 (N_16297,N_11313,N_13792);
or U16298 (N_16298,N_14867,N_12908);
and U16299 (N_16299,N_14582,N_14047);
and U16300 (N_16300,N_11635,N_11594);
nor U16301 (N_16301,N_13004,N_12639);
xnor U16302 (N_16302,N_11173,N_11375);
or U16303 (N_16303,N_13472,N_13341);
or U16304 (N_16304,N_14936,N_14976);
or U16305 (N_16305,N_12913,N_13361);
nor U16306 (N_16306,N_10360,N_13918);
xor U16307 (N_16307,N_12857,N_12732);
and U16308 (N_16308,N_13585,N_14695);
nor U16309 (N_16309,N_12972,N_13901);
or U16310 (N_16310,N_11010,N_11349);
nand U16311 (N_16311,N_11446,N_12524);
and U16312 (N_16312,N_11009,N_12180);
or U16313 (N_16313,N_10943,N_12033);
and U16314 (N_16314,N_14064,N_10408);
xor U16315 (N_16315,N_11412,N_10389);
or U16316 (N_16316,N_13714,N_13066);
nor U16317 (N_16317,N_10442,N_10286);
nor U16318 (N_16318,N_13229,N_10672);
or U16319 (N_16319,N_10901,N_12929);
or U16320 (N_16320,N_11847,N_12372);
and U16321 (N_16321,N_14713,N_12744);
and U16322 (N_16322,N_13363,N_11925);
or U16323 (N_16323,N_11715,N_13400);
nor U16324 (N_16324,N_13909,N_12757);
nor U16325 (N_16325,N_13068,N_10960);
nor U16326 (N_16326,N_11395,N_12834);
and U16327 (N_16327,N_11959,N_14957);
nor U16328 (N_16328,N_10606,N_14502);
nand U16329 (N_16329,N_11569,N_14354);
nor U16330 (N_16330,N_14778,N_11283);
nand U16331 (N_16331,N_11339,N_11247);
nand U16332 (N_16332,N_12912,N_14016);
and U16333 (N_16333,N_14746,N_12292);
or U16334 (N_16334,N_10301,N_11991);
nand U16335 (N_16335,N_11124,N_10232);
or U16336 (N_16336,N_11471,N_12600);
nand U16337 (N_16337,N_14579,N_14940);
or U16338 (N_16338,N_13292,N_11298);
and U16339 (N_16339,N_11099,N_12689);
and U16340 (N_16340,N_11193,N_13026);
or U16341 (N_16341,N_12481,N_11668);
nor U16342 (N_16342,N_13722,N_14263);
or U16343 (N_16343,N_12790,N_12705);
nor U16344 (N_16344,N_11651,N_12911);
or U16345 (N_16345,N_10522,N_11030);
xor U16346 (N_16346,N_10198,N_10792);
and U16347 (N_16347,N_11634,N_11995);
or U16348 (N_16348,N_10084,N_12221);
nand U16349 (N_16349,N_11988,N_11428);
and U16350 (N_16350,N_14984,N_12741);
xnor U16351 (N_16351,N_14846,N_13406);
or U16352 (N_16352,N_12342,N_13187);
xnor U16353 (N_16353,N_13088,N_12657);
nor U16354 (N_16354,N_13017,N_11271);
or U16355 (N_16355,N_13542,N_10570);
nor U16356 (N_16356,N_13389,N_13327);
nor U16357 (N_16357,N_10329,N_11465);
xnor U16358 (N_16358,N_10530,N_12125);
nand U16359 (N_16359,N_14114,N_11750);
nor U16360 (N_16360,N_14711,N_12088);
nand U16361 (N_16361,N_14760,N_13097);
or U16362 (N_16362,N_11217,N_13084);
nand U16363 (N_16363,N_14177,N_11877);
or U16364 (N_16364,N_11032,N_11290);
nor U16365 (N_16365,N_13593,N_14437);
or U16366 (N_16366,N_13012,N_10686);
nand U16367 (N_16367,N_13911,N_11695);
and U16368 (N_16368,N_11268,N_13987);
xnor U16369 (N_16369,N_11801,N_12512);
or U16370 (N_16370,N_13060,N_14245);
or U16371 (N_16371,N_10803,N_12598);
and U16372 (N_16372,N_11854,N_11891);
and U16373 (N_16373,N_11414,N_11834);
nand U16374 (N_16374,N_12295,N_11786);
and U16375 (N_16375,N_14679,N_11403);
nor U16376 (N_16376,N_12607,N_11381);
and U16377 (N_16377,N_10488,N_13225);
xnor U16378 (N_16378,N_13956,N_10044);
or U16379 (N_16379,N_12076,N_10628);
and U16380 (N_16380,N_12873,N_11561);
or U16381 (N_16381,N_14015,N_11760);
nand U16382 (N_16382,N_13115,N_13907);
nor U16383 (N_16383,N_14431,N_13868);
or U16384 (N_16384,N_12630,N_14041);
nand U16385 (N_16385,N_10768,N_10848);
or U16386 (N_16386,N_10665,N_13890);
nor U16387 (N_16387,N_12956,N_11615);
and U16388 (N_16388,N_13773,N_10151);
nor U16389 (N_16389,N_13605,N_11527);
xnor U16390 (N_16390,N_14822,N_14500);
xnor U16391 (N_16391,N_14655,N_14364);
or U16392 (N_16392,N_12014,N_10846);
or U16393 (N_16393,N_14921,N_11619);
or U16394 (N_16394,N_13114,N_12435);
or U16395 (N_16395,N_13186,N_14312);
or U16396 (N_16396,N_13771,N_12265);
or U16397 (N_16397,N_14199,N_13064);
nand U16398 (N_16398,N_11302,N_14506);
nand U16399 (N_16399,N_10603,N_14399);
nor U16400 (N_16400,N_13912,N_11684);
nand U16401 (N_16401,N_11242,N_14298);
or U16402 (N_16402,N_10227,N_12530);
xnor U16403 (N_16403,N_13708,N_13827);
or U16404 (N_16404,N_14308,N_12949);
nand U16405 (N_16405,N_12264,N_13003);
and U16406 (N_16406,N_12560,N_12987);
nor U16407 (N_16407,N_14601,N_10694);
or U16408 (N_16408,N_11253,N_13262);
or U16409 (N_16409,N_10473,N_13673);
xor U16410 (N_16410,N_13630,N_14749);
or U16411 (N_16411,N_11181,N_13856);
and U16412 (N_16412,N_10841,N_10077);
nor U16413 (N_16413,N_12410,N_11508);
nor U16414 (N_16414,N_11650,N_13401);
nor U16415 (N_16415,N_12062,N_12000);
nand U16416 (N_16416,N_11701,N_10999);
nand U16417 (N_16417,N_14111,N_10572);
nand U16418 (N_16418,N_11571,N_11982);
and U16419 (N_16419,N_13236,N_13787);
nand U16420 (N_16420,N_13749,N_10656);
and U16421 (N_16421,N_10778,N_13686);
nor U16422 (N_16422,N_13515,N_13378);
or U16423 (N_16423,N_12099,N_14835);
or U16424 (N_16424,N_10542,N_12932);
nor U16425 (N_16425,N_12776,N_14924);
and U16426 (N_16426,N_10357,N_12916);
nor U16427 (N_16427,N_14008,N_12023);
and U16428 (N_16428,N_11862,N_10988);
or U16429 (N_16429,N_14397,N_11374);
and U16430 (N_16430,N_14466,N_10320);
nor U16431 (N_16431,N_14473,N_10956);
xor U16432 (N_16432,N_12336,N_14717);
xor U16433 (N_16433,N_13052,N_13543);
nor U16434 (N_16434,N_14259,N_12869);
nor U16435 (N_16435,N_13434,N_11439);
and U16436 (N_16436,N_13994,N_12635);
and U16437 (N_16437,N_10796,N_10162);
nor U16438 (N_16438,N_10294,N_11758);
and U16439 (N_16439,N_11440,N_10324);
or U16440 (N_16440,N_12195,N_13402);
or U16441 (N_16441,N_12789,N_11319);
or U16442 (N_16442,N_14766,N_10391);
nand U16443 (N_16443,N_10167,N_11306);
or U16444 (N_16444,N_11017,N_13158);
and U16445 (N_16445,N_11609,N_10062);
or U16446 (N_16446,N_12443,N_10850);
nand U16447 (N_16447,N_14955,N_12377);
or U16448 (N_16448,N_13445,N_14543);
nor U16449 (N_16449,N_12178,N_10023);
and U16450 (N_16450,N_10017,N_10702);
or U16451 (N_16451,N_12733,N_12704);
or U16452 (N_16452,N_12672,N_11192);
and U16453 (N_16453,N_10624,N_14445);
xnor U16454 (N_16454,N_10709,N_10056);
or U16455 (N_16455,N_12959,N_14555);
nor U16456 (N_16456,N_11098,N_12246);
nor U16457 (N_16457,N_12203,N_13460);
or U16458 (N_16458,N_14461,N_11163);
xnor U16459 (N_16459,N_14608,N_14880);
and U16460 (N_16460,N_13449,N_12553);
and U16461 (N_16461,N_13461,N_12343);
or U16462 (N_16462,N_12006,N_10967);
nand U16463 (N_16463,N_10209,N_11091);
nand U16464 (N_16464,N_11102,N_11146);
nand U16465 (N_16465,N_12898,N_11136);
nand U16466 (N_16466,N_13045,N_12736);
nand U16467 (N_16467,N_11149,N_12229);
or U16468 (N_16468,N_12259,N_10096);
or U16469 (N_16469,N_12886,N_11441);
and U16470 (N_16470,N_11802,N_10148);
or U16471 (N_16471,N_13446,N_10444);
nand U16472 (N_16472,N_13294,N_14013);
and U16473 (N_16473,N_13000,N_13078);
nor U16474 (N_16474,N_14671,N_10580);
and U16475 (N_16475,N_11544,N_11792);
nand U16476 (N_16476,N_12239,N_11748);
and U16477 (N_16477,N_12760,N_10599);
nor U16478 (N_16478,N_14076,N_10591);
nor U16479 (N_16479,N_13062,N_10475);
xor U16480 (N_16480,N_14617,N_10363);
or U16481 (N_16481,N_12830,N_13731);
nand U16482 (N_16482,N_14571,N_13002);
or U16483 (N_16483,N_10448,N_11022);
or U16484 (N_16484,N_13962,N_12623);
or U16485 (N_16485,N_13725,N_13473);
xnor U16486 (N_16486,N_13594,N_12059);
xnor U16487 (N_16487,N_10233,N_14526);
and U16488 (N_16488,N_14232,N_11866);
or U16489 (N_16489,N_11045,N_12332);
nand U16490 (N_16490,N_10015,N_13972);
nor U16491 (N_16491,N_14017,N_13616);
nor U16492 (N_16492,N_12041,N_10425);
or U16493 (N_16493,N_11692,N_10325);
nor U16494 (N_16494,N_11076,N_10636);
nor U16495 (N_16495,N_14492,N_10028);
nor U16496 (N_16496,N_11399,N_12112);
nor U16497 (N_16497,N_13739,N_14521);
nor U16498 (N_16498,N_13305,N_14159);
nand U16499 (N_16499,N_10298,N_11887);
or U16500 (N_16500,N_14594,N_14504);
nor U16501 (N_16501,N_10859,N_12452);
nor U16502 (N_16502,N_14768,N_12498);
or U16503 (N_16503,N_10689,N_11261);
or U16504 (N_16504,N_11762,N_11815);
nor U16505 (N_16505,N_10963,N_13291);
and U16506 (N_16506,N_14572,N_14583);
or U16507 (N_16507,N_11379,N_10366);
and U16508 (N_16508,N_14377,N_11817);
xnor U16509 (N_16509,N_12660,N_12390);
nand U16510 (N_16510,N_12063,N_10842);
xnor U16511 (N_16511,N_13497,N_12339);
and U16512 (N_16512,N_10754,N_10797);
and U16513 (N_16513,N_12272,N_11885);
or U16514 (N_16514,N_14001,N_12728);
and U16515 (N_16515,N_13479,N_14942);
or U16516 (N_16516,N_14449,N_13604);
and U16517 (N_16517,N_12082,N_14972);
xnor U16518 (N_16518,N_14185,N_11879);
and U16519 (N_16519,N_13684,N_10344);
nor U16520 (N_16520,N_11948,N_11890);
and U16521 (N_16521,N_10076,N_10118);
nor U16522 (N_16522,N_13598,N_11549);
nand U16523 (N_16523,N_13589,N_14751);
nand U16524 (N_16524,N_11671,N_14830);
nor U16525 (N_16525,N_10295,N_12690);
nand U16526 (N_16526,N_14290,N_11354);
xnor U16527 (N_16527,N_13289,N_12297);
nand U16528 (N_16528,N_13049,N_11825);
xor U16529 (N_16529,N_14712,N_13794);
or U16530 (N_16530,N_10703,N_13675);
nor U16531 (N_16531,N_10586,N_11365);
and U16532 (N_16532,N_12224,N_14438);
nand U16533 (N_16533,N_13641,N_10812);
nor U16534 (N_16534,N_14469,N_12210);
and U16535 (N_16535,N_14249,N_12649);
nor U16536 (N_16536,N_14160,N_12590);
nand U16537 (N_16537,N_10102,N_14282);
xor U16538 (N_16538,N_13306,N_11627);
and U16539 (N_16539,N_11505,N_13454);
or U16540 (N_16540,N_12606,N_13545);
nand U16541 (N_16541,N_12950,N_11353);
nand U16542 (N_16542,N_14460,N_10217);
nand U16543 (N_16543,N_10007,N_11437);
nor U16544 (N_16544,N_13489,N_14200);
nor U16545 (N_16545,N_14565,N_11956);
nand U16546 (N_16546,N_12893,N_10878);
or U16547 (N_16547,N_10387,N_14965);
nand U16548 (N_16548,N_12319,N_10166);
nor U16549 (N_16549,N_10482,N_13674);
nand U16550 (N_16550,N_11317,N_11670);
nand U16551 (N_16551,N_13780,N_11983);
or U16552 (N_16552,N_11327,N_12144);
or U16553 (N_16553,N_13825,N_13754);
or U16554 (N_16554,N_12812,N_14121);
nor U16555 (N_16555,N_11546,N_10427);
or U16556 (N_16556,N_13549,N_14518);
nand U16557 (N_16557,N_14155,N_13655);
nor U16558 (N_16558,N_13041,N_14937);
nand U16559 (N_16559,N_11389,N_12941);
nor U16560 (N_16560,N_12416,N_12572);
and U16561 (N_16561,N_12684,N_14401);
and U16562 (N_16562,N_14130,N_10695);
or U16563 (N_16563,N_14350,N_10713);
or U16564 (N_16564,N_10930,N_12551);
or U16565 (N_16565,N_13228,N_12315);
nand U16566 (N_16566,N_12773,N_13521);
nand U16567 (N_16567,N_11513,N_12191);
or U16568 (N_16568,N_12905,N_13751);
xnor U16569 (N_16569,N_11999,N_12681);
nand U16570 (N_16570,N_12591,N_10204);
nand U16571 (N_16571,N_13344,N_11432);
xnor U16572 (N_16572,N_13800,N_10126);
nand U16573 (N_16573,N_10714,N_13493);
and U16574 (N_16574,N_13897,N_10937);
nand U16575 (N_16575,N_13111,N_11250);
nor U16576 (N_16576,N_10361,N_12140);
and U16577 (N_16577,N_13756,N_14873);
or U16578 (N_16578,N_14464,N_11775);
or U16579 (N_16579,N_14738,N_13029);
xnor U16580 (N_16580,N_11323,N_14540);
nand U16581 (N_16581,N_14661,N_10027);
nor U16582 (N_16582,N_12601,N_12973);
and U16583 (N_16583,N_14286,N_12747);
or U16584 (N_16584,N_12890,N_12090);
and U16585 (N_16585,N_10845,N_14109);
and U16586 (N_16586,N_10717,N_10649);
and U16587 (N_16587,N_12832,N_13332);
xor U16588 (N_16588,N_10343,N_12262);
nor U16589 (N_16589,N_14194,N_14895);
or U16590 (N_16590,N_10428,N_13379);
nand U16591 (N_16591,N_14095,N_11540);
nand U16592 (N_16592,N_12926,N_14264);
nor U16593 (N_16593,N_14560,N_14628);
nor U16594 (N_16594,N_11523,N_12438);
or U16595 (N_16595,N_14903,N_12582);
nor U16596 (N_16596,N_11194,N_12351);
and U16597 (N_16597,N_11721,N_14735);
or U16598 (N_16598,N_13051,N_12691);
nor U16599 (N_16599,N_12399,N_10961);
xor U16600 (N_16600,N_11071,N_13562);
and U16601 (N_16601,N_13501,N_14559);
nand U16602 (N_16602,N_12933,N_14801);
and U16603 (N_16603,N_12675,N_12683);
nor U16604 (N_16604,N_12065,N_13006);
nand U16605 (N_16605,N_13234,N_10191);
nand U16606 (N_16606,N_10681,N_10673);
or U16607 (N_16607,N_12818,N_12296);
nor U16608 (N_16608,N_11883,N_14799);
and U16609 (N_16609,N_13643,N_11214);
or U16610 (N_16610,N_13350,N_12300);
and U16611 (N_16611,N_10353,N_11387);
nand U16612 (N_16612,N_13397,N_10638);
nand U16613 (N_16613,N_13009,N_11516);
and U16614 (N_16614,N_10687,N_11109);
xnor U16615 (N_16615,N_14226,N_12030);
nand U16616 (N_16616,N_14169,N_12086);
nand U16617 (N_16617,N_11153,N_13638);
nand U16618 (N_16618,N_11100,N_10266);
nand U16619 (N_16619,N_10078,N_10173);
nor U16620 (N_16620,N_13138,N_13629);
or U16621 (N_16621,N_11062,N_14945);
nor U16622 (N_16622,N_14851,N_13149);
nand U16623 (N_16623,N_11229,N_14024);
nor U16624 (N_16624,N_11575,N_12527);
xor U16625 (N_16625,N_12290,N_14620);
nor U16626 (N_16626,N_13448,N_14708);
or U16627 (N_16627,N_12917,N_12126);
and U16628 (N_16628,N_13634,N_12896);
or U16629 (N_16629,N_14475,N_11568);
nand U16630 (N_16630,N_10210,N_11470);
nand U16631 (N_16631,N_12131,N_11492);
xnor U16632 (N_16632,N_10022,N_12457);
nand U16633 (N_16633,N_10314,N_11849);
nor U16634 (N_16634,N_10281,N_13761);
and U16635 (N_16635,N_14522,N_14113);
and U16636 (N_16636,N_12516,N_14567);
nor U16637 (N_16637,N_11291,N_11402);
or U16638 (N_16638,N_13620,N_11559);
and U16639 (N_16639,N_13170,N_14349);
or U16640 (N_16640,N_14409,N_10925);
or U16641 (N_16641,N_12266,N_13556);
xnor U16642 (N_16642,N_10521,N_10633);
nand U16643 (N_16643,N_10480,N_13280);
or U16644 (N_16644,N_11714,N_12154);
or U16645 (N_16645,N_11233,N_14478);
xor U16646 (N_16646,N_11462,N_13896);
nor U16647 (N_16647,N_12120,N_12783);
nand U16648 (N_16648,N_10562,N_14706);
nand U16649 (N_16649,N_12686,N_11264);
or U16650 (N_16650,N_11106,N_14374);
nor U16651 (N_16651,N_14167,N_11148);
nand U16652 (N_16652,N_10091,N_13959);
or U16653 (N_16653,N_10996,N_14353);
or U16654 (N_16654,N_13672,N_10083);
xnor U16655 (N_16655,N_12208,N_10534);
or U16656 (N_16656,N_13939,N_13927);
nand U16657 (N_16657,N_11642,N_13308);
nand U16658 (N_16658,N_12204,N_11333);
nor U16659 (N_16659,N_12123,N_14005);
nand U16660 (N_16660,N_14659,N_10893);
nand U16661 (N_16661,N_11251,N_11493);
or U16662 (N_16662,N_12386,N_12346);
nor U16663 (N_16663,N_10516,N_13468);
nor U16664 (N_16664,N_11351,N_12823);
and U16665 (N_16665,N_10908,N_10113);
or U16666 (N_16666,N_13710,N_10648);
nor U16667 (N_16667,N_10460,N_12634);
or U16668 (N_16668,N_14667,N_14425);
nor U16669 (N_16669,N_11243,N_10646);
and U16670 (N_16670,N_14547,N_10131);
nand U16671 (N_16671,N_14971,N_12337);
xor U16672 (N_16672,N_13865,N_10014);
nand U16673 (N_16673,N_13452,N_10696);
nand U16674 (N_16674,N_11016,N_13140);
nor U16675 (N_16675,N_10423,N_10528);
nand U16676 (N_16676,N_12084,N_10244);
nor U16677 (N_16677,N_12658,N_13682);
nor U16678 (N_16678,N_13921,N_11500);
nor U16679 (N_16679,N_14137,N_10251);
nor U16680 (N_16680,N_11597,N_11357);
or U16681 (N_16681,N_11218,N_10505);
xor U16682 (N_16682,N_14178,N_13757);
nor U16683 (N_16683,N_13916,N_11204);
and U16684 (N_16684,N_13092,N_13886);
nor U16685 (N_16685,N_11664,N_10230);
and U16686 (N_16686,N_13303,N_14622);
nand U16687 (N_16687,N_14411,N_13247);
xor U16688 (N_16688,N_12957,N_13196);
nor U16689 (N_16689,N_13957,N_14675);
nand U16690 (N_16690,N_12842,N_13526);
or U16691 (N_16691,N_12644,N_13476);
or U16692 (N_16692,N_12179,N_13697);
xor U16693 (N_16693,N_12153,N_12685);
nand U16694 (N_16694,N_13762,N_14068);
or U16695 (N_16695,N_12856,N_11515);
and U16696 (N_16696,N_13028,N_11618);
or U16697 (N_16697,N_14663,N_13377);
nand U16698 (N_16698,N_10823,N_10629);
and U16699 (N_16699,N_12482,N_10551);
or U16700 (N_16700,N_12143,N_13135);
nand U16701 (N_16701,N_10066,N_14511);
nand U16702 (N_16702,N_14293,N_13847);
nand U16703 (N_16703,N_11228,N_14807);
nand U16704 (N_16704,N_11423,N_11739);
and U16705 (N_16705,N_14931,N_11480);
xnor U16706 (N_16706,N_13221,N_10401);
xnor U16707 (N_16707,N_10192,N_10634);
or U16708 (N_16708,N_12197,N_14887);
nand U16709 (N_16709,N_12085,N_13993);
nor U16710 (N_16710,N_11297,N_14973);
xnor U16711 (N_16711,N_12105,N_11981);
or U16712 (N_16712,N_11888,N_10820);
or U16713 (N_16713,N_13053,N_13619);
and U16714 (N_16714,N_14453,N_14069);
nand U16715 (N_16715,N_11105,N_12169);
nand U16716 (N_16716,N_10864,N_14919);
nand U16717 (N_16717,N_13365,N_13529);
and U16718 (N_16718,N_11903,N_13679);
nor U16719 (N_16719,N_13950,N_11860);
or U16720 (N_16720,N_13860,N_14035);
nor U16721 (N_16721,N_13208,N_12402);
or U16722 (N_16722,N_11155,N_13418);
and U16723 (N_16723,N_11344,N_12198);
nor U16724 (N_16724,N_12374,N_14176);
or U16725 (N_16725,N_11653,N_14301);
xnor U16726 (N_16726,N_12434,N_14384);
or U16727 (N_16727,N_14520,N_12027);
and U16728 (N_16728,N_10250,N_11494);
nor U16729 (N_16729,N_14382,N_13747);
or U16730 (N_16730,N_11909,N_11055);
and U16731 (N_16731,N_10872,N_12284);
and U16732 (N_16732,N_14009,N_10853);
nor U16733 (N_16733,N_11215,N_12070);
nor U16734 (N_16734,N_12479,N_10178);
and U16735 (N_16735,N_11726,N_14688);
or U16736 (N_16736,N_11073,N_14611);
nand U16737 (N_16737,N_12723,N_14139);
nand U16738 (N_16738,N_10088,N_11150);
or U16739 (N_16739,N_14651,N_11944);
or U16740 (N_16740,N_10784,N_10742);
nand U16741 (N_16741,N_10128,N_10117);
nand U16742 (N_16742,N_11567,N_13793);
or U16743 (N_16743,N_10139,N_13968);
xnor U16744 (N_16744,N_13311,N_14699);
and U16745 (N_16745,N_10465,N_12170);
or U16746 (N_16746,N_12444,N_10682);
and U16747 (N_16747,N_14036,N_14784);
and U16748 (N_16748,N_10054,N_14234);
nand U16749 (N_16749,N_11928,N_12940);
nor U16750 (N_16750,N_11164,N_12183);
or U16751 (N_16751,N_12378,N_14097);
nor U16752 (N_16752,N_12748,N_10826);
nand U16753 (N_16753,N_11476,N_14336);
nand U16754 (N_16754,N_12546,N_11814);
or U16755 (N_16755,N_11803,N_12914);
nor U16756 (N_16756,N_11560,N_11159);
or U16757 (N_16757,N_11330,N_10632);
xnor U16758 (N_16758,N_11921,N_13456);
or U16759 (N_16759,N_10262,N_10018);
nand U16760 (N_16760,N_13644,N_11818);
and U16761 (N_16761,N_14056,N_11142);
and U16762 (N_16762,N_10237,N_14932);
nor U16763 (N_16763,N_11657,N_12472);
xor U16764 (N_16764,N_12798,N_12536);
nand U16765 (N_16765,N_13733,N_13275);
nor U16766 (N_16766,N_14906,N_12422);
and U16767 (N_16767,N_14771,N_12750);
nand U16768 (N_16768,N_11095,N_11372);
and U16769 (N_16769,N_10840,N_13963);
nor U16770 (N_16770,N_12699,N_14051);
and U16771 (N_16771,N_10092,N_10885);
or U16772 (N_16772,N_14011,N_10279);
or U16773 (N_16773,N_13600,N_13803);
and U16774 (N_16774,N_11685,N_11595);
or U16775 (N_16775,N_10604,N_12310);
or U16776 (N_16776,N_13804,N_13511);
and U16777 (N_16777,N_10441,N_13192);
nor U16778 (N_16778,N_11474,N_14539);
or U16779 (N_16779,N_10783,N_10949);
nand U16780 (N_16780,N_12730,N_10759);
xnor U16781 (N_16781,N_11998,N_12515);
or U16782 (N_16782,N_12803,N_13917);
nor U16783 (N_16783,N_13047,N_11552);
and U16784 (N_16784,N_10267,N_13298);
and U16785 (N_16785,N_12226,N_14950);
or U16786 (N_16786,N_13966,N_12115);
and U16787 (N_16787,N_11273,N_10212);
or U16788 (N_16788,N_11773,N_14994);
nand U16789 (N_16789,N_14889,N_10112);
or U16790 (N_16790,N_11935,N_10965);
or U16791 (N_16791,N_13241,N_10154);
xor U16792 (N_16792,N_11997,N_13395);
or U16793 (N_16793,N_14089,N_12270);
nand U16794 (N_16794,N_11341,N_13130);
and U16795 (N_16795,N_10001,N_12055);
xnor U16796 (N_16796,N_13117,N_11363);
or U16797 (N_16797,N_13370,N_14432);
or U16798 (N_16798,N_13835,N_12232);
or U16799 (N_16799,N_12267,N_12793);
nor U16800 (N_16800,N_13482,N_13252);
nand U16801 (N_16801,N_14151,N_10582);
nor U16802 (N_16802,N_10986,N_13813);
and U16803 (N_16803,N_14189,N_10903);
and U16804 (N_16804,N_13498,N_10086);
nand U16805 (N_16805,N_10654,N_12275);
or U16806 (N_16806,N_10554,N_13971);
and U16807 (N_16807,N_13271,N_13544);
xnor U16808 (N_16808,N_10860,N_12631);
or U16809 (N_16809,N_12273,N_11930);
nand U16810 (N_16810,N_10055,N_14369);
xor U16811 (N_16811,N_11669,N_11565);
nor U16812 (N_16812,N_14070,N_14552);
nand U16813 (N_16813,N_10164,N_11551);
nand U16814 (N_16814,N_10995,N_10587);
and U16815 (N_16815,N_13903,N_12016);
nand U16816 (N_16816,N_14480,N_14158);
or U16817 (N_16817,N_11931,N_14561);
xor U16818 (N_16818,N_12981,N_12825);
nand U16819 (N_16819,N_10600,N_10187);
or U16820 (N_16820,N_13284,N_14681);
nand U16821 (N_16821,N_13660,N_10177);
or U16822 (N_16822,N_10466,N_11799);
or U16823 (N_16823,N_14098,N_14307);
or U16824 (N_16824,N_13670,N_11112);
nor U16825 (N_16825,N_13692,N_13174);
nor U16826 (N_16826,N_13202,N_10469);
nand U16827 (N_16827,N_11391,N_11162);
nand U16828 (N_16828,N_11007,N_12764);
or U16829 (N_16829,N_13923,N_11518);
nor U16830 (N_16830,N_14501,N_10087);
nand U16831 (N_16831,N_12168,N_14550);
xnor U16832 (N_16832,N_13738,N_12755);
and U16833 (N_16833,N_12701,N_11369);
nor U16834 (N_16834,N_14549,N_14519);
or U16835 (N_16835,N_14088,N_11449);
nor U16836 (N_16836,N_14958,N_12771);
nand U16837 (N_16837,N_11892,N_13758);
and U16838 (N_16838,N_11972,N_14703);
or U16839 (N_16839,N_12286,N_11129);
nand U16840 (N_16840,N_10560,N_11157);
nor U16841 (N_16841,N_10806,N_11415);
nor U16842 (N_16842,N_11734,N_10095);
or U16843 (N_16843,N_12891,N_14085);
nor U16844 (N_16844,N_11083,N_12282);
or U16845 (N_16845,N_14935,N_13176);
nand U16846 (N_16846,N_12603,N_13437);
or U16847 (N_16847,N_13254,N_14358);
nor U16848 (N_16848,N_10327,N_11025);
or U16849 (N_16849,N_12739,N_10517);
nand U16850 (N_16850,N_14721,N_14562);
nand U16851 (N_16851,N_11816,N_10833);
nor U16852 (N_16852,N_11947,N_13188);
nand U16853 (N_16853,N_13947,N_10941);
nor U16854 (N_16854,N_13989,N_12165);
nor U16855 (N_16855,N_12985,N_10490);
nor U16856 (N_16856,N_12919,N_14728);
or U16857 (N_16857,N_10909,N_12804);
and U16858 (N_16858,N_12231,N_14666);
nand U16859 (N_16859,N_10832,N_13157);
or U16860 (N_16860,N_13879,N_10578);
xnor U16861 (N_16861,N_12866,N_10081);
nand U16862 (N_16862,N_13326,N_11843);
nor U16863 (N_16863,N_12233,N_14883);
or U16864 (N_16864,N_14090,N_14954);
nand U16865 (N_16865,N_13011,N_13741);
nand U16866 (N_16866,N_11623,N_12408);
or U16867 (N_16867,N_11125,N_11422);
or U16868 (N_16868,N_11275,N_10989);
nor U16869 (N_16869,N_12619,N_13477);
nand U16870 (N_16870,N_10330,N_10287);
and U16871 (N_16871,N_10454,N_10743);
and U16872 (N_16872,N_10500,N_10891);
and U16873 (N_16873,N_11487,N_10341);
nand U16874 (N_16874,N_13375,N_11580);
and U16875 (N_16875,N_12700,N_14454);
and U16876 (N_16876,N_13859,N_14979);
or U16877 (N_16877,N_12706,N_12860);
or U16878 (N_16878,N_14393,N_10031);
nand U16879 (N_16879,N_12117,N_14484);
or U16880 (N_16880,N_11417,N_14120);
and U16881 (N_16881,N_10731,N_12046);
xnor U16882 (N_16882,N_11707,N_11652);
nand U16883 (N_16883,N_12632,N_13755);
xor U16884 (N_16884,N_14223,N_14156);
or U16885 (N_16885,N_10935,N_14302);
and U16886 (N_16886,N_13955,N_11137);
nor U16887 (N_16887,N_14495,N_13882);
nor U16888 (N_16888,N_10589,N_14597);
nand U16889 (N_16889,N_11821,N_10228);
nor U16890 (N_16890,N_13914,N_13736);
and U16891 (N_16891,N_13823,N_13805);
nor U16892 (N_16892,N_13245,N_11147);
and U16893 (N_16893,N_10042,N_10615);
nand U16894 (N_16894,N_13689,N_12968);
nand U16895 (N_16895,N_13946,N_14876);
or U16896 (N_16896,N_11993,N_14563);
and U16897 (N_16897,N_14481,N_10484);
nor U16898 (N_16898,N_12819,N_13852);
xor U16899 (N_16899,N_11755,N_10174);
xor U16900 (N_16900,N_12749,N_12709);
nand U16901 (N_16901,N_11355,N_13680);
nor U16902 (N_16902,N_13840,N_12175);
or U16903 (N_16903,N_12015,N_13333);
and U16904 (N_16904,N_11889,N_13866);
nor U16905 (N_16905,N_11478,N_11024);
nor U16906 (N_16906,N_13952,N_12369);
xor U16907 (N_16907,N_10899,N_10529);
xnor U16908 (N_16908,N_14012,N_11675);
or U16909 (N_16909,N_14690,N_12676);
or U16910 (N_16910,N_10026,N_12581);
and U16911 (N_16911,N_10477,N_13203);
or U16912 (N_16912,N_13067,N_11769);
nand U16913 (N_16913,N_14253,N_11305);
and U16914 (N_16914,N_12218,N_11761);
nor U16915 (N_16915,N_13032,N_12892);
nor U16916 (N_16916,N_11485,N_11901);
nor U16917 (N_16917,N_11677,N_12205);
and U16918 (N_16918,N_11839,N_12149);
and U16919 (N_16919,N_14525,N_14686);
or U16920 (N_16920,N_13089,N_14995);
or U16921 (N_16921,N_13977,N_10939);
and U16922 (N_16922,N_12432,N_10045);
nor U16923 (N_16923,N_12629,N_14485);
or U16924 (N_16924,N_14654,N_11212);
xnor U16925 (N_16925,N_13257,N_12872);
nor U16926 (N_16926,N_10959,N_14465);
xor U16927 (N_16927,N_13612,N_13038);
xor U16928 (N_16928,N_13746,N_10216);
nand U16929 (N_16929,N_11061,N_14319);
nor U16930 (N_16930,N_10003,N_13877);
nand U16931 (N_16931,N_14756,N_10393);
nor U16932 (N_16932,N_14866,N_11542);
or U16933 (N_16933,N_12335,N_12622);
or U16934 (N_16934,N_13359,N_12743);
or U16935 (N_16935,N_12217,N_12312);
or U16936 (N_16936,N_13777,N_14456);
nand U16937 (N_16937,N_10149,N_10755);
and U16938 (N_16938,N_11202,N_10046);
and U16939 (N_16939,N_14351,N_10218);
nor U16940 (N_16940,N_12520,N_11593);
nor U16941 (N_16941,N_14261,N_13724);
nor U16942 (N_16942,N_11356,N_10627);
nand U16943 (N_16943,N_13079,N_14229);
and U16944 (N_16944,N_14414,N_13118);
nor U16945 (N_16945,N_10776,N_13387);
xor U16946 (N_16946,N_11086,N_11197);
and U16947 (N_16947,N_14060,N_14516);
or U16948 (N_16948,N_13127,N_10381);
and U16949 (N_16949,N_12060,N_13748);
or U16950 (N_16950,N_12321,N_12663);
nand U16951 (N_16951,N_11370,N_13103);
nand U16952 (N_16952,N_12002,N_12017);
or U16953 (N_16953,N_14163,N_11213);
and U16954 (N_16954,N_11996,N_10874);
nor U16955 (N_16955,N_10144,N_13273);
or U16956 (N_16956,N_12162,N_12393);
nor U16957 (N_16957,N_13770,N_11867);
and U16958 (N_16958,N_10724,N_14853);
or U16959 (N_16959,N_14879,N_13412);
nand U16960 (N_16960,N_13842,N_12324);
nor U16961 (N_16961,N_11135,N_14285);
nor U16962 (N_16962,N_11973,N_10057);
nand U16963 (N_16963,N_13525,N_11757);
xor U16964 (N_16964,N_10608,N_12459);
or U16965 (N_16965,N_11443,N_13416);
and U16966 (N_16966,N_14623,N_11713);
nor U16967 (N_16967,N_10769,N_11467);
and U16968 (N_16968,N_14993,N_10892);
or U16969 (N_16969,N_12305,N_11553);
and U16970 (N_16970,N_12327,N_13681);
nor U16971 (N_16971,N_10030,N_10137);
nor U16972 (N_16972,N_11405,N_13518);
or U16973 (N_16973,N_14503,N_10337);
and U16974 (N_16974,N_11245,N_13936);
nor U16975 (N_16975,N_10365,N_13920);
nor U16976 (N_16976,N_11165,N_13403);
or U16977 (N_16977,N_11346,N_12562);
nand U16978 (N_16978,N_13293,N_10037);
and U16979 (N_16979,N_10752,N_11539);
or U16980 (N_16980,N_10652,N_13388);
nor U16981 (N_16981,N_11292,N_14104);
nand U16982 (N_16982,N_14910,N_11608);
xnor U16983 (N_16983,N_14817,N_11267);
nand U16984 (N_16984,N_12888,N_10927);
xnor U16985 (N_16985,N_11249,N_11394);
xor U16986 (N_16986,N_13484,N_10815);
and U16987 (N_16987,N_14683,N_11237);
nand U16988 (N_16988,N_13904,N_12806);
and U16989 (N_16989,N_11858,N_10008);
or U16990 (N_16990,N_12796,N_11296);
nand U16991 (N_16991,N_10356,N_10052);
and U16992 (N_16992,N_10675,N_13483);
nor U16993 (N_16993,N_11004,N_11272);
or U16994 (N_16994,N_14217,N_10059);
nand U16995 (N_16995,N_14213,N_14508);
and U16996 (N_16996,N_13367,N_11224);
and U16997 (N_16997,N_10569,N_12364);
or U16998 (N_16998,N_13021,N_14497);
or U16999 (N_16999,N_13967,N_11706);
nand U17000 (N_17000,N_14859,N_12609);
xnor U17001 (N_17001,N_13707,N_11876);
nor U17002 (N_17002,N_13285,N_13155);
xnor U17003 (N_17003,N_13123,N_12550);
nor U17004 (N_17004,N_10097,N_12510);
nand U17005 (N_17005,N_13668,N_12827);
and U17006 (N_17006,N_14584,N_11190);
and U17007 (N_17007,N_12083,N_10122);
nor U17008 (N_17008,N_11829,N_13313);
and U17009 (N_17009,N_10103,N_13471);
and U17010 (N_17010,N_11882,N_11771);
nand U17011 (N_17011,N_14977,N_12251);
nor U17012 (N_17012,N_11285,N_13737);
and U17013 (N_17013,N_10405,N_13018);
nor U17014 (N_17014,N_14826,N_10510);
and U17015 (N_17015,N_12817,N_14419);
or U17016 (N_17016,N_13824,N_13005);
or U17017 (N_17017,N_11994,N_13960);
and U17018 (N_17018,N_13425,N_11364);
or U17019 (N_17019,N_13357,N_11426);
xor U17020 (N_17020,N_14884,N_11036);
and U17021 (N_17021,N_11358,N_10169);
nor U17022 (N_17022,N_13249,N_12977);
or U17023 (N_17023,N_13706,N_11293);
or U17024 (N_17024,N_13146,N_10429);
nor U17025 (N_17025,N_12302,N_12588);
xor U17026 (N_17026,N_14428,N_12189);
and U17027 (N_17027,N_12349,N_11498);
nor U17028 (N_17028,N_10915,N_13381);
nor U17029 (N_17029,N_10786,N_12778);
xnor U17030 (N_17030,N_11507,N_14433);
nor U17031 (N_17031,N_11248,N_13538);
nand U17032 (N_17032,N_14814,N_14860);
or U17033 (N_17033,N_12424,N_13189);
nor U17034 (N_17034,N_13565,N_10447);
and U17035 (N_17035,N_11287,N_13270);
nand U17036 (N_17036,N_11964,N_12735);
xor U17037 (N_17037,N_14837,N_10992);
nand U17038 (N_17038,N_10526,N_14410);
xnor U17039 (N_17039,N_11481,N_11751);
and U17040 (N_17040,N_14443,N_12258);
nor U17041 (N_17041,N_10146,N_13494);
xor U17042 (N_17042,N_12109,N_12147);
or U17043 (N_17043,N_14418,N_13913);
nor U17044 (N_17044,N_12626,N_10268);
nand U17045 (N_17045,N_11853,N_12237);
nor U17046 (N_17046,N_13640,N_13074);
or U17047 (N_17047,N_10593,N_12426);
or U17048 (N_17048,N_12508,N_12470);
xnor U17049 (N_17049,N_14292,N_11046);
or U17050 (N_17050,N_12967,N_10274);
xor U17051 (N_17051,N_13652,N_11927);
or U17052 (N_17052,N_14797,N_10779);
nor U17053 (N_17053,N_13837,N_10650);
or U17054 (N_17054,N_12163,N_14648);
xnor U17055 (N_17055,N_13366,N_10079);
nor U17056 (N_17056,N_14072,N_14668);
or U17057 (N_17057,N_13120,N_11881);
or U17058 (N_17058,N_10025,N_10050);
nor U17059 (N_17059,N_10424,N_14370);
and U17060 (N_17060,N_13124,N_11779);
xnor U17061 (N_17061,N_11438,N_11029);
or U17062 (N_17062,N_12485,N_14922);
nor U17063 (N_17063,N_12874,N_13774);
nor U17064 (N_17064,N_14018,N_13321);
nand U17065 (N_17065,N_11875,N_12291);
nor U17066 (N_17066,N_10501,N_10933);
xor U17067 (N_17067,N_13261,N_13628);
xor U17068 (N_17068,N_14265,N_10161);
nand U17069 (N_17069,N_13752,N_14718);
nand U17070 (N_17070,N_10777,N_14315);
or U17071 (N_17071,N_10229,N_11070);
xnor U17072 (N_17072,N_13915,N_14227);
or U17073 (N_17073,N_14632,N_12250);
nor U17074 (N_17074,N_10311,N_13352);
nand U17075 (N_17075,N_13584,N_11424);
or U17076 (N_17076,N_13217,N_13376);
and U17077 (N_17077,N_11869,N_11324);
xnor U17078 (N_17078,N_14865,N_13260);
nor U17079 (N_17079,N_14247,N_14750);
xor U17080 (N_17080,N_10553,N_13531);
nand U17081 (N_17081,N_13133,N_14960);
nand U17082 (N_17082,N_11139,N_10905);
nand U17083 (N_17083,N_11919,N_14239);
nor U17084 (N_17084,N_13136,N_10748);
and U17085 (N_17085,N_13695,N_14780);
nor U17086 (N_17086,N_11128,N_10775);
nand U17087 (N_17087,N_13723,N_14742);
nor U17088 (N_17088,N_12156,N_12475);
or U17089 (N_17089,N_14093,N_11087);
nand U17090 (N_17090,N_14040,N_12061);
or U17091 (N_17091,N_14978,N_12924);
nand U17092 (N_17092,N_13809,N_10543);
or U17093 (N_17093,N_12078,N_14855);
or U17094 (N_17094,N_14306,N_13364);
or U17095 (N_17095,N_13453,N_11318);
or U17096 (N_17096,N_12942,N_10954);
nor U17097 (N_17097,N_12397,N_11065);
nand U17098 (N_17098,N_11043,N_10753);
nor U17099 (N_17099,N_11836,N_10358);
or U17100 (N_17100,N_10422,N_12653);
nand U17101 (N_17101,N_11733,N_12079);
or U17102 (N_17102,N_12811,N_11081);
or U17103 (N_17103,N_12054,N_11266);
nand U17104 (N_17104,N_11263,N_14505);
nand U17105 (N_17105,N_10090,N_11660);
nor U17106 (N_17106,N_14231,N_10333);
or U17107 (N_17107,N_12782,N_14926);
or U17108 (N_17108,N_12927,N_10549);
nor U17109 (N_17109,N_14327,N_13632);
and U17110 (N_17110,N_11097,N_14262);
or U17111 (N_17111,N_14755,N_13279);
and U17112 (N_17112,N_11460,N_12326);
nand U17113 (N_17113,N_14864,N_11126);
or U17114 (N_17114,N_11610,N_11656);
and U17115 (N_17115,N_12329,N_10876);
nor U17116 (N_17116,N_11975,N_10788);
and U17117 (N_17117,N_10668,N_14658);
nand U17118 (N_17118,N_13024,N_12040);
and U17119 (N_17119,N_10819,N_11850);
nor U17120 (N_17120,N_13656,N_11182);
or U17121 (N_17121,N_13025,N_11703);
or U17122 (N_17122,N_10993,N_13336);
nand U17123 (N_17123,N_11647,N_13175);
and U17124 (N_17124,N_10468,N_11027);
nand U17125 (N_17125,N_11390,N_10886);
nand U17126 (N_17126,N_11957,N_12122);
xor U17127 (N_17127,N_13834,N_13816);
nor U17128 (N_17128,N_12518,N_10431);
or U17129 (N_17129,N_13580,N_12368);
nand U17130 (N_17130,N_11920,N_11765);
and U17131 (N_17131,N_11918,N_12785);
xnor U17132 (N_17132,N_10012,N_10179);
or U17133 (N_17133,N_13031,N_13661);
nor U17134 (N_17134,N_11479,N_10292);
nor U17135 (N_17135,N_12441,N_13742);
and U17136 (N_17136,N_14614,N_10895);
or U17137 (N_17137,N_14303,N_13677);
and U17138 (N_17138,N_11884,N_10835);
nand U17139 (N_17139,N_11209,N_14420);
nand U17140 (N_17140,N_10997,N_11530);
or U17141 (N_17141,N_12960,N_12446);
nand U17142 (N_17142,N_13147,N_11789);
and U17143 (N_17143,N_10732,N_14857);
nand U17144 (N_17144,N_12604,N_12026);
or U17145 (N_17145,N_12740,N_11114);
and U17146 (N_17146,N_13618,N_10811);
nand U17147 (N_17147,N_13537,N_13324);
nor U17148 (N_17148,N_11506,N_14710);
nand U17149 (N_17149,N_12849,N_11630);
or U17150 (N_17150,N_13832,N_14557);
nor U17151 (N_17151,N_10494,N_14753);
and U17152 (N_17152,N_13509,N_10159);
or U17153 (N_17153,N_11326,N_13044);
or U17154 (N_17154,N_13597,N_10035);
nor U17155 (N_17155,N_10440,N_11689);
or U17156 (N_17156,N_13614,N_12884);
nor U17157 (N_17157,N_12288,N_10080);
or U17158 (N_17158,N_13166,N_10680);
nand U17159 (N_17159,N_10818,N_12128);
and U17160 (N_17160,N_14996,N_14943);
nor U17161 (N_17161,N_13602,N_12930);
or U17162 (N_17162,N_13540,N_11556);
nor U17163 (N_17163,N_14692,N_14482);
xor U17164 (N_17164,N_14953,N_12129);
nor U17165 (N_17165,N_13591,N_13310);
nor U17166 (N_17166,N_14898,N_10197);
nand U17167 (N_17167,N_10644,N_11337);
xnor U17168 (N_17168,N_12311,N_13996);
nand U17169 (N_17169,N_14283,N_13653);
and U17170 (N_17170,N_12328,N_13790);
and U17171 (N_17171,N_14916,N_12483);
nand U17172 (N_17172,N_13269,N_11289);
nand U17173 (N_17173,N_14053,N_10374);
and U17174 (N_17174,N_12243,N_11719);
or U17175 (N_17175,N_12067,N_10436);
nor U17176 (N_17176,N_14610,N_14138);
or U17177 (N_17177,N_12395,N_10403);
nor U17178 (N_17178,N_10181,N_14693);
or U17179 (N_17179,N_11231,N_12097);
or U17180 (N_17180,N_12436,N_13609);
nand U17181 (N_17181,N_10975,N_13394);
and U17182 (N_17182,N_12671,N_11084);
or U17183 (N_17183,N_10541,N_12222);
or U17184 (N_17184,N_10024,N_12826);
and U17185 (N_17185,N_12194,N_11795);
or U17186 (N_17186,N_13648,N_11785);
and U17187 (N_17187,N_14757,N_12779);
nand U17188 (N_17188,N_10917,N_13557);
nor U17189 (N_17189,N_12454,N_12614);
or U17190 (N_17190,N_11582,N_14959);
and U17191 (N_17191,N_13814,N_13726);
nor U17192 (N_17192,N_10968,N_13559);
and U17193 (N_17193,N_14118,N_13191);
nor U17194 (N_17194,N_11187,N_12468);
nor U17195 (N_17195,N_13975,N_12044);
or U17196 (N_17196,N_14084,N_14800);
nand U17197 (N_17197,N_12570,N_11077);
and U17198 (N_17198,N_14033,N_14843);
and U17199 (N_17199,N_12953,N_13274);
or U17200 (N_17200,N_10058,N_12729);
or U17201 (N_17201,N_11929,N_14548);
nand U17202 (N_17202,N_13301,N_10705);
nor U17203 (N_17203,N_11466,N_10834);
or U17204 (N_17204,N_14743,N_14422);
nand U17205 (N_17205,N_10143,N_12341);
or U17206 (N_17206,N_10145,N_11543);
and U17207 (N_17207,N_11178,N_12157);
nor U17208 (N_17208,N_13796,N_14235);
nor U17209 (N_17209,N_10489,N_13296);
nand U17210 (N_17210,N_11809,N_10506);
nand U17211 (N_17211,N_13862,N_11483);
or U17212 (N_17212,N_10780,N_14643);
or U17213 (N_17213,N_14773,N_12392);
and U17214 (N_17214,N_12072,N_10116);
nor U17215 (N_17215,N_14787,N_12298);
nand U17216 (N_17216,N_12994,N_14720);
and U17217 (N_17217,N_13786,N_11127);
nand U17218 (N_17218,N_11039,N_10339);
nor U17219 (N_17219,N_12132,N_12278);
and U17220 (N_17220,N_12726,N_10620);
nor U17221 (N_17221,N_11536,N_10384);
or U17222 (N_17222,N_12474,N_10020);
and U17223 (N_17223,N_10653,N_11636);
nand U17224 (N_17224,N_13657,N_10382);
or U17225 (N_17225,N_12938,N_14266);
xnor U17226 (N_17226,N_13709,N_12469);
nand U17227 (N_17227,N_11037,N_14002);
nor U17228 (N_17228,N_14871,N_10019);
xor U17229 (N_17229,N_11170,N_12955);
and U17230 (N_17230,N_13844,N_13256);
nand U17231 (N_17231,N_12445,N_14186);
nor U17232 (N_17232,N_14909,N_14233);
nor U17233 (N_17233,N_12260,N_11764);
nor U17234 (N_17234,N_13063,N_13554);
and U17235 (N_17235,N_12007,N_12753);
or U17236 (N_17236,N_10873,N_12937);
and U17237 (N_17237,N_10435,N_12376);
or U17238 (N_17238,N_13926,N_10866);
and U17239 (N_17239,N_14210,N_11968);
nand U17240 (N_17240,N_10016,N_10814);
nor U17241 (N_17241,N_10546,N_10310);
nor U17242 (N_17242,N_14587,N_10168);
nor U17243 (N_17243,N_10172,N_12382);
xor U17244 (N_17244,N_13297,N_12661);
and U17245 (N_17245,N_10847,N_14000);
or U17246 (N_17246,N_14025,N_11072);
nor U17247 (N_17247,N_10556,N_13110);
and U17248 (N_17248,N_13351,N_11301);
or U17249 (N_17249,N_11628,N_11210);
nor U17250 (N_17250,N_12148,N_10745);
or U17251 (N_17251,N_14783,N_13940);
xnor U17252 (N_17252,N_14694,N_11006);
and U17253 (N_17253,N_13719,N_11545);
or U17254 (N_17254,N_14774,N_10132);
and U17255 (N_17255,N_13523,N_12539);
or U17256 (N_17256,N_14295,N_12979);
xnor U17257 (N_17257,N_11564,N_10952);
nor U17258 (N_17258,N_14168,N_10781);
or U17259 (N_17259,N_12220,N_10155);
and U17260 (N_17260,N_13331,N_10987);
nor U17261 (N_17261,N_14479,N_13438);
nor U17262 (N_17262,N_12997,N_10707);
xor U17263 (N_17263,N_14809,N_13508);
nand U17264 (N_17264,N_13015,N_12037);
nand U17265 (N_17265,N_14030,N_12746);
or U17266 (N_17266,N_12405,N_10085);
nand U17267 (N_17267,N_12453,N_14106);
or U17268 (N_17268,N_10994,N_13784);
nor U17269 (N_17269,N_14802,N_14006);
nand U17270 (N_17270,N_12215,N_14441);
and U17271 (N_17271,N_10067,N_14451);
or U17272 (N_17272,N_12010,N_10645);
nand U17273 (N_17273,N_14054,N_12522);
or U17274 (N_17274,N_14459,N_11579);
and U17275 (N_17275,N_10701,N_14537);
nand U17276 (N_17276,N_12028,N_13642);
nor U17277 (N_17277,N_11367,N_12794);
and U17278 (N_17278,N_13169,N_14948);
and U17279 (N_17279,N_14125,N_13093);
or U17280 (N_17280,N_11132,N_14362);
and U17281 (N_17281,N_14080,N_14849);
nor U17282 (N_17282,N_14553,N_13716);
or U17283 (N_17283,N_14215,N_11945);
nand U17284 (N_17284,N_12712,N_12287);
and U17285 (N_17285,N_10299,N_11434);
and U17286 (N_17286,N_10900,N_13873);
nand U17287 (N_17287,N_14032,N_11900);
nor U17288 (N_17288,N_13487,N_13945);
or U17289 (N_17289,N_11787,N_12784);
nand U17290 (N_17290,N_10407,N_14344);
nor U17291 (N_17291,N_14219,N_13573);
xnor U17292 (N_17292,N_12531,N_14820);
nand U17293 (N_17293,N_12387,N_12902);
and U17294 (N_17294,N_14847,N_13646);
nand U17295 (N_17295,N_11980,N_10280);
xnor U17296 (N_17296,N_13463,N_11486);
nor U17297 (N_17297,N_11951,N_12714);
nor U17298 (N_17298,N_10452,N_14709);
nand U17299 (N_17299,N_14195,N_14831);
and U17300 (N_17300,N_10175,N_10254);
xnor U17301 (N_17301,N_14395,N_14255);
nand U17302 (N_17302,N_12765,N_11519);
nor U17303 (N_17303,N_14145,N_12879);
nor U17304 (N_17304,N_12616,N_14631);
xnor U17305 (N_17305,N_12160,N_13179);
and U17306 (N_17306,N_10278,N_10884);
and U17307 (N_17307,N_10774,N_13345);
and U17308 (N_17308,N_12840,N_12380);
nand U17309 (N_17309,N_14702,N_14471);
or U17310 (N_17310,N_12276,N_10520);
nor U17311 (N_17311,N_12398,N_11131);
nor U17312 (N_17312,N_10605,N_11103);
nand U17313 (N_17313,N_12389,N_14676);
xor U17314 (N_17314,N_14116,N_14161);
or U17315 (N_17315,N_10446,N_12877);
or U17316 (N_17316,N_14662,N_13970);
or U17317 (N_17317,N_11404,N_11397);
and U17318 (N_17318,N_14021,N_14982);
nor U17319 (N_17319,N_12655,N_10880);
and U17320 (N_17320,N_10269,N_11121);
nor U17321 (N_17321,N_12412,N_10767);
nor U17322 (N_17322,N_11599,N_14119);
or U17323 (N_17323,N_12774,N_14938);
nor U17324 (N_17324,N_11510,N_10919);
nand U17325 (N_17325,N_12853,N_14010);
or U17326 (N_17326,N_10453,N_11453);
nor U17327 (N_17327,N_10622,N_14381);
nand U17328 (N_17328,N_12316,N_13592);
nor U17329 (N_17329,N_14134,N_11971);
or U17330 (N_17330,N_14135,N_13715);
nor U17331 (N_17331,N_14316,N_12813);
and U17332 (N_17332,N_13791,N_13263);
nand U17333 (N_17333,N_13016,N_13346);
nand U17334 (N_17334,N_12317,N_13082);
nor U17335 (N_17335,N_12897,N_13447);
nor U17336 (N_17336,N_14515,N_12242);
nand U17337 (N_17337,N_12280,N_12092);
nand U17338 (N_17338,N_10662,N_11376);
or U17339 (N_17339,N_10547,N_14489);
nor U17340 (N_17340,N_12080,N_10235);
nand U17341 (N_17341,N_10584,N_14103);
nand U17342 (N_17342,N_14225,N_12802);
nand U17343 (N_17343,N_14477,N_13464);
and U17344 (N_17344,N_11343,N_12401);
and U17345 (N_17345,N_10208,N_13595);
and U17346 (N_17346,N_10898,N_14868);
xnor U17347 (N_17347,N_13607,N_10631);
nor U17348 (N_17348,N_11089,N_10307);
xnor U17349 (N_17349,N_10640,N_12810);
and U17350 (N_17350,N_11189,N_12019);
nor U17351 (N_17351,N_13745,N_14621);
nand U17352 (N_17352,N_10319,N_14154);
or U17353 (N_17353,N_14509,N_14413);
or U17354 (N_17354,N_13258,N_10375);
nand U17355 (N_17355,N_14535,N_10625);
or U17356 (N_17356,N_11873,N_12638);
nor U17357 (N_17357,N_10514,N_10010);
nor U17358 (N_17358,N_11563,N_13922);
nor U17359 (N_17359,N_13663,N_11852);
nor U17360 (N_17360,N_13734,N_14407);
and U17361 (N_17361,N_14650,N_11448);
nor U17362 (N_17362,N_11117,N_13150);
or U17363 (N_17363,N_10376,N_12836);
or U17364 (N_17364,N_13662,N_14913);
xnor U17365 (N_17365,N_13073,N_12142);
or U17366 (N_17366,N_12907,N_14429);
or U17367 (N_17367,N_14082,N_14074);
and U17368 (N_17368,N_10108,N_11172);
nand U17369 (N_17369,N_10974,N_11175);
xor U17370 (N_17370,N_13895,N_12567);
nor U17371 (N_17371,N_13334,N_11451);
and U17372 (N_17372,N_13122,N_11681);
nor U17373 (N_17373,N_11794,N_14230);
or U17374 (N_17374,N_12322,N_13567);
and U17375 (N_17375,N_13013,N_13210);
or U17376 (N_17376,N_13506,N_11962);
or U17377 (N_17377,N_10072,N_10213);
nand U17378 (N_17378,N_10414,N_13104);
nor U17379 (N_17379,N_10011,N_11111);
nor U17380 (N_17380,N_12240,N_11749);
or U17381 (N_17381,N_13159,N_12244);
nand U17382 (N_17382,N_11940,N_12011);
or U17383 (N_17383,N_12673,N_13581);
or U17384 (N_17384,N_13831,N_14646);
or U17385 (N_17385,N_13622,N_10508);
and U17386 (N_17386,N_13033,N_11687);
nor U17387 (N_17387,N_11807,N_13678);
or U17388 (N_17388,N_12056,N_14881);
or U17389 (N_17389,N_10661,N_14698);
xnor U17390 (N_17390,N_10926,N_10336);
or U17391 (N_17391,N_14524,N_12064);
or U17392 (N_17392,N_10246,N_13080);
nand U17393 (N_17393,N_14131,N_12174);
nand U17394 (N_17394,N_12904,N_10978);
nor U17395 (N_17395,N_12354,N_11473);
nor U17396 (N_17396,N_11622,N_11199);
nand U17397 (N_17397,N_13564,N_13061);
xnor U17398 (N_17398,N_13587,N_11134);
nor U17399 (N_17399,N_14517,N_13869);
nand U17400 (N_17400,N_13596,N_14727);
nor U17401 (N_17401,N_13474,N_10944);
or U17402 (N_17402,N_10782,N_12181);
or U17403 (N_17403,N_11682,N_12865);
nor U17404 (N_17404,N_10476,N_13696);
and U17405 (N_17405,N_12946,N_11547);
nand U17406 (N_17406,N_11922,N_14446);
nand U17407 (N_17407,N_11038,N_12150);
and U17408 (N_17408,N_11254,N_12050);
xor U17409 (N_17409,N_12731,N_11056);
or U17410 (N_17410,N_12073,N_11880);
and U17411 (N_17411,N_14498,N_12135);
and U17412 (N_17412,N_13908,N_13239);
and U17413 (N_17413,N_12362,N_12248);
nand U17414 (N_17414,N_12137,N_11855);
and U17415 (N_17415,N_12384,N_10658);
nor U17416 (N_17416,N_11708,N_11328);
nor U17417 (N_17417,N_11912,N_10306);
nor U17418 (N_17418,N_11590,N_14839);
nor U17419 (N_17419,N_11184,N_12502);
xnor U17420 (N_17420,N_11299,N_14019);
and U17421 (N_17421,N_10119,N_12211);
nand U17422 (N_17422,N_12763,N_10867);
xor U17423 (N_17423,N_11308,N_11241);
nor U17424 (N_17424,N_12428,N_12958);
and U17425 (N_17425,N_14494,N_14603);
and U17426 (N_17426,N_12534,N_14112);
nand U17427 (N_17427,N_12133,N_10053);
and U17428 (N_17428,N_12216,N_12777);
nor U17429 (N_17429,N_13238,N_12697);
or U17430 (N_17430,N_12991,N_14529);
or U17431 (N_17431,N_10602,N_12529);
xnor U17432 (N_17432,N_14166,N_10406);
xor U17433 (N_17433,N_10261,N_12612);
nor U17434 (N_17434,N_12196,N_14042);
or U17435 (N_17435,N_12800,N_12594);
or U17436 (N_17436,N_11110,N_10773);
nand U17437 (N_17437,N_14462,N_13265);
xnor U17438 (N_17438,N_11613,N_10271);
nor U17439 (N_17439,N_12227,N_12042);
nor U17440 (N_17440,N_13077,N_13615);
or U17441 (N_17441,N_11573,N_10334);
nor U17442 (N_17442,N_14963,N_10515);
nand U17443 (N_17443,N_10462,N_13944);
nand U17444 (N_17444,N_12670,N_11368);
nor U17445 (N_17445,N_12400,N_14152);
and U17446 (N_17446,N_10347,N_10699);
nor U17447 (N_17447,N_10243,N_13978);
xnor U17448 (N_17448,N_12637,N_14697);
nor U17449 (N_17449,N_11188,N_10138);
and U17450 (N_17450,N_13390,N_10048);
nor U17451 (N_17451,N_12219,N_12720);
xnor U17452 (N_17452,N_13850,N_11693);
nand U17453 (N_17453,N_11388,N_12366);
nor U17454 (N_17454,N_11667,N_12617);
or U17455 (N_17455,N_14383,N_14450);
and U17456 (N_17456,N_10897,N_10976);
xnor U17457 (N_17457,N_10639,N_10338);
and U17458 (N_17458,N_14339,N_13071);
or U17459 (N_17459,N_12095,N_11729);
nor U17460 (N_17460,N_10991,N_10844);
and U17461 (N_17461,N_14877,N_12303);
and U17462 (N_17462,N_13181,N_11658);
or U17463 (N_17463,N_11491,N_10304);
nor U17464 (N_17464,N_14144,N_10856);
nor U17465 (N_17465,N_11140,N_10739);
xnor U17466 (N_17466,N_11517,N_12268);
nand U17467 (N_17467,N_14237,N_14842);
xor U17468 (N_17468,N_14192,N_11464);
or U17469 (N_17469,N_11895,N_14528);
or U17470 (N_17470,N_14191,N_14246);
and U17471 (N_17471,N_12456,N_12682);
nand U17472 (N_17472,N_11746,N_11094);
nor U17473 (N_17473,N_10272,N_10221);
nand U17474 (N_17474,N_11161,N_13507);
nor U17475 (N_17475,N_14586,N_13151);
nand U17476 (N_17476,N_13462,N_14280);
xnor U17477 (N_17477,N_14513,N_12895);
or U17478 (N_17478,N_12464,N_13812);
or U17479 (N_17479,N_11340,N_13469);
xor U17480 (N_17480,N_10511,N_10877);
nor U17481 (N_17481,N_10770,N_10372);
nand U17482 (N_17482,N_13095,N_10497);
nor U17483 (N_17483,N_12039,N_11662);
nor U17484 (N_17484,N_10184,N_14740);
or U17485 (N_17485,N_11342,N_10945);
or U17486 (N_17486,N_14573,N_10300);
and U17487 (N_17487,N_11606,N_12130);
nor U17488 (N_17488,N_11938,N_14544);
or U17489 (N_17489,N_14635,N_14463);
nand U17490 (N_17490,N_13268,N_13266);
and U17491 (N_17491,N_12952,N_12855);
xor U17492 (N_17492,N_11620,N_10575);
nor U17493 (N_17493,N_10737,N_10955);
nor U17494 (N_17494,N_13338,N_10074);
nand U17495 (N_17495,N_10032,N_14256);
and U17496 (N_17496,N_12245,N_14468);
nand U17497 (N_17497,N_14949,N_13177);
nand U17498 (N_17498,N_11269,N_10400);
or U17499 (N_17499,N_11574,N_11060);
xnor U17500 (N_17500,N_14347,N_13002);
nor U17501 (N_17501,N_11079,N_12626);
and U17502 (N_17502,N_13335,N_14965);
and U17503 (N_17503,N_14055,N_10158);
nand U17504 (N_17504,N_13294,N_12733);
or U17505 (N_17505,N_11350,N_12288);
and U17506 (N_17506,N_10627,N_13072);
xnor U17507 (N_17507,N_10066,N_11714);
and U17508 (N_17508,N_11656,N_11703);
nand U17509 (N_17509,N_11504,N_12520);
nor U17510 (N_17510,N_11726,N_14454);
nand U17511 (N_17511,N_13173,N_12988);
nor U17512 (N_17512,N_12409,N_10865);
nand U17513 (N_17513,N_14153,N_14135);
nor U17514 (N_17514,N_10515,N_11900);
xnor U17515 (N_17515,N_11280,N_13625);
nand U17516 (N_17516,N_14018,N_14945);
nand U17517 (N_17517,N_12707,N_10121);
nor U17518 (N_17518,N_14311,N_12137);
nor U17519 (N_17519,N_11793,N_12469);
or U17520 (N_17520,N_12497,N_10953);
nand U17521 (N_17521,N_11859,N_11938);
and U17522 (N_17522,N_11218,N_12186);
nand U17523 (N_17523,N_10589,N_13541);
nand U17524 (N_17524,N_13942,N_10863);
and U17525 (N_17525,N_14284,N_11571);
nand U17526 (N_17526,N_11835,N_11559);
nand U17527 (N_17527,N_11272,N_13941);
and U17528 (N_17528,N_12687,N_10989);
or U17529 (N_17529,N_14382,N_13714);
or U17530 (N_17530,N_13139,N_10700);
xor U17531 (N_17531,N_12904,N_13514);
and U17532 (N_17532,N_14413,N_10521);
nand U17533 (N_17533,N_12190,N_14184);
xnor U17534 (N_17534,N_11763,N_13862);
nand U17535 (N_17535,N_14870,N_10817);
nor U17536 (N_17536,N_11794,N_10250);
or U17537 (N_17537,N_10534,N_14978);
nor U17538 (N_17538,N_13404,N_10554);
and U17539 (N_17539,N_12342,N_14438);
and U17540 (N_17540,N_11016,N_14544);
nand U17541 (N_17541,N_13989,N_10691);
and U17542 (N_17542,N_14827,N_10667);
nand U17543 (N_17543,N_11447,N_13400);
nor U17544 (N_17544,N_13082,N_13535);
or U17545 (N_17545,N_12398,N_10297);
nor U17546 (N_17546,N_11978,N_12610);
nor U17547 (N_17547,N_10645,N_13616);
nand U17548 (N_17548,N_10244,N_14202);
nor U17549 (N_17549,N_10855,N_14257);
nand U17550 (N_17550,N_11001,N_13909);
nand U17551 (N_17551,N_10334,N_11472);
and U17552 (N_17552,N_13894,N_13732);
and U17553 (N_17553,N_14832,N_10999);
and U17554 (N_17554,N_14122,N_13052);
or U17555 (N_17555,N_12380,N_10804);
xor U17556 (N_17556,N_13502,N_10771);
xnor U17557 (N_17557,N_13949,N_11053);
and U17558 (N_17558,N_10232,N_10951);
nand U17559 (N_17559,N_13002,N_14225);
and U17560 (N_17560,N_13017,N_14669);
nor U17561 (N_17561,N_10195,N_14752);
xor U17562 (N_17562,N_10762,N_13868);
nor U17563 (N_17563,N_12617,N_10286);
and U17564 (N_17564,N_13167,N_14057);
xor U17565 (N_17565,N_12497,N_12280);
nand U17566 (N_17566,N_10344,N_11609);
and U17567 (N_17567,N_12749,N_14571);
nor U17568 (N_17568,N_10662,N_10056);
xnor U17569 (N_17569,N_12041,N_10048);
nor U17570 (N_17570,N_13300,N_13063);
or U17571 (N_17571,N_14185,N_13966);
nand U17572 (N_17572,N_11942,N_10193);
nand U17573 (N_17573,N_12645,N_14948);
and U17574 (N_17574,N_14989,N_10457);
nand U17575 (N_17575,N_13078,N_10547);
xor U17576 (N_17576,N_13820,N_11865);
or U17577 (N_17577,N_12792,N_10675);
nand U17578 (N_17578,N_13999,N_10336);
nor U17579 (N_17579,N_13035,N_14368);
and U17580 (N_17580,N_11074,N_13789);
or U17581 (N_17581,N_12879,N_10038);
or U17582 (N_17582,N_13469,N_11447);
nand U17583 (N_17583,N_13948,N_14838);
or U17584 (N_17584,N_14706,N_13084);
nor U17585 (N_17585,N_11457,N_11828);
xor U17586 (N_17586,N_14635,N_12345);
or U17587 (N_17587,N_14258,N_13912);
nor U17588 (N_17588,N_13358,N_12545);
and U17589 (N_17589,N_10111,N_13583);
xnor U17590 (N_17590,N_11666,N_12037);
nand U17591 (N_17591,N_13634,N_14992);
xor U17592 (N_17592,N_11629,N_13791);
or U17593 (N_17593,N_12844,N_14667);
nand U17594 (N_17594,N_10874,N_10370);
or U17595 (N_17595,N_11631,N_12729);
nand U17596 (N_17596,N_11009,N_10200);
nor U17597 (N_17597,N_12385,N_11821);
nand U17598 (N_17598,N_13423,N_10962);
nand U17599 (N_17599,N_12223,N_10510);
nor U17600 (N_17600,N_10838,N_14728);
and U17601 (N_17601,N_13984,N_14017);
and U17602 (N_17602,N_11032,N_13419);
and U17603 (N_17603,N_11356,N_11062);
or U17604 (N_17604,N_10747,N_10535);
or U17605 (N_17605,N_14362,N_10064);
and U17606 (N_17606,N_11472,N_12030);
and U17607 (N_17607,N_10094,N_10471);
and U17608 (N_17608,N_12623,N_10320);
and U17609 (N_17609,N_12050,N_10549);
nor U17610 (N_17610,N_10003,N_14160);
nor U17611 (N_17611,N_10806,N_13743);
and U17612 (N_17612,N_13990,N_12749);
or U17613 (N_17613,N_10307,N_10024);
nand U17614 (N_17614,N_11751,N_14966);
or U17615 (N_17615,N_12051,N_14458);
and U17616 (N_17616,N_14176,N_12302);
and U17617 (N_17617,N_13410,N_10567);
nor U17618 (N_17618,N_14700,N_12255);
and U17619 (N_17619,N_14700,N_13542);
xor U17620 (N_17620,N_12951,N_12135);
and U17621 (N_17621,N_11057,N_14753);
and U17622 (N_17622,N_14706,N_10138);
nand U17623 (N_17623,N_13713,N_12485);
nand U17624 (N_17624,N_10955,N_12258);
or U17625 (N_17625,N_10237,N_12192);
nand U17626 (N_17626,N_10752,N_10174);
nor U17627 (N_17627,N_14151,N_11128);
and U17628 (N_17628,N_10519,N_10752);
or U17629 (N_17629,N_10717,N_13067);
or U17630 (N_17630,N_12871,N_11194);
nor U17631 (N_17631,N_10742,N_11152);
nor U17632 (N_17632,N_10474,N_11419);
or U17633 (N_17633,N_14394,N_13863);
nand U17634 (N_17634,N_10806,N_13264);
nand U17635 (N_17635,N_11219,N_11862);
or U17636 (N_17636,N_10141,N_11617);
nand U17637 (N_17637,N_10462,N_10185);
nand U17638 (N_17638,N_14742,N_12660);
nor U17639 (N_17639,N_11221,N_14923);
or U17640 (N_17640,N_11893,N_11748);
and U17641 (N_17641,N_13608,N_14851);
or U17642 (N_17642,N_11575,N_13287);
nand U17643 (N_17643,N_11911,N_14267);
nand U17644 (N_17644,N_10633,N_10962);
nand U17645 (N_17645,N_14637,N_13549);
xor U17646 (N_17646,N_10247,N_13704);
nor U17647 (N_17647,N_12025,N_12105);
or U17648 (N_17648,N_13873,N_14608);
nand U17649 (N_17649,N_12203,N_11515);
or U17650 (N_17650,N_13991,N_11568);
and U17651 (N_17651,N_13764,N_13733);
nor U17652 (N_17652,N_10683,N_12851);
or U17653 (N_17653,N_10853,N_12742);
or U17654 (N_17654,N_12260,N_14530);
or U17655 (N_17655,N_12833,N_10914);
nor U17656 (N_17656,N_12415,N_14050);
nand U17657 (N_17657,N_14327,N_12883);
nand U17658 (N_17658,N_13280,N_14424);
nand U17659 (N_17659,N_13092,N_10112);
and U17660 (N_17660,N_13143,N_13927);
or U17661 (N_17661,N_10340,N_12105);
xor U17662 (N_17662,N_10283,N_12022);
nand U17663 (N_17663,N_11488,N_10481);
nor U17664 (N_17664,N_10340,N_14232);
or U17665 (N_17665,N_10144,N_11126);
and U17666 (N_17666,N_11151,N_11034);
nand U17667 (N_17667,N_14950,N_11731);
and U17668 (N_17668,N_14173,N_11622);
nand U17669 (N_17669,N_10300,N_12180);
or U17670 (N_17670,N_14285,N_14812);
and U17671 (N_17671,N_11731,N_11218);
nor U17672 (N_17672,N_14091,N_13502);
or U17673 (N_17673,N_14092,N_10529);
nand U17674 (N_17674,N_10164,N_10706);
or U17675 (N_17675,N_10627,N_13423);
nor U17676 (N_17676,N_11167,N_14523);
and U17677 (N_17677,N_12737,N_12546);
or U17678 (N_17678,N_14328,N_10321);
nor U17679 (N_17679,N_14861,N_12606);
nor U17680 (N_17680,N_10922,N_14136);
nand U17681 (N_17681,N_11049,N_13325);
nand U17682 (N_17682,N_14419,N_10606);
nand U17683 (N_17683,N_11176,N_10368);
nor U17684 (N_17684,N_12251,N_10626);
and U17685 (N_17685,N_14205,N_14954);
nand U17686 (N_17686,N_12241,N_14966);
nor U17687 (N_17687,N_14088,N_12862);
and U17688 (N_17688,N_11531,N_13283);
or U17689 (N_17689,N_13947,N_14402);
nand U17690 (N_17690,N_10691,N_14267);
or U17691 (N_17691,N_12483,N_14403);
xor U17692 (N_17692,N_12013,N_11517);
and U17693 (N_17693,N_11589,N_10162);
and U17694 (N_17694,N_10584,N_13811);
nor U17695 (N_17695,N_11909,N_12401);
or U17696 (N_17696,N_12509,N_10844);
nor U17697 (N_17697,N_13952,N_12800);
xor U17698 (N_17698,N_14436,N_11923);
and U17699 (N_17699,N_11350,N_11906);
nor U17700 (N_17700,N_12839,N_14780);
nand U17701 (N_17701,N_13664,N_12965);
or U17702 (N_17702,N_13116,N_14023);
nand U17703 (N_17703,N_14804,N_11242);
or U17704 (N_17704,N_10586,N_12112);
or U17705 (N_17705,N_13650,N_11415);
and U17706 (N_17706,N_13992,N_14145);
or U17707 (N_17707,N_10453,N_13185);
xnor U17708 (N_17708,N_10156,N_11441);
nor U17709 (N_17709,N_14586,N_14567);
and U17710 (N_17710,N_13260,N_11738);
xnor U17711 (N_17711,N_14850,N_11213);
nor U17712 (N_17712,N_10991,N_10306);
xor U17713 (N_17713,N_13156,N_13486);
and U17714 (N_17714,N_11476,N_10637);
and U17715 (N_17715,N_10993,N_14014);
and U17716 (N_17716,N_14734,N_12543);
or U17717 (N_17717,N_11786,N_14228);
nand U17718 (N_17718,N_11334,N_14563);
or U17719 (N_17719,N_14076,N_12780);
nand U17720 (N_17720,N_13368,N_14965);
or U17721 (N_17721,N_14630,N_10834);
nand U17722 (N_17722,N_13498,N_13568);
nor U17723 (N_17723,N_13972,N_14205);
and U17724 (N_17724,N_10035,N_13448);
and U17725 (N_17725,N_14436,N_11129);
nand U17726 (N_17726,N_11502,N_14800);
nor U17727 (N_17727,N_13167,N_14493);
and U17728 (N_17728,N_13513,N_10902);
nor U17729 (N_17729,N_13850,N_12135);
nand U17730 (N_17730,N_13286,N_11000);
nor U17731 (N_17731,N_10209,N_10060);
nor U17732 (N_17732,N_13172,N_12930);
nor U17733 (N_17733,N_10884,N_11744);
nand U17734 (N_17734,N_11847,N_11027);
nor U17735 (N_17735,N_14953,N_14272);
nand U17736 (N_17736,N_14575,N_12931);
nor U17737 (N_17737,N_13384,N_14829);
nor U17738 (N_17738,N_10184,N_10630);
nand U17739 (N_17739,N_14654,N_13936);
and U17740 (N_17740,N_14132,N_14787);
and U17741 (N_17741,N_10259,N_11893);
nand U17742 (N_17742,N_11931,N_10819);
or U17743 (N_17743,N_12318,N_13481);
nand U17744 (N_17744,N_14353,N_13573);
and U17745 (N_17745,N_10332,N_14626);
or U17746 (N_17746,N_10990,N_13030);
and U17747 (N_17747,N_10838,N_14312);
or U17748 (N_17748,N_11053,N_12885);
nor U17749 (N_17749,N_10985,N_11440);
nand U17750 (N_17750,N_12872,N_14078);
nand U17751 (N_17751,N_12378,N_14611);
nor U17752 (N_17752,N_13934,N_14503);
nand U17753 (N_17753,N_12435,N_11028);
or U17754 (N_17754,N_13234,N_10236);
nand U17755 (N_17755,N_11476,N_11934);
or U17756 (N_17756,N_12551,N_11662);
and U17757 (N_17757,N_12902,N_10088);
and U17758 (N_17758,N_14049,N_10179);
and U17759 (N_17759,N_11926,N_11794);
nand U17760 (N_17760,N_13296,N_12562);
and U17761 (N_17761,N_12851,N_14509);
nor U17762 (N_17762,N_10404,N_13073);
nor U17763 (N_17763,N_12277,N_10272);
nand U17764 (N_17764,N_13011,N_12436);
or U17765 (N_17765,N_11132,N_13168);
and U17766 (N_17766,N_11347,N_10531);
nand U17767 (N_17767,N_14766,N_10329);
and U17768 (N_17768,N_10441,N_11742);
nand U17769 (N_17769,N_14278,N_12456);
or U17770 (N_17770,N_14157,N_12788);
and U17771 (N_17771,N_13139,N_10046);
nor U17772 (N_17772,N_13978,N_13251);
or U17773 (N_17773,N_13421,N_10095);
xnor U17774 (N_17774,N_10027,N_10213);
and U17775 (N_17775,N_10169,N_12476);
nor U17776 (N_17776,N_13114,N_13974);
nor U17777 (N_17777,N_12887,N_10588);
nor U17778 (N_17778,N_11419,N_11433);
and U17779 (N_17779,N_11477,N_11534);
and U17780 (N_17780,N_10030,N_13819);
or U17781 (N_17781,N_12098,N_13954);
nor U17782 (N_17782,N_12016,N_11807);
nand U17783 (N_17783,N_14959,N_10848);
and U17784 (N_17784,N_11859,N_13074);
and U17785 (N_17785,N_10988,N_14066);
nor U17786 (N_17786,N_12427,N_10171);
nand U17787 (N_17787,N_13695,N_12805);
nor U17788 (N_17788,N_10089,N_13756);
and U17789 (N_17789,N_12568,N_10591);
nor U17790 (N_17790,N_13868,N_13519);
or U17791 (N_17791,N_14188,N_13983);
nor U17792 (N_17792,N_14065,N_13045);
nor U17793 (N_17793,N_13610,N_10061);
and U17794 (N_17794,N_12596,N_12210);
xnor U17795 (N_17795,N_11513,N_10097);
or U17796 (N_17796,N_14907,N_12965);
and U17797 (N_17797,N_13221,N_14758);
nand U17798 (N_17798,N_10251,N_14493);
nor U17799 (N_17799,N_10007,N_14370);
nand U17800 (N_17800,N_10457,N_14453);
nor U17801 (N_17801,N_10299,N_11487);
and U17802 (N_17802,N_10845,N_12780);
or U17803 (N_17803,N_10108,N_10561);
or U17804 (N_17804,N_10092,N_10162);
or U17805 (N_17805,N_13143,N_14170);
and U17806 (N_17806,N_12257,N_13552);
nand U17807 (N_17807,N_11316,N_13743);
nand U17808 (N_17808,N_11484,N_14876);
and U17809 (N_17809,N_12401,N_10726);
or U17810 (N_17810,N_12080,N_14705);
nor U17811 (N_17811,N_14785,N_10575);
and U17812 (N_17812,N_11332,N_10949);
or U17813 (N_17813,N_14925,N_13669);
nor U17814 (N_17814,N_11276,N_14799);
nor U17815 (N_17815,N_10215,N_14225);
nor U17816 (N_17816,N_12296,N_13110);
or U17817 (N_17817,N_10370,N_12498);
and U17818 (N_17818,N_13212,N_14733);
nor U17819 (N_17819,N_12657,N_10766);
nor U17820 (N_17820,N_13039,N_12515);
and U17821 (N_17821,N_12175,N_11950);
nor U17822 (N_17822,N_10382,N_13187);
nor U17823 (N_17823,N_10105,N_12230);
nand U17824 (N_17824,N_11895,N_12428);
or U17825 (N_17825,N_12570,N_12992);
nand U17826 (N_17826,N_11533,N_13063);
or U17827 (N_17827,N_12442,N_14030);
and U17828 (N_17828,N_12979,N_11170);
nor U17829 (N_17829,N_14023,N_12072);
nor U17830 (N_17830,N_11262,N_14889);
xor U17831 (N_17831,N_13972,N_10005);
nand U17832 (N_17832,N_12959,N_14809);
or U17833 (N_17833,N_13061,N_14422);
nand U17834 (N_17834,N_12781,N_12448);
nor U17835 (N_17835,N_10191,N_14549);
or U17836 (N_17836,N_12017,N_12275);
or U17837 (N_17837,N_13296,N_14697);
nor U17838 (N_17838,N_14981,N_14170);
or U17839 (N_17839,N_10595,N_12080);
and U17840 (N_17840,N_12575,N_12018);
xor U17841 (N_17841,N_12474,N_12666);
and U17842 (N_17842,N_11799,N_10756);
nand U17843 (N_17843,N_14442,N_13389);
nor U17844 (N_17844,N_11856,N_14011);
nor U17845 (N_17845,N_13781,N_10904);
nand U17846 (N_17846,N_12879,N_12829);
and U17847 (N_17847,N_13770,N_13538);
and U17848 (N_17848,N_14220,N_12324);
nor U17849 (N_17849,N_10257,N_12667);
and U17850 (N_17850,N_14573,N_12867);
and U17851 (N_17851,N_11927,N_14004);
xnor U17852 (N_17852,N_14413,N_12630);
nor U17853 (N_17853,N_14868,N_14519);
xnor U17854 (N_17854,N_13435,N_12661);
nand U17855 (N_17855,N_10275,N_11565);
nand U17856 (N_17856,N_11435,N_13361);
and U17857 (N_17857,N_14112,N_14077);
nor U17858 (N_17858,N_11312,N_10094);
or U17859 (N_17859,N_14304,N_13583);
xor U17860 (N_17860,N_12299,N_14029);
and U17861 (N_17861,N_11584,N_14432);
nor U17862 (N_17862,N_14707,N_12021);
nor U17863 (N_17863,N_14080,N_14379);
and U17864 (N_17864,N_14375,N_13397);
nand U17865 (N_17865,N_14553,N_14803);
nand U17866 (N_17866,N_11339,N_12317);
or U17867 (N_17867,N_12082,N_13929);
and U17868 (N_17868,N_13724,N_12219);
nand U17869 (N_17869,N_10169,N_14019);
or U17870 (N_17870,N_10251,N_14179);
nor U17871 (N_17871,N_13093,N_10771);
and U17872 (N_17872,N_12464,N_12031);
xor U17873 (N_17873,N_12923,N_13080);
or U17874 (N_17874,N_11981,N_14647);
nor U17875 (N_17875,N_13190,N_11331);
nand U17876 (N_17876,N_13302,N_11602);
nor U17877 (N_17877,N_10414,N_13651);
or U17878 (N_17878,N_14250,N_13237);
nor U17879 (N_17879,N_12684,N_13230);
or U17880 (N_17880,N_13924,N_10911);
nor U17881 (N_17881,N_12050,N_10592);
and U17882 (N_17882,N_11330,N_13656);
and U17883 (N_17883,N_12880,N_12692);
and U17884 (N_17884,N_13120,N_11669);
or U17885 (N_17885,N_11167,N_10095);
nand U17886 (N_17886,N_11903,N_11009);
xor U17887 (N_17887,N_14738,N_11367);
xnor U17888 (N_17888,N_11040,N_12876);
or U17889 (N_17889,N_14644,N_12446);
nor U17890 (N_17890,N_13667,N_13817);
nand U17891 (N_17891,N_14152,N_14724);
nand U17892 (N_17892,N_12351,N_12015);
nand U17893 (N_17893,N_11264,N_11000);
nand U17894 (N_17894,N_13264,N_10600);
xnor U17895 (N_17895,N_10387,N_11646);
or U17896 (N_17896,N_12191,N_13795);
or U17897 (N_17897,N_12397,N_13531);
and U17898 (N_17898,N_10483,N_13227);
nor U17899 (N_17899,N_12380,N_14475);
nor U17900 (N_17900,N_10611,N_10457);
or U17901 (N_17901,N_10388,N_13219);
and U17902 (N_17902,N_12227,N_13560);
nand U17903 (N_17903,N_13899,N_12642);
nor U17904 (N_17904,N_11922,N_10045);
and U17905 (N_17905,N_11034,N_13957);
nand U17906 (N_17906,N_12311,N_14915);
nor U17907 (N_17907,N_14143,N_12550);
and U17908 (N_17908,N_12610,N_13643);
nor U17909 (N_17909,N_11315,N_13290);
or U17910 (N_17910,N_11016,N_14975);
nand U17911 (N_17911,N_12974,N_13115);
nor U17912 (N_17912,N_13353,N_10198);
nor U17913 (N_17913,N_13417,N_14799);
nor U17914 (N_17914,N_11617,N_12066);
nor U17915 (N_17915,N_10544,N_10821);
nor U17916 (N_17916,N_11845,N_11377);
nor U17917 (N_17917,N_13357,N_13933);
and U17918 (N_17918,N_13643,N_11906);
nor U17919 (N_17919,N_10604,N_13468);
xor U17920 (N_17920,N_10802,N_14961);
and U17921 (N_17921,N_13037,N_10831);
nor U17922 (N_17922,N_11419,N_11170);
nand U17923 (N_17923,N_14632,N_11573);
nand U17924 (N_17924,N_13746,N_14550);
nand U17925 (N_17925,N_13671,N_10235);
or U17926 (N_17926,N_13612,N_14537);
or U17927 (N_17927,N_13466,N_11979);
nor U17928 (N_17928,N_12000,N_12610);
and U17929 (N_17929,N_14697,N_13084);
and U17930 (N_17930,N_10138,N_10937);
nand U17931 (N_17931,N_11920,N_14061);
nand U17932 (N_17932,N_12373,N_10884);
or U17933 (N_17933,N_11301,N_12622);
nor U17934 (N_17934,N_13721,N_14882);
nor U17935 (N_17935,N_14773,N_12928);
and U17936 (N_17936,N_14128,N_10846);
and U17937 (N_17937,N_13531,N_12196);
and U17938 (N_17938,N_10647,N_13365);
and U17939 (N_17939,N_10513,N_13559);
and U17940 (N_17940,N_13123,N_10514);
or U17941 (N_17941,N_11916,N_11748);
or U17942 (N_17942,N_10176,N_11535);
or U17943 (N_17943,N_11898,N_11626);
nor U17944 (N_17944,N_14875,N_10499);
and U17945 (N_17945,N_11175,N_12685);
xor U17946 (N_17946,N_10125,N_14212);
nand U17947 (N_17947,N_10375,N_10006);
xnor U17948 (N_17948,N_10726,N_14326);
or U17949 (N_17949,N_10187,N_12971);
and U17950 (N_17950,N_10812,N_10209);
nor U17951 (N_17951,N_10544,N_13334);
and U17952 (N_17952,N_11936,N_14373);
nand U17953 (N_17953,N_11843,N_13291);
or U17954 (N_17954,N_10389,N_10818);
and U17955 (N_17955,N_10835,N_13773);
nand U17956 (N_17956,N_11842,N_12086);
nand U17957 (N_17957,N_11511,N_13295);
nand U17958 (N_17958,N_14228,N_12194);
or U17959 (N_17959,N_10376,N_12560);
xor U17960 (N_17960,N_11456,N_10834);
or U17961 (N_17961,N_12861,N_12997);
and U17962 (N_17962,N_10806,N_13471);
or U17963 (N_17963,N_13541,N_13138);
or U17964 (N_17964,N_14015,N_13932);
nor U17965 (N_17965,N_12464,N_12202);
and U17966 (N_17966,N_13039,N_11603);
and U17967 (N_17967,N_13303,N_12069);
nand U17968 (N_17968,N_11286,N_14719);
or U17969 (N_17969,N_10948,N_12455);
nand U17970 (N_17970,N_14171,N_13888);
and U17971 (N_17971,N_12094,N_14614);
or U17972 (N_17972,N_13723,N_12466);
nor U17973 (N_17973,N_14485,N_12097);
or U17974 (N_17974,N_10524,N_10126);
and U17975 (N_17975,N_14593,N_14559);
or U17976 (N_17976,N_14691,N_10867);
xnor U17977 (N_17977,N_12787,N_14885);
and U17978 (N_17978,N_10547,N_10794);
xnor U17979 (N_17979,N_13053,N_10633);
nor U17980 (N_17980,N_11439,N_12000);
nand U17981 (N_17981,N_10569,N_13336);
or U17982 (N_17982,N_11036,N_12474);
nand U17983 (N_17983,N_12592,N_13043);
nor U17984 (N_17984,N_14385,N_10151);
xnor U17985 (N_17985,N_13904,N_13043);
and U17986 (N_17986,N_14781,N_10659);
xnor U17987 (N_17987,N_11952,N_10640);
nor U17988 (N_17988,N_11034,N_13464);
xnor U17989 (N_17989,N_11079,N_11937);
xnor U17990 (N_17990,N_13899,N_10672);
nand U17991 (N_17991,N_10010,N_10831);
xnor U17992 (N_17992,N_14717,N_13401);
nand U17993 (N_17993,N_10256,N_10797);
and U17994 (N_17994,N_14346,N_10555);
or U17995 (N_17995,N_13772,N_13028);
nand U17996 (N_17996,N_13226,N_14312);
nand U17997 (N_17997,N_11106,N_12436);
and U17998 (N_17998,N_10600,N_13493);
nand U17999 (N_17999,N_10224,N_11398);
and U18000 (N_18000,N_13961,N_13823);
and U18001 (N_18001,N_10995,N_12299);
nand U18002 (N_18002,N_13713,N_13449);
nor U18003 (N_18003,N_11916,N_11347);
or U18004 (N_18004,N_10091,N_14360);
and U18005 (N_18005,N_13704,N_13389);
or U18006 (N_18006,N_11841,N_14063);
and U18007 (N_18007,N_12099,N_12420);
nand U18008 (N_18008,N_14232,N_11618);
or U18009 (N_18009,N_10543,N_11990);
or U18010 (N_18010,N_14118,N_11062);
xnor U18011 (N_18011,N_12654,N_12271);
xor U18012 (N_18012,N_11557,N_12083);
nand U18013 (N_18013,N_13514,N_11928);
nand U18014 (N_18014,N_10167,N_11615);
xnor U18015 (N_18015,N_13745,N_11244);
nor U18016 (N_18016,N_12326,N_14752);
or U18017 (N_18017,N_13191,N_14485);
xor U18018 (N_18018,N_12939,N_10225);
nand U18019 (N_18019,N_11530,N_13716);
or U18020 (N_18020,N_10250,N_12481);
nand U18021 (N_18021,N_11039,N_11744);
and U18022 (N_18022,N_11293,N_10507);
nor U18023 (N_18023,N_10002,N_12679);
and U18024 (N_18024,N_10182,N_10538);
and U18025 (N_18025,N_13166,N_14311);
or U18026 (N_18026,N_12790,N_11103);
or U18027 (N_18027,N_12655,N_14643);
nor U18028 (N_18028,N_14994,N_13969);
nor U18029 (N_18029,N_12811,N_10655);
or U18030 (N_18030,N_11738,N_14019);
nor U18031 (N_18031,N_10487,N_14505);
and U18032 (N_18032,N_12787,N_10040);
and U18033 (N_18033,N_14278,N_11106);
and U18034 (N_18034,N_10012,N_10756);
and U18035 (N_18035,N_12794,N_10586);
and U18036 (N_18036,N_11378,N_13329);
xnor U18037 (N_18037,N_12651,N_13737);
nor U18038 (N_18038,N_14639,N_10373);
nand U18039 (N_18039,N_14271,N_14372);
and U18040 (N_18040,N_11331,N_10943);
xor U18041 (N_18041,N_13310,N_12701);
and U18042 (N_18042,N_14003,N_13276);
xor U18043 (N_18043,N_12285,N_12166);
xor U18044 (N_18044,N_12898,N_10873);
nand U18045 (N_18045,N_12805,N_11706);
nor U18046 (N_18046,N_14930,N_11475);
or U18047 (N_18047,N_11336,N_13174);
xor U18048 (N_18048,N_13469,N_12948);
nor U18049 (N_18049,N_11145,N_12239);
nor U18050 (N_18050,N_14823,N_12393);
and U18051 (N_18051,N_10128,N_14211);
nand U18052 (N_18052,N_10426,N_12371);
and U18053 (N_18053,N_14083,N_13032);
nor U18054 (N_18054,N_11187,N_13170);
or U18055 (N_18055,N_13342,N_10412);
and U18056 (N_18056,N_13587,N_12996);
or U18057 (N_18057,N_14425,N_12395);
xor U18058 (N_18058,N_12579,N_11029);
xor U18059 (N_18059,N_11104,N_14843);
nand U18060 (N_18060,N_10053,N_12962);
xnor U18061 (N_18061,N_11524,N_14283);
nand U18062 (N_18062,N_14425,N_10453);
nand U18063 (N_18063,N_10767,N_10342);
nor U18064 (N_18064,N_14299,N_11896);
xnor U18065 (N_18065,N_12322,N_12969);
nand U18066 (N_18066,N_14251,N_13074);
nand U18067 (N_18067,N_14318,N_14075);
and U18068 (N_18068,N_13714,N_11268);
and U18069 (N_18069,N_10297,N_12133);
and U18070 (N_18070,N_14933,N_13770);
or U18071 (N_18071,N_11233,N_13103);
nor U18072 (N_18072,N_13592,N_14488);
and U18073 (N_18073,N_12699,N_12868);
nand U18074 (N_18074,N_11545,N_14102);
nand U18075 (N_18075,N_13818,N_12321);
and U18076 (N_18076,N_10410,N_11212);
nand U18077 (N_18077,N_14932,N_12713);
and U18078 (N_18078,N_14490,N_13080);
or U18079 (N_18079,N_12813,N_11525);
nand U18080 (N_18080,N_10183,N_12238);
or U18081 (N_18081,N_14326,N_12220);
and U18082 (N_18082,N_12169,N_10126);
or U18083 (N_18083,N_11013,N_13136);
nor U18084 (N_18084,N_12644,N_12277);
and U18085 (N_18085,N_14569,N_14561);
nor U18086 (N_18086,N_13249,N_13460);
nand U18087 (N_18087,N_10440,N_14638);
or U18088 (N_18088,N_14398,N_14694);
nand U18089 (N_18089,N_11798,N_13919);
nand U18090 (N_18090,N_10836,N_12672);
and U18091 (N_18091,N_12938,N_10472);
nor U18092 (N_18092,N_13390,N_14393);
and U18093 (N_18093,N_10891,N_10106);
and U18094 (N_18094,N_12684,N_14419);
nor U18095 (N_18095,N_12652,N_13052);
nand U18096 (N_18096,N_11624,N_14658);
and U18097 (N_18097,N_11201,N_10985);
or U18098 (N_18098,N_12414,N_11624);
or U18099 (N_18099,N_10502,N_12701);
or U18100 (N_18100,N_11038,N_13663);
nor U18101 (N_18101,N_13179,N_10961);
nand U18102 (N_18102,N_14989,N_12448);
nor U18103 (N_18103,N_12768,N_14792);
nand U18104 (N_18104,N_12997,N_10655);
nor U18105 (N_18105,N_10115,N_10900);
xnor U18106 (N_18106,N_10113,N_10477);
nand U18107 (N_18107,N_14309,N_14238);
or U18108 (N_18108,N_13502,N_12009);
nor U18109 (N_18109,N_11518,N_13586);
and U18110 (N_18110,N_10769,N_13264);
xnor U18111 (N_18111,N_12647,N_13722);
nand U18112 (N_18112,N_11299,N_14421);
or U18113 (N_18113,N_13216,N_13881);
and U18114 (N_18114,N_13020,N_13436);
and U18115 (N_18115,N_12323,N_13320);
or U18116 (N_18116,N_12504,N_10335);
and U18117 (N_18117,N_11375,N_11980);
and U18118 (N_18118,N_12743,N_11444);
nor U18119 (N_18119,N_11872,N_11935);
and U18120 (N_18120,N_10001,N_14986);
and U18121 (N_18121,N_14318,N_14265);
and U18122 (N_18122,N_14170,N_12983);
and U18123 (N_18123,N_11008,N_14860);
nand U18124 (N_18124,N_14614,N_12065);
nand U18125 (N_18125,N_13266,N_14390);
and U18126 (N_18126,N_13690,N_10865);
and U18127 (N_18127,N_11398,N_11810);
nand U18128 (N_18128,N_14648,N_12956);
nand U18129 (N_18129,N_12540,N_13927);
or U18130 (N_18130,N_11847,N_13050);
nand U18131 (N_18131,N_11182,N_12729);
nor U18132 (N_18132,N_11555,N_10310);
or U18133 (N_18133,N_12319,N_14780);
nand U18134 (N_18134,N_11724,N_12979);
and U18135 (N_18135,N_12101,N_11188);
nor U18136 (N_18136,N_10913,N_12628);
xor U18137 (N_18137,N_10193,N_12242);
nand U18138 (N_18138,N_13065,N_14312);
nand U18139 (N_18139,N_12896,N_13487);
xnor U18140 (N_18140,N_13161,N_10067);
nand U18141 (N_18141,N_12664,N_12283);
nand U18142 (N_18142,N_12400,N_11902);
nor U18143 (N_18143,N_10531,N_13707);
nand U18144 (N_18144,N_13627,N_14930);
nand U18145 (N_18145,N_12890,N_13971);
or U18146 (N_18146,N_13147,N_11260);
nand U18147 (N_18147,N_12489,N_10535);
or U18148 (N_18148,N_11578,N_14253);
and U18149 (N_18149,N_13436,N_10204);
or U18150 (N_18150,N_13341,N_13244);
xnor U18151 (N_18151,N_14248,N_12468);
and U18152 (N_18152,N_10892,N_13311);
nor U18153 (N_18153,N_10512,N_13041);
and U18154 (N_18154,N_10564,N_13549);
xnor U18155 (N_18155,N_10335,N_14543);
or U18156 (N_18156,N_14967,N_11591);
and U18157 (N_18157,N_12607,N_13941);
xnor U18158 (N_18158,N_12571,N_10601);
nand U18159 (N_18159,N_13608,N_10510);
xnor U18160 (N_18160,N_13917,N_12649);
nor U18161 (N_18161,N_12396,N_10655);
nor U18162 (N_18162,N_13536,N_10027);
nand U18163 (N_18163,N_13170,N_14342);
xnor U18164 (N_18164,N_11815,N_14538);
xor U18165 (N_18165,N_12201,N_13279);
nor U18166 (N_18166,N_10092,N_13434);
or U18167 (N_18167,N_13973,N_10968);
nor U18168 (N_18168,N_14802,N_14037);
and U18169 (N_18169,N_11261,N_14626);
and U18170 (N_18170,N_11375,N_13139);
xor U18171 (N_18171,N_14908,N_14614);
and U18172 (N_18172,N_12821,N_10845);
nand U18173 (N_18173,N_14116,N_10838);
nand U18174 (N_18174,N_11888,N_13277);
or U18175 (N_18175,N_10241,N_10083);
or U18176 (N_18176,N_14216,N_11991);
nor U18177 (N_18177,N_11718,N_11411);
nand U18178 (N_18178,N_11987,N_11030);
nor U18179 (N_18179,N_14275,N_13776);
nor U18180 (N_18180,N_13261,N_14013);
and U18181 (N_18181,N_12271,N_10111);
or U18182 (N_18182,N_12589,N_13974);
nand U18183 (N_18183,N_14129,N_12746);
or U18184 (N_18184,N_12010,N_14798);
or U18185 (N_18185,N_12154,N_14329);
or U18186 (N_18186,N_11579,N_10082);
nor U18187 (N_18187,N_11590,N_11739);
and U18188 (N_18188,N_14548,N_13004);
or U18189 (N_18189,N_14836,N_11580);
nor U18190 (N_18190,N_10661,N_11901);
and U18191 (N_18191,N_12466,N_11195);
nor U18192 (N_18192,N_12912,N_12479);
nand U18193 (N_18193,N_13782,N_11531);
and U18194 (N_18194,N_10339,N_14689);
nor U18195 (N_18195,N_10515,N_13257);
nand U18196 (N_18196,N_13379,N_14709);
nand U18197 (N_18197,N_14970,N_11996);
and U18198 (N_18198,N_11820,N_11979);
nand U18199 (N_18199,N_11061,N_10229);
or U18200 (N_18200,N_14567,N_14678);
or U18201 (N_18201,N_10791,N_11859);
nand U18202 (N_18202,N_13253,N_14674);
nor U18203 (N_18203,N_14758,N_13229);
xor U18204 (N_18204,N_10833,N_11784);
and U18205 (N_18205,N_12569,N_11080);
nor U18206 (N_18206,N_12758,N_12068);
nor U18207 (N_18207,N_13684,N_11117);
xnor U18208 (N_18208,N_14392,N_12061);
nor U18209 (N_18209,N_12629,N_10083);
nor U18210 (N_18210,N_10509,N_14998);
and U18211 (N_18211,N_13372,N_11197);
or U18212 (N_18212,N_12597,N_13915);
and U18213 (N_18213,N_12926,N_12236);
xnor U18214 (N_18214,N_11284,N_11102);
nor U18215 (N_18215,N_13066,N_12548);
or U18216 (N_18216,N_13264,N_11617);
and U18217 (N_18217,N_12757,N_13982);
and U18218 (N_18218,N_14230,N_10505);
xor U18219 (N_18219,N_10478,N_11754);
and U18220 (N_18220,N_10243,N_10770);
nand U18221 (N_18221,N_13258,N_13961);
and U18222 (N_18222,N_11154,N_14303);
nand U18223 (N_18223,N_14595,N_11846);
and U18224 (N_18224,N_11638,N_10438);
and U18225 (N_18225,N_13229,N_12687);
nor U18226 (N_18226,N_11188,N_11267);
or U18227 (N_18227,N_12353,N_10451);
nand U18228 (N_18228,N_13638,N_10785);
and U18229 (N_18229,N_10706,N_12288);
xor U18230 (N_18230,N_10882,N_13028);
nor U18231 (N_18231,N_10427,N_12995);
nand U18232 (N_18232,N_10786,N_11665);
nand U18233 (N_18233,N_14065,N_10776);
xnor U18234 (N_18234,N_14000,N_11391);
nor U18235 (N_18235,N_10435,N_13560);
nor U18236 (N_18236,N_11301,N_13088);
nor U18237 (N_18237,N_12426,N_14438);
nand U18238 (N_18238,N_10191,N_14712);
or U18239 (N_18239,N_13738,N_14203);
nand U18240 (N_18240,N_14279,N_13980);
and U18241 (N_18241,N_11111,N_14338);
xor U18242 (N_18242,N_11046,N_14364);
nand U18243 (N_18243,N_12811,N_12351);
nand U18244 (N_18244,N_14440,N_10081);
nand U18245 (N_18245,N_11197,N_11557);
and U18246 (N_18246,N_11277,N_12574);
or U18247 (N_18247,N_12329,N_10513);
nor U18248 (N_18248,N_13459,N_11435);
xnor U18249 (N_18249,N_12177,N_12280);
nand U18250 (N_18250,N_11789,N_13977);
nor U18251 (N_18251,N_13168,N_12972);
and U18252 (N_18252,N_12633,N_13328);
or U18253 (N_18253,N_14566,N_12435);
nand U18254 (N_18254,N_10302,N_14364);
xor U18255 (N_18255,N_10740,N_13083);
nand U18256 (N_18256,N_14677,N_13964);
xnor U18257 (N_18257,N_13099,N_13188);
nand U18258 (N_18258,N_13192,N_12631);
nor U18259 (N_18259,N_14571,N_13625);
and U18260 (N_18260,N_12964,N_12634);
nand U18261 (N_18261,N_10227,N_14314);
and U18262 (N_18262,N_11950,N_11399);
or U18263 (N_18263,N_11400,N_14448);
nand U18264 (N_18264,N_10127,N_12912);
and U18265 (N_18265,N_12028,N_14281);
and U18266 (N_18266,N_11682,N_13678);
nor U18267 (N_18267,N_10201,N_10712);
or U18268 (N_18268,N_13402,N_11517);
or U18269 (N_18269,N_10087,N_10430);
nor U18270 (N_18270,N_10644,N_11021);
or U18271 (N_18271,N_10280,N_11200);
nor U18272 (N_18272,N_10301,N_11673);
or U18273 (N_18273,N_12631,N_13943);
or U18274 (N_18274,N_10758,N_14757);
and U18275 (N_18275,N_14200,N_11986);
nand U18276 (N_18276,N_13654,N_12727);
or U18277 (N_18277,N_14733,N_10408);
and U18278 (N_18278,N_13469,N_12177);
nand U18279 (N_18279,N_12951,N_13530);
or U18280 (N_18280,N_14554,N_10462);
and U18281 (N_18281,N_13092,N_14143);
xor U18282 (N_18282,N_11437,N_12130);
nand U18283 (N_18283,N_12277,N_10948);
nand U18284 (N_18284,N_14953,N_12189);
nand U18285 (N_18285,N_10528,N_12762);
nor U18286 (N_18286,N_10581,N_13635);
nor U18287 (N_18287,N_13423,N_14182);
nor U18288 (N_18288,N_11303,N_12283);
nand U18289 (N_18289,N_12696,N_14860);
and U18290 (N_18290,N_12894,N_11163);
xnor U18291 (N_18291,N_11037,N_13986);
and U18292 (N_18292,N_11965,N_12840);
and U18293 (N_18293,N_11421,N_10790);
and U18294 (N_18294,N_13369,N_14635);
nor U18295 (N_18295,N_14149,N_14300);
nor U18296 (N_18296,N_12612,N_10864);
and U18297 (N_18297,N_10059,N_12532);
nand U18298 (N_18298,N_10117,N_10642);
and U18299 (N_18299,N_12512,N_11890);
nand U18300 (N_18300,N_14522,N_10805);
and U18301 (N_18301,N_12332,N_11726);
nand U18302 (N_18302,N_13333,N_14492);
or U18303 (N_18303,N_14250,N_10571);
or U18304 (N_18304,N_10565,N_11073);
nand U18305 (N_18305,N_11319,N_13155);
or U18306 (N_18306,N_10208,N_14276);
and U18307 (N_18307,N_10506,N_10175);
nand U18308 (N_18308,N_12262,N_12188);
nand U18309 (N_18309,N_10581,N_13587);
and U18310 (N_18310,N_13365,N_14275);
nor U18311 (N_18311,N_13931,N_10005);
xor U18312 (N_18312,N_11263,N_11215);
and U18313 (N_18313,N_10850,N_10821);
xor U18314 (N_18314,N_12482,N_11289);
xor U18315 (N_18315,N_12093,N_11048);
or U18316 (N_18316,N_13227,N_12550);
nand U18317 (N_18317,N_13848,N_12316);
and U18318 (N_18318,N_12737,N_12119);
nand U18319 (N_18319,N_12082,N_10831);
nor U18320 (N_18320,N_13667,N_10876);
or U18321 (N_18321,N_14976,N_14697);
nand U18322 (N_18322,N_14320,N_10661);
and U18323 (N_18323,N_14835,N_10054);
xor U18324 (N_18324,N_14148,N_13232);
nand U18325 (N_18325,N_12805,N_10948);
nor U18326 (N_18326,N_13653,N_12450);
nand U18327 (N_18327,N_10267,N_14025);
nor U18328 (N_18328,N_13585,N_10728);
or U18329 (N_18329,N_14824,N_10355);
nor U18330 (N_18330,N_13660,N_10066);
and U18331 (N_18331,N_13629,N_13077);
nand U18332 (N_18332,N_11218,N_14350);
or U18333 (N_18333,N_12918,N_12334);
and U18334 (N_18334,N_13072,N_12316);
nand U18335 (N_18335,N_12817,N_14788);
and U18336 (N_18336,N_11794,N_11048);
nand U18337 (N_18337,N_14072,N_12639);
and U18338 (N_18338,N_13882,N_11147);
xnor U18339 (N_18339,N_12080,N_13146);
nand U18340 (N_18340,N_14268,N_13011);
nor U18341 (N_18341,N_11319,N_11314);
nand U18342 (N_18342,N_10253,N_14569);
and U18343 (N_18343,N_14896,N_12247);
nor U18344 (N_18344,N_10042,N_12550);
nor U18345 (N_18345,N_11606,N_11751);
nor U18346 (N_18346,N_11180,N_12859);
and U18347 (N_18347,N_10235,N_13036);
and U18348 (N_18348,N_12462,N_14019);
nand U18349 (N_18349,N_11328,N_14929);
and U18350 (N_18350,N_14511,N_10511);
nor U18351 (N_18351,N_12106,N_14107);
and U18352 (N_18352,N_11659,N_13377);
nor U18353 (N_18353,N_12485,N_10108);
nor U18354 (N_18354,N_13212,N_11541);
and U18355 (N_18355,N_13337,N_11179);
or U18356 (N_18356,N_10598,N_12722);
nand U18357 (N_18357,N_13825,N_10221);
nor U18358 (N_18358,N_11868,N_11475);
and U18359 (N_18359,N_10014,N_12085);
xor U18360 (N_18360,N_13451,N_11450);
and U18361 (N_18361,N_10786,N_13711);
nand U18362 (N_18362,N_14128,N_14076);
nand U18363 (N_18363,N_11434,N_10401);
nand U18364 (N_18364,N_10497,N_10648);
nor U18365 (N_18365,N_10374,N_14422);
or U18366 (N_18366,N_10053,N_11894);
nand U18367 (N_18367,N_14518,N_10054);
and U18368 (N_18368,N_10406,N_13546);
and U18369 (N_18369,N_10874,N_14382);
or U18370 (N_18370,N_14259,N_12064);
and U18371 (N_18371,N_14358,N_11096);
or U18372 (N_18372,N_11346,N_14635);
and U18373 (N_18373,N_14040,N_10517);
nand U18374 (N_18374,N_13334,N_11217);
nor U18375 (N_18375,N_13215,N_13499);
xor U18376 (N_18376,N_13835,N_12297);
xnor U18377 (N_18377,N_11836,N_13884);
nor U18378 (N_18378,N_14079,N_14520);
and U18379 (N_18379,N_11072,N_13916);
xnor U18380 (N_18380,N_14596,N_13177);
nor U18381 (N_18381,N_13186,N_10034);
nor U18382 (N_18382,N_10076,N_12185);
nand U18383 (N_18383,N_14877,N_10037);
nor U18384 (N_18384,N_10604,N_11483);
or U18385 (N_18385,N_14470,N_12947);
or U18386 (N_18386,N_14159,N_10342);
nor U18387 (N_18387,N_13331,N_10840);
nor U18388 (N_18388,N_11803,N_12734);
or U18389 (N_18389,N_10891,N_12848);
and U18390 (N_18390,N_13318,N_13778);
nor U18391 (N_18391,N_12431,N_12566);
xnor U18392 (N_18392,N_12664,N_12867);
nand U18393 (N_18393,N_14158,N_10041);
xor U18394 (N_18394,N_12125,N_13052);
nor U18395 (N_18395,N_12562,N_12591);
xnor U18396 (N_18396,N_13018,N_10094);
nor U18397 (N_18397,N_10321,N_12663);
and U18398 (N_18398,N_10931,N_10299);
or U18399 (N_18399,N_10179,N_12850);
nor U18400 (N_18400,N_13935,N_10958);
and U18401 (N_18401,N_11413,N_10918);
nor U18402 (N_18402,N_10793,N_13667);
or U18403 (N_18403,N_13300,N_10712);
or U18404 (N_18404,N_13826,N_13527);
nor U18405 (N_18405,N_10887,N_10662);
and U18406 (N_18406,N_13920,N_12205);
xnor U18407 (N_18407,N_12962,N_11381);
nand U18408 (N_18408,N_10414,N_13210);
or U18409 (N_18409,N_13229,N_13647);
or U18410 (N_18410,N_14737,N_10591);
or U18411 (N_18411,N_10742,N_14080);
and U18412 (N_18412,N_12375,N_10593);
xnor U18413 (N_18413,N_13281,N_11846);
nor U18414 (N_18414,N_10019,N_12729);
xnor U18415 (N_18415,N_13259,N_12659);
or U18416 (N_18416,N_12095,N_14782);
or U18417 (N_18417,N_12766,N_13726);
and U18418 (N_18418,N_11335,N_11223);
or U18419 (N_18419,N_11534,N_10173);
nand U18420 (N_18420,N_12308,N_10411);
and U18421 (N_18421,N_11222,N_13273);
and U18422 (N_18422,N_13960,N_14660);
nor U18423 (N_18423,N_10759,N_12315);
nand U18424 (N_18424,N_13661,N_10079);
nor U18425 (N_18425,N_14074,N_10585);
nor U18426 (N_18426,N_12599,N_10364);
and U18427 (N_18427,N_10386,N_13203);
nand U18428 (N_18428,N_13746,N_14175);
nand U18429 (N_18429,N_12844,N_10052);
or U18430 (N_18430,N_11216,N_12815);
or U18431 (N_18431,N_10952,N_12485);
nand U18432 (N_18432,N_12396,N_12282);
nand U18433 (N_18433,N_11353,N_14673);
nor U18434 (N_18434,N_13655,N_11192);
nor U18435 (N_18435,N_12302,N_11347);
nor U18436 (N_18436,N_10128,N_12876);
nand U18437 (N_18437,N_14590,N_14084);
nor U18438 (N_18438,N_11006,N_13726);
and U18439 (N_18439,N_11209,N_13805);
and U18440 (N_18440,N_12067,N_12829);
nor U18441 (N_18441,N_10159,N_13950);
or U18442 (N_18442,N_10526,N_14549);
nor U18443 (N_18443,N_13736,N_14120);
and U18444 (N_18444,N_13625,N_10726);
nor U18445 (N_18445,N_12676,N_10726);
nor U18446 (N_18446,N_14183,N_10794);
nand U18447 (N_18447,N_13810,N_11631);
or U18448 (N_18448,N_10276,N_11212);
nand U18449 (N_18449,N_13778,N_10067);
nand U18450 (N_18450,N_11595,N_14258);
nor U18451 (N_18451,N_12505,N_11170);
or U18452 (N_18452,N_12960,N_10107);
nor U18453 (N_18453,N_13976,N_10936);
or U18454 (N_18454,N_10419,N_13669);
and U18455 (N_18455,N_14783,N_11027);
nand U18456 (N_18456,N_10586,N_12698);
or U18457 (N_18457,N_10665,N_10021);
nor U18458 (N_18458,N_10985,N_13088);
nor U18459 (N_18459,N_10627,N_10622);
or U18460 (N_18460,N_14166,N_13002);
nand U18461 (N_18461,N_11215,N_10613);
nand U18462 (N_18462,N_13789,N_14039);
or U18463 (N_18463,N_14591,N_12227);
nand U18464 (N_18464,N_10759,N_13324);
and U18465 (N_18465,N_11505,N_12671);
nand U18466 (N_18466,N_14936,N_11276);
and U18467 (N_18467,N_13079,N_10634);
nor U18468 (N_18468,N_13102,N_10260);
and U18469 (N_18469,N_10111,N_10613);
or U18470 (N_18470,N_10782,N_13680);
or U18471 (N_18471,N_13828,N_10181);
nor U18472 (N_18472,N_11058,N_10558);
nand U18473 (N_18473,N_11086,N_14994);
or U18474 (N_18474,N_10892,N_13206);
and U18475 (N_18475,N_10894,N_14669);
nand U18476 (N_18476,N_14015,N_14270);
and U18477 (N_18477,N_14726,N_12372);
nand U18478 (N_18478,N_14473,N_13422);
or U18479 (N_18479,N_13166,N_13970);
nand U18480 (N_18480,N_12609,N_11128);
nor U18481 (N_18481,N_11157,N_11164);
and U18482 (N_18482,N_10435,N_11098);
nand U18483 (N_18483,N_13043,N_13804);
and U18484 (N_18484,N_12214,N_11398);
nand U18485 (N_18485,N_10682,N_11812);
nand U18486 (N_18486,N_12779,N_12768);
xor U18487 (N_18487,N_14350,N_13260);
and U18488 (N_18488,N_13888,N_10133);
xnor U18489 (N_18489,N_14696,N_12682);
nor U18490 (N_18490,N_14826,N_14304);
or U18491 (N_18491,N_11547,N_11786);
nand U18492 (N_18492,N_12697,N_12986);
nand U18493 (N_18493,N_12713,N_13058);
and U18494 (N_18494,N_10617,N_11607);
or U18495 (N_18495,N_12434,N_10527);
and U18496 (N_18496,N_13007,N_12368);
or U18497 (N_18497,N_11833,N_14030);
or U18498 (N_18498,N_14078,N_13925);
or U18499 (N_18499,N_12698,N_11532);
nor U18500 (N_18500,N_14027,N_14976);
nand U18501 (N_18501,N_13866,N_10380);
nor U18502 (N_18502,N_10637,N_11541);
nand U18503 (N_18503,N_13348,N_12611);
nand U18504 (N_18504,N_10029,N_14880);
nor U18505 (N_18505,N_14168,N_11480);
or U18506 (N_18506,N_14771,N_10943);
xnor U18507 (N_18507,N_11888,N_14340);
nor U18508 (N_18508,N_10580,N_11292);
nor U18509 (N_18509,N_10288,N_10859);
nand U18510 (N_18510,N_12767,N_11909);
nor U18511 (N_18511,N_10426,N_14183);
and U18512 (N_18512,N_13237,N_12125);
and U18513 (N_18513,N_13584,N_11676);
nor U18514 (N_18514,N_13028,N_11703);
and U18515 (N_18515,N_13196,N_11784);
and U18516 (N_18516,N_13117,N_14712);
and U18517 (N_18517,N_12552,N_13012);
or U18518 (N_18518,N_14395,N_10591);
nor U18519 (N_18519,N_10158,N_11241);
xnor U18520 (N_18520,N_11801,N_13409);
nor U18521 (N_18521,N_11073,N_11866);
nand U18522 (N_18522,N_13100,N_14507);
and U18523 (N_18523,N_10785,N_14090);
and U18524 (N_18524,N_11809,N_13082);
or U18525 (N_18525,N_14712,N_13504);
nor U18526 (N_18526,N_12794,N_14683);
nand U18527 (N_18527,N_13616,N_12811);
nand U18528 (N_18528,N_13894,N_10406);
nor U18529 (N_18529,N_13173,N_10310);
nand U18530 (N_18530,N_12356,N_13796);
nand U18531 (N_18531,N_10360,N_14789);
and U18532 (N_18532,N_14146,N_10558);
xor U18533 (N_18533,N_10750,N_14923);
and U18534 (N_18534,N_12747,N_12245);
xnor U18535 (N_18535,N_10475,N_14433);
and U18536 (N_18536,N_13633,N_13608);
or U18537 (N_18537,N_13326,N_13313);
nand U18538 (N_18538,N_14475,N_11482);
nor U18539 (N_18539,N_11819,N_13436);
nand U18540 (N_18540,N_12582,N_10815);
nor U18541 (N_18541,N_12604,N_12066);
xnor U18542 (N_18542,N_13247,N_12639);
or U18543 (N_18543,N_11745,N_10815);
or U18544 (N_18544,N_10633,N_12979);
nand U18545 (N_18545,N_12387,N_12455);
xor U18546 (N_18546,N_11279,N_11566);
nor U18547 (N_18547,N_10628,N_12031);
nor U18548 (N_18548,N_14886,N_11079);
and U18549 (N_18549,N_12780,N_12727);
nand U18550 (N_18550,N_13011,N_11058);
nor U18551 (N_18551,N_12577,N_13749);
and U18552 (N_18552,N_10166,N_13777);
or U18553 (N_18553,N_11693,N_12521);
nor U18554 (N_18554,N_13172,N_12018);
nor U18555 (N_18555,N_13074,N_12204);
nor U18556 (N_18556,N_11918,N_11443);
nor U18557 (N_18557,N_10036,N_12748);
or U18558 (N_18558,N_14074,N_10531);
or U18559 (N_18559,N_14245,N_13889);
and U18560 (N_18560,N_11434,N_10616);
and U18561 (N_18561,N_12478,N_12127);
nor U18562 (N_18562,N_11910,N_11382);
nor U18563 (N_18563,N_12908,N_14948);
or U18564 (N_18564,N_11658,N_11516);
and U18565 (N_18565,N_10976,N_13581);
nand U18566 (N_18566,N_11283,N_10732);
and U18567 (N_18567,N_11202,N_14013);
nor U18568 (N_18568,N_14847,N_13277);
nand U18569 (N_18569,N_11735,N_14262);
nor U18570 (N_18570,N_14041,N_13922);
and U18571 (N_18571,N_13109,N_12064);
nand U18572 (N_18572,N_11576,N_10710);
and U18573 (N_18573,N_10626,N_10384);
and U18574 (N_18574,N_13339,N_11275);
and U18575 (N_18575,N_10602,N_10772);
and U18576 (N_18576,N_14204,N_12803);
nor U18577 (N_18577,N_11694,N_10033);
xnor U18578 (N_18578,N_10855,N_12910);
and U18579 (N_18579,N_14394,N_13295);
and U18580 (N_18580,N_13672,N_12488);
nand U18581 (N_18581,N_11983,N_14459);
xor U18582 (N_18582,N_12075,N_13113);
or U18583 (N_18583,N_13429,N_11035);
and U18584 (N_18584,N_10895,N_10682);
or U18585 (N_18585,N_10100,N_11798);
and U18586 (N_18586,N_14715,N_10328);
and U18587 (N_18587,N_14058,N_11909);
nor U18588 (N_18588,N_12663,N_14068);
nand U18589 (N_18589,N_12407,N_11300);
xnor U18590 (N_18590,N_10810,N_12690);
nor U18591 (N_18591,N_14843,N_11669);
or U18592 (N_18592,N_10676,N_11925);
nand U18593 (N_18593,N_13670,N_14760);
and U18594 (N_18594,N_14274,N_14715);
and U18595 (N_18595,N_14864,N_10515);
or U18596 (N_18596,N_13110,N_14580);
and U18597 (N_18597,N_10204,N_14009);
nand U18598 (N_18598,N_14357,N_14290);
xnor U18599 (N_18599,N_10449,N_10855);
and U18600 (N_18600,N_10742,N_11238);
nand U18601 (N_18601,N_12690,N_10557);
nor U18602 (N_18602,N_10378,N_14470);
and U18603 (N_18603,N_12113,N_11644);
nand U18604 (N_18604,N_10711,N_12045);
nor U18605 (N_18605,N_12819,N_12016);
nand U18606 (N_18606,N_10034,N_13453);
nand U18607 (N_18607,N_10222,N_13769);
and U18608 (N_18608,N_10616,N_11728);
nand U18609 (N_18609,N_10634,N_10834);
or U18610 (N_18610,N_10117,N_12777);
nand U18611 (N_18611,N_14036,N_12829);
nand U18612 (N_18612,N_14646,N_10860);
and U18613 (N_18613,N_10846,N_12380);
nor U18614 (N_18614,N_13804,N_11418);
and U18615 (N_18615,N_14769,N_14781);
nor U18616 (N_18616,N_14873,N_14439);
nand U18617 (N_18617,N_12620,N_13160);
or U18618 (N_18618,N_13600,N_12692);
nor U18619 (N_18619,N_10162,N_14750);
or U18620 (N_18620,N_12793,N_12146);
xnor U18621 (N_18621,N_12889,N_11561);
and U18622 (N_18622,N_12282,N_13108);
nand U18623 (N_18623,N_12228,N_14945);
and U18624 (N_18624,N_13618,N_10938);
nor U18625 (N_18625,N_13659,N_11176);
and U18626 (N_18626,N_12275,N_14393);
nand U18627 (N_18627,N_10614,N_13815);
and U18628 (N_18628,N_12611,N_14121);
xor U18629 (N_18629,N_10197,N_12403);
and U18630 (N_18630,N_14012,N_11123);
nand U18631 (N_18631,N_10358,N_14074);
or U18632 (N_18632,N_13061,N_14384);
nand U18633 (N_18633,N_10053,N_12630);
nand U18634 (N_18634,N_11768,N_12367);
or U18635 (N_18635,N_14530,N_13795);
and U18636 (N_18636,N_10462,N_13043);
nor U18637 (N_18637,N_14131,N_11602);
and U18638 (N_18638,N_11884,N_14312);
nor U18639 (N_18639,N_14038,N_13141);
and U18640 (N_18640,N_10333,N_13852);
and U18641 (N_18641,N_11503,N_12565);
and U18642 (N_18642,N_14192,N_10684);
or U18643 (N_18643,N_11682,N_12593);
or U18644 (N_18644,N_13783,N_13506);
and U18645 (N_18645,N_10112,N_14091);
nor U18646 (N_18646,N_12540,N_13157);
and U18647 (N_18647,N_12405,N_11230);
nand U18648 (N_18648,N_12188,N_14225);
and U18649 (N_18649,N_11745,N_12415);
and U18650 (N_18650,N_10160,N_11465);
nand U18651 (N_18651,N_10659,N_12435);
nor U18652 (N_18652,N_11976,N_12703);
or U18653 (N_18653,N_10173,N_14486);
nand U18654 (N_18654,N_11562,N_13469);
or U18655 (N_18655,N_12658,N_14190);
and U18656 (N_18656,N_10013,N_14393);
or U18657 (N_18657,N_12118,N_12186);
and U18658 (N_18658,N_12322,N_14047);
and U18659 (N_18659,N_11857,N_12664);
nor U18660 (N_18660,N_14966,N_11565);
nor U18661 (N_18661,N_13287,N_10488);
and U18662 (N_18662,N_13543,N_13953);
or U18663 (N_18663,N_13141,N_14326);
or U18664 (N_18664,N_14638,N_13206);
xor U18665 (N_18665,N_11825,N_14439);
or U18666 (N_18666,N_14293,N_13509);
and U18667 (N_18667,N_11190,N_12561);
nor U18668 (N_18668,N_10798,N_14753);
nand U18669 (N_18669,N_14048,N_10913);
nor U18670 (N_18670,N_13514,N_12843);
or U18671 (N_18671,N_13611,N_12433);
and U18672 (N_18672,N_10671,N_10737);
or U18673 (N_18673,N_12931,N_11307);
xnor U18674 (N_18674,N_13790,N_12874);
or U18675 (N_18675,N_13643,N_13998);
and U18676 (N_18676,N_10607,N_13481);
and U18677 (N_18677,N_14992,N_12524);
xor U18678 (N_18678,N_10339,N_10835);
or U18679 (N_18679,N_10611,N_14709);
nand U18680 (N_18680,N_10922,N_14656);
nor U18681 (N_18681,N_12388,N_11587);
or U18682 (N_18682,N_11698,N_14606);
nor U18683 (N_18683,N_10835,N_11160);
nand U18684 (N_18684,N_12955,N_11755);
and U18685 (N_18685,N_13992,N_12019);
nand U18686 (N_18686,N_11609,N_10595);
xnor U18687 (N_18687,N_12741,N_12298);
nand U18688 (N_18688,N_13805,N_14938);
and U18689 (N_18689,N_12091,N_11874);
and U18690 (N_18690,N_10838,N_13815);
nor U18691 (N_18691,N_12535,N_12588);
and U18692 (N_18692,N_10980,N_11329);
and U18693 (N_18693,N_12409,N_12427);
and U18694 (N_18694,N_10543,N_12383);
nand U18695 (N_18695,N_10465,N_12808);
or U18696 (N_18696,N_10897,N_11969);
or U18697 (N_18697,N_10883,N_13171);
nor U18698 (N_18698,N_13304,N_14916);
or U18699 (N_18699,N_10129,N_11461);
nand U18700 (N_18700,N_13625,N_13661);
or U18701 (N_18701,N_11173,N_10018);
nand U18702 (N_18702,N_12522,N_11893);
nor U18703 (N_18703,N_13052,N_12457);
nand U18704 (N_18704,N_12932,N_13602);
xor U18705 (N_18705,N_11964,N_10881);
nor U18706 (N_18706,N_14836,N_14358);
and U18707 (N_18707,N_10116,N_12005);
and U18708 (N_18708,N_10802,N_11923);
nor U18709 (N_18709,N_11103,N_11752);
xnor U18710 (N_18710,N_12478,N_10868);
nand U18711 (N_18711,N_13751,N_11227);
and U18712 (N_18712,N_10417,N_11840);
or U18713 (N_18713,N_10929,N_13606);
or U18714 (N_18714,N_12497,N_13194);
and U18715 (N_18715,N_10344,N_13567);
and U18716 (N_18716,N_12342,N_12281);
xor U18717 (N_18717,N_11495,N_14870);
or U18718 (N_18718,N_10247,N_10931);
nor U18719 (N_18719,N_13994,N_12568);
nor U18720 (N_18720,N_11750,N_12075);
nor U18721 (N_18721,N_11480,N_11134);
or U18722 (N_18722,N_14555,N_10804);
and U18723 (N_18723,N_13855,N_12525);
and U18724 (N_18724,N_14712,N_13262);
nor U18725 (N_18725,N_11335,N_10510);
or U18726 (N_18726,N_14358,N_14775);
nand U18727 (N_18727,N_11686,N_12919);
nor U18728 (N_18728,N_11476,N_12453);
xnor U18729 (N_18729,N_12020,N_11225);
nand U18730 (N_18730,N_11706,N_13649);
or U18731 (N_18731,N_11695,N_12963);
nor U18732 (N_18732,N_12295,N_14681);
nand U18733 (N_18733,N_12148,N_11504);
and U18734 (N_18734,N_11825,N_11313);
and U18735 (N_18735,N_13447,N_13357);
nand U18736 (N_18736,N_11881,N_14887);
nand U18737 (N_18737,N_11077,N_12819);
nor U18738 (N_18738,N_12686,N_14994);
xnor U18739 (N_18739,N_12547,N_13427);
nand U18740 (N_18740,N_10440,N_13646);
xor U18741 (N_18741,N_12250,N_11764);
or U18742 (N_18742,N_12297,N_14847);
and U18743 (N_18743,N_11142,N_10807);
and U18744 (N_18744,N_13828,N_11154);
and U18745 (N_18745,N_12348,N_11672);
nand U18746 (N_18746,N_10818,N_12357);
or U18747 (N_18747,N_14911,N_14703);
nor U18748 (N_18748,N_13216,N_12635);
or U18749 (N_18749,N_14917,N_10388);
nor U18750 (N_18750,N_11563,N_10063);
or U18751 (N_18751,N_13981,N_10937);
or U18752 (N_18752,N_14606,N_13665);
xor U18753 (N_18753,N_13754,N_11756);
nor U18754 (N_18754,N_14321,N_12008);
xor U18755 (N_18755,N_11729,N_12430);
nor U18756 (N_18756,N_13517,N_11135);
nor U18757 (N_18757,N_10567,N_10193);
and U18758 (N_18758,N_14527,N_11401);
nand U18759 (N_18759,N_10487,N_10462);
or U18760 (N_18760,N_10094,N_13313);
nand U18761 (N_18761,N_11528,N_14520);
nand U18762 (N_18762,N_11299,N_11903);
nand U18763 (N_18763,N_11259,N_12184);
xor U18764 (N_18764,N_13401,N_12436);
or U18765 (N_18765,N_10523,N_13214);
or U18766 (N_18766,N_14446,N_14704);
nor U18767 (N_18767,N_10868,N_14337);
or U18768 (N_18768,N_10390,N_14653);
or U18769 (N_18769,N_10290,N_12713);
nor U18770 (N_18770,N_11656,N_11673);
nor U18771 (N_18771,N_13759,N_10093);
nor U18772 (N_18772,N_14677,N_12653);
or U18773 (N_18773,N_11571,N_13446);
or U18774 (N_18774,N_10408,N_10461);
and U18775 (N_18775,N_12837,N_10899);
or U18776 (N_18776,N_10297,N_10906);
nor U18777 (N_18777,N_13064,N_10997);
and U18778 (N_18778,N_11086,N_12440);
nor U18779 (N_18779,N_12719,N_14560);
and U18780 (N_18780,N_11984,N_10245);
nand U18781 (N_18781,N_11375,N_14224);
nand U18782 (N_18782,N_10552,N_14719);
nand U18783 (N_18783,N_11206,N_12677);
nor U18784 (N_18784,N_14854,N_12123);
or U18785 (N_18785,N_11971,N_11748);
nor U18786 (N_18786,N_12662,N_12658);
and U18787 (N_18787,N_14996,N_11761);
nor U18788 (N_18788,N_11179,N_12415);
xnor U18789 (N_18789,N_13699,N_12258);
or U18790 (N_18790,N_12116,N_14344);
xnor U18791 (N_18791,N_10609,N_12637);
nand U18792 (N_18792,N_14010,N_14283);
nor U18793 (N_18793,N_14662,N_11338);
xor U18794 (N_18794,N_13708,N_11477);
or U18795 (N_18795,N_14931,N_11321);
nand U18796 (N_18796,N_10811,N_12463);
nand U18797 (N_18797,N_14120,N_10596);
and U18798 (N_18798,N_13164,N_14164);
nor U18799 (N_18799,N_14914,N_14987);
nor U18800 (N_18800,N_11117,N_14844);
nor U18801 (N_18801,N_11451,N_10984);
nor U18802 (N_18802,N_12652,N_11165);
or U18803 (N_18803,N_12515,N_11895);
nor U18804 (N_18804,N_14453,N_11242);
and U18805 (N_18805,N_13035,N_14014);
or U18806 (N_18806,N_12181,N_11443);
nand U18807 (N_18807,N_14309,N_12906);
nand U18808 (N_18808,N_13491,N_13906);
and U18809 (N_18809,N_10166,N_11312);
nor U18810 (N_18810,N_12201,N_12649);
nand U18811 (N_18811,N_12331,N_14394);
or U18812 (N_18812,N_14837,N_14745);
and U18813 (N_18813,N_14514,N_12287);
nand U18814 (N_18814,N_12152,N_10729);
or U18815 (N_18815,N_10741,N_12047);
nor U18816 (N_18816,N_14003,N_14382);
and U18817 (N_18817,N_14869,N_12413);
or U18818 (N_18818,N_14507,N_13329);
and U18819 (N_18819,N_10118,N_13238);
and U18820 (N_18820,N_12056,N_12899);
nand U18821 (N_18821,N_10085,N_12317);
or U18822 (N_18822,N_11944,N_11393);
nand U18823 (N_18823,N_14197,N_13206);
nand U18824 (N_18824,N_10655,N_12647);
and U18825 (N_18825,N_10475,N_12519);
nand U18826 (N_18826,N_11365,N_10598);
or U18827 (N_18827,N_10884,N_14674);
or U18828 (N_18828,N_11500,N_14817);
and U18829 (N_18829,N_13438,N_10785);
nand U18830 (N_18830,N_10169,N_11327);
xor U18831 (N_18831,N_10659,N_13160);
nand U18832 (N_18832,N_12227,N_13363);
and U18833 (N_18833,N_12517,N_14332);
or U18834 (N_18834,N_10013,N_10007);
and U18835 (N_18835,N_11701,N_11174);
xnor U18836 (N_18836,N_13860,N_12717);
nor U18837 (N_18837,N_13996,N_13419);
nor U18838 (N_18838,N_14400,N_14519);
nor U18839 (N_18839,N_10346,N_14021);
nand U18840 (N_18840,N_11019,N_10034);
nand U18841 (N_18841,N_11475,N_12097);
and U18842 (N_18842,N_10360,N_10682);
nand U18843 (N_18843,N_11180,N_12543);
xnor U18844 (N_18844,N_10854,N_10087);
xor U18845 (N_18845,N_14810,N_10957);
nand U18846 (N_18846,N_10278,N_12873);
nor U18847 (N_18847,N_10146,N_10992);
xnor U18848 (N_18848,N_14145,N_12676);
nand U18849 (N_18849,N_11038,N_12576);
or U18850 (N_18850,N_11102,N_12485);
nand U18851 (N_18851,N_14172,N_13046);
xor U18852 (N_18852,N_13945,N_10799);
or U18853 (N_18853,N_13733,N_14785);
nand U18854 (N_18854,N_13813,N_10047);
or U18855 (N_18855,N_10257,N_14580);
nand U18856 (N_18856,N_13489,N_11440);
nand U18857 (N_18857,N_11400,N_12641);
or U18858 (N_18858,N_10557,N_10751);
and U18859 (N_18859,N_14468,N_10599);
nand U18860 (N_18860,N_12861,N_11909);
nand U18861 (N_18861,N_14913,N_10048);
and U18862 (N_18862,N_13886,N_12938);
nor U18863 (N_18863,N_13275,N_11552);
nor U18864 (N_18864,N_10496,N_14852);
or U18865 (N_18865,N_13338,N_13350);
or U18866 (N_18866,N_12630,N_13689);
nor U18867 (N_18867,N_12090,N_12529);
and U18868 (N_18868,N_14583,N_10286);
xor U18869 (N_18869,N_11555,N_10716);
and U18870 (N_18870,N_13384,N_10522);
nand U18871 (N_18871,N_12785,N_14178);
nor U18872 (N_18872,N_11156,N_12236);
nor U18873 (N_18873,N_14039,N_13917);
nor U18874 (N_18874,N_11150,N_12041);
nand U18875 (N_18875,N_11068,N_12859);
nand U18876 (N_18876,N_11881,N_12572);
nor U18877 (N_18877,N_14555,N_14823);
nand U18878 (N_18878,N_11126,N_10311);
nor U18879 (N_18879,N_14686,N_13953);
xor U18880 (N_18880,N_11875,N_14097);
xnor U18881 (N_18881,N_11279,N_10723);
nand U18882 (N_18882,N_10162,N_11861);
nand U18883 (N_18883,N_11427,N_12915);
and U18884 (N_18884,N_14562,N_11267);
nand U18885 (N_18885,N_12784,N_14619);
nand U18886 (N_18886,N_11962,N_10007);
nor U18887 (N_18887,N_10173,N_12403);
nand U18888 (N_18888,N_14210,N_13307);
xor U18889 (N_18889,N_10195,N_12895);
or U18890 (N_18890,N_13270,N_12512);
or U18891 (N_18891,N_10561,N_13367);
xor U18892 (N_18892,N_11125,N_10962);
or U18893 (N_18893,N_11731,N_10963);
and U18894 (N_18894,N_10391,N_11812);
nand U18895 (N_18895,N_13754,N_13976);
nor U18896 (N_18896,N_13872,N_11647);
nor U18897 (N_18897,N_10585,N_11710);
and U18898 (N_18898,N_13407,N_11181);
and U18899 (N_18899,N_11626,N_11309);
or U18900 (N_18900,N_11997,N_10781);
xnor U18901 (N_18901,N_10425,N_12649);
nand U18902 (N_18902,N_13787,N_14402);
and U18903 (N_18903,N_14697,N_13939);
nor U18904 (N_18904,N_10954,N_13384);
nor U18905 (N_18905,N_12599,N_11562);
nor U18906 (N_18906,N_10390,N_14806);
nor U18907 (N_18907,N_14050,N_14674);
nand U18908 (N_18908,N_13617,N_12804);
xnor U18909 (N_18909,N_11641,N_14626);
nand U18910 (N_18910,N_13804,N_10113);
or U18911 (N_18911,N_11269,N_13650);
and U18912 (N_18912,N_12947,N_13110);
nor U18913 (N_18913,N_14475,N_12675);
nand U18914 (N_18914,N_10091,N_12476);
nand U18915 (N_18915,N_14970,N_12735);
nand U18916 (N_18916,N_10899,N_13009);
nand U18917 (N_18917,N_13386,N_11320);
and U18918 (N_18918,N_10698,N_11457);
nand U18919 (N_18919,N_10811,N_13633);
nand U18920 (N_18920,N_12473,N_14802);
xnor U18921 (N_18921,N_12081,N_14443);
nand U18922 (N_18922,N_12774,N_12132);
nor U18923 (N_18923,N_12419,N_10999);
nor U18924 (N_18924,N_11850,N_11019);
nor U18925 (N_18925,N_14253,N_13320);
or U18926 (N_18926,N_12933,N_10562);
nand U18927 (N_18927,N_10679,N_14428);
and U18928 (N_18928,N_14451,N_13901);
and U18929 (N_18929,N_10688,N_10975);
and U18930 (N_18930,N_12513,N_10546);
or U18931 (N_18931,N_12063,N_14511);
nand U18932 (N_18932,N_11304,N_11831);
nor U18933 (N_18933,N_10164,N_10299);
nor U18934 (N_18934,N_11873,N_11067);
xor U18935 (N_18935,N_14389,N_14794);
nand U18936 (N_18936,N_11665,N_11334);
and U18937 (N_18937,N_14556,N_14343);
or U18938 (N_18938,N_10218,N_12654);
nand U18939 (N_18939,N_10110,N_13572);
nand U18940 (N_18940,N_10828,N_13311);
nand U18941 (N_18941,N_11598,N_14208);
and U18942 (N_18942,N_13574,N_10177);
nand U18943 (N_18943,N_14015,N_10944);
nand U18944 (N_18944,N_10381,N_13111);
and U18945 (N_18945,N_12688,N_10726);
or U18946 (N_18946,N_14270,N_12519);
nor U18947 (N_18947,N_11805,N_12111);
or U18948 (N_18948,N_11179,N_12450);
or U18949 (N_18949,N_14219,N_13952);
and U18950 (N_18950,N_12409,N_11982);
nand U18951 (N_18951,N_13151,N_12962);
or U18952 (N_18952,N_13535,N_11106);
xor U18953 (N_18953,N_13228,N_12391);
nor U18954 (N_18954,N_12330,N_13316);
or U18955 (N_18955,N_11470,N_13120);
and U18956 (N_18956,N_10760,N_12332);
or U18957 (N_18957,N_14706,N_11278);
and U18958 (N_18958,N_13147,N_14496);
nor U18959 (N_18959,N_11959,N_12200);
or U18960 (N_18960,N_11690,N_11298);
nand U18961 (N_18961,N_13364,N_10914);
nand U18962 (N_18962,N_14915,N_14605);
or U18963 (N_18963,N_11763,N_11417);
nor U18964 (N_18964,N_12032,N_11549);
or U18965 (N_18965,N_13120,N_13955);
and U18966 (N_18966,N_14899,N_10484);
and U18967 (N_18967,N_10317,N_14770);
or U18968 (N_18968,N_12057,N_14754);
or U18969 (N_18969,N_10893,N_14765);
and U18970 (N_18970,N_13476,N_11905);
nand U18971 (N_18971,N_11411,N_13137);
and U18972 (N_18972,N_10348,N_12761);
and U18973 (N_18973,N_12851,N_11916);
or U18974 (N_18974,N_12930,N_14830);
nor U18975 (N_18975,N_13857,N_11837);
nand U18976 (N_18976,N_13460,N_13897);
and U18977 (N_18977,N_14620,N_14164);
and U18978 (N_18978,N_14111,N_12584);
and U18979 (N_18979,N_12410,N_14818);
nor U18980 (N_18980,N_14926,N_14665);
xnor U18981 (N_18981,N_10100,N_13474);
xor U18982 (N_18982,N_13244,N_11796);
nor U18983 (N_18983,N_13892,N_11506);
or U18984 (N_18984,N_14746,N_12092);
xnor U18985 (N_18985,N_12180,N_13447);
or U18986 (N_18986,N_11908,N_11398);
nor U18987 (N_18987,N_10766,N_10633);
or U18988 (N_18988,N_12663,N_10612);
and U18989 (N_18989,N_13969,N_14886);
and U18990 (N_18990,N_14953,N_10742);
or U18991 (N_18991,N_13442,N_11016);
nor U18992 (N_18992,N_14435,N_14797);
or U18993 (N_18993,N_10879,N_10083);
or U18994 (N_18994,N_14844,N_13168);
nor U18995 (N_18995,N_14965,N_10191);
or U18996 (N_18996,N_14553,N_10762);
nand U18997 (N_18997,N_10308,N_12448);
and U18998 (N_18998,N_12935,N_12612);
or U18999 (N_18999,N_12869,N_12802);
nand U19000 (N_19000,N_11496,N_13517);
or U19001 (N_19001,N_11484,N_11062);
xor U19002 (N_19002,N_10725,N_11288);
nand U19003 (N_19003,N_12379,N_14385);
nand U19004 (N_19004,N_11925,N_11050);
nor U19005 (N_19005,N_14648,N_14536);
xor U19006 (N_19006,N_10576,N_14946);
or U19007 (N_19007,N_13134,N_13251);
nor U19008 (N_19008,N_13904,N_11537);
nor U19009 (N_19009,N_10935,N_12933);
nor U19010 (N_19010,N_12184,N_10553);
nand U19011 (N_19011,N_13996,N_11291);
nand U19012 (N_19012,N_12760,N_13192);
or U19013 (N_19013,N_13992,N_10909);
nand U19014 (N_19014,N_11983,N_13814);
nor U19015 (N_19015,N_14487,N_12566);
nor U19016 (N_19016,N_10426,N_12503);
or U19017 (N_19017,N_13448,N_10325);
nor U19018 (N_19018,N_11303,N_12119);
and U19019 (N_19019,N_14771,N_10049);
or U19020 (N_19020,N_13710,N_13001);
and U19021 (N_19021,N_14527,N_10703);
and U19022 (N_19022,N_11196,N_10132);
nor U19023 (N_19023,N_13652,N_10182);
xnor U19024 (N_19024,N_13987,N_14522);
or U19025 (N_19025,N_13312,N_12814);
and U19026 (N_19026,N_13644,N_14410);
or U19027 (N_19027,N_11654,N_14774);
nand U19028 (N_19028,N_11294,N_11915);
or U19029 (N_19029,N_10947,N_11051);
xnor U19030 (N_19030,N_14140,N_13128);
nand U19031 (N_19031,N_14219,N_11306);
nand U19032 (N_19032,N_13110,N_12664);
or U19033 (N_19033,N_10250,N_10218);
nand U19034 (N_19034,N_13414,N_12759);
nand U19035 (N_19035,N_10098,N_13700);
nand U19036 (N_19036,N_13126,N_10089);
and U19037 (N_19037,N_11298,N_12476);
nor U19038 (N_19038,N_14972,N_10594);
or U19039 (N_19039,N_11790,N_14973);
nor U19040 (N_19040,N_12005,N_11198);
and U19041 (N_19041,N_12785,N_14802);
nor U19042 (N_19042,N_10041,N_12262);
and U19043 (N_19043,N_14612,N_12360);
or U19044 (N_19044,N_14541,N_14375);
nor U19045 (N_19045,N_13112,N_12586);
or U19046 (N_19046,N_12138,N_10844);
or U19047 (N_19047,N_12761,N_13712);
nor U19048 (N_19048,N_10448,N_11544);
nor U19049 (N_19049,N_12756,N_14911);
nand U19050 (N_19050,N_13973,N_13444);
or U19051 (N_19051,N_11106,N_11790);
nand U19052 (N_19052,N_12070,N_13763);
nand U19053 (N_19053,N_11662,N_13058);
and U19054 (N_19054,N_11001,N_14712);
nor U19055 (N_19055,N_14182,N_10796);
xor U19056 (N_19056,N_13847,N_13281);
xnor U19057 (N_19057,N_11209,N_13827);
nand U19058 (N_19058,N_12829,N_10027);
nand U19059 (N_19059,N_14880,N_13814);
and U19060 (N_19060,N_10681,N_11191);
nor U19061 (N_19061,N_11178,N_10367);
nor U19062 (N_19062,N_10341,N_14909);
or U19063 (N_19063,N_12067,N_14202);
or U19064 (N_19064,N_14479,N_13970);
xor U19065 (N_19065,N_11198,N_11498);
nand U19066 (N_19066,N_12411,N_13834);
nand U19067 (N_19067,N_13719,N_13189);
and U19068 (N_19068,N_10556,N_13291);
or U19069 (N_19069,N_13825,N_14536);
nand U19070 (N_19070,N_10170,N_14816);
nor U19071 (N_19071,N_12174,N_13162);
or U19072 (N_19072,N_12157,N_12310);
nand U19073 (N_19073,N_12358,N_14463);
nor U19074 (N_19074,N_12941,N_12967);
and U19075 (N_19075,N_13262,N_12484);
and U19076 (N_19076,N_13383,N_11490);
xnor U19077 (N_19077,N_14026,N_13695);
nor U19078 (N_19078,N_10296,N_12609);
nand U19079 (N_19079,N_10131,N_10042);
nand U19080 (N_19080,N_13417,N_13890);
and U19081 (N_19081,N_14690,N_12345);
and U19082 (N_19082,N_11483,N_14737);
nand U19083 (N_19083,N_13967,N_10743);
and U19084 (N_19084,N_13571,N_13232);
and U19085 (N_19085,N_13454,N_11418);
nor U19086 (N_19086,N_10472,N_11282);
nor U19087 (N_19087,N_13338,N_12980);
and U19088 (N_19088,N_10998,N_12022);
nand U19089 (N_19089,N_12540,N_13837);
and U19090 (N_19090,N_13250,N_12619);
nor U19091 (N_19091,N_11709,N_14877);
xor U19092 (N_19092,N_10188,N_13544);
nand U19093 (N_19093,N_14806,N_10925);
nor U19094 (N_19094,N_10952,N_11360);
or U19095 (N_19095,N_13467,N_13516);
and U19096 (N_19096,N_11358,N_12887);
nor U19097 (N_19097,N_11853,N_13092);
or U19098 (N_19098,N_13900,N_13279);
and U19099 (N_19099,N_12532,N_10117);
xor U19100 (N_19100,N_12928,N_12495);
xor U19101 (N_19101,N_10017,N_13588);
and U19102 (N_19102,N_11050,N_13429);
and U19103 (N_19103,N_13113,N_10524);
nor U19104 (N_19104,N_13139,N_11274);
nor U19105 (N_19105,N_11419,N_11360);
nand U19106 (N_19106,N_10677,N_14141);
nor U19107 (N_19107,N_11498,N_14930);
or U19108 (N_19108,N_12787,N_12983);
nor U19109 (N_19109,N_10338,N_14245);
xnor U19110 (N_19110,N_14648,N_14892);
nor U19111 (N_19111,N_13408,N_10448);
nand U19112 (N_19112,N_13022,N_10735);
or U19113 (N_19113,N_13591,N_13899);
or U19114 (N_19114,N_14872,N_11437);
nor U19115 (N_19115,N_14719,N_14878);
xnor U19116 (N_19116,N_13065,N_14776);
nor U19117 (N_19117,N_14615,N_10697);
and U19118 (N_19118,N_14235,N_14923);
and U19119 (N_19119,N_10525,N_10752);
xor U19120 (N_19120,N_14391,N_10815);
or U19121 (N_19121,N_12495,N_14408);
or U19122 (N_19122,N_12414,N_11587);
or U19123 (N_19123,N_12494,N_10058);
and U19124 (N_19124,N_11765,N_12961);
nor U19125 (N_19125,N_14485,N_10719);
nor U19126 (N_19126,N_10253,N_12227);
and U19127 (N_19127,N_12100,N_13913);
nand U19128 (N_19128,N_14949,N_12815);
nor U19129 (N_19129,N_14589,N_12437);
nor U19130 (N_19130,N_11646,N_14254);
nand U19131 (N_19131,N_14410,N_12352);
nand U19132 (N_19132,N_13950,N_13010);
nor U19133 (N_19133,N_14250,N_11123);
nand U19134 (N_19134,N_10952,N_13857);
or U19135 (N_19135,N_13774,N_13058);
and U19136 (N_19136,N_13767,N_11293);
nor U19137 (N_19137,N_13082,N_11652);
nand U19138 (N_19138,N_10540,N_11740);
nand U19139 (N_19139,N_13550,N_14470);
and U19140 (N_19140,N_10653,N_14616);
nor U19141 (N_19141,N_12118,N_14812);
nand U19142 (N_19142,N_14698,N_10567);
or U19143 (N_19143,N_10258,N_11365);
or U19144 (N_19144,N_13892,N_13439);
nand U19145 (N_19145,N_13739,N_13284);
nand U19146 (N_19146,N_12354,N_14041);
nand U19147 (N_19147,N_14440,N_14273);
nor U19148 (N_19148,N_11174,N_10372);
or U19149 (N_19149,N_13960,N_10340);
and U19150 (N_19150,N_14298,N_12374);
or U19151 (N_19151,N_12129,N_13871);
and U19152 (N_19152,N_14935,N_13017);
nor U19153 (N_19153,N_10187,N_14108);
nor U19154 (N_19154,N_12777,N_14649);
nand U19155 (N_19155,N_12213,N_14985);
nor U19156 (N_19156,N_13375,N_11651);
nand U19157 (N_19157,N_14781,N_10542);
or U19158 (N_19158,N_11082,N_11742);
or U19159 (N_19159,N_13981,N_12656);
nor U19160 (N_19160,N_10681,N_13252);
nor U19161 (N_19161,N_12772,N_11343);
and U19162 (N_19162,N_13021,N_13333);
and U19163 (N_19163,N_11377,N_14375);
and U19164 (N_19164,N_14417,N_14582);
or U19165 (N_19165,N_10197,N_11782);
and U19166 (N_19166,N_11475,N_11043);
xor U19167 (N_19167,N_14544,N_12311);
and U19168 (N_19168,N_10630,N_10755);
nand U19169 (N_19169,N_12710,N_13153);
nor U19170 (N_19170,N_10854,N_12797);
nor U19171 (N_19171,N_14895,N_14496);
nand U19172 (N_19172,N_11194,N_13076);
and U19173 (N_19173,N_14024,N_10355);
and U19174 (N_19174,N_11817,N_12090);
or U19175 (N_19175,N_10795,N_14639);
or U19176 (N_19176,N_11757,N_11088);
nor U19177 (N_19177,N_10198,N_14604);
or U19178 (N_19178,N_11742,N_12322);
or U19179 (N_19179,N_11335,N_14428);
nor U19180 (N_19180,N_11384,N_11928);
nor U19181 (N_19181,N_11106,N_13859);
nor U19182 (N_19182,N_12023,N_11634);
or U19183 (N_19183,N_13468,N_13083);
nand U19184 (N_19184,N_12632,N_12040);
nor U19185 (N_19185,N_13726,N_13401);
nand U19186 (N_19186,N_10098,N_13181);
and U19187 (N_19187,N_11437,N_14148);
and U19188 (N_19188,N_11790,N_10559);
and U19189 (N_19189,N_13144,N_14403);
and U19190 (N_19190,N_11502,N_10846);
or U19191 (N_19191,N_10820,N_10071);
and U19192 (N_19192,N_13307,N_14195);
or U19193 (N_19193,N_13064,N_11210);
nor U19194 (N_19194,N_10025,N_11442);
and U19195 (N_19195,N_13565,N_11804);
nand U19196 (N_19196,N_10715,N_13082);
nand U19197 (N_19197,N_10684,N_10669);
or U19198 (N_19198,N_14965,N_14599);
nor U19199 (N_19199,N_12497,N_14194);
or U19200 (N_19200,N_13317,N_11294);
and U19201 (N_19201,N_12258,N_11513);
xnor U19202 (N_19202,N_12992,N_14450);
xnor U19203 (N_19203,N_11803,N_14614);
xnor U19204 (N_19204,N_11082,N_12813);
or U19205 (N_19205,N_13201,N_10663);
or U19206 (N_19206,N_14706,N_11783);
nand U19207 (N_19207,N_13855,N_14744);
or U19208 (N_19208,N_11655,N_13365);
xor U19209 (N_19209,N_11326,N_10029);
and U19210 (N_19210,N_13838,N_12247);
nor U19211 (N_19211,N_12553,N_11277);
and U19212 (N_19212,N_11138,N_14621);
nor U19213 (N_19213,N_14679,N_14032);
or U19214 (N_19214,N_13781,N_12115);
xnor U19215 (N_19215,N_11978,N_13525);
or U19216 (N_19216,N_11991,N_12843);
nand U19217 (N_19217,N_10529,N_10349);
or U19218 (N_19218,N_13274,N_14252);
or U19219 (N_19219,N_10164,N_13679);
nand U19220 (N_19220,N_11268,N_11519);
or U19221 (N_19221,N_13827,N_12900);
nor U19222 (N_19222,N_13451,N_10250);
or U19223 (N_19223,N_10573,N_11175);
or U19224 (N_19224,N_10342,N_14153);
or U19225 (N_19225,N_12889,N_11492);
or U19226 (N_19226,N_11984,N_10923);
or U19227 (N_19227,N_10344,N_11191);
nor U19228 (N_19228,N_13981,N_12734);
nand U19229 (N_19229,N_10786,N_12562);
nor U19230 (N_19230,N_12793,N_10791);
nand U19231 (N_19231,N_10000,N_10918);
or U19232 (N_19232,N_12995,N_10507);
and U19233 (N_19233,N_11657,N_12585);
nor U19234 (N_19234,N_13230,N_10728);
nor U19235 (N_19235,N_13249,N_14276);
xnor U19236 (N_19236,N_13347,N_12024);
nand U19237 (N_19237,N_14591,N_14184);
or U19238 (N_19238,N_11741,N_13261);
nor U19239 (N_19239,N_14891,N_12976);
and U19240 (N_19240,N_12007,N_10107);
nand U19241 (N_19241,N_12262,N_10062);
or U19242 (N_19242,N_12825,N_11397);
nor U19243 (N_19243,N_14930,N_14810);
or U19244 (N_19244,N_10579,N_11959);
and U19245 (N_19245,N_13205,N_12518);
or U19246 (N_19246,N_11849,N_13749);
or U19247 (N_19247,N_10834,N_14803);
nor U19248 (N_19248,N_11629,N_14164);
nor U19249 (N_19249,N_13201,N_14649);
nor U19250 (N_19250,N_11676,N_12096);
or U19251 (N_19251,N_10648,N_13298);
nor U19252 (N_19252,N_14908,N_14082);
and U19253 (N_19253,N_10632,N_13622);
and U19254 (N_19254,N_13368,N_11166);
or U19255 (N_19255,N_13108,N_13305);
nor U19256 (N_19256,N_10119,N_13289);
or U19257 (N_19257,N_12178,N_12401);
nand U19258 (N_19258,N_14297,N_12445);
xor U19259 (N_19259,N_13838,N_13209);
nor U19260 (N_19260,N_10273,N_14450);
nand U19261 (N_19261,N_13079,N_11798);
nand U19262 (N_19262,N_14508,N_11709);
xnor U19263 (N_19263,N_14541,N_12818);
or U19264 (N_19264,N_11170,N_10376);
xnor U19265 (N_19265,N_10934,N_13265);
or U19266 (N_19266,N_14994,N_13891);
nand U19267 (N_19267,N_12994,N_11079);
or U19268 (N_19268,N_11612,N_14415);
nand U19269 (N_19269,N_14750,N_14754);
or U19270 (N_19270,N_14895,N_11503);
or U19271 (N_19271,N_10747,N_14996);
nand U19272 (N_19272,N_11658,N_10684);
and U19273 (N_19273,N_13449,N_13057);
and U19274 (N_19274,N_11305,N_12121);
nand U19275 (N_19275,N_10488,N_11547);
nand U19276 (N_19276,N_13820,N_11480);
nand U19277 (N_19277,N_14682,N_14066);
nor U19278 (N_19278,N_10548,N_14557);
nand U19279 (N_19279,N_13223,N_12751);
and U19280 (N_19280,N_12643,N_12880);
nand U19281 (N_19281,N_13099,N_10171);
nand U19282 (N_19282,N_10455,N_11908);
nand U19283 (N_19283,N_14347,N_11192);
and U19284 (N_19284,N_11668,N_10928);
nand U19285 (N_19285,N_11582,N_11957);
nand U19286 (N_19286,N_14211,N_14310);
nor U19287 (N_19287,N_13366,N_12278);
nand U19288 (N_19288,N_14292,N_13237);
nand U19289 (N_19289,N_13014,N_12903);
nor U19290 (N_19290,N_11081,N_14003);
xor U19291 (N_19291,N_11754,N_12969);
or U19292 (N_19292,N_13439,N_13617);
xnor U19293 (N_19293,N_14338,N_13959);
nand U19294 (N_19294,N_10669,N_13754);
and U19295 (N_19295,N_13873,N_13491);
nor U19296 (N_19296,N_11712,N_11515);
nor U19297 (N_19297,N_12762,N_12119);
and U19298 (N_19298,N_10144,N_12014);
nor U19299 (N_19299,N_10354,N_11235);
or U19300 (N_19300,N_14838,N_10480);
and U19301 (N_19301,N_10274,N_14544);
nor U19302 (N_19302,N_10177,N_10420);
nor U19303 (N_19303,N_13547,N_14535);
or U19304 (N_19304,N_10460,N_11122);
nand U19305 (N_19305,N_13767,N_11044);
and U19306 (N_19306,N_13283,N_14930);
and U19307 (N_19307,N_14926,N_14256);
nor U19308 (N_19308,N_12257,N_12379);
nand U19309 (N_19309,N_11397,N_11675);
and U19310 (N_19310,N_14275,N_11718);
or U19311 (N_19311,N_12327,N_11176);
nand U19312 (N_19312,N_11820,N_13121);
and U19313 (N_19313,N_10732,N_11999);
nor U19314 (N_19314,N_14362,N_10831);
xnor U19315 (N_19315,N_11688,N_10397);
and U19316 (N_19316,N_10292,N_12565);
nand U19317 (N_19317,N_14429,N_12718);
nand U19318 (N_19318,N_11972,N_11074);
or U19319 (N_19319,N_13652,N_11252);
nand U19320 (N_19320,N_10303,N_12871);
and U19321 (N_19321,N_10976,N_10399);
nor U19322 (N_19322,N_12088,N_11021);
or U19323 (N_19323,N_14055,N_12830);
nor U19324 (N_19324,N_11533,N_12204);
or U19325 (N_19325,N_10777,N_11606);
xor U19326 (N_19326,N_14232,N_13936);
and U19327 (N_19327,N_14839,N_14841);
xnor U19328 (N_19328,N_10886,N_11870);
nor U19329 (N_19329,N_13820,N_14732);
nand U19330 (N_19330,N_12541,N_13822);
xor U19331 (N_19331,N_11802,N_14442);
nand U19332 (N_19332,N_10490,N_12492);
nand U19333 (N_19333,N_10228,N_11126);
nor U19334 (N_19334,N_14659,N_13770);
nor U19335 (N_19335,N_10373,N_11970);
xnor U19336 (N_19336,N_11311,N_13931);
and U19337 (N_19337,N_10897,N_13948);
and U19338 (N_19338,N_11238,N_14920);
or U19339 (N_19339,N_11480,N_11247);
or U19340 (N_19340,N_10836,N_14612);
or U19341 (N_19341,N_11301,N_10575);
and U19342 (N_19342,N_14988,N_12444);
nor U19343 (N_19343,N_10854,N_10986);
xor U19344 (N_19344,N_13064,N_11961);
xor U19345 (N_19345,N_11625,N_11248);
nor U19346 (N_19346,N_14477,N_14178);
nor U19347 (N_19347,N_14862,N_14876);
and U19348 (N_19348,N_11816,N_14955);
and U19349 (N_19349,N_13207,N_14684);
nor U19350 (N_19350,N_14950,N_14827);
nand U19351 (N_19351,N_12231,N_12428);
xor U19352 (N_19352,N_11567,N_14032);
and U19353 (N_19353,N_10844,N_13720);
nor U19354 (N_19354,N_14246,N_13638);
nor U19355 (N_19355,N_14552,N_11245);
and U19356 (N_19356,N_10183,N_13126);
nand U19357 (N_19357,N_12566,N_13312);
nand U19358 (N_19358,N_13760,N_12782);
and U19359 (N_19359,N_14362,N_13535);
and U19360 (N_19360,N_11905,N_11609);
and U19361 (N_19361,N_12542,N_10679);
and U19362 (N_19362,N_12150,N_14631);
and U19363 (N_19363,N_10142,N_10063);
xor U19364 (N_19364,N_11730,N_14300);
xor U19365 (N_19365,N_10769,N_13327);
and U19366 (N_19366,N_12301,N_12878);
and U19367 (N_19367,N_10370,N_12785);
nand U19368 (N_19368,N_10731,N_12780);
nor U19369 (N_19369,N_11599,N_11940);
nand U19370 (N_19370,N_14576,N_12128);
nand U19371 (N_19371,N_11345,N_10330);
or U19372 (N_19372,N_14394,N_10795);
nand U19373 (N_19373,N_12500,N_10185);
or U19374 (N_19374,N_12758,N_13205);
or U19375 (N_19375,N_12347,N_11561);
nand U19376 (N_19376,N_13543,N_13073);
or U19377 (N_19377,N_13933,N_13936);
xnor U19378 (N_19378,N_13144,N_14405);
and U19379 (N_19379,N_11379,N_10681);
or U19380 (N_19380,N_12557,N_14757);
and U19381 (N_19381,N_11525,N_11567);
or U19382 (N_19382,N_12535,N_12672);
or U19383 (N_19383,N_11453,N_14572);
and U19384 (N_19384,N_14324,N_13291);
or U19385 (N_19385,N_14360,N_13407);
and U19386 (N_19386,N_14403,N_12197);
and U19387 (N_19387,N_12116,N_11464);
or U19388 (N_19388,N_13223,N_11055);
nor U19389 (N_19389,N_12298,N_10506);
or U19390 (N_19390,N_13119,N_11132);
nor U19391 (N_19391,N_13725,N_12974);
xor U19392 (N_19392,N_10819,N_12163);
nor U19393 (N_19393,N_10176,N_12909);
nor U19394 (N_19394,N_10195,N_13651);
nand U19395 (N_19395,N_11439,N_11480);
nor U19396 (N_19396,N_14497,N_13308);
xor U19397 (N_19397,N_12002,N_14482);
nand U19398 (N_19398,N_11363,N_13997);
nor U19399 (N_19399,N_13990,N_11507);
nand U19400 (N_19400,N_13086,N_13893);
xnor U19401 (N_19401,N_11665,N_13426);
or U19402 (N_19402,N_14582,N_13424);
or U19403 (N_19403,N_10278,N_12354);
or U19404 (N_19404,N_10263,N_12810);
nor U19405 (N_19405,N_14129,N_13674);
and U19406 (N_19406,N_12106,N_11325);
or U19407 (N_19407,N_14619,N_14010);
nor U19408 (N_19408,N_12139,N_10586);
and U19409 (N_19409,N_14268,N_14520);
or U19410 (N_19410,N_10656,N_14945);
nor U19411 (N_19411,N_12359,N_11355);
or U19412 (N_19412,N_13046,N_11963);
nand U19413 (N_19413,N_12034,N_13409);
or U19414 (N_19414,N_10232,N_13938);
and U19415 (N_19415,N_11787,N_14757);
and U19416 (N_19416,N_12689,N_11934);
xnor U19417 (N_19417,N_11517,N_13145);
nand U19418 (N_19418,N_13676,N_14763);
and U19419 (N_19419,N_11171,N_12304);
and U19420 (N_19420,N_14535,N_10012);
nand U19421 (N_19421,N_13822,N_14337);
and U19422 (N_19422,N_12262,N_10968);
nand U19423 (N_19423,N_12630,N_11903);
nor U19424 (N_19424,N_14577,N_13183);
or U19425 (N_19425,N_12148,N_11814);
and U19426 (N_19426,N_14575,N_14058);
or U19427 (N_19427,N_11490,N_14393);
and U19428 (N_19428,N_12451,N_12229);
or U19429 (N_19429,N_12522,N_13467);
or U19430 (N_19430,N_14313,N_11570);
nor U19431 (N_19431,N_13899,N_10386);
nand U19432 (N_19432,N_11352,N_10910);
nor U19433 (N_19433,N_13385,N_11689);
nor U19434 (N_19434,N_10744,N_11322);
nand U19435 (N_19435,N_13648,N_11547);
or U19436 (N_19436,N_11009,N_13308);
nand U19437 (N_19437,N_13719,N_14878);
nor U19438 (N_19438,N_14270,N_12332);
or U19439 (N_19439,N_13450,N_10481);
nor U19440 (N_19440,N_14101,N_10259);
nor U19441 (N_19441,N_11976,N_11120);
nand U19442 (N_19442,N_14589,N_14392);
and U19443 (N_19443,N_13729,N_12529);
nand U19444 (N_19444,N_12974,N_14816);
nand U19445 (N_19445,N_11980,N_10146);
and U19446 (N_19446,N_11909,N_11408);
nor U19447 (N_19447,N_11598,N_10783);
nor U19448 (N_19448,N_11630,N_13334);
nor U19449 (N_19449,N_10050,N_11060);
nand U19450 (N_19450,N_10982,N_13047);
or U19451 (N_19451,N_13804,N_10866);
or U19452 (N_19452,N_10757,N_10293);
or U19453 (N_19453,N_10587,N_10291);
and U19454 (N_19454,N_14713,N_10029);
or U19455 (N_19455,N_14690,N_12865);
nor U19456 (N_19456,N_11559,N_14606);
nor U19457 (N_19457,N_13562,N_12992);
nor U19458 (N_19458,N_13739,N_11247);
nand U19459 (N_19459,N_13225,N_12458);
nand U19460 (N_19460,N_12671,N_10517);
nand U19461 (N_19461,N_11500,N_10593);
nor U19462 (N_19462,N_13608,N_14187);
nand U19463 (N_19463,N_10207,N_13590);
xor U19464 (N_19464,N_12893,N_14473);
or U19465 (N_19465,N_11505,N_12632);
nor U19466 (N_19466,N_13055,N_10727);
nor U19467 (N_19467,N_14053,N_13293);
nor U19468 (N_19468,N_11842,N_10323);
nor U19469 (N_19469,N_13441,N_12901);
nand U19470 (N_19470,N_11426,N_10313);
or U19471 (N_19471,N_11641,N_11341);
nand U19472 (N_19472,N_10697,N_12537);
or U19473 (N_19473,N_11771,N_10287);
xnor U19474 (N_19474,N_11315,N_13267);
and U19475 (N_19475,N_11679,N_11044);
nor U19476 (N_19476,N_13592,N_13102);
nor U19477 (N_19477,N_14089,N_11099);
or U19478 (N_19478,N_11071,N_11964);
nand U19479 (N_19479,N_12312,N_10230);
and U19480 (N_19480,N_10205,N_10651);
and U19481 (N_19481,N_12707,N_12496);
xnor U19482 (N_19482,N_14918,N_13415);
nand U19483 (N_19483,N_11683,N_13303);
nor U19484 (N_19484,N_13422,N_13491);
nand U19485 (N_19485,N_12569,N_10247);
nor U19486 (N_19486,N_14359,N_10289);
or U19487 (N_19487,N_14005,N_13368);
nand U19488 (N_19488,N_14869,N_12138);
xnor U19489 (N_19489,N_13271,N_13201);
nor U19490 (N_19490,N_10903,N_11012);
nor U19491 (N_19491,N_10035,N_10401);
nor U19492 (N_19492,N_12690,N_12817);
and U19493 (N_19493,N_11094,N_13479);
and U19494 (N_19494,N_10653,N_13837);
and U19495 (N_19495,N_12460,N_12608);
nor U19496 (N_19496,N_13979,N_12089);
and U19497 (N_19497,N_14117,N_11598);
or U19498 (N_19498,N_12615,N_11612);
xor U19499 (N_19499,N_14887,N_11376);
or U19500 (N_19500,N_11673,N_10178);
xor U19501 (N_19501,N_10351,N_10494);
and U19502 (N_19502,N_11841,N_13649);
nand U19503 (N_19503,N_13500,N_14849);
and U19504 (N_19504,N_11144,N_13955);
nand U19505 (N_19505,N_14001,N_14298);
nor U19506 (N_19506,N_14881,N_14643);
and U19507 (N_19507,N_13028,N_11823);
nand U19508 (N_19508,N_13722,N_14516);
or U19509 (N_19509,N_12653,N_13439);
and U19510 (N_19510,N_14347,N_13827);
nand U19511 (N_19511,N_12317,N_13629);
and U19512 (N_19512,N_10266,N_14672);
nand U19513 (N_19513,N_14350,N_12473);
nand U19514 (N_19514,N_13575,N_13503);
or U19515 (N_19515,N_11160,N_10105);
nor U19516 (N_19516,N_11360,N_10630);
xor U19517 (N_19517,N_11503,N_11110);
or U19518 (N_19518,N_13006,N_13700);
xnor U19519 (N_19519,N_11521,N_14250);
nand U19520 (N_19520,N_12360,N_12919);
xor U19521 (N_19521,N_11170,N_14125);
nor U19522 (N_19522,N_14117,N_14392);
or U19523 (N_19523,N_12660,N_10800);
or U19524 (N_19524,N_10761,N_11458);
nor U19525 (N_19525,N_14992,N_13518);
nor U19526 (N_19526,N_14016,N_13715);
nor U19527 (N_19527,N_10644,N_14859);
and U19528 (N_19528,N_12191,N_10584);
nor U19529 (N_19529,N_13861,N_14246);
or U19530 (N_19530,N_12728,N_14713);
xor U19531 (N_19531,N_11039,N_14543);
and U19532 (N_19532,N_11524,N_13617);
nand U19533 (N_19533,N_10267,N_11504);
or U19534 (N_19534,N_11096,N_13282);
nor U19535 (N_19535,N_13948,N_11346);
xor U19536 (N_19536,N_14710,N_13717);
nor U19537 (N_19537,N_14936,N_13502);
nand U19538 (N_19538,N_11146,N_11927);
xnor U19539 (N_19539,N_11594,N_13632);
nand U19540 (N_19540,N_10026,N_10216);
nand U19541 (N_19541,N_12375,N_13676);
or U19542 (N_19542,N_10830,N_12353);
nor U19543 (N_19543,N_12432,N_12455);
and U19544 (N_19544,N_10296,N_14984);
or U19545 (N_19545,N_13619,N_14402);
nor U19546 (N_19546,N_12613,N_10857);
or U19547 (N_19547,N_12881,N_14680);
xor U19548 (N_19548,N_12452,N_11527);
or U19549 (N_19549,N_12179,N_14242);
nor U19550 (N_19550,N_13411,N_12428);
nand U19551 (N_19551,N_14792,N_12140);
or U19552 (N_19552,N_12913,N_11922);
and U19553 (N_19553,N_12757,N_12662);
or U19554 (N_19554,N_12182,N_13530);
nand U19555 (N_19555,N_14727,N_13597);
nor U19556 (N_19556,N_11308,N_13718);
xnor U19557 (N_19557,N_12663,N_13835);
or U19558 (N_19558,N_14734,N_13158);
nor U19559 (N_19559,N_11031,N_12500);
nor U19560 (N_19560,N_12414,N_12408);
nor U19561 (N_19561,N_13294,N_11619);
or U19562 (N_19562,N_10035,N_10662);
nor U19563 (N_19563,N_14504,N_12225);
nand U19564 (N_19564,N_10646,N_14084);
and U19565 (N_19565,N_12957,N_11141);
xor U19566 (N_19566,N_13127,N_11619);
nor U19567 (N_19567,N_12889,N_11571);
or U19568 (N_19568,N_13918,N_11579);
xnor U19569 (N_19569,N_11439,N_10382);
nand U19570 (N_19570,N_11315,N_13747);
and U19571 (N_19571,N_13650,N_13031);
nor U19572 (N_19572,N_10936,N_13370);
or U19573 (N_19573,N_14053,N_10054);
nor U19574 (N_19574,N_12934,N_11730);
nor U19575 (N_19575,N_13243,N_13937);
nor U19576 (N_19576,N_12765,N_14403);
and U19577 (N_19577,N_11298,N_11254);
and U19578 (N_19578,N_10208,N_11257);
nand U19579 (N_19579,N_14231,N_13745);
nand U19580 (N_19580,N_12692,N_12362);
xnor U19581 (N_19581,N_13360,N_13396);
or U19582 (N_19582,N_12000,N_10728);
or U19583 (N_19583,N_10185,N_14290);
and U19584 (N_19584,N_11528,N_14685);
nand U19585 (N_19585,N_13721,N_14711);
or U19586 (N_19586,N_12769,N_10320);
nand U19587 (N_19587,N_12586,N_14338);
nand U19588 (N_19588,N_10142,N_10718);
nor U19589 (N_19589,N_10345,N_12774);
nand U19590 (N_19590,N_13859,N_11903);
or U19591 (N_19591,N_11594,N_13704);
or U19592 (N_19592,N_11445,N_11114);
nor U19593 (N_19593,N_13145,N_10503);
and U19594 (N_19594,N_13762,N_11065);
or U19595 (N_19595,N_14319,N_11319);
xor U19596 (N_19596,N_13395,N_14123);
xor U19597 (N_19597,N_10800,N_14308);
nand U19598 (N_19598,N_14739,N_13333);
xnor U19599 (N_19599,N_11786,N_10863);
nor U19600 (N_19600,N_13085,N_11568);
xor U19601 (N_19601,N_13211,N_13041);
and U19602 (N_19602,N_10624,N_11857);
nand U19603 (N_19603,N_10194,N_11815);
xnor U19604 (N_19604,N_13732,N_12788);
xor U19605 (N_19605,N_13841,N_14339);
or U19606 (N_19606,N_10224,N_13750);
and U19607 (N_19607,N_13903,N_14937);
nand U19608 (N_19608,N_13040,N_13656);
xnor U19609 (N_19609,N_11792,N_12521);
or U19610 (N_19610,N_13970,N_11228);
nand U19611 (N_19611,N_13031,N_10612);
xnor U19612 (N_19612,N_11433,N_11157);
or U19613 (N_19613,N_12293,N_13653);
nand U19614 (N_19614,N_11688,N_13515);
or U19615 (N_19615,N_10574,N_12501);
nor U19616 (N_19616,N_13830,N_13401);
nand U19617 (N_19617,N_14390,N_14321);
or U19618 (N_19618,N_10182,N_10196);
or U19619 (N_19619,N_10617,N_13116);
or U19620 (N_19620,N_11175,N_14215);
and U19621 (N_19621,N_13714,N_12866);
nor U19622 (N_19622,N_11615,N_14308);
or U19623 (N_19623,N_12386,N_13144);
nor U19624 (N_19624,N_11669,N_13890);
nand U19625 (N_19625,N_11002,N_12808);
and U19626 (N_19626,N_10699,N_10770);
nand U19627 (N_19627,N_12284,N_10459);
or U19628 (N_19628,N_12980,N_12984);
nor U19629 (N_19629,N_10587,N_12121);
nand U19630 (N_19630,N_11588,N_12435);
or U19631 (N_19631,N_13769,N_13764);
nand U19632 (N_19632,N_10856,N_10718);
and U19633 (N_19633,N_14877,N_12386);
and U19634 (N_19634,N_12886,N_10066);
nor U19635 (N_19635,N_11861,N_13929);
and U19636 (N_19636,N_10006,N_13800);
nor U19637 (N_19637,N_10747,N_12875);
nand U19638 (N_19638,N_14672,N_13609);
nand U19639 (N_19639,N_11586,N_14505);
and U19640 (N_19640,N_10909,N_13509);
nand U19641 (N_19641,N_10082,N_10306);
and U19642 (N_19642,N_14895,N_11238);
or U19643 (N_19643,N_13717,N_12210);
nor U19644 (N_19644,N_10339,N_11096);
nor U19645 (N_19645,N_12289,N_11698);
xor U19646 (N_19646,N_13431,N_10357);
nor U19647 (N_19647,N_13294,N_14478);
nor U19648 (N_19648,N_14905,N_12499);
or U19649 (N_19649,N_14713,N_11687);
xor U19650 (N_19650,N_10666,N_12014);
and U19651 (N_19651,N_12317,N_11657);
nand U19652 (N_19652,N_12514,N_10066);
nand U19653 (N_19653,N_11580,N_11944);
nor U19654 (N_19654,N_12277,N_11499);
or U19655 (N_19655,N_11797,N_11642);
or U19656 (N_19656,N_11906,N_10193);
or U19657 (N_19657,N_13609,N_10823);
nor U19658 (N_19658,N_10790,N_11445);
nor U19659 (N_19659,N_10828,N_11690);
nor U19660 (N_19660,N_12741,N_14040);
xnor U19661 (N_19661,N_11767,N_11313);
nand U19662 (N_19662,N_14624,N_13520);
or U19663 (N_19663,N_10697,N_10339);
or U19664 (N_19664,N_12054,N_12329);
or U19665 (N_19665,N_13286,N_12472);
nor U19666 (N_19666,N_14910,N_13372);
xnor U19667 (N_19667,N_12204,N_12684);
nor U19668 (N_19668,N_12744,N_14569);
nor U19669 (N_19669,N_12628,N_10530);
or U19670 (N_19670,N_14474,N_10725);
or U19671 (N_19671,N_12402,N_13219);
or U19672 (N_19672,N_14486,N_10706);
nand U19673 (N_19673,N_13919,N_10031);
or U19674 (N_19674,N_14396,N_13310);
nand U19675 (N_19675,N_10563,N_12853);
xor U19676 (N_19676,N_12455,N_14049);
and U19677 (N_19677,N_11593,N_14082);
nor U19678 (N_19678,N_14693,N_11102);
nor U19679 (N_19679,N_13726,N_12491);
nor U19680 (N_19680,N_12531,N_14524);
or U19681 (N_19681,N_13586,N_12345);
and U19682 (N_19682,N_13767,N_11909);
or U19683 (N_19683,N_13210,N_11597);
and U19684 (N_19684,N_11698,N_14336);
or U19685 (N_19685,N_11871,N_14422);
nor U19686 (N_19686,N_14296,N_11387);
xor U19687 (N_19687,N_12477,N_10331);
and U19688 (N_19688,N_12002,N_14901);
nand U19689 (N_19689,N_11597,N_10050);
xor U19690 (N_19690,N_14628,N_13122);
or U19691 (N_19691,N_13749,N_12712);
and U19692 (N_19692,N_10469,N_14081);
nor U19693 (N_19693,N_11290,N_13907);
and U19694 (N_19694,N_14059,N_12383);
nor U19695 (N_19695,N_10499,N_10234);
nand U19696 (N_19696,N_13745,N_14048);
and U19697 (N_19697,N_13860,N_13177);
nor U19698 (N_19698,N_13195,N_11916);
or U19699 (N_19699,N_10559,N_12278);
and U19700 (N_19700,N_14120,N_10784);
or U19701 (N_19701,N_11034,N_14788);
and U19702 (N_19702,N_12308,N_14276);
and U19703 (N_19703,N_13543,N_11087);
nor U19704 (N_19704,N_13949,N_11757);
and U19705 (N_19705,N_10040,N_10389);
nand U19706 (N_19706,N_12284,N_13813);
and U19707 (N_19707,N_13214,N_12037);
xnor U19708 (N_19708,N_14296,N_10137);
nor U19709 (N_19709,N_10356,N_12453);
or U19710 (N_19710,N_14214,N_12796);
and U19711 (N_19711,N_11759,N_12966);
or U19712 (N_19712,N_12550,N_14112);
nand U19713 (N_19713,N_13246,N_14122);
nor U19714 (N_19714,N_12263,N_10272);
or U19715 (N_19715,N_10229,N_12462);
and U19716 (N_19716,N_10016,N_12157);
and U19717 (N_19717,N_13251,N_13306);
or U19718 (N_19718,N_14460,N_14218);
nor U19719 (N_19719,N_12444,N_13193);
or U19720 (N_19720,N_12372,N_11495);
nand U19721 (N_19721,N_10657,N_10052);
and U19722 (N_19722,N_12346,N_14893);
nor U19723 (N_19723,N_12850,N_13576);
or U19724 (N_19724,N_14921,N_11805);
and U19725 (N_19725,N_12341,N_11650);
nor U19726 (N_19726,N_10024,N_12026);
nor U19727 (N_19727,N_10378,N_12267);
or U19728 (N_19728,N_10832,N_10212);
and U19729 (N_19729,N_10873,N_12382);
nor U19730 (N_19730,N_10790,N_13301);
nand U19731 (N_19731,N_13647,N_12392);
nor U19732 (N_19732,N_12711,N_14657);
or U19733 (N_19733,N_14152,N_12494);
and U19734 (N_19734,N_12920,N_10669);
or U19735 (N_19735,N_10629,N_10691);
nor U19736 (N_19736,N_10755,N_11838);
nor U19737 (N_19737,N_12280,N_12869);
nand U19738 (N_19738,N_12609,N_11211);
nand U19739 (N_19739,N_10514,N_12079);
nand U19740 (N_19740,N_13161,N_13315);
nor U19741 (N_19741,N_12938,N_12834);
nand U19742 (N_19742,N_13787,N_12812);
and U19743 (N_19743,N_10830,N_12623);
and U19744 (N_19744,N_14957,N_13480);
nor U19745 (N_19745,N_14870,N_13211);
xor U19746 (N_19746,N_12682,N_12390);
nor U19747 (N_19747,N_13221,N_14268);
nand U19748 (N_19748,N_11216,N_13320);
or U19749 (N_19749,N_13658,N_13783);
and U19750 (N_19750,N_13392,N_12121);
and U19751 (N_19751,N_11716,N_14688);
or U19752 (N_19752,N_10181,N_10368);
or U19753 (N_19753,N_11787,N_10720);
and U19754 (N_19754,N_12294,N_14277);
nand U19755 (N_19755,N_11310,N_13100);
and U19756 (N_19756,N_14404,N_10314);
nor U19757 (N_19757,N_10514,N_14369);
nor U19758 (N_19758,N_11659,N_14208);
nor U19759 (N_19759,N_11546,N_10320);
nand U19760 (N_19760,N_11591,N_11084);
nand U19761 (N_19761,N_12137,N_10391);
xnor U19762 (N_19762,N_12381,N_11893);
nand U19763 (N_19763,N_11231,N_12686);
nand U19764 (N_19764,N_12232,N_12111);
xnor U19765 (N_19765,N_12306,N_12416);
nor U19766 (N_19766,N_13683,N_12592);
nand U19767 (N_19767,N_12893,N_10565);
and U19768 (N_19768,N_10238,N_14984);
nand U19769 (N_19769,N_11900,N_11395);
nand U19770 (N_19770,N_11618,N_11117);
or U19771 (N_19771,N_12222,N_11648);
nand U19772 (N_19772,N_13507,N_11961);
nand U19773 (N_19773,N_11953,N_12701);
xnor U19774 (N_19774,N_13308,N_13498);
nor U19775 (N_19775,N_10342,N_14993);
nand U19776 (N_19776,N_14994,N_13748);
nor U19777 (N_19777,N_14851,N_11745);
and U19778 (N_19778,N_12674,N_12083);
xor U19779 (N_19779,N_14051,N_10561);
nor U19780 (N_19780,N_11028,N_11931);
nor U19781 (N_19781,N_14551,N_13625);
xnor U19782 (N_19782,N_10907,N_14360);
xor U19783 (N_19783,N_13216,N_11628);
and U19784 (N_19784,N_13427,N_11473);
xor U19785 (N_19785,N_12941,N_14496);
nand U19786 (N_19786,N_13284,N_14454);
nor U19787 (N_19787,N_12785,N_11697);
nand U19788 (N_19788,N_14285,N_13048);
nand U19789 (N_19789,N_13904,N_10823);
and U19790 (N_19790,N_10468,N_10487);
nand U19791 (N_19791,N_10267,N_10608);
xor U19792 (N_19792,N_11444,N_13797);
nand U19793 (N_19793,N_11885,N_14435);
nand U19794 (N_19794,N_10845,N_12096);
xnor U19795 (N_19795,N_14437,N_13275);
and U19796 (N_19796,N_11555,N_12238);
and U19797 (N_19797,N_10558,N_12209);
and U19798 (N_19798,N_13354,N_13395);
and U19799 (N_19799,N_13208,N_14172);
nor U19800 (N_19800,N_10753,N_14460);
nand U19801 (N_19801,N_12464,N_14371);
nor U19802 (N_19802,N_14706,N_10928);
nand U19803 (N_19803,N_13854,N_14819);
or U19804 (N_19804,N_10553,N_12885);
nor U19805 (N_19805,N_10566,N_12310);
or U19806 (N_19806,N_14622,N_11857);
nand U19807 (N_19807,N_11444,N_11055);
and U19808 (N_19808,N_11035,N_14271);
xor U19809 (N_19809,N_13201,N_14863);
xor U19810 (N_19810,N_10798,N_13753);
nor U19811 (N_19811,N_14858,N_10235);
nand U19812 (N_19812,N_14618,N_12154);
nand U19813 (N_19813,N_12336,N_13992);
xnor U19814 (N_19814,N_11026,N_12477);
or U19815 (N_19815,N_14576,N_11583);
or U19816 (N_19816,N_13324,N_14311);
and U19817 (N_19817,N_13238,N_13127);
or U19818 (N_19818,N_13720,N_10116);
and U19819 (N_19819,N_13847,N_14570);
and U19820 (N_19820,N_13783,N_12633);
nor U19821 (N_19821,N_12874,N_10090);
or U19822 (N_19822,N_12433,N_12712);
nor U19823 (N_19823,N_12497,N_10511);
nor U19824 (N_19824,N_10295,N_12430);
xnor U19825 (N_19825,N_13609,N_14057);
and U19826 (N_19826,N_11654,N_11260);
nor U19827 (N_19827,N_11240,N_11484);
nand U19828 (N_19828,N_12840,N_10436);
or U19829 (N_19829,N_12591,N_10992);
and U19830 (N_19830,N_10959,N_11460);
nor U19831 (N_19831,N_11991,N_13440);
or U19832 (N_19832,N_14912,N_12982);
nor U19833 (N_19833,N_10407,N_10261);
nand U19834 (N_19834,N_10115,N_11880);
and U19835 (N_19835,N_11254,N_10312);
and U19836 (N_19836,N_10672,N_14359);
nor U19837 (N_19837,N_14495,N_13438);
nand U19838 (N_19838,N_13109,N_13399);
or U19839 (N_19839,N_14116,N_11593);
and U19840 (N_19840,N_11021,N_13625);
nor U19841 (N_19841,N_11787,N_12808);
and U19842 (N_19842,N_13279,N_11428);
and U19843 (N_19843,N_11376,N_11605);
nand U19844 (N_19844,N_10704,N_14625);
xnor U19845 (N_19845,N_12351,N_11122);
and U19846 (N_19846,N_10171,N_13405);
xnor U19847 (N_19847,N_13734,N_10414);
or U19848 (N_19848,N_14920,N_13873);
and U19849 (N_19849,N_14564,N_10926);
nand U19850 (N_19850,N_14245,N_11898);
xnor U19851 (N_19851,N_13103,N_13536);
nand U19852 (N_19852,N_13554,N_12248);
and U19853 (N_19853,N_12764,N_12496);
nor U19854 (N_19854,N_10644,N_14025);
nand U19855 (N_19855,N_12897,N_10526);
xnor U19856 (N_19856,N_10796,N_14187);
nand U19857 (N_19857,N_13230,N_13811);
or U19858 (N_19858,N_13707,N_13720);
or U19859 (N_19859,N_14223,N_12693);
nand U19860 (N_19860,N_11603,N_13757);
and U19861 (N_19861,N_13654,N_12200);
and U19862 (N_19862,N_11925,N_12052);
nand U19863 (N_19863,N_11222,N_12324);
nor U19864 (N_19864,N_11159,N_11104);
nand U19865 (N_19865,N_13582,N_14999);
and U19866 (N_19866,N_14602,N_13835);
nand U19867 (N_19867,N_10710,N_10702);
nor U19868 (N_19868,N_14314,N_14546);
and U19869 (N_19869,N_10042,N_12039);
nor U19870 (N_19870,N_12186,N_11945);
and U19871 (N_19871,N_10511,N_14605);
and U19872 (N_19872,N_13125,N_14216);
and U19873 (N_19873,N_13048,N_13389);
and U19874 (N_19874,N_13030,N_14704);
nand U19875 (N_19875,N_14844,N_10559);
nand U19876 (N_19876,N_12732,N_10448);
nor U19877 (N_19877,N_11620,N_11733);
nor U19878 (N_19878,N_12494,N_10780);
nand U19879 (N_19879,N_12374,N_14925);
xnor U19880 (N_19880,N_10385,N_10110);
and U19881 (N_19881,N_13672,N_12273);
or U19882 (N_19882,N_14668,N_13432);
nand U19883 (N_19883,N_11166,N_12648);
nor U19884 (N_19884,N_10353,N_14929);
or U19885 (N_19885,N_10371,N_12690);
or U19886 (N_19886,N_11726,N_10140);
nand U19887 (N_19887,N_12316,N_11843);
nor U19888 (N_19888,N_11558,N_14162);
or U19889 (N_19889,N_12456,N_11883);
nor U19890 (N_19890,N_12465,N_11712);
nand U19891 (N_19891,N_14379,N_11534);
nand U19892 (N_19892,N_12779,N_11600);
nand U19893 (N_19893,N_14198,N_10092);
and U19894 (N_19894,N_11442,N_13905);
nand U19895 (N_19895,N_10830,N_13203);
nor U19896 (N_19896,N_10536,N_14982);
nand U19897 (N_19897,N_13660,N_11491);
or U19898 (N_19898,N_11358,N_10833);
or U19899 (N_19899,N_14248,N_12031);
nand U19900 (N_19900,N_11250,N_13014);
xor U19901 (N_19901,N_12367,N_14071);
nor U19902 (N_19902,N_10706,N_13415);
nand U19903 (N_19903,N_12275,N_10448);
nand U19904 (N_19904,N_14425,N_13999);
and U19905 (N_19905,N_13298,N_11900);
and U19906 (N_19906,N_13814,N_11513);
nor U19907 (N_19907,N_12897,N_13036);
nor U19908 (N_19908,N_14587,N_12104);
or U19909 (N_19909,N_12486,N_11515);
nand U19910 (N_19910,N_13064,N_13851);
nor U19911 (N_19911,N_14364,N_12511);
nand U19912 (N_19912,N_10863,N_14625);
nor U19913 (N_19913,N_11309,N_14026);
nand U19914 (N_19914,N_14273,N_12121);
or U19915 (N_19915,N_12252,N_10028);
xnor U19916 (N_19916,N_11326,N_11131);
nand U19917 (N_19917,N_12367,N_13526);
and U19918 (N_19918,N_14282,N_11243);
nor U19919 (N_19919,N_13469,N_13916);
and U19920 (N_19920,N_10894,N_12902);
nand U19921 (N_19921,N_14661,N_14276);
nor U19922 (N_19922,N_11888,N_10300);
xor U19923 (N_19923,N_12927,N_14806);
and U19924 (N_19924,N_13759,N_12664);
or U19925 (N_19925,N_10921,N_14916);
and U19926 (N_19926,N_11769,N_13448);
nor U19927 (N_19927,N_10318,N_12535);
xor U19928 (N_19928,N_10055,N_13904);
and U19929 (N_19929,N_14918,N_11457);
and U19930 (N_19930,N_13087,N_13191);
nand U19931 (N_19931,N_13490,N_14778);
nand U19932 (N_19932,N_13692,N_10120);
nand U19933 (N_19933,N_14013,N_11460);
nand U19934 (N_19934,N_12581,N_13141);
nor U19935 (N_19935,N_14723,N_12252);
nand U19936 (N_19936,N_12912,N_14662);
or U19937 (N_19937,N_10982,N_13084);
nand U19938 (N_19938,N_12366,N_10231);
nand U19939 (N_19939,N_13196,N_14953);
nor U19940 (N_19940,N_13234,N_10572);
and U19941 (N_19941,N_13294,N_10006);
and U19942 (N_19942,N_11074,N_12640);
or U19943 (N_19943,N_11177,N_12966);
nand U19944 (N_19944,N_12726,N_12366);
and U19945 (N_19945,N_10822,N_12618);
or U19946 (N_19946,N_14936,N_14462);
and U19947 (N_19947,N_10044,N_11444);
and U19948 (N_19948,N_13149,N_13109);
nand U19949 (N_19949,N_12412,N_10963);
nor U19950 (N_19950,N_13231,N_14461);
nand U19951 (N_19951,N_12054,N_13863);
or U19952 (N_19952,N_14681,N_10851);
nor U19953 (N_19953,N_10478,N_11795);
and U19954 (N_19954,N_13599,N_14815);
and U19955 (N_19955,N_13312,N_12052);
and U19956 (N_19956,N_12925,N_11835);
nor U19957 (N_19957,N_12162,N_13507);
nand U19958 (N_19958,N_14129,N_14293);
or U19959 (N_19959,N_11336,N_11290);
and U19960 (N_19960,N_13439,N_10150);
nand U19961 (N_19961,N_13948,N_12054);
nor U19962 (N_19962,N_14410,N_10770);
nor U19963 (N_19963,N_10572,N_10970);
and U19964 (N_19964,N_13565,N_11943);
and U19965 (N_19965,N_12219,N_14175);
nor U19966 (N_19966,N_13015,N_13277);
nor U19967 (N_19967,N_13012,N_13609);
xnor U19968 (N_19968,N_13178,N_10950);
or U19969 (N_19969,N_11999,N_10602);
nor U19970 (N_19970,N_14679,N_10479);
and U19971 (N_19971,N_10093,N_10160);
nor U19972 (N_19972,N_14432,N_11064);
or U19973 (N_19973,N_13067,N_14591);
and U19974 (N_19974,N_13141,N_13937);
xnor U19975 (N_19975,N_10783,N_10452);
and U19976 (N_19976,N_13768,N_10601);
and U19977 (N_19977,N_10913,N_11585);
and U19978 (N_19978,N_11468,N_10993);
nor U19979 (N_19979,N_12345,N_14423);
nor U19980 (N_19980,N_12668,N_14362);
nand U19981 (N_19981,N_14338,N_12669);
nand U19982 (N_19982,N_11372,N_12339);
nand U19983 (N_19983,N_12722,N_13953);
or U19984 (N_19984,N_10497,N_14158);
nand U19985 (N_19985,N_12005,N_12466);
nor U19986 (N_19986,N_10113,N_12353);
nor U19987 (N_19987,N_12434,N_10572);
nand U19988 (N_19988,N_14052,N_12784);
nor U19989 (N_19989,N_14685,N_10952);
xnor U19990 (N_19990,N_14977,N_10885);
and U19991 (N_19991,N_12877,N_14020);
or U19992 (N_19992,N_12837,N_12349);
nor U19993 (N_19993,N_10620,N_11378);
nor U19994 (N_19994,N_13514,N_13841);
and U19995 (N_19995,N_11585,N_11058);
and U19996 (N_19996,N_10972,N_12005);
nand U19997 (N_19997,N_14463,N_13652);
or U19998 (N_19998,N_10475,N_11657);
and U19999 (N_19999,N_14878,N_12368);
and UO_0 (O_0,N_16855,N_16170);
nor UO_1 (O_1,N_16542,N_19746);
or UO_2 (O_2,N_18778,N_16452);
nand UO_3 (O_3,N_19828,N_19320);
or UO_4 (O_4,N_15838,N_17360);
or UO_5 (O_5,N_17538,N_18283);
and UO_6 (O_6,N_18391,N_16498);
nor UO_7 (O_7,N_19816,N_17509);
xnor UO_8 (O_8,N_17397,N_18518);
nand UO_9 (O_9,N_17846,N_16196);
or UO_10 (O_10,N_17553,N_18953);
or UO_11 (O_11,N_19046,N_19059);
xnor UO_12 (O_12,N_16526,N_17441);
nor UO_13 (O_13,N_18715,N_15177);
or UO_14 (O_14,N_16784,N_16928);
and UO_15 (O_15,N_19571,N_19726);
nand UO_16 (O_16,N_15604,N_16535);
and UO_17 (O_17,N_18884,N_19885);
nand UO_18 (O_18,N_18871,N_16415);
nand UO_19 (O_19,N_19891,N_16358);
nor UO_20 (O_20,N_18030,N_19245);
nand UO_21 (O_21,N_19097,N_17202);
or UO_22 (O_22,N_18207,N_15511);
or UO_23 (O_23,N_18968,N_16681);
or UO_24 (O_24,N_15529,N_19590);
and UO_25 (O_25,N_18098,N_16128);
nand UO_26 (O_26,N_17077,N_19566);
nor UO_27 (O_27,N_16878,N_15718);
and UO_28 (O_28,N_19584,N_18134);
xor UO_29 (O_29,N_19485,N_15446);
or UO_30 (O_30,N_15612,N_16854);
nand UO_31 (O_31,N_17948,N_19294);
or UO_32 (O_32,N_18370,N_16625);
nor UO_33 (O_33,N_16605,N_19112);
xnor UO_34 (O_34,N_17548,N_16617);
nor UO_35 (O_35,N_16748,N_17409);
or UO_36 (O_36,N_18297,N_17103);
and UO_37 (O_37,N_16611,N_16538);
nand UO_38 (O_38,N_18656,N_15104);
and UO_39 (O_39,N_19692,N_15664);
nand UO_40 (O_40,N_15912,N_19183);
or UO_41 (O_41,N_18474,N_17781);
nor UO_42 (O_42,N_15115,N_16081);
and UO_43 (O_43,N_16040,N_19626);
nand UO_44 (O_44,N_16959,N_15433);
nor UO_45 (O_45,N_18050,N_18442);
nor UO_46 (O_46,N_18709,N_16810);
nand UO_47 (O_47,N_17107,N_15903);
nand UO_48 (O_48,N_15130,N_17101);
or UO_49 (O_49,N_15083,N_19738);
or UO_50 (O_50,N_16824,N_19090);
or UO_51 (O_51,N_15327,N_19895);
nor UO_52 (O_52,N_15830,N_16127);
nand UO_53 (O_53,N_16754,N_17765);
or UO_54 (O_54,N_17938,N_19897);
nand UO_55 (O_55,N_16390,N_17182);
nand UO_56 (O_56,N_17297,N_16279);
and UO_57 (O_57,N_17008,N_15404);
nand UO_58 (O_58,N_17779,N_19005);
and UO_59 (O_59,N_18914,N_19964);
nor UO_60 (O_60,N_18460,N_17542);
and UO_61 (O_61,N_16378,N_16125);
nor UO_62 (O_62,N_15198,N_16494);
nor UO_63 (O_63,N_19954,N_19055);
nand UO_64 (O_64,N_16946,N_19727);
and UO_65 (O_65,N_16579,N_18482);
nand UO_66 (O_66,N_17595,N_19283);
nor UO_67 (O_67,N_16235,N_16168);
nand UO_68 (O_68,N_17573,N_17447);
xnor UO_69 (O_69,N_17823,N_19280);
nor UO_70 (O_70,N_19741,N_18363);
and UO_71 (O_71,N_19711,N_15532);
xnor UO_72 (O_72,N_15243,N_16471);
nor UO_73 (O_73,N_18171,N_17139);
nand UO_74 (O_74,N_16155,N_17651);
and UO_75 (O_75,N_15591,N_18492);
and UO_76 (O_76,N_17104,N_18885);
xnor UO_77 (O_77,N_19596,N_16961);
nand UO_78 (O_78,N_15753,N_19036);
xor UO_79 (O_79,N_16366,N_15242);
nand UO_80 (O_80,N_15008,N_17115);
nor UO_81 (O_81,N_19884,N_17195);
or UO_82 (O_82,N_17418,N_18429);
and UO_83 (O_83,N_18570,N_15096);
and UO_84 (O_84,N_17493,N_15970);
nor UO_85 (O_85,N_15452,N_18372);
or UO_86 (O_86,N_19969,N_17567);
nor UO_87 (O_87,N_19017,N_17436);
xnor UO_88 (O_88,N_16757,N_15963);
and UO_89 (O_89,N_16334,N_18658);
or UO_90 (O_90,N_17124,N_15190);
or UO_91 (O_91,N_19344,N_15081);
or UO_92 (O_92,N_17731,N_19122);
or UO_93 (O_93,N_17109,N_16112);
and UO_94 (O_94,N_17970,N_18143);
nand UO_95 (O_95,N_18589,N_17535);
xnor UO_96 (O_96,N_16315,N_18137);
nand UO_97 (O_97,N_16372,N_16092);
and UO_98 (O_98,N_15809,N_18354);
nand UO_99 (O_99,N_15229,N_17140);
nand UO_100 (O_100,N_17400,N_16259);
nand UO_101 (O_101,N_16407,N_18996);
nand UO_102 (O_102,N_15748,N_18959);
xor UO_103 (O_103,N_16889,N_18619);
nand UO_104 (O_104,N_16003,N_16276);
nor UO_105 (O_105,N_17749,N_17971);
and UO_106 (O_106,N_18291,N_18802);
and UO_107 (O_107,N_19247,N_17677);
nand UO_108 (O_108,N_17772,N_19671);
and UO_109 (O_109,N_15364,N_18052);
or UO_110 (O_110,N_18287,N_19364);
nor UO_111 (O_111,N_15867,N_16693);
nor UO_112 (O_112,N_17399,N_18168);
nand UO_113 (O_113,N_18866,N_18870);
nor UO_114 (O_114,N_18795,N_16565);
nor UO_115 (O_115,N_19502,N_15413);
or UO_116 (O_116,N_17836,N_19603);
or UO_117 (O_117,N_17078,N_17773);
nor UO_118 (O_118,N_17009,N_18558);
nor UO_119 (O_119,N_18334,N_15031);
and UO_120 (O_120,N_19213,N_19299);
or UO_121 (O_121,N_17830,N_16570);
and UO_122 (O_122,N_15667,N_19306);
nand UO_123 (O_123,N_17189,N_17745);
nor UO_124 (O_124,N_16786,N_18002);
or UO_125 (O_125,N_16422,N_15799);
and UO_126 (O_126,N_19988,N_17430);
nand UO_127 (O_127,N_16489,N_16432);
nor UO_128 (O_128,N_16661,N_16894);
nand UO_129 (O_129,N_15567,N_18095);
nor UO_130 (O_130,N_19693,N_16343);
or UO_131 (O_131,N_15510,N_19417);
nor UO_132 (O_132,N_16266,N_18780);
and UO_133 (O_133,N_19889,N_15235);
and UO_134 (O_134,N_17964,N_17648);
and UO_135 (O_135,N_18472,N_19553);
nor UO_136 (O_136,N_18629,N_18853);
and UO_137 (O_137,N_16572,N_19825);
nor UO_138 (O_138,N_15998,N_16180);
and UO_139 (O_139,N_17983,N_19781);
and UO_140 (O_140,N_16865,N_18874);
nor UO_141 (O_141,N_17005,N_15589);
nor UO_142 (O_142,N_15048,N_16553);
nor UO_143 (O_143,N_18265,N_18009);
and UO_144 (O_144,N_19117,N_17105);
xor UO_145 (O_145,N_17456,N_15440);
and UO_146 (O_146,N_16727,N_16654);
or UO_147 (O_147,N_15714,N_18100);
nor UO_148 (O_148,N_19953,N_16778);
and UO_149 (O_149,N_15683,N_17741);
nand UO_150 (O_150,N_15142,N_17294);
xnor UO_151 (O_151,N_17564,N_19611);
nand UO_152 (O_152,N_16253,N_19794);
nor UO_153 (O_153,N_19841,N_19628);
nand UO_154 (O_154,N_16598,N_18110);
or UO_155 (O_155,N_15794,N_19922);
xnor UO_156 (O_156,N_19893,N_17697);
or UO_157 (O_157,N_17874,N_17762);
nand UO_158 (O_158,N_19854,N_19676);
nand UO_159 (O_159,N_16591,N_17556);
nand UO_160 (O_160,N_16876,N_19312);
or UO_161 (O_161,N_15425,N_15249);
nand UO_162 (O_162,N_16059,N_17114);
nand UO_163 (O_163,N_18652,N_16873);
and UO_164 (O_164,N_15315,N_16183);
and UO_165 (O_165,N_19965,N_17261);
or UO_166 (O_166,N_17803,N_19718);
nand UO_167 (O_167,N_18484,N_19303);
nor UO_168 (O_168,N_17166,N_19109);
or UO_169 (O_169,N_19548,N_16020);
or UO_170 (O_170,N_19388,N_15611);
nor UO_171 (O_171,N_15196,N_17081);
nor UO_172 (O_172,N_16545,N_15194);
nand UO_173 (O_173,N_19957,N_16157);
xor UO_174 (O_174,N_19955,N_16387);
nor UO_175 (O_175,N_15947,N_19175);
nand UO_176 (O_176,N_15145,N_15497);
nand UO_177 (O_177,N_19785,N_15221);
xnor UO_178 (O_178,N_16822,N_16408);
and UO_179 (O_179,N_16462,N_16463);
nand UO_180 (O_180,N_16846,N_18441);
nor UO_181 (O_181,N_16507,N_19119);
nand UO_182 (O_182,N_18341,N_15864);
and UO_183 (O_183,N_16706,N_16672);
xnor UO_184 (O_184,N_15493,N_17171);
or UO_185 (O_185,N_19398,N_18663);
or UO_186 (O_186,N_15318,N_16690);
nand UO_187 (O_187,N_15162,N_17882);
and UO_188 (O_188,N_19982,N_15778);
nand UO_189 (O_189,N_15080,N_19899);
or UO_190 (O_190,N_18607,N_16521);
nand UO_191 (O_191,N_16658,N_19807);
and UO_192 (O_192,N_15985,N_19077);
xnor UO_193 (O_193,N_15870,N_17528);
nor UO_194 (O_194,N_17723,N_15164);
xor UO_195 (O_195,N_18163,N_17704);
or UO_196 (O_196,N_17522,N_19185);
nor UO_197 (O_197,N_19260,N_15905);
and UO_198 (O_198,N_15747,N_19100);
and UO_199 (O_199,N_15739,N_15442);
nand UO_200 (O_200,N_15924,N_18231);
nand UO_201 (O_201,N_18108,N_18478);
or UO_202 (O_202,N_19522,N_16513);
xor UO_203 (O_203,N_18085,N_17513);
xor UO_204 (O_204,N_17067,N_17079);
or UO_205 (O_205,N_15795,N_17233);
and UO_206 (O_206,N_19883,N_18670);
or UO_207 (O_207,N_15948,N_16512);
nor UO_208 (O_208,N_19057,N_16476);
and UO_209 (O_209,N_18621,N_19406);
and UO_210 (O_210,N_19428,N_15934);
and UO_211 (O_211,N_18964,N_16499);
nand UO_212 (O_212,N_17386,N_18318);
xnor UO_213 (O_213,N_17552,N_19072);
and UO_214 (O_214,N_18587,N_18872);
nand UO_215 (O_215,N_18299,N_16599);
or UO_216 (O_216,N_16838,N_18602);
and UO_217 (O_217,N_17226,N_16163);
nor UO_218 (O_218,N_17636,N_17933);
xor UO_219 (O_219,N_17444,N_17724);
or UO_220 (O_220,N_15876,N_19208);
and UO_221 (O_221,N_16234,N_19882);
xor UO_222 (O_222,N_15102,N_15895);
and UO_223 (O_223,N_19351,N_18149);
nand UO_224 (O_224,N_16009,N_15919);
and UO_225 (O_225,N_15393,N_17678);
or UO_226 (O_226,N_15369,N_15270);
nand UO_227 (O_227,N_15922,N_17328);
nand UO_228 (O_228,N_15129,N_15615);
nand UO_229 (O_229,N_18854,N_15660);
or UO_230 (O_230,N_16045,N_19652);
and UO_231 (O_231,N_18244,N_16531);
or UO_232 (O_232,N_17517,N_19219);
nor UO_233 (O_233,N_15681,N_15676);
or UO_234 (O_234,N_15940,N_17318);
and UO_235 (O_235,N_15853,N_15548);
nor UO_236 (O_236,N_16472,N_16501);
and UO_237 (O_237,N_15889,N_16042);
and UO_238 (O_238,N_17032,N_15251);
nor UO_239 (O_239,N_17639,N_15370);
or UO_240 (O_240,N_17946,N_17342);
or UO_241 (O_241,N_19371,N_17738);
and UO_242 (O_242,N_16899,N_17034);
and UO_243 (O_243,N_17985,N_18400);
nand UO_244 (O_244,N_18029,N_18850);
and UO_245 (O_245,N_18876,N_15451);
or UO_246 (O_246,N_17931,N_18295);
nand UO_247 (O_247,N_19875,N_16887);
nor UO_248 (O_248,N_17381,N_19284);
xnor UO_249 (O_249,N_16615,N_18827);
nand UO_250 (O_250,N_17742,N_18366);
nor UO_251 (O_251,N_18298,N_19707);
or UO_252 (O_252,N_19871,N_18503);
or UO_253 (O_253,N_17799,N_16038);
and UO_254 (O_254,N_17138,N_19941);
nor UO_255 (O_255,N_16711,N_18490);
nand UO_256 (O_256,N_17488,N_18397);
nand UO_257 (O_257,N_16431,N_17625);
nor UO_258 (O_258,N_15518,N_17841);
nor UO_259 (O_259,N_18459,N_15419);
nor UO_260 (O_260,N_18627,N_15205);
and UO_261 (O_261,N_15768,N_19649);
and UO_262 (O_262,N_17039,N_18903);
nor UO_263 (O_263,N_19654,N_16340);
and UO_264 (O_264,N_16919,N_18965);
nor UO_265 (O_265,N_19866,N_17217);
or UO_266 (O_266,N_15473,N_17133);
and UO_267 (O_267,N_15720,N_15568);
and UO_268 (O_268,N_19124,N_15628);
nor UO_269 (O_269,N_15844,N_19602);
nor UO_270 (O_270,N_16115,N_19639);
and UO_271 (O_271,N_18594,N_17770);
and UO_272 (O_272,N_17987,N_18378);
and UO_273 (O_273,N_19322,N_17581);
nor UO_274 (O_274,N_15028,N_17520);
and UO_275 (O_275,N_16016,N_19385);
or UO_276 (O_276,N_15295,N_18173);
or UO_277 (O_277,N_17241,N_19135);
nor UO_278 (O_278,N_17144,N_15043);
and UO_279 (O_279,N_16644,N_16160);
and UO_280 (O_280,N_18346,N_19058);
or UO_281 (O_281,N_18606,N_17110);
nor UO_282 (O_282,N_15290,N_16060);
or UO_283 (O_283,N_18937,N_16424);
or UO_284 (O_284,N_18189,N_18909);
nand UO_285 (O_285,N_17972,N_15647);
nor UO_286 (O_286,N_17685,N_16816);
nor UO_287 (O_287,N_15523,N_18062);
nand UO_288 (O_288,N_15161,N_16187);
and UO_289 (O_289,N_19047,N_16212);
or UO_290 (O_290,N_19715,N_18421);
or UO_291 (O_291,N_19706,N_18025);
xor UO_292 (O_292,N_15042,N_16568);
nor UO_293 (O_293,N_19802,N_16121);
or UO_294 (O_294,N_18286,N_19297);
or UO_295 (O_295,N_19926,N_17051);
and UO_296 (O_296,N_19818,N_15685);
or UO_297 (O_297,N_19958,N_17827);
and UO_298 (O_298,N_18464,N_17661);
xor UO_299 (O_299,N_15749,N_18177);
or UO_300 (O_300,N_17525,N_16525);
nor UO_301 (O_301,N_19222,N_19452);
or UO_302 (O_302,N_15967,N_16371);
or UO_303 (O_303,N_15731,N_15301);
or UO_304 (O_304,N_18784,N_15779);
nor UO_305 (O_305,N_16169,N_19780);
nor UO_306 (O_306,N_18593,N_18008);
or UO_307 (O_307,N_15391,N_19483);
and UO_308 (O_308,N_17997,N_15521);
nand UO_309 (O_309,N_19609,N_17240);
or UO_310 (O_310,N_15513,N_19979);
nor UO_311 (O_311,N_19186,N_17563);
xor UO_312 (O_312,N_16954,N_18772);
and UO_313 (O_313,N_16971,N_16627);
nor UO_314 (O_314,N_19325,N_16646);
or UO_315 (O_315,N_15132,N_18340);
nand UO_316 (O_316,N_17206,N_19973);
xnor UO_317 (O_317,N_17879,N_15535);
or UO_318 (O_318,N_15773,N_15276);
xnor UO_319 (O_319,N_15422,N_16692);
nor UO_320 (O_320,N_15597,N_17196);
and UO_321 (O_321,N_15756,N_17490);
nor UO_322 (O_322,N_16006,N_18385);
nor UO_323 (O_323,N_15605,N_15524);
nor UO_324 (O_324,N_17900,N_16732);
nand UO_325 (O_325,N_15530,N_17868);
nand UO_326 (O_326,N_16963,N_18691);
nor UO_327 (O_327,N_15849,N_16058);
nand UO_328 (O_328,N_15209,N_16455);
nand UO_329 (O_329,N_17376,N_18529);
nand UO_330 (O_330,N_18382,N_16540);
or UO_331 (O_331,N_16523,N_18091);
nand UO_332 (O_332,N_15296,N_15197);
and UO_333 (O_333,N_16186,N_19387);
and UO_334 (O_334,N_19352,N_17809);
or UO_335 (O_335,N_17960,N_18338);
and UO_336 (O_336,N_15593,N_18146);
or UO_337 (O_337,N_18960,N_16241);
nor UO_338 (O_338,N_18605,N_15434);
and UO_339 (O_339,N_16219,N_18610);
nor UO_340 (O_340,N_17185,N_18407);
nor UO_341 (O_341,N_17062,N_19220);
xnor UO_342 (O_342,N_16544,N_15661);
and UO_343 (O_343,N_16725,N_16301);
nor UO_344 (O_344,N_17251,N_16292);
nor UO_345 (O_345,N_15491,N_17084);
and UO_346 (O_346,N_16709,N_19085);
or UO_347 (O_347,N_19053,N_17843);
or UO_348 (O_348,N_19856,N_17693);
or UO_349 (O_349,N_18159,N_19797);
or UO_350 (O_350,N_19233,N_19468);
nor UO_351 (O_351,N_16328,N_18535);
xnor UO_352 (O_352,N_17808,N_15498);
nor UO_353 (O_353,N_19674,N_19632);
or UO_354 (O_354,N_18786,N_15536);
nor UO_355 (O_355,N_19678,N_16960);
nand UO_356 (O_356,N_18426,N_18682);
nor UO_357 (O_357,N_16638,N_18153);
or UO_358 (O_358,N_16685,N_18268);
or UO_359 (O_359,N_19365,N_19688);
or UO_360 (O_360,N_15514,N_15744);
and UO_361 (O_361,N_19310,N_19917);
and UO_362 (O_362,N_16450,N_17918);
nand UO_363 (O_363,N_19273,N_17794);
and UO_364 (O_364,N_18505,N_19145);
xor UO_365 (O_365,N_15317,N_17130);
and UO_366 (O_366,N_19240,N_15519);
or UO_367 (O_367,N_17375,N_17953);
nand UO_368 (O_368,N_17249,N_19616);
or UO_369 (O_369,N_16309,N_17224);
nand UO_370 (O_370,N_19537,N_16091);
or UO_371 (O_371,N_15014,N_18015);
nand UO_372 (O_372,N_18816,N_16430);
nor UO_373 (O_373,N_18465,N_16468);
nor UO_374 (O_374,N_17001,N_16316);
and UO_375 (O_375,N_19892,N_18413);
nor UO_376 (O_376,N_19939,N_16392);
nand UO_377 (O_377,N_15231,N_16594);
xnor UO_378 (O_378,N_17432,N_17650);
and UO_379 (O_379,N_18563,N_16319);
nand UO_380 (O_380,N_19140,N_15976);
and UO_381 (O_381,N_15850,N_16400);
nand UO_382 (O_382,N_19834,N_17006);
and UO_383 (O_383,N_15707,N_18046);
nand UO_384 (O_384,N_15193,N_15121);
nand UO_385 (O_385,N_16214,N_15623);
and UO_386 (O_386,N_15657,N_15721);
or UO_387 (O_387,N_18625,N_16660);
or UO_388 (O_388,N_19441,N_18929);
nor UO_389 (O_389,N_19378,N_16204);
xor UO_390 (O_390,N_17915,N_17305);
or UO_391 (O_391,N_15960,N_17621);
and UO_392 (O_392,N_19111,N_16659);
and UO_393 (O_393,N_15813,N_18281);
and UO_394 (O_394,N_17368,N_15856);
xnor UO_395 (O_395,N_15280,N_15846);
nand UO_396 (O_396,N_19677,N_16027);
or UO_397 (O_397,N_15199,N_15291);
or UO_398 (O_398,N_15026,N_15163);
nand UO_399 (O_399,N_17851,N_18186);
nor UO_400 (O_400,N_19493,N_19154);
xnor UO_401 (O_401,N_16662,N_19811);
and UO_402 (O_402,N_15949,N_17292);
nor UO_403 (O_403,N_18527,N_18998);
nor UO_404 (O_404,N_16274,N_19712);
and UO_405 (O_405,N_19268,N_16588);
nor UO_406 (O_406,N_19092,N_15150);
nand UO_407 (O_407,N_17994,N_17024);
and UO_408 (O_408,N_19510,N_17740);
nand UO_409 (O_409,N_17792,N_16067);
and UO_410 (O_410,N_18679,N_15892);
nor UO_411 (O_411,N_16518,N_18637);
nor UO_412 (O_412,N_18399,N_18684);
or UO_413 (O_413,N_15557,N_17690);
nand UO_414 (O_414,N_17887,N_16571);
xor UO_415 (O_415,N_18302,N_17390);
nand UO_416 (O_416,N_18845,N_15978);
nand UO_417 (O_417,N_19102,N_18056);
and UO_418 (O_418,N_16687,N_18775);
nand UO_419 (O_419,N_16098,N_18211);
or UO_420 (O_420,N_18865,N_16191);
nor UO_421 (O_421,N_17603,N_17478);
or UO_422 (O_422,N_16554,N_15839);
and UO_423 (O_423,N_19429,N_19855);
or UO_424 (O_424,N_15283,N_18925);
nor UO_425 (O_425,N_17268,N_17939);
nand UO_426 (O_426,N_17486,N_15835);
nand UO_427 (O_427,N_18991,N_17036);
or UO_428 (O_428,N_19424,N_15805);
nor UO_429 (O_429,N_19132,N_17949);
nand UO_430 (O_430,N_19164,N_17545);
nand UO_431 (O_431,N_15979,N_16557);
nor UO_432 (O_432,N_15137,N_18512);
or UO_433 (O_433,N_16859,N_19859);
xor UO_434 (O_434,N_16326,N_17755);
nor UO_435 (O_435,N_18516,N_17820);
nor UO_436 (O_436,N_19874,N_18181);
nand UO_437 (O_437,N_15929,N_17052);
nor UO_438 (O_438,N_18183,N_16852);
and UO_439 (O_439,N_15148,N_19971);
or UO_440 (O_440,N_15981,N_18248);
or UO_441 (O_441,N_19471,N_16368);
or UO_442 (O_442,N_16425,N_17637);
xor UO_443 (O_443,N_15138,N_16596);
xor UO_444 (O_444,N_15737,N_17529);
nand UO_445 (O_445,N_17952,N_15560);
nand UO_446 (O_446,N_19809,N_16350);
and UO_447 (O_447,N_18258,N_17439);
or UO_448 (O_448,N_17413,N_19760);
xnor UO_449 (O_449,N_19497,N_15176);
or UO_450 (O_450,N_16381,N_17445);
xnor UO_451 (O_451,N_15117,N_18723);
and UO_452 (O_452,N_19403,N_15174);
xnor UO_453 (O_453,N_15995,N_15011);
and UO_454 (O_454,N_16741,N_16825);
or UO_455 (O_455,N_18436,N_18238);
nor UO_456 (O_456,N_15050,N_18567);
and UO_457 (O_457,N_19836,N_16307);
nand UO_458 (O_458,N_18113,N_15622);
nor UO_459 (O_459,N_17274,N_19435);
or UO_460 (O_460,N_17613,N_18841);
and UO_461 (O_461,N_16473,N_17569);
nand UO_462 (O_462,N_17726,N_18790);
and UO_463 (O_463,N_18350,N_17254);
and UO_464 (O_464,N_16103,N_16797);
or UO_465 (O_465,N_18881,N_19585);
xor UO_466 (O_466,N_17287,N_16289);
xor UO_467 (O_467,N_15468,N_19679);
or UO_468 (O_468,N_19838,N_15165);
xnor UO_469 (O_469,N_16395,N_15499);
xnor UO_470 (O_470,N_15687,N_19901);
or UO_471 (O_471,N_15294,N_18351);
nand UO_472 (O_472,N_15341,N_19949);
or UO_473 (O_473,N_18020,N_19642);
nor UO_474 (O_474,N_17824,N_16656);
nor UO_475 (O_475,N_18840,N_17134);
and UO_476 (O_476,N_15377,N_16978);
or UO_477 (O_477,N_15006,N_18767);
nand UO_478 (O_478,N_17551,N_15952);
nor UO_479 (O_479,N_17911,N_18393);
or UO_480 (O_480,N_19717,N_17168);
or UO_481 (O_481,N_15845,N_19749);
or UO_482 (O_482,N_17424,N_17408);
nand UO_483 (O_483,N_17605,N_19501);
nand UO_484 (O_484,N_16586,N_15246);
or UO_485 (O_485,N_15910,N_15217);
nor UO_486 (O_486,N_15658,N_15486);
xor UO_487 (O_487,N_15307,N_19568);
xnor UO_488 (O_488,N_19350,N_15269);
nor UO_489 (O_489,N_15760,N_17201);
and UO_490 (O_490,N_15801,N_19120);
or UO_491 (O_491,N_15938,N_17627);
nor UO_492 (O_492,N_18126,N_16920);
xnor UO_493 (O_493,N_15860,N_15420);
or UO_494 (O_494,N_18481,N_18751);
or UO_495 (O_495,N_19486,N_15527);
or UO_496 (O_496,N_15001,N_16161);
and UO_497 (O_497,N_18657,N_17256);
xnor UO_498 (O_498,N_19752,N_19755);
xor UO_499 (O_499,N_18349,N_15030);
nand UO_500 (O_500,N_15668,N_17363);
nand UO_501 (O_501,N_17974,N_16198);
nand UO_502 (O_502,N_19198,N_16769);
or UO_503 (O_503,N_17301,N_19581);
nand UO_504 (O_504,N_19230,N_18038);
nor UO_505 (O_505,N_18463,N_16404);
nor UO_506 (O_506,N_17326,N_17574);
and UO_507 (O_507,N_19160,N_16994);
and UO_508 (O_508,N_19239,N_19014);
nand UO_509 (O_509,N_18860,N_19205);
nand UO_510 (O_510,N_18285,N_16700);
nand UO_511 (O_511,N_16771,N_16213);
nor UO_512 (O_512,N_16321,N_18107);
nand UO_513 (O_513,N_17165,N_17620);
nand UO_514 (O_514,N_18158,N_16434);
nor UO_515 (O_515,N_19808,N_19031);
or UO_516 (O_516,N_15828,N_19149);
xnor UO_517 (O_517,N_17875,N_17718);
xnor UO_518 (O_518,N_17589,N_19075);
nor UO_519 (O_519,N_15201,N_15909);
and UO_520 (O_520,N_15114,N_19324);
nor UO_521 (O_521,N_16634,N_17054);
nor UO_522 (O_522,N_17664,N_16753);
nand UO_523 (O_523,N_15103,N_18104);
xnor UO_524 (O_524,N_17435,N_17989);
or UO_525 (O_525,N_19863,N_18092);
or UO_526 (O_526,N_17502,N_15215);
nand UO_527 (O_527,N_15070,N_16975);
or UO_528 (O_528,N_16389,N_18249);
or UO_529 (O_529,N_17239,N_16666);
and UO_530 (O_530,N_19975,N_18722);
nand UO_531 (O_531,N_16017,N_16010);
nor UO_532 (O_532,N_16829,N_18916);
and UO_533 (O_533,N_15184,N_17056);
and UO_534 (O_534,N_15621,N_19697);
or UO_535 (O_535,N_17163,N_18076);
nand UO_536 (O_536,N_17750,N_16880);
nand UO_537 (O_537,N_18669,N_18668);
xor UO_538 (O_538,N_17208,N_19728);
nand UO_539 (O_539,N_16379,N_15454);
or UO_540 (O_540,N_18209,N_19383);
nand UO_541 (O_541,N_17854,N_17072);
xor UO_542 (O_542,N_19173,N_15840);
nor UO_543 (O_543,N_18147,N_18331);
xnor UO_544 (O_544,N_18498,N_16299);
xnor UO_545 (O_545,N_18733,N_18510);
nor UO_546 (O_546,N_18761,N_16775);
nor UO_547 (O_547,N_17370,N_19594);
and UO_548 (O_548,N_18940,N_19264);
and UO_549 (O_549,N_18405,N_16719);
xnor UO_550 (O_550,N_17607,N_19912);
or UO_551 (O_551,N_15577,N_17920);
and UO_552 (O_552,N_19474,N_18748);
xnor UO_553 (O_553,N_18986,N_17066);
or UO_554 (O_554,N_15616,N_15427);
nor UO_555 (O_555,N_19333,N_15515);
or UO_556 (O_556,N_17469,N_15256);
or UO_557 (O_557,N_16923,N_16718);
and UO_558 (O_558,N_16765,N_16745);
nor UO_559 (O_559,N_18043,N_17757);
or UO_560 (O_560,N_19577,N_19083);
and UO_561 (O_561,N_15695,N_16867);
or UO_562 (O_562,N_16064,N_18264);
or UO_563 (O_563,N_19007,N_15918);
nor UO_564 (O_564,N_15677,N_17540);
or UO_565 (O_565,N_16273,N_16674);
nor UO_566 (O_566,N_17463,N_17956);
nor UO_567 (O_567,N_17756,N_15466);
nand UO_568 (O_568,N_18650,N_18404);
nor UO_569 (O_569,N_15858,N_17711);
nand UO_570 (O_570,N_16364,N_16005);
or UO_571 (O_571,N_17819,N_16014);
or UO_572 (O_572,N_19504,N_17069);
xnor UO_573 (O_573,N_19684,N_15097);
and UO_574 (O_574,N_18501,N_18167);
or UO_575 (O_575,N_17106,N_19106);
nand UO_576 (O_576,N_18868,N_17341);
or UO_577 (O_577,N_17074,N_15599);
xnor UO_578 (O_578,N_19595,N_19918);
nor UO_579 (O_579,N_16497,N_16509);
nand UO_580 (O_580,N_16226,N_15418);
nand UO_581 (O_581,N_19263,N_16135);
nor UO_582 (O_582,N_15550,N_16981);
or UO_583 (O_583,N_17720,N_17560);
nand UO_584 (O_584,N_15285,N_18475);
nor UO_585 (O_585,N_19399,N_17132);
nor UO_586 (O_586,N_15262,N_19362);
or UO_587 (O_587,N_18419,N_18217);
and UO_588 (O_588,N_19232,N_15358);
nand UO_589 (O_589,N_18275,N_19757);
nor UO_590 (O_590,N_17591,N_18757);
and UO_591 (O_591,N_15426,N_17571);
nand UO_592 (O_592,N_15832,N_18476);
nor UO_593 (O_593,N_19870,N_15338);
and UO_594 (O_594,N_17406,N_18852);
nor UO_595 (O_595,N_17020,N_17771);
nor UO_596 (O_596,N_17505,N_19888);
nor UO_597 (O_597,N_15202,N_17282);
nor UO_598 (O_598,N_15694,N_15182);
and UO_599 (O_599,N_17706,N_19550);
and UO_600 (O_600,N_17991,N_19721);
xor UO_601 (O_601,N_19987,N_15712);
or UO_602 (O_602,N_19125,N_18164);
nand UO_603 (O_603,N_18622,N_15153);
or UO_604 (O_604,N_18253,N_16766);
nand UO_605 (O_605,N_15093,N_15287);
and UO_606 (O_606,N_17500,N_16367);
nor UO_607 (O_607,N_18918,N_15408);
and UO_608 (O_608,N_16788,N_15396);
or UO_609 (O_609,N_18202,N_17684);
or UO_610 (O_610,N_19906,N_19691);
and UO_611 (O_611,N_17371,N_18383);
and UO_612 (O_612,N_15987,N_17713);
nor UO_613 (O_613,N_17472,N_16013);
nand UO_614 (O_614,N_18648,N_18863);
nor UO_615 (O_615,N_17147,N_15808);
nand UO_616 (O_616,N_19037,N_16134);
and UO_617 (O_617,N_16088,N_17531);
nand UO_618 (O_618,N_15053,N_17818);
nor UO_619 (O_619,N_19894,N_19521);
xor UO_620 (O_620,N_18178,N_15797);
or UO_621 (O_621,N_15461,N_18749);
xnor UO_622 (O_622,N_19215,N_18674);
nor UO_623 (O_623,N_19361,N_19934);
or UO_624 (O_624,N_17362,N_16385);
nor UO_625 (O_625,N_18993,N_19207);
or UO_626 (O_626,N_16021,N_18132);
or UO_627 (O_627,N_17908,N_15482);
or UO_628 (O_628,N_19159,N_17884);
nand UO_629 (O_629,N_15169,N_15401);
and UO_630 (O_630,N_19323,N_18572);
or UO_631 (O_631,N_17895,N_18196);
and UO_632 (O_632,N_19475,N_19465);
or UO_633 (O_633,N_16500,N_17252);
or UO_634 (O_634,N_16739,N_17060);
nand UO_635 (O_635,N_16222,N_18241);
nor UO_636 (O_636,N_17099,N_15941);
nand UO_637 (O_637,N_16791,N_17903);
nand UO_638 (O_638,N_15613,N_17783);
or UO_639 (O_639,N_17981,N_18787);
or UO_640 (O_640,N_18212,N_16870);
or UO_641 (O_641,N_18844,N_19443);
or UO_642 (O_642,N_17187,N_15820);
xor UO_643 (O_643,N_17592,N_15073);
or UO_644 (O_644,N_18859,N_18348);
and UO_645 (O_645,N_16451,N_18080);
nand UO_646 (O_646,N_16171,N_19588);
or UO_647 (O_647,N_15409,N_15319);
nand UO_648 (O_648,N_18039,N_15818);
xnor UO_649 (O_649,N_18078,N_17068);
or UO_650 (O_650,N_17098,N_15310);
nor UO_651 (O_651,N_18396,N_18829);
xor UO_652 (O_652,N_18583,N_19601);
nor UO_653 (O_653,N_17683,N_15554);
or UO_654 (O_654,N_17446,N_19065);
nand UO_655 (O_655,N_19731,N_16881);
nor UO_656 (O_656,N_18855,N_16426);
nand UO_657 (O_657,N_19449,N_18667);
nand UO_658 (O_658,N_16914,N_16137);
nand UO_659 (O_659,N_15303,N_17480);
xnor UO_660 (O_660,N_18087,N_17299);
nor UO_661 (O_661,N_17387,N_18288);
nand UO_662 (O_662,N_16696,N_16877);
nand UO_663 (O_663,N_19166,N_16339);
and UO_664 (O_664,N_16550,N_19835);
or UO_665 (O_665,N_18409,N_19898);
nor UO_666 (O_666,N_18195,N_17336);
nand UO_667 (O_667,N_18276,N_15716);
nand UO_668 (O_668,N_19402,N_18105);
and UO_669 (O_669,N_18966,N_15826);
or UO_670 (O_670,N_15516,N_16229);
and UO_671 (O_671,N_15352,N_16823);
nor UO_672 (O_672,N_19082,N_17532);
nor UO_673 (O_673,N_16976,N_18592);
and UO_674 (O_674,N_16536,N_17668);
nor UO_675 (O_675,N_16872,N_16728);
and UO_676 (O_676,N_19038,N_15578);
nor UO_677 (O_677,N_18458,N_17448);
nor UO_678 (O_678,N_17385,N_19942);
xor UO_679 (O_679,N_16720,N_16396);
or UO_680 (O_680,N_15717,N_17585);
or UO_681 (O_681,N_19784,N_15172);
or UO_682 (O_682,N_16835,N_17283);
nand UO_683 (O_683,N_16190,N_18913);
nand UO_684 (O_684,N_16917,N_17638);
and UO_685 (O_685,N_18278,N_17536);
nor UO_686 (O_686,N_19187,N_18234);
xnor UO_687 (O_687,N_17675,N_19622);
nor UO_688 (O_688,N_15379,N_16635);
and UO_689 (O_689,N_17247,N_15387);
nand UO_690 (O_690,N_17507,N_16441);
and UO_691 (O_691,N_18321,N_15500);
nand UO_692 (O_692,N_15843,N_18023);
nand UO_693 (O_693,N_15821,N_15090);
nor UO_694 (O_694,N_16148,N_15881);
nor UO_695 (O_695,N_18701,N_16294);
nor UO_696 (O_696,N_15106,N_19454);
nand UO_697 (O_697,N_15774,N_15783);
and UO_698 (O_698,N_16107,N_17998);
or UO_699 (O_699,N_16200,N_15733);
nor UO_700 (O_700,N_15738,N_16388);
nor UO_701 (O_701,N_17481,N_18438);
or UO_702 (O_702,N_15973,N_17654);
nand UO_703 (O_703,N_17954,N_16141);
nor UO_704 (O_704,N_18608,N_19578);
or UO_705 (O_705,N_17026,N_15241);
and UO_706 (O_706,N_19758,N_15204);
xnor UO_707 (O_707,N_15356,N_15052);
nand UO_708 (O_708,N_18537,N_19305);
xnor UO_709 (O_709,N_19513,N_15018);
xnor UO_710 (O_710,N_17351,N_18127);
and UO_711 (O_711,N_16584,N_19913);
and UO_712 (O_712,N_18536,N_15983);
xnor UO_713 (O_713,N_17951,N_19009);
and UO_714 (O_714,N_19314,N_16290);
nor UO_715 (O_715,N_18386,N_15888);
nand UO_716 (O_716,N_15305,N_15388);
or UO_717 (O_717,N_16109,N_15098);
nor UO_718 (O_718,N_15920,N_18204);
and UO_719 (O_719,N_16030,N_19617);
nor UO_720 (O_720,N_17788,N_18362);
nand UO_721 (O_721,N_15447,N_16344);
xor UO_722 (O_722,N_18461,N_15289);
nor UO_723 (O_723,N_17966,N_17372);
or UO_724 (O_724,N_18812,N_16142);
or UO_725 (O_725,N_15430,N_16743);
nand UO_726 (O_726,N_17590,N_15619);
nor UO_727 (O_727,N_16490,N_19153);
nor UO_728 (O_728,N_19703,N_18097);
or UO_729 (O_729,N_16131,N_17304);
nor UO_730 (O_730,N_17611,N_18815);
or UO_731 (O_731,N_19517,N_16435);
nor UO_732 (O_732,N_19282,N_19804);
xnor UO_733 (O_733,N_19410,N_16906);
nor UO_734 (O_734,N_18358,N_15371);
and UO_735 (O_735,N_16514,N_16491);
and UO_736 (O_736,N_15107,N_17291);
nand UO_737 (O_737,N_16601,N_16158);
nand UO_738 (O_738,N_16149,N_16298);
nor UO_739 (O_739,N_17673,N_18497);
xor UO_740 (O_740,N_19747,N_17129);
nand UO_741 (O_741,N_18361,N_19060);
nand UO_742 (O_742,N_18151,N_15384);
nand UO_743 (O_743,N_15882,N_17225);
and UO_744 (O_744,N_16011,N_19234);
nor UO_745 (O_745,N_16145,N_18706);
xor UO_746 (O_746,N_19086,N_19028);
nor UO_747 (O_747,N_19401,N_17877);
or UO_748 (O_748,N_15261,N_18553);
or UO_749 (O_749,N_18365,N_18979);
nor UO_750 (O_750,N_19347,N_16529);
or UO_751 (O_751,N_19156,N_17979);
nand UO_752 (O_752,N_19141,N_16174);
or UO_753 (O_753,N_15049,N_15742);
and UO_754 (O_754,N_17193,N_15782);
nand UO_755 (O_755,N_17703,N_18969);
and UO_756 (O_756,N_19089,N_17035);
nand UO_757 (O_757,N_16244,N_15453);
or UO_758 (O_758,N_15133,N_16933);
nor UO_759 (O_759,N_19565,N_17999);
nor UO_760 (O_760,N_18205,N_18216);
or UO_761 (O_761,N_19848,N_17046);
or UO_762 (O_762,N_19536,N_16247);
nand UO_763 (O_763,N_19985,N_19938);
nand UO_764 (O_764,N_18737,N_18686);
and UO_765 (O_765,N_15110,N_16236);
nor UO_766 (O_766,N_18811,N_19342);
xor UO_767 (O_767,N_17045,N_16772);
nor UO_768 (O_768,N_17198,N_17250);
or UO_769 (O_769,N_15373,N_19190);
nand UO_770 (O_770,N_15708,N_18388);
or UO_771 (O_771,N_16549,N_16256);
xnor UO_772 (O_772,N_16543,N_18473);
and UO_773 (O_773,N_18373,N_16844);
nor UO_774 (O_774,N_19743,N_18797);
nor UO_775 (O_775,N_17656,N_17941);
nor UO_776 (O_776,N_17121,N_15361);
nor UO_777 (O_777,N_18839,N_17753);
nor UO_778 (O_778,N_17159,N_19646);
or UO_779 (O_779,N_17317,N_17452);
nand UO_780 (O_780,N_17038,N_17366);
or UO_781 (O_781,N_17412,N_15609);
or UO_782 (O_782,N_15438,N_19641);
and UO_783 (O_783,N_19908,N_17963);
or UO_784 (O_784,N_17245,N_18005);
nor UO_785 (O_785,N_19608,N_17265);
nor UO_786 (O_786,N_18316,N_15435);
nand UO_787 (O_787,N_17857,N_16414);
or UO_788 (O_788,N_17393,N_18034);
or UO_789 (O_789,N_15206,N_18905);
nand UO_790 (O_790,N_15732,N_16248);
and UO_791 (O_791,N_16285,N_19904);
nand UO_792 (O_792,N_15012,N_15395);
or UO_793 (O_793,N_19636,N_18626);
nor UO_794 (O_794,N_16237,N_17961);
xor UO_795 (O_795,N_16188,N_15139);
nor UO_796 (O_796,N_18301,N_19249);
nand UO_797 (O_797,N_17804,N_19408);
nand UO_798 (O_798,N_16304,N_19194);
nor UO_799 (O_799,N_17930,N_15259);
or UO_800 (O_800,N_16726,N_19852);
or UO_801 (O_801,N_15456,N_16403);
or UO_802 (O_802,N_17150,N_16034);
or UO_803 (O_803,N_17995,N_18891);
nand UO_804 (O_804,N_15381,N_15471);
or UO_805 (O_805,N_16488,N_17735);
nand UO_806 (O_806,N_19461,N_19455);
nor UO_807 (O_807,N_15044,N_18014);
and UO_808 (O_808,N_15542,N_17641);
or UO_809 (O_809,N_18500,N_16902);
and UO_810 (O_810,N_19191,N_15640);
and UO_811 (O_811,N_17323,N_18462);
or UO_812 (O_812,N_17440,N_19242);
nor UO_813 (O_813,N_15375,N_17028);
and UO_814 (O_814,N_18242,N_18449);
and UO_815 (O_815,N_18934,N_15595);
or UO_816 (O_816,N_18735,N_17324);
xnor UO_817 (O_817,N_17349,N_15281);
or UO_818 (O_818,N_16173,N_15309);
nand UO_819 (O_819,N_15101,N_19337);
nor UO_820 (O_820,N_18193,N_18696);
nor UO_821 (O_821,N_17761,N_15023);
or UO_822 (O_822,N_15702,N_19946);
nor UO_823 (O_823,N_16546,N_19393);
nor UO_824 (O_824,N_18339,N_17117);
nand UO_825 (O_825,N_16922,N_18817);
xor UO_826 (O_826,N_16159,N_19573);
or UO_827 (O_827,N_17806,N_18644);
and UO_828 (O_828,N_19488,N_16773);
nor UO_829 (O_829,N_17572,N_18398);
or UO_830 (O_830,N_18522,N_18374);
xnor UO_831 (O_831,N_18044,N_17403);
and UO_832 (O_832,N_17727,N_15766);
and UO_833 (O_833,N_15762,N_17511);
and UO_834 (O_834,N_19627,N_19287);
nor UO_835 (O_835,N_16516,N_15549);
and UO_836 (O_836,N_19063,N_19332);
and UO_837 (O_837,N_18642,N_17310);
nand UO_838 (O_838,N_19800,N_16445);
and UO_839 (O_839,N_18886,N_16461);
and UO_840 (O_840,N_15054,N_17826);
xor UO_841 (O_841,N_19340,N_16792);
or UO_842 (O_842,N_19700,N_17805);
and UO_843 (O_843,N_19621,N_16801);
and UO_844 (O_844,N_16813,N_18628);
nor UO_845 (O_845,N_17758,N_15581);
or UO_846 (O_846,N_17815,N_17680);
or UO_847 (O_847,N_16866,N_15741);
nor UO_848 (O_848,N_16903,N_19651);
and UO_849 (O_849,N_18170,N_16761);
or UO_850 (O_850,N_19777,N_16998);
and UO_851 (O_851,N_19551,N_17976);
nor UO_852 (O_852,N_17610,N_19152);
nand UO_853 (O_853,N_16080,N_17978);
or UO_854 (O_854,N_18304,N_18513);
nand UO_855 (O_855,N_16506,N_17033);
nand UO_856 (O_856,N_16827,N_18615);
or UO_857 (O_857,N_19887,N_17148);
nor UO_858 (O_858,N_16444,N_19224);
or UO_859 (O_859,N_16924,N_19231);
or UO_860 (O_860,N_17322,N_15538);
or UO_861 (O_861,N_17616,N_16483);
and UO_862 (O_862,N_16311,N_15279);
nor UO_863 (O_863,N_19583,N_18920);
and UO_864 (O_864,N_15293,N_16086);
nor UO_865 (O_865,N_16802,N_15815);
or UO_866 (O_866,N_17498,N_16151);
nor UO_867 (O_867,N_18208,N_17280);
nand UO_868 (O_868,N_16900,N_18831);
and UO_869 (O_869,N_16798,N_17797);
and UO_870 (O_870,N_17319,N_19307);
and UO_871 (O_871,N_19511,N_16327);
nand UO_872 (O_872,N_17747,N_18114);
and UO_873 (O_873,N_17389,N_18310);
nor UO_874 (O_874,N_19543,N_17180);
nor UO_875 (O_875,N_16679,N_18342);
and UO_876 (O_876,N_18324,N_16032);
and UO_877 (O_877,N_15806,N_17583);
and UO_878 (O_878,N_19801,N_19661);
nor UO_879 (O_879,N_19004,N_17044);
or UO_880 (O_880,N_19034,N_18922);
or UO_881 (O_881,N_17344,N_17210);
or UO_882 (O_882,N_15669,N_15033);
or UO_883 (O_883,N_16410,N_19480);
nand UO_884 (O_884,N_18542,N_16028);
and UO_885 (O_885,N_17449,N_15796);
and UO_886 (O_886,N_18257,N_15158);
nand UO_887 (O_887,N_17160,N_18071);
and UO_888 (O_888,N_18942,N_17721);
or UO_889 (O_889,N_19528,N_15417);
or UO_890 (O_890,N_15005,N_16375);
or UO_891 (O_891,N_16853,N_18272);
xnor UO_892 (O_892,N_18992,N_19623);
and UO_893 (O_893,N_15208,N_19318);
or UO_894 (O_894,N_17442,N_16480);
and UO_895 (O_895,N_17212,N_19246);
nand UO_896 (O_896,N_19567,N_15617);
xnor UO_897 (O_897,N_18215,N_19634);
and UO_898 (O_898,N_19861,N_18004);
nand UO_899 (O_899,N_15900,N_19359);
nor UO_900 (O_900,N_18243,N_19235);
and UO_901 (O_901,N_18744,N_17688);
and UO_902 (O_902,N_18717,N_16632);
nor UO_903 (O_903,N_16969,N_18832);
or UO_904 (O_904,N_19670,N_18889);
xnor UO_905 (O_905,N_17913,N_18836);
or UO_906 (O_906,N_19538,N_16023);
nor UO_907 (O_907,N_19795,N_18676);
or UO_908 (O_908,N_16988,N_19236);
or UO_909 (O_909,N_17021,N_17215);
nor UO_910 (O_910,N_18957,N_18824);
nand UO_911 (O_911,N_16552,N_15936);
or UO_912 (O_912,N_16678,N_15351);
and UO_913 (O_913,N_18368,N_17156);
and UO_914 (O_914,N_17888,N_18791);
nor UO_915 (O_915,N_19256,N_18948);
nand UO_916 (O_916,N_17059,N_19150);
nand UO_917 (O_917,N_17306,N_17227);
xnor UO_918 (O_918,N_15735,N_16090);
and UO_919 (O_919,N_16329,N_17179);
and UO_920 (O_920,N_15684,N_18552);
nor UO_921 (O_921,N_15745,N_19555);
nor UO_922 (O_922,N_16893,N_18814);
nor UO_923 (O_923,N_19881,N_16228);
xnor UO_924 (O_924,N_16879,N_18511);
xnor UO_925 (O_925,N_16053,N_19788);
and UO_926 (O_926,N_19540,N_19139);
and UO_927 (O_927,N_16948,N_16493);
xnor UO_928 (O_928,N_19115,N_15638);
or UO_929 (O_929,N_17969,N_17694);
and UO_930 (O_930,N_17003,N_16111);
and UO_931 (O_931,N_19559,N_16555);
nand UO_932 (O_932,N_18624,N_18054);
xnor UO_933 (O_933,N_16087,N_17510);
nand UO_934 (O_934,N_16812,N_17766);
nor UO_935 (O_935,N_16310,N_17491);
and UO_936 (O_936,N_18418,N_17262);
and UO_937 (O_937,N_16755,N_19659);
or UO_938 (O_938,N_17228,N_19737);
nand UO_939 (O_939,N_15725,N_18308);
or UO_940 (O_940,N_18466,N_17634);
or UO_941 (O_941,N_16708,N_17615);
nand UO_942 (O_942,N_18539,N_16001);
or UO_943 (O_943,N_15402,N_17267);
or UO_944 (O_944,N_17016,N_17234);
nand UO_945 (O_945,N_17496,N_18103);
or UO_946 (O_946,N_18422,N_18277);
nand UO_947 (O_947,N_15330,N_16856);
and UO_948 (O_948,N_15944,N_18967);
or UO_949 (O_949,N_19998,N_15896);
nand UO_950 (O_950,N_17730,N_17460);
nor UO_951 (O_951,N_16947,N_17834);
xnor UO_952 (O_952,N_17512,N_16225);
and UO_953 (O_953,N_17473,N_15673);
and UO_954 (O_954,N_15879,N_18156);
nand UO_955 (O_955,N_19210,N_18760);
nand UO_956 (O_956,N_17565,N_15181);
or UO_957 (O_957,N_15916,N_15982);
or UO_958 (O_958,N_15666,N_16181);
nor UO_959 (O_959,N_17521,N_17925);
or UO_960 (O_960,N_17373,N_19631);
nor UO_961 (O_961,N_19572,N_17898);
nand UO_962 (O_962,N_18861,N_19593);
nand UO_963 (O_963,N_17137,N_15061);
and UO_964 (O_964,N_16713,N_19791);
nand UO_965 (O_965,N_16478,N_15576);
xor UO_966 (O_966,N_15841,N_16336);
nor UO_967 (O_967,N_17082,N_18982);
or UO_968 (O_968,N_18525,N_19722);
nand UO_969 (O_969,N_15155,N_17142);
nand UO_970 (O_970,N_18976,N_18947);
xor UO_971 (O_971,N_17343,N_16282);
and UO_972 (O_972,N_18515,N_16730);
xor UO_973 (O_973,N_18225,N_18566);
nor UO_974 (O_974,N_15357,N_17733);
and UO_975 (O_975,N_19733,N_19772);
nor UO_976 (O_976,N_19790,N_18743);
nor UO_977 (O_977,N_15112,N_15227);
nor UO_978 (O_978,N_15955,N_16442);
or UO_979 (O_979,N_18541,N_18908);
nand UO_980 (O_980,N_18131,N_19999);
nor UO_981 (O_981,N_15131,N_15335);
nor UO_982 (O_982,N_15772,N_16936);
nand UO_983 (O_983,N_16650,N_15974);
nand UO_984 (O_984,N_15816,N_17313);
and UO_985 (O_985,N_19561,N_19579);
or UO_986 (O_986,N_17128,N_15533);
nor UO_987 (O_987,N_15068,N_15496);
nor UO_988 (O_988,N_17853,N_17923);
and UO_989 (O_989,N_16456,N_16636);
nor UO_990 (O_990,N_18150,N_18089);
and UO_991 (O_991,N_18864,N_18065);
nor UO_992 (O_992,N_17764,N_15598);
nor UO_993 (O_993,N_17734,N_15273);
nor UO_994 (O_994,N_17300,N_18381);
and UO_995 (O_995,N_17027,N_15618);
or UO_996 (O_996,N_18336,N_16937);
nor UO_997 (O_997,N_18756,N_19052);
nand UO_998 (O_998,N_15629,N_16055);
xnor UO_999 (O_999,N_15233,N_17296);
and UO_1000 (O_1000,N_19886,N_18142);
nor UO_1001 (O_1001,N_16245,N_18818);
and UO_1002 (O_1002,N_16794,N_16729);
and UO_1003 (O_1003,N_15789,N_18896);
xor UO_1004 (O_1004,N_19490,N_15585);
or UO_1005 (O_1005,N_15428,N_18379);
and UO_1006 (O_1006,N_16052,N_17582);
nand UO_1007 (O_1007,N_18237,N_17852);
xnor UO_1008 (O_1008,N_15728,N_15062);
nand UO_1009 (O_1009,N_16063,N_16901);
nand UO_1010 (O_1010,N_15047,N_19381);
nor UO_1011 (O_1011,N_17484,N_17314);
nor UO_1012 (O_1012,N_15091,N_16556);
or UO_1013 (O_1013,N_19924,N_19087);
nor UO_1014 (O_1014,N_18770,N_19556);
nor UO_1015 (O_1015,N_18997,N_17232);
nand UO_1016 (O_1016,N_18483,N_19104);
nor UO_1017 (O_1017,N_15706,N_15656);
and UO_1018 (O_1018,N_16915,N_15411);
and UO_1019 (O_1019,N_16637,N_16166);
nand UO_1020 (O_1020,N_16318,N_19315);
or UO_1021 (O_1021,N_17379,N_18582);
nor UO_1022 (O_1022,N_15862,N_17698);
or UO_1023 (O_1023,N_19013,N_16830);
or UO_1024 (O_1024,N_19614,N_17643);
nor UO_1025 (O_1025,N_17575,N_16616);
and UO_1026 (O_1026,N_16789,N_15997);
nand UO_1027 (O_1027,N_18213,N_18394);
nor UO_1028 (O_1028,N_16302,N_18785);
or UO_1029 (O_1029,N_16966,N_16215);
and UO_1030 (O_1030,N_16548,N_17508);
and UO_1031 (O_1031,N_18402,N_15013);
nor UO_1032 (O_1032,N_19327,N_19740);
or UO_1033 (O_1033,N_17599,N_17492);
and UO_1034 (O_1034,N_15171,N_18911);
or UO_1035 (O_1035,N_16860,N_16639);
xnor UO_1036 (O_1036,N_19262,N_19719);
or UO_1037 (O_1037,N_19162,N_18945);
and UO_1038 (O_1038,N_17149,N_15002);
and UO_1039 (O_1039,N_16749,N_16044);
nand UO_1040 (O_1040,N_17327,N_18262);
or UO_1041 (O_1041,N_18221,N_19151);
xnor UO_1042 (O_1042,N_19050,N_19766);
nand UO_1043 (O_1043,N_19062,N_17272);
and UO_1044 (O_1044,N_19961,N_15902);
or UO_1045 (O_1045,N_18480,N_18470);
or UO_1046 (O_1046,N_17186,N_17752);
or UO_1047 (O_1047,N_15320,N_19890);
or UO_1048 (O_1048,N_15300,N_18878);
or UO_1049 (O_1049,N_18254,N_15614);
nand UO_1050 (O_1050,N_15195,N_17333);
nor UO_1051 (O_1051,N_19366,N_16515);
and UO_1052 (O_1052,N_19181,N_19499);
nand UO_1053 (O_1053,N_18526,N_16858);
and UO_1054 (O_1054,N_17671,N_19586);
nand UO_1055 (O_1055,N_15159,N_16626);
or UO_1056 (O_1056,N_16073,N_18042);
and UO_1057 (O_1057,N_17010,N_18603);
nor UO_1058 (O_1058,N_15965,N_18588);
and UO_1059 (O_1059,N_16593,N_18963);
or UO_1060 (O_1060,N_18021,N_19696);
nand UO_1061 (O_1061,N_18636,N_19575);
nand UO_1062 (O_1062,N_18888,N_19905);
or UO_1063 (O_1063,N_19168,N_15448);
nand UO_1064 (O_1064,N_16578,N_18632);
or UO_1065 (O_1065,N_15219,N_16809);
nor UO_1066 (O_1066,N_16892,N_15272);
nor UO_1067 (O_1067,N_19557,N_18517);
nand UO_1068 (O_1068,N_19519,N_17687);
and UO_1069 (O_1069,N_15087,N_16502);
or UO_1070 (O_1070,N_18027,N_19289);
or UO_1071 (O_1071,N_17594,N_18804);
nor UO_1072 (O_1072,N_18246,N_17092);
nand UO_1073 (O_1073,N_17847,N_18692);
xnor UO_1074 (O_1074,N_18201,N_16288);
and UO_1075 (O_1075,N_18962,N_15348);
and UO_1076 (O_1076,N_18741,N_15149);
nand UO_1077 (O_1077,N_18387,N_19200);
and UO_1078 (O_1078,N_15004,N_15036);
nand UO_1079 (O_1079,N_18467,N_15526);
or UO_1080 (O_1080,N_15534,N_18267);
nor UO_1081 (O_1081,N_18578,N_16985);
nand UO_1082 (O_1082,N_18328,N_16698);
xnor UO_1083 (O_1083,N_16380,N_18591);
nor UO_1084 (O_1084,N_16360,N_19425);
or UO_1085 (O_1085,N_17588,N_18486);
or UO_1086 (O_1086,N_18162,N_19357);
or UO_1087 (O_1087,N_16440,N_15883);
or UO_1088 (O_1088,N_15152,N_18573);
or UO_1089 (O_1089,N_18453,N_16194);
nor UO_1090 (O_1090,N_17043,N_15874);
nand UO_1091 (O_1091,N_16655,N_18064);
nand UO_1092 (O_1092,N_16211,N_16438);
nor UO_1093 (O_1093,N_18732,N_19329);
or UO_1094 (O_1094,N_16722,N_17566);
or UO_1095 (O_1095,N_18654,N_19960);
xor UO_1096 (O_1096,N_17866,N_16991);
nand UO_1097 (O_1097,N_18647,N_15547);
or UO_1098 (O_1098,N_19765,N_16308);
xor UO_1099 (O_1099,N_17850,N_17655);
or UO_1100 (O_1100,N_19970,N_15798);
nor UO_1101 (O_1101,N_17977,N_15378);
nand UO_1102 (O_1102,N_15216,N_18671);
or UO_1103 (O_1103,N_18559,N_16560);
and UO_1104 (O_1104,N_17993,N_15340);
and UO_1105 (O_1105,N_18115,N_15663);
or UO_1106 (O_1106,N_18641,N_19473);
xnor UO_1107 (O_1107,N_18135,N_19206);
nor UO_1108 (O_1108,N_16436,N_16799);
nor UO_1109 (O_1109,N_17587,N_16803);
nor UO_1110 (O_1110,N_15562,N_19250);
and UO_1111 (O_1111,N_17712,N_18700);
and UO_1112 (O_1112,N_18116,N_18433);
and UO_1113 (O_1113,N_17519,N_15116);
and UO_1114 (O_1114,N_16293,N_17019);
and UO_1115 (O_1115,N_16817,N_18988);
nand UO_1116 (O_1116,N_19101,N_19664);
or UO_1117 (O_1117,N_18943,N_15551);
or UO_1118 (O_1118,N_18160,N_17011);
and UO_1119 (O_1119,N_19792,N_17364);
nand UO_1120 (O_1120,N_17796,N_19492);
and UO_1121 (O_1121,N_19003,N_19839);
xnor UO_1122 (O_1122,N_17063,N_19447);
or UO_1123 (O_1123,N_16648,N_16096);
or UO_1124 (O_1124,N_18122,N_17482);
nor UO_1125 (O_1125,N_17916,N_15025);
nand UO_1126 (O_1126,N_17205,N_17242);
or UO_1127 (O_1127,N_19867,N_16069);
nand UO_1128 (O_1128,N_19767,N_18718);
and UO_1129 (O_1129,N_16093,N_15966);
and UO_1130 (O_1130,N_16897,N_19940);
nor UO_1131 (O_1131,N_19070,N_15994);
nand UO_1132 (O_1132,N_19826,N_18075);
nor UO_1133 (O_1133,N_17701,N_15484);
nand UO_1134 (O_1134,N_17352,N_19444);
nor UO_1135 (O_1135,N_15540,N_17119);
nand UO_1136 (O_1136,N_19683,N_15752);
nand UO_1137 (O_1137,N_19001,N_17118);
xnor UO_1138 (O_1138,N_18835,N_19411);
nor UO_1139 (O_1139,N_15322,N_16165);
nor UO_1140 (O_1140,N_15890,N_19769);
nor UO_1141 (O_1141,N_19515,N_15688);
nor UO_1142 (O_1142,N_15863,N_15321);
or UO_1143 (O_1143,N_19687,N_16429);
nand UO_1144 (O_1144,N_16806,N_18468);
nand UO_1145 (O_1145,N_19709,N_18376);
or UO_1146 (O_1146,N_17798,N_16409);
nor UO_1147 (O_1147,N_19993,N_18293);
and UO_1148 (O_1148,N_15443,N_16271);
nor UO_1149 (O_1149,N_19079,N_15460);
xor UO_1150 (O_1150,N_19562,N_19370);
nand UO_1151 (O_1151,N_16949,N_19831);
nand UO_1152 (O_1152,N_17257,N_16845);
or UO_1153 (O_1153,N_18185,N_16474);
or UO_1154 (O_1154,N_16581,N_18708);
and UO_1155 (O_1155,N_19660,N_16428);
nor UO_1156 (O_1156,N_16363,N_15630);
xor UO_1157 (O_1157,N_18609,N_18705);
nand UO_1158 (O_1158,N_19073,N_19857);
nor UO_1159 (O_1159,N_17737,N_19843);
nor UO_1160 (O_1160,N_15958,N_15689);
nor UO_1161 (O_1161,N_15703,N_18018);
or UO_1162 (O_1162,N_17934,N_18445);
and UO_1163 (O_1163,N_18528,N_19662);
or UO_1164 (O_1164,N_15871,N_19293);
nor UO_1165 (O_1165,N_18834,N_18935);
nand UO_1166 (O_1166,N_18069,N_16567);
and UO_1167 (O_1167,N_15812,N_15959);
or UO_1168 (O_1168,N_18012,N_18961);
or UO_1169 (O_1169,N_15672,N_19876);
nor UO_1170 (O_1170,N_18543,N_15927);
nor UO_1171 (O_1171,N_18423,N_17197);
nor UO_1172 (O_1172,N_16386,N_17791);
and UO_1173 (O_1173,N_19197,N_19742);
nand UO_1174 (O_1174,N_18873,N_18994);
and UO_1175 (O_1175,N_18047,N_17812);
nor UO_1176 (O_1176,N_19389,N_18282);
nor UO_1177 (O_1177,N_19019,N_16233);
nand UO_1178 (O_1178,N_19328,N_15367);
and UO_1179 (O_1179,N_17580,N_16871);
nor UO_1180 (O_1180,N_19774,N_16907);
nand UO_1181 (O_1181,N_15455,N_16721);
or UO_1182 (O_1182,N_19404,N_17527);
or UO_1183 (O_1183,N_17308,N_16482);
or UO_1184 (O_1184,N_19656,N_16417);
or UO_1185 (O_1185,N_17213,N_16699);
or UO_1186 (O_1186,N_18499,N_16078);
and UO_1187 (O_1187,N_19981,N_18932);
xnor UO_1188 (O_1188,N_19878,N_17899);
and UO_1189 (O_1189,N_18540,N_16982);
nor UO_1190 (O_1190,N_19847,N_18848);
or UO_1191 (O_1191,N_16944,N_19896);
and UO_1192 (O_1192,N_17111,N_19355);
or UO_1193 (O_1193,N_19134,N_19451);
nor UO_1194 (O_1194,N_17450,N_17459);
and UO_1195 (O_1195,N_17216,N_16603);
and UO_1196 (O_1196,N_18545,N_15641);
or UO_1197 (O_1197,N_18090,N_15007);
and UO_1198 (O_1198,N_16814,N_18611);
or UO_1199 (O_1199,N_16776,N_18094);
nor UO_1200 (O_1200,N_16774,N_16905);
and UO_1201 (O_1201,N_15817,N_16913);
nor UO_1202 (O_1202,N_15776,N_18773);
or UO_1203 (O_1203,N_18119,N_15823);
and UO_1204 (O_1204,N_15099,N_18312);
or UO_1205 (O_1205,N_15344,N_16821);
nor UO_1206 (O_1206,N_17175,N_19430);
nand UO_1207 (O_1207,N_17660,N_16864);
and UO_1208 (O_1208,N_17696,N_18547);
or UO_1209 (O_1209,N_16714,N_18455);
or UO_1210 (O_1210,N_19422,N_15740);
xor UO_1211 (O_1211,N_17031,N_15991);
nor UO_1212 (O_1212,N_15898,N_17609);
and UO_1213 (O_1213,N_16220,N_17859);
xor UO_1214 (O_1214,N_17736,N_19103);
and UO_1215 (O_1215,N_19302,N_19384);
and UO_1216 (O_1216,N_17787,N_19130);
or UO_1217 (O_1217,N_15088,N_16759);
nand UO_1218 (O_1218,N_18892,N_15017);
and UO_1219 (O_1219,N_18454,N_19827);
and UO_1220 (O_1220,N_18769,N_17173);
nand UO_1221 (O_1221,N_16099,N_17401);
and UO_1222 (O_1222,N_18620,N_17483);
nor UO_1223 (O_1223,N_16847,N_16670);
or UO_1224 (O_1224,N_17672,N_15650);
xnor UO_1225 (O_1225,N_18377,N_15167);
or UO_1226 (O_1226,N_18200,N_17910);
nor UO_1227 (O_1227,N_17485,N_17417);
nand UO_1228 (O_1228,N_17624,N_18007);
nand UO_1229 (O_1229,N_16260,N_17479);
nor UO_1230 (O_1230,N_18296,N_18899);
or UO_1231 (O_1231,N_15126,N_17248);
nor UO_1232 (O_1232,N_16102,N_16178);
nor UO_1233 (O_1233,N_18569,N_17312);
nor UO_1234 (O_1234,N_15730,N_15306);
and UO_1235 (O_1235,N_19962,N_15302);
or UO_1236 (O_1236,N_17880,N_15010);
and UO_1237 (O_1237,N_16815,N_15386);
nand UO_1238 (O_1238,N_19335,N_18792);
and UO_1239 (O_1239,N_19274,N_15037);
xnor UO_1240 (O_1240,N_19533,N_17414);
nor UO_1241 (O_1241,N_15489,N_19921);
and UO_1242 (O_1242,N_16071,N_19880);
or UO_1243 (O_1243,N_18530,N_15807);
nor UO_1244 (O_1244,N_17968,N_17462);
nor UO_1245 (O_1245,N_17909,N_17471);
nand UO_1246 (O_1246,N_15039,N_15470);
nand UO_1247 (O_1247,N_15154,N_18053);
nand UO_1248 (O_1248,N_16996,N_15353);
xnor UO_1249 (O_1249,N_16252,N_15407);
and UO_1250 (O_1250,N_16682,N_15483);
and UO_1251 (O_1251,N_19056,N_18788);
and UO_1252 (O_1252,N_16939,N_19027);
and UO_1253 (O_1253,N_16533,N_16573);
nand UO_1254 (O_1254,N_19386,N_15365);
or UO_1255 (O_1255,N_17849,N_19225);
or UO_1256 (O_1256,N_15328,N_16849);
nor UO_1257 (O_1257,N_18655,N_16886);
nand UO_1258 (O_1258,N_19439,N_15094);
and UO_1259 (O_1259,N_18631,N_15825);
nand UO_1260 (O_1260,N_15913,N_15746);
xnor UO_1261 (O_1261,N_15990,N_16036);
nor UO_1262 (O_1262,N_16393,N_17988);
nor UO_1263 (O_1263,N_18900,N_19730);
nor UO_1264 (O_1264,N_17955,N_17869);
or UO_1265 (O_1265,N_16883,N_19710);
nand UO_1266 (O_1266,N_15678,N_19754);
nor UO_1267 (O_1267,N_19278,N_16793);
xnor UO_1268 (O_1268,N_15346,N_17339);
or UO_1269 (O_1269,N_16250,N_16608);
nor UO_1270 (O_1270,N_18155,N_15931);
or UO_1271 (O_1271,N_17839,N_16606);
xor UO_1272 (O_1272,N_16710,N_16689);
or UO_1273 (O_1273,N_18157,N_16423);
nand UO_1274 (O_1274,N_18138,N_17167);
and UO_1275 (O_1275,N_19607,N_18356);
nand UO_1276 (O_1276,N_16790,N_15478);
nand UO_1277 (O_1277,N_16750,N_18443);
nor UO_1278 (O_1278,N_19218,N_19275);
nand UO_1279 (O_1279,N_17211,N_17169);
and UO_1280 (O_1280,N_15923,N_15626);
nand UO_1281 (O_1281,N_16065,N_18332);
or UO_1282 (O_1282,N_16496,N_19546);
and UO_1283 (O_1283,N_16989,N_15123);
nand UO_1284 (O_1284,N_18601,N_18124);
and UO_1285 (O_1285,N_17596,N_19255);
nand UO_1286 (O_1286,N_17334,N_16079);
and UO_1287 (O_1287,N_18250,N_19334);
and UO_1288 (O_1288,N_18049,N_18495);
or UO_1289 (O_1289,N_18226,N_18838);
and UO_1290 (O_1290,N_16383,N_16018);
nand UO_1291 (O_1291,N_15814,N_19252);
nand UO_1292 (O_1292,N_18082,N_17246);
and UO_1293 (O_1293,N_15847,N_18673);
nor UO_1294 (O_1294,N_15187,N_16120);
nand UO_1295 (O_1295,N_19518,N_18890);
nand UO_1296 (O_1296,N_19860,N_16677);
or UO_1297 (O_1297,N_18917,N_16683);
nand UO_1298 (O_1298,N_16508,N_15334);
nand UO_1299 (O_1299,N_17838,N_16094);
xnor UO_1300 (O_1300,N_19698,N_18058);
nand UO_1301 (O_1301,N_17238,N_17454);
nor UO_1302 (O_1302,N_19984,N_15127);
nand UO_1303 (O_1303,N_15699,N_18726);
and UO_1304 (O_1304,N_19331,N_15467);
nor UO_1305 (O_1305,N_17894,N_15727);
or UO_1306 (O_1306,N_15851,N_15855);
and UO_1307 (O_1307,N_17064,N_15260);
nor UO_1308 (O_1308,N_17667,N_15897);
or UO_1309 (O_1309,N_16649,N_15751);
nand UO_1310 (O_1310,N_19910,N_16231);
xor UO_1311 (O_1311,N_18415,N_16114);
nor UO_1312 (O_1312,N_16629,N_19420);
and UO_1313 (O_1313,N_16861,N_16592);
nand UO_1314 (O_1314,N_16733,N_15583);
nor UO_1315 (O_1315,N_17608,N_19394);
nor UO_1316 (O_1316,N_16206,N_17813);
or UO_1317 (O_1317,N_19285,N_19496);
xor UO_1318 (O_1318,N_19237,N_16811);
or UO_1319 (O_1319,N_15600,N_19931);
xnor UO_1320 (O_1320,N_16820,N_19012);
or UO_1321 (O_1321,N_19044,N_17746);
nand UO_1322 (O_1322,N_18035,N_18678);
nor UO_1323 (O_1323,N_15416,N_17943);
nor UO_1324 (O_1324,N_18022,N_16620);
xor UO_1325 (O_1325,N_19994,N_18712);
nor UO_1326 (O_1326,N_17645,N_18983);
or UO_1327 (O_1327,N_15964,N_17223);
or UO_1328 (O_1328,N_16356,N_16580);
and UO_1329 (O_1329,N_18677,N_19516);
or UO_1330 (O_1330,N_19261,N_18521);
or UO_1331 (O_1331,N_15584,N_18031);
or UO_1332 (O_1332,N_17315,N_18972);
or UO_1333 (O_1333,N_18616,N_16950);
nor UO_1334 (O_1334,N_16118,N_17855);
nand UO_1335 (O_1335,N_19093,N_19547);
nor UO_1336 (O_1336,N_16819,N_18597);
and UO_1337 (O_1337,N_15792,N_18251);
nand UO_1338 (O_1338,N_15877,N_18758);
nor UO_1339 (O_1339,N_17665,N_15793);
or UO_1340 (O_1340,N_17524,N_15019);
and UO_1341 (O_1341,N_15213,N_15571);
nor UO_1342 (O_1342,N_15298,N_16943);
nor UO_1343 (O_1343,N_16049,N_16201);
nand UO_1344 (O_1344,N_15758,N_19489);
nand UO_1345 (O_1345,N_19668,N_19944);
nand UO_1346 (O_1346,N_19123,N_19950);
or UO_1347 (O_1347,N_18565,N_18633);
and UO_1348 (O_1348,N_17619,N_16207);
and UO_1349 (O_1349,N_16577,N_16243);
nor UO_1350 (O_1350,N_15490,N_18081);
and UO_1351 (O_1351,N_17722,N_17259);
or UO_1352 (O_1352,N_19576,N_16564);
nor UO_1353 (O_1353,N_19126,N_15183);
or UO_1354 (O_1354,N_18440,N_17992);
and UO_1355 (O_1355,N_19041,N_18843);
nor UO_1356 (O_1356,N_19653,N_18659);
nor UO_1357 (O_1357,N_18010,N_18939);
and UO_1358 (O_1358,N_18879,N_15403);
nand UO_1359 (O_1359,N_19773,N_17769);
and UO_1360 (O_1360,N_16095,N_18921);
nor UO_1361 (O_1361,N_16195,N_16640);
and UO_1362 (O_1362,N_16595,N_19990);
nand UO_1363 (O_1363,N_15643,N_18067);
nor UO_1364 (O_1364,N_16305,N_17049);
nor UO_1365 (O_1365,N_16022,N_16458);
xnor UO_1366 (O_1366,N_17112,N_19978);
or UO_1367 (O_1367,N_15119,N_16756);
and UO_1368 (O_1368,N_15697,N_15715);
nand UO_1369 (O_1369,N_18488,N_19423);
or UO_1370 (O_1370,N_19209,N_16117);
nor UO_1371 (O_1371,N_17143,N_17145);
nand UO_1372 (O_1372,N_16734,N_18660);
and UO_1373 (O_1373,N_15852,N_19936);
and UO_1374 (O_1374,N_19695,N_16374);
nor UO_1375 (O_1375,N_15337,N_15502);
or UO_1376 (O_1376,N_18245,N_15210);
nor UO_1377 (O_1377,N_16446,N_16139);
and UO_1378 (O_1378,N_16416,N_19373);
and UO_1379 (O_1379,N_15191,N_18319);
nor UO_1380 (O_1380,N_16590,N_18825);
or UO_1381 (O_1381,N_17353,N_17466);
nand UO_1382 (O_1382,N_18313,N_16138);
and UO_1383 (O_1383,N_19446,N_18725);
xnor UO_1384 (O_1384,N_18165,N_18789);
xor UO_1385 (O_1385,N_15105,N_15777);
nand UO_1386 (O_1386,N_18901,N_17816);
nand UO_1387 (O_1387,N_17831,N_18531);
nor UO_1388 (O_1388,N_18425,N_15464);
nor UO_1389 (O_1389,N_15479,N_16479);
and UO_1390 (O_1390,N_15268,N_15648);
nor UO_1391 (O_1391,N_17061,N_17311);
xor UO_1392 (O_1392,N_16671,N_16286);
nor UO_1393 (O_1393,N_16833,N_15950);
xnor UO_1394 (O_1394,N_18984,N_19832);
nor UO_1395 (O_1395,N_16717,N_17886);
or UO_1396 (O_1396,N_16349,N_17100);
and UO_1397 (O_1397,N_19574,N_16481);
nand UO_1398 (O_1398,N_16312,N_15880);
or UO_1399 (O_1399,N_17929,N_15022);
nand UO_1400 (O_1400,N_16323,N_18759);
xor UO_1401 (O_1401,N_17237,N_19095);
and UO_1402 (O_1402,N_15003,N_15248);
or UO_1403 (O_1403,N_15819,N_18006);
nor UO_1404 (O_1404,N_15076,N_17178);
and UO_1405 (O_1405,N_18096,N_17922);
or UO_1406 (O_1406,N_19269,N_16563);
or UO_1407 (O_1407,N_19229,N_15034);
or UO_1408 (O_1408,N_17919,N_17055);
nand UO_1409 (O_1409,N_17844,N_19610);
xor UO_1410 (O_1410,N_18218,N_17464);
and UO_1411 (O_1411,N_19704,N_19813);
nand UO_1412 (O_1412,N_19545,N_19976);
and UO_1413 (O_1413,N_16313,N_16925);
or UO_1414 (O_1414,N_16651,N_18730);
and UO_1415 (O_1415,N_19436,N_16657);
nand UO_1416 (O_1416,N_15986,N_19498);
nor UO_1417 (O_1417,N_16203,N_19348);
nand UO_1418 (O_1418,N_18895,N_15962);
and UO_1419 (O_1419,N_18017,N_16623);
nand UO_1420 (O_1420,N_17188,N_17965);
nor UO_1421 (O_1421,N_16705,N_15633);
xor UO_1422 (O_1422,N_18970,N_18214);
or UO_1423 (O_1423,N_18688,N_17058);
and UO_1424 (O_1424,N_16394,N_19432);
nor UO_1425 (O_1425,N_17378,N_19534);
or UO_1426 (O_1426,N_16841,N_18072);
nor UO_1427 (O_1427,N_18716,N_19810);
or UO_1428 (O_1428,N_18148,N_17967);
nand UO_1429 (O_1429,N_17926,N_19858);
or UO_1430 (O_1430,N_16164,N_19416);
nand UO_1431 (O_1431,N_19763,N_16800);
nor UO_1432 (O_1432,N_16272,N_19458);
xnor UO_1433 (O_1433,N_17014,N_17896);
xnor UO_1434 (O_1434,N_19529,N_19724);
nand UO_1435 (O_1435,N_17832,N_18041);
nor UO_1436 (O_1436,N_18057,N_17183);
or UO_1437 (O_1437,N_19155,N_17277);
nand UO_1438 (O_1438,N_18763,N_19354);
nor UO_1439 (O_1439,N_17048,N_17236);
and UO_1440 (O_1440,N_16039,N_18206);
nand UO_1441 (O_1441,N_16910,N_15553);
xor UO_1442 (O_1442,N_18000,N_15423);
xor UO_1443 (O_1443,N_15556,N_16126);
nor UO_1444 (O_1444,N_18070,N_17095);
xor UO_1445 (O_1445,N_18576,N_16382);
and UO_1446 (O_1446,N_17906,N_16024);
xor UO_1447 (O_1447,N_16527,N_15977);
nand UO_1448 (O_1448,N_18083,N_15827);
and UO_1449 (O_1449,N_15886,N_15546);
nor UO_1450 (O_1450,N_15563,N_18136);
nand UO_1451 (O_1451,N_18403,N_18048);
nor UO_1452 (O_1452,N_18001,N_18434);
and UO_1453 (O_1453,N_19288,N_17881);
and UO_1454 (O_1454,N_16694,N_17425);
and UO_1455 (O_1455,N_15462,N_19932);
or UO_1456 (O_1456,N_18869,N_18228);
nor UO_1457 (O_1457,N_19643,N_15066);
and UO_1458 (O_1458,N_17695,N_18777);
or UO_1459 (O_1459,N_18424,N_19554);
nand UO_1460 (O_1460,N_18220,N_19916);
and UO_1461 (O_1461,N_15946,N_19356);
or UO_1462 (O_1462,N_15907,N_15655);
or UO_1463 (O_1463,N_18906,N_18284);
or UO_1464 (O_1464,N_17382,N_18406);
or UO_1465 (O_1465,N_16249,N_19459);
nor UO_1466 (O_1466,N_19532,N_16133);
and UO_1467 (O_1467,N_15405,N_15921);
and UO_1468 (O_1468,N_19783,N_19837);
nand UO_1469 (O_1469,N_18783,N_18882);
and UO_1470 (O_1470,N_17136,N_18364);
nand UO_1471 (O_1471,N_18508,N_18523);
nand UO_1472 (O_1472,N_17822,N_19633);
nand UO_1473 (O_1473,N_16783,N_15021);
or UO_1474 (O_1474,N_19945,N_18973);
nand UO_1475 (O_1475,N_19947,N_18981);
nand UO_1476 (O_1476,N_19243,N_16391);
or UO_1477 (O_1477,N_18649,N_17455);
and UO_1478 (O_1478,N_17091,N_16147);
nor UO_1479 (O_1479,N_19199,N_16997);
nand UO_1480 (O_1480,N_15469,N_18561);
nand UO_1481 (O_1481,N_15980,N_18033);
or UO_1482 (O_1482,N_18750,N_16487);
nand UO_1483 (O_1483,N_19951,N_16119);
nor UO_1484 (O_1484,N_17396,N_16144);
nor UO_1485 (O_1485,N_16345,N_19503);
nand UO_1486 (O_1486,N_17597,N_17642);
nor UO_1487 (O_1487,N_19180,N_18662);
and UO_1488 (O_1488,N_15928,N_17093);
nand UO_1489 (O_1489,N_18026,N_18390);
and UO_1490 (O_1490,N_15784,N_17330);
xnor UO_1491 (O_1491,N_15463,N_17422);
xor UO_1492 (O_1492,N_19686,N_15214);
nor UO_1493 (O_1493,N_17682,N_16208);
nor UO_1494 (O_1494,N_17647,N_19226);
nor UO_1495 (O_1495,N_16322,N_16621);
or UO_1496 (O_1496,N_16007,N_16398);
nor UO_1497 (O_1497,N_16731,N_17204);
and UO_1498 (O_1498,N_19172,N_18395);
and UO_1499 (O_1499,N_16804,N_16077);
and UO_1500 (O_1500,N_15588,N_16530);
and UO_1501 (O_1501,N_15654,N_15596);
and UO_1502 (O_1502,N_18745,N_15238);
and UO_1503 (O_1503,N_16760,N_17814);
xor UO_1504 (O_1504,N_15775,N_16702);
xnor UO_1505 (O_1505,N_18809,N_18235);
nand UO_1506 (O_1506,N_15682,N_19756);
and UO_1507 (O_1507,N_17790,N_16882);
nor UO_1508 (O_1508,N_17288,N_19074);
and UO_1509 (O_1509,N_17374,N_15060);
or UO_1510 (O_1510,N_19830,N_18190);
or UO_1511 (O_1511,N_19427,N_17229);
xnor UO_1512 (O_1512,N_15624,N_16205);
nand UO_1513 (O_1513,N_15041,N_17708);
or UO_1514 (O_1514,N_17957,N_19983);
nor UO_1515 (O_1515,N_17487,N_16539);
nor UO_1516 (O_1516,N_16486,N_17088);
nand UO_1517 (O_1517,N_19744,N_15465);
nand UO_1518 (O_1518,N_17901,N_16043);
nor UO_1519 (O_1519,N_15925,N_17271);
nand UO_1520 (O_1520,N_17155,N_15503);
and UO_1521 (O_1521,N_18417,N_16172);
or UO_1522 (O_1522,N_16295,N_17405);
and UO_1523 (O_1523,N_17557,N_15275);
and UO_1524 (O_1524,N_16184,N_19986);
xnor UO_1525 (O_1525,N_19142,N_18697);
nor UO_1526 (O_1526,N_19846,N_17732);
or UO_1527 (O_1527,N_17022,N_15559);
or UO_1528 (O_1528,N_15570,N_16239);
xnor UO_1529 (O_1529,N_15288,N_18329);
nand UO_1530 (O_1530,N_16618,N_19267);
and UO_1531 (O_1531,N_15058,N_16402);
nor UO_1532 (O_1532,N_19535,N_19195);
and UO_1533 (O_1533,N_17541,N_16335);
nor UO_1534 (O_1534,N_19374,N_16324);
nand UO_1535 (O_1535,N_16227,N_16089);
and UO_1536 (O_1536,N_19873,N_15859);
and UO_1537 (O_1537,N_16357,N_17157);
nor UO_1538 (O_1538,N_19996,N_16770);
nor UO_1539 (O_1539,N_16015,N_16938);
and UO_1540 (O_1540,N_18729,N_15188);
nor UO_1541 (O_1541,N_17878,N_19257);
xor UO_1542 (O_1542,N_15000,N_15224);
and UO_1543 (O_1543,N_15675,N_16874);
nor UO_1544 (O_1544,N_18175,N_15316);
and UO_1545 (O_1545,N_16418,N_17800);
xnor UO_1546 (O_1546,N_17714,N_17593);
nor UO_1547 (O_1547,N_16105,N_15935);
nand UO_1548 (O_1548,N_19911,N_18414);
nor UO_1549 (O_1549,N_16129,N_16341);
nor UO_1550 (O_1550,N_15255,N_15333);
xor UO_1551 (O_1551,N_18604,N_17153);
nor UO_1552 (O_1552,N_19035,N_17782);
and UO_1553 (O_1553,N_15757,N_19966);
or UO_1554 (O_1554,N_15311,N_19127);
nor UO_1555 (O_1555,N_17161,N_16955);
nor UO_1556 (O_1556,N_17928,N_17927);
nor UO_1557 (O_1557,N_16278,N_18066);
nor UO_1558 (O_1558,N_19176,N_17601);
and UO_1559 (O_1559,N_15449,N_19300);
or UO_1560 (O_1560,N_18919,N_18203);
nor UO_1561 (O_1561,N_15324,N_18024);
or UO_1562 (O_1562,N_15366,N_19644);
and UO_1563 (O_1563,N_18793,N_16074);
or UO_1564 (O_1564,N_15284,N_15239);
nor UO_1565 (O_1565,N_15035,N_17065);
nand UO_1566 (O_1566,N_16737,N_16645);
and UO_1567 (O_1567,N_18638,N_17047);
and UO_1568 (O_1568,N_17598,N_19114);
or UO_1569 (O_1569,N_17617,N_15067);
and UO_1570 (O_1570,N_17431,N_18345);
and UO_1571 (O_1571,N_15444,N_19472);
or UO_1572 (O_1572,N_18013,N_19589);
xnor UO_1573 (O_1573,N_15698,N_16085);
nand UO_1574 (O_1574,N_18259,N_16376);
or UO_1575 (O_1575,N_15528,N_15173);
xor UO_1576 (O_1576,N_16569,N_19476);
and UO_1577 (O_1577,N_15701,N_17434);
nand UO_1578 (O_1578,N_15057,N_18803);
and UO_1579 (O_1579,N_16154,N_19648);
or UO_1580 (O_1580,N_18857,N_16317);
nand UO_1581 (O_1581,N_15885,N_17907);
or UO_1582 (O_1582,N_15914,N_18702);
nor UO_1583 (O_1583,N_18118,N_18930);
xnor UO_1584 (O_1584,N_18946,N_15143);
nand UO_1585 (O_1585,N_17600,N_17942);
and UO_1586 (O_1586,N_19597,N_18822);
or UO_1587 (O_1587,N_15822,N_17763);
or UO_1588 (O_1588,N_17398,N_18431);
xnor UO_1589 (O_1589,N_17354,N_16862);
or UO_1590 (O_1590,N_16230,N_16707);
and UO_1591 (O_1591,N_19613,N_18477);
nor UO_1592 (O_1592,N_19026,N_19084);
nor UO_1593 (O_1593,N_17276,N_15645);
and UO_1594 (O_1594,N_17437,N_16909);
nor UO_1595 (O_1595,N_19375,N_17122);
nand UO_1596 (O_1596,N_15180,N_19015);
or UO_1597 (O_1597,N_16875,N_15234);
nor UO_1598 (O_1598,N_16986,N_19637);
nand UO_1599 (O_1599,N_16524,N_16143);
and UO_1600 (O_1600,N_15230,N_17559);
and UO_1601 (O_1601,N_15937,N_19750);
and UO_1602 (O_1602,N_17705,N_19010);
or UO_1603 (O_1603,N_15244,N_16097);
nor UO_1604 (O_1604,N_16012,N_17359);
or UO_1605 (O_1605,N_16828,N_19481);
or UO_1606 (O_1606,N_17025,N_16460);
nand UO_1607 (O_1607,N_18837,N_18675);
and UO_1608 (O_1608,N_18375,N_18435);
nand UO_1609 (O_1609,N_16742,N_15200);
nor UO_1610 (O_1610,N_17116,N_17944);
nor UO_1611 (O_1611,N_16898,N_19500);
nand UO_1612 (O_1612,N_18695,N_17544);
and UO_1613 (O_1613,N_15056,N_15894);
nand UO_1614 (O_1614,N_19241,N_17890);
nor UO_1615 (O_1615,N_15625,N_18279);
nand UO_1616 (O_1616,N_16412,N_19479);
xnor UO_1617 (O_1617,N_15226,N_17729);
and UO_1618 (O_1618,N_19202,N_16002);
or UO_1619 (O_1619,N_17973,N_16805);
or UO_1620 (O_1620,N_18987,N_18152);
or UO_1621 (O_1621,N_15541,N_15857);
or UO_1622 (O_1622,N_15398,N_19196);
nand UO_1623 (O_1623,N_17663,N_16911);
nor UO_1624 (O_1624,N_18571,N_15185);
xor UO_1625 (O_1625,N_19615,N_17780);
or UO_1626 (O_1626,N_17451,N_18274);
xnor UO_1627 (O_1627,N_15247,N_17286);
and UO_1628 (O_1628,N_17785,N_16965);
nand UO_1629 (O_1629,N_17793,N_17453);
nor UO_1630 (O_1630,N_18915,N_18727);
or UO_1631 (O_1631,N_16628,N_19419);
and UO_1632 (O_1632,N_17194,N_16503);
or UO_1633 (O_1633,N_18233,N_19380);
nand UO_1634 (O_1634,N_15545,N_19098);
and UO_1635 (O_1635,N_18270,N_18867);
or UO_1636 (O_1636,N_19276,N_18766);
or UO_1637 (O_1637,N_17670,N_15906);
and UO_1638 (O_1638,N_18819,N_19456);
nor UO_1639 (O_1639,N_16958,N_17644);
nor UO_1640 (O_1640,N_15679,N_18801);
nand UO_1641 (O_1641,N_15829,N_19736);
nand UO_1642 (O_1642,N_18776,N_18851);
or UO_1643 (O_1643,N_17337,N_16868);
or UO_1644 (O_1644,N_19167,N_18432);
nand UO_1645 (O_1645,N_16047,N_18408);
nor UO_1646 (O_1646,N_16037,N_15421);
or UO_1647 (O_1647,N_19570,N_15345);
nor UO_1648 (O_1648,N_18504,N_18457);
and UO_1649 (O_1649,N_19542,N_19685);
or UO_1650 (O_1650,N_15232,N_19699);
and UO_1651 (O_1651,N_15988,N_18731);
or UO_1652 (O_1652,N_15450,N_19563);
and UO_1653 (O_1653,N_19762,N_19729);
nand UO_1654 (O_1654,N_19799,N_18444);
or UO_1655 (O_1655,N_17096,N_18640);
nand UO_1656 (O_1656,N_16990,N_18509);
nor UO_1657 (O_1657,N_17828,N_17214);
or UO_1658 (O_1658,N_18826,N_17000);
or UO_1659 (O_1659,N_15078,N_17199);
nand UO_1660 (O_1660,N_18223,N_15429);
nand UO_1661 (O_1661,N_17863,N_18427);
xor UO_1662 (O_1662,N_15218,N_18416);
nor UO_1663 (O_1663,N_19771,N_16983);
nand UO_1664 (O_1664,N_17516,N_15686);
nor UO_1665 (O_1665,N_18359,N_18280);
nor UO_1666 (O_1666,N_16528,N_19438);
nor UO_1667 (O_1667,N_19650,N_18653);
and UO_1668 (O_1668,N_19484,N_17940);
or UO_1669 (O_1669,N_15790,N_16807);
or UO_1670 (O_1670,N_15476,N_19021);
and UO_1671 (O_1671,N_17309,N_19296);
nor UO_1672 (O_1672,N_18036,N_15118);
xnor UO_1673 (O_1673,N_17912,N_17495);
nor UO_1674 (O_1674,N_19775,N_15024);
or UO_1675 (O_1675,N_19720,N_15445);
nand UO_1676 (O_1676,N_18596,N_15015);
or UO_1677 (O_1677,N_19170,N_19822);
or UO_1678 (O_1678,N_16642,N_17523);
nand UO_1679 (O_1679,N_15211,N_16979);
or UO_1680 (O_1680,N_16369,N_17612);
and UO_1681 (O_1681,N_16101,N_18060);
or UO_1682 (O_1682,N_16916,N_15587);
and UO_1683 (O_1683,N_18897,N_18028);
nand UO_1684 (O_1684,N_17506,N_15397);
nand UO_1685 (O_1685,N_17570,N_19254);
and UO_1686 (O_1686,N_18894,N_15160);
or UO_1687 (O_1687,N_15392,N_18479);
or UO_1688 (O_1688,N_19787,N_18232);
nand UO_1689 (O_1689,N_18666,N_15674);
or UO_1690 (O_1690,N_17759,N_17833);
xor UO_1691 (O_1691,N_15800,N_19675);
or UO_1692 (O_1692,N_16232,N_19258);
nand UO_1693 (O_1693,N_18229,N_19174);
or UO_1694 (O_1694,N_15606,N_19339);
xor UO_1695 (O_1695,N_16413,N_18016);
nand UO_1696 (O_1696,N_18550,N_18847);
and UO_1697 (O_1697,N_19523,N_16202);
nor UO_1698 (O_1698,N_18337,N_18485);
or UO_1699 (O_1699,N_19193,N_15415);
nand UO_1700 (O_1700,N_17578,N_17817);
xnor UO_1701 (O_1701,N_15354,N_18273);
nor UO_1702 (O_1702,N_19002,N_17123);
and UO_1703 (O_1703,N_19330,N_15670);
and UO_1704 (O_1704,N_15355,N_17626);
nand UO_1705 (O_1705,N_15786,N_15304);
nand UO_1706 (O_1706,N_19110,N_19188);
nor UO_1707 (O_1707,N_18714,N_15237);
nor UO_1708 (O_1708,N_16122,N_16576);
nor UO_1709 (O_1709,N_17184,N_19992);
nor UO_1710 (O_1710,N_19526,N_15586);
nand UO_1711 (O_1711,N_16370,N_16008);
nand UO_1712 (O_1712,N_16686,N_17789);
nand UO_1713 (O_1713,N_18117,N_18269);
nor UO_1714 (O_1714,N_16384,N_15868);
xor UO_1715 (O_1715,N_16209,N_18311);
nor UO_1716 (O_1716,N_16884,N_16457);
nor UO_1717 (O_1717,N_17692,N_15764);
and UO_1718 (O_1718,N_15704,N_18880);
or UO_1719 (O_1719,N_16918,N_16890);
or UO_1720 (O_1720,N_17090,N_18325);
or UO_1721 (O_1721,N_17530,N_16929);
and UO_1722 (O_1722,N_17394,N_16465);
or UO_1723 (O_1723,N_16767,N_18980);
and UO_1724 (O_1724,N_18197,N_16609);
and UO_1725 (O_1725,N_18808,N_17628);
or UO_1726 (O_1726,N_18532,N_18307);
or UO_1727 (O_1727,N_19514,N_18634);
nand UO_1728 (O_1728,N_18051,N_18133);
and UO_1729 (O_1729,N_17269,N_16351);
or UO_1730 (O_1730,N_18446,N_17810);
or UO_1731 (O_1731,N_17845,N_18451);
nand UO_1732 (O_1732,N_17358,N_16575);
or UO_1733 (O_1733,N_18055,N_17013);
nand UO_1734 (O_1734,N_15069,N_16267);
or UO_1735 (O_1735,N_19040,N_17860);
and UO_1736 (O_1736,N_17220,N_15810);
or UO_1737 (O_1737,N_16264,N_15326);
xor UO_1738 (O_1738,N_15517,N_15662);
and UO_1739 (O_1739,N_17795,N_18549);
and UO_1740 (O_1740,N_19223,N_19369);
or UO_1741 (O_1741,N_19051,N_17258);
and UO_1742 (O_1742,N_16342,N_18555);
or UO_1743 (O_1743,N_15565,N_18584);
and UO_1744 (O_1744,N_17885,N_15147);
xnor UO_1745 (O_1745,N_16747,N_18369);
nand UO_1746 (O_1746,N_15653,N_15724);
nor UO_1747 (O_1747,N_15374,N_15512);
and UO_1748 (O_1748,N_19203,N_15331);
xor UO_1749 (O_1749,N_19877,N_16406);
and UO_1750 (O_1750,N_16421,N_18719);
nand UO_1751 (O_1751,N_19764,N_18199);
or UO_1752 (O_1752,N_15992,N_16597);
or UO_1753 (O_1753,N_16029,N_15108);
nand UO_1754 (O_1754,N_19360,N_18577);
and UO_1755 (O_1755,N_18491,N_16263);
and UO_1756 (O_1756,N_18941,N_16781);
and UO_1757 (O_1757,N_15257,N_15431);
nand UO_1758 (O_1758,N_16255,N_19346);
or UO_1759 (O_1759,N_19713,N_15743);
and UO_1760 (O_1760,N_17151,N_19216);
or UO_1761 (O_1761,N_17935,N_19980);
nand UO_1762 (O_1762,N_16330,N_19326);
nand UO_1763 (O_1763,N_19204,N_15009);
nor UO_1764 (O_1764,N_19182,N_17936);
and UO_1765 (O_1765,N_19580,N_18734);
nand UO_1766 (O_1766,N_18661,N_19400);
or UO_1767 (O_1767,N_17235,N_19694);
nand UO_1768 (O_1768,N_16331,N_19376);
and UO_1769 (O_1769,N_19798,N_16782);
and UO_1770 (O_1770,N_17801,N_15968);
or UO_1771 (O_1771,N_17270,N_19201);
nor UO_1772 (O_1772,N_19920,N_19833);
nor UO_1773 (O_1773,N_15362,N_18736);
nor UO_1774 (O_1774,N_18389,N_17335);
nand UO_1775 (O_1775,N_16283,N_18128);
nor UO_1776 (O_1776,N_18227,N_15376);
or UO_1777 (O_1777,N_17539,N_19024);
nand UO_1778 (O_1778,N_18579,N_18645);
nor UO_1779 (O_1779,N_16470,N_17357);
nand UO_1780 (O_1780,N_17775,N_19409);
nor UO_1781 (O_1781,N_15834,N_15264);
and UO_1782 (O_1782,N_16942,N_16970);
or UO_1783 (O_1783,N_15939,N_17945);
nand UO_1784 (O_1784,N_17222,N_17260);
or UO_1785 (O_1785,N_16176,N_15086);
or UO_1786 (O_1786,N_16162,N_19177);
nor UO_1787 (O_1787,N_17320,N_17658);
xnor UO_1788 (O_1788,N_17774,N_16287);
nand UO_1789 (O_1789,N_19645,N_15250);
nor UO_1790 (O_1790,N_16130,N_15282);
or UO_1791 (O_1791,N_16785,N_15178);
nand UO_1792 (O_1792,N_18084,N_15943);
and UO_1793 (O_1793,N_19270,N_17778);
and UO_1794 (O_1794,N_19778,N_16668);
xor UO_1795 (O_1795,N_19157,N_18290);
xor UO_1796 (O_1796,N_16224,N_17073);
nor UO_1797 (O_1797,N_15475,N_18635);
or UO_1798 (O_1798,N_18912,N_15051);
and UO_1799 (O_1799,N_18219,N_18830);
nor UO_1800 (O_1800,N_18771,N_19512);
or UO_1801 (O_1801,N_19029,N_15833);
nand UO_1802 (O_1802,N_16083,N_15136);
nand UO_1803 (O_1803,N_19914,N_15804);
nor UO_1804 (O_1804,N_18927,N_18494);
or UO_1805 (O_1805,N_15124,N_15642);
and UO_1806 (O_1806,N_19591,N_16353);
nand UO_1807 (O_1807,N_19624,N_17338);
and UO_1808 (O_1808,N_15389,N_19392);
nor UO_1809 (O_1809,N_15349,N_17423);
nand UO_1810 (O_1810,N_19630,N_19011);
nor UO_1811 (O_1811,N_17162,N_19907);
and UO_1812 (O_1812,N_18951,N_17568);
and UO_1813 (O_1813,N_17499,N_17623);
and UO_1814 (O_1814,N_17632,N_16475);
or UO_1815 (O_1815,N_16104,N_19701);
xnor UO_1816 (O_1816,N_15552,N_18799);
xnor UO_1817 (O_1817,N_17618,N_19793);
nor UO_1818 (O_1818,N_18950,N_17154);
or UO_1819 (O_1819,N_17902,N_17904);
and UO_1820 (O_1820,N_19604,N_19148);
nor UO_1821 (O_1821,N_19963,N_16477);
or UO_1822 (O_1822,N_18975,N_17709);
xnor UO_1823 (O_1823,N_17932,N_18958);
or UO_1824 (O_1824,N_18101,N_16931);
nor UO_1825 (O_1825,N_17307,N_17108);
and UO_1826 (O_1826,N_17543,N_16050);
nor UO_1827 (O_1827,N_15865,N_15038);
and UO_1828 (O_1828,N_17275,N_17754);
nand UO_1829 (O_1829,N_18681,N_15084);
nor UO_1830 (O_1830,N_16957,N_17420);
or UO_1831 (O_1831,N_16361,N_18833);
xor UO_1832 (O_1832,N_18210,N_16146);
nor UO_1833 (O_1833,N_15665,N_17325);
or UO_1834 (O_1834,N_18614,N_19291);
nand UO_1835 (O_1835,N_19311,N_15170);
nand UO_1836 (O_1836,N_16934,N_17865);
or UO_1837 (O_1837,N_16551,N_15543);
or UO_1838 (O_1838,N_18437,N_16070);
nor UO_1839 (O_1839,N_17864,N_17192);
and UO_1840 (O_1840,N_16895,N_19076);
or UO_1841 (O_1841,N_15861,N_17699);
nor UO_1842 (O_1842,N_18710,N_18764);
and UO_1843 (O_1843,N_15831,N_17263);
and UO_1844 (O_1844,N_18003,N_16156);
nor UO_1845 (O_1845,N_17786,N_17120);
and UO_1846 (O_1846,N_17837,N_16116);
nand UO_1847 (O_1847,N_18063,N_15755);
or UO_1848 (O_1848,N_19248,N_19927);
nor UO_1849 (O_1849,N_19667,N_15636);
nor UO_1850 (O_1850,N_15372,N_16744);
nor UO_1851 (O_1851,N_18487,N_18144);
or UO_1852 (O_1852,N_19067,N_19259);
and UO_1853 (O_1853,N_17562,N_18355);
nand UO_1854 (O_1854,N_16614,N_19869);
nand UO_1855 (O_1855,N_17776,N_19358);
or UO_1856 (O_1856,N_18687,N_19524);
nor UO_1857 (O_1857,N_19782,N_19309);
and UO_1858 (O_1858,N_17347,N_15400);
nor UO_1859 (O_1859,N_16888,N_19925);
nor UO_1860 (O_1860,N_19705,N_17584);
nor UO_1861 (O_1861,N_18317,N_16647);
xor UO_1862 (O_1862,N_15336,N_15579);
and UO_1863 (O_1863,N_16048,N_18502);
nor UO_1864 (O_1864,N_16968,N_16185);
nor UO_1865 (O_1865,N_17558,N_17577);
nand UO_1866 (O_1866,N_16362,N_18685);
or UO_1867 (O_1867,N_19395,N_16066);
nor UO_1868 (O_1868,N_18326,N_19989);
nor UO_1869 (O_1869,N_17674,N_17428);
and UO_1870 (O_1870,N_15761,N_16152);
or UO_1871 (O_1871,N_18194,N_15263);
nor UO_1872 (O_1872,N_19470,N_18740);
xor UO_1873 (O_1873,N_18129,N_17549);
and UO_1874 (O_1874,N_17255,N_15151);
xnor UO_1875 (O_1875,N_17102,N_19032);
nand UO_1876 (O_1876,N_19146,N_16041);
or UO_1877 (O_1877,N_15771,N_17402);
nand UO_1878 (O_1878,N_19094,N_15971);
nor UO_1879 (O_1879,N_17458,N_16972);
nand UO_1880 (O_1880,N_15292,N_15811);
nand UO_1881 (O_1881,N_18774,N_19714);
xor UO_1882 (O_1882,N_17332,N_16987);
xor UO_1883 (O_1883,N_16999,N_19113);
nor UO_1884 (O_1884,N_15767,N_15696);
and UO_1885 (O_1885,N_16561,N_17835);
nand UO_1886 (O_1886,N_18936,N_15722);
and UO_1887 (O_1887,N_17411,N_16359);
nor UO_1888 (O_1888,N_19845,N_15252);
or UO_1889 (O_1889,N_16265,N_18995);
and UO_1890 (O_1890,N_18040,N_16401);
nand UO_1891 (O_1891,N_15113,N_19915);
nand UO_1892 (O_1892,N_19552,N_16604);
nand UO_1893 (O_1893,N_17203,N_18977);
and UO_1894 (O_1894,N_15993,N_16701);
and UO_1895 (O_1895,N_18401,N_17622);
nor UO_1896 (O_1896,N_18506,N_16631);
and UO_1897 (O_1897,N_16269,N_16467);
and UO_1898 (O_1898,N_17924,N_19163);
nor UO_1899 (O_1899,N_15602,N_15077);
and UO_1900 (O_1900,N_19158,N_18174);
nor UO_1901 (O_1901,N_16246,N_19509);
nand UO_1902 (O_1902,N_17383,N_17404);
xor UO_1903 (O_1903,N_17986,N_15710);
nor UO_1904 (O_1904,N_18600,N_15956);
nand UO_1905 (O_1905,N_15414,N_15436);
and UO_1906 (O_1906,N_19048,N_15240);
and UO_1907 (O_1907,N_19681,N_17475);
and UO_1908 (O_1908,N_19768,N_18493);
and UO_1909 (O_1909,N_18720,N_19539);
and UO_1910 (O_1910,N_18011,N_17369);
nand UO_1911 (O_1911,N_18989,N_18807);
or UO_1912 (O_1912,N_15128,N_16453);
nand UO_1913 (O_1913,N_18256,N_17872);
nor UO_1914 (O_1914,N_15329,N_17554);
nor UO_1915 (O_1915,N_17380,N_18575);
nand UO_1916 (O_1916,N_18439,N_19192);
or UO_1917 (O_1917,N_17126,N_19000);
or UO_1918 (O_1918,N_19016,N_18672);
or UO_1919 (O_1919,N_19853,N_17635);
and UO_1920 (O_1920,N_19418,N_18335);
nand UO_1921 (O_1921,N_16724,N_18711);
nor UO_1922 (O_1922,N_18806,N_16238);
and UO_1923 (O_1923,N_17725,N_17040);
or UO_1924 (O_1924,N_15933,N_19279);
nand UO_1925 (O_1925,N_18910,N_15901);
and UO_1926 (O_1926,N_19006,N_15580);
and UO_1927 (O_1927,N_16464,N_19491);
xnor UO_1928 (O_1928,N_17080,N_19943);
nor UO_1929 (O_1929,N_18309,N_16673);
nand UO_1930 (O_1930,N_18990,N_18327);
or UO_1931 (O_1931,N_18112,N_16495);
xnor UO_1932 (O_1932,N_16680,N_16826);
or UO_1933 (O_1933,N_17653,N_15477);
and UO_1934 (O_1934,N_18045,N_18887);
nand UO_1935 (O_1935,N_15631,N_19527);
or UO_1936 (O_1936,N_15836,N_18224);
and UO_1937 (O_1937,N_15225,N_16113);
nand UO_1938 (O_1938,N_18428,N_16704);
nand UO_1939 (O_1939,N_18412,N_15399);
xor UO_1940 (O_1940,N_18893,N_15508);
nor UO_1941 (O_1941,N_19042,N_15212);
nor UO_1942 (O_1942,N_19868,N_19061);
nor UO_1943 (O_1943,N_19598,N_18598);
nand UO_1944 (O_1944,N_19178,N_15607);
nand UO_1945 (O_1945,N_18755,N_15394);
or UO_1946 (O_1946,N_16140,N_19820);
nand UO_1947 (O_1947,N_16891,N_15342);
nand UO_1948 (O_1948,N_19666,N_18680);
and UO_1949 (O_1949,N_19469,N_15652);
xor UO_1950 (O_1950,N_15100,N_16167);
and UO_1951 (O_1951,N_17053,N_17962);
xor UO_1952 (O_1952,N_15639,N_16216);
and UO_1953 (O_1953,N_19599,N_17094);
nand UO_1954 (O_1954,N_19806,N_18564);
and UO_1955 (O_1955,N_15360,N_15899);
nor UO_1956 (O_1956,N_15332,N_18489);
nand UO_1957 (O_1957,N_16558,N_19948);
and UO_1958 (O_1958,N_19372,N_19391);
nand UO_1959 (O_1959,N_19272,N_15299);
or UO_1960 (O_1960,N_17316,N_17984);
or UO_1961 (O_1961,N_18800,N_15075);
or UO_1962 (O_1962,N_15520,N_15492);
xor UO_1963 (O_1963,N_15713,N_18247);
or UO_1964 (O_1964,N_17002,N_17856);
and UO_1965 (O_1965,N_19508,N_17172);
or UO_1966 (O_1966,N_17377,N_16373);
nand UO_1967 (O_1967,N_19786,N_19673);
nor UO_1968 (O_1968,N_17012,N_18574);
and UO_1969 (O_1969,N_19045,N_15040);
nand UO_1970 (O_1970,N_16084,N_17384);
nor UO_1971 (O_1971,N_15363,N_18944);
xnor UO_1972 (O_1972,N_17433,N_19972);
or UO_1973 (O_1973,N_17018,N_17996);
or UO_1974 (O_1974,N_19054,N_18192);
or UO_1975 (O_1975,N_15951,N_15961);
and UO_1976 (O_1976,N_17861,N_19657);
nor UO_1977 (O_1977,N_15765,N_15770);
nor UO_1978 (O_1978,N_17367,N_15531);
and UO_1979 (O_1979,N_18842,N_16352);
and UO_1980 (O_1980,N_15610,N_19482);
nand UO_1981 (O_1981,N_16768,N_15505);
and UO_1982 (O_1982,N_15166,N_15719);
and UO_1983 (O_1983,N_15312,N_19991);
or UO_1984 (O_1984,N_17497,N_15659);
or UO_1985 (O_1985,N_17662,N_15474);
and UO_1986 (O_1986,N_17889,N_19968);
nand UO_1987 (O_1987,N_17207,N_15711);
and UO_1988 (O_1988,N_19313,N_19725);
nor UO_1989 (O_1989,N_18752,N_15064);
nand UO_1990 (O_1990,N_19702,N_19081);
nor UO_1991 (O_1991,N_16932,N_18534);
or UO_1992 (O_1992,N_18768,N_19520);
and UO_1993 (O_1993,N_16399,N_19732);
xor UO_1994 (O_1994,N_19025,N_16930);
and UO_1995 (O_1995,N_19640,N_17518);
and UO_1996 (O_1996,N_16622,N_18093);
nand UO_1997 (O_1997,N_19080,N_18111);
nand UO_1998 (O_1998,N_17470,N_19477);
nor UO_1999 (O_1999,N_17007,N_16532);
xor UO_2000 (O_2000,N_15071,N_15872);
nand UO_2001 (O_2001,N_18252,N_18061);
nor UO_2002 (O_2002,N_17550,N_17125);
nand UO_2003 (O_2003,N_15016,N_16547);
and UO_2004 (O_2004,N_19544,N_17777);
or UO_2005 (O_2005,N_16912,N_15709);
xnor UO_2006 (O_2006,N_15111,N_15271);
nand UO_2007 (O_2007,N_18862,N_18239);
nor UO_2008 (O_2008,N_19849,N_15203);
and UO_2009 (O_2009,N_16941,N_19850);
or UO_2010 (O_2010,N_19974,N_18300);
nand UO_2011 (O_2011,N_15109,N_17004);
and UO_2012 (O_2012,N_16182,N_17633);
nand UO_2013 (O_2013,N_18952,N_16051);
nor UO_2014 (O_2014,N_17744,N_19803);
nor UO_2015 (O_2015,N_15186,N_16653);
or UO_2016 (O_2016,N_19286,N_19440);
or UO_2017 (O_2017,N_15592,N_17657);
nor UO_2018 (O_2018,N_17355,N_17883);
nor UO_2019 (O_2019,N_18747,N_16365);
and UO_2020 (O_2020,N_17652,N_19118);
or UO_2021 (O_2021,N_18255,N_17230);
nand UO_2022 (O_2022,N_19069,N_18754);
nor UO_2023 (O_2023,N_19457,N_19796);
nor UO_2024 (O_2024,N_16325,N_16676);
xnor UO_2025 (O_2025,N_16652,N_15680);
and UO_2026 (O_2026,N_17174,N_19478);
nand UO_2027 (O_2027,N_18699,N_17649);
and UO_2028 (O_2028,N_15027,N_17076);
nand UO_2029 (O_2029,N_19862,N_17870);
nor UO_2030 (O_2030,N_19295,N_15634);
nor UO_2031 (O_2031,N_16715,N_16297);
and UO_2032 (O_2032,N_19821,N_19464);
nor UO_2033 (O_2033,N_16448,N_17158);
or UO_2034 (O_2034,N_18938,N_16935);
nand UO_2035 (O_2035,N_17089,N_15932);
or UO_2036 (O_2036,N_18556,N_19995);
or UO_2037 (O_2037,N_18411,N_15691);
nor UO_2038 (O_2038,N_17244,N_19745);
or UO_2039 (O_2039,N_19426,N_15984);
nor UO_2040 (O_2040,N_16712,N_19133);
or UO_2041 (O_2041,N_17586,N_15385);
and UO_2042 (O_2042,N_15637,N_17017);
nor UO_2043 (O_2043,N_16834,N_17717);
or UO_2044 (O_2044,N_16848,N_16857);
or UO_2045 (O_2045,N_16075,N_17152);
nand UO_2046 (O_2046,N_16210,N_18694);
xnor UO_2047 (O_2047,N_16738,N_17748);
xnor UO_2048 (O_2048,N_16057,N_15085);
or UO_2049 (O_2049,N_18856,N_19929);
and UO_2050 (O_2050,N_19043,N_15700);
nand UO_2051 (O_2051,N_17361,N_15134);
xor UO_2052 (O_2052,N_18471,N_18877);
or UO_2053 (O_2053,N_17164,N_16242);
nand UO_2054 (O_2054,N_17767,N_19221);
xor UO_2055 (O_2055,N_15608,N_15671);
nor UO_2056 (O_2056,N_16510,N_18707);
or UO_2057 (O_2057,N_19495,N_19462);
or UO_2058 (O_2058,N_19506,N_15509);
nor UO_2059 (O_2059,N_16752,N_17576);
nor UO_2060 (O_2060,N_15590,N_17914);
and UO_2061 (O_2061,N_19415,N_18125);
nand UO_2062 (O_2062,N_19564,N_17893);
or UO_2063 (O_2063,N_17231,N_16612);
nor UO_2064 (O_2064,N_15146,N_15236);
nand UO_2065 (O_2065,N_18746,N_16240);
and UO_2066 (O_2066,N_16842,N_18182);
xor UO_2067 (O_2067,N_17921,N_15594);
nor UO_2068 (O_2068,N_19169,N_19020);
nor UO_2069 (O_2069,N_17340,N_18261);
nor UO_2070 (O_2070,N_15065,N_17659);
nor UO_2071 (O_2071,N_15278,N_19952);
nor UO_2072 (O_2072,N_19442,N_19251);
or UO_2073 (O_2073,N_19690,N_18145);
or UO_2074 (O_2074,N_16062,N_17848);
xnor UO_2075 (O_2075,N_17646,N_18169);
nor UO_2076 (O_2076,N_16723,N_19211);
xnor UO_2077 (O_2077,N_18166,N_19107);
nand UO_2078 (O_2078,N_15522,N_19505);
nand UO_2079 (O_2079,N_16189,N_18176);
or UO_2080 (O_2080,N_16610,N_17476);
or UO_2081 (O_2081,N_16281,N_19319);
nor UO_2082 (O_2082,N_16124,N_18384);
or UO_2083 (O_2083,N_18172,N_19467);
or UO_2084 (O_2084,N_18643,N_16885);
or UO_2085 (O_2085,N_16840,N_15878);
and UO_2086 (O_2086,N_16218,N_17176);
or UO_2087 (O_2087,N_17802,N_16839);
or UO_2088 (O_2088,N_16419,N_16061);
or UO_2089 (O_2089,N_16851,N_16832);
or UO_2090 (O_2090,N_17640,N_16443);
and UO_2091 (O_2091,N_17037,N_16251);
and UO_2092 (O_2092,N_19658,N_19108);
nand UO_2093 (O_2093,N_15156,N_18933);
and UO_2094 (O_2094,N_19431,N_19716);
nor UO_2095 (O_2095,N_17691,N_18303);
or UO_2096 (O_2096,N_15848,N_19217);
or UO_2097 (O_2097,N_17873,N_18260);
and UO_2098 (O_2098,N_19531,N_16268);
nand UO_2099 (O_2099,N_16992,N_17982);
nor UO_2100 (O_2100,N_18420,N_19407);
nand UO_2101 (O_2101,N_16338,N_18665);
nor UO_2102 (O_2102,N_17862,N_17135);
nor UO_2103 (O_2103,N_17395,N_18949);
and UO_2104 (O_2104,N_18580,N_19600);
and UO_2105 (O_2105,N_19824,N_17331);
nor UO_2106 (O_2106,N_15032,N_16280);
or UO_2107 (O_2107,N_15785,N_16697);
nand UO_2108 (O_2108,N_17113,N_15314);
nand UO_2109 (O_2109,N_17293,N_18639);
nand UO_2110 (O_2110,N_15265,N_16695);
nor UO_2111 (O_2111,N_17858,N_19466);
or UO_2112 (O_2112,N_18323,N_15769);
or UO_2113 (O_2113,N_19105,N_19928);
nor UO_2114 (O_2114,N_15168,N_19336);
and UO_2115 (O_2115,N_15157,N_17461);
or UO_2116 (O_2116,N_18180,N_19138);
nor UO_2117 (O_2117,N_19147,N_17681);
nand UO_2118 (O_2118,N_16031,N_15079);
nor UO_2119 (O_2119,N_19689,N_16665);
nor UO_2120 (O_2120,N_18765,N_19128);
and UO_2121 (O_2121,N_19397,N_19569);
nor UO_2122 (O_2122,N_16254,N_17348);
or UO_2123 (O_2123,N_19844,N_18796);
and UO_2124 (O_2124,N_18907,N_19620);
or UO_2125 (O_2125,N_18762,N_17515);
nor UO_2126 (O_2126,N_17457,N_16908);
nand UO_2127 (O_2127,N_16447,N_19238);
nand UO_2128 (O_2128,N_15046,N_16132);
nand UO_2129 (O_2129,N_18077,N_15228);
nand UO_2130 (O_2130,N_18738,N_18955);
and UO_2131 (O_2131,N_15953,N_18292);
or UO_2132 (O_2132,N_18689,N_15975);
and UO_2133 (O_2133,N_15601,N_16613);
nand UO_2134 (O_2134,N_16993,N_16000);
nand UO_2135 (O_2135,N_17679,N_19930);
nand UO_2136 (O_2136,N_18191,N_15082);
and UO_2137 (O_2137,N_16275,N_19066);
or UO_2138 (O_2138,N_17329,N_16663);
and UO_2139 (O_2139,N_17264,N_16534);
nand UO_2140 (O_2140,N_18410,N_19815);
and UO_2141 (O_2141,N_17950,N_16763);
nand UO_2142 (O_2142,N_17346,N_15787);
nor UO_2143 (O_2143,N_18617,N_15074);
xnor UO_2144 (O_2144,N_18121,N_18507);
and UO_2145 (O_2145,N_19071,N_17190);
nor UO_2146 (O_2146,N_15996,N_16520);
and UO_2147 (O_2147,N_17041,N_18698);
or UO_2148 (O_2148,N_15437,N_16777);
and UO_2149 (O_2149,N_17392,N_15222);
nand UO_2150 (O_2150,N_19629,N_18294);
nand UO_2151 (O_2151,N_19739,N_15441);
or UO_2152 (O_2152,N_18139,N_16346);
nor UO_2153 (O_2153,N_18828,N_16449);
and UO_2154 (O_2154,N_16333,N_15539);
nor UO_2155 (O_2155,N_15690,N_15837);
or UO_2156 (O_2156,N_15620,N_16123);
or UO_2157 (O_2157,N_15480,N_18452);
or UO_2158 (O_2158,N_18978,N_16193);
or UO_2159 (O_2159,N_17474,N_15501);
nand UO_2160 (O_2160,N_19304,N_19363);
nand UO_2161 (O_2161,N_18032,N_17669);
and UO_2162 (O_2162,N_17546,N_18161);
xor UO_2163 (O_2163,N_16397,N_19379);
nand UO_2164 (O_2164,N_17429,N_17273);
and UO_2165 (O_2165,N_15729,N_19761);
and UO_2166 (O_2166,N_19997,N_19865);
nand UO_2167 (O_2167,N_19525,N_17959);
or UO_2168 (O_2168,N_15380,N_15472);
nor UO_2169 (O_2169,N_15245,N_19096);
and UO_2170 (O_2170,N_19805,N_16332);
nand UO_2171 (O_2171,N_16199,N_15564);
or UO_2172 (O_2172,N_17501,N_15555);
nand UO_2173 (O_2173,N_18333,N_19450);
and UO_2174 (O_2174,N_18813,N_16735);
nand UO_2175 (O_2175,N_16624,N_17281);
xor UO_2176 (O_2176,N_15487,N_15189);
nand UO_2177 (O_2177,N_19587,N_19842);
nand UO_2178 (O_2178,N_15763,N_18353);
nor UO_2179 (O_2179,N_15999,N_17284);
or UO_2180 (O_2180,N_17825,N_15412);
nor UO_2181 (O_2181,N_18630,N_19819);
nand UO_2182 (O_2182,N_19161,N_17023);
nand UO_2183 (O_2183,N_16973,N_17477);
xnor UO_2184 (O_2184,N_19625,N_16433);
nand UO_2185 (O_2185,N_17534,N_17365);
and UO_2186 (O_2186,N_17388,N_19064);
nand UO_2187 (O_2187,N_16505,N_16921);
or UO_2188 (O_2188,N_17350,N_19405);
nor UO_2189 (O_2189,N_18306,N_17489);
nand UO_2190 (O_2190,N_15424,N_19281);
nor UO_2191 (O_2191,N_19619,N_15323);
nor UO_2192 (O_2192,N_15644,N_16348);
and UO_2193 (O_2193,N_17917,N_17181);
nand UO_2194 (O_2194,N_15308,N_16150);
nand UO_2195 (O_2195,N_18548,N_16836);
or UO_2196 (O_2196,N_15368,N_15759);
nand UO_2197 (O_2197,N_19618,N_18392);
or UO_2198 (O_2198,N_15382,N_15432);
or UO_2199 (O_2199,N_19605,N_18924);
xnor UO_2200 (O_2200,N_18742,N_15635);
nand UO_2201 (O_2201,N_18130,N_16046);
nand UO_2202 (O_2202,N_17892,N_15406);
nor UO_2203 (O_2203,N_18141,N_16537);
nor UO_2204 (O_2204,N_18123,N_17533);
nand UO_2205 (O_2205,N_18612,N_15972);
nor UO_2206 (O_2206,N_19277,N_17415);
or UO_2207 (O_2207,N_18849,N_17219);
nor UO_2208 (O_2208,N_16054,N_18683);
nor UO_2209 (O_2209,N_16217,N_18448);
and UO_2210 (O_2210,N_16684,N_16019);
and UO_2211 (O_2211,N_17784,N_17494);
or UO_2212 (O_2212,N_18187,N_16320);
xor UO_2213 (O_2213,N_18240,N_19789);
or UO_2214 (O_2214,N_19448,N_15488);
and UO_2215 (O_2215,N_19116,N_18544);
nor UO_2216 (O_2216,N_16589,N_16762);
and UO_2217 (O_2217,N_18703,N_19377);
and UO_2218 (O_2218,N_19171,N_18088);
or UO_2219 (O_2219,N_16354,N_18721);
nand UO_2220 (O_2220,N_17905,N_15842);
nor UO_2221 (O_2221,N_17719,N_16964);
and UO_2222 (O_2222,N_15507,N_15891);
nand UO_2223 (O_2223,N_16485,N_19817);
or UO_2224 (O_2224,N_18560,N_17980);
nand UO_2225 (O_2225,N_16740,N_17426);
and UO_2226 (O_2226,N_18898,N_16995);
and UO_2227 (O_2227,N_19367,N_15537);
xnor UO_2228 (O_2228,N_19560,N_17821);
or UO_2229 (O_2229,N_18956,N_15942);
xor UO_2230 (O_2230,N_18858,N_15627);
xnor UO_2231 (O_2231,N_19463,N_18059);
nor UO_2232 (O_2232,N_16633,N_19433);
nand UO_2233 (O_2233,N_16940,N_15485);
nor UO_2234 (O_2234,N_16504,N_16984);
nand UO_2235 (O_2235,N_15297,N_17295);
and UO_2236 (O_2236,N_17467,N_16377);
nand UO_2237 (O_2237,N_15573,N_15582);
nand UO_2238 (O_2238,N_19663,N_16607);
nand UO_2239 (O_2239,N_19099,N_16967);
or UO_2240 (O_2240,N_15494,N_16796);
nor UO_2241 (O_2241,N_17243,N_16033);
or UO_2242 (O_2242,N_19638,N_18520);
or UO_2243 (O_2243,N_18557,N_16926);
nor UO_2244 (O_2244,N_18923,N_15911);
and UO_2245 (O_2245,N_17015,N_16484);
or UO_2246 (O_2246,N_15179,N_16296);
and UO_2247 (O_2247,N_17811,N_18931);
xnor UO_2248 (O_2248,N_17716,N_16585);
xor UO_2249 (O_2249,N_19184,N_15089);
nand UO_2250 (O_2250,N_15072,N_16951);
and UO_2251 (O_2251,N_17937,N_16314);
and UO_2252 (O_2252,N_15267,N_15120);
or UO_2253 (O_2253,N_17416,N_18102);
or UO_2254 (O_2254,N_18713,N_19776);
nand UO_2255 (O_2255,N_18581,N_19708);
nand UO_2256 (O_2256,N_15930,N_18568);
nand UO_2257 (O_2257,N_16808,N_19292);
or UO_2258 (O_2258,N_18883,N_15339);
nor UO_2259 (O_2259,N_16405,N_15904);
and UO_2260 (O_2260,N_17279,N_17947);
or UO_2261 (O_2261,N_16667,N_15649);
or UO_2262 (O_2262,N_18551,N_18140);
or UO_2263 (O_2263,N_17751,N_17177);
nand UO_2264 (O_2264,N_16306,N_16587);
or UO_2265 (O_2265,N_19049,N_16303);
or UO_2266 (O_2266,N_16688,N_19341);
nand UO_2267 (O_2267,N_18533,N_15277);
nand UO_2268 (O_2268,N_19635,N_18821);
nor UO_2269 (O_2269,N_15045,N_16574);
xor UO_2270 (O_2270,N_18904,N_19494);
nand UO_2271 (O_2271,N_15788,N_17579);
and UO_2272 (O_2272,N_17127,N_15207);
nor UO_2273 (O_2273,N_15175,N_15561);
nor UO_2274 (O_2274,N_16437,N_17468);
or UO_2275 (O_2275,N_19753,N_17891);
nand UO_2276 (O_2276,N_19933,N_17345);
nand UO_2277 (O_2277,N_15736,N_15572);
or UO_2278 (O_2278,N_15632,N_19214);
or UO_2279 (O_2279,N_17842,N_16582);
nand UO_2280 (O_2280,N_17666,N_17356);
xnor UO_2281 (O_2281,N_15495,N_16439);
and UO_2282 (O_2282,N_18447,N_17097);
nand UO_2283 (O_2283,N_18037,N_17421);
and UO_2284 (O_2284,N_16056,N_17676);
xor UO_2285 (O_2285,N_18496,N_16100);
or UO_2286 (O_2286,N_18810,N_16197);
or UO_2287 (O_2287,N_18086,N_16004);
xor UO_2288 (O_2288,N_18074,N_17029);
nand UO_2289 (O_2289,N_19507,N_18724);
and UO_2290 (O_2290,N_19851,N_16746);
xor UO_2291 (O_2291,N_17278,N_15957);
nor UO_2292 (O_2292,N_19018,N_15253);
and UO_2293 (O_2293,N_19413,N_18079);
and UO_2294 (O_2294,N_18753,N_16522);
nor UO_2295 (O_2295,N_19558,N_17503);
nor UO_2296 (O_2296,N_15439,N_15989);
and UO_2297 (O_2297,N_15803,N_15734);
nor UO_2298 (O_2298,N_19723,N_19068);
nand UO_2299 (O_2299,N_15286,N_18198);
nor UO_2300 (O_2300,N_15125,N_16221);
nor UO_2301 (O_2301,N_16736,N_19033);
and UO_2302 (O_2302,N_16691,N_18820);
nand UO_2303 (O_2303,N_17614,N_19244);
nor UO_2304 (O_2304,N_19437,N_18739);
or UO_2305 (O_2305,N_17715,N_16843);
nor UO_2306 (O_2306,N_17876,N_19606);
or UO_2307 (O_2307,N_16517,N_17131);
nand UO_2308 (O_2308,N_16035,N_17057);
and UO_2309 (O_2309,N_17218,N_15383);
or UO_2310 (O_2310,N_18690,N_18184);
or UO_2311 (O_2311,N_18109,N_18781);
nor UO_2312 (O_2312,N_16831,N_18371);
nor UO_2313 (O_2313,N_16837,N_19088);
and UO_2314 (O_2314,N_18357,N_16068);
and UO_2315 (O_2315,N_16454,N_17302);
nand UO_2316 (O_2316,N_15651,N_19301);
nor UO_2317 (O_2317,N_16643,N_16175);
or UO_2318 (O_2318,N_19144,N_19137);
nand UO_2319 (O_2319,N_19421,N_15873);
nor UO_2320 (O_2320,N_16583,N_17443);
or UO_2321 (O_2321,N_16291,N_16896);
and UO_2322 (O_2322,N_18798,N_18875);
and UO_2323 (O_2323,N_18651,N_16469);
or UO_2324 (O_2324,N_17604,N_19228);
nor UO_2325 (O_2325,N_16780,N_19165);
or UO_2326 (O_2326,N_19682,N_15603);
nor UO_2327 (O_2327,N_19655,N_18926);
and UO_2328 (O_2328,N_19919,N_19902);
xnor UO_2329 (O_2329,N_19647,N_18782);
and UO_2330 (O_2330,N_17537,N_19022);
nor UO_2331 (O_2331,N_16703,N_16779);
nor UO_2332 (O_2332,N_15347,N_16179);
and UO_2333 (O_2333,N_17146,N_18450);
nor UO_2334 (O_2334,N_16675,N_15791);
and UO_2335 (O_2335,N_17514,N_15754);
xor UO_2336 (O_2336,N_18846,N_19909);
and UO_2337 (O_2337,N_19734,N_15506);
or UO_2338 (O_2338,N_19023,N_17629);
nor UO_2339 (O_2339,N_16869,N_18330);
and UO_2340 (O_2340,N_18704,N_19879);
nand UO_2341 (O_2341,N_17438,N_17700);
or UO_2342 (O_2342,N_19937,N_16716);
nor UO_2343 (O_2343,N_18546,N_19212);
nor UO_2344 (O_2344,N_16136,N_18271);
xnor UO_2345 (O_2345,N_19434,N_16355);
nand UO_2346 (O_2346,N_18263,N_18380);
nand UO_2347 (O_2347,N_17083,N_15144);
or UO_2348 (O_2348,N_16562,N_19091);
nand UO_2349 (O_2349,N_16177,N_17419);
xor UO_2350 (O_2350,N_16262,N_18073);
xor UO_2351 (O_2351,N_16427,N_18289);
nor UO_2352 (O_2352,N_19829,N_16511);
nor UO_2353 (O_2353,N_18693,N_18664);
and UO_2354 (O_2354,N_17030,N_18019);
and UO_2355 (O_2355,N_18524,N_19189);
nand UO_2356 (O_2356,N_15780,N_18367);
nand UO_2357 (O_2357,N_15254,N_15781);
or UO_2358 (O_2358,N_19121,N_18106);
or UO_2359 (O_2359,N_16751,N_17410);
nor UO_2360 (O_2360,N_17760,N_19541);
or UO_2361 (O_2361,N_17702,N_15343);
or UO_2362 (O_2362,N_15481,N_17085);
nand UO_2363 (O_2363,N_16850,N_19396);
and UO_2364 (O_2364,N_18538,N_16818);
nor UO_2365 (O_2365,N_18230,N_18154);
or UO_2366 (O_2366,N_16082,N_15575);
xor UO_2367 (O_2367,N_15258,N_18099);
xor UO_2368 (O_2368,N_18352,N_18646);
nand UO_2369 (O_2369,N_17840,N_16641);
nand UO_2370 (O_2370,N_19008,N_16277);
and UO_2371 (O_2371,N_15693,N_18585);
nor UO_2372 (O_2372,N_17871,N_19129);
nor UO_2373 (O_2373,N_18599,N_18120);
xnor UO_2374 (O_2374,N_16270,N_19665);
or UO_2375 (O_2375,N_18068,N_15458);
xor UO_2376 (O_2376,N_19136,N_16559);
nor UO_2377 (O_2377,N_18595,N_15723);
and UO_2378 (O_2378,N_18613,N_15726);
nor UO_2379 (O_2379,N_18320,N_15692);
and UO_2380 (O_2380,N_15869,N_19349);
or UO_2381 (O_2381,N_17829,N_17391);
or UO_2382 (O_2382,N_15558,N_19271);
and UO_2383 (O_2383,N_18343,N_15059);
nand UO_2384 (O_2384,N_19414,N_18902);
xor UO_2385 (O_2385,N_17427,N_17728);
nand UO_2386 (O_2386,N_15926,N_19265);
nor UO_2387 (O_2387,N_19368,N_17897);
xnor UO_2388 (O_2388,N_18360,N_19592);
nand UO_2389 (O_2389,N_16459,N_16664);
and UO_2390 (O_2390,N_18985,N_19582);
nand UO_2391 (O_2391,N_15274,N_18179);
or UO_2392 (O_2392,N_16347,N_15915);
or UO_2393 (O_2393,N_15135,N_19316);
xor UO_2394 (O_2394,N_17087,N_17689);
nor UO_2395 (O_2395,N_18971,N_15824);
nor UO_2396 (O_2396,N_16411,N_19823);
nor UO_2397 (O_2397,N_16619,N_16492);
and UO_2398 (O_2398,N_16795,N_15141);
nand UO_2399 (O_2399,N_15917,N_17200);
nor UO_2400 (O_2400,N_17070,N_16110);
or UO_2401 (O_2401,N_16300,N_19445);
or UO_2402 (O_2402,N_19412,N_17707);
nor UO_2403 (O_2403,N_19390,N_17743);
nor UO_2404 (O_2404,N_17606,N_19290);
or UO_2405 (O_2405,N_17739,N_19680);
and UO_2406 (O_2406,N_15390,N_19735);
and UO_2407 (O_2407,N_19967,N_15504);
xor UO_2408 (O_2408,N_19864,N_16764);
or UO_2409 (O_2409,N_15092,N_18188);
and UO_2410 (O_2410,N_18805,N_17686);
or UO_2411 (O_2411,N_15122,N_15854);
nand UO_2412 (O_2412,N_19751,N_17191);
and UO_2413 (O_2413,N_16758,N_16600);
nor UO_2414 (O_2414,N_19039,N_16192);
or UO_2415 (O_2415,N_15457,N_15325);
nand UO_2416 (O_2416,N_18314,N_16466);
nand UO_2417 (O_2417,N_19872,N_15359);
and UO_2418 (O_2418,N_15566,N_19935);
or UO_2419 (O_2419,N_19812,N_17602);
xor UO_2420 (O_2420,N_19669,N_16541);
nand UO_2421 (O_2421,N_15525,N_18222);
nor UO_2422 (O_2422,N_19030,N_19672);
and UO_2423 (O_2423,N_18999,N_18514);
and UO_2424 (O_2424,N_15802,N_18519);
and UO_2425 (O_2425,N_16076,N_16261);
nand UO_2426 (O_2426,N_18236,N_17465);
or UO_2427 (O_2427,N_16952,N_19923);
nor UO_2428 (O_2428,N_19253,N_17710);
nor UO_2429 (O_2429,N_19266,N_16337);
or UO_2430 (O_2430,N_18823,N_18928);
nand UO_2431 (O_2431,N_16026,N_15192);
xnor UO_2432 (O_2432,N_18779,N_16153);
and UO_2433 (O_2433,N_15055,N_18344);
xnor UO_2434 (O_2434,N_19343,N_18469);
nand UO_2435 (O_2435,N_17141,N_18266);
and UO_2436 (O_2436,N_17630,N_19612);
and UO_2437 (O_2437,N_15954,N_15893);
or UO_2438 (O_2438,N_19179,N_15866);
nand UO_2439 (O_2439,N_16977,N_17266);
nand UO_2440 (O_2440,N_15544,N_17990);
nand UO_2441 (O_2441,N_16519,N_15945);
and UO_2442 (O_2442,N_17631,N_16962);
and UO_2443 (O_2443,N_17768,N_17526);
and UO_2444 (O_2444,N_15646,N_19345);
nor UO_2445 (O_2445,N_18590,N_19298);
nand UO_2446 (O_2446,N_16953,N_17555);
and UO_2447 (O_2447,N_16258,N_16927);
nand UO_2448 (O_2448,N_15569,N_18456);
or UO_2449 (O_2449,N_18347,N_16223);
or UO_2450 (O_2450,N_15969,N_15029);
and UO_2451 (O_2451,N_15313,N_17561);
nand UO_2452 (O_2452,N_17221,N_16072);
or UO_2453 (O_2453,N_15884,N_19748);
nor UO_2454 (O_2454,N_16025,N_17086);
nor UO_2455 (O_2455,N_17958,N_16257);
xor UO_2456 (O_2456,N_15063,N_18430);
nand UO_2457 (O_2457,N_19353,N_19530);
and UO_2458 (O_2458,N_15875,N_19382);
and UO_2459 (O_2459,N_19903,N_16669);
and UO_2460 (O_2460,N_15266,N_15223);
and UO_2461 (O_2461,N_16284,N_18623);
and UO_2462 (O_2462,N_15887,N_16566);
and UO_2463 (O_2463,N_19321,N_15410);
nor UO_2464 (O_2464,N_17289,N_17071);
nand UO_2465 (O_2465,N_15574,N_18554);
nor UO_2466 (O_2466,N_15140,N_16904);
and UO_2467 (O_2467,N_17042,N_16787);
nor UO_2468 (O_2468,N_19131,N_19959);
nand UO_2469 (O_2469,N_17050,N_19460);
and UO_2470 (O_2470,N_19956,N_18322);
xnor UO_2471 (O_2471,N_19840,N_17290);
or UO_2472 (O_2472,N_18305,N_16863);
and UO_2473 (O_2473,N_19143,N_17867);
nor UO_2474 (O_2474,N_18728,N_16945);
nor UO_2475 (O_2475,N_17504,N_16108);
nor UO_2476 (O_2476,N_18586,N_19227);
xor UO_2477 (O_2477,N_16974,N_15750);
or UO_2478 (O_2478,N_19900,N_17303);
nand UO_2479 (O_2479,N_19308,N_18562);
nand UO_2480 (O_2480,N_19814,N_16602);
nand UO_2481 (O_2481,N_17298,N_17253);
or UO_2482 (O_2482,N_17075,N_17807);
or UO_2483 (O_2483,N_19770,N_18794);
nor UO_2484 (O_2484,N_17209,N_17285);
xnor UO_2485 (O_2485,N_15020,N_15459);
and UO_2486 (O_2486,N_19487,N_16980);
or UO_2487 (O_2487,N_15220,N_17975);
xnor UO_2488 (O_2488,N_19317,N_18315);
nand UO_2489 (O_2489,N_15350,N_19977);
and UO_2490 (O_2490,N_19779,N_18974);
or UO_2491 (O_2491,N_17547,N_16956);
nand UO_2492 (O_2492,N_15705,N_19453);
nor UO_2493 (O_2493,N_15908,N_19549);
and UO_2494 (O_2494,N_17407,N_19078);
nor UO_2495 (O_2495,N_19338,N_15095);
and UO_2496 (O_2496,N_18618,N_18954);
nor UO_2497 (O_2497,N_17321,N_16420);
or UO_2498 (O_2498,N_19759,N_17170);
or UO_2499 (O_2499,N_16630,N_16106);
endmodule